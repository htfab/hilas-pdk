VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_li2m2
  CLASS BLOCK ;
  FOREIGN sky130_hilas_li2m2 ;
  ORIGIN 0.140 0.150 ;
  SIZE 0.340 BY 0.330 ;
  OBS
      LAYER li1 ;
        RECT -0.130 0.100 0.190 0.140 ;
        RECT -0.130 -0.090 0.200 0.100 ;
        RECT -0.130 -0.120 0.190 -0.090 ;
      LAYER mcon ;
        RECT -0.070 -0.080 0.100 0.090 ;
      LAYER met1 ;
        RECT -0.140 -0.150 0.180 0.170 ;
      LAYER via ;
        RECT -0.110 -0.120 0.150 0.140 ;
      LAYER met2 ;
        RECT -0.140 -0.150 0.170 0.180 ;
  END
END sky130_hilas_li2m2
END LIBRARY

