VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_TgateSingle01Part2
  CLASS BLOCK ;
  FOREIGN /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_TgateSingle01Part2 ;
  ORIGIN 0.670 1.810 ;
  SIZE 1.630 BY 1.430 ;
  OBS
      LAYER nwell ;
        RECT -0.670 -1.810 0.960 -0.970 ;
      LAYER li1 ;
        RECT -0.270 -1.670 0.960 -0.700 ;
      LAYER met1 ;
        RECT -0.280 -1.700 0.950 -0.470 ;
      LAYER met2 ;
        RECT -0.670 -1.710 0.960 -0.500 ;
  END
END /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_TgateSingle01Part2
END LIBRARY

