* NGSPICE file created from /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_pFETLargePart1.ext - technology: sky130A

.subckt sky130_hilas_pFETmed a_440_n8# w_294_n44# $SUB a_330_n8#
X0 a_440_n8# a_388_n34# a_330_n8# w_294_n44# sky130_fd_pr__pfet_01v8 w=2.51e+06u l=260000u
.ends


* Top level circuit /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_pFETLargePart1

Xsky130_hilas_pFETmed_0 sky130_hilas_pFETmed_1/a_330_n8# sky130_hilas_pFETmed_4/w_294_n44#
+ $SUB sky130_hilas_pFETmed_4/a_440_n8# sky130_hilas_pFETmed
Xsky130_hilas_pFETmed_2 sky130_hilas_pFETmed_3/a_330_n8# sky130_hilas_pFETmed_4/w_294_n44#
+ $SUB sky130_hilas_pFETmed_2/a_330_n8# sky130_hilas_pFETmed
Xsky130_hilas_pFETmed_1 sky130_hilas_pFETmed_2/a_330_n8# sky130_hilas_pFETmed_4/w_294_n44#
+ $SUB sky130_hilas_pFETmed_1/a_330_n8# sky130_hilas_pFETmed
Xsky130_hilas_pFETmed_3 sky130_hilas_pFETmed_3/a_440_n8# sky130_hilas_pFETmed_4/w_294_n44#
+ $SUB sky130_hilas_pFETmed_3/a_330_n8# sky130_hilas_pFETmed
Xsky130_hilas_pFETmed_4 sky130_hilas_pFETmed_4/a_440_n8# sky130_hilas_pFETmed_4/w_294_n44#
+ $SUB sky130_hilas_pFETmed_4/a_330_n8# sky130_hilas_pFETmed
.end

