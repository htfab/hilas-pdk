* NGSPICE file created from /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_CapModule03.ext - technology: sky130A


* Top level circuit /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_CapModule03

X0 c1_n664_n410# m3_n784_n490# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=3.22e+06u
.end

