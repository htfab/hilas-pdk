magic
tech sky130A
timestamp 1632494644
<< error_s >>
rect -1025 555 -1009 569
rect -984 555 -965 569
rect -826 513 -805 530
rect -805 342 -784 359
rect -817 319 -800 322
rect -817 308 -803 319
rect -997 279 -966 282
rect -957 279 -949 282
rect -1025 264 -1009 278
rect -997 274 -944 279
rect -997 269 -941 274
rect -997 268 -961 269
rect -997 265 -984 268
rect -982 265 -961 268
rect -997 264 -994 265
rect -982 257 -969 264
rect -966 262 -961 265
rect -954 266 -941 269
rect -954 265 -944 266
rect -954 264 -949 265
rect -954 262 -944 264
rect -966 257 -944 262
rect -973 244 -970 254
rect -957 252 -944 257
rect -957 249 -949 252
rect -817 206 -802 210
rect -826 193 -802 206
rect -826 189 -805 193
rect -805 17 -784 34
rect -1025 -42 -1009 -28
rect -984 -42 -965 -28
<< nwell >>
rect -1101 561 -805 562
rect -1101 546 -1060 561
rect -532 552 -494 562
rect -129 548 -89 562
rect -1101 545 -1042 546
rect -1101 369 -1060 545
rect -1112 327 -1060 369
rect -1112 307 -1061 327
rect -1112 254 -1060 307
rect -1101 -42 -1060 254
<< poly >>
rect 209 516 229 589
rect 209 -61 229 -18
<< locali >>
rect -1115 -25 -1097 67
<< metal1 >>
rect -1025 555 -1009 562
rect -984 555 -965 562
rect -944 555 -928 562
rect -532 552 -494 562
rect -129 534 -89 562
rect 131 516 154 589
rect 257 516 280 589
rect -782 430 -761 504
rect -1112 254 -1091 369
rect -784 93 -768 243
rect 257 127 280 132
rect 253 126 281 127
rect 253 124 283 126
rect 253 97 254 124
rect 281 97 283 124
rect 253 94 283 97
rect -532 -43 -494 -33
rect 131 -61 154 -18
rect 257 -61 280 -18
<< via1 >>
rect 254 97 281 124
<< metal2 >>
rect -1116 515 -1043 533
rect -758 512 7 531
rect -758 510 24 512
rect -14 491 24 510
rect -65 490 -51 491
rect -1112 427 -1097 469
rect -65 457 -50 490
rect -65 437 56 457
rect -1112 418 -785 427
rect 170 426 296 442
rect -1112 412 -769 418
rect -799 402 -769 412
rect -1114 352 -1082 379
rect -54 371 66 381
rect -55 363 66 371
rect 38 351 66 363
rect 38 349 41 351
rect -1119 320 -1061 338
rect 170 333 296 349
rect -791 304 -768 305
rect -791 301 -34 304
rect -791 284 -28 301
rect -791 274 -767 284
rect -1112 256 -767 274
rect -47 264 24 284
rect -1112 254 -775 256
rect -777 234 -32 236
rect -777 214 24 234
rect -777 213 -745 214
rect -1116 191 -1061 209
rect -1118 118 -1098 168
rect -56 152 44 168
rect 170 149 296 165
rect 251 124 284 125
rect -1118 98 -763 118
rect 251 116 254 124
rect -384 99 254 116
rect 251 97 254 99
rect 281 97 284 124
rect 251 96 284 97
rect -1119 47 -1091 74
rect -55 54 45 71
rect 172 56 296 72
rect -55 53 39 54
rect -1118 -5 -1061 13
rect -32 8 23 9
rect -790 -14 23 8
rect -790 -15 -31 -14
rect -790 -16 -713 -15
rect -1114 -33 -1080 -20
rect -790 -33 -766 -16
rect -1114 -41 -766 -33
rect -1103 -57 -766 -41
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1632488964
transform 1 0 -1102 0 1 -37
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1632488964
transform 1 0 -1107 0 1 59
box -14 -15 20 18
use sky130_hilas_m12m2  sky130_hilas_m12m2_5
timestamp 1629420194
transform 1 0 -791 0 1 103
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1629420194
transform 1 0 -1107 0 1 258
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_3
timestamp 1629420194
transform 1 0 -1105 0 1 359
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1629420194
transform 1 0 -776 0 1 514
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_2
timestamp 1629420194
transform 1 0 -778 0 1 409
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_4
timestamp 1629420194
transform 1 0 -778 0 1 221
box -9 -10 23 22
use sky130_hilas_WTA4stage01  sky130_hilas_WTA4stage01_0
timestamp 1632494644
transform 1 0 67 0 1 -19
box -54 1 229 535
use sky130_hilas_swc4x1BiasCelld3  sky130_hilas_swc4x1BiasCelld3_0
timestamp 1632494644
transform -1 0 -317 0 1 339
box -264 -400 749 250
<< labels >>
rlabel metal2 289 426 296 442 0 OUTPUT1
port 4 nsew analog default
rlabel metal2 291 333 296 349 0 OUTPUT2
port 5 nsew analog default
rlabel metal2 291 149 296 165 0 OUTPUT3
port 6 nsew analog default
rlabel metal2 291 56 296 72 0 OUTPUT4
port 7 nsew analog default
rlabel metal1 257 556 280 562 0 VGND
port 1 nsew ground default
rlabel metal1 257 -43 280 -37 0 VGND
port 1 nsew ground default
rlabel metal2 -1112 449 -1097 469 0 INPUT1
port 8 nsew analog default
rlabel metal2 -1112 352 -1086 378 0 INPUT2
port 9 nsew analog default
rlabel metal2 -1118 151 -1098 168 0 INPUT3
port 10 nsew analog default
rlabel metal2 -1119 47 -1091 74 0 INPUT4
port 11 nsew analog default
rlabel metal1 -531 552 -495 562 0 GATE1
port 16 nsew
rlabel metal1 -129 548 -89 562 0 VTUN
port 17 nsew
rlabel metal1 131 -43 154 -37 0 WTAMIDDLENODE
port 18 nsew
rlabel metal1 131 556 154 562 0 WTAMIDDLENODE
port 18 nsew
rlabel metal1 -984 555 -965 562 0 COLSEL1
port 19 nsew
rlabel metal1 -1025 555 -1009 562 0 VINJ
port 21 nsew
rlabel metal1 -944 555 -928 562 0 VPWR
port 20 nsew
rlabel metal2 -1116 515 -1107 533 0 DRAIN1
port 12 nsew
rlabel metal2 -1119 320 -1110 338 0 DRAIN2
port 22 nsew
rlabel metal2 -1116 191 -1107 209 0 DRAIN3
port 23 nsew
rlabel metal2 -1118 -5 -1109 13 0 DRAIN4
port 24 nsew
<< end >>
