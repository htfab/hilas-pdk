magic
tech sky130A
timestamp 1628704254
<< checkpaint >>
rect -557 -538 1076 751
rect -366 -599 1030 -538
rect -253 -600 1030 -599
<< error_s >>
rect 125 127 165 132
rect 351 127 391 134
rect 125 85 165 90
rect 351 85 391 92
rect 201 60 241 66
rect 351 60 391 66
rect 201 18 241 24
rect 351 18 391 24
<< nwell >>
rect 12 84 288 161
rect 12 67 211 84
rect 12 5 210 67
rect 12 0 288 5
<< pmos >>
rect 125 90 165 127
<< pdiff >>
rect 96 115 125 127
rect 96 98 102 115
rect 119 98 125 115
rect 96 90 125 98
rect 165 115 193 127
rect 165 98 171 115
rect 188 98 193 115
rect 165 90 193 98
<< pdiffc >>
rect 102 98 119 115
rect 171 98 188 115
<< nsubdiff >>
rect 36 56 68 69
rect 36 39 43 56
rect 60 39 68 56
rect 36 27 68 39
<< nsubdiffcont >>
rect 43 39 60 56
<< poly >>
rect 29 135 288 150
rect 125 127 165 135
rect 211 103 244 109
rect 125 68 165 90
rect 211 86 219 103
rect 236 86 244 103
rect 211 74 244 86
<< polycont >>
rect 219 86 236 103
<< locali >>
rect 162 115 288 116
rect 92 103 102 115
rect 75 98 102 103
rect 119 98 127 115
rect 162 98 171 115
rect 188 103 288 115
rect 188 98 219 103
rect 75 90 94 98
rect 73 87 94 90
rect 72 86 94 87
rect 211 86 219 98
rect 236 98 288 103
rect 236 86 244 98
rect 60 81 94 86
rect 47 78 94 81
rect 43 75 94 78
rect 43 69 92 75
rect 43 64 77 69
rect 43 62 69 64
rect 43 60 66 62
rect 43 56 64 60
rect 43 28 60 39
<< metal1 >>
rect 74 0 94 161
rect 425 157 444 161
rect 425 0 444 5
<< metal2 >>
rect 0 114 61 134
rect 469 114 476 134
rect 87 36 199 37
rect 0 16 199 36
rect 87 15 199 16
use sky130_hilas_li2m1  sky130_hilas_li2m1_2
timestamp 1628285143
transform 1 0 83 0 1 100
box -10 -8 13 21
use sky130_hilas_poly2m1  sky130_hilas_poly2m1_0
timestamp 1628704241
transform 1 0 27 0 1 121
box 0 0 33 51
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1628285143
transform 1 0 38 0 1 124
box -9 -10 23 22
use sky130_hilas_TgateSingle01Part1  sky130_hilas_TgateSingle01Part1_0
timestamp 1628285143
transform 1 0 31 0 1 186
box 257 -181 445 -29
use sky130_hilas_TgateSingle01Part2  sky130_hilas_TgateSingle01Part2_0
timestamp 1628285143
transform 1 0 192 0 1 186
box -67 -181 96 -38
<< labels >>
rlabel metal2 0 114 9 134 0 Select
rlabel metal2 0 16 9 36 0 Input
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
