magic
tech sky130A
timestamp 1629420194
<< poly >>
rect 142 506 162 535
rect 141 229 162 308
rect 142 1 162 30
<< metal1 >>
rect 64 258 87 278
rect 190 258 213 279
use sky130_hilas_WTAsinglestage01  sky130_hilas_WTAsinglestage01_3
timestamp 1629420194
transform 1 0 54 0 1 354
box -108 -76 175 67
use sky130_hilas_WTAsinglestage01  sky130_hilas_WTAsinglestage01_2
timestamp 1629420194
transform 1 0 54 0 -1 459
box -108 -76 175 67
use sky130_hilas_WTAsinglestage01  sky130_hilas_WTAsinglestage01_1
timestamp 1629420194
transform 1 0 54 0 -1 182
box -108 -76 175 67
use sky130_hilas_WTAsinglestage01  sky130_hilas_WTAsinglestage01_0
timestamp 1629420194
transform 1 0 54 0 1 77
box -108 -76 175 67
<< end >>
