magic
tech sky130A
timestamp 1628178864
<< error_s >>
rect 1135 598 1185 603
rect 1275 598 1325 604
rect 1455 598 1505 603
rect 1135 556 1185 561
rect 1275 556 1325 562
rect 1455 556 1505 561
rect 1135 531 1185 537
rect 1455 531 1505 537
rect 1135 489 1185 495
rect 1455 489 1505 495
rect 1135 428 1185 434
rect 1455 428 1505 434
rect 1135 386 1185 392
rect 1455 386 1505 392
rect 1135 362 1185 367
rect 1275 361 1325 367
rect 1455 362 1505 367
rect 1135 320 1185 325
rect 1275 319 1325 325
rect 1455 320 1505 325
rect 1135 278 1185 283
rect 1275 278 1325 284
rect 1455 278 1505 283
rect 1135 236 1185 241
rect 1275 236 1325 242
rect 1455 236 1505 241
rect 1135 211 1185 217
rect 1455 211 1505 217
rect 1135 169 1185 175
rect 1455 169 1505 175
rect 1135 108 1185 114
rect 1455 108 1505 114
rect 1135 66 1185 72
rect 1455 66 1505 72
rect 1135 42 1185 47
rect 1275 41 1325 47
rect 1455 42 1505 47
rect 1135 0 1185 5
rect 1275 -1 1325 5
rect 1455 0 1505 5
<< nwell >>
rect 1050 461 1392 462
rect 1050 140 1392 142
<< metal1 >>
rect 1108 603 1133 610
rect 1407 603 1430 610
rect 1542 605 1561 610
rect 1108 461 1133 462
rect 1108 141 1133 142
rect 1407 5 1430 13
rect 1542 5 1561 12
<< metal2 >>
rect 1050 567 1228 585
rect 1614 517 1622 540
rect 1607 383 1622 407
rect 1050 337 1228 353
rect 1050 258 1107 259
rect 1050 257 1177 258
rect 1050 241 1250 257
rect 1614 197 1622 220
rect 1613 63 1622 86
rect 1050 15 1228 32
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_3
timestamp 1628178864
transform 1 0 1282 0 -1 266
box -232 -45 336 125
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_2
timestamp 1628178864
transform 1 0 1282 0 1 17
box -232 -45 336 125
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_0
timestamp 1628178864
transform 1 0 1282 0 1 337
box -232 -45 336 125
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_1
timestamp 1628178864
transform 1 0 1282 0 -1 586
box -232 -45 336 125
<< labels >>
rlabel space 1107 356 1112 374 0 DRAIN2
port 3 nsew analog default
rlabel metal2 1107 241 1112 258 0 DRAIN3
port 2 nsew
rlabel metal1 1108 603 1133 610 0 VINJ
port 9 nsew power default
rlabel metal1 1407 603 1430 610 0 DRAIN_MUX
port 10 nsew analog default
rlabel metal1 1407 5 1430 13 0 DRAIN_MUX
port 10 nsew analog default
rlabel metal1 1542 5 1561 12 0 VGND
port 11 nsew ground default
rlabel metal1 1542 605 1561 610 0 VGND
port 11 nsew ground default
rlabel metal2 1611 384 1622 407 0 SELECT2
port 14 nsew
rlabel metal2 1614 517 1622 540 0 SELECT1
port 15 nsew
rlabel metal2 1614 197 1622 220 0 SELECT3
port 16 nsew
rlabel metal2 1613 63 1622 86 0 SELECT4
port 17 nsew
<< end >>
