magic
tech sky130A
magscale 1 2
timestamp 1627063652
<< error_s >>
rect 134 1906 234 1928
rect 278 1906 378 1928
rect 5798 1906 5898 1928
rect 5942 1906 6042 1928
rect 378 1844 446 1845
rect 5730 1844 5798 1845
rect 134 1822 234 1844
rect 278 1822 378 1844
rect 5798 1822 5898 1844
rect 5942 1822 6042 1844
rect 263 1781 280 1784
rect 382 1781 446 1784
rect 510 1781 588 1784
rect 780 1781 860 1784
rect 5316 1781 5396 1784
rect 5588 1781 5666 1784
rect 5730 1781 5794 1784
rect 5896 1781 5913 1784
rect 224 1572 233 1653
rect 504 1630 510 1730
rect 588 1630 594 1730
rect 776 1630 780 1730
rect 860 1630 864 1730
rect 5312 1630 5316 1730
rect 5396 1630 5400 1730
rect 5582 1630 5588 1730
rect 5666 1630 5672 1730
rect 5943 1606 5952 1653
rect 5990 1572 5999 1606
rect 504 1472 510 1572
rect 588 1472 594 1572
rect 776 1472 780 1572
rect 860 1472 864 1572
rect 5312 1472 5316 1572
rect 5396 1472 5400 1572
rect 5582 1472 5588 1572
rect 5666 1472 5672 1572
rect 224 1176 232 1210
rect 224 1132 233 1176
rect 504 1166 510 1266
rect 536 1210 662 1464
rect 790 1278 1176 1376
rect 780 1266 1176 1278
rect 576 1206 662 1210
rect 776 1230 1176 1266
rect 5284 1278 5348 1314
rect 5284 1266 5396 1278
rect 776 1208 1148 1230
rect 776 1206 894 1208
rect 920 1206 922 1208
rect 588 1166 594 1206
rect 776 1166 780 1206
rect 830 1146 998 1206
rect 1008 1146 1148 1208
rect 1318 1188 1360 1216
rect 1412 1194 1450 1222
rect 1494 1198 1536 1226
rect 1740 1210 1746 1224
rect 3888 1194 3934 1222
rect 3940 1166 3962 1238
rect 5030 1222 5166 1230
rect 5284 1222 5400 1266
rect 5030 1206 5168 1222
rect 5192 1194 5230 1222
rect 5280 1210 5400 1222
rect 5514 1241 5602 1460
rect 5514 1210 5661 1241
rect 5284 1160 5661 1210
rect 5666 1194 5672 1266
rect 5890 1244 5896 1306
rect 5910 1244 5952 1278
rect 5890 1222 5952 1244
rect 5284 1146 5624 1160
rect 5682 1154 5694 1160
rect 5678 1148 5694 1154
rect 920 1118 922 1146
rect 5382 1112 5464 1146
rect 5570 1144 5624 1146
rect 5570 1142 5612 1144
rect 5682 1142 5694 1148
rect 5562 1138 5612 1142
rect 5562 1130 5614 1138
rect 5562 1120 5660 1130
rect 5710 1124 5722 1132
rect 5562 1112 5614 1120
rect 5710 1114 5726 1124
rect 504 1008 510 1108
rect 588 1008 594 1108
rect 776 1008 780 1108
rect 790 1074 818 1110
rect 5382 1108 5465 1112
rect 5611 1108 5612 1109
rect 5673 1108 5688 1112
rect 5730 1108 5748 1172
rect 5890 1154 5980 1222
rect 6034 1180 6110 1222
rect 6122 1180 6128 1238
rect 6150 1180 6156 1210
rect 6016 1166 6150 1180
rect 5995 1154 6150 1166
rect 860 1008 864 1108
rect 5312 1008 5316 1108
rect 5382 1008 5512 1108
rect 5612 1107 5613 1108
rect 5666 1107 5688 1108
rect 5660 1096 5688 1107
rect 5610 1086 5688 1096
rect 5626 1062 5688 1086
rect 5864 1090 5952 1154
rect 5980 1136 6150 1154
rect 5980 1114 6034 1136
rect 5980 1099 6030 1114
rect 6042 1099 6150 1136
rect 5980 1090 6150 1099
rect 5864 1084 6150 1090
rect 5710 1068 5752 1070
rect 5926 1068 5984 1084
rect 5998 1070 6022 1084
rect 6030 1070 6042 1084
rect 5710 1066 5756 1068
rect 5666 1042 5688 1062
rect 5744 1053 5756 1066
rect 5758 1053 5778 1056
rect 5782 1053 5794 1068
rect 5896 1056 5984 1068
rect 5666 1039 5724 1042
rect 5615 1038 5724 1039
rect 5615 1028 5688 1038
rect 5610 1008 5688 1028
rect 5382 993 5465 1008
rect 5610 994 5660 1008
rect 5382 957 5464 993
rect 5610 962 5644 994
rect 5673 993 5688 1008
rect 5710 982 5722 1034
rect 5744 1022 5873 1053
rect 5896 1038 6022 1056
rect 5926 1022 6022 1038
rect 6030 1036 6060 1070
rect 6124 1048 6128 1084
rect 6110 1036 6150 1048
rect 6030 1022 6150 1036
rect 5744 1008 5952 1022
rect 5730 1006 5952 1008
rect 5980 1007 6150 1022
rect 5730 958 5756 1006
rect 5758 958 5778 1006
rect 5782 972 5952 1006
rect 5730 957 5748 958
rect 5782 957 5812 972
rect 263 954 280 957
rect 382 954 446 957
rect 510 954 588 957
rect 780 954 860 957
rect 5316 954 5465 957
rect 134 894 234 916
rect 278 894 378 916
rect 378 893 446 894
rect 5382 892 5422 954
rect 5450 942 5465 954
rect 5673 942 5688 957
rect 5730 956 5812 957
rect 5864 962 5952 972
rect 5984 967 6030 1007
rect 6042 967 6150 1007
rect 5980 962 6150 967
rect 5730 954 5794 956
rect 5864 954 6150 962
rect 5864 953 5913 954
rect 5926 953 6150 954
rect 5864 952 6150 953
rect 5450 908 5512 942
rect 5612 908 5688 942
rect 5926 926 5980 952
rect 5984 926 6022 952
rect 6042 948 6110 952
rect 5450 893 5465 908
rect 5670 894 5688 908
rect 5826 894 5864 916
rect 5673 893 5688 894
rect 5730 893 5798 894
rect 5730 885 5748 893
rect 5730 882 5873 885
rect 6124 884 6128 952
rect 5730 878 5906 882
rect 5680 840 5682 866
rect 5702 864 5906 878
rect 5926 878 5942 884
rect 6110 878 6150 884
rect 5702 862 5873 864
rect 5724 858 5873 862
rect 5926 858 6150 878
rect 5724 840 6110 858
rect 5730 838 6110 840
rect 134 810 234 832
rect 278 810 378 832
rect 5678 812 5682 838
rect 5724 834 6110 838
rect 5724 832 5748 834
rect 5767 832 6110 834
rect 5724 812 5730 832
rect 5748 810 5898 832
rect 5748 804 5798 810
rect 5836 802 5898 810
rect 5864 794 5879 802
rect 5980 800 6042 832
rect 6042 794 6110 800
rect 5796 789 6110 794
rect 6124 789 6150 858
rect 5796 788 6150 789
rect 5796 766 6110 788
rect 6124 764 6128 788
rect 5926 726 5980 740
rect 6152 736 6156 1180
rect 6332 1128 6366 1137
rect 5926 642 5980 656
rect 5926 562 5980 576
rect 5926 478 5980 492
rect 5926 430 5980 444
rect 5926 346 5980 360
rect 5926 266 5980 280
rect 5926 182 5980 196
rect 790 100 818 136
rect 5926 134 5980 148
rect 6285 122 6332 131
rect 5926 50 5980 64
rect 1320 2 1366 30
rect 5192 0 5230 28
rect 5280 0 5336 28
<< nwell >>
rect 790 1208 1452 1210
rect 5384 1208 5652 1210
rect 830 1146 894 1206
rect 5284 1146 5348 1206
rect 6154 1174 6410 1210
rect 6154 0 6410 38
<< metal1 >>
rect 862 1206 894 1210
rect 830 1202 894 1206
rect 830 1150 836 1202
rect 888 1150 894 1202
rect 944 1198 982 1210
rect 1318 1188 1360 1210
rect 1412 1194 1450 1210
rect 1494 1198 1536 1210
rect 1710 1196 1746 1210
rect 2942 1180 3026 1210
rect 3148 1180 3232 1210
rect 3888 1194 3934 1210
rect 5192 1194 5230 1210
rect 5280 1206 5336 1210
rect 5280 1202 5348 1206
rect 5280 1194 5290 1202
rect 2942 1152 3232 1180
rect 830 1146 894 1150
rect 5284 1150 5290 1194
rect 5342 1150 5348 1202
rect 6018 1182 6086 1210
rect 6150 1180 6206 1210
rect 5284 1146 5348 1150
rect 5712 96 5776 100
rect 2474 66 2538 70
rect 1320 2 1366 26
rect 2474 14 2480 66
rect 2532 14 2538 66
rect 2474 10 2538 14
rect 3634 66 3698 70
rect 3634 14 3640 66
rect 3692 14 3698 66
rect 5712 44 5718 96
rect 5770 44 5776 96
rect 5712 40 5776 44
rect 5712 38 6020 40
rect 5712 28 6086 38
rect 3634 10 3698 14
rect 5722 12 6086 28
rect 5192 0 5230 10
rect 5280 0 5336 10
rect 6018 0 6086 12
rect 6152 0 6206 42
<< via1 >>
rect 836 1150 888 1202
rect 5290 1150 5342 1202
rect 2480 14 2532 66
rect 3640 14 3692 66
rect 5718 44 5770 96
<< metal2 >>
rect 830 1202 894 1206
rect 830 1150 836 1202
rect 888 1182 894 1202
rect 5284 1202 5348 1206
rect 5284 1182 5290 1202
rect 888 1150 5290 1182
rect 5342 1150 5348 1202
rect 5504 1156 5566 1204
rect 830 1146 5348 1150
rect 790 1074 806 1110
rect 5726 1030 5770 1034
rect 5716 962 5770 1030
rect 5368 862 5438 906
rect 5730 848 5770 850
rect 3092 764 4690 804
rect 5730 782 5774 848
rect 5734 780 5774 782
rect 4410 628 4454 630
rect 3094 578 4460 628
rect 4646 620 4690 764
rect 5520 622 5584 670
rect 6388 668 6410 714
rect 3094 394 3796 432
rect 3750 274 3796 394
rect 4402 344 4460 578
rect 4640 612 4690 620
rect 4640 484 4692 612
rect 6388 504 6410 548
rect 4640 442 5466 484
rect 5424 414 5466 442
rect 5424 372 5798 414
rect 4402 300 4980 344
rect 4402 298 4460 300
rect 3750 244 3794 274
rect 4624 244 5798 254
rect 3750 212 5798 244
rect 3750 200 4702 212
rect 790 100 806 136
rect 5712 96 5776 100
rect 5712 70 5718 96
rect 2474 66 5718 70
rect 2474 14 2480 66
rect 2532 40 3640 66
rect 2532 14 2538 40
rect 2474 10 2538 14
rect 3634 14 3640 40
rect 3692 44 5718 66
rect 5770 44 5776 96
rect 3692 40 5776 44
rect 3692 14 3698 40
rect 3634 10 3698 14
use sky130_hilas_FGBias2x1cell  sky130_hilas_FGBias2x1cell_0
timestamp 1627063299
transform 1 0 3870 0 1 764
box 0 0 2306 1210
use sky130_hilas_FGtrans2x1cell  sky130_hilas_FGtrans2x1cell_0
timestamp 1627063299
transform -1 0 2304 0 1 764
box 0 0 2304 1210
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1608384750
transform 1 0 5116 0 -1 330
box 266 -880 640 330
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1608069483
transform 1 0 6100 0 1 82
box -344 -44 310 1100
<< labels >>
rlabel metal1 6018 1198 6086 1210 0 VGND
port 11 nsew
rlabel metal1 6150 1198 6206 1210 0 VPWR
port 10 nsew
rlabel metal1 6152 0 6206 12 0 VPWR
port 10 nsew
rlabel metal1 6018 0 6086 12 0 VGND
port 11 nsew
rlabel metal2 5520 622 5584 670 0 VIN21
port 9 nsew
rlabel metal2 5504 1156 5566 1204 1 VIN22
port 8 n
rlabel metal1 1320 2 1366 26 0 VIN12
port 18 nsew
rlabel metal1 1318 1188 1360 1210 0 VIN11
port 5 nsew
rlabel metal1 3148 1196 3232 1210 0 VTUN
port 1 nsew
rlabel metal1 2942 1196 3026 1210 0 VTUN
rlabel metal1 1494 1198 1536 1210 0 PROG
port 3 nsew
rlabel metal1 862 1198 894 1210 0 VINJ
port 6 nsew
rlabel metal1 5280 1194 5336 1210 0 VINJ
port 6 nsew
rlabel metal2 6388 668 6410 714 0 OUTPUT1
port 13 nsew
rlabel metal2 6388 504 6410 548 0 OUTPUT2
port 12 nsew
rlabel metal1 944 1198 982 1210 0 GATESEL1
port 14 nsew
rlabel metal1 5192 0 5230 10 0 GATESEL2
port 15 nsew
rlabel metal1 5280 0 5336 10 0 VINJ
port 6 nsew
rlabel metal1 5192 1194 5230 1210 0 GATESEL2
port 15 nsew
rlabel metal2 790 1074 806 1110 0 DRAIN1
port 16 nsew
rlabel metal2 790 100 806 136 0 DRAIN2
port 17 nsew
rlabel metal1 3888 1194 3934 1210 0 GATE1
port 4 nsew
rlabel metal1 1412 1194 1450 1210 0 GATE2
port 19 nsew
rlabel metal1 1710 1196 1746 1210 0 RUN
port 20 nsew
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
