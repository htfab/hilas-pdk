magic
tech sky130A
timestamp 1628704319
<< checkpaint >>
rect 49 1240 1565 1246
rect -351 1227 1565 1240
rect -580 -613 1565 1227
rect -351 -625 1565 -613
rect 49 -630 1565 -625
<< error_s >>
rect 100 579 129 597
rect 346 577 375 593
rect 425 577 454 593
rect 504 577 533 593
rect 583 577 612 593
rect 100 547 101 548
rect 128 547 129 548
rect 50 518 68 547
rect 99 546 130 547
rect 100 537 129 546
rect 100 528 110 537
rect 119 528 129 537
rect 100 519 129 528
rect 99 518 130 519
rect 161 518 179 547
rect 346 543 347 544
rect 374 543 375 544
rect 425 543 426 544
rect 453 543 454 544
rect 504 543 505 544
rect 532 543 533 544
rect 583 543 584 544
rect 611 543 612 544
rect 100 517 101 518
rect 128 517 129 518
rect 296 514 314 543
rect 345 542 376 543
rect 424 542 455 543
rect 503 542 534 543
rect 582 542 613 543
rect 346 535 375 542
rect 425 535 454 542
rect 504 535 533 542
rect 583 535 612 542
rect 346 521 356 535
rect 603 521 612 535
rect 346 515 375 521
rect 425 515 454 521
rect 504 515 533 521
rect 583 515 612 521
rect 345 514 376 515
rect 424 514 455 515
rect 503 514 534 515
rect 582 514 613 515
rect 645 514 662 543
rect 679 521 681 522
rect 346 513 347 514
rect 374 513 375 514
rect 425 513 426 514
rect 453 513 454 514
rect 504 513 505 514
rect 532 513 533 514
rect 583 513 584 514
rect 611 513 612 514
rect 100 468 129 486
rect 346 464 375 479
rect 425 464 454 479
rect 504 464 533 479
rect 583 464 612 479
rect 100 427 129 445
rect 346 430 375 446
rect 425 430 454 446
rect 504 430 533 446
rect 583 430 612 446
rect 346 396 347 397
rect 374 396 375 397
rect 425 396 426 397
rect 453 396 454 397
rect 504 396 505 397
rect 532 396 533 397
rect 583 396 584 397
rect 611 396 612 397
rect 100 395 101 396
rect 128 395 129 396
rect 50 366 68 395
rect 99 394 130 395
rect 100 385 129 394
rect 100 376 110 385
rect 119 376 129 385
rect 100 367 129 376
rect 99 366 130 367
rect 161 366 179 395
rect 296 367 314 396
rect 345 395 376 396
rect 424 395 455 396
rect 503 395 534 396
rect 582 395 613 396
rect 346 388 375 395
rect 425 388 454 395
rect 504 388 533 395
rect 583 388 612 395
rect 346 374 356 388
rect 603 374 612 388
rect 346 368 375 374
rect 425 368 454 374
rect 504 368 533 374
rect 583 368 612 374
rect 345 367 376 368
rect 424 367 455 368
rect 503 367 534 368
rect 582 367 613 368
rect 645 367 662 396
rect 674 370 687 374
rect 688 370 701 375
rect 674 367 701 370
rect 346 366 347 367
rect 374 366 375 367
rect 425 366 426 367
rect 453 366 454 367
rect 504 366 505 367
rect 532 366 533 367
rect 583 366 584 367
rect 611 366 612 367
rect 100 365 101 366
rect 128 365 129 366
rect 100 316 129 334
rect 346 317 375 332
rect 425 317 454 332
rect 504 317 533 332
rect 583 317 612 332
rect 100 282 129 300
rect 346 283 375 299
rect 425 283 454 299
rect 504 283 533 299
rect 583 283 612 299
rect 100 250 101 251
rect 128 250 129 251
rect 50 221 68 250
rect 99 249 130 250
rect 100 240 129 249
rect 100 231 110 240
rect 119 231 129 240
rect 100 222 129 231
rect 99 221 130 222
rect 161 221 179 250
rect 346 249 347 250
rect 374 249 375 250
rect 425 249 426 250
rect 453 249 454 250
rect 504 249 505 250
rect 532 249 533 250
rect 583 249 584 250
rect 611 249 612 250
rect 100 220 101 221
rect 128 220 129 221
rect 296 220 314 249
rect 345 248 376 249
rect 424 248 455 249
rect 503 248 534 249
rect 582 248 613 249
rect 346 241 375 248
rect 425 241 454 248
rect 504 241 533 248
rect 583 241 612 248
rect 346 227 356 241
rect 603 227 612 241
rect 346 221 375 227
rect 425 221 454 227
rect 504 221 533 227
rect 583 221 612 227
rect 345 220 376 221
rect 424 220 455 221
rect 503 220 534 221
rect 582 220 613 221
rect 645 220 662 249
rect 346 219 347 220
rect 374 219 375 220
rect 425 219 426 220
rect 453 219 454 220
rect 504 219 505 220
rect 532 219 533 220
rect 583 219 584 220
rect 611 219 612 220
rect 100 171 129 189
rect 346 170 375 185
rect 425 170 454 185
rect 504 170 533 185
rect 583 170 612 185
rect 100 128 129 146
rect 346 136 375 152
rect 425 136 454 152
rect 504 136 533 152
rect 583 136 612 152
rect 346 102 347 103
rect 374 102 375 103
rect 425 102 426 103
rect 453 102 454 103
rect 504 102 505 103
rect 532 102 533 103
rect 583 102 584 103
rect 611 102 612 103
rect 100 96 101 97
rect 128 96 129 97
rect 50 67 68 96
rect 99 95 130 96
rect 100 86 129 95
rect 100 77 110 86
rect 119 77 129 86
rect 100 68 129 77
rect 99 67 130 68
rect 161 67 179 96
rect 296 73 314 102
rect 345 101 376 102
rect 424 101 455 102
rect 503 101 534 102
rect 582 101 613 102
rect 346 94 375 101
rect 425 94 454 101
rect 504 94 533 101
rect 583 94 612 101
rect 346 80 356 94
rect 603 80 612 94
rect 346 74 375 80
rect 425 74 454 80
rect 504 74 533 80
rect 583 74 612 80
rect 345 73 376 74
rect 424 73 455 74
rect 503 73 534 74
rect 582 73 613 74
rect 645 73 662 102
rect 346 72 347 73
rect 374 72 375 73
rect 425 72 426 73
rect 453 72 454 73
rect 504 72 505 73
rect 532 72 533 73
rect 583 72 584 73
rect 611 72 612 73
rect 100 66 101 67
rect 128 66 129 67
rect 100 17 129 35
rect 346 23 375 38
rect 425 23 454 38
rect 504 23 533 38
rect 583 23 612 38
<< nwell >>
rect 823 315 858 316
rect 823 299 840 315
rect 857 299 858 315
<< poly >>
rect 660 534 680 538
rect 172 501 321 525
rect 660 522 679 534
rect 172 392 319 416
rect 660 378 679 395
rect 840 315 858 316
rect 856 299 858 315
rect 172 212 321 236
rect 660 220 679 237
rect 172 92 323 116
rect 660 78 679 95
<< polycont >>
rect 823 299 840 316
<< locali >>
rect 814 299 823 316
<< viali >>
rect 840 299 858 316
<< metal1 >>
rect 101 5 128 610
rect 845 319 858 321
rect 837 316 861 319
rect 837 299 840 316
rect 858 299 861 316
rect 837 296 861 299
rect 847 292 858 296
<< metal2 >>
rect 0 553 688 560
rect 0 542 691 553
rect 0 499 901 517
rect 0 411 688 417
rect 0 399 691 411
rect 0 367 687 374
rect 0 356 691 367
rect 0 241 691 258
rect 0 199 691 216
rect 0 101 691 118
rect 0 57 691 74
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_3
timestamp 1628704317
transform 1 0 112 0 1 60
box 0 0 129 129
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_2
timestamp 1628704317
transform 1 0 112 0 1 214
box 0 0 129 129
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_3
timestamp 1628704281
transform 1 0 800 0 1 59
box 0 0 400 164
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_2
timestamp 1628704281
transform 1 0 800 0 1 206
box 0 0 400 164
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_1
timestamp 1628704305
transform 1 0 968 0 1 -41
box -289 41 -33 232
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_2
timestamp 1628704305
transform 1 0 968 0 -1 356
box -289 41 -33 232
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_1
timestamp 1628704317
transform 1 0 112 0 1 359
box 0 0 129 129
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_1
timestamp 1628704281
transform 1 0 800 0 1 353
box 0 0 400 164
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_0
timestamp 1628704305
transform 1 0 968 0 1 259
box -289 41 -33 232
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_0
timestamp 1628704317
transform 1 0 112 0 1 511
box 0 0 129 129
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_0
timestamp 1628704281
transform 1 0 800 0 1 500
box 0 0 400 164
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_3
timestamp 1628704305
transform 1 0 968 0 -1 657
box -289 41 -33 232
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
