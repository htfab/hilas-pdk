magic
tech sky130A
timestamp 1632251432
<< nwell >>
rect 0 165 271 169
rect 0 0 272 165
<< mvvaractor >>
rect 104 58 215 108
<< mvnsubdiff >>
rect 33 115 215 134
rect 33 93 55 115
rect 104 108 215 115
rect 51 76 55 93
rect 33 43 55 76
rect 104 33 215 58
<< mvnsubdiffcont >>
rect 33 76 51 93
<< poly >>
rect 64 58 104 108
rect 215 58 256 108
<< locali >>
rect 30 117 53 121
rect 30 100 33 117
rect 50 100 53 117
rect 30 93 53 100
rect 30 76 33 93
rect 51 76 53 93
rect 30 72 53 76
rect 30 55 33 72
rect 50 55 53 72
rect 30 52 53 55
<< viali >>
rect 33 100 50 117
rect 33 55 50 72
<< metal1 >>
rect 28 117 54 126
rect 28 100 33 117
rect 50 100 54 117
rect 28 72 54 100
rect 28 55 33 72
rect 50 55 54 72
rect 28 47 54 55
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
