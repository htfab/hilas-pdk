magic
tech sky130A
timestamp 1628704307
<< checkpaint >>
rect -894 1680 539 2080
rect -894 1468 1615 1680
rect -894 1207 1990 1468
rect -894 1139 2365 1207
rect -894 170 2380 1139
rect -630 -230 2380 170
rect -73 -519 2380 -230
rect -73 -525 2365 -519
rect -68 -587 2365 -525
rect -68 -621 1226 -587
<< error_s >>
rect 684 616 734 622
rect 756 616 806 622
rect 684 574 734 580
rect 756 574 806 580
rect 756 547 806 553
rect 756 505 806 511
rect 756 464 806 470
rect 756 422 806 428
rect 684 395 734 401
rect 756 395 806 401
rect 684 353 734 359
rect 756 353 806 359
rect 684 292 734 298
rect 756 292 806 298
rect 684 250 734 256
rect 756 250 806 256
rect 756 223 806 229
rect 756 181 806 187
rect 756 139 806 145
rect 756 97 806 103
rect 684 70 734 76
rect 756 70 806 76
rect 684 28 734 34
rect 756 28 806 34
<< nwell >>
rect 577 622 873 623
rect 577 607 618 622
rect 1146 613 1184 623
rect 1549 609 1589 623
rect 577 606 636 607
rect 577 430 618 606
rect 566 388 618 430
rect 566 368 617 388
rect 566 315 618 368
rect 577 19 618 315
<< poly >>
rect 1887 577 1907 623
rect 1887 18 1907 43
<< locali >>
rect 563 36 581 128
<< metal1 >>
rect 653 616 669 623
rect 694 616 713 623
rect 734 616 750 623
rect 1146 613 1184 623
rect 1549 595 1589 623
rect 1809 577 1832 623
rect 1935 577 1958 623
rect 896 491 917 565
rect 566 315 587 430
rect 894 154 910 304
rect 1935 188 1958 193
rect 1931 187 1959 188
rect 1931 185 1961 187
rect 1931 158 1932 185
rect 1959 158 1961 185
rect 1931 155 1961 158
rect 1146 18 1184 28
rect 1809 18 1832 43
rect 1935 18 1958 43
<< via1 >>
rect 1932 158 1959 185
<< metal2 >>
rect 562 576 635 594
rect 920 573 1685 592
rect 920 571 1702 573
rect 1664 552 1702 571
rect 1613 551 1627 552
rect 566 488 581 530
rect 1613 518 1628 551
rect 1613 498 1734 518
rect 566 479 893 488
rect 1848 487 1974 503
rect 566 473 909 479
rect 879 463 909 473
rect 564 413 596 440
rect 1624 432 1744 442
rect 1623 424 1744 432
rect 1716 412 1744 424
rect 1716 410 1719 412
rect 559 381 617 399
rect 1848 394 1974 410
rect 887 365 910 366
rect 887 362 1644 365
rect 887 345 1650 362
rect 887 335 911 345
rect 566 317 911 335
rect 1631 325 1702 345
rect 566 315 903 317
rect 901 295 1646 297
rect 901 275 1702 295
rect 901 274 933 275
rect 562 252 617 270
rect 560 179 580 229
rect 1622 213 1722 229
rect 1848 210 1974 226
rect 1929 185 1962 186
rect 560 159 915 179
rect 1929 177 1932 185
rect 1294 160 1932 177
rect 1929 158 1932 160
rect 1959 158 1962 185
rect 1929 157 1962 158
rect 559 108 587 135
rect 1623 115 1723 132
rect 1850 117 1974 133
rect 1623 114 1717 115
rect 560 56 617 74
rect 1646 69 1701 70
rect 888 47 1701 69
rect 888 46 1647 47
rect 888 45 965 46
rect 564 28 598 41
rect 888 28 912 45
rect 564 20 912 28
rect 575 4 912 20
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628704305
transform 1 0 571 0 1 120
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628704305
transform 1 0 576 0 1 24
box 0 0 34 33
use sky130_hilas_m12m2  sky130_hilas_m12m2_4
timestamp 1628285143
transform 1 0 900 0 1 282
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_2
timestamp 1628285143
transform 1 0 900 0 1 470
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1628285143
transform 1 0 902 0 1 575
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_3
timestamp 1628285143
transform 1 0 573 0 1 420
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1628285143
transform 1 0 571 0 1 319
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_5
timestamp 1628285143
transform 1 0 887 0 1 164
box -9 -10 23 22
use sky130_hilas_WTA4stage01  sky130_hilas_WTA4stage01_0
timestamp 1628704305
transform 1 0 1745 0 1 42
box -54 1 229 535
use sky130_hilas_swc4x1BiasCell  sky130_hilas_swc4x1BiasCell_0
timestamp 1628704305
transform -1 0 1361 0 1 400
box 0 0 1625 1050
<< labels >>
rlabel metal2 1967 487 1974 503 0 OUTPUT1
port 4 nsew analog default
rlabel metal2 1969 394 1974 410 0 OUTPUT2
port 5 nsew analog default
rlabel metal2 1969 210 1974 226 0 OUTPUT3
port 6 nsew analog default
rlabel metal2 1969 117 1974 133 0 OUTPUT4
port 7 nsew analog default
rlabel metal1 1935 617 1958 623 0 VGND
port 1 nsew ground default
rlabel metal1 1935 18 1958 24 0 VGND
port 1 nsew ground default
rlabel metal2 566 510 581 530 0 INPUT1
port 8 nsew analog default
rlabel metal2 566 413 592 439 0 INPUT2
port 9 nsew analog default
rlabel metal2 560 212 580 229 0 INPUT3
port 10 nsew analog default
rlabel metal2 559 108 587 135 0 INPUT4
port 11 nsew analog default
rlabel metal1 1147 613 1183 623 0 GATE1
port 16 nsew
rlabel metal1 1549 609 1589 623 0 VTUN
port 17 nsew
rlabel metal1 1809 18 1832 24 0 WTAMIDDLENODE
port 18 nsew
rlabel metal1 1809 617 1832 623 0 WTAMIDDLENODE
port 18 nsew
rlabel metal1 694 616 713 623 0 COLSEL1
port 19 nsew
rlabel metal1 653 616 669 623 0 VINJ
port 21 nsew
rlabel metal1 734 616 750 623 0 VPWR
port 20 nsew
rlabel metal2 562 576 571 594 0 DRAIN1
port 12 nsew
rlabel metal2 559 381 568 399 0 DRAIN2
port 22 nsew
rlabel metal2 562 252 571 270 0 DRAIN3
port 23 nsew
rlabel metal2 560 56 569 74 0 DRAIN4
port 24 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
