magic
tech sky130A
timestamp 1627218289
<< error_p >>
rect -1394 -283 -1388 -277
rect -1341 -283 -1335 -277
rect -1400 -333 -1394 -327
rect -1335 -333 -1329 -327
<< nwell >>
rect -1451 -400 -1278 -210
<< mvvaractor >>
rect -1394 -333 -1335 -283
<< mvnsubdiff >>
rect -1394 -283 -1335 -247
rect -1394 -367 -1335 -333
<< poly >>
rect -1436 -333 -1394 -283
rect -1335 -333 -1293 -283
<< end >>
