VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_ta2cell_nofg
  CLASS BLOCK ;
  FOREIGN sky130_hilas_ta2cell_nofg ;
  ORIGIN 14.730 -1.400 ;
  SIZE 17.920 BY 6.050 ;
  OBS
      LAYER nwell ;
        RECT 1.920 7.270 3.190 7.450 ;
        RECT -3.280 5.710 -1.620 5.930 ;
        RECT -2.820 4.100 -2.540 4.340 ;
        RECT 1.910 1.400 3.190 1.590 ;
      LAYER met1 ;
        RECT -4.160 7.370 -3.970 7.450 ;
        RECT -3.720 7.370 -3.440 7.450 ;
        RECT 1.230 7.310 1.570 7.450 ;
        RECT 1.900 7.300 2.170 7.450 ;
        RECT 1.230 1.400 1.570 1.590 ;
        RECT 1.900 1.400 2.170 1.610 ;
      LAYER met2 ;
        RECT -1.300 7.180 -1.050 7.440 ;
        RECT -0.240 6.200 0.010 6.570 ;
        RECT -3.280 5.710 -1.620 5.930 ;
        RECT -0.210 5.350 0.000 5.640 ;
        RECT 3.040 4.740 3.190 4.960 ;
        RECT -1.260 4.510 -1.010 4.740 ;
        RECT -2.820 4.100 -2.540 4.340 ;
        RECT 3.040 3.920 3.190 4.140 ;
        RECT -1.770 3.270 0.000 3.470 ;
        RECT -3.340 2.780 -3.180 3.180 ;
        RECT -2.060 2.460 0.000 2.670 ;
        RECT -2.860 1.420 -2.600 1.670 ;
  END
END sky130_hilas_ta2cell_nofg
END LIBRARY

