magic
tech sky130A
timestamp 1608384750
<< error_s >>
rect -338 150 -332 156
rect -285 150 -279 156
rect -344 100 -338 106
rect -279 100 -273 106
rect 85 91 91 97
rect 190 91 196 97
rect 79 41 85 47
rect 196 41 202 47
rect 85 -210 91 -204
rect 190 -210 196 -204
rect -338 -264 -332 -258
rect -285 -264 -279 -258
rect 79 -260 85 -254
rect 196 -260 202 -254
rect -344 -314 -338 -308
rect -279 -314 -273 -308
<< nwell >>
rect 426 222 757 223
rect -337 -242 -281 0
<< psubdiff >>
rect -95 -42 -70 121
rect -95 -59 -92 -42
rect -73 -59 -70 -42
rect -95 -72 -70 -59
rect -95 -75 267 -72
rect -95 -76 146 -75
rect -95 -93 -71 -76
rect -52 -93 -28 -76
rect -9 -93 16 -76
rect 35 -93 56 -76
rect 75 -93 100 -76
rect 119 -92 146 -76
rect 165 -76 267 -75
rect 165 -92 190 -76
rect 119 -93 190 -92
rect 209 -93 236 -76
rect 255 -93 267 -76
rect -95 -97 267 -93
rect -95 -110 -70 -97
rect -95 -127 -92 -110
rect -73 -127 -70 -110
rect -95 -281 -70 -127
<< mvnsubdiff >>
rect -337 -242 -281 0
<< psubdiffcont >>
rect -92 -59 -73 -42
rect -71 -93 -52 -76
rect -28 -93 -9 -76
rect 16 -93 35 -76
rect 56 -93 75 -76
rect 100 -93 119 -76
rect 146 -92 165 -75
rect 190 -93 209 -76
rect 236 -93 255 -76
rect -92 -127 -73 -110
<< poly >>
rect -237 134 332 151
rect -237 126 -185 134
rect 45 91 64 134
rect 220 90 237 134
rect 46 -293 63 -260
rect 220 -293 237 -260
rect -280 -310 331 -293
<< locali >>
rect 467 28 470 45
rect -92 -42 -73 -34
rect 467 -51 472 -34
rect -92 -75 -73 -59
rect -92 -76 146 -75
rect -92 -93 -71 -76
rect -52 -93 -28 -76
rect -9 -93 16 -76
rect 35 -93 56 -76
rect 75 -93 100 -76
rect 119 -92 146 -76
rect 165 -76 263 -75
rect 165 -92 190 -76
rect 119 -93 190 -92
rect 209 -93 236 -76
rect 255 -93 263 -76
rect -92 -110 -73 -93
rect 474 -108 491 -51
rect 467 -125 469 -108
rect -92 -135 -73 -127
rect 11 -197 34 -193
rect 467 -204 470 -187
<< metal1 >>
rect -361 -382 -319 223
rect -113 -382 -90 223
rect 9 -382 32 223
rect 661 222 680 223
rect 661 -382 680 -377
rect 705 -382 733 223
<< metal2 >>
rect 484 173 516 175
rect -396 155 516 173
rect 554 49 757 71
rect 622 -98 740 -63
rect 553 -226 757 -205
rect 510 -315 526 -313
rect -396 -320 526 -315
rect -396 -330 514 -320
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_3
timestamp 1608066871
transform 1 0 1056 0 1 433
box -1451 -400 -1278 -210
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_1
timestamp 1608066871
transform 1 0 1056 0 1 19
box -1451 -400 -1278 -210
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1607179295
transform 1 0 -103 0 1 -92
box -10 -8 13 21
use sky130_hilas_wellContact  sky130_hilas_wellContact_1
timestamp 1606753443
transform 1 0 1054 0 1 404
box -1449 -441 -1275 -255
use sky130_hilas_wellContact  sky130_hilas_wellContact_0
timestamp 1606753443
transform 1 0 1054 0 1 231
box -1449 -441 -1275 -255
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_0
timestamp 1606868103
transform 1 0 986 0 1 62
box -1005 -380 -733 -211
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_2
timestamp 1606868103
transform 1 0 986 0 -1 -231
box -1005 -380 -733 -211
use sky130_hilas_horizTransCell01  sky130_hilas_horizTransCell01_1
timestamp 1607269823
transform 1 0 790 0 -1 270
box -476 48 -33 359
use sky130_hilas_horizTransCell01  sky130_hilas_horizTransCell01_0
timestamp 1607269823
transform 1 0 790 0 1 -429
box -476 48 -33 359
use sky130_hilas_m12m2  sky130_hilas_m12m2_2
timestamp 1607949437
transform 1 0 721 0 1 -84
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1607949437
transform 1 0 627 0 1 -56
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1607949437
transform 1 0 627 0 1 -116
box -9 -10 23 22
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1607089160
transform 1 0 538 0 1 -216
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1607089160
transform 1 0 538 0 1 60
box -14 -15 20 18
<< labels >>
rlabel metal1 -361 216 -319 223 0 VTUN
port 1 nsew analog default
rlabel metal1 -113 216 -90 223 0 VGND
port 2 nsew ground default
rlabel metal1 9 215 32 223 0 GATE_CONTROL
port 3 nsew analog default
rlabel metal1 705 216 733 223 0 VINJ
port 7 nsew power default
rlabel metal2 749 49 757 71 0 OUTPUT1
port 8 nsew analog default
rlabel metal2 750 -226 757 -205 0 OUTPUT2
port 9 nsew analog default
rlabel space 661 219 680 223 0 gateColSelect
rlabel metal1 -361 -382 -319 -370 0 VTUN
port 1 nsew analog default
rlabel metal1 9 -382 32 -376 0 GATE_CONTROL
port 4 nsew analog default
rlabel metal1 -113 -382 -90 -376 0 VGND
port 2 nsew ground default
rlabel metal2 -396 155 -389 173 0 DRAIN1
port 5 nsew analog default
rlabel metal2 -396 -330 -390 -315 0 DRAIN4
port 6 nsew analog default
rlabel metal1 661 -382 680 -377 0 GateColSelect
rlabel metal1 705 -382 733 -377 0 VINJ
<< end >>
