magic
tech sky130A
timestamp 1627219129
<< error_p >>
rect -500 -276 -494 -270
rect 350 -276 357 -270
rect -506 -742 -500 -736
rect 356 -742 362 -736
<< nwell >>
rect -556 -677 413 -217
rect -556 -816 473 -677
<< mvvaractor >>
rect -500 -742 356 -276
<< mvnsubdiff >>
rect -500 -276 357 -250
rect 404 -727 440 -710
rect -500 -766 356 -742
rect 404 -744 410 -727
rect 427 -744 440 -727
rect 404 -761 440 -744
rect 404 -766 410 -761
rect -500 -778 410 -766
rect 427 -778 440 -761
rect -500 -783 440 -778
<< mvnsubdiffcont >>
rect 410 -744 427 -727
rect 410 -778 427 -761
<< poly >>
rect -540 -742 -500 -276
rect 356 -742 395 -276
<< locali >>
rect 410 -727 427 -719
rect 410 -786 427 -778
<< viali >>
rect 410 -761 427 -744
<< metal1 >>
rect 407 -744 431 -734
rect 407 -761 410 -744
rect 427 -761 431 -744
rect 407 -770 431 -761
<< end >>
