* NGSPICE file created from /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_swc4x1BiasCell.ext - technology: sky130A

.subckt sky130_hilas_TunCap01 VSUBS a_n2872_n666# w_n2902_n800#
X0 a_n2872_n666# w_n2902_n800# w_n2902_n800# sky130_fd_pr__cap_var w=590000u l=500000u
.ends

.subckt sky130_hilas_horizPcell01 VSUBS a_n502_286# a_n508_162# w_n578_94# a_n578_238#
+ m1_n258_94# a_n300_94# a_n344_286#
X0 w_n578_94# a_n300_94# a_n344_162# w_n578_94# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
X1 a_n344_286# a_n578_238# a_n502_286# w_n578_94# sky130_fd_pr__pfet_g5v0d10v5 w=300000u l=500000u
X2 a_n344_162# a_n578_238# a_n508_162# w_n578_94# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
.ends

.subckt sky130_hilas_FGVaractorCapacitor VSUBS m1_n1784_n790# a_n1882_n672# w_n1914_n790#
X0 a_n1882_n672# w_n1914_n790# w_n1914_n790# sky130_fd_pr__cap_var w=1.11e+06u l=640000u
.ends

.subckt home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_swc4x1BiasCell
+ bias1 bias2 bias3 bias4 Vtun Gate Vinj Vdd GateSelect drain1 drain2 drain3 drain4
Xsky130_hilas_TunCap01_0 VSUBS a_640_n334# Vtun sky130_hilas_TunCap01
Xsky130_hilas_TunCap01_1 VSUBS a_640_n618# Vtun sky130_hilas_TunCap01
Xsky130_hilas_TunCap01_2 VSUBS a_n214_10# Vtun sky130_hilas_TunCap01
Xsky130_hilas_TunCap01_3 VSUBS a_638_270# Vtun sky130_hilas_TunCap01
Xsky130_hilas_horizPcell01_0 VSUBS bias2 drain2 Vinj a_n214_10# GateSelect GateSelect
+ Vdd sky130_hilas_horizPcell01
Xsky130_hilas_horizPcell01_1 VSUBS bias4 drain4 Vinj a_640_n618# GateSelect GateSelect
+ Vdd sky130_hilas_horizPcell01
Xsky130_hilas_horizPcell01_2 VSUBS bias3 drain3 Vinj a_640_n334# GateSelect GateSelect
+ Vdd sky130_hilas_horizPcell01
Xsky130_hilas_horizPcell01_3 VSUBS bias1 drain1 Vinj a_638_270# GateSelect GateSelect
+ Vdd sky130_hilas_horizPcell01
Xsky130_hilas_FGVaractorCapacitor_0 VSUBS Gate a_640_n618# Gate sky130_hilas_FGVaractorCapacitor
Xsky130_hilas_FGVaractorCapacitor_2 VSUBS Gate a_n214_10# Gate sky130_hilas_FGVaractorCapacitor
Xsky130_hilas_FGVaractorCapacitor_1 VSUBS Gate a_640_n334# Gate sky130_hilas_FGVaractorCapacitor
Xsky130_hilas_FGVaractorCapacitor_3 VSUBS Gate a_638_270# Gate sky130_hilas_FGVaractorCapacitor
.ends

