magic
tech sky130A
timestamp 1629420194
<< error_s >>
rect 52 825 81 841
rect 131 825 160 841
rect 210 825 239 841
rect 289 825 318 841
rect 52 791 53 792
rect 80 791 81 792
rect 131 791 132 792
rect 159 791 160 792
rect 210 791 211 792
rect 238 791 239 792
rect 289 791 290 792
rect 317 791 318 792
rect 2 762 20 791
rect 51 790 82 791
rect 130 790 161 791
rect 209 790 240 791
rect 288 790 319 791
rect 52 783 81 790
rect 131 783 160 790
rect 210 783 239 790
rect 289 783 318 790
rect 52 769 62 783
rect 309 769 318 783
rect 52 763 81 769
rect 131 763 160 769
rect 210 763 239 769
rect 289 763 318 769
rect 51 762 82 763
rect 130 762 161 763
rect 209 762 240 763
rect 288 762 319 763
rect 351 762 368 791
rect 52 761 53 762
rect 80 761 81 762
rect 131 761 132 762
rect 159 761 160 762
rect 210 761 211 762
rect 238 761 239 762
rect 289 761 290 762
rect 317 761 318 762
rect 52 712 81 727
rect 131 712 160 727
rect 210 712 239 727
rect 289 712 318 727
rect 52 545 81 561
rect 131 545 160 561
rect 210 545 239 561
rect 289 545 318 561
rect 52 511 53 512
rect 80 511 81 512
rect 131 511 132 512
rect 159 511 160 512
rect 210 511 211 512
rect 238 511 239 512
rect 289 511 290 512
rect 317 511 318 512
rect 2 482 20 511
rect 51 510 82 511
rect 130 510 161 511
rect 209 510 240 511
rect 288 510 319 511
rect 52 503 81 510
rect 131 503 160 510
rect 210 503 239 510
rect 289 503 318 510
rect 52 489 62 503
rect 309 489 318 503
rect 52 483 81 489
rect 131 483 160 489
rect 210 483 239 489
rect 289 483 318 489
rect 51 482 82 483
rect 130 482 161 483
rect 209 482 240 483
rect 288 482 319 483
rect 351 482 368 511
rect 52 481 53 482
rect 80 481 81 482
rect 131 481 132 482
rect 159 481 160 482
rect 210 481 211 482
rect 238 481 239 482
rect 289 481 290 482
rect 317 481 318 482
rect -807 463 -778 481
rect 52 432 81 447
rect 131 432 160 447
rect 210 432 239 447
rect 289 432 318 447
rect -807 431 -806 432
rect -779 431 -778 432
rect -857 402 -839 431
rect -808 430 -777 431
rect -807 421 -778 430
rect -807 412 -797 421
rect -788 412 -778 421
rect -807 403 -778 412
rect -808 402 -777 403
rect -746 402 -728 431
rect -807 401 -806 402
rect -779 401 -778 402
rect 52 390 81 406
rect 131 390 160 406
rect 210 390 239 406
rect 289 390 318 406
rect -807 352 -778 370
rect 52 356 53 357
rect 80 356 81 357
rect 131 356 132 357
rect 159 356 160 357
rect 210 356 211 357
rect 238 356 239 357
rect 289 356 290 357
rect 317 356 318 357
rect 2 327 20 356
rect 51 355 82 356
rect 130 355 161 356
rect 209 355 240 356
rect 288 355 319 356
rect 52 348 81 355
rect 131 348 160 355
rect 210 348 239 355
rect 289 348 318 355
rect 52 334 62 348
rect 309 334 318 348
rect 52 328 81 334
rect 131 328 160 334
rect 210 328 239 334
rect 289 328 318 334
rect 51 327 82 328
rect 130 327 161 328
rect 209 327 240 328
rect 288 327 319 328
rect 351 327 368 356
rect 52 326 53 327
rect 80 326 81 327
rect 131 326 132 327
rect 159 326 160 327
rect 210 326 211 327
rect 238 326 239 327
rect 289 326 290 327
rect 317 326 318 327
rect 52 277 81 292
rect 131 277 160 292
rect 210 277 239 292
rect 289 277 318 292
<< nwell >>
rect 4 697 119 714
rect 123 697 174 714
rect -15 579 385 697
rect -15 578 174 579
rect 306 578 385 579
rect 4 559 119 578
rect 123 558 174 578
rect 279 559 306 577
rect 1799 509 2073 859
rect -409 427 -387 438
<< mvnmos >>
rect 1688 764 1751 814
rect 1688 542 1751 592
rect 1688 375 1750 452
rect 1833 375 1897 430
rect 1975 375 2039 430
<< mvpmos >>
rect 1836 738 1896 793
rect 1976 738 2036 793
rect 1836 571 1896 626
rect 1976 571 2036 626
<< mvndiff >>
rect 1688 837 1751 841
rect 1688 820 1694 837
rect 1711 820 1728 837
rect 1745 820 1751 837
rect 1688 814 1751 820
rect 1688 751 1751 764
rect 1689 736 1718 737
rect 1688 621 1718 736
rect 1688 592 1751 597
rect 1688 536 1751 542
rect 1688 519 1693 536
rect 1710 519 1727 536
rect 1744 519 1751 536
rect 1688 513 1751 519
rect 1688 475 1750 483
rect 1688 458 1693 475
rect 1710 458 1727 475
rect 1744 458 1750 475
rect 1688 452 1750 458
rect 1833 453 1897 460
rect 1833 436 1840 453
rect 1857 436 1874 453
rect 1891 436 1897 453
rect 1833 430 1897 436
rect 1975 453 2039 459
rect 1975 436 1981 453
rect 1998 436 2015 453
rect 2032 436 2039 453
rect 1975 430 2039 436
rect 1688 369 1750 375
rect 1688 352 1692 369
rect 1709 352 1726 369
rect 1743 352 1750 369
rect 1688 345 1750 352
rect 1833 369 1897 375
rect 1833 352 1840 369
rect 1857 352 1874 369
rect 1891 352 1897 369
rect 1833 345 1897 352
rect 1975 369 2039 375
rect 1975 352 1981 369
rect 1998 352 2015 369
rect 2032 352 2039 369
rect 1975 346 2039 352
<< mvpdiff >>
rect 1836 816 1896 822
rect 1836 799 1840 816
rect 1857 799 1874 816
rect 1891 799 1896 816
rect 1836 793 1896 799
rect 1976 816 2036 822
rect 1976 799 1981 816
rect 1998 799 2015 816
rect 2032 799 2036 816
rect 1976 793 2036 799
rect 1836 731 1896 738
rect 1836 714 1840 731
rect 1857 714 1874 731
rect 1891 714 1896 731
rect 1836 697 1896 714
rect 1836 649 1896 667
rect 1836 632 1840 649
rect 1857 632 1874 649
rect 1891 632 1896 649
rect 1836 626 1896 632
rect 1976 731 2036 738
rect 1976 714 1981 731
rect 1998 714 2015 731
rect 2032 714 2036 731
rect 1976 697 2036 714
rect 1976 649 2036 667
rect 1976 632 1981 649
rect 1998 632 2015 649
rect 2032 632 2036 649
rect 1976 626 2036 632
rect 1836 565 1896 571
rect 1836 548 1840 565
rect 1857 548 1874 565
rect 1891 548 1896 565
rect 1836 542 1896 548
rect 1976 565 2036 571
rect 1976 548 1981 565
rect 1998 548 2015 565
rect 2032 548 2036 565
rect 1976 542 2036 548
<< mvndiffc >>
rect 1694 820 1711 837
rect 1728 820 1745 837
rect 1693 519 1710 536
rect 1727 519 1744 536
rect 1693 458 1710 475
rect 1727 458 1744 475
rect 1840 436 1857 453
rect 1874 436 1891 453
rect 1981 436 1998 453
rect 2015 436 2032 453
rect 1692 352 1709 369
rect 1726 352 1743 369
rect 1840 352 1857 369
rect 1874 352 1891 369
rect 1981 352 1998 369
rect 2015 352 2032 369
<< mvpdiffc >>
rect 1840 799 1857 816
rect 1874 799 1891 816
rect 1981 799 1998 816
rect 2015 799 2032 816
rect 1840 714 1857 731
rect 1874 714 1891 731
rect 1840 632 1857 649
rect 1874 632 1891 649
rect 1981 714 1998 731
rect 2015 714 2032 731
rect 1981 632 1998 649
rect 2015 632 2032 649
rect 1840 548 1857 565
rect 1874 548 1891 565
rect 1981 548 1998 565
rect 2015 548 2032 565
<< psubdiff >>
rect -533 637 -199 642
rect -533 620 -493 637
rect -476 620 -459 637
rect -442 620 -425 637
rect -408 620 -391 637
rect -374 620 -357 637
rect -340 620 -323 637
rect -306 620 -289 637
rect -272 620 -255 637
rect -238 620 -199 637
rect -533 616 -199 620
rect -533 597 -504 616
rect -533 580 -527 597
rect -510 580 -504 597
rect -533 568 -504 580
rect -649 563 -504 568
rect -649 555 -527 563
rect -649 538 -629 555
rect -612 538 -595 555
rect -578 538 -561 555
rect -544 546 -527 555
rect -510 546 -504 563
rect -544 538 -504 546
rect -649 530 -504 538
rect -533 529 -504 530
rect -533 512 -527 529
rect -510 512 -504 529
rect -533 495 -504 512
rect -533 478 -527 495
rect -510 478 -504 495
rect -533 461 -504 478
rect -533 444 -527 461
rect -510 444 -504 461
rect -533 427 -504 444
rect 448 603 487 636
rect 448 586 460 603
rect 477 586 487 603
rect 448 557 487 586
rect 448 540 460 557
rect 477 540 487 557
rect 448 519 487 540
rect 448 502 460 519
rect 477 502 487 519
rect 448 476 487 502
rect 448 459 460 476
rect 477 459 487 476
rect -533 410 -527 427
rect -510 410 -504 427
rect -533 393 -504 410
rect -533 376 -527 393
rect -510 376 -504 393
rect -533 359 -504 376
rect -533 342 -527 359
rect -510 342 -504 359
rect 448 421 487 459
rect 448 404 460 421
rect 477 404 487 421
rect 448 381 487 404
rect 448 364 460 381
rect 477 364 487 381
rect -533 330 -504 342
rect 448 345 487 364
rect 448 328 460 345
rect 477 328 487 345
rect 448 307 487 328
rect 448 290 459 307
rect 476 290 487 307
rect 448 274 487 290
<< mvpsubdiff >>
rect 1689 302 2043 308
rect 1689 301 1769 302
rect 1689 284 1701 301
rect 1718 284 1735 301
rect 1752 285 1769 301
rect 1786 285 1805 302
rect 1822 285 1841 302
rect 1858 285 1875 302
rect 1892 285 1909 302
rect 1926 285 1943 302
rect 1960 285 1977 302
rect 1994 285 2011 302
rect 2028 285 2043 302
rect 1752 284 2043 285
rect 1689 278 2043 284
<< mvnsubdiff >>
rect 311 688 352 696
rect 311 671 323 688
rect 340 671 352 688
rect 311 654 352 671
rect 311 637 323 654
rect 340 637 352 654
rect 311 620 352 637
rect 311 603 323 620
rect 340 603 352 620
rect 311 598 352 603
rect 312 594 352 598
rect 1836 690 1896 697
rect 1836 673 1857 690
rect 1874 673 1896 690
rect 1836 667 1896 673
rect 1976 690 2036 697
rect 1976 673 1997 690
rect 2014 673 2036 690
rect 1976 667 2036 673
rect -409 427 -387 438
<< psubdiffcont >>
rect -493 620 -476 637
rect -459 620 -442 637
rect -425 620 -408 637
rect -391 620 -374 637
rect -357 620 -340 637
rect -323 620 -306 637
rect -289 620 -272 637
rect -255 620 -238 637
rect -527 580 -510 597
rect -629 538 -612 555
rect -595 538 -578 555
rect -561 538 -544 555
rect -527 546 -510 563
rect -527 512 -510 529
rect -527 478 -510 495
rect -527 444 -510 461
rect 460 586 477 603
rect 460 540 477 557
rect 460 502 477 519
rect 460 459 477 476
rect -527 410 -510 427
rect -527 376 -510 393
rect -527 342 -510 359
rect 460 404 477 421
rect 460 364 477 381
rect 460 328 477 345
rect 459 290 476 307
<< mvpsubdiffcont >>
rect 1701 284 1718 301
rect 1735 284 1752 301
rect 1769 285 1786 302
rect 1805 285 1822 302
rect 1841 285 1858 302
rect 1875 285 1892 302
rect 1909 285 1926 302
rect 1943 285 1960 302
rect 1977 285 1994 302
rect 2011 285 2028 302
<< mvnsubdiffcont >>
rect 323 671 340 688
rect 323 637 340 654
rect 323 603 340 620
rect 1857 673 1874 690
rect 1997 673 2014 690
<< poly >>
rect -708 746 -680 796
rect -705 679 -680 746
rect -186 716 -137 803
rect 1477 801 1688 814
rect -186 714 8 716
rect 291 714 342 715
rect 365 714 561 801
rect 1476 764 1688 801
rect 1751 764 1764 814
rect 1912 815 1920 831
rect 1912 793 1932 815
rect 2053 814 2062 831
rect 2050 793 2068 814
rect 1476 750 1530 764
rect 1822 738 1836 793
rect 1896 738 1932 793
rect 1960 738 1976 793
rect 2036 738 2068 793
rect -186 679 160 714
rect -817 655 160 679
rect -817 476 -779 655
rect -186 559 160 655
rect 1734 658 1781 692
rect 1765 592 1781 658
rect 1912 626 1932 738
rect 2051 626 2068 738
rect 291 577 342 578
rect 279 559 342 577
rect -186 558 8 559
rect 109 558 160 559
rect -186 433 -137 558
rect 1673 542 1688 592
rect 1751 542 1781 592
rect 1822 571 1836 626
rect 1896 571 1932 626
rect 1962 571 1976 626
rect 2036 571 2068 626
rect 1776 495 1814 496
rect -186 404 103 433
rect 1758 457 1814 495
rect 1758 452 1779 457
rect -186 349 -137 404
rect 1673 375 1688 452
rect 1750 437 1779 452
rect 1750 375 1764 437
rect 1817 375 1833 430
rect 1897 375 1975 430
rect 2039 375 2052 430
<< locali >>
rect 1686 820 1694 837
rect 1745 820 1753 837
rect 1916 816 1924 831
rect 2053 817 2062 831
rect 1973 816 2073 817
rect 1832 799 1840 816
rect 1891 799 1933 816
rect 1973 799 1981 816
rect 2032 799 2073 816
rect 1832 714 1840 731
rect 1891 714 1981 731
rect 2032 714 2040 731
rect 323 688 340 696
rect 1840 673 1857 690
rect 1891 673 1980 690
rect 2014 673 2022 690
rect 323 661 340 671
rect 323 654 383 661
rect -527 637 -510 639
rect 340 637 383 654
rect -527 620 -493 637
rect -476 620 -459 637
rect -442 620 -425 637
rect -408 620 -391 637
rect -374 620 -357 637
rect -340 620 -323 637
rect -306 620 -289 637
rect -272 620 -255 637
rect -238 620 -221 637
rect 323 635 383 637
rect 323 620 340 635
rect 1832 632 1840 649
rect 1891 632 1981 649
rect 2032 632 2040 649
rect -527 597 -510 620
rect 323 595 340 603
rect 460 603 477 614
rect -527 563 -510 580
rect -637 538 -629 555
rect -612 538 -595 555
rect -578 538 -561 555
rect -544 546 -527 555
rect -544 538 -510 546
rect -527 529 -510 538
rect -527 495 -510 512
rect -527 461 -510 478
rect -527 427 -510 444
rect -527 393 -510 410
rect -527 359 -510 376
rect 460 557 477 586
rect 1832 548 1840 565
rect 1891 548 1900 565
rect 1973 548 1981 565
rect 2032 548 2040 565
rect 460 519 477 540
rect 1685 519 1693 536
rect 1710 519 1727 536
rect 1744 519 1799 536
rect 460 476 477 502
rect 460 421 477 459
rect 1685 458 1693 475
rect 1744 458 1752 475
rect 1832 436 1840 453
rect 1891 436 1920 453
rect 1973 436 1981 453
rect 2032 436 2040 453
rect 460 381 477 404
rect 460 349 477 364
rect 1683 352 1692 369
rect 1709 352 1726 369
rect 1743 352 1840 369
rect 1857 352 1874 369
rect 1891 352 1981 369
rect 1998 352 2015 369
rect 2032 352 2041 369
rect -527 297 -510 342
rect 459 345 477 349
rect 459 328 460 345
rect 459 307 477 328
rect 476 290 477 307
rect 1710 302 1778 307
rect 1710 301 1769 302
rect 459 276 477 290
rect 1693 284 1701 301
rect 1718 284 1735 301
rect 1752 285 1769 301
rect 1786 285 1805 302
rect 1822 285 1841 302
rect 1858 285 1875 302
rect 1892 285 1909 302
rect 1926 285 1943 302
rect 1960 285 1977 302
rect 1994 285 2011 302
rect 2028 285 2036 302
rect 1752 284 1778 285
<< viali >>
rect 1711 820 1728 837
rect 1857 799 1874 816
rect 1998 799 2015 816
rect 1857 714 1874 731
rect 1998 714 2015 731
rect 1874 673 1891 690
rect 1980 673 1997 690
rect 1857 632 1874 649
rect 1998 632 2015 649
rect 1857 548 1874 565
rect 1998 548 2015 565
rect 1710 458 1727 475
rect 1857 436 1874 453
rect 1998 436 2015 453
<< metal1 >>
rect -884 775 -858 864
rect -414 739 -387 864
rect 173 823 197 864
rect 1705 837 1734 840
rect 1705 820 1711 837
rect 1728 820 1734 837
rect 1705 817 1734 820
rect 1781 816 1884 824
rect 1781 799 1857 816
rect 1874 799 1884 816
rect 1781 793 1884 799
rect 1987 816 2025 824
rect 1987 799 1998 816
rect 2015 799 2025 816
rect 1987 793 2025 799
rect 1706 748 1733 761
rect 1697 739 1733 748
rect 1697 719 1739 739
rect 1697 625 1720 719
rect 1697 607 1733 625
rect -805 277 -780 464
rect -806 259 -780 277
rect -415 259 -384 518
rect 1706 478 1733 607
rect 1781 516 1805 793
rect 1854 731 1877 737
rect 1854 714 1857 731
rect 1874 714 1877 731
rect 1994 731 2018 737
rect 1994 714 1998 731
rect 2015 714 2018 731
rect 1849 690 2024 714
rect 1849 673 1874 690
rect 1891 673 1980 690
rect 1997 673 2024 690
rect 1849 649 2024 673
rect 1849 648 1857 649
rect 1854 632 1857 648
rect 1874 648 1998 649
rect 1874 632 1877 648
rect 1854 626 1877 632
rect 1994 632 1998 648
rect 2015 648 2024 649
rect 2015 632 2018 648
rect 1994 626 2018 632
rect 1854 565 1877 571
rect 1854 548 1857 565
rect 1874 548 1877 565
rect 1700 475 1733 478
rect 1700 458 1710 475
rect 1727 458 1733 475
rect 1700 455 1733 458
rect 1854 453 1877 548
rect 174 259 198 447
rect 1854 436 1857 453
rect 1874 436 1877 453
rect 1854 430 1877 436
rect 1995 565 2018 571
rect 1995 548 1998 565
rect 2015 548 2018 565
rect 1995 453 2018 548
rect 1995 436 1998 453
rect 2015 436 2018 453
rect 1995 430 2018 436
rect 1505 259 1534 365
<< metal2 >>
rect 1704 817 1993 841
rect 351 718 1816 731
rect 351 710 2083 718
rect 174 640 204 686
rect 247 641 277 687
rect 385 643 409 710
rect 1802 693 2083 710
rect 1738 559 1765 687
rect 1816 642 2083 693
rect 1738 558 2017 559
rect 1738 536 2083 558
rect 1790 535 2083 536
rect 2021 487 2083 519
rect 1780 448 2083 471
rect 1695 321 2083 354
rect 1694 312 2083 321
rect 1695 305 2083 312
rect 1719 287 1763 305
rect -531 266 1792 287
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_1
timestamp 1629420194
transform 1 0 563 0 1 1073
box -1005 -380 -733 -211
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_2
timestamp 1629420194
transform 1 0 563 0 1 774
box -1005 -380 -733 -211
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_0
timestamp 1629420194
transform 1 0 563 0 1 673
box -1005 -380 -733 -211
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_0
timestamp 1629420194
transform 1 0 -795 0 1 395
box -62 -43 67 86
use sky130_hilas_FGVaractorTunnelCap01  sky130_hilas_FGVaractorTunnelCap01_0
timestamp 1629420194
transform 1 0 93 0 1 1068
box -1005 -380 -783 -211
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_0
timestamp 1629420194
transform 1 0 506 0 1 748
box -521 -54 -121 110
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_2
timestamp 1629420194
transform 1 0 506 0 1 313
box -521 -54 -121 110
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_1
timestamp 1629420194
transform 1 0 506 0 1 468
box -521 -54 -121 110
use sky130_hilas_li2m2  sky130_hilas_li2m2_14
timestamp 1629420194
transform 1 0 -520 0 1 283
box -14 -15 20 18
use sky130_hilas_FGHugeVaractorCapacitor01  sky130_hilas_FGHugeVaractorCapacitor01_0
timestamp 1629420194
transform 1 0 1099 0 1 1077
box -556 -816 473 -217
use sky130_hilas_pFETdevice01w1  sky130_hilas_pFETdevice01w1_0
timestamp 1629420194
transform 1 0 224 0 1 655
box -79 -78 82 43
use sky130_hilas_li2m2  sky130_hilas_li2m2_11
timestamp 1629420194
transform 1 0 394 0 1 647
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_12
timestamp 1629420194
transform 1 0 258 0 1 655
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_13
timestamp 1629420194
transform 1 0 189 0 1 654
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1629420194
transform 1 0 466 0 1 281
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_9
timestamp 1629420194
transform 1 0 1706 0 1 298
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_6
timestamp 1629420194
transform 1 0 1851 0 1 299
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_5
timestamp 1629420194
transform 1 0 1777 0 1 299
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_4
timestamp 1629420194
transform 1 0 1792 0 1 359
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_8
timestamp 1629420194
transform 1 0 2014 0 1 299
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_7
timestamp 1629420194
transform 1 0 1921 0 1 299
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1629420194
transform 1 0 1935 0 1 357
box -14 -15 20 18
use sky130_hilas_poly2li  sky130_hilas_poly2li_5
timestamp 1629420194
transform -1 0 1805 0 -1 480
box -9 -14 18 19
use sky130_hilas_li2m2  sky130_hilas_li2m2_10
timestamp 1629420194
transform -1 0 1795 0 -1 479
box -14 -15 20 18
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1629420194
transform 1 0 1791 0 1 524
box -10 -8 13 21
use sky130_hilas_poly2li  sky130_hilas_poly2li_3
timestamp 1629420194
transform 1 0 1921 0 1 440
box -9 -14 18 19
use sky130_hilas_m12m2  sky130_hilas_m12m2_9
timestamp 1629420194
transform 1 0 2000 0 1 497
box -9 -10 23 22
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_0
timestamp 1629420194
transform 1 0 1743 0 1 666
box -9 -26 24 29
use sky130_hilas_nDiffThOxContact  sky130_hilas_nDiffThOxContact_3
timestamp 1629420194
transform 1 0 1712 0 1 580
box -26 13 41 42
use sky130_hilas_m12m2  sky130_hilas_m12m2_6
timestamp 1629420194
transform 1 0 1859 0 1 720
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_4
timestamp 1629420194
transform 1 0 1857 0 1 634
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1629420194
transform 1 0 1859 0 1 676
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_3
timestamp 1629420194
transform 1 0 2000 0 1 632
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_2
timestamp 1629420194
transform 1 0 2000 0 1 719
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1629420194
transform 1 0 2000 0 1 674
box -9 -10 23 22
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1629420194
transform 1 0 1933 0 1 721
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1629420194
transform 1 0 1933 0 1 637
box -14 -15 20 18
use sky130_hilas_nDiffThOxContact  sky130_hilas_nDiffThOxContact_0
timestamp 1629420194
transform 1 0 1712 0 1 723
box -26 13 41 42
use sky130_hilas_m12m2  sky130_hilas_m12m2_10
timestamp 1629420194
transform 1 0 1713 0 1 827
box -9 -10 23 22
use sky130_hilas_poly2li  sky130_hilas_poly2li_1
timestamp 1629420194
transform 1 0 1924 0 1 828
box -9 -14 18 19
use sky130_hilas_m12m2  sky130_hilas_m12m2_7
timestamp 1629420194
transform 1 0 1999 0 1 822
box -9 -10 23 22
use sky130_hilas_poly2li  sky130_hilas_poly2li_4
timestamp 1629420194
transform 1 0 2064 0 1 828
box -9 -14 18 19
<< labels >>
rlabel metal2 2077 305 2083 354 0 VGND
port 8 nsew ground default
rlabel metal2 2077 487 2083 519 0 OUTPUT
port 10 nsew analog default
rlabel metal2 2076 642 2083 718 0 VINJ
port 9 nsew power default
rlabel metal2 2077 448 2083 471 0 VBIAS
port 12 nsew analog default
rlabel metal2 2077 535 2083 558 0 VREF
port 11 nsew analog default
rlabel metal1 1505 261 1534 266 0 LARGECAPACITOR
port 7 nsew analog default
rlabel metal1 173 858 197 864 0 GATE3
port 3 nsew analog default
rlabel metal1 174 259 198 266 0 GATE4
port 6 nsew analog default
rlabel metal1 -415 259 -384 266 0 GATE2
port 5 nsew analog default
rlabel metal1 -414 855 -387 864 0 GATE1
port 2 nsew analog default
rlabel metal1 -806 259 -780 269 0 VTUNOVERLAP01
port 4 nsew analog default
rlabel metal1 -884 857 -858 864 0 VTUN
port 1 nsew analog default
rlabel metal2 174 675 204 686 0 DRAIN1
port 13 nsew
rlabel metal2 247 676 276 687 0 SOURCE1
port 14 nsew
<< end >>
