magic
tech sky130A
timestamp 1628698485
<< checkpaint >>
rect -1933 -709 334 1201
<< error_s >>
rect -872 485 -866 491
rect -767 485 -761 491
rect -1246 475 -1240 481
rect -1193 475 -1187 481
rect -1252 425 -1246 431
rect -1187 425 -1181 431
rect -878 421 -872 427
rect -761 421 -755 427
rect -1246 366 -1240 372
rect -1193 366 -1187 372
rect -872 368 -866 374
rect -767 368 -761 374
rect -1252 316 -1246 322
rect -1187 316 -1181 322
rect -878 304 -872 310
rect -761 304 -755 310
rect 2331 228 2333 256
rect -872 183 -866 189
rect -767 183 -761 189
rect -1246 177 -1240 183
rect -1193 177 -1187 183
rect -1252 127 -1246 133
rect -1187 127 -1181 133
rect -878 119 -872 125
rect -761 119 -755 125
rect -872 67 -866 73
rect -767 67 -761 73
rect -1246 60 -1240 66
rect -1193 60 -1187 66
rect -1252 10 -1246 16
rect -1187 10 -1181 16
rect -878 3 -872 9
rect -761 3 -755 9
<< nwell >>
rect -297 547 2238 548
rect -296 540 2238 547
rect -1303 480 -1292 498
rect -1304 294 -1292 312
rect -1302 -5 -1292 12
rect -298 -51 2238 540
rect -297 -56 2238 -51
rect -104 -57 2238 -56
<< metal1 >>
rect -1268 534 -1228 548
rect -1024 542 -1000 548
rect -862 540 -825 548
rect -631 541 -607 548
rect -392 543 -373 548
rect -348 543 -332 548
rect -863 535 -825 540
rect -864 -44 -863 -42
rect -1268 -57 -1229 -45
rect -1024 -57 -1000 -50
rect -864 -56 -825 -44
rect -864 -57 -863 -56
rect -631 -57 -607 -50
rect -429 -56 -413 -50
rect -392 -56 -373 -50
rect -348 -56 -332 -50
<< metal2 >>
rect -230 545 -179 548
rect -230 543 -137 545
rect -230 536 -174 543
rect -416 517 -174 536
rect -187 515 -174 517
rect -146 515 -137 543
rect -1303 480 -1292 498
rect -406 480 2366 498
rect -412 437 2366 455
rect -406 337 2366 355
rect 2265 312 2366 313
rect -1304 294 -1292 312
rect -410 294 2366 312
rect 2297 256 2366 263
rect 2297 228 2304 256
rect 2333 228 2366 256
rect 2297 222 2366 228
rect -1302 179 -1292 196
rect -427 179 2366 196
rect -417 137 2366 154
rect -419 39 2366 56
rect -1302 -5 -1292 12
rect -423 -5 2366 12
<< via2 >>
rect -174 515 -146 543
rect 2304 228 2333 256
<< metal3 >>
rect -179 543 -141 546
rect -179 517 -174 543
rect -187 515 -174 517
rect -146 517 -141 543
rect -146 515 -133 517
rect -187 392 -133 515
rect 2219 256 2334 327
rect 2219 228 2304 256
rect 2333 228 2334 256
rect -267 143 -249 173
rect 2219 163 2334 228
rect 2264 162 2334 163
rect -158 22 -140 52
<< metal4 >>
rect -25 481 385 511
rect -194 420 76 431
rect -194 390 97 420
rect 46 356 97 390
rect 347 361 385 481
rect 631 364 959 394
rect -263 318 -127 348
rect -157 262 -127 318
rect 631 262 661 364
rect 929 262 959 364
rect -157 232 959 262
rect 1199 362 2088 392
rect 67 173 386 176
rect 631 173 661 176
rect -267 143 953 173
rect 67 106 97 143
rect 356 109 386 143
rect 631 109 661 143
rect 356 106 661 109
rect 923 106 953 143
rect 67 76 953 106
rect 1199 110 1229 362
rect 1482 359 1793 362
rect 1482 110 1512 359
rect 1763 110 1793 359
rect 2058 110 2088 362
rect 1199 80 2094 110
rect 1763 79 2094 80
rect -170 22 -119 52
rect -149 -2 -119 22
rect 2064 -2 2094 79
rect -149 -32 2094 -2
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_1
timestamp 1628285143
transform 1 0 -1040 0 1 325
box -263 -404 744 246
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_0
timestamp 1628285143
transform 1 0 -1040 0 1 325
box -263 -404 744 246
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1628285143
transform 1 0 -428 0 1 524
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1628285143
transform 1 0 -428 0 1 524
box -9 -10 23 22
use sky130_hilas_m22m4  sky130_hilas_m22m4_3
timestamp 1607701799
transform 1 0 -197 0 1 52
box -36 -36 43 39
use sky130_hilas_m22m4  sky130_hilas_m22m4_2
timestamp 1607701799
transform 1 0 -306 0 1 139
box -36 -36 43 39
use sky130_hilas_m22m4  sky130_hilas_m22m4_1
timestamp 1607701799
transform 1 0 -302 0 1 348
box -36 -36 43 39
<< labels >>
rlabel metal2 2354 222 2366 263 0 CAPTERM2
port 1 nsew analog default
rlabel metal2 -230 535 -179 548 0 CAPTERM1
port 2 nsew analog default
rlabel metal1 -392 543 -373 548 0 GATESELECT
port 4 nsew
rlabel metal1 -348 543 -332 548 0 VINJ
port 3 nsew power default
rlabel metal1 -862 535 -825 548 0 GATE
port 6 nsew analog default
rlabel metal1 -1268 534 -1228 548 0 VTUN
port 5 nsew
rlabel metal1 -1268 -57 -1229 -45 0 VTUN
port 5 nsew
rlabel metal1 -864 -56 -825 -44 0 GATE
port 6 nsew
rlabel metal1 -348 -56 -332 -50 0 VINJ
rlabel metal1 -429 -56 -413 -50 0 CAPTERM1
rlabel metal1 -392 -56 -373 -50 0 GATESELECT
rlabel metal2 -1303 480 -1292 498 0 DRAIN1
port 8 nsew
rlabel metal2 -1304 294 -1292 312 0 DRAIN2
port 7 nsew
rlabel metal2 2356 -5 2366 12 0 DRAIN4
port 10 nsew
rlabel metal2 2356 480 2366 498 0 DRAIN1
port 8 nsew
rlabel metal2 2355 294 2366 313 0 DRAIN2
port 7 nsew
rlabel metal2 2355 179 2366 196 0 DRAIN3
port 11 nsew
rlabel metal2 -1302 179 -1292 196 0 DRAIN3
port 11 nsew
rlabel metal2 -1302 -5 -1292 12 0 DRAIN4
port 10 nsew
rlabel metal1 -1024 542 -1000 548 0 VGND
port 12 nsew
rlabel metal1 -631 541 -607 548 0 VGND
port 12 nsew
rlabel metal1 -1024 -57 -1000 -50 0 VGND
port 12 nsew
rlabel metal1 -631 -57 -607 -50 0 VGND
port 12 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
