magic
tech sky130A
timestamp 1629137209
<< checkpaint >>
rect -630 -592 913 1126
<< poly >>
rect 88 505 108 534
rect 87 228 108 307
rect 88 0 108 29
<< metal1 >>
rect 10 257 33 277
rect 136 257 159 278
use sky130_hilas_WTAsinglestage01  sky130_hilas_WTAsinglestage01_0
timestamp 1629137201
transform 1 0 0 0 1 76
box 0 0 283 143
use sky130_hilas_WTAsinglestage01  sky130_hilas_WTAsinglestage01_1
timestamp 1629137201
transform 1 0 0 0 -1 181
box 0 0 283 143
use sky130_hilas_WTAsinglestage01  sky130_hilas_WTAsinglestage01_2
timestamp 1629137201
transform 1 0 0 0 -1 458
box 0 0 283 143
use sky130_hilas_WTAsinglestage01  sky130_hilas_WTAsinglestage01_3
timestamp 1629137201
transform 1 0 0 0 1 353
box 0 0 283 143
<< end >>
