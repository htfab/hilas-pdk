magic
tech sky130A
timestamp 1628616713
<< checkpaint >>
rect 1412 46462 4052 47207
rect 1412 39646 4200 46462
rect 963 39423 37101 39646
rect 961 38023 37101 39423
rect -505 37951 37101 38023
rect -505 36917 37790 37951
rect -505 8035 4200 36917
rect 11272 30331 26709 36917
rect 11272 30093 26351 30331
rect 12066 29538 26351 30093
rect 35302 29981 37790 36917
rect 35302 16678 40002 29981
rect -505 -404 1987 8035
rect 37426 7963 40002 16678
<< error_s >>
rect 14842 37094 14871 37110
rect 14921 37094 14950 37110
rect 15000 37094 15029 37110
rect 15079 37094 15108 37110
rect 14966 37071 14983 37072
rect 14842 37060 14843 37061
rect 14870 37060 14871 37061
rect 14921 37060 14922 37061
rect 14949 37060 14950 37061
rect 15000 37060 15001 37061
rect 15028 37060 15029 37061
rect 15079 37060 15080 37061
rect 15107 37060 15108 37061
rect 14792 37031 14809 37060
rect 14841 37059 14872 37060
rect 14920 37059 14951 37060
rect 14999 37059 15030 37060
rect 15078 37059 15109 37060
rect 14842 37052 14871 37059
rect 14921 37052 14950 37059
rect 14966 37052 14983 37053
rect 15000 37052 15029 37059
rect 15079 37052 15108 37059
rect 14842 37038 14851 37052
rect 15098 37038 15108 37052
rect 14842 37032 14871 37038
rect 14921 37032 14950 37038
rect 14966 37036 14983 37038
rect 15000 37032 15029 37038
rect 15079 37032 15108 37038
rect 14841 37031 14872 37032
rect 14920 37031 14951 37032
rect 14999 37031 15030 37032
rect 15078 37031 15109 37032
rect 15140 37031 15158 37060
rect 14842 37030 14843 37031
rect 14870 37030 14871 37031
rect 14921 37030 14922 37031
rect 14949 37030 14950 37031
rect 15000 37030 15001 37031
rect 15028 37030 15029 37031
rect 15079 37030 15080 37031
rect 15107 37030 15108 37031
rect 14966 37017 14983 37019
rect 14842 36981 14871 36996
rect 14921 36981 14950 36996
rect 15000 36981 15029 36996
rect 15079 36981 15108 36996
rect 14915 36944 14954 36947
rect 14915 36902 14954 36905
rect 14842 36814 14871 36830
rect 14921 36814 14950 36830
rect 15000 36814 15029 36830
rect 15079 36814 15108 36830
rect 14966 36791 14983 36792
rect 14842 36780 14843 36781
rect 14870 36780 14871 36781
rect 14921 36780 14922 36781
rect 14949 36780 14950 36781
rect 15000 36780 15001 36781
rect 15028 36780 15029 36781
rect 15079 36780 15080 36781
rect 15107 36780 15108 36781
rect 14792 36751 14809 36780
rect 14841 36779 14872 36780
rect 14920 36779 14951 36780
rect 14999 36779 15030 36780
rect 15078 36779 15109 36780
rect 14842 36772 14871 36779
rect 14921 36772 14950 36779
rect 14966 36772 14983 36773
rect 15000 36772 15029 36779
rect 15079 36772 15108 36779
rect 14842 36758 14851 36772
rect 15098 36758 15108 36772
rect 14842 36752 14871 36758
rect 14921 36752 14950 36758
rect 14966 36756 14983 36758
rect 15000 36752 15029 36758
rect 15079 36752 15108 36758
rect 14841 36751 14872 36752
rect 14920 36751 14951 36752
rect 14999 36751 15030 36752
rect 15078 36751 15109 36752
rect 15140 36751 15158 36780
rect 14842 36750 14843 36751
rect 14870 36750 14871 36751
rect 14921 36750 14922 36751
rect 14949 36750 14950 36751
rect 15000 36750 15001 36751
rect 15028 36750 15029 36751
rect 15079 36750 15080 36751
rect 15107 36750 15108 36751
rect 14966 36737 14983 36739
rect 15938 36732 15967 36750
rect 14842 36701 14871 36716
rect 14921 36701 14950 36716
rect 15000 36701 15029 36716
rect 15079 36701 15108 36716
rect 15938 36700 15939 36701
rect 15966 36700 15967 36701
rect 14842 36659 14871 36675
rect 14921 36659 14950 36675
rect 15000 36659 15029 36675
rect 15079 36659 15108 36675
rect 15888 36671 15906 36700
rect 15937 36699 15968 36700
rect 15938 36690 15967 36699
rect 15938 36681 15948 36690
rect 15957 36681 15967 36690
rect 15938 36672 15967 36681
rect 15937 36671 15968 36672
rect 15999 36671 16017 36700
rect 15938 36670 15939 36671
rect 15966 36670 15967 36671
rect 14966 36636 14983 36637
rect 14842 36625 14843 36626
rect 14870 36625 14871 36626
rect 14921 36625 14922 36626
rect 14949 36625 14950 36626
rect 15000 36625 15001 36626
rect 15028 36625 15029 36626
rect 15079 36625 15080 36626
rect 15107 36625 15108 36626
rect 14792 36596 14809 36625
rect 14841 36624 14872 36625
rect 14920 36624 14951 36625
rect 14999 36624 15030 36625
rect 15078 36624 15109 36625
rect 14842 36617 14871 36624
rect 14921 36617 14950 36624
rect 14966 36617 14983 36618
rect 15000 36617 15029 36624
rect 15079 36617 15108 36624
rect 14842 36603 14851 36617
rect 15098 36603 15108 36617
rect 14842 36597 14871 36603
rect 14921 36597 14950 36603
rect 14966 36601 14983 36603
rect 15000 36597 15029 36603
rect 15079 36597 15108 36603
rect 14841 36596 14872 36597
rect 14920 36596 14951 36597
rect 14999 36596 15030 36597
rect 15078 36596 15109 36597
rect 15140 36596 15158 36625
rect 15938 36621 15967 36639
rect 14842 36595 14843 36596
rect 14870 36595 14871 36596
rect 14921 36595 14922 36596
rect 14949 36595 14950 36596
rect 15000 36595 15001 36596
rect 15028 36595 15029 36596
rect 15079 36595 15080 36596
rect 15107 36595 15108 36596
rect 14966 36582 14983 36584
rect 14842 36546 14871 36561
rect 14921 36546 14950 36561
rect 15000 36546 15029 36561
rect 15079 36546 15108 36561
rect 16710 35907 16738 35923
rect 16852 35907 16880 35923
rect 16987 35913 17037 35922
rect 17320 35916 17370 35927
rect 16956 35907 16987 35913
rect 17286 35910 17320 35916
rect 16764 35881 16769 35886
rect 16710 35865 16738 35881
rect 16852 35865 16880 35881
rect 16987 35871 17037 35880
rect 17204 35873 17221 35878
rect 17320 35874 17370 35885
rect 17377 35865 17394 35866
rect 16661 35844 16689 35861
rect 16901 35844 16929 35861
rect 17058 35845 17109 35855
rect 17249 35854 17299 35865
rect 17377 35846 17394 35847
rect 17122 35840 17141 35845
rect 16661 35802 16689 35819
rect 16901 35802 16929 35819
rect 17027 35813 17058 35819
rect 17136 35813 17141 35840
rect 17217 35823 17249 35828
rect 17058 35803 17109 35813
rect 17249 35812 17299 35823
rect 16710 35752 16738 35768
rect 16852 35752 16880 35768
rect 16987 35758 17037 35767
rect 17320 35761 17370 35772
rect 16956 35752 16987 35758
rect 17286 35755 17320 35761
rect 16764 35726 16769 35731
rect 16710 35710 16738 35726
rect 16852 35710 16880 35726
rect 16987 35716 17037 35725
rect 17204 35718 17221 35723
rect 17320 35719 17370 35730
rect 17377 35710 17394 35711
rect 16661 35689 16689 35706
rect 16901 35689 16929 35706
rect 17058 35690 17109 35700
rect 17249 35699 17299 35710
rect 17377 35691 17394 35692
rect 17122 35685 17141 35690
rect 14525 35645 14552 35652
rect 16661 35647 16689 35664
rect 16901 35647 16929 35664
rect 17027 35658 17058 35664
rect 17136 35658 17141 35685
rect 17217 35668 17249 35673
rect 17058 35648 17109 35658
rect 17249 35657 17299 35668
rect 14525 35603 14552 35610
rect 16710 35597 16738 35613
rect 16852 35597 16880 35613
rect 16987 35603 17037 35612
rect 17320 35606 17370 35617
rect 18164 35608 18214 35619
rect 18236 35608 18286 35619
rect 20205 35608 20255 35619
rect 20277 35608 20327 35619
rect 20665 35614 20692 35621
rect 16956 35597 16987 35603
rect 17286 35600 17320 35606
rect 20868 35601 20885 35606
rect 18286 35577 18320 35578
rect 20171 35577 20205 35578
rect 16764 35571 16769 35576
rect 14525 35553 14552 35560
rect 16710 35555 16738 35571
rect 16852 35555 16880 35571
rect 16987 35561 17037 35570
rect 17204 35563 17221 35568
rect 17320 35564 17370 35575
rect 18164 35566 18214 35577
rect 18236 35566 18286 35577
rect 20205 35566 20255 35577
rect 20277 35566 20327 35577
rect 20665 35572 20692 35579
rect 17377 35555 17394 35556
rect 16661 35534 16689 35551
rect 16901 35534 16929 35551
rect 17058 35535 17109 35545
rect 17249 35544 17299 35555
rect 20665 35548 20692 35555
rect 18228 35545 18237 35547
rect 18288 35545 18320 35547
rect 18352 35545 18391 35547
rect 18487 35545 18527 35547
rect 19964 35545 20004 35547
rect 20100 35545 20139 35547
rect 20171 35545 20203 35547
rect 20254 35545 20263 35547
rect 17377 35536 17394 35537
rect 17122 35530 17141 35535
rect 14525 35511 14552 35518
rect 16661 35492 16689 35509
rect 16901 35492 16929 35509
rect 17027 35503 17058 35509
rect 17136 35503 17141 35530
rect 17217 35513 17249 35518
rect 17058 35493 17109 35503
rect 17249 35502 17299 35513
rect 14525 35461 14552 35468
rect 16710 35442 16738 35458
rect 16852 35442 16880 35458
rect 16987 35448 17037 35457
rect 17320 35451 17370 35462
rect 16956 35442 16987 35448
rect 17286 35445 17320 35451
rect 18209 35441 18214 35482
rect 18349 35470 18352 35520
rect 18391 35470 18394 35520
rect 18485 35470 18487 35520
rect 18527 35470 18529 35520
rect 19962 35470 19964 35520
rect 20004 35470 20006 35520
rect 20097 35470 20100 35520
rect 20139 35470 20142 35520
rect 20665 35506 20692 35513
rect 20277 35458 20282 35482
rect 20665 35466 20692 35473
rect 20301 35441 20306 35458
rect 14525 35419 14552 35426
rect 16764 35416 16769 35421
rect 16710 35400 16738 35416
rect 16852 35400 16880 35416
rect 16987 35406 17037 35415
rect 17204 35408 17221 35413
rect 17320 35409 17370 35420
rect 17377 35400 17394 35401
rect 16661 35379 16689 35396
rect 16901 35379 16929 35396
rect 17058 35380 17109 35390
rect 17249 35389 17299 35400
rect 18349 35391 18352 35441
rect 18391 35391 18394 35441
rect 18485 35391 18487 35441
rect 18527 35391 18529 35441
rect 19962 35391 19964 35441
rect 20004 35391 20006 35441
rect 20097 35391 20100 35441
rect 20139 35391 20142 35441
rect 20665 35424 20692 35431
rect 20665 35400 20692 35407
rect 17377 35381 17394 35382
rect 17122 35375 17141 35380
rect 14517 35355 14556 35358
rect 16661 35337 16689 35354
rect 16901 35337 16929 35354
rect 17027 35348 17058 35354
rect 17136 35348 17141 35375
rect 17217 35358 17249 35363
rect 20665 35358 20692 35365
rect 17058 35338 17109 35348
rect 17249 35347 17299 35358
rect 23423 35348 23463 35359
rect 23573 35348 23613 35359
rect 20665 35318 20692 35325
rect 14517 35313 14556 35316
rect 23423 35306 23463 35317
rect 23573 35306 23613 35317
rect 16661 35287 16689 35304
rect 16901 35287 16929 35304
rect 17058 35293 17109 35303
rect 17027 35287 17058 35293
rect 17136 35266 17141 35293
rect 17249 35283 17299 35294
rect 17217 35278 17249 35283
rect 17574 35268 17624 35279
rect 17754 35268 17804 35279
rect 17894 35268 17944 35278
rect 14517 35259 14556 35262
rect 16661 35245 16689 35262
rect 16788 35244 16793 35249
rect 16901 35245 16929 35262
rect 17122 35261 17141 35266
rect 17058 35251 17109 35261
rect 17377 35259 17394 35260
rect 17217 35252 17245 35257
rect 17990 35256 18007 35258
rect 17249 35241 17299 35252
rect 16710 35225 16738 35241
rect 16852 35225 16880 35241
rect 17377 35240 17394 35241
rect 17804 35237 17834 35241
rect 16987 35226 17037 35235
rect 17320 35221 17370 35232
rect 17574 35226 17624 35237
rect 17754 35226 17804 35237
rect 17864 35236 17869 35241
rect 17990 35237 18007 35239
rect 17894 35226 17944 35236
rect 17990 35222 18007 35224
rect 18209 35221 18214 35262
rect 18349 35238 18352 35288
rect 18391 35238 18394 35288
rect 18485 35238 18487 35288
rect 18527 35238 18529 35288
rect 19962 35238 19964 35288
rect 20004 35238 20006 35288
rect 20097 35238 20100 35288
rect 20139 35238 20142 35288
rect 23347 35287 23387 35297
rect 23573 35285 23613 35297
rect 20665 35276 20692 35283
rect 20277 35238 20282 35262
rect 20665 35252 20692 35259
rect 23347 35245 23387 35255
rect 23573 35243 23613 35255
rect 20301 35221 20306 35238
rect 14517 35217 14556 35220
rect 17574 35206 17624 35217
rect 17840 35206 17845 35217
rect 17894 35206 17944 35217
rect 20665 35210 20692 35217
rect 17864 35200 17869 35206
rect 17990 35203 18007 35205
rect 16710 35183 16738 35199
rect 16852 35183 16880 35199
rect 16956 35193 16987 35199
rect 16987 35184 17037 35193
rect 17286 35190 17320 35196
rect 17320 35179 17370 35190
rect 17546 35175 17574 35181
rect 17624 35175 17652 35181
rect 17864 35175 17894 35181
rect 14517 35163 14556 35166
rect 17574 35164 17624 35175
rect 17894 35164 17944 35175
rect 18349 35159 18352 35209
rect 18391 35159 18394 35209
rect 18485 35159 18487 35209
rect 18527 35159 18529 35209
rect 19962 35159 19964 35209
rect 20004 35159 20006 35209
rect 20097 35159 20100 35209
rect 20139 35159 20142 35209
rect 23347 35186 23387 35196
rect 23573 35186 23613 35198
rect 20665 35170 20692 35177
rect 16661 35132 16689 35149
rect 16901 35132 16929 35149
rect 17058 35138 17109 35148
rect 23347 35144 23387 35154
rect 23573 35144 23613 35156
rect 17027 35132 17058 35138
rect 14517 35121 14556 35124
rect 17136 35111 17141 35138
rect 17249 35128 17299 35139
rect 18228 35132 18237 35134
rect 18288 35132 18320 35134
rect 18352 35132 18391 35134
rect 18487 35132 18527 35134
rect 19964 35132 20004 35134
rect 20100 35132 20139 35134
rect 20171 35132 20203 35134
rect 20254 35132 20263 35134
rect 20665 35128 20692 35135
rect 17217 35123 17249 35128
rect 17574 35115 17624 35126
rect 17894 35115 17944 35126
rect 23423 35124 23463 35135
rect 23573 35124 23613 35135
rect 16661 35090 16689 35107
rect 16788 35089 16793 35094
rect 16901 35090 16929 35107
rect 17122 35106 17141 35111
rect 17546 35109 17574 35115
rect 17624 35109 17652 35115
rect 17864 35109 17894 35115
rect 17058 35096 17109 35106
rect 17377 35104 17394 35105
rect 17217 35097 17245 35102
rect 17249 35086 17299 35097
rect 16710 35070 16738 35086
rect 16852 35070 16880 35086
rect 17377 35085 17394 35086
rect 17864 35084 17869 35109
rect 18164 35102 18214 35113
rect 18236 35102 18286 35113
rect 20205 35102 20255 35113
rect 20277 35102 20327 35113
rect 20665 35104 20692 35111
rect 18286 35101 18320 35102
rect 20171 35101 20205 35102
rect 20844 35098 20868 35103
rect 17990 35085 18007 35087
rect 16987 35071 17037 35080
rect 17320 35066 17370 35077
rect 17574 35073 17624 35084
rect 17840 35077 17845 35078
rect 17828 35073 17845 35077
rect 17894 35073 17944 35084
rect 23423 35082 23463 35093
rect 23573 35082 23613 35093
rect 17990 35066 18007 35068
rect 17574 35053 17624 35064
rect 17754 35053 17804 35064
rect 17894 35054 17944 35064
rect 18164 35060 18214 35071
rect 18236 35060 18286 35071
rect 20205 35060 20255 35071
rect 20277 35060 20327 35071
rect 20665 35062 20692 35069
rect 17990 35051 18007 35053
rect 23423 35046 23463 35057
rect 23573 35046 23613 35057
rect 16710 35028 16738 35044
rect 16852 35028 16880 35044
rect 16956 35038 16987 35044
rect 16987 35029 17037 35038
rect 17286 35035 17320 35041
rect 17320 35024 17370 35035
rect 17990 35032 18007 35034
rect 17574 35011 17624 35022
rect 17754 35011 17804 35022
rect 17894 35012 17944 35022
rect 18165 35005 18215 35016
rect 18237 35005 18287 35016
rect 20205 35005 20255 35016
rect 20277 35005 20327 35016
rect 20665 35011 20692 35018
rect 23423 35004 23463 35015
rect 23573 35004 23613 35015
rect 20868 34998 20885 35003
rect 16661 34977 16689 34994
rect 16901 34977 16929 34994
rect 17058 34983 17109 34993
rect 17027 34977 17058 34983
rect 17136 34956 17141 34983
rect 17249 34973 17299 34984
rect 17574 34975 17624 34986
rect 17754 34975 17804 34986
rect 23347 34985 23387 34995
rect 17894 34975 17944 34985
rect 23573 34983 23613 34995
rect 18287 34974 18321 34975
rect 20171 34974 20205 34975
rect 17217 34968 17249 34973
rect 17990 34963 18007 34965
rect 18165 34963 18215 34974
rect 18237 34963 18287 34974
rect 20205 34963 20255 34974
rect 20277 34963 20327 34974
rect 20665 34969 20692 34976
rect 16661 34935 16689 34952
rect 16788 34934 16793 34939
rect 16901 34935 16929 34952
rect 17122 34951 17141 34956
rect 17058 34941 17109 34951
rect 17377 34949 17394 34950
rect 17217 34942 17245 34947
rect 17804 34944 17834 34948
rect 17249 34931 17299 34942
rect 17574 34933 17624 34944
rect 17754 34933 17804 34944
rect 17864 34943 17869 34948
rect 17990 34944 18007 34946
rect 20665 34945 20692 34952
rect 17894 34933 17944 34943
rect 18229 34942 18238 34944
rect 18289 34942 18321 34944
rect 18353 34942 18392 34944
rect 18488 34942 18528 34944
rect 19964 34942 20004 34944
rect 20100 34942 20139 34944
rect 20171 34942 20203 34944
rect 20254 34942 20263 34944
rect 23347 34943 23387 34953
rect 18526 34934 18528 34942
rect 23573 34941 23613 34953
rect 16710 34915 16738 34931
rect 16852 34915 16880 34931
rect 17377 34930 17394 34931
rect 17990 34929 18007 34931
rect 16987 34916 17037 34925
rect 17320 34911 17370 34922
rect 17574 34913 17624 34924
rect 17840 34913 17845 34924
rect 17894 34913 17944 34924
rect 17864 34907 17869 34913
rect 17990 34910 18007 34912
rect 16710 34873 16738 34889
rect 16852 34873 16880 34889
rect 16956 34883 16987 34889
rect 16987 34874 17037 34883
rect 17286 34880 17320 34886
rect 17546 34882 17574 34888
rect 17624 34882 17652 34888
rect 17864 34882 17894 34888
rect 17320 34869 17370 34880
rect 17574 34871 17624 34882
rect 17894 34871 17944 34882
rect 16661 34822 16689 34839
rect 16901 34822 16929 34839
rect 18210 34838 18215 34879
rect 18350 34867 18353 34917
rect 18392 34867 18395 34917
rect 18486 34867 18488 34917
rect 18528 34867 18530 34917
rect 19962 34867 19964 34917
rect 20004 34867 20006 34917
rect 20097 34867 20100 34917
rect 20139 34867 20142 34917
rect 20665 34903 20692 34910
rect 23347 34884 23387 34894
rect 23573 34884 23613 34896
rect 20277 34855 20282 34879
rect 20665 34863 20692 34870
rect 20301 34838 20306 34855
rect 23347 34842 23387 34852
rect 23573 34842 23613 34854
rect 17058 34828 17109 34838
rect 17027 34822 17058 34828
rect 17136 34801 17141 34828
rect 17249 34818 17299 34829
rect 17574 34822 17624 34833
rect 17894 34822 17944 34833
rect 17217 34813 17249 34818
rect 17546 34816 17574 34822
rect 17624 34816 17652 34822
rect 17864 34816 17894 34822
rect 16661 34780 16689 34797
rect 16788 34779 16793 34784
rect 16901 34780 16929 34797
rect 17122 34796 17141 34801
rect 17058 34786 17109 34796
rect 17377 34794 17394 34795
rect 17217 34787 17245 34792
rect 17864 34791 17869 34816
rect 17990 34792 18007 34794
rect 17249 34776 17299 34787
rect 17574 34780 17624 34791
rect 17840 34784 17845 34785
rect 17828 34780 17845 34784
rect 17894 34780 17944 34791
rect 18350 34788 18353 34838
rect 18392 34788 18395 34838
rect 18486 34788 18488 34838
rect 18528 34788 18530 34838
rect 19962 34788 19964 34838
rect 20004 34788 20006 34838
rect 20097 34788 20100 34838
rect 20139 34788 20142 34838
rect 20665 34821 20692 34828
rect 23423 34822 23463 34833
rect 23573 34822 23613 34833
rect 20665 34797 20692 34804
rect 23423 34780 23463 34791
rect 23573 34780 23613 34791
rect 16710 34760 16738 34776
rect 16852 34760 16880 34776
rect 17377 34775 17394 34776
rect 17990 34773 18007 34775
rect 16987 34761 17037 34770
rect 17320 34756 17370 34767
rect 17574 34760 17624 34771
rect 17754 34760 17804 34771
rect 17894 34761 17944 34771
rect 17990 34758 18007 34760
rect 18948 34757 18965 34758
rect 19527 34757 19544 34758
rect 20665 34755 20692 34762
rect 17990 34739 18007 34741
rect 18948 34738 18965 34739
rect 19527 34738 19544 34739
rect 16710 34718 16738 34734
rect 16852 34718 16880 34734
rect 16956 34728 16987 34734
rect 16987 34719 17037 34728
rect 17286 34725 17320 34731
rect 17320 34714 17370 34725
rect 17574 34718 17624 34729
rect 17754 34718 17804 34729
rect 17894 34719 17944 34729
rect 18948 34722 18965 34724
rect 19527 34722 19544 34724
rect 20665 34715 20692 34722
rect 18949 34703 18966 34705
rect 19527 34703 19544 34705
rect 18210 34618 18215 34659
rect 18350 34635 18353 34685
rect 18392 34635 18395 34685
rect 18486 34635 18488 34685
rect 18528 34635 18530 34685
rect 19962 34635 19964 34685
rect 20004 34635 20006 34685
rect 20097 34635 20100 34685
rect 20139 34635 20142 34685
rect 20665 34673 20692 34680
rect 20277 34635 20282 34659
rect 20665 34649 20692 34656
rect 20301 34618 20306 34635
rect 20665 34607 20692 34614
rect 18350 34556 18353 34606
rect 18392 34556 18395 34606
rect 18486 34556 18488 34606
rect 18528 34556 18530 34606
rect 19962 34556 19964 34606
rect 20004 34556 20006 34606
rect 20097 34556 20100 34606
rect 20139 34556 20142 34606
rect 20665 34567 20692 34574
rect 18229 34529 18238 34531
rect 18289 34529 18321 34531
rect 18353 34529 18392 34531
rect 18488 34529 18528 34531
rect 19964 34529 20004 34531
rect 20100 34529 20139 34531
rect 20171 34529 20203 34531
rect 20254 34529 20263 34531
rect 20665 34525 20692 34532
rect 18165 34499 18215 34510
rect 18237 34499 18287 34510
rect 20205 34499 20255 34510
rect 20277 34499 20327 34510
rect 20665 34501 20692 34508
rect 18287 34498 18321 34499
rect 20171 34498 20205 34499
rect 20844 34495 20868 34500
rect 18165 34457 18215 34468
rect 18237 34457 18287 34468
rect 20205 34457 20255 34468
rect 20277 34457 20327 34468
rect 20665 34459 20692 34466
rect 16661 34274 16689 34291
rect 16901 34274 16929 34291
rect 17058 34280 17109 34290
rect 17027 34274 17058 34280
rect 17136 34253 17141 34280
rect 17249 34270 17299 34281
rect 17217 34265 17249 34270
rect 17574 34261 17624 34272
rect 17754 34261 17804 34272
rect 17894 34261 17944 34271
rect 18309 34270 18359 34281
rect 18381 34270 18431 34281
rect 20065 34270 20115 34281
rect 20137 34270 20187 34281
rect 16661 34232 16689 34249
rect 16788 34231 16793 34236
rect 16901 34232 16929 34249
rect 17122 34248 17141 34253
rect 17990 34249 18007 34251
rect 17058 34238 17109 34248
rect 17377 34246 17394 34247
rect 17217 34239 17245 34244
rect 18431 34239 18463 34240
rect 20033 34239 20065 34240
rect 17249 34228 17299 34239
rect 17804 34230 17834 34234
rect 16710 34212 16738 34228
rect 16852 34212 16880 34228
rect 17377 34227 17394 34228
rect 16987 34213 17037 34222
rect 17574 34219 17624 34230
rect 17754 34219 17804 34230
rect 17864 34229 17869 34234
rect 17990 34230 18007 34232
rect 17894 34219 17944 34229
rect 18309 34228 18359 34239
rect 18381 34228 18431 34239
rect 20065 34228 20115 34239
rect 20137 34228 20187 34239
rect 17320 34208 17370 34219
rect 17990 34215 18007 34217
rect 17574 34199 17624 34210
rect 17840 34199 17845 34210
rect 17894 34199 17944 34210
rect 18381 34208 18431 34220
rect 20065 34208 20115 34220
rect 17864 34193 17869 34199
rect 17990 34196 18007 34198
rect 16710 34170 16738 34186
rect 16852 34170 16880 34186
rect 16956 34180 16987 34186
rect 16987 34171 17037 34180
rect 17286 34177 17320 34183
rect 18350 34178 18354 34208
rect 18431 34207 18460 34208
rect 20036 34207 20065 34208
rect 20142 34178 20146 34208
rect 17320 34166 17370 34177
rect 17546 34168 17574 34174
rect 17624 34168 17652 34174
rect 17864 34168 17894 34174
rect 17574 34157 17624 34168
rect 17894 34157 17944 34168
rect 18381 34166 18431 34178
rect 20065 34166 20115 34178
rect 18556 34162 18573 34164
rect 18950 34163 18967 34165
rect 19529 34163 19546 34165
rect 19923 34162 19940 34164
rect 18556 34143 18573 34145
rect 18950 34144 18967 34146
rect 19529 34144 19546 34146
rect 19923 34143 19940 34145
rect 16661 34119 16689 34136
rect 16901 34119 16929 34136
rect 17058 34125 17109 34135
rect 18381 34126 18431 34138
rect 20065 34126 20115 34138
rect 17027 34119 17058 34125
rect 17136 34098 17141 34125
rect 17249 34115 17299 34126
rect 17217 34110 17249 34115
rect 17574 34108 17624 34119
rect 17894 34108 17944 34119
rect 17546 34102 17574 34108
rect 17624 34102 17652 34108
rect 17864 34102 17894 34108
rect 16661 34077 16689 34094
rect 16788 34076 16793 34081
rect 16901 34077 16929 34094
rect 17122 34093 17141 34098
rect 17058 34083 17109 34093
rect 17377 34091 17394 34092
rect 17217 34084 17245 34089
rect 17249 34073 17299 34084
rect 17864 34077 17869 34102
rect 18350 34096 18354 34126
rect 18431 34096 18460 34097
rect 20036 34096 20065 34097
rect 20142 34096 20146 34126
rect 18381 34084 18431 34096
rect 20065 34084 20115 34096
rect 17990 34078 18007 34080
rect 16710 34057 16738 34073
rect 16852 34057 16880 34073
rect 17377 34072 17394 34073
rect 16987 34058 17037 34067
rect 17574 34066 17624 34077
rect 17840 34070 17845 34071
rect 17828 34066 17845 34070
rect 17894 34066 17944 34077
rect 18309 34065 18359 34076
rect 18381 34065 18431 34076
rect 20065 34065 20115 34076
rect 20137 34065 20187 34076
rect 18431 34064 18463 34065
rect 20033 34064 20065 34065
rect 17320 34053 17370 34064
rect 17990 34059 18007 34061
rect 17574 34046 17624 34057
rect 17754 34046 17804 34057
rect 17894 34047 17944 34057
rect 17990 34044 18007 34046
rect 16710 34015 16738 34031
rect 16852 34015 16880 34031
rect 16956 34025 16987 34031
rect 16987 34016 17037 34025
rect 17286 34022 17320 34028
rect 17990 34025 18007 34027
rect 18309 34023 18359 34034
rect 18381 34023 18431 34034
rect 20065 34023 20115 34034
rect 20137 34023 20187 34034
rect 17320 34011 17370 34022
rect 18949 34017 18966 34019
rect 19530 34017 19547 34019
rect 17574 34004 17624 34015
rect 17754 34004 17804 34015
rect 17894 34005 17944 34015
rect 18556 34003 18573 34005
rect 19923 34003 19940 34005
rect 18949 33998 18966 34000
rect 19530 33998 19547 34000
rect 18556 33984 18573 33986
rect 19923 33984 19940 33986
rect 16661 33964 16689 33981
rect 16901 33964 16929 33981
rect 17058 33970 17109 33980
rect 17027 33964 17058 33970
rect 17136 33943 17141 33970
rect 17249 33960 17299 33971
rect 17574 33968 17624 33979
rect 17754 33968 17804 33979
rect 17894 33968 17944 33978
rect 18309 33969 18359 33980
rect 18381 33969 18431 33980
rect 20065 33969 20115 33980
rect 20137 33969 20187 33980
rect 17217 33955 17249 33960
rect 17990 33956 18007 33958
rect 16661 33922 16689 33939
rect 16788 33921 16793 33926
rect 16901 33922 16929 33939
rect 17122 33938 17141 33943
rect 17058 33928 17109 33938
rect 17804 33937 17834 33941
rect 17377 33936 17394 33937
rect 17217 33929 17245 33934
rect 17249 33918 17299 33929
rect 17574 33926 17624 33937
rect 17754 33926 17804 33937
rect 17864 33936 17869 33941
rect 17990 33937 18007 33939
rect 18431 33938 18463 33939
rect 20033 33938 20065 33939
rect 17894 33926 17944 33936
rect 18309 33927 18359 33938
rect 18381 33927 18431 33938
rect 20065 33927 20115 33938
rect 20137 33927 20187 33938
rect 17990 33922 18007 33924
rect 16710 33902 16738 33918
rect 16852 33902 16880 33918
rect 17377 33917 17394 33918
rect 16987 33903 17037 33912
rect 17320 33898 17370 33909
rect 17574 33906 17624 33917
rect 17840 33906 17845 33917
rect 17894 33906 17944 33917
rect 18381 33907 18431 33919
rect 20065 33907 20115 33919
rect 17864 33900 17869 33906
rect 17990 33903 18007 33905
rect 16710 33860 16738 33876
rect 16852 33860 16880 33876
rect 16956 33870 16987 33876
rect 17546 33875 17574 33881
rect 17624 33875 17652 33881
rect 17864 33875 17894 33881
rect 18350 33877 18354 33907
rect 18431 33906 18460 33907
rect 20036 33906 20065 33907
rect 20142 33877 20146 33907
rect 16987 33861 17037 33870
rect 17286 33867 17320 33873
rect 17320 33856 17370 33867
rect 17574 33864 17624 33875
rect 17894 33864 17944 33875
rect 18381 33865 18431 33877
rect 20065 33865 20115 33877
rect 18381 33826 18431 33838
rect 20065 33826 20115 33838
rect 16661 33809 16689 33826
rect 16901 33809 16929 33826
rect 17058 33815 17109 33825
rect 17027 33809 17058 33815
rect 17136 33788 17141 33815
rect 17249 33805 17299 33816
rect 17574 33815 17624 33826
rect 17894 33815 17944 33826
rect 17546 33809 17574 33815
rect 17624 33809 17652 33815
rect 17864 33809 17894 33815
rect 17217 33800 17249 33805
rect 16661 33767 16689 33784
rect 16788 33766 16793 33771
rect 16901 33767 16929 33784
rect 17122 33783 17141 33788
rect 17864 33784 17869 33809
rect 18350 33796 18354 33826
rect 18431 33796 18460 33797
rect 20036 33796 20065 33797
rect 20142 33796 20146 33826
rect 17990 33785 18007 33787
rect 18381 33784 18431 33796
rect 20065 33784 20115 33796
rect 17058 33773 17109 33783
rect 17377 33781 17394 33782
rect 17217 33774 17245 33779
rect 17249 33763 17299 33774
rect 17574 33773 17624 33784
rect 17840 33777 17845 33778
rect 17828 33773 17845 33777
rect 17894 33773 17944 33784
rect 17990 33766 18007 33768
rect 18309 33765 18359 33776
rect 18381 33765 18431 33776
rect 20065 33765 20115 33776
rect 20137 33765 20187 33776
rect 18431 33764 18463 33765
rect 20033 33764 20065 33765
rect 16710 33747 16738 33763
rect 16852 33747 16880 33763
rect 17377 33762 17394 33763
rect 16987 33748 17037 33757
rect 17320 33743 17370 33754
rect 17574 33753 17624 33764
rect 17754 33753 17804 33764
rect 17894 33754 17944 33764
rect 17990 33751 18007 33753
rect 17990 33732 18007 33734
rect 18309 33723 18359 33734
rect 18381 33723 18431 33734
rect 20065 33723 20115 33734
rect 20137 33723 20187 33734
rect 16710 33705 16738 33721
rect 16852 33705 16880 33721
rect 16956 33715 16987 33721
rect 16987 33706 17037 33715
rect 17286 33712 17320 33718
rect 17320 33701 17370 33712
rect 17574 33711 17624 33722
rect 17754 33711 17804 33722
rect 17894 33712 17944 33722
rect 16661 33297 16689 33314
rect 16901 33297 16929 33314
rect 17058 33303 17109 33313
rect 17027 33297 17058 33303
rect 17136 33276 17141 33303
rect 17249 33293 17299 33304
rect 17217 33288 17249 33293
rect 17574 33285 17624 33296
rect 17754 33285 17804 33296
rect 17894 33285 17944 33295
rect 18309 33292 18359 33303
rect 18381 33292 18431 33303
rect 16661 33255 16689 33272
rect 16788 33254 16793 33259
rect 16901 33255 16929 33272
rect 17122 33271 17141 33276
rect 17990 33273 18007 33275
rect 17058 33261 17109 33271
rect 17377 33269 17394 33270
rect 17217 33262 17245 33267
rect 17249 33251 17299 33262
rect 18431 33261 18463 33262
rect 17804 33254 17834 33258
rect 16710 33235 16738 33251
rect 16852 33235 16880 33251
rect 17377 33250 17394 33251
rect 16987 33236 17037 33245
rect 17574 33243 17624 33254
rect 17754 33243 17804 33254
rect 17864 33253 17869 33258
rect 17990 33254 18007 33256
rect 17894 33243 17944 33253
rect 18309 33250 18359 33261
rect 18381 33250 18431 33261
rect 17320 33231 17370 33242
rect 17990 33239 18007 33241
rect 17574 33223 17624 33234
rect 17840 33223 17845 33234
rect 17894 33223 17944 33234
rect 18381 33230 18431 33242
rect 17864 33217 17869 33223
rect 17990 33220 18007 33222
rect 16710 33193 16738 33209
rect 16852 33193 16880 33209
rect 16956 33203 16987 33209
rect 16987 33194 17037 33203
rect 17286 33200 17320 33206
rect 18350 33200 18354 33230
rect 18431 33229 18460 33230
rect 17320 33189 17370 33200
rect 17546 33192 17574 33198
rect 17624 33192 17652 33198
rect 17864 33192 17894 33198
rect 17574 33181 17624 33192
rect 17894 33181 17944 33192
rect 18381 33188 18431 33200
rect 18971 33185 18988 33187
rect 18569 33182 18586 33184
rect 18971 33166 18988 33168
rect 18569 33163 18586 33165
rect 16661 33142 16689 33159
rect 16901 33142 16929 33159
rect 17058 33148 17109 33158
rect 17027 33142 17058 33148
rect 17136 33121 17141 33148
rect 17249 33138 17299 33149
rect 18381 33148 18431 33160
rect 17217 33133 17249 33138
rect 17574 33132 17624 33143
rect 17894 33132 17944 33143
rect 17546 33126 17574 33132
rect 17624 33126 17652 33132
rect 17864 33126 17894 33132
rect 16661 33100 16689 33117
rect 16788 33099 16793 33104
rect 16901 33100 16929 33117
rect 17122 33116 17141 33121
rect 17058 33106 17109 33116
rect 17377 33114 17394 33115
rect 17217 33107 17245 33112
rect 17249 33096 17299 33107
rect 17864 33101 17869 33126
rect 18350 33118 18354 33148
rect 18431 33118 18460 33119
rect 18381 33106 18431 33118
rect 17990 33102 18007 33104
rect 16710 33080 16738 33096
rect 16852 33080 16880 33096
rect 17377 33095 17394 33096
rect 17574 33090 17624 33101
rect 17840 33094 17845 33095
rect 17828 33090 17845 33094
rect 17894 33090 17944 33101
rect 16987 33081 17037 33090
rect 18309 33087 18359 33098
rect 18381 33087 18431 33098
rect 17320 33076 17370 33087
rect 18431 33086 18463 33087
rect 17990 33083 18007 33085
rect 17574 33070 17624 33081
rect 17754 33070 17804 33081
rect 17894 33071 17944 33081
rect 17990 33068 18007 33070
rect 18568 33064 18585 33066
rect 18970 33058 18987 33060
rect 16710 33038 16738 33054
rect 16852 33038 16880 33054
rect 16956 33048 16987 33054
rect 16987 33039 17037 33048
rect 17286 33045 17320 33051
rect 17990 33049 18007 33051
rect 18309 33045 18359 33056
rect 18381 33045 18431 33056
rect 18568 33045 18585 33047
rect 17320 33034 17370 33045
rect 18970 33039 18987 33041
rect 17574 33028 17624 33039
rect 17754 33028 17804 33039
rect 17894 33029 17944 33039
rect 18568 33030 18585 33032
rect 18970 33024 18987 33026
rect 18568 33011 18585 33013
rect 18970 33005 18987 33007
rect 16661 32987 16689 33004
rect 16901 32987 16929 33004
rect 17058 32993 17109 33003
rect 17027 32987 17058 32993
rect 17136 32966 17141 32993
rect 17249 32983 17299 32994
rect 17574 32992 17624 33003
rect 17754 32992 17804 33003
rect 17894 32992 17944 33002
rect 18309 32991 18359 33002
rect 18381 32991 18431 33002
rect 18568 32996 18585 32998
rect 18970 32990 18987 32992
rect 17217 32978 17249 32983
rect 17990 32980 18007 32982
rect 18568 32977 18585 32979
rect 18970 32971 18987 32973
rect 16661 32945 16689 32962
rect 16788 32944 16793 32949
rect 16901 32945 16929 32962
rect 17122 32961 17141 32966
rect 17804 32961 17834 32965
rect 17058 32951 17109 32961
rect 17377 32959 17394 32960
rect 17217 32952 17245 32957
rect 17249 32941 17299 32952
rect 17574 32950 17624 32961
rect 17754 32950 17804 32961
rect 17864 32960 17869 32965
rect 17990 32961 18007 32963
rect 18431 32960 18463 32961
rect 17894 32950 17944 32960
rect 18309 32949 18359 32960
rect 18381 32949 18431 32960
rect 18970 32956 18987 32958
rect 17990 32946 18007 32948
rect 16710 32925 16738 32941
rect 16852 32925 16880 32941
rect 17377 32940 17394 32941
rect 16987 32926 17037 32935
rect 17320 32921 17370 32932
rect 17574 32930 17624 32941
rect 17840 32930 17845 32941
rect 17894 32930 17944 32941
rect 17864 32924 17869 32930
rect 18381 32929 18431 32941
rect 17990 32927 18007 32929
rect 17546 32899 17574 32905
rect 17624 32899 17652 32905
rect 17864 32899 17894 32905
rect 18350 32899 18354 32929
rect 18431 32928 18460 32929
rect 16710 32883 16738 32899
rect 16852 32883 16880 32899
rect 16956 32893 16987 32899
rect 16987 32884 17037 32893
rect 17286 32890 17320 32896
rect 17320 32879 17370 32890
rect 17574 32888 17624 32899
rect 17894 32888 17944 32899
rect 18381 32887 18431 32899
rect 16661 32832 16689 32849
rect 16901 32832 16929 32849
rect 17058 32838 17109 32848
rect 17574 32839 17624 32850
rect 17894 32839 17944 32850
rect 18381 32848 18431 32860
rect 17027 32832 17058 32838
rect 17136 32811 17141 32838
rect 17249 32828 17299 32839
rect 17546 32833 17574 32839
rect 17624 32833 17652 32839
rect 17864 32833 17894 32839
rect 17217 32823 17249 32828
rect 16661 32790 16689 32807
rect 16788 32789 16793 32794
rect 16901 32790 16929 32807
rect 17122 32806 17141 32811
rect 17864 32808 17869 32833
rect 18350 32818 18354 32848
rect 18431 32818 18460 32819
rect 17990 32809 18007 32811
rect 17058 32796 17109 32806
rect 17377 32804 17394 32805
rect 17217 32797 17245 32802
rect 17574 32797 17624 32808
rect 17840 32801 17845 32802
rect 17828 32797 17845 32801
rect 17894 32797 17944 32808
rect 18381 32806 18431 32818
rect 17249 32786 17299 32797
rect 17990 32790 18007 32792
rect 16710 32770 16738 32786
rect 16852 32770 16880 32786
rect 17377 32785 17394 32786
rect 16987 32771 17037 32780
rect 17574 32777 17624 32788
rect 17754 32777 17804 32788
rect 17894 32778 17944 32788
rect 18309 32787 18359 32798
rect 18381 32787 18431 32798
rect 18431 32786 18463 32787
rect 17320 32766 17370 32777
rect 17990 32775 18007 32777
rect 17990 32756 18007 32758
rect 16710 32728 16738 32744
rect 16852 32728 16880 32744
rect 16956 32738 16987 32744
rect 16987 32729 17037 32738
rect 17286 32735 17320 32741
rect 17574 32735 17624 32746
rect 17754 32735 17804 32746
rect 17894 32736 17944 32746
rect 18309 32745 18359 32756
rect 18381 32745 18431 32756
rect 17320 32724 17370 32735
rect 22937 31860 22940 31899
rect 22979 31860 22982 31899
rect 23033 31860 23036 31899
rect 23075 31860 23078 31899
rect 23129 31860 23132 31899
rect 23171 31860 23174 31899
rect 23225 31860 23228 31899
rect 23267 31860 23270 31899
rect 23321 31860 23324 31899
rect 23363 31860 23366 31899
rect 23417 31860 23420 31899
rect 23459 31860 23462 31899
rect 22937 31699 22940 31738
rect 22979 31699 22982 31738
rect 23033 31698 23036 31737
rect 23075 31698 23078 31737
rect 23129 31698 23132 31737
rect 23171 31698 23174 31737
rect 23225 31698 23228 31737
rect 23267 31698 23270 31737
rect 23321 31698 23324 31737
rect 23363 31698 23366 31737
rect 23417 31699 23420 31738
rect 23459 31699 23462 31738
rect 22937 31538 22940 31577
rect 22979 31538 22982 31577
rect 23033 31537 23036 31576
rect 23075 31537 23078 31576
rect 23129 31537 23132 31576
rect 23171 31537 23174 31576
rect 23225 31537 23228 31576
rect 23267 31537 23270 31576
rect 23321 31537 23324 31576
rect 23363 31537 23366 31576
rect 23417 31538 23420 31577
rect 23459 31538 23462 31577
rect 23509 31471 23513 31503
rect 23523 31457 23527 31517
rect 22937 31377 22940 31416
rect 22979 31377 22982 31416
rect 23033 31376 23036 31415
rect 23075 31376 23078 31415
rect 23129 31376 23132 31415
rect 23171 31376 23174 31415
rect 23225 31376 23228 31415
rect 23267 31376 23270 31415
rect 23321 31376 23324 31415
rect 23363 31376 23366 31415
rect 23417 31377 23420 31416
rect 23459 31377 23462 31416
rect 23039 31349 23075 31354
rect 23509 31310 23513 31342
rect 23523 31296 23527 31356
rect 22937 31216 22940 31255
rect 22979 31216 22982 31255
rect 23033 31215 23036 31254
rect 23075 31215 23078 31254
rect 23129 31215 23132 31254
rect 23171 31215 23174 31254
rect 23225 31215 23228 31254
rect 23267 31215 23270 31254
rect 23321 31215 23324 31254
rect 23363 31215 23366 31254
rect 23417 31216 23420 31255
rect 23459 31216 23462 31255
rect 23205 31165 23209 31166
rect 23508 31149 23512 31181
rect 23522 31135 23526 31195
rect 22937 31055 22940 31094
rect 22979 31055 22982 31094
rect 23033 31054 23036 31093
rect 23075 31054 23078 31093
rect 23129 31054 23132 31093
rect 23171 31054 23174 31093
rect 23225 31054 23228 31093
rect 23267 31054 23270 31093
rect 23321 31054 23324 31093
rect 23363 31054 23366 31093
rect 23417 31055 23420 31094
rect 23459 31055 23462 31094
rect 23508 30987 23513 31019
rect 23522 30973 23527 31033
rect 22937 30894 22940 30933
rect 22979 30894 22982 30933
rect 23033 30893 23036 30932
rect 23075 30893 23078 30932
rect 23129 30893 23132 30932
rect 23171 30893 23174 30932
rect 23225 30893 23228 30932
rect 23267 30893 23270 30932
rect 23321 30893 23324 30932
rect 23363 30893 23366 30932
rect 23417 30894 23420 30933
rect 23459 30894 23462 30933
rect 23508 30826 23512 30858
rect 23522 30812 23526 30872
rect 22937 30733 22940 30772
rect 22979 30733 22982 30772
rect 23033 30732 23036 30771
rect 23075 30732 23078 30771
rect 23129 30732 23132 30771
rect 23171 30732 23174 30771
rect 23225 30732 23228 30771
rect 23267 30732 23270 30771
rect 23321 30732 23324 30771
rect 23363 30732 23366 30771
rect 23417 30733 23420 30772
rect 23459 30733 23462 30772
rect 22937 30572 22940 30611
rect 22979 30572 22982 30611
rect 23033 30571 23036 30610
rect 23075 30571 23078 30610
rect 23129 30571 23132 30610
rect 23171 30571 23174 30610
rect 23225 30571 23228 30610
rect 23267 30571 23270 30610
rect 23321 30571 23324 30610
rect 23363 30571 23366 30610
rect 23417 30572 23420 30611
rect 23459 30572 23462 30611
rect 23509 30506 23512 30538
rect 23523 30492 23526 30552
rect 22937 30411 22940 30450
rect 22979 30411 22982 30450
rect 23033 30411 23036 30450
rect 23075 30411 23078 30450
rect 23129 30411 23132 30450
rect 23171 30411 23174 30450
rect 23225 30411 23228 30450
rect 23267 30411 23270 30450
rect 23321 30411 23324 30450
rect 23363 30411 23366 30450
rect 23417 30411 23420 30450
rect 23459 30411 23462 30450
<< metal1 >>
rect 2362 38791 2751 38908
rect 5221 38790 5610 38907
rect 8080 38790 8469 38907
rect 12270 38793 12659 38910
rect 16482 38791 16871 38908
rect 19341 38791 19730 38908
rect 22201 38791 22590 38908
rect 25060 38791 25449 38908
rect 27919 38791 28308 38908
rect 30778 38790 31167 38907
rect 33637 38790 34026 38907
rect 2914 36559 3237 37870
rect 5773 36900 6096 37870
rect 8632 37329 8955 37870
rect 9886 37649 9903 37661
rect 8589 37298 8972 37329
rect 8589 37073 8632 37298
rect 8955 37073 8972 37298
rect 8589 37055 8972 37073
rect 9851 36993 9903 37649
rect 9845 36982 9910 36993
rect 9845 36945 9851 36982
rect 9903 36945 9910 36982
rect 9845 36942 9910 36945
rect 5757 36849 6107 36900
rect 5757 36624 5773 36849
rect 6096 36624 6107 36849
rect 5757 36611 6107 36624
rect 2697 36520 3237 36559
rect 2697 36197 2731 36520
rect 2956 36197 3237 36520
rect 1453 36189 1792 36196
rect 1356 36180 1792 36189
rect 1033 35857 1578 36180
rect 1764 35857 1792 36180
rect 2697 36179 2991 36197
rect 9851 36174 9903 36942
rect 10191 36551 10232 37672
rect 12902 37472 13018 37663
rect 12902 37359 15638 37472
rect 12902 37339 15657 37359
rect 15505 37199 15638 37339
rect 17034 37248 17357 37871
rect 18198 37663 18259 37677
rect 18196 37467 18314 37663
rect 18116 37376 18314 37467
rect 18116 37358 18297 37376
rect 18640 37360 18712 37746
rect 18116 37289 18189 37358
rect 19893 37248 20216 37870
rect 22752 37248 23075 37870
rect 23645 37609 23664 37610
rect 24358 37609 24430 37746
rect 23645 37574 24430 37609
rect 23645 37361 23664 37574
rect 25611 37555 25934 37870
rect 25535 37527 25934 37555
rect 25533 37507 25934 37527
rect 25515 37410 25950 37507
rect 25515 37204 25611 37410
rect 25934 37204 25950 37410
rect 25515 37137 25950 37204
rect 28470 37089 28793 37870
rect 28440 37045 28795 37089
rect 28440 36715 28470 37045
rect 28676 36715 28795 37045
rect 28440 36684 28795 36715
rect 10179 36548 10232 36551
rect 10179 36507 10185 36548
rect 10226 36507 10232 36548
rect 31329 36526 31652 37870
rect 10179 36504 10232 36507
rect 9831 36165 9903 36174
rect 9831 36113 9837 36165
rect 9889 36113 9903 36165
rect 9831 36101 9903 36113
rect 1356 35789 1792 35857
rect 0 35305 125 35694
rect 2370 33321 2596 33325
rect 1033 32998 2383 33321
rect 2591 32998 2596 33321
rect 2370 32994 2596 32998
rect 1 32447 126 32836
rect 9851 32566 9903 36101
rect 10191 36079 10232 36504
rect 31309 36496 31668 36526
rect 31309 36290 31329 36496
rect 31652 36290 31668 36496
rect 31309 36273 31668 36290
rect 34188 36177 34511 37870
rect 10177 36069 10239 36079
rect 10177 36028 10190 36069
rect 10231 36028 10239 36069
rect 10177 36020 10239 36028
rect 34157 36054 34533 36177
rect 9843 32563 9906 32566
rect 9843 32511 9847 32563
rect 9899 32511 9906 32563
rect 9843 32506 9906 32511
rect 10191 32464 10232 36020
rect 34157 35849 34188 36054
rect 34511 35849 34533 36054
rect 34157 35815 34533 35849
rect 35592 36108 35933 36140
rect 35592 35785 35622 36108
rect 35821 35785 36256 36108
rect 26424 35719 26866 35780
rect 35592 35736 35933 35785
rect 26424 35687 26448 35719
rect 26670 35687 26866 35719
rect 26424 32769 26866 35687
rect 37160 35235 37285 35624
rect 34751 33249 34983 33257
rect 34751 32926 34767 33249
rect 34976 32926 36255 33249
rect 34751 32920 34983 32926
rect 26421 32757 26868 32769
rect 26421 32648 26432 32757
rect 26860 32648 26868 32757
rect 26421 32637 26868 32648
rect 10186 32461 10234 32464
rect 10186 32417 10190 32461
rect 10231 32417 10234 32461
rect 10186 32414 10234 32417
rect 2761 30462 2984 30470
rect 1034 30139 2773 30462
rect 2981 30139 2984 30462
rect 2761 30124 2984 30139
rect 0 29587 125 29976
rect 3212 27603 3453 27613
rect 1033 27280 3236 27603
rect 3444 27280 3453 27603
rect 3212 27270 3453 27280
rect 2 26728 127 27117
rect 3668 24744 3895 24751
rect 1034 24421 3677 24744
rect 3885 24421 3895 24744
rect 3668 24411 3895 24421
rect 1 23870 126 24259
rect 4104 21885 4329 21891
rect 1033 21562 4111 21885
rect 4319 21562 4329 21885
rect 4104 21554 4329 21562
rect 0 21010 125 21399
rect 4536 19026 4761 19037
rect 1033 18703 4776 19026
rect 4536 18692 4761 18703
rect 1 18152 126 18541
rect 26424 16507 26866 32637
rect 37159 32375 37284 32764
rect 34334 30390 34570 30403
rect 34334 30067 34342 30390
rect 34551 30067 36257 30390
rect 34334 30057 34570 30067
rect 37159 29515 37284 29904
rect 33933 27531 34161 27547
rect 33933 27208 33944 27531
rect 34153 27208 36255 27531
rect 33933 27197 34161 27208
rect 37160 26659 37285 27048
rect 33503 24672 33745 24684
rect 33503 24349 33519 24672
rect 33728 24349 36255 24672
rect 33503 24333 33745 24349
rect 37158 23798 37283 24187
rect 33114 21813 33341 21824
rect 33114 21490 33125 21813
rect 33334 21490 36256 21813
rect 33114 21477 33341 21490
rect 37160 20940 37285 21329
rect 32674 18954 32904 18962
rect 32674 18631 36256 18954
rect 32674 18621 32904 18631
rect 37160 18079 37285 18468
rect 26332 16496 26866 16507
rect 4942 16167 5183 16177
rect 1033 15844 4965 16167
rect 5173 15844 5183 16167
rect 26332 16054 26350 16496
rect 26792 16133 26866 16496
rect 26792 16054 26808 16133
rect 26332 16037 26808 16054
rect 4942 15826 5183 15844
rect 4 15294 129 15683
rect 5370 13308 5616 13315
rect 1033 12985 5616 13308
rect 5370 12980 5616 12985
rect 2 12433 127 12822
rect 5807 10449 6047 10463
rect 1032 10126 5827 10449
rect 6035 10126 6047 10449
rect 5807 10116 6047 10126
rect 1 9574 126 9963
rect 6201 7590 6450 7598
rect 1032 7267 6224 7590
rect 6432 7267 6450 7590
rect 6201 7248 6450 7267
rect 1 6715 126 7104
rect 6648 4731 6883 4741
rect 1034 4408 6668 4731
rect 6876 4408 6883 4731
rect 6648 4395 6883 4408
rect 2 3856 127 4245
rect 7048 1872 7319 1878
rect 1034 1549 7098 1872
rect 7306 1549 7319 1872
rect 7048 1537 7319 1549
rect 2 998 127 1387
<< via1 >>
rect 8632 37073 8955 37298
rect 9851 36945 9903 36982
rect 5773 36624 6096 36849
rect 2731 36197 2956 36520
rect 1578 35857 1764 36180
rect 25611 37204 25934 37410
rect 28470 36715 28676 37045
rect 10185 36507 10226 36548
rect 9837 36113 9889 36165
rect 2383 32998 2591 33321
rect 31329 36290 31652 36496
rect 10190 36028 10231 36069
rect 9847 32511 9899 32563
rect 34188 35849 34511 36054
rect 35622 35785 35821 36108
rect 26448 35687 26670 35719
rect 34767 32926 34976 33249
rect 26432 32648 26860 32757
rect 10190 32417 10231 32461
rect 2773 30139 2981 30462
rect 3236 27280 3444 27603
rect 3677 24421 3885 24744
rect 4111 21562 4319 21885
rect 34342 30067 34551 30390
rect 33944 27208 34153 27531
rect 33519 24349 33728 24672
rect 33125 21490 33334 21813
rect 4965 15844 5173 16167
rect 26350 16054 26792 16496
rect 5827 10126 6035 10449
rect 6224 7267 6432 7590
rect 6668 4408 6876 4731
rect 7098 1549 7306 1872
<< metal2 >>
rect 36849 38502 36968 38503
rect 342 38501 1635 38502
rect 329 38362 1635 38501
rect 35669 38450 36968 38502
rect 35648 38374 36968 38450
rect 329 38210 558 38362
rect 374 38206 558 38210
rect 418 37354 558 38206
rect 36752 38242 36968 38374
rect 1045 37725 1620 37865
rect 35584 37732 36251 37872
rect 1045 37253 1185 37725
rect 25496 37410 25976 37490
rect 8576 37324 8985 37349
rect 8576 37298 12773 37324
rect 8576 37073 8632 37298
rect 8955 37099 12773 37298
rect 25496 37281 25611 37410
rect 24326 37204 25611 37281
rect 25934 37281 25976 37410
rect 25934 37204 25981 37281
rect 8955 37073 8985 37099
rect 24326 37075 25981 37204
rect 36110 37181 36250 37732
rect 36752 37319 36880 38242
rect 36804 37245 36880 37319
rect 8576 37039 8985 37073
rect 28455 37045 28786 37074
rect 9846 36988 9908 36990
rect 9846 36982 12761 36988
rect 9846 36945 9851 36982
rect 9903 36951 12761 36982
rect 9903 36945 9908 36951
rect 9846 36944 9908 36945
rect 5764 36875 6102 36886
rect 5723 36849 12773 36875
rect 28455 36868 28470 37045
rect 5723 36650 5773 36849
rect 5764 36624 5773 36650
rect 6096 36650 12773 36849
rect 24326 36715 28470 36868
rect 28676 36868 28786 37045
rect 28676 36715 28818 36868
rect 24326 36662 28818 36715
rect 6096 36624 6102 36650
rect 5764 36618 6102 36624
rect 10181 36548 10229 36549
rect 2710 36520 2974 36544
rect 2710 36426 2731 36520
rect 2702 36201 2731 36426
rect 2710 36197 2731 36201
rect 2956 36426 2974 36520
rect 10181 36507 10185 36548
rect 10226 36546 10229 36548
rect 10226 36508 12760 36546
rect 10226 36507 10229 36508
rect 10181 36506 10229 36507
rect 31294 36496 31687 36505
rect 31294 36460 31329 36496
rect 2956 36201 12733 36426
rect 24326 36290 31329 36460
rect 31652 36290 31687 36496
rect 24326 36254 31687 36290
rect 31294 36253 31687 36254
rect 2956 36197 2974 36201
rect 1487 36180 1776 36188
rect 2710 36184 2974 36197
rect 1487 35992 1578 36180
rect 1484 35857 1578 35992
rect 1764 35992 1776 36180
rect 9834 36165 9896 36168
rect 9834 36113 9837 36165
rect 9889 36159 9896 36165
rect 9889 36118 12728 36159
rect 9889 36113 9896 36118
rect 9834 36109 9896 36113
rect 35344 36108 35915 36183
rect 10181 36069 10235 36072
rect 10181 36028 10190 36069
rect 10231 36028 12724 36069
rect 34174 36054 34524 36080
rect 10181 36024 10235 36028
rect 34174 36026 34188 36054
rect 1764 35857 12696 35992
rect 1484 35806 12696 35857
rect 24326 35849 34188 36026
rect 34511 36026 34524 36054
rect 34511 35849 34533 36026
rect 24326 35821 34533 35849
rect 35344 35785 35622 36108
rect 35821 35785 35915 36108
rect 24344 35719 26677 35724
rect 24344 35687 26448 35719
rect 26670 35687 26677 35719
rect 24344 35681 26677 35687
rect 35344 35619 35915 35785
rect 35300 35615 35915 35619
rect 24326 35569 35915 35615
rect 2373 35340 12725 35548
rect 24326 35379 35899 35569
rect 2373 33329 2581 35340
rect 34766 35141 34975 35159
rect 2789 34852 12773 35060
rect 24326 34932 34975 35141
rect 2366 33321 2600 33329
rect 2366 32998 2383 33321
rect 2591 32998 2600 33321
rect 2366 32992 2600 32998
rect 2373 32905 2581 32992
rect 2789 30469 2997 34852
rect 2767 30462 2997 30469
rect 2767 30139 2773 30462
rect 2981 30139 2997 30462
rect 2767 30128 2997 30139
rect 2789 30095 2997 30128
rect 3223 34370 12773 34578
rect 24326 34392 34561 34601
rect 3223 27621 3431 34370
rect 3677 33900 12773 34108
rect 24326 33904 34153 34113
rect 3202 27603 3459 27621
rect 3202 27280 3236 27603
rect 3444 27280 3459 27603
rect 3202 27261 3459 27280
rect 3223 27257 3431 27261
rect 3677 24759 3885 33900
rect 4112 33474 12773 33682
rect 3661 24744 3900 24759
rect 3661 24421 3677 24744
rect 3885 24421 3900 24744
rect 3661 24402 3900 24421
rect 3677 24349 3885 24402
rect 4112 21898 4320 33474
rect 24326 33384 33744 33593
rect 4546 33067 12773 33275
rect 4094 21885 4339 21898
rect 4094 21562 4111 21885
rect 4319 21562 4339 21885
rect 4094 21546 4339 21562
rect 4112 21534 4320 21546
rect 4546 19047 4754 33067
rect 24326 32880 33331 33089
rect 4962 32652 12773 32860
rect 26423 32758 26876 32766
rect 24354 32757 26883 32758
rect 4521 18674 4781 19047
rect 4546 18641 4754 18674
rect 4962 16184 5170 32652
rect 24354 32648 26432 32757
rect 26860 32648 26883 32757
rect 24354 32643 26883 32648
rect 26423 32641 26876 32643
rect 9844 32563 9904 32564
rect 9844 32511 9847 32563
rect 9899 32559 9904 32563
rect 9899 32515 12778 32559
rect 9899 32511 9904 32515
rect 9844 32508 9904 32511
rect 10187 32461 10233 32462
rect 10187 32417 10190 32461
rect 10231 32417 12774 32461
rect 10187 32415 10233 32417
rect 5387 32137 12773 32345
rect 24358 32329 32907 32538
rect 4920 16167 5191 16184
rect 4920 15844 4965 16167
rect 5173 15844 5191 16167
rect 4920 15817 5191 15844
rect 4962 15745 5170 15817
rect 5387 13322 5595 32137
rect 5813 31711 12773 31919
rect 5354 12974 5628 13322
rect 5387 12893 5595 12974
rect 5813 10493 6021 31711
rect 6228 31207 12773 31415
rect 5791 10449 6070 10493
rect 5791 10126 5827 10449
rect 6035 10126 6070 10449
rect 5791 10088 6070 10126
rect 5813 10060 6021 10088
rect 6228 7615 6436 31207
rect 6663 30646 12773 30854
rect 6179 7590 6462 7615
rect 6179 7267 6224 7590
rect 6432 7267 6462 7590
rect 6179 7237 6462 7267
rect 6228 7181 6436 7237
rect 6663 4757 6871 30646
rect 7079 30176 12773 30384
rect 6628 4731 6893 4757
rect 6628 4408 6668 4731
rect 6876 4408 6893 4731
rect 6628 4385 6893 4408
rect 6663 4384 6871 4385
rect 7079 1887 7287 30176
rect 7060 1872 7327 1887
rect 7060 1549 7098 1872
rect 7306 1549 7327 1872
rect 7060 1534 7327 1549
rect 13233 951 13567 30190
rect 14199 521 14401 30180
rect 14605 678 14807 30180
rect 14605 522 14808 678
rect 15002 677 15204 30180
rect 15402 677 15604 30180
rect 14605 521 14807 522
rect 15001 521 15204 677
rect 15401 521 15604 677
rect 15807 521 16009 30180
rect 16208 678 16410 30180
rect 16207 522 16410 678
rect 16208 521 16410 522
rect 16608 521 16810 30180
rect 17017 521 17219 30180
rect 17430 677 17632 30180
rect 17830 677 18032 30180
rect 18226 677 18428 30180
rect 17429 521 17632 677
rect 17829 521 18032 677
rect 18225 521 18428 677
rect 18631 678 18833 30180
rect 18631 522 18834 678
rect 18631 521 18833 522
rect 19040 521 19242 30180
rect 19441 676 19643 30180
rect 19845 677 20047 30180
rect 19441 521 19644 676
rect 19845 521 20048 677
rect 20254 675 20456 30180
rect 20254 521 20457 675
rect 20659 521 20861 30180
rect 21056 521 21258 30180
rect 21468 521 21670 30180
rect 19442 520 19644 521
rect 20255 519 20457 521
rect 21881 520 22083 30180
rect 22282 521 22484 30180
rect 22683 689 22885 30180
rect 22683 523 22887 689
rect 23092 687 23294 30180
rect 23092 521 23295 687
rect 23509 521 23711 30180
rect 23909 687 24111 30180
rect 24310 687 24512 30180
rect 24706 687 24908 30180
rect 23909 521 24112 687
rect 24307 521 24512 687
rect 24705 521 24908 687
rect 25111 687 25313 30180
rect 25517 687 25719 30180
rect 32698 19186 32907 32329
rect 33122 21833 33331 32880
rect 33535 24681 33744 33384
rect 33944 27558 34153 33904
rect 34352 30408 34561 34392
rect 34766 33264 34975 34932
rect 34746 33249 34989 33264
rect 34746 32926 34767 33249
rect 34976 32926 34989 33249
rect 34746 32910 34989 32926
rect 34766 32843 34975 32910
rect 34328 30390 34579 30408
rect 34328 30067 34342 30390
rect 34551 30067 34579 30390
rect 34328 30051 34579 30067
rect 33924 27531 34176 27558
rect 33924 27208 33944 27531
rect 34153 27208 34176 27531
rect 33924 27187 34176 27208
rect 33944 27184 34153 27187
rect 33508 24672 33744 24681
rect 33508 24349 33519 24672
rect 33728 24349 33744 24672
rect 33508 24339 33744 24349
rect 33535 24268 33744 24339
rect 33105 21813 33348 21833
rect 33105 21490 33125 21813
rect 33334 21490 33348 21813
rect 33105 21462 33348 21490
rect 32699 18996 32907 19186
rect 32699 18984 32908 18996
rect 32688 18978 32908 18984
rect 32662 18610 32915 18978
rect 32688 18608 32897 18610
rect 36806 17339 36880 17373
rect 36108 17236 36248 17314
rect 36740 17299 36881 17339
rect 36107 17224 36248 17236
rect 36742 17230 36880 17299
rect 36106 17209 36248 17224
rect 36106 17119 36247 17209
rect 36741 17113 36881 17230
rect 26339 16496 26799 16501
rect 26339 16054 26350 16496
rect 26792 16423 26799 16496
rect 26792 16255 36254 16423
rect 26792 16126 36267 16255
rect 26792 16054 26799 16126
rect 26339 16044 26799 16054
rect 25111 521 25315 687
rect 25517 521 25721 687
rect 415 33 555 230
rect 1045 0 1185 366
use sky130_hilas_LeftProtection  sky130_hilas_LeftProtection_0
timestamp 1628616568
transform 1 0 2190 0 1 8665
box 0 0 1380 37167
use sky130_hilas_TopLevelTextStructure  sky130_hilas_TopLevelTextStructure_0
timestamp 1628616711
transform 1 0 12478 0 1 30961
box 0 0 13573 7816
use sky130_hilas_TopProtection  sky130_hilas_TopProtection_0
timestamp 1628616684
transform 1 0 1593 0 1 37623
box 0 0 34133 1393
use sky130_hilas_RightProtection  sky130_hilas_RightProtection_0
timestamp 1628616667
transform 1 0 37986 0 1 8593
box 0 0 1386 20013
<< labels >>
rlabel metal1 37160 18079 37285 18468 0 IO07
port 1 nsew
rlabel metal1 37160 20940 37285 21329 0 IO08
port 2 nsew
rlabel metal1 37158 23798 37283 24187 0 IO09
port 3 nsew
rlabel metal1 37160 26659 37285 27048 0 IO10
port 4 nsew
rlabel metal1 37159 29515 37284 29904 0 IO11
port 5 nsew
rlabel metal1 37159 32375 37284 32764 0 IO12
port 6 nsew
rlabel metal1 37160 35235 37285 35624 0 IO13
port 7 nsew
rlabel metal1 0 35305 125 35694 0 IO25
port 8 nsew
rlabel metal1 1 32447 126 32836 0 IO26
port 9 nsew
rlabel metal1 0 29587 125 29976 0 IO27
port 10 nsew
rlabel metal1 2 26728 127 27117 0 IO28
port 11 nsew
rlabel metal1 1 23870 126 24259 0 IO29
port 12 nsew
rlabel metal1 0 21010 125 21399 0 IO30
port 13 nsew
rlabel metal1 1 18152 126 18541 0 IO31
port 14 nsew
rlabel metal1 4 15294 129 15683 0 IO32
port 15 nsew
rlabel metal1 2 12433 127 12822 0 IO33
port 16 nsew
rlabel metal1 1 9574 126 9963 0 IO34
port 17 nsew
rlabel metal1 1 6715 126 7104 0 IO35
port 18 nsew
rlabel metal1 2 3856 127 4245 0 IO36
port 19 nsew
rlabel metal1 2 998 127 1387 0 IO37
port 20 nsew
rlabel metal2 329 38210 497 38501 0 VSSA1
port 21 nsew
rlabel metal1 2362 38791 2751 38908 0 ANALOG10
port 22 nsew
rlabel metal1 5221 38790 5610 38907 0 ANALOG09
port 23 nsew
rlabel metal1 8080 38790 8469 38907 0 ANALOG08
port 24 nsew
rlabel metal1 12270 38793 12659 38910 0 ANALOG07
port 25 nsew
rlabel metal1 16482 38791 16871 38908 0 ANALOG06
port 26 nsew
rlabel metal1 19341 38791 19730 38908 0 ANALOG05
port 27 nsew
rlabel metal1 22201 38791 22590 38908 0 ANALOG04
port 28 nsew
rlabel metal1 25060 38791 25449 38908 0 ANALOG03
port 29 nsew
rlabel metal1 27919 38791 28308 38908 0 ANALOG02
port 30 nsew
rlabel metal1 30778 38790 31167 38907 0 ANALOG01
port 31 nsew
rlabel metal1 33637 38790 34026 38907 0 ANALOG00
port 32 nsew
rlabel metal2 36849 38245 36968 38503 0 VSSA1
port 33 nsew
rlabel metal2 1045 0 1185 140 0 VDDA1
port 34 nsew
rlabel metal2 415 33 555 173 0 VSSA1
port 33 nsew
rlabel metal2 36107 17119 36247 17236 0 VDDA1
port 34 nsew
rlabel metal2 36741 17113 36881 17230 0 VSSA1
port 33 nsew
rlabel metal2 14199 521 14401 677 0 LADATAOUT00
port 36 nsew
rlabel metal2 14606 522 14808 678 0 LADATAOUT01
port 35 nsew
rlabel metal2 15001 521 15203 677 0 LADATAOUT02
port 37 nsew
rlabel metal2 15401 521 15603 677 0 LADATAOUT03
port 38 nsew
rlabel metal2 15807 521 16009 677 0 LADATAOUT04
port 39 nsew
rlabel metal2 16207 522 16409 678 0 LADATAOUT05
port 40 nsew
rlabel metal2 16608 521 16810 677 0 LADATAOUT06
port 41 nsew
rlabel metal2 17017 521 17219 677 0 LADATAOUT07
port 42 nsew
rlabel metal2 17429 521 17631 677 0 LADATAOUT08
port 43 nsew
rlabel metal2 17829 521 18031 677 0 LADATAOUT09
port 44 nsew
rlabel metal2 18225 521 18427 677 0 LADATAOUT10
port 45 nsew
rlabel metal2 18632 522 18834 678 0 LADATAOUT11
port 46 nsew
rlabel metal2 19040 521 19242 677 0 LADATAOUT12
port 47 nsew
rlabel metal2 19442 520 19644 676 0 LADATAOUT13
port 48 nsew
rlabel metal2 19846 521 20048 677 0 LADATAOUT14
port 49 nsew
rlabel metal2 20255 519 20457 675 0 LADATAOUT15
port 50 nsew
rlabel metal2 20659 521 20861 677 0 LADATA16
port 51 nsew
rlabel metal2 21056 521 21258 677 0 LADATAOUT17
port 52 nsew
rlabel metal2 21468 522 21670 678 0 LADATAOUT18
port 53 nsew
rlabel metal2 21881 520 22083 676 0 LADATAOUT19
port 54 nsew
rlabel metal2 22282 521 22484 677 0 LADATAOUT20
port 55 nsew
rlabel metal2 22683 523 22887 689 0 LADATAOUT21
port 56 nsew
rlabel metal2 23092 521 23295 687 0 LADATAOUT22
port 57 nsew
rlabel metal2 23507 521 23710 687 0 LADATAOUT23
port 58 nsew
rlabel metal2 23909 521 24112 687 0 LADATAOUT24
port 59 nsew
rlabel metal2 24307 521 24510 687 0 LADATAIN00
port 60 nsew
rlabel metal2 24705 521 24908 687 0 LADATAIN01
port 61 nsew
rlabel metal2 25112 521 25315 687 0 LADATAIN02
port 62 nsew
rlabel metal2 25518 521 25721 687 0 LADATAIN03
port 63 nsew
rlabel metal2 36151 16126 36267 16252 0 VCCA
port 64 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
