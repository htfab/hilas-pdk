magic
tech sky130A
timestamp 1607261501
<< error_p >>
rect -454 77 -425 93
rect -375 77 -346 93
rect -296 77 -267 93
rect -217 77 -188 93
rect -454 43 -453 44
rect -426 43 -425 44
rect -375 43 -374 44
rect -347 43 -346 44
rect -296 43 -295 44
rect -268 43 -267 44
rect -217 43 -216 44
rect -189 43 -188 44
rect -504 14 -486 43
rect -455 42 -424 43
rect -376 42 -345 43
rect -297 42 -266 43
rect -218 42 -187 43
rect -454 35 -425 42
rect -375 35 -346 42
rect -296 35 -267 42
rect -217 35 -188 42
rect -454 21 -444 35
rect -197 21 -188 35
rect -454 15 -425 21
rect -375 15 -346 21
rect -296 15 -267 21
rect -217 15 -188 21
rect -455 14 -424 15
rect -376 14 -345 15
rect -297 14 -266 15
rect -218 14 -187 15
rect -155 14 -138 43
rect -454 13 -453 14
rect -426 13 -425 14
rect -375 13 -374 14
rect -347 13 -346 14
rect -296 13 -295 14
rect -268 13 -267 14
rect -217 13 -216 14
rect -189 13 -188 14
rect -454 -36 -425 -21
rect -375 -36 -346 -21
rect -296 -36 -267 -21
rect -217 -36 -188 -21
<< nwell >>
rect -521 -54 -121 110
<< mvpmos >>
rect -486 43 -155 77
rect -486 14 -454 43
rect -425 14 -375 43
rect -346 14 -296 43
rect -267 14 -217 43
rect -188 14 -155 43
rect -486 -21 -155 14
<< mvpdiff >>
rect -454 37 -425 43
rect -454 20 -448 37
rect -431 20 -425 37
rect -454 14 -425 20
rect -375 37 -346 43
rect -375 20 -369 37
rect -352 20 -346 37
rect -375 14 -346 20
rect -296 37 -267 43
rect -296 20 -290 37
rect -273 20 -267 37
rect -296 14 -267 20
rect -217 37 -188 43
rect -217 20 -211 37
rect -194 20 -188 37
rect -217 14 -188 20
<< mvpdiffc >>
rect -448 20 -431 37
rect -369 20 -352 37
rect -290 20 -273 37
rect -211 20 -194 37
<< poly >>
rect -502 77 -140 91
rect -502 -21 -486 77
rect -155 -21 -140 77
rect -502 -35 -140 -21
<< locali >>
rect -486 71 -155 77
rect -486 54 -329 71
rect -312 54 -155 71
rect -486 37 -155 54
rect -486 20 -448 37
rect -431 20 -369 37
rect -352 36 -290 37
rect -352 20 -329 36
rect -486 19 -329 20
rect -312 20 -290 36
rect -273 20 -211 37
rect -194 20 -155 37
rect -312 19 -155 20
rect -486 2 -155 19
rect -486 -15 -329 2
rect -312 -15 -155 2
rect -486 -21 -155 -15
<< viali >>
rect -329 54 -312 71
rect -329 19 -312 36
rect -329 -15 -312 2
<< metal1 >>
rect -333 71 -309 77
rect -333 54 -329 71
rect -312 54 -309 71
rect -333 36 -309 54
rect -333 19 -329 36
rect -312 19 -309 36
rect -333 13 -309 19
rect -332 2 -309 13
rect -332 -15 -329 2
rect -312 -13 -309 2
rect -312 -15 -308 -13
rect -332 -35 -308 -15
<< end >>
