magic
tech sky130A
timestamp 1627744303
<< error_s >>
rect 568 189 618 200
rect 640 189 690 200
rect 534 158 568 159
rect 568 147 618 158
rect 640 147 690 158
rect 327 126 367 128
rect 463 126 502 128
rect 534 126 566 128
rect 617 126 626 128
rect 325 51 327 101
rect 367 51 369 101
rect 460 51 463 101
rect 502 51 505 101
rect 640 39 645 63
rect 664 22 669 39
rect 325 -28 327 22
rect 367 -28 369 22
rect 460 -28 463 22
rect 502 -28 505 22
rect 325 -181 327 -131
rect 367 -181 369 -131
rect 460 -181 463 -131
rect 502 -181 505 -131
rect 640 -181 645 -157
rect 664 -198 669 -181
rect 325 -260 327 -210
rect 367 -260 369 -210
rect 460 -260 463 -210
rect 502 -260 505 -210
rect 327 -287 367 -285
rect 463 -287 502 -285
rect 534 -287 566 -285
rect 617 -287 626 -285
rect 568 -317 618 -306
rect 640 -317 690 -306
rect 534 -318 568 -317
rect 568 -359 618 -348
rect 640 -359 690 -348
<< nwell >>
rect -337 -242 -281 0
rect -361 -381 -319 -374
<< psubdiff >>
rect -95 -42 -70 121
rect -95 -59 -92 -42
rect -73 -59 -70 -42
rect -95 -72 -70 -59
rect -95 -75 268 -72
rect -95 -76 146 -75
rect -95 -93 -71 -76
rect -52 -93 -28 -76
rect -9 -93 16 -76
rect 35 -93 56 -76
rect 75 -93 100 -76
rect 119 -92 146 -76
rect 165 -76 268 -75
rect 165 -92 190 -76
rect 119 -93 190 -92
rect 209 -93 236 -76
rect 255 -93 268 -76
rect -95 -97 268 -93
rect -95 -110 -70 -97
rect -95 -127 -92 -110
rect -73 -127 -70 -110
rect -95 -281 -70 -127
<< mvnsubdiff >>
rect -337 -242 -281 0
<< psubdiffcont >>
rect -92 -59 -73 -42
rect -71 -93 -52 -76
rect -28 -93 -9 -76
rect 16 -93 35 -76
rect 56 -93 75 -76
rect 100 -93 119 -76
rect 146 -92 165 -75
rect 190 -93 209 -76
rect 236 -93 255 -76
rect -92 -127 -73 -110
<< poly >>
rect -237 134 331 151
rect -237 126 -185 134
rect -2 91 20 134
rect 166 91 188 134
rect 276 51 314 101
rect 276 -210 291 51
rect 384 -28 398 -27
rect 384 -131 406 -28
rect 276 -233 316 -210
rect 272 -238 316 -233
rect 272 -255 280 -238
rect 297 -255 316 -238
rect 272 -260 316 -255
rect -3 -293 17 -260
rect 169 -293 189 -260
rect 272 -263 300 -260
rect -280 -310 331 -293
<< polycont >>
rect 280 -255 297 -238
<< locali >>
rect 386 163 474 180
rect 386 124 403 163
rect 364 107 403 124
rect 444 107 466 124
rect 221 28 329 45
rect 362 28 470 45
rect -92 -42 -73 -34
rect 464 -51 472 -34
rect -92 -75 -73 -59
rect -92 -76 146 -75
rect -92 -93 -71 -76
rect -52 -93 -28 -76
rect -9 -93 16 -76
rect 35 -93 56 -76
rect 75 -93 100 -76
rect 119 -92 146 -76
rect 165 -76 263 -75
rect 165 -92 190 -76
rect 119 -93 190 -92
rect 209 -93 236 -76
rect 255 -93 263 -76
rect -92 -110 -73 -93
rect 338 -108 355 -51
rect 356 -111 364 -110
rect 422 -111 427 -110
rect 356 -115 427 -111
rect 354 -119 427 -115
rect -92 -135 -73 -127
rect 347 -131 431 -119
rect 464 -125 469 -108
rect 206 -204 330 -187
rect 362 -204 470 -187
rect 280 -236 297 -230
rect 280 -264 297 -257
rect 364 -267 410 -266
rect 363 -282 410 -267
rect 364 -283 410 -282
rect 445 -283 466 -266
rect 391 -317 410 -283
rect 391 -335 487 -317
<< viali >>
rect 278 -238 299 -236
rect 278 -255 280 -238
rect 280 -255 297 -238
rect 297 -255 299 -238
rect 278 -257 299 -255
<< metal1 >>
rect -361 -382 -319 223
rect -113 -382 -90 223
rect 279 -230 297 223
rect 274 -236 303 -230
rect 274 -257 278 -236
rect 299 -257 303 -236
rect 274 -264 303 -257
rect 279 -382 297 -264
rect 384 -382 405 223
rect 427 -382 446 223
rect 472 -56 493 223
rect 661 217 680 223
rect 705 218 721 223
rect 621 -101 645 -59
rect 472 -332 491 -107
rect 522 -332 523 -331
rect 469 -382 492 -332
rect 661 -382 680 -377
rect 705 -382 721 -377
<< metal2 >>
rect 484 173 516 175
rect -395 155 516 173
rect 749 155 757 173
rect -395 0 576 19
rect -395 -73 621 -69
rect -395 -92 622 -73
rect -395 -186 577 -167
rect 510 -315 526 -313
rect -395 -320 526 -315
rect -395 -330 514 -320
rect 749 -332 757 -314
use sky130_hilas_wellContact  sky130_hilas_wellContact_1
timestamp 1627744303
transform 1 0 1054 0 1 404
box -1449 -441 -1275 -255
use sky130_hilas_wellContact  sky130_hilas_wellContact_0
timestamp 1627744303
transform 1 0 1054 0 1 231
box -1449 -441 -1275 -255
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_1
timestamp 1627744303
transform 1 0 1056 0 1 19
box -1451 -400 -1278 -210
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_3
timestamp 1627744303
transform 1 0 1056 0 1 433
box -1451 -400 -1278 -210
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1627744303
transform 1 0 -103 0 1 -92
box -10 -8 13 21
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_2
timestamp 1627744303
transform -1 0 -752 0 -1 -231
box -1005 -380 -733 -211
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_0
timestamp 1627744303
transform -1 0 -752 0 1 62
box -1005 -380 -733 -211
use sky130_hilas_poly2m1  sky130_hilas_poly2m1_0
timestamp 1627744303
transform 1 0 389 0 1 -74
box -9 -26 24 25
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1627744303
transform 1 0 434 0 1 -123
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_3
timestamp 1627744303
transform 1 0 480 0 1 -141
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_2
timestamp 1627744303
transform 1 0 435 0 1 -281
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_5
timestamp 1627744303
transform 1 0 478 0 1 -332
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_6
timestamp 1627744303
transform 1 0 481 0 1 165
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_4
timestamp 1627744303
transform 1 0 434 0 1 109
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_7
timestamp 1627744303
transform 1 0 481 0 1 -34
box -10 -8 13 21
use sky130_hilas_horizTransCell01  sky130_hilas_horizTransCell01_0
timestamp 1627744303
transform 1 0 790 0 1 -429
box -476 48 -33 359
use sky130_hilas_horizTransCell01  sky130_hilas_horizTransCell01_1
timestamp 1627744303
transform 1 0 790 0 -1 270
box -476 48 -33 359
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1627744303
transform 1 0 562 0 1 3
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1627744303
transform 1 0 563 0 1 -166
box -14 -15 20 18
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1627744303
transform 1 0 628 0 1 -85
box -9 -10 23 22
<< labels >>
rlabel metal1 -361 216 -319 223 0 VTUN
port 11 nsew analog default
rlabel metal1 -113 216 -90 223 0 VGND
port 10 nsew ground default
rlabel space 705 217 721 222 0 VINJ
port 2 nsew analog default
rlabel metal2 -395 -330 -391 -315 3 DRAIN2
port 12 e analog default
rlabel metal2 -395 155 -389 173 0 DRAIN1
port 15 nsew analog default
rlabel metal1 427 217 446 223 0 GATE1
port 9 nsew analog default
rlabel metal1 469 -381 492 -357 0 VIN2
port 7 nsew analog default
rlabel metal1 279 -382 297 -375 0 RUN
port 6 nsew analog default
rlabel metal1 384 -382 405 -375 0 PROG
port 5 nsew analog default
rlabel metal1 279 216 297 223 0 RUN
port 6 nsew analog default
rlabel metal1 384 217 405 223 0 PROG
port 5 nsew analog default
rlabel metal1 472 191 493 222 0 VIN1
port 8 nsew analog default
rlabel metal1 661 217 680 223 0 COLSEL1
port 1 nsew analog default
rlabel metal1 661 -382 680 -377 0 COLSEL1
port 1 nsew analog default
rlabel metal1 705 -382 721 -377 0 VINJ
port 2 nsew analog default
rlabel metal2 749 155 757 173 0 DRAIN1
port 3 nsew analog default
rlabel metal2 749 -332 757 -314 0 DRAIN2
port 4 nsew analog default
rlabel metal1 427 -381 446 -376 0 GATE1
port 9 nsew analog default
rlabel metal1 -113 -382 -90 -375 0 VGND
port 10 nsew ground default
rlabel metal1 -361 -381 -319 -374 0 VTUN
port 11 nsew analog default
rlabel metal2 -395 -92 -389 -69 0 COL1
port 16 nsew
rlabel metal2 -395 0 -389 19 0 ROW1
port 17 nsew
rlabel metal2 -395 -186 -389 -167 0 ROW2
port 18 nsew
<< end >>
