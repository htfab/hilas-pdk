magic
tech sky130A
timestamp 1627737364
<< metal1 >>
rect -898 27122 -834 27516
rect -2065 26640 -1984 27030
rect -898 24264 -834 24658
rect -2065 23781 -1984 24171
rect -897 21403 -833 21797
rect -2065 20922 -1984 21312
rect -898 18545 -834 18939
rect -2064 18063 -1983 18453
rect -897 15687 -833 16081
rect -2065 15204 -1984 15594
rect -898 12828 -834 13222
rect -2065 12345 -1984 12735
rect -898 9969 -834 10363
rect -2065 9487 -1984 9877
rect -898 7109 -834 7503
rect -2063 6628 -1982 7018
rect -898 4250 -834 4644
rect -2064 3768 -1983 4158
rect -899 1393 -835 1787
rect -2064 909 -1983 1299
rect -899 -1467 -835 -1073
rect -2064 -1950 -1983 -1560
rect -897 -4327 -833 -3933
rect -2063 -4809 -1982 -4419
rect -897 -7184 -833 -6790
rect -2065 -7668 -1984 -7278
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_0
timestamp 1627735001
transform 0 -1 -1126 1 0 -7694
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_1
timestamp 1627735001
transform 0 -1 -1126 1 0 -4835
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_2
timestamp 1627735001
transform 0 -1 -1126 1 0 -1976
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_3
timestamp 1627735001
transform 0 -1 -1126 1 0 883
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_4
timestamp 1627735001
transform 0 -1 -1126 1 0 3742
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_6
timestamp 1627735001
transform 0 -1 -1126 1 0 6601
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_9
timestamp 1627735001
transform 0 -1 -1126 1 0 9460
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_7
timestamp 1627735001
transform 0 -1 -1126 1 0 12319
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_8
timestamp 1627735001
transform 0 -1 -1126 1 0 15178
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_5
timestamp 1627735001
transform 0 -1 -1126 1 0 18037
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_10
timestamp 1627735001
transform 0 -1 -1126 1 0 20896
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_11
timestamp 1627735001
transform 0 -1 -1126 1 0 23755
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_12
timestamp 1627735001
transform 0 -1 -1126 1 0 26614
box -745 -229 2114 858
<< labels >>
rlabel metal1 -2065 26640 -1984 27030 0 IO25
port 1 nsew
rlabel metal1 -2065 23781 -1984 24171 0 IO26
port 2 nsew
rlabel metal1 -2065 20922 -1984 21312 0 IO27
port 3 nsew
rlabel metal1 -2064 18063 -1983 18453 0 IO28
port 4 nsew
rlabel metal1 -2065 15204 -1984 15594 0 IO29
port 5 nsew
rlabel metal1 -2065 12345 -1984 12735 0 IO30
port 6 nsew
rlabel metal1 -2065 9487 -1984 9877 0 IO31
port 7 nsew
rlabel metal1 -2063 6628 -1982 7018 0 IO32
port 8 nsew
rlabel metal1 -2064 3768 -1983 4158 0 IO33
port 9 nsew
rlabel metal1 -2064 909 -1983 1299 0 IO34
port 10 nsew
rlabel metal1 -2064 -1950 -1983 -1560 0 IO35
port 11 nsew
rlabel metal1 -2063 -4809 -1982 -4419 0 IO36
port 12 nsew
rlabel metal1 -2065 -7668 -1984 -7278 0 IO37
port 13 nsew
rlabel metal1 -898 27122 -834 27516 0 PIN1
port 14 nsew
rlabel metal1 -898 24264 -834 24658 0 PIN2
port 15 nsew
rlabel metal1 -897 21403 -833 21797 0 PIN3
rlabel metal1 -898 18545 -834 18939 0 PIN4
port 16 nsew
rlabel metal1 -897 15687 -833 16081 0 PIN5
port 17 nsew
rlabel metal1 -898 12828 -834 13222 0 PIN6
port 18 nsew
rlabel metal1 -898 9969 -834 10363 0 PIN7
port 19 nsew
rlabel metal1 -898 7109 -834 7503 0 PIN8
port 20 nsew
rlabel metal1 -898 4250 -834 4644 0 PIN9
port 21 nsew
rlabel metal1 -899 1393 -835 1787 0 PIN10
port 22 nsew
rlabel metal1 -899 -1467 -835 -1073 0 PIN11
port 23 nsew
rlabel metal1 -897 -4327 -833 -3933 0 PIN12
port 24 nsew
rlabel metal1 -897 -7184 -833 -6790 0 PIN13
port 25 nsew
<< end >>
