magic
tech sky130A
timestamp 1634057722
<< checkpaint >>
rect -607 -548 687 745
<< nwell >>
rect 0 0 256 191
<< mvpmos >>
rect 67 85 117 139
<< mvpdiff >>
rect 38 133 67 139
rect 38 91 42 133
rect 60 91 67 133
rect 38 85 67 91
rect 117 128 147 139
rect 117 111 123 128
rect 142 111 147 128
rect 117 85 147 111
<< mvpdiffc >>
rect 42 91 60 133
rect 123 111 142 128
<< nsubdiff >>
rect 147 128 192 139
rect 147 111 161 128
rect 180 111 192 128
rect 147 84 192 111
<< nsubdiffcont >>
rect 161 111 180 128
<< poly >>
rect 67 139 117 152
rect 67 76 117 85
rect 0 59 117 76
<< locali >>
rect 34 133 68 135
rect 34 91 42 133
rect 60 91 68 133
rect 123 128 183 136
rect 142 111 161 128
rect 180 111 183 128
rect 123 97 183 111
rect 123 80 124 97
rect 141 80 162 97
rect 179 80 183 97
rect 123 76 183 80
<< viali >>
rect 124 80 141 97
rect 162 80 179 97
<< metal1 >>
rect 123 153 139 191
rect 123 100 182 153
rect 121 97 182 100
rect 121 80 124 97
rect 141 80 162 97
rect 179 80 182 97
rect 121 76 182 80
rect 123 74 182 76
rect 123 1 139 74
<< metal2 >>
rect 0 99 9 117
rect 39 99 256 117
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1634057699
transform 1 0 23 0 -1 115
box 0 0 34 33
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
