* Copyright 2020 The Hilas PDK Authors
* 
* This file is part of HILAS.
* 
* HILAS is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published by
* the Free Software Foundation, version 3 of the License.
* 
* HILAS is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
* 
* You should have received a copy of the GNU Lesser General Public License
* along with HILAS.  If not, see <https://www.gnu.org/licenses/>.
* 
* Licensed under the Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
* https://www.gnu.org/licenses/lgpl-3.0.en.html
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
* SPDX-License-Identifier: LGPL-3.0
* 
* 

* NGSPICE file created from sky130_hilas_TAcoreblock.ext - technology: sky130A

.subckt sky130_hilas_TACoreBlock2 $SUB
X0 w_n122_224# a_n106_328# a_n106_328# w_n122_224# sky130_fd_pr__pfet_01v8 w=680000u l=300000u
X1 $SUB a_n66_n378# a_n66_n378# $SUB sky130_fd_pr__nfet_01v8 w=330000u l=290000u
X2 a_n106_328# a_n66_n378# $SUB $SUB sky130_fd_pr__nfet_01v8 w=330000u l=290000u
X3 a_128_272# a_124_n238# $SUB $SUB sky130_fd_pr__nfet_01v8 w=330000u l=290000u
X4 w_n122_224# a_n106_328# a_128_272# w_n122_224# sky130_fd_pr__pfet_01v8 w=680000u l=300000u
X5 $SUB a_124_n238# a_124_n238# $SUB sky130_fd_pr__nfet_01v8 w=330000u l=290000u
.ends


* Top level circuit sky130_hilas_TAcoreblock

Xsky130_hilas_TACoreBlock2_0 $SUB sky130_hilas_TACoreBlock2
.end

