* Qucs 0.0.22 /home/ubuntu/.qucs/Hilas_prj/nFETLarge.sch
* Qucs 0.0.22  /home/ubuntu/.qucs/Hilas_prj/nFETLarge.sch
M1 Drain1n  Gate1n  Source1n  0 MOSN
.control
echo "" > spice4qucs.cir.noise
echo "" > spice4qucs.cir.pz
exit
.endc
.END
