magic
tech sky130A
timestamp 1629137146
<< locali >>
rect 1 25 33 29
rect 1 24 34 25
rect 1 7 7 24
rect 24 7 34 24
rect 1 6 34 7
rect 1 3 33 6
<< viali >>
rect 7 7 24 24
<< metal1 >>
rect 0 29 32 32
rect 0 3 3 29
rect 29 3 32 29
rect 0 0 32 3
<< via1 >>
rect 3 24 29 29
rect 3 7 7 24
rect 7 7 24 24
rect 24 7 29 24
rect 3 3 29 7
<< metal2 >>
rect 0 29 31 33
rect 0 3 3 29
rect 29 3 31 29
rect 0 0 31 3
<< end >>
