magic
tech sky130A
timestamp 1632251396
<< checkpaint >>
rect -603 781 690 797
rect -603 776 700 781
rect -603 775 1156 776
rect -603 754 1260 775
rect -603 -514 1318 754
rect -601 -521 1318 -514
rect -547 -535 1318 -521
rect -520 -583 1272 -535
rect -385 -597 1272 -583
rect -385 -604 1231 -597
rect -385 -619 1217 -604
rect -385 -620 909 -619
<< nwell >>
rect 12 0 359 152
<< nmos >>
rect 583 87 623 117
rect 440 24 480 55
rect 583 24 623 55
<< pmos >>
rect 125 85 165 117
rect 125 24 165 55
rect 272 24 312 55
<< ndiff >>
rect 554 111 583 117
rect 554 94 559 111
rect 576 94 583 111
rect 554 87 583 94
rect 623 111 654 117
rect 623 94 630 111
rect 647 94 654 111
rect 623 87 654 94
rect 408 47 440 55
rect 408 30 414 47
rect 431 30 440 47
rect 408 24 440 30
rect 480 47 512 55
rect 480 30 488 47
rect 505 30 512 47
rect 480 24 512 30
rect 554 48 583 55
rect 554 31 560 48
rect 577 31 583 48
rect 554 24 583 31
rect 623 48 653 55
rect 623 31 629 48
rect 646 31 653 48
rect 623 24 653 31
<< pdiff >>
rect 96 110 125 117
rect 96 93 102 110
rect 119 93 125 110
rect 96 85 125 93
rect 165 110 193 117
rect 165 93 171 110
rect 188 93 193 110
rect 165 85 193 93
rect 95 47 125 55
rect 95 30 102 47
rect 119 30 125 47
rect 95 24 125 30
rect 165 47 192 55
rect 165 30 171 47
rect 188 30 192 47
rect 165 24 192 30
rect 243 48 272 55
rect 243 31 249 48
rect 266 31 272 48
rect 243 24 272 31
rect 312 48 341 55
rect 312 31 318 48
rect 335 31 341 48
rect 312 24 341 31
<< ndiffc >>
rect 559 94 576 111
rect 630 94 647 111
rect 414 30 431 47
rect 488 30 505 47
rect 560 31 577 48
rect 629 31 646 48
<< pdiffc >>
rect 102 93 119 110
rect 171 93 188 110
rect 102 30 119 47
rect 171 30 188 47
rect 249 31 266 48
rect 318 31 335 48
<< psubdiff >>
rect 680 47 703 59
rect 680 30 683 47
rect 700 30 703 47
rect 680 18 703 30
<< nsubdiff >>
rect 36 51 68 64
rect 36 34 43 51
rect 60 34 68 51
rect 36 22 68 34
<< psubdiffcont >>
rect 683 30 700 47
<< nsubdiffcont >>
rect 43 34 60 51
<< poly >>
rect 29 125 623 141
rect 125 117 165 125
rect 583 117 623 125
rect 211 98 244 104
rect 125 55 165 85
rect 211 81 219 98
rect 236 81 244 98
rect 211 78 244 81
rect 211 63 480 78
rect 272 55 312 63
rect 440 55 480 63
rect 583 55 623 87
rect 125 11 165 24
rect 272 11 312 24
rect 440 11 480 24
rect 583 11 623 24
<< polycont >>
rect 219 81 236 98
<< locali >>
rect 162 110 559 111
rect 92 98 102 110
rect 75 93 102 98
rect 119 93 127 110
rect 162 93 171 110
rect 188 98 559 110
rect 188 93 219 98
rect 75 85 94 93
rect 73 82 94 85
rect 72 81 94 82
rect 211 81 219 93
rect 236 94 559 98
rect 576 94 584 111
rect 622 94 630 111
rect 647 94 657 111
rect 236 93 584 94
rect 236 81 244 93
rect 675 90 700 110
rect 60 76 94 81
rect 47 73 94 76
rect 43 70 94 73
rect 43 64 92 70
rect 43 59 77 64
rect 43 57 69 59
rect 171 57 187 71
rect 43 55 66 57
rect 43 51 64 55
rect 111 47 129 51
rect 43 23 60 34
rect 94 30 102 47
rect 119 30 129 47
rect 171 47 188 57
rect 171 22 188 30
rect 249 48 266 56
rect 249 26 266 31
rect 318 48 335 57
rect 318 22 335 31
rect 414 47 431 52
rect 414 22 431 30
rect 488 47 505 59
rect 488 21 505 30
rect 560 48 577 56
rect 626 31 629 48
rect 646 31 655 48
rect 683 47 700 90
rect 560 26 577 31
rect 683 22 700 30
<< metal1 >>
rect 74 0 94 152
rect 172 74 189 101
rect 317 76 334 103
rect 489 73 506 107
rect 609 53 628 128
rect 657 0 676 152
<< metal2 >>
rect 0 109 61 129
rect 170 109 708 129
rect 0 59 437 79
rect 0 11 577 31
use sky130_hilas_poly2m1  sky130_hilas_poly2m1_0
timestamp 1632251319
transform 1 0 27 0 1 116
box 0 0 33 51
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1632251372
transform 1 0 38 0 1 119
box 0 0 32 32
use sky130_hilas_li2m1  sky130_hilas_li2m1_2
timestamp 1632251332
transform 1 0 83 0 1 95
box 0 0 23 29
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1632251356
transform 1 0 124 0 1 62
box 0 0 34 33
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1632251372
transform 1 0 177 0 1 111
box 0 0 32 32
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1632251332
transform 1 0 180 0 1 54
box 0 0 23 29
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1632251356
transform 1 0 259 0 1 25
box 0 0 34 33
use sky130_hilas_m12m2  sky130_hilas_m12m2_2
timestamp 1632251372
transform 1 0 319 0 1 112
box 0 0 32 32
use sky130_hilas_li2m1  sky130_hilas_li2m1_3
timestamp 1632251332
transform 1 0 325 0 1 56
box 0 0 23 29
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1632251356
transform 1 0 416 0 1 62
box 0 0 34 33
use sky130_hilas_m12m2  sky130_hilas_m12m2_4
timestamp 1632251372
transform 1 0 494 0 1 114
box 0 0 32 32
use sky130_hilas_li2m1  sky130_hilas_li2m1_4
timestamp 1632251332
transform 1 0 496 0 1 55
box 0 0 23 29
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1632251356
transform 1 0 567 0 1 26
box 0 0 34 33
use sky130_hilas_m12m2  sky130_hilas_m12m2_3
timestamp 1632251372
transform 1 0 598 0 1 113
box 0 0 32 32
use sky130_hilas_li2m1  sky130_hilas_li2m1_5
timestamp 1632251332
transform 1 0 619 0 1 33
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1632251332
transform 1 0 665 0 1 95
box 0 0 23 29
<< labels >>
rlabel metal2 702 109 708 129 0 output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
