magic
tech sky130A
timestamp 1628617015
<< checkpaint >>
rect -454 714 840 715
rect -563 699 840 714
rect -577 -578 840 699
rect -577 -593 826 -578
rect -577 -594 717 -593
<< nmos >>
rect 111 35 138 77
<< ndiff >>
rect 80 61 111 77
rect 80 44 85 61
rect 105 44 111 61
rect 80 35 111 44
rect 138 61 169 77
rect 138 44 144 61
rect 164 44 169 61
rect 138 35 169 44
<< ndiffc >>
rect 85 44 105 61
rect 144 44 164 61
<< poly >>
rect 111 77 138 90
rect 111 27 138 35
rect 30 22 138 27
rect 30 5 38 22
rect 55 12 138 22
rect 55 5 63 12
rect 30 0 63 5
<< polycont >>
rect 38 5 55 22
<< locali >>
rect 85 61 105 69
rect 85 36 105 44
rect 144 61 164 69
rect 144 36 164 44
rect 30 5 38 22
rect 55 5 63 22
<< metal2 >>
rect 0 43 60 60
rect 186 44 208 61
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628616992
transform 1 0 67 0 1 51
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628616992
transform 1 0 176 0 1 52
box 0 0 34 33
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
