magic
tech sky130A
timestamp 1628616977
<< checkpaint >>
rect -630 1796 9207 2023
rect 13490 1853 34763 2023
rect 9947 1796 34763 1853
rect -630 1794 34763 1796
rect -1375 -324 34763 1794
rect -1375 -553 34018 -324
<< metal1 >>
rect 26 1164 415 1244
rect 2885 1164 3274 1244
rect 5744 1164 6133 1244
rect 9934 1166 10323 1246
rect 14146 1164 14535 1244
rect 17005 1164 17394 1244
rect 19865 1164 20254 1244
rect 22724 1164 23113 1244
rect 25582 1164 25971 1244
rect 28441 1164 28830 1244
rect 31301 1164 31690 1244
rect 508 0 903 77
rect 3368 0 3763 77
rect 6226 0 6621 77
rect 10503 0 10751 77
rect 14628 1 15023 78
rect 17487 0 17882 77
rect 20346 0 20741 77
rect 23205 0 23600 77
rect 26065 0 26460 77
rect 28923 0 29318 77
rect 31782 0 32177 77
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_1
timestamp 1628616751
transform 1 0 2859 0 1 306
box 0 0 2859 1087
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_0
timestamp 1628616751
transform 1 0 0 0 1 306
box 0 0 2859 1087
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_2
timestamp 1628616751
transform 1 0 5718 0 1 306
box 0 0 2859 1087
use sky130_hilas_polyresistorGND  sky130_hilas_polyresistorGND_0
timestamp 1628616684
transform 1 0 10577 0 1 134
box 0 0 5547 1089
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_3
timestamp 1628616751
transform 1 0 14120 0 1 306
box 0 0 2859 1087
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_4
timestamp 1628616751
transform 1 0 16979 0 1 306
box 0 0 2859 1087
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_5
timestamp 1628616751
transform 1 0 19838 0 1 306
box 0 0 2859 1087
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_6
timestamp 1628616751
transform 1 0 22697 0 1 306
box 0 0 2859 1087
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_9
timestamp 1628616751
transform 1 0 25556 0 1 306
box 0 0 2859 1087
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_7
timestamp 1628616751
transform 1 0 28415 0 1 306
box 0 0 2859 1087
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_8
timestamp 1628616751
transform 1 0 31274 0 1 306
box 0 0 2859 1087
<< labels >>
rlabel metal1 31301 1164 31690 1244 0 ANALOG00
port 1 nsew
rlabel metal1 28441 1164 28830 1244 0 ANALOG01
port 2 nsew
rlabel metal1 25582 1164 25971 1244 0 ANALOG02
port 3 nsew
rlabel metal1 22724 1164 23113 1244 0 ANALOG03
port 4 nsew
rlabel metal1 19865 1164 20254 1244 0 ANALOG04
port 5 nsew
rlabel metal1 17005 1164 17394 1244 0 ANALOG05
port 6 nsew
rlabel metal1 14146 1164 14535 1244 0 ANALOG06
port 7 nsew
rlabel metal1 9934 1166 10323 1246 0 ANALOG07
port 8 nsew
rlabel metal1 5744 1164 6133 1244 0 ANALOG08
port 9 nsew
rlabel metal1 2885 1164 3274 1244 0 ANALOG09
port 10 nsew
rlabel metal1 26 1164 415 1244 0 ANALOG10
port 11 nsew
rlabel metal1 31782 0 32177 77 0 PIN1
port 12 nsew
rlabel metal1 28923 0 29318 77 0 PIN2
port 13 nsew
rlabel metal1 26065 0 26460 77 0 PIN3
port 14 nsew
rlabel metal1 23205 0 23600 77 0 PIN4
port 15 nsew
rlabel metal1 20346 0 20741 77 0 PIN5
port 16 nsew
rlabel metal1 17487 0 17882 77 0 PIN6
port 17 nsew
rlabel metal1 14628 1 15023 78 0 PIN7
port 18 nsew
rlabel metal1 6226 0 6621 77 0 PIN8
port 19 nsew
rlabel metal1 3368 0 3763 77 0 PIN9
port 20 nsew
rlabel metal1 508 0 903 77 0 PIN10
port 21 nsew
rlabel metal1 10503 0 10751 77 0 VTUN
port 22 nsew
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
