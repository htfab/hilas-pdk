VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_tunvaractorcapcitor
  CLASS BLOCK ;
  FOREIGN sky130_hilas_tunvaractorcapcitor ;
  ORIGIN 14.660 4.420 ;
  SIZE 10.430 BY 7.010 ;
  OBS
      LAYER nwell ;
        RECT -14.660 1.750 -12.750 2.260 ;
        RECT -14.650 -4.400 -12.750 1.750 ;
        RECT -9.920 0.260 -7.130 2.240 ;
        RECT -9.940 -2.530 -7.120 0.260 ;
        RECT -9.900 -4.400 -7.120 -2.530 ;
        RECT -5.720 -4.400 -4.250 2.260 ;
        RECT -5.070 -4.420 -4.250 -4.400 ;
      LAYER li1 ;
        RECT -5.230 1.720 -4.890 1.890 ;
        RECT -5.230 0.930 -4.890 1.100 ;
        RECT -5.230 0.360 -4.890 0.530 ;
        RECT -5.240 -1.170 -4.890 -1.000 ;
        RECT -5.230 -2.690 -4.890 -2.520 ;
        RECT -5.230 -3.250 -4.890 -3.080 ;
        RECT -13.790 -3.950 -13.510 -3.520 ;
        RECT -6.600 -3.780 -6.260 -3.610 ;
        RECT -5.230 -4.040 -4.890 -3.870 ;
  END
END sky130_hilas_tunvaractorcapcitor
END LIBRARY

