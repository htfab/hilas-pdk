magic
tech sky130A
timestamp 1629137262
<< checkpaint >>
rect -611 1157 821 1253
rect -612 1126 821 1157
rect -612 -320 839 1126
rect -612 -512 810 -320
rect -611 -608 810 -512
<< error_s >>
rect 1 522 40 525
rect 1 480 40 483
rect 0 426 39 429
rect 0 384 39 387
rect 0 330 39 333
rect 0 288 39 291
rect 0 234 39 237
rect 0 192 39 195
rect 0 138 39 141
rect 0 96 39 99
rect 1 42 40 45
rect 1 0 40 3
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_0
timestamp 1629137183
transform 1 0 18 0 1 118
box 0 0 161 121
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_4
timestamp 1629137183
transform 1 0 18 0 1 214
box 0 0 161 121
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_6
timestamp 1629137183
transform 1 0 18 0 1 406
box 0 0 161 121
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_0
timestamp 1629137127
transform 1 0 19 0 1 502
box 0 0 172 121
use sky130_hilas_pFETdevice01a  sky130_hilas_pFETdevice01a_0
timestamp 1629137174
transform 1 0 19 0 1 22
box 0 0 161 85
use sky130_hilas_pFETdevice01d  sky130_hilas_pFETdevice01d_0
timestamp 1629137210
transform 1 0 18 0 1 310
box 0 0 191 186
<< end >>
