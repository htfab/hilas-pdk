magic
tech sky130A
timestamp 1628707314
<< checkpaint >>
rect 338 1287 1854 1328
rect 49 1281 1854 1287
rect -351 1268 1854 1281
rect -580 -572 1854 1268
rect -351 -584 1854 -572
rect 49 -589 1854 -584
rect 338 -630 1854 -589
<< error_s >>
rect 100 620 129 638
rect 346 618 375 634
rect 425 618 454 634
rect 504 618 533 634
rect 583 618 612 634
rect 100 588 101 589
rect 128 588 129 589
rect 50 559 68 588
rect 99 587 130 588
rect 100 578 129 587
rect 100 569 110 578
rect 119 569 129 578
rect 100 560 129 569
rect 99 559 130 560
rect 161 559 179 588
rect 346 584 347 585
rect 374 584 375 585
rect 425 584 426 585
rect 453 584 454 585
rect 504 584 505 585
rect 532 584 533 585
rect 583 584 584 585
rect 611 584 612 585
rect 100 558 101 559
rect 128 558 129 559
rect 296 555 314 584
rect 345 583 376 584
rect 424 583 455 584
rect 503 583 534 584
rect 582 583 613 584
rect 346 576 375 583
rect 425 576 454 583
rect 504 576 533 583
rect 583 576 612 583
rect 346 562 356 576
rect 603 562 612 576
rect 346 556 375 562
rect 425 556 454 562
rect 504 556 533 562
rect 583 556 612 562
rect 345 555 376 556
rect 424 555 455 556
rect 503 555 534 556
rect 582 555 613 556
rect 645 555 662 584
rect 679 562 681 563
rect 346 554 347 555
rect 374 554 375 555
rect 425 554 426 555
rect 453 554 454 555
rect 504 554 505 555
rect 532 554 533 555
rect 583 554 584 555
rect 611 554 612 555
rect 100 509 129 527
rect 346 505 375 520
rect 425 505 454 520
rect 504 505 533 520
rect 583 505 612 520
rect 100 468 129 486
rect 346 471 375 487
rect 425 471 454 487
rect 504 471 533 487
rect 583 471 612 487
rect 346 437 347 438
rect 374 437 375 438
rect 425 437 426 438
rect 453 437 454 438
rect 504 437 505 438
rect 532 437 533 438
rect 583 437 584 438
rect 611 437 612 438
rect 100 436 101 437
rect 128 436 129 437
rect 50 407 68 436
rect 99 435 130 436
rect 100 426 129 435
rect 100 417 110 426
rect 119 417 129 426
rect 100 408 129 417
rect 99 407 130 408
rect 161 407 179 436
rect 296 408 314 437
rect 345 436 376 437
rect 424 436 455 437
rect 503 436 534 437
rect 582 436 613 437
rect 346 429 375 436
rect 425 429 454 436
rect 504 429 533 436
rect 583 429 612 436
rect 346 415 356 429
rect 603 415 612 429
rect 346 409 375 415
rect 425 409 454 415
rect 504 409 533 415
rect 583 409 612 415
rect 345 408 376 409
rect 424 408 455 409
rect 503 408 534 409
rect 582 408 613 409
rect 645 408 662 437
rect 674 411 687 415
rect 688 411 701 416
rect 674 408 701 411
rect 346 407 347 408
rect 374 407 375 408
rect 425 407 426 408
rect 453 407 454 408
rect 504 407 505 408
rect 532 407 533 408
rect 583 407 584 408
rect 611 407 612 408
rect 100 406 101 407
rect 128 406 129 407
rect 100 357 129 375
rect 346 358 375 373
rect 425 358 454 373
rect 504 358 533 373
rect 583 358 612 373
rect 100 323 129 341
rect 346 324 375 340
rect 425 324 454 340
rect 504 324 533 340
rect 583 324 612 340
rect 100 291 101 292
rect 128 291 129 292
rect 50 262 68 291
rect 99 290 130 291
rect 100 281 129 290
rect 100 272 110 281
rect 119 272 129 281
rect 100 263 129 272
rect 99 262 130 263
rect 161 262 179 291
rect 346 290 347 291
rect 374 290 375 291
rect 425 290 426 291
rect 453 290 454 291
rect 504 290 505 291
rect 532 290 533 291
rect 583 290 584 291
rect 611 290 612 291
rect 100 261 101 262
rect 128 261 129 262
rect 296 261 314 290
rect 345 289 376 290
rect 424 289 455 290
rect 503 289 534 290
rect 582 289 613 290
rect 346 282 375 289
rect 425 282 454 289
rect 504 282 533 289
rect 583 282 612 289
rect 346 268 356 282
rect 603 268 612 282
rect 346 262 375 268
rect 425 262 454 268
rect 504 262 533 268
rect 583 262 612 268
rect 345 261 376 262
rect 424 261 455 262
rect 503 261 534 262
rect 582 261 613 262
rect 645 261 662 290
rect 346 260 347 261
rect 374 260 375 261
rect 425 260 426 261
rect 453 260 454 261
rect 504 260 505 261
rect 532 260 533 261
rect 583 260 584 261
rect 611 260 612 261
rect 100 212 129 230
rect 346 211 375 226
rect 425 211 454 226
rect 504 211 533 226
rect 583 211 612 226
rect 100 169 129 187
rect 346 177 375 193
rect 425 177 454 193
rect 504 177 533 193
rect 583 177 612 193
rect 346 143 347 144
rect 374 143 375 144
rect 425 143 426 144
rect 453 143 454 144
rect 504 143 505 144
rect 532 143 533 144
rect 583 143 584 144
rect 611 143 612 144
rect 100 137 101 138
rect 128 137 129 138
rect 50 108 68 137
rect 99 136 130 137
rect 100 127 129 136
rect 100 118 110 127
rect 119 118 129 127
rect 100 109 129 118
rect 99 108 130 109
rect 161 108 179 137
rect 296 114 314 143
rect 345 142 376 143
rect 424 142 455 143
rect 503 142 534 143
rect 582 142 613 143
rect 346 135 375 142
rect 425 135 454 142
rect 504 135 533 142
rect 583 135 612 142
rect 346 121 356 135
rect 603 121 612 135
rect 346 115 375 121
rect 425 115 454 121
rect 504 115 533 121
rect 583 115 612 121
rect 345 114 376 115
rect 424 114 455 115
rect 503 114 534 115
rect 582 114 613 115
rect 645 114 662 143
rect 346 113 347 114
rect 374 113 375 114
rect 425 113 426 114
rect 453 113 454 114
rect 504 113 505 114
rect 532 113 533 114
rect 583 113 584 114
rect 611 113 612 114
rect 100 107 101 108
rect 128 107 129 108
rect 100 58 129 76
rect 346 64 375 79
rect 425 64 454 79
rect 504 64 533 79
rect 583 64 612 79
<< nwell >>
rect 823 356 858 357
rect 823 340 840 356
rect 857 340 858 356
<< poly >>
rect 660 575 680 579
rect 172 542 321 566
rect 660 563 679 575
rect 172 433 319 457
rect 660 419 679 436
rect 840 356 858 357
rect 856 340 858 356
rect 172 253 321 277
rect 660 261 679 278
rect 172 133 323 157
rect 660 119 679 136
<< polycont >>
rect 823 340 840 357
<< locali >>
rect 814 340 823 357
<< viali >>
rect 840 340 858 357
<< metal1 >>
rect 101 46 128 651
rect 845 360 858 362
rect 837 357 861 360
rect 837 340 840 357
rect 858 340 861 357
rect 837 337 861 340
rect 847 333 858 337
<< metal2 >>
rect 0 594 688 601
rect 0 583 691 594
rect 0 540 901 558
rect 0 452 688 458
rect 0 440 691 452
rect 0 408 687 415
rect 0 397 691 408
rect 0 282 691 299
rect 0 240 691 257
rect 0 142 691 159
rect 0 98 691 115
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_3
timestamp 1628707313
transform 1 0 112 0 1 101
box 0 0 129 129
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_3
timestamp 1628707295
transform 1 0 800 0 1 100
box 0 0 400 164
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_1
timestamp 1628707307
transform 1 0 968 0 1 0
box 0 0 256 191
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_2
timestamp 1628707313
transform 1 0 112 0 1 255
box 0 0 129 129
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_2
timestamp 1628707295
transform 1 0 800 0 1 247
box 0 0 400 164
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_2
timestamp 1628707307
transform 1 0 968 0 -1 397
box 0 0 256 191
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_0
timestamp 1628707307
transform 1 0 968 0 1 300
box 0 0 256 191
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_1
timestamp 1628707313
transform 1 0 112 0 1 400
box 0 0 129 129
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_0
timestamp 1628707313
transform 1 0 112 0 1 552
box 0 0 129 129
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_1
timestamp 1628707295
transform 1 0 800 0 1 394
box 0 0 400 164
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_0
timestamp 1628707295
transform 1 0 800 0 1 541
box 0 0 400 164
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_3
timestamp 1628707307
transform 1 0 968 0 -1 698
box 0 0 256 191
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
