magic
tech sky130A
timestamp 1627218289
<< nwell >>
rect 147 -22 266 265
<< pmos >>
rect 194 -4 220 247
<< pdiff >>
rect 165 223 194 247
rect 165 206 171 223
rect 188 206 194 223
rect 165 189 194 206
rect 165 172 171 189
rect 188 172 194 189
rect 165 155 194 172
rect 165 138 171 155
rect 188 138 194 155
rect 165 121 194 138
rect 165 104 171 121
rect 188 104 194 121
rect 165 87 194 104
rect 165 70 171 87
rect 188 70 194 87
rect 165 53 194 70
rect 165 36 171 53
rect 188 36 194 53
rect 165 19 194 36
rect 165 2 171 19
rect 188 2 194 19
rect 165 -4 194 2
rect 220 223 248 247
rect 220 206 226 223
rect 243 206 248 223
rect 220 189 248 206
rect 220 172 226 189
rect 243 172 248 189
rect 220 155 248 172
rect 220 138 226 155
rect 243 138 248 155
rect 220 121 248 138
rect 220 104 226 121
rect 243 104 248 121
rect 220 87 248 104
rect 220 70 226 87
rect 243 70 248 87
rect 220 53 248 70
rect 220 36 226 53
rect 243 36 248 53
rect 220 19 248 36
rect 220 2 226 19
rect 243 2 248 19
rect 220 -4 248 2
<< pdiffc >>
rect 171 206 188 223
rect 171 172 188 189
rect 171 138 188 155
rect 171 104 188 121
rect 171 70 188 87
rect 171 36 188 53
rect 171 2 188 19
rect 226 206 243 223
rect 226 172 243 189
rect 226 138 243 155
rect 226 104 243 121
rect 226 70 243 87
rect 226 36 243 53
rect 226 2 243 19
<< poly >>
rect 194 247 220 260
rect 194 -17 220 -4
<< locali >>
rect 171 223 188 242
rect 171 189 188 206
rect 171 155 188 172
rect 171 121 188 138
rect 171 87 188 104
rect 171 53 188 70
rect 171 19 188 36
rect 171 -7 188 2
rect 226 223 243 242
rect 226 189 243 206
rect 226 155 243 172
rect 226 121 243 138
rect 226 87 243 104
rect 226 53 243 70
rect 226 19 243 36
rect 226 -8 243 2
<< end >>
