VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_hilas_TA2Cell_1FG_Strong
  CLASS CORE ;
  FOREIGN sky130_hilas_TA2Cell_1FG_Strong ;
  ORIGIN 0.000 0.000 ;
  SIZE 32.820 BY 10.100 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VTUN
    ANTENNADIFFAREA 1.808400 ;
    PORT
      LAYER nwell ;
        RECT 16.180 1.780 17.910 5.350 ;
        RECT 16.750 1.450 17.310 1.780 ;
      LAYER met1 ;
        RECT 15.480 5.950 15.900 6.100 ;
        RECT 16.510 5.950 16.930 6.100 ;
        RECT 15.480 5.810 16.930 5.950 ;
        RECT 16.510 0.050 16.930 5.810 ;
    END
  END VTUN
  PIN PROG
    PORT
      LAYER met1 ;
        RECT 8.240 6.040 8.450 6.100 ;
    END
  END PROG
  PIN GATE1
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT 19.930 3.710 22.650 5.360 ;
        RECT 19.930 3.670 22.640 3.710 ;
        RECT 19.930 2.340 22.640 2.380 ;
        RECT 19.930 0.690 22.650 2.340 ;
      LAYER met1 ;
        RECT 20.210 4.890 20.440 6.100 ;
        RECT 20.210 4.100 20.470 4.890 ;
        RECT 20.210 1.950 20.440 4.100 ;
        RECT 20.210 1.160 20.470 1.950 ;
        RECT 20.210 0.050 20.440 1.160 ;
    END
  END GATE1
  PIN VIN11
    PORT
      LAYER met1 ;
        RECT 7.360 5.990 7.570 6.100 ;
    END
  END VIN11
  PIN VINJ
    ANTENNADIFFAREA 2.163200 ;
    PORT
      LAYER nwell ;
        RECT 24.380 6.100 27.690 6.150 ;
        RECT 24.380 6.090 29.030 6.100 ;
        RECT 24.380 3.100 27.690 6.090 ;
        RECT 24.380 3.030 29.540 3.100 ;
        RECT 24.380 0.000 27.690 3.030 ;
      LAYER met2 ;
        RECT 2.540 6.070 2.850 6.260 ;
        RECT 4.920 6.070 5.240 6.080 ;
        RECT 2.540 5.960 12.290 6.070 ;
        RECT 27.190 5.960 27.510 6.080 ;
        RECT 2.540 5.930 27.510 5.960 ;
        RECT 2.570 5.880 27.510 5.930 ;
        RECT 4.920 5.780 27.510 5.880 ;
        RECT 26.300 3.240 26.620 3.500 ;
        RECT 26.340 3.220 27.520 3.240 ;
        RECT 26.340 2.960 27.560 3.220 ;
        RECT 26.340 2.900 27.520 2.960 ;
        RECT 26.300 2.890 27.520 2.900 ;
        RECT 26.300 2.640 26.620 2.890 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.170 6.080 27.450 6.100 ;
        RECT 27.170 5.780 27.510 6.080 ;
        RECT 27.170 5.450 27.450 5.780 ;
        RECT 27.060 4.850 27.450 5.450 ;
        RECT 27.170 3.250 27.450 4.850 ;
        RECT 27.170 2.930 27.530 3.250 ;
        RECT 27.170 1.300 27.450 2.930 ;
        RECT 27.060 0.700 27.450 1.300 ;
        RECT 27.170 0.050 27.450 0.700 ;
      LAYER via ;
        RECT 27.220 5.800 27.480 6.060 ;
        RECT 27.270 2.960 27.530 3.220 ;
    END
  END VINJ
  PIN VIN22
    PORT
      LAYER met2 ;
        RECT 28.930 6.080 29.240 6.090 ;
        RECT 28.360 6.070 29.240 6.080 ;
        RECT 28.290 5.830 29.240 6.070 ;
        RECT 28.930 5.760 29.240 5.830 ;
    END
  END VIN22
  PIN VIN21
    PORT
      LAYER met2 ;
        RECT 28.690 3.400 29.000 3.440 ;
        RECT 28.370 3.390 29.030 3.400 ;
        RECT 28.370 3.160 29.470 3.390 ;
        RECT 28.690 3.110 29.000 3.160 ;
    END
  END VIN21
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 31.620 6.020 31.930 6.100 ;
        RECT 31.620 5.790 32.820 6.020 ;
        RECT 31.620 5.770 31.930 5.790 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.530 0.050 31.800 0.260 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 30.860 5.960 31.200 6.100 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.330 0.400 29.650 0.550 ;
        RECT 13.140 0.250 29.650 0.400 ;
        RECT 13.140 0.100 13.460 0.250 ;
        RECT 18.940 0.100 19.260 0.250 ;
    END
  END VGND
  PIN OUTPUT2
    PORT
      LAYER met2 ;
        RECT 32.710 2.570 32.820 2.790 ;
    END
  END OUTPUT2
  PIN OUTPUT1
    PORT
      LAYER met2 ;
        RECT 32.710 3.390 32.820 3.620 ;
    END
  END OUTPUT1
  PIN GATESEL1
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER met1 ;
        RECT 5.370 6.100 5.550 9.970 ;
        RECT 5.370 6.040 5.680 6.100 ;
        RECT 5.370 5.440 5.550 6.040 ;
        RECT 5.310 5.100 5.600 5.440 ;
        RECT 5.370 3.920 5.550 5.100 ;
    END
  END GATESEL1
  PIN GATESEL2
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT 26.730 4.640 26.920 6.100 ;
        RECT 26.730 4.610 26.950 4.640 ;
        RECT 26.710 4.340 26.960 4.610 ;
        RECT 26.720 4.330 26.960 4.340 ;
        RECT 26.720 4.090 26.950 4.330 ;
        RECT 26.760 2.060 26.920 4.090 ;
        RECT 26.720 1.820 26.950 2.060 ;
        RECT 26.720 1.810 26.960 1.820 ;
        RECT 26.710 1.540 26.960 1.810 ;
        RECT 26.730 1.510 26.950 1.540 ;
        RECT 26.730 0.050 26.920 1.510 ;
    END
  END GATESEL2
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 4.720 5.420 4.800 5.600 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 4.720 0.550 4.800 0.730 ;
    END
  END DRAIN2
  PIN VIN12
    PORT
      LAYER met1 ;
        RECT 7.370 0.060 7.600 0.180 ;
    END
  END VIN12
  PIN GATE2
    PORT
      LAYER met1 ;
        RECT 7.830 6.020 8.020 6.100 ;
    END
  END GATE2
  PIN RUN
    ANTENNADIFFAREA 1.850000 ;
    PORT
      LAYER met1 ;
        RECT 9.240 7.110 9.470 9.970 ;
        RECT 9.140 6.820 9.470 7.110 ;
        RECT 9.240 6.100 9.470 6.820 ;
        RECT 9.240 6.030 9.500 6.100 ;
        RECT 9.240 3.920 9.470 6.030 ;
    END
  END RUN
  OBS
      LAYER nwell ;
        RECT 0.770 3.870 4.080 10.020 ;
        RECT 5.810 7.580 8.530 9.230 ;
        RECT 5.810 7.540 8.520 7.580 ;
        RECT 5.810 6.210 8.520 6.250 ;
        RECT 5.810 6.100 8.530 6.210 ;
        RECT 4.720 6.090 8.530 6.100 ;
        RECT 4.920 5.780 5.240 6.080 ;
        RECT 5.810 4.560 8.530 6.090 ;
        RECT 10.550 5.650 12.280 9.220 ;
        RECT 30.680 8.200 32.410 10.100 ;
        RECT 31.540 5.960 32.820 6.100 ;
        RECT 30.680 5.920 32.820 5.960 ;
        RECT 11.150 5.320 11.710 5.650 ;
        RECT 30.680 4.060 32.410 5.920 ;
        RECT 11.530 3.930 11.950 4.000 ;
        RECT 29.020 3.160 29.470 3.390 ;
        RECT 31.310 0.000 32.820 1.650 ;
      LAYER li1 ;
        RECT 1.170 9.290 1.370 9.640 ;
        RECT 2.650 9.390 3.180 9.560 ;
        RECT 3.320 9.420 3.510 9.650 ;
        RECT 3.600 9.370 4.480 9.540 ;
        RECT 1.160 9.260 1.370 9.290 ;
        RECT 1.160 8.680 1.380 9.260 ;
        RECT 1.160 8.670 1.370 8.680 ;
        RECT 1.540 8.500 1.730 8.510 ;
        RECT 1.530 8.210 1.730 8.500 ;
        RECT 1.470 7.880 1.740 8.210 ;
        RECT 1.930 7.400 2.100 9.010 ;
        RECT 2.760 7.910 2.930 9.000 ;
        RECT 3.790 8.980 3.980 9.090 ;
        RECT 3.350 8.860 3.980 8.980 ;
        RECT 4.310 8.980 4.480 9.370 ;
        RECT 3.350 8.810 3.900 8.860 ;
        RECT 4.310 8.810 5.050 8.980 ;
        RECT 6.110 8.190 6.340 8.710 ;
        RECT 3.350 8.020 6.340 8.190 ;
        RECT 2.530 7.870 2.930 7.910 ;
        RECT 2.520 7.680 2.930 7.870 ;
        RECT 11.310 7.830 11.860 8.260 ;
        RECT 2.530 7.650 2.930 7.680 ;
        RECT 1.920 7.210 2.100 7.400 ;
        RECT 2.760 7.310 2.930 7.650 ;
        RECT 3.320 7.430 3.510 7.660 ;
        RECT 3.350 7.230 3.700 7.400 ;
        RECT 4.180 7.080 4.390 7.510 ;
        RECT 4.700 7.230 5.040 7.400 ;
        RECT 4.200 7.060 4.370 7.080 ;
        RECT 1.920 6.490 2.100 6.680 ;
        RECT 3.350 6.590 3.700 6.660 ;
        RECT 1.470 5.680 1.740 6.010 ;
        RECT 1.530 5.390 1.730 5.680 ;
        RECT 1.540 5.380 1.730 5.390 ;
        RECT 1.160 5.210 1.370 5.220 ;
        RECT 1.160 4.630 1.380 5.210 ;
        RECT 1.930 4.880 2.100 6.490 ;
        RECT 2.760 6.220 2.930 6.580 ;
        RECT 3.330 6.490 3.700 6.590 ;
        RECT 3.790 6.540 3.980 6.770 ;
        RECT 4.790 6.660 4.960 7.230 ;
        RECT 9.070 7.080 9.260 7.400 ;
        RECT 9.070 6.990 9.350 7.080 ;
        RECT 5.710 6.850 9.350 6.990 ;
        RECT 5.710 6.810 9.260 6.850 ;
        RECT 4.070 6.630 4.120 6.640 ;
        RECT 4.700 6.630 5.040 6.660 ;
        RECT 4.070 6.550 5.040 6.630 ;
        RECT 4.030 6.490 5.040 6.550 ;
        RECT 3.330 6.360 3.520 6.490 ;
        RECT 4.030 6.430 4.870 6.490 ;
        RECT 9.070 6.390 9.260 6.810 ;
        RECT 2.520 6.180 2.930 6.220 ;
        RECT 2.510 5.990 2.930 6.180 ;
        RECT 11.310 6.100 11.860 6.530 ;
        RECT 2.520 5.960 2.930 5.990 ;
        RECT 2.760 4.890 2.930 5.960 ;
        RECT 28.670 6.050 28.840 6.100 ;
        RECT 31.860 6.060 32.060 6.100 ;
        RECT 3.350 5.770 6.280 5.870 ;
        RECT 28.670 5.790 29.230 6.050 ;
        RECT 31.630 5.800 32.060 6.060 ;
        RECT 28.670 5.770 28.840 5.790 ;
        RECT 31.860 5.770 32.060 5.800 ;
        RECT 3.350 5.700 6.340 5.770 ;
        RECT 5.370 5.380 5.540 5.440 ;
        RECT 3.780 5.080 3.970 5.190 ;
        RECT 5.350 5.170 5.560 5.380 ;
        RECT 5.370 5.100 5.540 5.170 ;
        RECT 6.110 5.080 6.340 5.700 ;
        RECT 25.280 5.520 25.810 5.690 ;
        RECT 27.090 5.420 27.290 5.770 ;
        RECT 27.090 5.390 27.300 5.420 ;
        RECT 3.350 4.960 3.970 5.080 ;
        RECT 3.350 4.910 3.890 4.960 ;
        RECT 4.240 4.910 5.050 5.080 ;
        RECT 1.160 4.600 1.370 4.630 ;
        RECT 1.170 4.250 1.370 4.600 ;
        RECT 3.350 4.570 3.540 4.680 ;
        RECT 4.240 4.570 4.430 4.910 ;
        RECT 2.650 4.330 3.180 4.500 ;
        RECT 3.350 4.450 4.430 4.570 ;
        RECT 3.470 4.390 4.430 4.450 ;
        RECT 16.600 3.960 17.150 4.390 ;
        RECT 20.230 4.150 20.460 4.840 ;
        RECT 25.530 4.610 25.700 5.130 ;
        RECT 25.370 4.350 25.700 4.610 ;
        RECT 19.200 3.210 19.390 3.530 ;
        RECT 25.530 3.440 25.700 4.350 ;
        RECT 26.360 3.530 26.530 5.140 ;
        RECT 27.080 4.810 27.300 5.390 ;
        RECT 31.450 5.410 31.620 5.450 ;
        RECT 31.860 5.410 32.060 5.440 ;
        RECT 29.070 5.220 29.150 5.360 ;
        RECT 29.060 5.180 29.380 5.220 ;
        RECT 29.050 4.990 29.380 5.180 ;
        RECT 31.450 5.150 32.060 5.410 ;
        RECT 31.450 5.120 31.620 5.150 ;
        RECT 31.860 5.110 32.060 5.150 ;
        RECT 32.450 5.110 32.820 6.100 ;
        RECT 29.060 4.960 29.380 4.990 ;
        RECT 27.090 4.800 27.300 4.810 ;
        RECT 27.970 4.660 28.290 4.690 ;
        RECT 26.730 4.630 26.920 4.640 ;
        RECT 26.730 4.340 26.930 4.630 ;
        RECT 27.970 4.470 28.300 4.660 ;
        RECT 31.450 4.560 31.620 4.590 ;
        RECT 31.860 4.560 32.060 4.600 ;
        RECT 27.970 4.430 28.290 4.470 ;
        RECT 26.720 4.010 27.010 4.340 ;
        RECT 31.450 4.300 32.060 4.560 ;
        RECT 31.450 4.260 31.620 4.300 ;
        RECT 31.860 4.270 32.060 4.300 ;
        RECT 31.860 3.910 32.060 3.940 ;
        RECT 31.630 3.650 32.060 3.910 ;
        RECT 26.360 3.340 26.540 3.530 ;
        RECT 19.110 3.120 19.390 3.210 ;
        RECT 19.110 2.980 22.750 3.120 ;
        RECT 19.200 2.940 22.750 2.980 ;
        RECT 16.600 2.230 17.150 2.660 ;
        RECT 19.200 2.520 19.390 2.940 ;
        RECT 20.230 1.210 20.460 1.940 ;
        RECT 25.530 1.850 25.700 2.710 ;
        RECT 25.370 1.590 25.700 1.850 ;
        RECT 25.530 1.020 25.700 1.590 ;
        RECT 26.360 2.620 26.540 2.810 ;
        RECT 26.360 1.010 26.530 2.620 ;
        RECT 28.090 2.560 28.270 3.620 ;
        RECT 31.860 3.610 32.060 3.650 ;
        RECT 32.450 3.610 32.820 4.600 ;
        RECT 28.700 3.380 29.020 3.410 ;
        RECT 28.700 3.190 29.030 3.380 ;
        RECT 28.700 3.150 29.020 3.190 ;
        RECT 28.700 3.070 28.870 3.150 ;
        RECT 28.650 2.900 28.870 3.070 ;
        RECT 31.860 3.060 32.060 3.100 ;
        RECT 28.650 2.740 28.820 2.900 ;
        RECT 31.630 2.800 32.060 3.060 ;
        RECT 31.860 2.770 32.060 2.800 ;
        RECT 29.140 2.400 29.220 2.480 ;
        RECT 29.280 2.400 29.470 2.520 ;
        RECT 29.140 2.310 29.470 2.400 ;
        RECT 29.280 2.290 29.470 2.310 ;
        RECT 31.450 2.410 31.620 2.450 ;
        RECT 31.860 2.410 32.060 2.440 ;
        RECT 31.450 2.150 32.060 2.410 ;
        RECT 26.720 1.810 27.010 2.140 ;
        RECT 31.450 2.120 31.620 2.150 ;
        RECT 31.860 2.110 32.060 2.150 ;
        RECT 32.450 2.110 32.820 3.100 ;
        RECT 26.730 1.520 26.930 1.810 ;
        RECT 31.450 1.560 31.620 1.590 ;
        RECT 31.860 1.560 32.060 1.600 ;
        RECT 26.730 1.510 26.920 1.520 ;
        RECT 27.090 1.340 27.300 1.350 ;
        RECT 27.080 0.760 27.300 1.340 ;
        RECT 31.450 1.300 32.060 1.560 ;
        RECT 31.450 1.260 31.620 1.300 ;
        RECT 31.860 1.270 32.060 1.300 ;
        RECT 31.720 0.940 31.900 1.180 ;
        RECT 31.720 0.910 32.060 0.940 ;
        RECT 27.090 0.730 27.300 0.760 ;
        RECT 25.280 0.460 25.810 0.630 ;
        RECT 27.090 0.380 27.290 0.730 ;
        RECT 31.630 0.650 32.060 0.910 ;
        RECT 31.720 0.610 32.060 0.650 ;
        RECT 32.450 0.610 32.820 1.600 ;
        RECT 31.720 0.000 31.900 0.610 ;
        RECT 32.530 0.000 32.700 0.610 ;
      LAYER mcon ;
        RECT 3.000 9.390 3.180 9.560 ;
        RECT 3.330 9.450 3.500 9.620 ;
        RECT 1.190 9.090 1.360 9.260 ;
        RECT 1.540 8.250 1.720 8.440 ;
        RECT 3.800 8.890 3.970 9.060 ;
        RECT 6.140 8.510 6.310 8.680 ;
        RECT 6.140 8.060 6.310 8.230 ;
        RECT 2.620 7.690 2.790 7.860 ;
        RECT 11.590 7.910 11.860 8.180 ;
        RECT 3.330 7.460 3.500 7.630 ;
        RECT 1.540 5.450 1.720 5.640 ;
        RECT 3.340 6.390 3.510 6.560 ;
        RECT 3.800 6.570 3.970 6.740 ;
        RECT 9.170 6.880 9.340 7.050 ;
        RECT 2.610 6.000 2.780 6.170 ;
        RECT 11.590 6.180 11.860 6.450 ;
        RECT 29.000 5.830 29.170 6.000 ;
        RECT 31.690 5.840 31.860 6.010 ;
        RECT 6.140 5.560 6.310 5.730 ;
        RECT 32.770 5.600 32.820 5.770 ;
        RECT 3.790 4.990 3.960 5.160 ;
        RECT 6.140 5.110 6.310 5.280 ;
        RECT 27.100 5.220 27.270 5.390 ;
        RECT 1.190 4.630 1.360 4.800 ;
        RECT 3.000 4.330 3.180 4.500 ;
        RECT 3.360 4.480 3.530 4.650 ;
        RECT 20.260 4.640 20.430 4.810 ;
        RECT 16.600 4.040 16.870 4.310 ;
        RECT 20.260 4.190 20.430 4.360 ;
        RECT 25.430 4.390 25.600 4.560 ;
        RECT 29.150 5.000 29.320 5.170 ;
        RECT 31.640 5.190 31.810 5.360 ;
        RECT 26.740 4.380 26.920 4.570 ;
        RECT 28.030 4.480 28.200 4.650 ;
        RECT 31.640 4.350 31.810 4.520 ;
        RECT 32.770 3.940 32.820 4.110 ;
        RECT 31.690 3.700 31.860 3.870 ;
        RECT 19.120 3.010 19.290 3.180 ;
        RECT 16.600 2.310 16.870 2.580 ;
        RECT 20.260 1.690 20.430 1.860 ;
        RECT 25.430 1.630 25.600 1.800 ;
        RECT 20.260 1.240 20.430 1.410 ;
        RECT 28.760 3.200 28.930 3.370 ;
        RECT 31.690 2.840 31.860 3.010 ;
        RECT 32.770 2.600 32.820 2.770 ;
        RECT 29.290 2.320 29.460 2.490 ;
        RECT 31.640 2.190 31.810 2.360 ;
        RECT 26.740 1.580 26.920 1.770 ;
        RECT 31.640 1.350 31.810 1.520 ;
        RECT 27.100 0.760 27.270 0.930 ;
        RECT 32.770 0.940 32.820 1.110 ;
        RECT 31.690 0.700 31.860 0.870 ;
      LAYER met1 ;
        RECT 1.130 9.320 1.290 9.970 ;
        RECT 1.130 8.770 1.400 9.320 ;
        RECT 1.120 8.720 1.400 8.770 ;
        RECT 1.120 8.630 1.290 8.720 ;
        RECT 1.130 5.260 1.290 8.630 ;
        RECT 1.540 8.510 1.730 9.970 ;
        RECT 3.410 9.680 3.620 9.970 ;
        RECT 2.940 9.150 3.250 9.590 ;
        RECT 3.300 9.390 3.620 9.680 ;
        RECT 1.510 8.480 1.730 8.510 ;
        RECT 1.500 8.210 1.750 8.480 ;
        RECT 1.500 8.200 1.740 8.210 ;
        RECT 1.510 7.960 1.740 8.200 ;
        RECT 1.540 5.930 1.700 7.960 ;
        RECT 2.540 7.620 2.860 7.940 ;
        RECT 3.410 7.690 3.620 9.390 ;
        RECT 3.880 9.120 4.070 9.970 ;
        RECT 3.770 8.830 4.070 9.120 ;
        RECT 1.890 7.110 2.130 7.530 ;
        RECT 3.300 7.400 3.620 7.690 ;
        RECT 3.410 7.180 3.620 7.400 ;
        RECT 1.860 6.790 2.130 7.110 ;
        RECT 3.880 6.800 4.070 8.830 ;
        RECT 4.290 7.510 4.500 9.970 ;
        RECT 6.090 7.970 6.350 8.760 ;
        RECT 4.170 7.000 4.500 7.510 ;
        RECT 1.890 6.360 2.130 6.790 ;
        RECT 3.430 6.620 3.620 6.670 ;
        RECT 3.310 6.330 3.620 6.620 ;
        RECT 3.770 6.510 4.070 6.800 ;
        RECT 2.530 5.930 2.850 6.250 ;
        RECT 1.510 5.690 1.740 5.930 ;
        RECT 1.500 5.680 1.740 5.690 ;
        RECT 1.500 5.410 1.750 5.680 ;
        RECT 1.510 5.380 1.730 5.410 ;
        RECT 1.120 5.170 1.290 5.260 ;
        RECT 1.120 5.120 1.400 5.170 ;
        RECT 1.130 4.570 1.400 5.120 ;
        RECT 1.130 3.920 1.290 4.570 ;
        RECT 1.540 3.920 1.730 5.380 ;
        RECT 2.940 4.300 3.250 4.740 ;
        RECT 3.430 4.710 3.620 6.330 ;
        RECT 3.880 5.220 4.070 6.510 ;
        RECT 3.760 4.930 4.070 5.220 ;
        RECT 3.330 4.420 3.620 4.710 ;
        RECT 3.420 3.920 3.650 4.420 ;
        RECT 3.880 3.920 4.070 4.930 ;
        RECT 4.290 3.920 4.500 7.000 ;
        RECT 5.080 6.080 5.240 6.100 ;
        RECT 4.920 5.780 5.240 6.080 ;
        RECT 6.090 5.030 6.350 5.820 ;
        RECT 11.530 3.920 11.950 9.970 ;
        RECT 18.990 3.240 19.220 6.100 ;
        RECT 31.520 6.090 31.800 6.100 ;
        RECT 28.920 5.760 29.240 6.080 ;
        RECT 31.520 5.950 31.940 6.090 ;
        RECT 31.620 5.770 31.940 5.950 ;
        RECT 25.210 5.280 25.520 5.720 ;
        RECT 29.070 4.930 29.390 5.250 ;
        RECT 31.570 5.120 31.890 5.440 ;
        RECT 25.360 4.320 25.680 4.640 ;
        RECT 27.960 4.400 28.280 4.720 ;
        RECT 29.180 4.240 29.390 4.350 ;
        RECT 31.570 4.270 31.890 4.590 ;
        RECT 29.160 3.920 29.420 4.240 ;
        RECT 26.330 3.530 26.570 3.660 ;
        RECT 18.990 2.950 19.320 3.240 ;
        RECT 26.330 3.210 26.590 3.530 ;
        RECT 28.690 3.120 29.010 3.440 ;
        RECT 18.990 0.400 19.220 2.950 ;
        RECT 26.330 2.610 26.590 2.930 ;
        RECT 26.330 2.490 26.570 2.610 ;
        RECT 29.180 2.580 29.390 3.920 ;
        RECT 31.620 3.620 31.940 3.940 ;
        RECT 31.620 2.770 31.940 3.090 ;
        RECT 29.260 2.260 29.490 2.550 ;
        RECT 31.570 2.120 31.890 2.440 ;
        RECT 25.360 1.560 25.680 1.880 ;
        RECT 31.570 1.270 31.890 1.590 ;
        RECT 25.210 0.430 25.520 0.870 ;
        RECT 31.620 0.620 31.940 0.940 ;
        RECT 13.140 0.100 13.460 0.400 ;
        RECT 18.940 0.100 19.260 0.400 ;
        RECT 29.330 0.250 29.650 0.550 ;
        RECT 32.580 0.500 32.820 6.220 ;
        RECT 29.330 0.220 29.760 0.250 ;
        RECT 30.360 0.240 30.870 0.250 ;
        RECT 30.360 0.220 31.200 0.240 ;
        RECT 29.330 0.190 31.200 0.220 ;
        RECT 29.480 0.140 31.200 0.190 ;
        RECT 29.510 0.110 31.200 0.140 ;
        RECT 18.990 0.050 19.220 0.100 ;
        RECT 29.540 0.090 31.200 0.110 ;
        RECT 29.610 0.080 30.570 0.090 ;
        RECT 30.860 0.050 31.200 0.090 ;
      LAYER via ;
        RECT 2.960 9.180 3.220 9.440 ;
        RECT 2.570 7.650 2.830 7.910 ;
        RECT 1.860 6.820 2.120 7.080 ;
        RECT 2.560 5.960 2.820 6.220 ;
        RECT 2.960 4.450 3.220 4.710 ;
        RECT 4.950 5.800 5.210 6.060 ;
        RECT 28.950 5.790 29.210 6.050 ;
        RECT 31.650 5.800 31.910 6.060 ;
        RECT 25.240 5.310 25.500 5.570 ;
        RECT 29.100 4.960 29.360 5.220 ;
        RECT 31.600 5.150 31.860 5.410 ;
        RECT 25.390 4.350 25.650 4.610 ;
        RECT 27.990 4.430 28.250 4.690 ;
        RECT 31.600 4.300 31.860 4.560 ;
        RECT 29.160 3.950 29.420 4.210 ;
        RECT 26.330 3.240 26.590 3.500 ;
        RECT 28.720 3.150 28.980 3.410 ;
        RECT 26.330 2.640 26.590 2.900 ;
        RECT 31.650 3.650 31.910 3.910 ;
        RECT 31.650 2.800 31.910 3.060 ;
        RECT 31.600 2.150 31.860 2.410 ;
        RECT 25.390 1.590 25.650 1.850 ;
        RECT 31.600 1.300 31.860 1.560 ;
        RECT 25.240 0.580 25.500 0.840 ;
        RECT 31.650 0.650 31.910 0.910 ;
        RECT 13.170 0.120 13.430 0.380 ;
        RECT 18.970 0.120 19.230 0.380 ;
        RECT 29.360 0.270 29.620 0.530 ;
      LAYER met2 ;
        RECT 3.180 9.480 3.500 9.490 ;
        RECT 2.940 9.470 3.500 9.480 ;
        RECT 0.770 9.290 12.290 9.470 ;
        RECT 2.940 9.150 3.250 9.290 ;
        RECT 2.550 7.930 2.860 7.950 ;
        RECT 2.550 7.740 12.290 7.930 ;
        RECT 2.550 7.620 2.860 7.740 ;
        RECT 1.830 7.050 2.150 7.080 ;
        RECT 1.830 6.820 12.290 7.050 ;
        RECT 25.210 5.600 25.520 5.610 ;
        RECT 16.160 5.420 27.690 5.600 ;
        RECT 25.210 5.280 25.520 5.420 ;
        RECT 31.570 5.370 31.880 5.450 ;
        RECT 29.080 5.220 29.390 5.260 ;
        RECT 28.900 4.970 29.620 5.220 ;
        RECT 31.270 5.160 31.880 5.370 ;
        RECT 31.570 5.120 31.880 5.160 ;
        RECT 29.080 4.930 29.620 4.970 ;
        RECT 29.350 4.860 29.620 4.930 ;
        RECT 2.940 4.600 3.250 4.740 ;
        RECT 0.770 4.590 3.250 4.600 ;
        RECT 0.770 4.440 12.290 4.590 ;
        RECT 25.360 4.580 25.670 4.650 ;
        RECT 27.960 4.580 28.270 4.720 ;
        RECT 0.770 4.420 3.250 4.440 ;
        RECT 2.940 4.410 3.250 4.420 ;
        RECT 25.360 4.390 28.270 4.580 ;
        RECT 31.570 4.550 31.880 4.590 ;
        RECT 25.360 4.360 27.960 4.390 ;
        RECT 25.360 4.320 25.670 4.360 ;
        RECT 31.270 4.340 31.880 4.550 ;
        RECT 29.420 4.290 29.620 4.300 ;
        RECT 29.420 4.210 29.640 4.290 ;
        RECT 31.570 4.260 31.880 4.340 ;
        RECT 29.130 4.190 29.640 4.210 ;
        RECT 16.230 3.870 24.220 4.070 ;
        RECT 29.080 3.950 29.640 4.190 ;
        RECT 29.080 3.940 29.550 3.950 ;
        RECT 22.820 3.190 23.040 3.200 ;
        RECT 16.240 2.940 23.070 3.190 ;
        RECT 24.000 3.150 24.220 3.870 ;
        RECT 31.620 3.880 31.930 3.940 ;
        RECT 31.620 3.650 32.820 3.880 ;
        RECT 31.620 3.610 31.930 3.650 ;
        RECT 16.240 2.020 19.750 2.210 ;
        RECT 19.520 1.420 19.750 2.020 ;
        RECT 22.780 1.770 23.070 2.940 ;
        RECT 23.970 3.110 24.220 3.150 ;
        RECT 23.970 2.470 24.230 3.110 ;
        RECT 31.620 3.050 31.930 3.100 ;
        RECT 31.620 2.830 32.820 3.050 ;
        RECT 31.620 2.770 31.930 2.830 ;
        RECT 23.970 2.260 28.100 2.470 ;
        RECT 31.570 2.370 31.880 2.450 ;
        RECT 27.890 2.120 28.100 2.260 ;
        RECT 31.270 2.160 31.880 2.370 ;
        RECT 31.570 2.120 31.880 2.160 ;
        RECT 27.890 1.910 29.900 2.120 ;
        RECT 25.360 1.820 25.670 1.890 ;
        RECT 25.360 1.770 27.690 1.820 ;
        RECT 22.780 1.610 27.690 1.770 ;
        RECT 22.780 1.550 25.670 1.610 ;
        RECT 31.570 1.550 31.880 1.590 ;
        RECT 22.780 1.540 23.070 1.550 ;
        RECT 19.520 1.270 19.740 1.420 ;
        RECT 31.270 1.340 31.880 1.550 ;
        RECT 23.890 1.270 29.890 1.320 ;
        RECT 19.520 1.120 29.890 1.270 ;
        RECT 31.570 1.260 31.880 1.340 ;
        RECT 19.520 1.110 29.760 1.120 ;
        RECT 19.520 1.050 24.280 1.110 ;
        RECT 31.620 0.890 31.930 0.940 ;
        RECT 25.210 0.730 25.520 0.870 ;
        RECT 25.210 0.720 27.690 0.730 ;
        RECT 16.160 0.570 27.690 0.720 ;
        RECT 31.620 0.660 32.820 0.890 ;
        RECT 31.620 0.610 31.930 0.660 ;
        RECT 25.210 0.550 27.690 0.570 ;
        RECT 25.210 0.540 25.520 0.550 ;
  END
END sky130_hilas_TA2Cell_1FG_Strong

MACRO sky130_hilas_TA2Cell_NoFG
  CLASS CORE ;
  FOREIGN sky130_hilas_TA2Cell_NoFG ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 10.100 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN COLSEL1
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT 10.570 4.640 10.760 6.100 ;
        RECT 10.570 4.610 10.790 4.640 ;
        RECT 10.550 4.340 10.800 4.610 ;
        RECT 10.560 4.330 10.800 4.340 ;
        RECT 10.560 4.090 10.790 4.330 ;
        RECT 10.600 2.060 10.760 4.090 ;
        RECT 10.560 1.820 10.790 2.060 ;
        RECT 10.560 1.810 10.800 1.820 ;
        RECT 10.550 1.540 10.800 1.810 ;
        RECT 10.570 1.510 10.790 1.540 ;
        RECT 10.570 0.050 10.760 1.510 ;
    END
  END COLSEL1
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 12.470 0.320 12.780 0.390 ;
        RECT 11.870 0.070 12.780 0.320 ;
        RECT 12.470 0.060 12.780 0.070 ;
    END
  END VIN12
  PIN VIN21
    PORT
      LAYER met2 ;
        RECT 13.790 3.400 14.100 3.440 ;
        RECT 13.700 3.390 14.130 3.400 ;
        RECT 13.470 3.160 14.570 3.390 ;
        RECT 13.790 3.110 14.100 3.160 ;
    END
  END VIN21
  PIN VIN22
    PORT
      LAYER met2 ;
        RECT 13.430 6.080 13.680 6.090 ;
        RECT 14.030 6.080 14.340 6.090 ;
        RECT 13.430 5.830 14.340 6.080 ;
        RECT 14.030 5.760 14.340 5.830 ;
    END
  END VIN22
  PIN OUTPUT1
    ANTENNADIFFAREA 0.308800 ;
    PORT
      LAYER met2 ;
        RECT 15.000 2.790 15.310 2.840 ;
        RECT 17.290 2.790 17.600 2.920 ;
        RECT 15.000 2.570 17.920 2.790 ;
        RECT 15.000 2.510 15.310 2.570 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    ANTENNADIFFAREA 0.308800 ;
    PORT
      LAYER met2 ;
        RECT 15.000 3.620 15.310 3.680 ;
        RECT 17.300 3.620 17.610 3.640 ;
        RECT 15.000 3.390 17.920 3.620 ;
        RECT 15.000 3.350 15.310 3.390 ;
        RECT 17.300 3.310 17.610 3.390 ;
    END
  END OUTPUT2
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 15.960 4.650 16.300 4.740 ;
        RECT 13.610 4.460 16.300 4.650 ;
        RECT 13.610 3.890 13.800 4.460 ;
        RECT 15.960 4.410 16.300 4.460 ;
        RECT 2.820 3.700 13.800 3.890 ;
        RECT 2.820 3.520 3.010 3.700 ;
        RECT 2.800 2.530 3.150 3.520 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.960 0.050 16.300 6.100 ;
      LAYER via ;
        RECT 16.000 4.440 16.260 4.700 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 14.850 6.100 16.710 7.490 ;
        RECT 14.850 5.960 17.920 6.100 ;
        RECT 14.520 4.500 17.920 5.960 ;
        RECT 14.520 4.060 16.250 4.500 ;
        RECT 16.640 1.650 17.920 4.500 ;
        RECT 16.410 0.000 17.920 1.650 ;
      LAYER met2 ;
        RECT 15.000 5.760 15.310 5.840 ;
        RECT 17.250 5.760 17.560 5.860 ;
        RECT 15.000 5.530 17.560 5.760 ;
        RECT 15.000 5.510 15.310 5.530 ;
        RECT 14.180 5.220 14.490 5.260 ;
        RECT 14.000 5.110 14.740 5.220 ;
        RECT 14.950 5.110 15.260 5.190 ;
        RECT 14.000 4.970 15.260 5.110 ;
        RECT 14.180 4.930 15.260 4.970 ;
        RECT 14.490 4.900 15.260 4.930 ;
        RECT 14.490 4.850 14.740 4.900 ;
        RECT 14.950 4.860 15.260 4.900 ;
    END
    PORT
      LAYER met1 ;
        RECT 16.630 4.520 16.900 6.100 ;
        RECT 16.630 4.230 16.910 4.520 ;
        RECT 16.630 1.930 16.900 4.230 ;
        RECT 16.630 1.640 16.910 1.930 ;
        RECT 16.630 0.050 16.900 1.640 ;
    END
  END VPWR
  PIN DRAIN1
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 9.050 5.600 9.360 5.610 ;
        RECT 0.000 5.420 11.530 5.600 ;
        RECT 9.050 5.280 9.360 5.420 ;
    END
  END DRAIN1
  PIN DRAIN2
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 9.050 0.730 9.360 0.870 ;
        RECT 9.050 0.720 11.530 0.730 ;
        RECT 0.000 0.570 11.530 0.720 ;
        RECT 9.050 0.550 11.530 0.570 ;
        RECT 9.050 0.540 9.360 0.550 ;
    END
  END DRAIN2
  PIN VTUN
    ANTENNADIFFAREA 1.808400 ;
    PORT
      LAYER nwell ;
        RECT 0.020 1.780 1.750 5.350 ;
        RECT 0.590 1.450 1.150 1.780 ;
      LAYER met1 ;
        RECT 0.350 0.050 0.770 6.100 ;
    END
  END VTUN
  PIN GATE1
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT 3.770 3.710 6.490 5.360 ;
        RECT 3.770 3.670 6.480 3.710 ;
        RECT 3.770 2.340 6.480 2.380 ;
        RECT 3.770 0.690 6.490 2.340 ;
      LAYER met1 ;
        RECT 4.050 4.890 4.280 6.100 ;
        RECT 4.050 4.100 4.310 4.890 ;
        RECT 4.050 1.950 4.280 4.100 ;
        RECT 4.050 1.160 4.310 1.950 ;
        RECT 4.050 0.050 4.280 1.160 ;
    END
  END GATE1
  PIN VINJ
    ANTENNADIFFAREA 1.574400 ;
    PORT
      LAYER nwell ;
        RECT 8.220 4.580 11.530 6.150 ;
        RECT 8.220 4.360 13.110 4.580 ;
        RECT 8.220 3.120 11.530 4.360 ;
        RECT 8.220 3.100 13.080 3.120 ;
        RECT 8.220 3.050 14.640 3.100 ;
        RECT 8.220 0.000 11.530 3.050 ;
        RECT 12.780 3.030 14.640 3.050 ;
      LAYER met2 ;
        RECT 10.140 3.240 10.460 3.500 ;
        RECT 10.180 3.220 11.360 3.240 ;
        RECT 10.180 2.960 11.400 3.220 ;
        RECT 10.180 2.900 11.360 2.960 ;
        RECT 10.140 2.890 11.360 2.900 ;
        RECT 10.140 2.640 10.460 2.890 ;
    END
  END VINJ
  PIN VIN11
    PORT
      LAYER met2 ;
        RECT 12.230 2.990 12.540 3.040 ;
        RECT 11.910 2.760 13.010 2.990 ;
        RECT 11.910 2.750 12.570 2.760 ;
        RECT 12.230 2.710 12.540 2.750 ;
    END
  END VIN11
  OBS
      LAYER nwell ;
        RECT 14.520 8.200 16.710 10.100 ;
        RECT 14.850 7.550 16.710 8.200 ;
        RECT 14.120 3.160 14.570 3.390 ;
        RECT 11.910 2.750 12.190 2.990 ;
        RECT 12.560 2.760 13.010 2.990 ;
      LAYER li1 ;
        RECT 15.260 8.020 15.440 10.070 ;
        RECT 16.070 8.280 16.240 10.060 ;
        RECT 15.990 8.110 16.320 8.280 ;
        RECT 13.770 6.050 13.940 6.100 ;
        RECT 13.770 5.790 14.330 6.050 ;
        RECT 15.260 5.840 15.440 7.020 ;
        RECT 16.070 5.840 16.240 7.010 ;
        RECT 15.240 5.800 15.440 5.840 ;
        RECT 13.770 5.770 13.940 5.790 ;
        RECT 9.120 5.520 9.650 5.690 ;
        RECT 10.930 5.420 11.130 5.770 ;
        RECT 15.010 5.540 15.440 5.800 ;
        RECT 15.240 5.510 15.440 5.540 ;
        RECT 10.930 5.390 11.140 5.420 ;
        RECT 0.440 3.960 0.990 4.390 ;
        RECT 4.070 4.150 4.300 4.840 ;
        RECT 9.370 4.610 9.540 5.130 ;
        RECT 9.210 4.350 9.540 4.610 ;
        RECT 2.830 3.120 3.290 3.530 ;
        RECT 9.370 3.440 9.540 4.350 ;
        RECT 10.200 3.530 10.370 5.140 ;
        RECT 10.920 4.810 11.140 5.390 ;
        RECT 14.170 5.220 14.250 5.360 ;
        RECT 14.160 5.180 14.480 5.220 ;
        RECT 14.150 4.990 14.480 5.180 ;
        RECT 14.160 4.960 14.480 4.990 ;
        RECT 14.830 5.150 15.000 5.190 ;
        RECT 15.260 5.180 15.440 5.510 ;
        RECT 15.240 5.150 15.440 5.180 ;
        RECT 14.830 4.890 15.440 5.150 ;
        RECT 14.830 4.860 15.000 4.890 ;
        RECT 15.240 4.850 15.440 4.890 ;
        RECT 15.830 4.850 16.380 5.840 ;
        RECT 17.200 5.690 17.830 5.860 ;
        RECT 17.200 5.590 17.590 5.690 ;
        RECT 17.200 5.560 17.580 5.590 ;
        RECT 17.200 5.410 17.560 5.560 ;
        RECT 16.850 5.240 17.560 5.410 ;
        RECT 10.930 4.800 11.140 4.810 ;
        RECT 13.070 4.660 13.390 4.690 ;
        RECT 10.570 4.630 10.760 4.640 ;
        RECT 10.570 4.340 10.770 4.630 ;
        RECT 13.070 4.470 13.400 4.660 ;
        RECT 16.850 4.490 17.550 4.800 ;
        RECT 13.070 4.430 13.390 4.470 ;
        RECT 10.560 4.010 10.850 4.340 ;
        RECT 14.830 4.300 15.000 4.330 ;
        RECT 15.240 4.300 15.440 4.340 ;
        RECT 14.830 4.040 15.440 4.300 ;
        RECT 14.830 4.000 15.000 4.040 ;
        RECT 15.240 4.010 15.440 4.040 ;
        RECT 12.680 3.780 12.900 3.840 ;
        RECT 12.680 3.670 12.910 3.780 ;
        RECT 10.200 3.340 10.380 3.530 ;
        RECT 2.830 2.940 6.590 3.120 ;
        RECT 0.440 2.230 0.990 2.660 ;
        RECT 2.830 2.520 3.290 2.940 ;
        RECT 4.070 1.210 4.300 1.940 ;
        RECT 9.370 1.850 9.540 2.710 ;
        RECT 9.210 1.590 9.540 1.850 ;
        RECT 9.370 1.020 9.540 1.590 ;
        RECT 10.200 2.620 10.380 2.810 ;
        RECT 10.200 1.010 10.370 2.620 ;
        RECT 11.630 2.530 11.810 3.590 ;
        RECT 12.720 3.550 12.910 3.670 ;
        RECT 15.240 3.650 15.440 3.680 ;
        RECT 12.190 3.250 12.360 3.410 ;
        RECT 12.190 3.080 12.410 3.250 ;
        RECT 12.240 3.000 12.410 3.080 ;
        RECT 12.240 2.960 12.560 3.000 ;
        RECT 12.240 2.770 12.570 2.960 ;
        RECT 12.240 2.740 12.560 2.770 ;
        RECT 13.190 2.560 13.370 3.620 ;
        RECT 13.800 3.380 14.120 3.410 ;
        RECT 15.010 3.390 15.440 3.650 ;
        RECT 13.800 3.190 14.130 3.380 ;
        RECT 15.240 3.350 15.440 3.390 ;
        RECT 15.830 3.350 16.380 4.340 ;
        RECT 16.700 4.260 17.550 4.490 ;
        RECT 16.850 3.920 17.550 4.260 ;
        RECT 17.310 3.560 17.630 3.600 ;
        RECT 17.310 3.500 17.640 3.560 ;
        RECT 16.840 3.370 17.640 3.500 ;
        RECT 16.840 3.340 17.630 3.370 ;
        RECT 16.840 3.320 17.540 3.340 ;
        RECT 13.800 3.150 14.120 3.190 ;
        RECT 13.800 3.070 13.970 3.150 ;
        RECT 13.750 2.900 13.970 3.070 ;
        RECT 13.750 2.740 13.920 2.900 ;
        RECT 17.300 2.840 17.620 2.880 ;
        RECT 15.240 2.800 15.440 2.840 ;
        RECT 14.280 2.480 14.470 2.600 ;
        RECT 15.010 2.540 15.440 2.800 ;
        RECT 15.240 2.510 15.440 2.540 ;
        RECT 14.240 2.370 14.470 2.480 ;
        RECT 14.240 2.310 14.460 2.370 ;
        RECT 14.830 2.150 15.000 2.190 ;
        RECT 15.240 2.150 15.440 2.180 ;
        RECT 10.560 1.810 10.850 2.140 ;
        RECT 14.830 1.890 15.440 2.150 ;
        RECT 14.830 1.860 15.000 1.890 ;
        RECT 15.240 1.850 15.440 1.890 ;
        RECT 15.830 1.850 16.380 2.840 ;
        RECT 16.840 2.660 17.630 2.840 ;
        RECT 17.300 2.650 17.630 2.660 ;
        RECT 17.300 2.620 17.620 2.650 ;
        RECT 16.850 1.900 17.550 2.240 ;
        RECT 10.570 1.520 10.770 1.810 ;
        RECT 11.510 1.680 11.830 1.720 ;
        RECT 10.570 1.510 10.760 1.520 ;
        RECT 11.510 1.490 11.840 1.680 ;
        RECT 16.700 1.670 17.550 1.900 ;
        RECT 11.510 1.460 11.830 1.490 ;
        RECT 16.850 1.360 17.550 1.670 ;
        RECT 10.930 1.340 11.140 1.350 ;
        RECT 10.920 0.760 11.140 1.340 ;
        RECT 14.830 1.300 15.000 1.330 ;
        RECT 15.240 1.300 15.440 1.340 ;
        RECT 12.600 1.160 12.920 1.190 ;
        RECT 12.590 0.970 12.920 1.160 ;
        RECT 14.830 1.040 15.440 1.300 ;
        RECT 14.830 1.000 15.000 1.040 ;
        RECT 15.240 1.010 15.440 1.040 ;
        RECT 12.600 0.930 12.920 0.970 ;
        RECT 12.610 0.790 12.690 0.930 ;
        RECT 10.930 0.730 11.140 0.760 ;
        RECT 9.120 0.460 9.650 0.630 ;
        RECT 10.930 0.380 11.130 0.730 ;
        RECT 15.240 0.650 15.440 0.680 ;
        RECT 15.010 0.390 15.440 0.650 ;
        RECT 12.210 0.360 12.380 0.380 ;
        RECT 12.210 0.100 12.770 0.360 ;
        RECT 15.240 0.350 15.440 0.390 ;
        RECT 15.830 0.350 16.380 1.340 ;
        RECT 16.820 0.920 17.000 1.180 ;
        RECT 17.550 0.920 17.880 1.090 ;
        RECT 16.820 0.750 17.560 0.920 ;
        RECT 12.210 0.050 12.380 0.100 ;
        RECT 16.820 0.000 17.000 0.750 ;
        RECT 17.200 0.470 17.560 0.750 ;
        RECT 17.630 0.470 17.800 0.920 ;
        RECT 17.200 0.300 17.830 0.470 ;
        RECT 17.630 0.000 17.800 0.300 ;
      LAYER mcon ;
        RECT 14.100 5.830 14.270 6.000 ;
        RECT 15.070 5.580 15.240 5.750 ;
        RECT 10.940 5.220 11.110 5.390 ;
        RECT 4.100 4.640 4.270 4.810 ;
        RECT 0.440 4.040 0.710 4.310 ;
        RECT 4.100 4.190 4.270 4.360 ;
        RECT 9.270 4.390 9.440 4.560 ;
        RECT 14.250 5.000 14.420 5.170 ;
        RECT 15.020 4.930 15.190 5.100 ;
        RECT 16.050 5.260 16.220 5.430 ;
        RECT 17.320 5.600 17.490 5.770 ;
        RECT 10.580 4.380 10.760 4.570 ;
        RECT 13.130 4.480 13.300 4.650 ;
        RECT 15.020 4.090 15.190 4.260 ;
        RECT 16.710 4.290 16.880 4.460 ;
        RECT 2.860 3.270 3.030 3.440 ;
        RECT 2.860 2.930 3.030 3.100 ;
        RECT 0.440 2.310 0.710 2.580 ;
        RECT 2.860 2.580 3.030 2.750 ;
        RECT 4.100 1.690 4.270 1.860 ;
        RECT 9.270 1.630 9.440 1.800 ;
        RECT 4.100 1.240 4.270 1.410 ;
        RECT 12.730 3.580 12.900 3.750 ;
        RECT 16.050 3.760 16.220 3.930 ;
        RECT 12.300 2.780 12.470 2.950 ;
        RECT 15.070 3.440 15.240 3.610 ;
        RECT 13.860 3.200 14.030 3.370 ;
        RECT 17.370 3.380 17.540 3.550 ;
        RECT 14.290 2.400 14.460 2.570 ;
        RECT 15.070 2.580 15.240 2.750 ;
        RECT 17.360 2.660 17.530 2.830 ;
        RECT 16.050 2.260 16.220 2.430 ;
        RECT 15.020 1.930 15.190 2.100 ;
        RECT 10.580 1.580 10.760 1.770 ;
        RECT 16.710 1.700 16.880 1.870 ;
        RECT 11.570 1.500 11.740 1.670 ;
        RECT 12.690 0.980 12.860 1.150 ;
        RECT 15.020 1.090 15.190 1.260 ;
        RECT 10.940 0.760 11.110 0.930 ;
        RECT 16.050 0.760 16.220 0.930 ;
        RECT 15.070 0.440 15.240 0.610 ;
        RECT 12.540 0.150 12.710 0.320 ;
        RECT 17.280 0.410 17.450 0.580 ;
      LAYER met1 ;
        RECT 2.830 3.530 3.060 6.100 ;
        RECT 9.050 5.280 9.360 5.720 ;
        RECT 11.010 5.450 11.290 6.100 ;
        RECT 14.020 5.760 14.340 6.080 ;
        RECT 15.000 5.510 15.320 5.830 ;
        RECT 17.250 5.530 17.570 5.850 ;
        RECT 10.900 4.850 11.290 5.450 ;
        RECT 14.170 4.930 14.490 5.250 ;
        RECT 14.950 4.860 15.270 5.180 ;
        RECT 9.200 4.320 9.520 4.640 ;
        RECT 10.170 3.530 10.410 3.660 ;
        RECT 2.790 2.520 3.170 3.530 ;
        RECT 10.170 3.210 10.430 3.530 ;
        RECT 11.010 3.250 11.290 4.850 ;
        RECT 13.060 4.400 13.380 4.720 ;
        RECT 14.280 4.240 14.490 4.350 ;
        RECT 14.260 3.920 14.520 4.240 ;
        RECT 14.950 4.010 15.270 4.330 ;
        RECT 12.700 3.520 12.930 3.810 ;
        RECT 11.010 2.930 11.370 3.250 ;
        RECT 10.170 2.610 10.430 2.930 ;
        RECT 2.830 0.050 3.060 2.520 ;
        RECT 10.170 2.490 10.410 2.610 ;
        RECT 9.200 1.560 9.520 1.880 ;
        RECT 11.010 1.300 11.290 2.930 ;
        RECT 12.230 2.710 12.550 3.030 ;
        RECT 12.720 2.230 12.930 3.520 ;
        RECT 13.790 3.120 14.110 3.440 ;
        RECT 14.280 2.630 14.490 3.920 ;
        RECT 15.000 3.360 15.320 3.680 ;
        RECT 17.300 3.310 17.620 3.630 ;
        RECT 14.260 2.340 14.490 2.630 ;
        RECT 15.000 2.510 15.320 2.830 ;
        RECT 17.290 2.590 17.610 2.910 ;
        RECT 12.700 1.910 12.960 2.230 ;
        RECT 12.720 1.800 12.930 1.910 ;
        RECT 14.950 1.860 15.270 2.180 ;
        RECT 11.500 1.430 11.820 1.750 ;
        RECT 9.050 0.430 9.360 0.870 ;
        RECT 10.900 0.700 11.290 1.300 ;
        RECT 12.610 0.900 12.930 1.220 ;
        RECT 14.950 1.010 15.270 1.330 ;
        RECT 11.010 0.050 11.290 0.700 ;
        RECT 12.460 0.070 12.780 0.390 ;
        RECT 15.000 0.360 15.320 0.680 ;
        RECT 17.210 0.340 17.530 0.660 ;
      LAYER via ;
        RECT 9.080 5.310 9.340 5.570 ;
        RECT 14.050 5.790 14.310 6.050 ;
        RECT 15.030 5.540 15.290 5.800 ;
        RECT 17.280 5.560 17.540 5.820 ;
        RECT 14.200 4.960 14.460 5.220 ;
        RECT 14.980 4.890 15.240 5.150 ;
        RECT 9.230 4.350 9.490 4.610 ;
        RECT 2.830 2.560 3.120 3.490 ;
        RECT 10.170 3.240 10.430 3.500 ;
        RECT 13.090 4.430 13.350 4.690 ;
        RECT 14.260 3.950 14.520 4.210 ;
        RECT 14.980 4.040 15.240 4.300 ;
        RECT 11.110 2.960 11.370 3.220 ;
        RECT 10.170 2.640 10.430 2.900 ;
        RECT 9.230 1.590 9.490 1.850 ;
        RECT 12.260 2.740 12.520 3.000 ;
        RECT 13.820 3.150 14.080 3.410 ;
        RECT 15.030 3.390 15.290 3.650 ;
        RECT 17.330 3.340 17.590 3.600 ;
        RECT 15.030 2.540 15.290 2.800 ;
        RECT 17.320 2.620 17.580 2.880 ;
        RECT 12.700 1.940 12.960 2.200 ;
        RECT 14.980 1.890 15.240 2.150 ;
        RECT 11.530 1.460 11.790 1.720 ;
        RECT 9.080 0.580 9.340 0.840 ;
        RECT 12.640 0.930 12.900 1.190 ;
        RECT 14.980 1.040 15.240 1.300 ;
        RECT 15.030 0.390 15.290 0.650 ;
        RECT 17.240 0.370 17.500 0.630 ;
        RECT 12.490 0.100 12.750 0.360 ;
      LAYER met2 ;
        RECT 9.200 4.580 9.510 4.650 ;
        RECT 13.060 4.580 13.370 4.720 ;
        RECT 9.200 4.390 13.370 4.580 ;
        RECT 9.200 4.360 13.110 4.390 ;
        RECT 9.200 4.320 9.510 4.360 ;
        RECT 14.950 4.290 15.260 4.330 ;
        RECT 14.520 4.210 15.260 4.290 ;
        RECT 14.230 4.190 15.260 4.210 ;
        RECT 14.180 4.080 15.260 4.190 ;
        RECT 14.180 4.000 14.730 4.080 ;
        RECT 14.950 4.000 15.260 4.080 ;
        RECT 14.180 3.940 14.650 4.000 ;
        RECT 12.620 2.120 13.090 2.210 ;
        RECT 12.620 2.110 14.730 2.120 ;
        RECT 14.950 2.110 15.260 2.190 ;
        RECT 12.620 1.960 15.260 2.110 ;
        RECT 12.670 1.940 15.260 1.960 ;
        RECT 12.960 1.920 15.260 1.940 ;
        RECT 14.650 1.900 15.260 1.920 ;
        RECT 9.200 1.820 9.510 1.890 ;
        RECT 14.950 1.860 15.260 1.900 ;
        RECT 11.390 1.820 11.550 1.830 ;
        RECT 9.200 1.760 11.550 1.820 ;
        RECT 9.200 1.610 11.810 1.760 ;
        RECT 9.200 1.560 9.510 1.610 ;
        RECT 11.390 1.430 11.810 1.610 ;
        RECT 12.670 1.290 14.730 1.320 ;
        RECT 14.950 1.290 15.260 1.330 ;
        RECT 12.670 1.220 15.260 1.290 ;
        RECT 12.620 1.180 15.260 1.220 ;
        RECT 12.440 1.110 15.260 1.180 ;
        RECT 12.440 0.930 12.990 1.110 ;
        RECT 14.650 1.080 15.260 1.110 ;
        RECT 14.950 1.000 15.260 1.080 ;
        RECT 12.620 0.890 12.930 0.930 ;
        RECT 15.000 0.630 15.310 0.680 ;
        RECT 17.210 0.630 17.520 0.670 ;
        RECT 15.000 0.400 17.710 0.630 ;
        RECT 15.000 0.350 15.310 0.400 ;
        RECT 17.210 0.340 17.520 0.400 ;
  END
END sky130_hilas_TA2Cell_NoFG

MACRO sky130_hilas_TopLevelTextStructure
  CLASS CORE ;
  FOREIGN sky130_hilas_TopLevelTextStructure ;
  ORIGIN 0.000 0.000 ;
  SIZE 130.250 BY 75.780 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DIG24 
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 65.420 30.870 65.560 30.880 ;
        RECT 65.420 30.540 65.570 30.870 ;
        RECT 65.420 30.450 66.630 30.540 ;
        RECT 65.420 30.390 66.760 30.450 ;
        RECT 65.420 30.380 69.030 30.390 ;
        RECT 73.730 30.380 74.050 30.430 ;
        RECT 65.420 30.340 74.050 30.380 ;
        RECT 66.450 30.230 74.050 30.340 ;
        RECT 66.450 30.120 66.760 30.230 ;
        RECT 68.950 30.220 74.050 30.230 ;
        RECT 73.730 30.170 74.050 30.220 ;
        RECT 73.710 20.760 130.250 21.260 ;
        RECT 128.240 0.760 130.250 20.760 ;
        RECT 128.210 0.180 130.250 0.760 ;
        RECT 128.210 0.110 130.240 0.180 ;
    END
  END DIG24 
  PIN DIG23
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 65.530 29.680 66.730 29.780 ;
        RECT 65.520 29.600 66.730 29.680 ;
        RECT 66.450 29.570 66.730 29.600 ;
        RECT 66.450 29.460 66.760 29.570 ;
        RECT 66.450 29.450 69.030 29.460 ;
        RECT 73.210 29.450 73.530 29.500 ;
        RECT 66.450 29.300 73.530 29.450 ;
        RECT 66.450 29.240 66.760 29.300 ;
        RECT 68.950 29.290 73.530 29.300 ;
        RECT 73.210 29.240 73.530 29.290 ;
        RECT 124.150 20.360 126.160 20.380 ;
        RECT 73.170 19.860 126.160 20.360 ;
        RECT 124.150 0.740 126.160 19.860 ;
        RECT 124.150 0.090 126.190 0.740 ;
        RECT 124.150 0.010 126.160 0.090 ;
    END
  END DIG23
  PIN DIG22
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 66.450 27.650 66.760 27.680 ;
        RECT 65.510 27.620 66.760 27.650 ;
        RECT 65.510 27.610 69.030 27.620 ;
        RECT 72.740 27.610 73.060 27.660 ;
        RECT 65.510 27.490 73.060 27.610 ;
        RECT 66.450 27.460 73.060 27.490 ;
        RECT 66.450 27.350 66.760 27.460 ;
        RECT 68.950 27.450 73.060 27.460 ;
        RECT 72.740 27.400 73.060 27.450 ;
        RECT 72.700 19.440 121.970 19.460 ;
        RECT 72.700 18.960 122.080 19.440 ;
        RECT 120.070 0.760 122.080 18.960 ;
        RECT 120.070 0.110 122.140 0.760 ;
        RECT 120.070 0.070 122.080 0.110 ;
    END
  END DIG22
  PIN DIG21
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 66.450 26.690 66.760 26.800 ;
        RECT 66.450 26.680 69.030 26.690 ;
        RECT 72.240 26.680 72.560 26.730 ;
        RECT 65.520 26.530 72.560 26.680 ;
        RECT 65.520 26.500 66.760 26.530 ;
        RECT 68.950 26.520 72.560 26.530 ;
        RECT 66.450 26.470 66.760 26.500 ;
        RECT 72.240 26.470 72.560 26.520 ;
        RECT 72.220 18.550 118.010 18.560 ;
        RECT 72.220 18.060 118.220 18.550 ;
        RECT 116.210 0.760 118.220 18.060 ;
        RECT 116.150 0.240 118.220 0.760 ;
        RECT 116.150 0.110 118.180 0.240 ;
    END
  END DIG21
  PIN DIG29
    ANTENNAGATEAREA 2.944600 ;
    ANTENNADIFFAREA 0.128000 ;
    PORT
      LAYER met2 ;
        RECT 106.840 10.090 107.150 10.120 ;
        RECT 107.840 10.090 108.160 10.130 ;
        RECT 106.840 9.840 108.160 10.090 ;
        RECT 106.840 5.140 107.140 9.840 ;
        RECT 107.840 9.810 108.160 9.840 ;
        RECT 107.850 8.190 108.170 8.510 ;
        RECT 107.960 6.900 108.150 8.190 ;
        RECT 107.840 6.580 108.160 6.900 ;
        RECT 107.430 5.140 107.750 5.250 ;
        RECT 106.840 4.930 107.750 5.140 ;
        RECT 106.840 4.920 107.600 4.930 ;
        RECT 106.840 3.500 107.140 4.920 ;
        RECT 107.960 3.700 108.150 6.580 ;
        RECT 106.840 3.340 107.200 3.500 ;
        RECT 107.840 3.380 108.160 3.700 ;
        RECT 106.490 1.900 106.810 1.970 ;
        RECT 106.990 1.900 107.200 3.340 ;
        RECT 107.960 1.990 108.150 3.380 ;
        RECT 106.490 1.700 107.200 1.900 ;
        RECT 106.490 1.650 106.810 1.700 ;
        RECT 106.990 0.670 107.200 1.700 ;
        RECT 107.800 1.670 108.150 1.990 ;
        RECT 107.940 1.460 108.150 1.670 ;
        RECT 107.940 1.440 112.960 1.460 ;
        RECT 107.960 1.270 112.960 1.440 ;
        RECT 112.770 0.810 112.960 1.270 ;
        RECT 108.120 0.670 110.150 0.760 ;
        RECT 112.770 0.740 113.800 0.810 ;
        RECT 106.990 0.460 110.150 0.670 ;
        RECT 108.120 0.110 110.150 0.460 ;
        RECT 112.100 0.090 114.130 0.740 ;
    END
  END DIG29
  PIN DIG27
    ANTENNAGATEAREA 1.055900 ;
    ANTENNADIFFAREA 0.060000 ;
    PORT
      LAYER met2 ;
        RECT 105.060 11.740 107.870 11.750 ;
        RECT 105.060 11.550 108.170 11.740 ;
        RECT 105.060 0.760 105.270 11.550 ;
        RECT 107.850 11.420 108.170 11.550 ;
        RECT 103.940 0.110 105.970 0.760 ;
    END
  END DIG27
  PIN DIG26
    ANTENNAGATEAREA 0.323400 ;
    ANTENNADIFFAREA 0.082200 ;
    PORT
      LAYER met2 ;
        RECT 104.090 13.300 104.290 13.310 ;
        RECT 107.850 13.300 108.170 13.350 ;
        RECT 104.090 13.150 108.170 13.300 ;
        RECT 104.090 1.580 104.290 13.150 ;
        RECT 107.850 13.030 108.170 13.150 ;
        RECT 104.080 1.440 104.290 1.580 ;
        RECT 104.090 1.230 104.290 1.440 ;
        RECT 101.860 1.030 104.290 1.230 ;
        RECT 101.860 0.760 102.060 1.030 ;
        RECT 99.860 0.460 102.060 0.760 ;
        RECT 99.860 0.110 101.890 0.460 ;
    END
  END DIG26
  PIN DIG25
    PORT
      LAYER met2 ;
        RECT 102.940 9.700 103.200 10.020 ;
        RECT 102.970 1.640 103.170 9.700 ;
        RECT 96.930 1.440 103.170 1.640 ;
        RECT 96.930 0.760 97.130 1.440 ;
        RECT 95.840 0.110 97.870 0.760 ;
    END
  END DIG25
  PIN DIG20
    PORT
      LAYER met2 ;
        RECT 100.840 47.340 101.240 47.350 ;
        RECT 100.820 47.280 101.260 47.340 ;
        RECT 100.820 47.100 104.670 47.280 ;
        RECT 100.820 47.080 105.460 47.100 ;
        RECT 100.840 47.070 101.240 47.080 ;
        RECT 104.320 46.900 105.460 47.080 ;
        RECT 100.830 4.810 101.250 4.840 ;
        RECT 91.860 4.430 101.250 4.810 ;
        RECT 91.860 0.730 93.840 4.430 ;
        RECT 100.830 4.400 101.250 4.430 ;
        RECT 91.850 0.080 93.880 0.730 ;
    END
  END DIG20
  PIN DIG19
    ANTENNAGATEAREA 43.337997 ;
    ANTENNADIFFAREA 292.456207 ;
    PORT
      LAYER nwell ;
        RECT 18.390 49.700 20.420 52.670 ;
        RECT 19.210 49.650 19.750 49.700 ;
        RECT 19.030 49.200 19.750 49.650 ;
        RECT 17.180 49.020 19.750 49.200 ;
        RECT 39.250 44.520 41.020 58.630 ;
        RECT 44.890 44.520 47.390 58.630 ;
        RECT 80.950 52.710 84.260 57.310 ;
        RECT 85.990 54.870 88.710 56.520 ;
        RECT 85.990 54.830 88.700 54.870 ;
        RECT 85.990 53.500 88.700 53.540 ;
        RECT 85.990 53.390 88.710 53.500 ;
        RECT 84.900 53.380 88.710 53.390 ;
        RECT 50.060 51.660 53.370 52.630 ;
        RECT 54.010 51.660 54.040 51.670 ;
        RECT 49.910 51.360 54.040 51.660 ;
        RECT 49.910 51.320 54.010 51.360 ;
        RECT 49.910 48.710 54.020 51.320 ;
        RECT 55.100 50.190 57.820 51.840 ;
        RECT 79.970 51.160 84.260 52.710 ;
        RECT 85.990 51.850 88.710 53.380 ;
        RECT 90.730 52.940 92.460 56.510 ;
        RECT 104.560 53.390 107.870 53.440 ;
        RECT 108.370 53.390 111.130 54.070 ;
        RECT 104.560 53.380 111.130 53.390 ;
        RECT 91.330 52.610 91.890 52.940 ;
        RECT 79.970 50.810 81.700 51.160 ;
        RECT 100.110 51.000 102.830 52.650 ;
        RECT 100.110 50.960 102.820 51.000 ;
        RECT 55.110 50.150 57.820 50.190 ;
        RECT 104.560 50.390 107.870 53.380 ;
        RECT 108.370 53.250 111.130 53.380 ;
        RECT 111.720 53.250 113.000 53.390 ;
        RECT 108.370 53.210 113.000 53.250 ;
        RECT 108.370 52.460 112.590 53.210 ;
        RECT 110.860 51.950 112.590 52.460 ;
        RECT 108.370 51.350 112.590 51.950 ;
        RECT 108.370 50.390 111.130 51.350 ;
        RECT 104.560 50.320 111.130 50.390 ;
        RECT 100.110 49.630 102.820 49.670 ;
        RECT 55.110 48.820 57.820 48.860 ;
        RECT 55.100 48.710 57.820 48.820 ;
        RECT 49.910 48.700 57.820 48.710 ;
        RECT 49.910 48.210 54.020 48.700 ;
        RECT 49.910 48.030 54.090 48.210 ;
        RECT 49.910 45.180 54.020 48.030 ;
        RECT 55.100 47.170 57.820 48.700 ;
        RECT 73.670 48.710 76.980 48.760 ;
        RECT 73.670 48.700 78.450 48.710 ;
        RECT 49.260 45.070 54.020 45.180 ;
        RECT 73.670 45.710 76.980 48.700 ;
        RECT 77.220 48.170 77.780 48.700 ;
        RECT 100.110 47.980 102.830 49.630 ;
        RECT 104.560 47.290 107.870 50.320 ;
        RECT 108.370 49.260 111.130 50.320 ;
        RECT 73.670 45.640 78.830 45.710 ;
        RECT 39.250 34.390 41.020 41.390 ;
        RECT 44.890 39.860 47.390 41.390 ;
        RECT 49.260 41.190 50.990 45.070 ;
        RECT 73.670 42.610 76.980 45.640 ;
        RECT 44.890 34.390 48.380 39.860 ;
        RECT 49.260 38.690 53.310 41.190 ;
        RECT 49.890 35.860 53.310 38.690 ;
        RECT 49.890 34.600 55.380 35.860 ;
        RECT 55.430 35.850 57.990 41.190 ;
        RECT 55.430 34.690 59.140 35.850 ;
        RECT 72.990 34.690 75.550 41.190 ;
        RECT 46.650 33.360 48.380 34.390 ;
        RECT 39.210 25.330 40.980 32.330 ;
        RECT 44.850 25.330 47.350 32.330 ;
        RECT 52.820 31.920 55.380 34.600 ;
        RECT 49.920 31.590 55.380 31.920 ;
        RECT 56.910 31.590 59.140 34.690 ;
        RECT 49.920 31.580 59.140 31.590 ;
        RECT 49.920 31.430 55.470 31.580 ;
        RECT 49.920 31.420 55.650 31.430 ;
        RECT 49.920 29.240 55.470 31.420 ;
        RECT 56.910 29.360 59.140 31.580 ;
        RECT 49.920 29.040 55.460 29.240 ;
        RECT 49.920 25.550 55.470 29.040 ;
        RECT 49.920 25.520 56.340 25.550 ;
        RECT 49.920 25.330 53.340 25.520 ;
        RECT 55.460 25.360 56.340 25.520 ;
        RECT 57.230 24.080 65.070 24.090 ;
        RECT 55.220 24.060 65.070 24.080 ;
        RECT 47.420 18.390 65.070 24.060 ;
        RECT 47.420 18.360 55.260 18.390 ;
        RECT 103.590 17.740 108.640 18.710 ;
        RECT 103.590 17.100 109.210 17.740 ;
        RECT 107.860 16.820 109.210 17.100 ;
        RECT 107.860 16.020 110.380 16.820 ;
        RECT 12.660 8.670 16.580 14.370 ;
        RECT 103.950 11.990 110.380 16.020 ;
        RECT 103.950 11.470 109.210 11.990 ;
        RECT 102.210 11.190 109.210 11.470 ;
        RECT 102.210 8.250 106.900 11.190 ;
        RECT 107.140 7.970 107.210 11.190 ;
        RECT 107.430 9.050 109.210 11.190 ;
        RECT 107.860 8.770 109.210 9.050 ;
        RECT 107.860 7.970 110.380 8.770 ;
        RECT 103.950 4.220 110.380 7.970 ;
        RECT 103.590 3.940 110.380 4.220 ;
        RECT 103.590 2.610 109.210 3.940 ;
        RECT 107.860 2.270 109.210 2.610 ;
        RECT 107.850 1.800 109.210 2.270 ;
      LAYER met3 ;
        RECT 77.230 54.870 77.680 55.620 ;
        RECT 77.230 48.710 77.600 54.870 ;
        RECT 78.270 54.860 78.720 55.610 ;
        RECT 78.350 52.220 78.720 54.860 ;
        RECT 78.350 51.620 78.790 52.220 ;
        RECT 77.230 48.380 77.720 48.710 ;
        RECT 77.280 48.220 77.720 48.380 ;
        RECT 78.350 46.510 78.720 51.620 ;
        RECT 78.340 45.640 78.810 46.510 ;
    END
  END DIG19
  PIN DIG18
    ANTENNAGATEAREA 4.609400 ;
    ANTENNADIFFAREA 8.637700 ;
    PORT
      LAYER met2 ;
        RECT 115.950 54.450 116.310 54.460 ;
        RECT 102.100 54.270 102.400 54.290 ;
        RECT 115.390 54.270 116.310 54.450 ;
        RECT 102.090 54.170 116.310 54.270 ;
        RECT 102.090 53.850 116.350 54.170 ;
        RECT 102.100 53.830 102.400 53.850 ;
        RECT 108.540 53.800 108.860 53.850 ;
        RECT 110.810 53.800 111.130 53.820 ;
        RECT 111.820 53.800 112.140 53.830 ;
        RECT 108.250 53.600 108.860 53.800 ;
        RECT 110.760 53.600 113.010 53.800 ;
        RECT 110.810 53.560 111.130 53.600 ;
        RECT 111.820 53.570 112.140 53.600 ;
        RECT 115.390 53.510 116.350 53.850 ;
        RECT 111.800 53.310 112.110 53.390 ;
        RECT 114.050 53.310 114.360 53.410 ;
        RECT 111.800 53.080 114.360 53.310 ;
        RECT 111.800 53.060 112.110 53.080 ;
        RECT 109.890 52.830 110.200 52.950 ;
        RECT 109.120 52.820 110.240 52.830 ;
        RECT 111.460 52.820 111.770 52.950 ;
        RECT 108.250 52.740 111.770 52.820 ;
        RECT 108.250 52.620 112.060 52.740 ;
        RECT 109.120 52.610 110.240 52.620 ;
        RECT 110.310 52.470 110.380 52.620 ;
        RECT 111.450 52.450 112.060 52.620 ;
        RECT 111.750 52.410 112.060 52.450 ;
        RECT 115.450 52.080 116.350 53.510 ;
        RECT 105.540 51.870 105.850 51.940 ;
        RECT 108.140 51.870 108.450 52.010 ;
        RECT 105.540 51.790 108.450 51.870 ;
        RECT 109.120 51.790 110.240 51.800 ;
        RECT 110.310 51.790 110.380 51.940 ;
        RECT 111.750 51.840 112.060 51.880 ;
        RECT 111.450 51.790 112.060 51.840 ;
        RECT 105.540 51.680 112.060 51.790 ;
        RECT 105.540 51.650 108.140 51.680 ;
        RECT 105.540 51.610 105.850 51.650 ;
        RECT 108.250 51.590 112.060 51.680 ;
        RECT 109.120 51.580 110.240 51.590 ;
        RECT 109.600 51.500 109.820 51.580 ;
        RECT 109.310 51.480 109.820 51.500 ;
        RECT 87.480 51.210 95.690 51.430 ;
        RECT 95.470 49.330 95.690 51.210 ;
        RECT 96.410 51.160 104.400 51.360 ;
        RECT 109.260 51.240 109.820 51.480 ;
        RECT 109.890 51.460 110.200 51.580 ;
        RECT 111.460 51.550 112.060 51.590 ;
        RECT 111.460 51.460 111.770 51.550 ;
        RECT 109.260 51.230 109.730 51.240 ;
        RECT 98.090 50.950 98.550 51.080 ;
        RECT 104.180 51.030 104.400 51.160 ;
        RECT 111.800 51.170 112.110 51.230 ;
        RECT 114.100 51.170 114.410 51.190 ;
        RECT 104.180 50.950 105.460 51.030 ;
        RECT 98.090 50.830 105.460 50.950 ;
        RECT 109.820 50.830 111.540 51.030 ;
        RECT 111.800 50.940 114.720 51.170 ;
        RECT 111.800 50.900 112.110 50.940 ;
        RECT 98.090 50.750 104.670 50.830 ;
        RECT 109.820 50.810 111.530 50.830 ;
        RECT 111.820 50.810 112.140 50.840 ;
        RECT 112.890 50.810 113.000 50.910 ;
        RECT 114.100 50.860 114.410 50.940 ;
        RECT 98.090 50.630 98.550 50.750 ;
        RECT 103.000 50.480 103.220 50.490 ;
        RECT 96.420 50.300 103.250 50.480 ;
        RECT 104.180 50.440 104.400 50.750 ;
        RECT 108.250 50.690 108.860 50.810 ;
        RECT 109.820 50.750 113.010 50.810 ;
        RECT 108.870 50.690 109.180 50.730 ;
        RECT 108.250 50.680 109.210 50.690 ;
        RECT 108.250 50.610 109.650 50.680 ;
        RECT 110.760 50.610 113.010 50.750 ;
        RECT 108.540 50.600 109.650 50.610 ;
        RECT 110.810 50.600 111.130 50.610 ;
        RECT 111.330 50.600 111.530 50.610 ;
        RECT 111.820 50.600 112.140 50.610 ;
        RECT 104.150 50.400 104.400 50.440 ;
        RECT 108.250 50.450 109.650 50.600 ;
        RECT 108.250 50.400 108.860 50.450 ;
        RECT 108.870 50.400 109.180 50.450 ;
        RECT 110.760 50.400 113.010 50.600 ;
        RECT 104.150 50.300 104.410 50.400 ;
        RECT 110.810 50.360 111.130 50.400 ;
        RECT 111.330 50.300 111.530 50.400 ;
        RECT 111.820 50.390 112.140 50.400 ;
        RECT 96.420 50.230 105.460 50.300 ;
        RECT 99.100 50.100 105.460 50.230 ;
        RECT 109.820 50.100 111.530 50.300 ;
        RECT 99.100 49.980 99.460 50.100 ;
        RECT 96.420 49.330 99.930 49.500 ;
        RECT 95.470 49.320 99.930 49.330 ;
        RECT 102.960 49.320 103.250 50.100 ;
        RECT 104.150 49.760 104.410 50.100 ;
        RECT 104.150 49.620 108.280 49.760 ;
        RECT 111.330 49.750 111.530 50.100 ;
        RECT 111.800 50.370 112.140 50.390 ;
        RECT 111.800 50.340 112.110 50.370 ;
        RECT 114.090 50.340 114.400 50.470 ;
        RECT 111.800 50.120 114.720 50.340 ;
        RECT 111.800 50.060 112.110 50.120 ;
        RECT 109.890 49.630 110.200 49.750 ;
        RECT 111.330 49.740 111.770 49.750 ;
        RECT 109.120 49.620 110.240 49.630 ;
        RECT 111.330 49.620 112.060 49.740 ;
        RECT 104.150 49.550 112.060 49.620 ;
        RECT 108.070 49.420 112.060 49.550 ;
        RECT 108.070 49.410 108.280 49.420 ;
        RECT 109.120 49.410 110.240 49.420 ;
        RECT 95.470 49.120 105.460 49.320 ;
        RECT 108.070 49.200 110.080 49.410 ;
        RECT 110.310 49.270 110.380 49.420 ;
        RECT 95.470 49.110 97.070 49.120 ;
        RECT 99.700 48.910 99.930 49.120 ;
        RECT 102.960 49.060 103.250 49.120 ;
        RECT 105.540 49.110 105.850 49.180 ;
        RECT 105.540 49.060 107.870 49.110 ;
        RECT 102.960 48.910 107.870 49.060 ;
        RECT 87.480 48.900 107.870 48.910 ;
        RECT 111.330 49.050 111.530 49.420 ;
        RECT 111.750 49.410 112.060 49.420 ;
        RECT 115.420 49.050 116.320 49.720 ;
        RECT 87.480 48.840 105.850 48.900 ;
        RECT 87.480 48.810 104.670 48.840 ;
        RECT 87.480 48.710 105.460 48.810 ;
        RECT 99.700 48.560 99.920 48.710 ;
        RECT 104.370 48.610 105.460 48.710 ;
        RECT 105.620 48.610 105.680 48.740 ;
        RECT 104.070 48.600 110.070 48.610 ;
        RECT 104.070 48.590 110.240 48.600 ;
        RECT 110.310 48.590 110.380 48.740 ;
        RECT 111.330 48.620 116.320 49.050 ;
        RECT 111.330 48.590 111.530 48.620 ;
        RECT 111.750 48.590 112.060 48.620 ;
        RECT 104.070 48.560 112.060 48.590 ;
        RECT 99.700 48.550 112.060 48.560 ;
        RECT 99.700 48.400 111.770 48.550 ;
        RECT 99.700 48.340 104.460 48.400 ;
        RECT 108.250 48.390 111.770 48.400 ;
        RECT 109.120 48.380 110.240 48.390 ;
        RECT 109.890 48.260 110.200 48.380 ;
        RECT 111.330 48.260 111.770 48.390 ;
        RECT 100.020 48.040 100.410 48.060 ;
        RECT 100.010 48.010 100.420 48.040 ;
        RECT 105.390 48.020 105.700 48.160 ;
        RECT 105.390 48.010 107.870 48.020 ;
        RECT 96.340 47.860 107.870 48.010 ;
        RECT 111.330 47.930 111.530 48.260 ;
        RECT 100.010 47.830 104.670 47.860 ;
        RECT 105.390 47.840 107.870 47.860 ;
        RECT 109.820 47.840 111.530 47.930 ;
        RECT 111.800 48.180 112.110 48.230 ;
        RECT 114.010 48.180 114.320 48.220 ;
        RECT 111.800 47.950 114.510 48.180 ;
        RECT 111.800 47.900 112.110 47.950 ;
        RECT 114.010 47.890 114.320 47.950 ;
        RECT 105.390 47.830 105.700 47.840 ;
        RECT 100.010 47.730 105.460 47.830 ;
        RECT 100.010 47.690 100.420 47.730 ;
        RECT 104.440 47.690 105.460 47.730 ;
        RECT 105.620 47.690 105.670 47.760 ;
        RECT 109.510 47.690 111.530 47.840 ;
        RECT 93.320 47.630 111.530 47.690 ;
        RECT 93.320 47.540 109.830 47.630 ;
        RECT 110.810 47.610 111.130 47.630 ;
        RECT 111.330 47.610 111.530 47.630 ;
        RECT 111.820 47.610 112.140 47.640 ;
        RECT 115.420 47.630 116.320 48.620 ;
        RECT 93.320 47.390 93.640 47.540 ;
        RECT 99.120 47.390 99.440 47.540 ;
        RECT 108.250 47.410 108.860 47.540 ;
        RECT 110.760 47.410 113.010 47.610 ;
        RECT 108.540 47.320 108.860 47.410 ;
        RECT 110.810 47.390 111.130 47.410 ;
        RECT 111.330 47.280 111.530 47.410 ;
        RECT 111.820 47.380 112.140 47.410 ;
        RECT 109.820 47.100 111.530 47.280 ;
        RECT 109.760 46.960 111.530 47.100 ;
        RECT 109.760 46.900 111.520 46.960 ;
        RECT 98.170 7.240 98.600 7.260 ;
        RECT 79.670 7.210 81.630 7.240 ;
        RECT 98.150 7.210 98.610 7.240 ;
        RECT 79.670 6.860 98.610 7.210 ;
        RECT 79.670 0.760 81.630 6.860 ;
        RECT 98.150 6.840 98.610 6.860 ;
        RECT 98.170 6.830 98.600 6.840 ;
        RECT 99.070 6.430 99.500 6.450 ;
        RECT 99.060 6.420 99.510 6.430 ;
        RECT 83.600 6.040 99.510 6.420 ;
        RECT 79.640 0.110 81.670 0.760 ;
        RECT 83.600 0.740 85.560 6.040 ;
        RECT 99.070 6.020 99.500 6.040 ;
        RECT 99.990 5.600 100.440 5.610 ;
        RECT 87.750 5.220 100.440 5.600 ;
        RECT 87.750 0.760 89.730 5.220 ;
        RECT 83.590 0.090 85.620 0.740 ;
        RECT 87.710 0.110 89.740 0.760 ;
    END
  END DIG18
  PIN DIG16
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 38.690 57.310 39.150 57.380 ;
        RECT 38.300 57.140 39.150 57.310 ;
        RECT 37.330 56.580 37.720 56.670 ;
        RECT 38.300 56.580 38.470 57.140 ;
        RECT 38.690 57.060 39.150 57.140 ;
        RECT 37.330 56.410 38.480 56.580 ;
        RECT 37.310 7.700 37.730 7.710 ;
        RECT 37.310 7.450 77.580 7.700 ;
        RECT 37.310 7.370 77.590 7.450 ;
        RECT 37.310 7.360 37.730 7.370 ;
        RECT 71.550 7.350 77.590 7.370 ;
        RECT 75.650 6.850 77.590 7.350 ;
        RECT 75.650 0.780 77.580 6.850 ;
        RECT 75.560 0.000 77.590 0.780 ;
    END
  END DIG16
  PIN DIG15
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 38.690 55.480 39.150 55.630 ;
        RECT 38.300 55.310 39.150 55.480 ;
        RECT 36.730 55.040 37.060 55.050 ;
        RECT 36.710 54.940 37.080 55.040 ;
        RECT 38.300 54.940 38.470 55.310 ;
        RECT 36.710 54.770 38.470 54.940 ;
        RECT 36.710 54.660 37.080 54.770 ;
        RECT 38.300 54.760 38.470 54.770 ;
        RECT 36.710 7.080 37.090 7.090 ;
        RECT 36.710 6.750 73.510 7.080 ;
        RECT 36.710 6.740 37.090 6.750 ;
        RECT 67.440 6.740 73.510 6.750 ;
        RECT 71.550 6.420 73.510 6.740 ;
        RECT 71.550 0.760 73.500 6.420 ;
        RECT 71.490 0.110 73.520 0.760 ;
    END
  END DIG15
  PIN DIG14
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 38.690 53.750 39.150 53.880 ;
        RECT 38.260 53.580 39.150 53.750 ;
        RECT 36.130 53.460 36.520 53.560 ;
        RECT 38.260 53.460 38.430 53.580 ;
        RECT 38.690 53.560 39.150 53.580 ;
        RECT 36.130 53.290 38.430 53.460 ;
        RECT 36.130 53.190 36.520 53.290 ;
        RECT 36.070 6.450 36.490 6.460 ;
        RECT 36.070 6.120 69.430 6.450 ;
        RECT 36.070 6.110 36.490 6.120 ;
        RECT 67.440 0.760 69.430 6.120 ;
        RECT 67.440 0.110 69.470 0.760 ;
    END
  END DIG14
  PIN DIG13
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 38.690 52.030 39.150 52.130 ;
        RECT 35.490 51.860 35.880 51.950 ;
        RECT 38.430 51.860 39.150 52.030 ;
        RECT 35.490 51.810 39.150 51.860 ;
        RECT 35.490 51.690 39.060 51.810 ;
        RECT 35.490 51.600 35.880 51.690 ;
        RECT 38.430 51.670 38.600 51.690 ;
        RECT 35.480 5.810 35.880 5.830 ;
        RECT 35.480 5.480 65.420 5.810 ;
        RECT 35.480 5.470 35.880 5.480 ;
        RECT 63.460 0.760 65.410 5.480 ;
        RECT 63.410 0.110 65.440 0.760 ;
    END
  END DIG13
  PIN DIG12
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 34.850 51.290 35.240 51.400 ;
        RECT 38.690 51.290 39.150 51.340 ;
        RECT 34.850 51.120 39.150 51.290 ;
        RECT 34.850 51.020 35.240 51.120 ;
        RECT 38.690 51.020 39.150 51.120 ;
        RECT 34.820 5.140 35.230 5.150 ;
        RECT 34.810 4.810 61.330 5.140 ;
        RECT 34.820 4.790 35.230 4.810 ;
        RECT 59.420 0.740 61.330 4.810 ;
        RECT 59.340 0.090 61.370 0.740 ;
    END
  END DIG12
  PIN DIG11
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 34.240 49.720 34.630 49.820 ;
        RECT 34.240 49.590 39.060 49.720 ;
        RECT 34.240 49.550 39.150 49.590 ;
        RECT 34.240 49.450 34.630 49.550 ;
        RECT 38.510 49.390 39.150 49.550 ;
        RECT 38.690 49.270 39.150 49.390 ;
        RECT 34.240 4.520 34.650 4.530 ;
        RECT 34.240 4.500 57.310 4.520 ;
        RECT 34.240 4.190 57.320 4.500 ;
        RECT 34.240 4.180 34.650 4.190 ;
        RECT 55.320 0.810 57.320 4.190 ;
        RECT 55.290 0.110 57.320 0.810 ;
    END
  END DIG11
  PIN DIG10
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 33.610 48.190 34.030 48.280 ;
        RECT 33.610 48.020 38.510 48.190 ;
        RECT 33.610 47.930 34.030 48.020 ;
        RECT 38.340 47.840 38.510 48.020 ;
        RECT 38.340 47.670 39.150 47.840 ;
        RECT 38.690 47.520 39.150 47.670 ;
        RECT 33.640 3.870 34.030 3.880 ;
        RECT 33.640 3.550 53.330 3.870 ;
        RECT 33.740 3.540 53.330 3.550 ;
        RECT 51.340 0.830 53.330 3.540 ;
        RECT 51.330 0.080 53.360 0.830 ;
    END
  END DIG10
  PIN DIG09
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 33.050 46.620 33.440 46.710 ;
        RECT 33.050 46.450 38.420 46.620 ;
        RECT 33.050 46.360 33.440 46.450 ;
        RECT 38.260 46.340 38.420 46.450 ;
        RECT 38.260 46.040 38.430 46.340 ;
        RECT 38.690 46.040 39.150 46.090 ;
        RECT 38.260 45.870 39.150 46.040 ;
        RECT 38.690 45.770 39.150 45.870 ;
        RECT 33.060 3.260 33.450 3.310 ;
        RECT 33.060 2.980 49.420 3.260 ;
        RECT 33.320 2.930 49.420 2.980 ;
        RECT 47.350 0.110 49.380 2.930 ;
    END
  END DIG09
  PIN DIG08
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 32.440 41.150 32.810 41.270 ;
        RECT 38.690 41.150 39.150 41.210 ;
        RECT 32.440 40.980 39.150 41.150 ;
        RECT 32.440 40.870 32.810 40.980 ;
        RECT 38.690 40.890 39.150 40.980 ;
        RECT 32.480 2.290 45.220 2.620 ;
        RECT 43.170 0.990 45.200 2.290 ;
        RECT 43.170 0.700 45.210 0.990 ;
        RECT 43.180 0.090 45.210 0.700 ;
    END
  END DIG08
  PIN DIG07
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 31.800 39.560 32.190 39.650 ;
        RECT 31.800 39.460 38.760 39.560 ;
        RECT 31.800 39.390 39.150 39.460 ;
        RECT 31.800 39.300 32.190 39.390 ;
        RECT 38.470 39.270 39.150 39.390 ;
        RECT 38.690 39.140 39.150 39.270 ;
        RECT 39.090 1.990 41.110 2.010 ;
        RECT 31.930 1.980 41.140 1.990 ;
        RECT 31.830 1.660 41.140 1.980 ;
        RECT 31.830 1.650 32.220 1.660 ;
        RECT 39.060 0.110 41.140 1.660 ;
    END
  END DIG07
  PIN DIG06
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 31.180 38.010 31.570 38.090 ;
        RECT 31.180 37.840 38.360 38.010 ;
        RECT 31.180 37.760 31.570 37.840 ;
        RECT 38.210 37.770 38.360 37.840 ;
        RECT 38.210 37.660 38.380 37.770 ;
        RECT 38.690 37.660 39.150 37.710 ;
        RECT 38.210 37.490 39.150 37.660 ;
        RECT 38.690 37.390 39.150 37.490 ;
        RECT 31.190 1.000 37.170 1.340 ;
        RECT 35.140 0.740 37.180 1.000 ;
        RECT 35.130 0.080 37.180 0.740 ;
    END
  END DIG06
  PIN DIG05
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 30.570 36.530 30.990 36.620 ;
        RECT 30.570 36.360 38.380 36.530 ;
        RECT 30.570 36.260 30.990 36.360 ;
        RECT 38.210 35.870 38.380 36.360 ;
        RECT 38.690 35.870 39.150 35.960 ;
        RECT 38.210 35.700 39.150 35.870 ;
        RECT 38.690 35.640 39.150 35.700 ;
        RECT 30.580 0.750 31.130 0.770 ;
        RECT 30.580 0.320 33.130 0.750 ;
        RECT 31.100 0.090 33.130 0.320 ;
    END
  END DIG05
  PIN DIG04
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 38.650 32.070 39.110 32.150 ;
        RECT 38.400 31.830 39.110 32.070 ;
        RECT 38.400 31.800 38.780 31.830 ;
        RECT 38.400 31.580 38.680 31.800 ;
        RECT 29.930 31.360 30.340 31.460 ;
        RECT 38.400 31.360 38.670 31.580 ;
        RECT 29.930 31.190 38.670 31.360 ;
        RECT 29.930 31.100 30.340 31.190 ;
        RECT 38.400 31.180 38.570 31.190 ;
        RECT 29.080 0.770 29.730 0.780 ;
        RECT 27.050 0.140 29.730 0.770 ;
        RECT 27.050 0.110 29.080 0.140 ;
    END
  END DIG04
  PIN DIG03
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 38.650 30.310 39.110 30.400 ;
        RECT 38.340 30.140 39.110 30.310 ;
        RECT 29.270 29.790 29.660 29.900 ;
        RECT 38.340 29.850 38.510 30.140 ;
        RECT 38.650 30.080 39.110 30.140 ;
        RECT 38.340 29.790 38.500 29.850 ;
        RECT 29.270 29.630 38.500 29.790 ;
        RECT 29.270 29.620 38.150 29.630 ;
        RECT 29.270 29.520 29.660 29.620 ;
        RECT 29.250 1.400 29.740 1.600 ;
        RECT 23.640 1.380 29.740 1.400 ;
        RECT 23.070 1.100 29.740 1.380 ;
        RECT 23.070 1.000 29.650 1.100 ;
        RECT 23.070 0.770 25.050 1.000 ;
        RECT 23.050 0.110 25.080 0.770 ;
    END
  END DIG03
  PIN DIG02
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 38.650 28.500 39.110 28.650 ;
        RECT 38.260 28.330 39.110 28.500 ;
        RECT 38.260 28.290 38.430 28.330 ;
        RECT 28.660 28.250 29.030 28.260 ;
        RECT 38.260 28.250 38.420 28.290 ;
        RECT 28.660 28.080 38.420 28.250 ;
        RECT 28.660 27.870 29.030 28.080 ;
        RECT 28.570 2.210 29.110 2.280 ;
        RECT 19.140 1.780 29.110 2.210 ;
        RECT 19.140 0.770 21.120 1.780 ;
        RECT 19.090 0.110 21.120 0.770 ;
    END
  END DIG02
  PIN DIG01
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 27.970 26.710 28.360 26.810 ;
        RECT 38.650 26.780 39.110 26.900 ;
        RECT 38.170 26.710 39.110 26.780 ;
        RECT 27.970 26.610 39.110 26.710 ;
        RECT 27.970 26.540 38.460 26.610 ;
        RECT 38.650 26.580 39.110 26.610 ;
        RECT 27.970 26.440 28.360 26.540 ;
        RECT 38.290 26.520 38.460 26.540 ;
        RECT 27.920 3.050 28.460 3.090 ;
        RECT 15.090 3.010 28.460 3.050 ;
        RECT 15.040 2.620 28.460 3.010 ;
        RECT 15.040 0.740 17.050 2.620 ;
        RECT 27.920 2.590 28.460 2.620 ;
        RECT 15.020 0.080 17.050 0.740 ;
    END
  END DIG01
  PIN CAP2    
    ANTENNAGATEAREA 9.168500 ;
    ANTENNADIFFAREA 1.850000 ;
    PORT
      LAYER met2 ;
        RECT 25.160 59.220 25.480 59.230 ;
        RECT 89.590 59.220 90.120 59.250 ;
        RECT 25.160 58.990 90.120 59.220 ;
        RECT 25.160 58.930 25.480 58.990 ;
        RECT 89.590 58.640 90.120 58.990 ;
        RECT 89.440 22.750 90.040 22.800 ;
        RECT 115.850 22.750 117.950 23.690 ;
        RECT 89.440 22.280 117.950 22.750 ;
        RECT 89.440 22.240 90.040 22.280 ;
        RECT 115.850 21.610 117.950 22.280 ;
        RECT 115.870 21.600 116.640 21.610 ;
        RECT 65.190 18.550 65.790 19.040 ;
        RECT 65.180 18.220 65.790 18.550 ;
        RECT 65.070 14.400 65.590 14.420 ;
        RECT 71.570 14.400 72.170 14.830 ;
        RECT 89.560 14.400 90.120 14.410 ;
        RECT 65.070 13.940 90.210 14.400 ;
        RECT 65.070 13.890 65.600 13.940 ;
        RECT 65.070 13.840 65.590 13.890 ;
    END
  END CAP2    
  PIN GENERALGATE01   
    ANTENNAGATEAREA 35.608200 ;
    ANTENNADIFFAREA 263.195404 ;
    PORT
      LAYER met2 ;
        RECT 0.770 70.390 1.450 71.610 ;
        RECT 2.000 70.390 2.450 70.490 ;
        RECT 0.770 70.160 2.450 70.390 ;
        RECT 0.770 69.290 1.450 70.160 ;
        RECT 2.000 70.060 2.450 70.160 ;
        RECT 2.100 66.590 2.530 67.060 ;
        RECT 2.100 66.580 4.040 66.590 ;
        RECT 2.190 66.360 4.040 66.580 ;
        RECT 46.660 65.550 47.160 65.580 ;
        RECT 52.380 65.550 52.880 65.580 ;
        RECT 46.660 65.140 76.820 65.550 ;
        RECT 46.810 65.110 76.820 65.140 ;
        RECT 42.240 64.540 42.740 64.560 ;
        RECT 47.980 64.540 48.420 64.590 ;
        RECT 62.350 64.540 62.850 64.560 ;
        RECT 42.240 64.120 68.750 64.540 ;
        RECT 42.390 64.100 68.750 64.120 ;
        RECT 47.980 64.090 48.420 64.100 ;
        RECT 68.150 64.080 68.650 64.100 ;
        RECT 86.230 61.650 86.650 61.670 ;
        RECT 115.460 61.650 116.320 62.950 ;
        RECT 39.490 61.330 39.790 61.390 ;
        RECT 80.810 61.330 81.110 61.360 ;
        RECT 39.490 61.100 81.180 61.330 ;
        RECT 86.230 61.280 116.320 61.650 ;
        RECT 86.230 61.260 86.650 61.280 ;
        RECT 39.490 61.070 39.790 61.100 ;
        RECT 80.810 61.020 81.110 61.100 ;
        RECT 115.460 60.850 116.320 61.280 ;
        RECT 32.410 60.670 32.720 60.690 ;
        RECT 22.620 60.590 22.940 60.600 ;
        RECT 32.410 60.590 32.730 60.670 ;
        RECT 56.590 60.600 56.910 60.620 ;
        RECT 56.590 60.590 56.920 60.600 ;
        RECT 63.360 60.590 63.680 60.620 ;
        RECT 78.130 60.590 78.450 60.610 ;
        RECT 92.790 60.590 93.350 60.730 ;
        RECT 22.620 60.360 93.350 60.590 ;
        RECT 22.620 60.280 22.940 60.360 ;
        RECT 32.410 60.350 32.720 60.360 ;
        RECT 56.590 60.340 56.920 60.360 ;
        RECT 63.360 60.340 63.680 60.360 ;
        RECT 78.130 60.350 78.450 60.360 ;
        RECT 92.790 60.220 93.350 60.360 ;
        RECT 28.410 60.140 28.780 60.200 ;
        RECT 91.610 60.140 92.150 60.160 ;
        RECT 28.410 59.910 92.150 60.140 ;
        RECT 28.410 59.850 28.780 59.910 ;
        RECT 60.210 59.690 60.490 59.700 ;
        RECT 31.240 59.680 31.550 59.690 ;
        RECT 60.190 59.680 60.510 59.690 ;
        RECT 62.920 59.680 63.240 59.710 ;
        RECT 77.240 59.680 77.560 59.740 ;
        RECT 90.530 59.680 91.070 59.690 ;
        RECT 31.240 59.450 91.070 59.680 ;
        RECT 91.610 59.600 92.150 59.910 ;
        RECT 31.240 59.420 31.570 59.450 ;
        RECT 60.190 59.430 60.510 59.450 ;
        RECT 62.920 59.430 63.240 59.450 ;
        RECT 60.210 59.420 60.490 59.430 ;
        RECT 31.240 59.400 31.550 59.420 ;
        RECT 90.530 59.130 91.070 59.450 ;
        RECT 0.280 58.990 0.790 59.010 ;
        RECT 19.920 58.990 20.320 59.000 ;
        RECT 0.280 58.640 20.320 58.990 ;
        RECT 0.280 58.600 0.790 58.640 ;
        RECT 19.920 58.610 20.320 58.640 ;
        RECT 20.300 55.980 20.590 56.000 ;
        RECT 7.850 55.580 20.610 55.980 ;
        RECT 0.290 52.890 1.560 53.760 ;
        RECT 7.850 52.890 8.250 55.580 ;
        RECT 20.300 55.570 20.590 55.580 ;
        RECT 77.180 55.270 77.760 55.710 ;
        RECT 77.180 55.080 77.820 55.270 ;
        RECT 18.790 54.780 19.100 54.870 ;
        RECT 18.790 54.680 19.250 54.780 ;
        RECT 20.310 54.680 20.630 54.730 ;
        RECT 18.790 54.540 20.690 54.680 ;
        RECT 19.090 54.510 20.690 54.540 ;
        RECT 20.310 54.470 20.630 54.510 ;
        RECT 77.580 54.470 77.820 55.080 ;
        RECT 78.200 55.070 78.780 55.700 ;
        RECT 81.020 55.560 81.490 55.620 ;
        RECT 105.920 55.570 106.210 55.580 ;
        RECT 105.920 55.560 106.220 55.570 ;
        RECT 116.450 55.560 116.900 55.580 ;
        RECT 81.020 55.130 116.910 55.560 ;
        RECT 82.730 55.030 92.470 55.130 ;
        RECT 105.920 55.120 106.220 55.130 ;
        RECT 105.920 55.100 106.210 55.120 ;
        RECT 82.730 54.910 83.040 55.030 ;
        RECT 16.540 54.260 16.860 54.310 ;
        RECT 17.270 54.260 17.580 54.360 ;
        RECT 16.540 54.090 17.580 54.260 ;
        RECT 82.010 54.340 82.330 54.370 ;
        RECT 16.540 54.050 16.860 54.090 ;
        RECT 17.270 54.030 17.580 54.090 ;
        RECT 53.930 54.070 54.220 54.250 ;
        RECT 82.010 54.110 92.470 54.340 ;
        RECT 18.800 53.790 19.110 53.880 ;
        RECT 18.800 53.760 19.260 53.790 ;
        RECT 20.310 53.760 20.630 53.810 ;
        RECT 18.800 53.590 20.690 53.760 ;
        RECT 18.800 53.550 19.110 53.590 ;
        RECT 20.310 53.550 20.630 53.590 ;
        RECT 16.510 53.340 16.830 53.390 ;
        RECT 17.250 53.340 17.560 53.440 ;
        RECT 16.510 53.170 17.560 53.340 ;
        RECT 16.510 53.130 16.830 53.170 ;
        RECT 17.250 53.110 17.560 53.170 ;
        RECT 0.290 52.490 8.250 52.890 ;
        RECT 18.800 52.840 19.110 52.890 ;
        RECT 20.280 52.840 20.600 52.890 ;
        RECT 18.800 52.670 20.690 52.840 ;
        RECT 18.800 52.630 19.260 52.670 ;
        RECT 20.280 52.630 20.600 52.670 ;
        RECT 18.800 52.560 19.110 52.630 ;
        RECT 0.290 51.880 1.560 52.490 ;
        RECT 16.520 52.420 16.840 52.470 ;
        RECT 17.230 52.420 17.540 52.450 ;
        RECT 16.520 52.250 17.540 52.420 ;
        RECT 16.520 52.210 16.840 52.250 ;
        RECT 17.230 52.120 17.540 52.250 ;
        RECT 20.030 52.070 20.340 52.400 ;
        RECT 52.230 52.080 52.540 52.090 ;
        RECT 53.930 52.080 54.110 54.070 ;
        RECT 82.720 53.360 83.030 53.550 ;
        RECT 85.100 53.360 85.420 53.370 ;
        RECT 82.720 53.250 92.470 53.360 ;
        RECT 107.370 53.250 107.690 53.370 ;
        RECT 82.720 53.220 107.690 53.250 ;
        RECT 82.750 53.170 107.690 53.220 ;
        RECT 85.100 53.070 107.690 53.170 ;
        RECT 50.060 51.900 61.590 52.080 ;
        RECT 81.880 52.030 87.110 52.260 ;
        RECT 52.230 51.760 52.540 51.900 ;
        RECT 15.870 51.410 16.190 51.450 ;
        RECT 15.870 51.220 17.300 51.410 ;
        RECT 15.870 51.190 16.190 51.220 ;
        RECT 20.030 51.080 20.340 51.410 ;
        RECT 48.850 51.230 49.170 51.280 ;
        RECT 51.260 51.230 51.580 51.250 ;
        RECT 53.930 51.230 54.110 51.900 ;
        RECT 83.120 51.890 83.430 52.030 ;
        RECT 80.950 51.880 83.430 51.890 ;
        RECT 80.950 51.730 92.470 51.880 ;
        RECT 80.950 51.710 83.430 51.730 ;
        RECT 83.120 51.700 83.430 51.710 ;
        RECT 48.850 51.060 54.110 51.230 ;
        RECT 48.850 51.050 52.390 51.060 ;
        RECT 48.850 51.040 61.590 51.050 ;
        RECT 48.850 50.960 49.170 51.040 ;
        RECT 50.060 50.840 61.590 51.040 ;
        RECT 51.370 50.830 61.590 50.840 ;
        RECT 52.080 50.800 52.390 50.830 ;
        RECT 15.830 50.450 16.150 50.490 ;
        RECT 15.830 50.260 17.300 50.450 ;
        RECT 18.730 50.410 19.040 50.520 ;
        RECT 44.660 50.460 44.980 50.480 ;
        RECT 15.830 50.230 16.150 50.260 ;
        RECT 18.390 50.220 19.040 50.410 ;
        RECT 18.730 50.190 19.040 50.220 ;
        RECT 20.030 50.090 20.340 50.420 ;
        RECT 44.650 50.410 44.980 50.460 ;
        RECT 47.500 50.450 48.090 50.750 ;
        RECT 106.480 50.530 106.800 50.790 ;
        RECT 106.520 50.510 107.700 50.530 ;
        RECT 47.500 50.430 47.850 50.450 ;
        RECT 45.690 50.410 46.010 50.420 ;
        RECT 47.500 50.410 47.700 50.430 ;
        RECT 44.650 50.210 47.700 50.410 ;
        RECT 106.520 50.250 107.740 50.510 ;
        RECT 44.650 50.200 44.980 50.210 ;
        RECT 44.660 50.190 44.980 50.200 ;
        RECT 45.690 50.160 46.010 50.210 ;
        RECT 106.520 50.190 107.700 50.250 ;
        RECT 106.480 50.180 107.700 50.190 ;
        RECT 51.130 49.860 61.590 50.080 ;
        RECT 106.480 49.930 106.800 50.180 ;
        RECT 51.130 49.720 51.450 49.860 ;
        RECT 15.870 49.490 16.190 49.530 ;
        RECT 15.870 49.300 17.300 49.490 ;
        RECT 47.750 49.410 48.090 49.480 ;
        RECT 15.870 49.270 16.190 49.300 ;
        RECT 47.450 49.180 48.090 49.410 ;
        RECT 51.150 49.380 51.410 49.720 ;
        RECT 44.660 48.710 44.980 48.730 ;
        RECT 44.650 48.660 44.980 48.710 ;
        RECT 45.690 48.660 46.010 48.670 ;
        RECT 47.450 48.660 47.650 49.180 ;
        RECT 51.130 49.120 51.450 49.380 ;
        RECT 53.490 49.180 54.220 49.360 ;
        RECT 53.490 48.970 53.670 49.180 ;
        RECT 60.190 49.020 60.500 49.030 ;
        RECT 44.650 48.460 47.650 48.660 ;
        RECT 48.850 48.890 49.170 48.970 ;
        RECT 51.330 48.940 53.670 48.970 ;
        RECT 60.180 48.960 60.510 49.020 ;
        RECT 51.260 48.890 53.670 48.940 ;
        RECT 59.830 48.910 60.510 48.960 ;
        RECT 48.850 48.810 53.670 48.890 ;
        RECT 48.850 48.700 51.580 48.810 ;
        RECT 52.060 48.800 53.670 48.810 ;
        RECT 52.760 48.790 53.670 48.800 ;
        RECT 48.850 48.650 49.170 48.700 ;
        RECT 51.260 48.680 51.580 48.700 ;
        RECT 56.600 48.740 60.510 48.910 ;
        RECT 82.660 48.750 87.110 48.910 ;
        RECT 56.600 48.690 60.500 48.740 ;
        RECT 82.630 48.710 87.110 48.750 ;
        RECT 80.910 48.630 81.220 48.710 ;
        RECT 82.630 48.630 82.860 48.710 ;
        RECT 83.160 48.630 83.470 48.710 ;
        RECT 44.650 48.450 44.980 48.460 ;
        RECT 44.660 48.440 44.980 48.450 ;
        RECT 45.690 48.410 46.010 48.460 ;
        RECT 80.910 48.400 83.470 48.630 ;
        RECT 80.910 48.380 81.220 48.400 ;
        RECT 52.080 48.300 52.390 48.370 ;
        RECT 50.060 48.090 61.590 48.300 ;
        RECT 51.370 48.080 61.590 48.090 ;
        RECT 48.850 48.030 49.170 48.080 ;
        RECT 51.260 48.030 51.580 48.050 ;
        RECT 52.080 48.040 52.390 48.080 ;
        RECT 48.850 48.010 51.580 48.030 ;
        RECT 53.590 48.030 54.140 48.080 ;
        RECT 53.590 48.010 53.770 48.030 ;
        RECT 48.850 47.850 53.770 48.010 ;
        RECT 48.850 47.840 51.580 47.850 ;
        RECT 48.850 47.760 49.170 47.840 ;
        RECT 51.260 47.790 51.580 47.840 ;
        RECT 47.610 47.540 48.090 47.550 ;
        RECT 47.480 47.250 48.090 47.540 ;
        RECT 47.480 47.100 47.800 47.250 ;
        RECT 52.230 47.210 52.540 47.350 ;
        RECT 50.060 47.200 52.540 47.210 ;
        RECT 44.660 46.960 44.980 46.980 ;
        RECT 44.650 46.910 44.980 46.960 ;
        RECT 45.690 46.910 46.010 46.920 ;
        RECT 47.480 46.910 47.680 47.100 ;
        RECT 50.060 47.050 61.590 47.200 ;
        RECT 50.060 47.030 52.540 47.050 ;
        RECT 52.230 47.020 52.540 47.030 ;
        RECT 44.650 46.710 47.680 46.910 ;
        RECT 44.650 46.700 44.980 46.710 ;
        RECT 44.660 46.690 44.980 46.700 ;
        RECT 45.690 46.660 46.010 46.710 ;
        RECT 80.910 46.490 81.220 46.550 ;
        RECT 82.630 46.490 82.860 48.400 ;
        RECT 83.210 46.490 83.520 46.510 ;
        RECT 80.910 46.300 83.830 46.490 ;
        RECT 80.910 46.260 87.110 46.300 ;
        RECT 80.910 46.220 81.220 46.260 ;
        RECT 82.630 46.230 82.860 46.260 ;
        RECT 81.880 46.000 82.860 46.230 ;
        RECT 83.210 46.180 87.110 46.260 ;
        RECT 83.470 46.100 87.110 46.180 ;
        RECT 83.470 45.790 83.670 46.100 ;
        RECT 80.910 45.660 81.220 45.710 ;
        RECT 83.200 45.660 83.670 45.790 ;
        RECT 80.910 45.440 83.830 45.660 ;
        RECT 80.910 45.380 81.220 45.440 ;
        RECT 83.470 45.400 83.670 45.440 ;
        RECT 81.890 45.250 83.670 45.400 ;
        RECT 81.890 45.180 83.640 45.250 ;
        RECT 80.910 43.500 81.220 43.550 ;
        RECT 83.120 43.500 83.430 43.540 ;
        RECT 80.910 43.270 83.620 43.500 ;
        RECT 80.910 43.220 81.220 43.270 ;
        RECT 83.120 43.210 83.430 43.270 ;
        RECT 86.170 39.430 86.610 39.550 ;
        RECT 86.040 39.250 86.610 39.430 ;
        RECT 57.590 39.090 57.900 39.220 ;
        RECT 73.080 39.090 73.390 39.220 ;
        RECT 86.160 39.150 86.610 39.250 ;
        RECT 86.160 39.090 86.560 39.150 ;
        RECT 55.430 38.910 86.560 39.090 ;
        RECT 57.590 38.890 57.900 38.910 ;
        RECT 73.080 38.890 73.390 38.910 ;
        RECT 92.700 38.430 93.300 38.490 ;
        RECT 115.420 38.430 116.320 39.460 ;
        RECT 92.700 37.960 116.320 38.430 ;
        RECT 92.700 37.910 93.300 37.960 ;
        RECT 115.420 37.370 116.320 37.960 ;
        RECT 15.830 34.460 16.140 34.480 ;
        RECT 16.490 34.460 16.800 34.480 ;
        RECT 15.830 33.990 23.150 34.460 ;
        RECT 15.830 33.970 16.140 33.990 ;
        RECT 16.490 33.970 16.800 33.990 ;
        RECT 22.680 33.310 23.150 33.990 ;
        RECT 54.980 33.350 55.290 33.360 ;
        RECT 52.820 33.310 55.290 33.350 ;
        RECT 115.450 33.310 116.350 34.280 ;
        RECT 14.500 33.180 14.760 33.250 ;
        RECT 16.550 33.180 16.870 33.200 ;
        RECT 18.310 33.180 18.640 33.220 ;
        RECT 14.500 32.990 18.640 33.180 ;
        RECT 14.500 32.930 14.760 32.990 ;
        RECT 16.550 32.940 16.870 32.990 ;
        RECT 18.310 32.950 18.640 32.990 ;
        RECT 22.680 32.840 116.350 33.310 ;
        RECT 13.950 32.780 14.270 32.820 ;
        RECT 15.890 32.780 16.210 32.840 ;
        RECT 18.810 32.780 19.130 32.820 ;
        RECT 13.950 32.590 19.130 32.780 ;
        RECT 91.610 32.720 92.180 32.840 ;
        RECT 13.950 32.560 14.270 32.590 ;
        RECT 15.890 32.580 16.210 32.590 ;
        RECT 18.810 32.560 19.130 32.590 ;
        RECT 20.290 32.220 20.590 32.240 ;
        RECT 20.280 32.200 20.600 32.220 ;
        RECT 18.060 31.980 20.600 32.200 ;
        RECT 115.450 32.190 116.350 32.840 ;
        RECT 18.060 31.540 18.280 31.980 ;
        RECT 20.280 31.960 20.600 31.980 ;
        RECT 20.290 31.940 20.590 31.960 ;
        RECT 19.670 31.070 19.960 31.090 ;
        RECT 19.660 31.030 19.980 31.070 ;
        RECT 18.090 30.840 19.980 31.030 ;
        RECT 19.660 30.810 19.980 30.840 ;
        RECT 19.670 30.800 19.960 30.810 ;
        RECT 20.440 30.800 20.750 30.840 ;
        RECT 18.550 30.580 20.750 30.800 ;
        RECT 20.440 30.510 20.750 30.580 ;
        RECT 19.220 30.350 19.530 30.400 ;
        RECT 18.550 30.140 19.530 30.350 ;
        RECT 19.220 30.070 19.530 30.140 ;
        RECT 18.770 29.000 19.090 29.020 ;
        RECT 13.980 28.910 14.270 28.920 ;
        RECT 13.970 28.890 14.290 28.910 ;
        RECT 13.970 28.670 14.970 28.890 ;
        RECT 18.550 28.780 19.090 29.000 ;
        RECT 18.770 28.760 19.090 28.780 ;
        RECT 13.970 28.650 14.290 28.670 ;
        RECT 13.980 28.630 14.270 28.650 ;
        RECT 19.240 28.430 19.560 28.480 ;
        RECT 18.070 28.420 19.560 28.430 ;
        RECT 21.520 28.420 21.840 28.540 ;
        RECT 18.070 28.220 21.840 28.420 ;
        RECT 18.550 28.210 21.530 28.220 ;
        RECT 19.240 28.180 19.560 28.210 ;
        RECT 90.490 28.070 91.040 28.080 ;
        RECT 90.490 28.050 91.050 28.070 ;
        RECT 115.420 28.050 116.320 29.200 ;
        RECT 90.490 27.580 116.320 28.050 ;
        RECT 90.490 27.570 91.050 27.580 ;
        RECT 90.490 27.550 91.040 27.570 ;
        RECT 18.770 27.460 19.090 27.470 ;
        RECT 18.550 27.240 19.090 27.460 ;
        RECT 18.770 27.210 19.090 27.240 ;
        RECT 115.420 27.110 116.320 27.580 ;
        RECT 18.550 26.460 18.820 26.470 ;
        RECT 19.250 26.460 19.560 26.520 ;
        RECT 18.550 26.250 19.560 26.460 ;
        RECT 19.250 26.190 19.560 26.250 ;
        RECT 15.080 25.850 15.390 25.860 ;
        RECT 16.170 25.850 16.480 25.860 ;
        RECT 13.760 25.840 16.480 25.850 ;
        RECT 13.530 25.530 16.480 25.840 ;
        RECT 20.420 25.690 20.730 25.740 ;
        RECT 13.530 25.520 16.470 25.530 ;
        RECT 13.530 23.900 13.880 25.520 ;
        RECT 18.550 25.470 20.730 25.690 ;
        RECT 20.420 25.410 20.730 25.470 ;
        RECT 95.680 25.240 96.240 25.310 ;
        RECT 108.400 25.240 109.080 25.300 ;
        RECT 115.930 25.240 116.590 25.880 ;
        RECT 14.530 25.170 14.840 25.180 ;
        RECT 15.630 25.170 15.940 25.180 ;
        RECT 16.730 25.170 17.040 25.180 ;
        RECT 14.500 24.850 17.660 25.170 ;
        RECT 46.740 24.980 47.070 25.000 ;
        RECT 17.340 23.900 17.660 24.850 ;
        RECT 46.730 24.900 47.080 24.980 ;
        RECT 52.480 24.900 52.800 24.960 ;
        RECT 46.730 24.740 52.800 24.900 ;
        RECT 95.680 24.830 116.590 25.240 ;
        RECT 95.680 24.780 96.240 24.830 ;
        RECT 108.400 24.770 109.080 24.830 ;
        RECT 46.730 24.670 47.080 24.740 ;
        RECT 52.480 24.690 52.800 24.740 ;
        RECT 115.930 24.730 116.590 24.830 ;
        RECT 42.310 24.280 42.640 24.520 ;
        RECT 48.170 24.410 48.470 24.420 ;
        RECT 48.160 24.280 48.480 24.410 ;
        RECT 58.700 24.280 58.980 24.580 ;
        RECT 62.730 24.280 63.030 24.560 ;
        RECT 42.310 24.260 63.030 24.280 ;
        RECT 42.310 24.230 63.020 24.260 ;
        RECT 42.310 24.120 62.960 24.230 ;
        RECT 46.120 23.900 46.560 23.910 ;
        RECT 0.800 23.890 46.560 23.900 ;
        RECT 0.800 23.480 46.580 23.890 ;
        RECT 13.530 23.080 13.880 23.480 ;
        RECT 13.530 22.930 16.480 23.080 ;
        RECT 17.340 22.930 17.660 23.480 ;
        RECT 39.270 23.470 39.750 23.480 ;
        RECT 46.100 23.470 46.580 23.480 ;
        RECT 46.120 23.460 46.560 23.470 ;
        RECT 57.930 23.100 58.240 23.130 ;
        RECT 59.020 23.100 59.330 23.110 ;
        RECT 62.970 23.100 63.280 23.110 ;
        RECT 64.060 23.100 64.370 23.130 ;
        RECT 48.120 23.070 48.430 23.100 ;
        RECT 49.210 23.070 49.520 23.080 ;
        RECT 53.160 23.070 53.470 23.080 ;
        RECT 54.250 23.070 54.560 23.100 ;
        RECT 0.780 22.510 42.760 22.930 ;
        RECT 48.120 22.770 51.070 23.070 ;
        RECT 49.210 22.750 49.520 22.770 ;
        RECT 50.320 22.730 51.070 22.770 ;
        RECT 50.690 22.600 51.070 22.730 ;
        RECT 13.530 21.880 13.880 22.510 ;
        RECT 13.530 21.750 13.910 21.880 ;
        RECT 13.530 21.710 14.280 21.750 ;
        RECT 15.080 21.710 15.390 21.730 ;
        RECT 13.530 21.410 16.480 21.710 ;
        RECT 15.080 21.400 15.390 21.410 ;
        RECT 16.170 21.380 16.480 21.410 ;
        RECT 14.530 21.030 14.840 21.040 ;
        RECT 17.340 21.030 17.660 22.510 ;
        RECT 23.830 22.010 24.660 22.510 ;
        RECT 50.720 21.730 51.070 22.600 ;
        RECT 48.120 21.400 51.070 21.730 ;
        RECT 14.510 20.700 17.660 21.030 ;
        RECT 14.510 20.690 17.570 20.700 ;
        RECT 17.420 20.490 17.710 20.510 ;
        RECT 19.650 20.490 19.960 20.510 ;
        RECT 17.410 20.130 19.960 20.490 ;
        RECT 17.420 20.110 17.710 20.130 ;
        RECT 19.650 20.110 19.960 20.130 ;
        RECT 46.700 18.520 47.300 19.010 ;
        RECT 50.720 18.960 51.070 21.400 ;
        RECT 48.130 18.950 51.070 18.960 ;
        RECT 48.120 18.640 51.070 18.950 ;
        RECT 51.610 22.770 54.560 23.070 ;
        RECT 57.930 22.800 60.880 23.100 ;
        RECT 59.020 22.780 59.330 22.800 ;
        RECT 51.610 22.730 52.360 22.770 ;
        RECT 53.160 22.750 53.470 22.770 ;
        RECT 60.130 22.760 60.880 22.800 ;
        RECT 51.610 22.600 51.990 22.730 ;
        RECT 60.500 22.630 60.880 22.760 ;
        RECT 51.610 21.730 51.960 22.600 ;
        RECT 60.530 21.760 60.880 22.630 ;
        RECT 51.610 21.400 54.560 21.730 ;
        RECT 57.930 21.430 60.880 21.760 ;
        RECT 51.610 18.960 51.960 21.400 ;
        RECT 51.610 18.950 54.550 18.960 ;
        RECT 51.610 18.640 54.560 18.950 ;
        RECT 48.120 18.630 50.840 18.640 ;
        RECT 51.840 18.630 54.560 18.640 ;
        RECT 48.120 18.620 48.430 18.630 ;
        RECT 49.210 18.620 49.520 18.630 ;
        RECT 53.160 18.620 53.470 18.630 ;
        RECT 54.250 18.620 54.560 18.630 ;
        RECT 55.380 18.520 55.980 19.010 ;
        RECT 46.700 18.190 47.310 18.520 ;
        RECT 55.370 18.190 55.980 18.520 ;
        RECT 56.510 18.550 57.110 19.040 ;
        RECT 60.530 18.990 60.880 21.430 ;
        RECT 57.940 18.980 60.880 18.990 ;
        RECT 57.930 18.670 60.880 18.980 ;
        RECT 61.420 22.800 64.370 23.100 ;
        RECT 61.420 22.760 62.170 22.800 ;
        RECT 62.970 22.780 63.280 22.800 ;
        RECT 61.420 22.630 61.800 22.760 ;
        RECT 61.420 21.760 61.770 22.630 ;
        RECT 61.420 21.430 64.370 21.760 ;
        RECT 61.420 18.990 61.770 21.430 ;
        RECT 68.780 19.600 71.840 19.610 ;
        RECT 68.780 19.270 71.930 19.600 ;
        RECT 68.800 19.260 69.110 19.270 ;
        RECT 61.420 18.980 64.360 18.990 ;
        RECT 61.420 18.670 64.370 18.980 ;
        RECT 69.350 18.890 69.660 18.900 ;
        RECT 70.440 18.890 70.750 18.920 ;
        RECT 57.930 18.660 60.650 18.670 ;
        RECT 61.650 18.660 64.370 18.670 ;
        RECT 57.930 18.650 58.240 18.660 ;
        RECT 59.020 18.650 59.330 18.660 ;
        RECT 62.970 18.650 63.280 18.660 ;
        RECT 64.060 18.650 64.370 18.660 ;
        RECT 67.800 18.590 70.750 18.890 ;
        RECT 67.800 18.550 68.550 18.590 ;
        RECT 69.350 18.570 69.660 18.590 ;
        RECT 56.510 18.220 57.120 18.550 ;
        RECT 67.800 18.420 68.180 18.550 ;
        RECT 50.810 17.950 61.710 17.980 ;
        RECT 50.800 17.700 61.710 17.950 ;
        RECT 50.800 17.670 51.140 17.700 ;
        RECT 51.540 17.690 51.880 17.700 ;
        RECT 60.610 17.670 60.950 17.700 ;
        RECT 67.800 17.550 68.150 18.420 ;
        RECT 67.800 17.220 70.750 17.550 ;
        RECT 46.880 17.160 47.380 17.170 ;
        RECT 67.800 17.160 68.150 17.220 ;
        RECT 71.610 17.160 71.930 19.270 ;
        RECT 92.810 17.160 93.370 17.180 ;
        RECT 20.280 16.830 20.560 16.840 ;
        RECT 16.690 16.500 20.580 16.830 ;
        RECT 46.880 16.700 93.370 17.160 ;
        RECT 46.880 16.640 47.400 16.700 ;
        RECT 46.880 16.620 47.380 16.640 ;
        RECT 20.280 16.480 20.560 16.500 ;
        RECT 67.800 16.250 68.150 16.700 ;
        RECT 68.770 16.490 71.930 16.700 ;
        RECT 92.810 16.680 93.370 16.700 ;
        RECT 71.610 16.250 71.930 16.490 ;
        RECT 55.190 15.790 92.270 16.250 ;
        RECT 55.260 15.690 55.780 15.790 ;
        RECT 67.800 15.340 68.150 15.790 ;
        RECT 71.610 15.450 71.930 15.790 ;
        RECT 91.620 15.730 92.180 15.790 ;
        RECT 68.770 15.340 71.930 15.450 ;
        RECT 56.630 15.270 91.180 15.340 ;
        RECT 12.860 15.150 13.210 15.180 ;
        RECT 19.240 15.170 19.570 15.210 ;
        RECT 19.230 15.150 19.580 15.170 ;
        RECT 12.860 14.890 22.890 15.150 ;
        RECT 12.900 14.860 22.890 14.890 ;
        RECT 56.620 14.880 91.180 15.270 ;
        RECT 107.860 15.250 108.150 15.310 ;
        RECT 107.690 14.940 108.150 15.250 ;
        RECT 107.860 14.900 108.150 14.940 ;
        RECT 19.240 14.840 19.570 14.860 ;
        RECT 16.690 14.520 17.300 14.540 ;
        RECT 16.690 14.210 19.040 14.520 ;
        RECT 16.700 14.180 19.040 14.210 ;
        RECT 16.700 13.940 19.080 14.180 ;
        RECT 16.700 13.920 19.040 13.940 ;
        RECT 16.700 13.720 17.300 13.920 ;
        RECT 18.070 13.850 18.730 13.920 ;
        RECT 18.100 13.840 18.700 13.850 ;
        RECT 22.590 12.780 22.880 14.860 ;
        RECT 56.620 14.750 57.270 14.880 ;
        RECT 67.800 14.780 68.150 14.880 ;
        RECT 90.490 14.860 91.050 14.880 ;
        RECT 67.800 14.770 70.740 14.780 ;
        RECT 67.800 14.460 70.750 14.770 ;
        RECT 107.870 14.580 108.150 14.900 ;
        RECT 68.030 14.450 70.750 14.460 ;
        RECT 69.350 14.440 69.660 14.450 ;
        RECT 70.440 14.440 70.750 14.450 ;
        RECT 107.690 14.270 108.150 14.580 ;
        RECT 107.870 14.150 108.150 14.270 ;
        RECT 39.010 12.780 39.330 12.800 ;
        RECT 95.010 12.780 96.170 12.810 ;
        RECT 22.400 11.660 96.170 12.780 ;
        RECT 39.010 11.640 39.330 11.660 ;
        RECT 50.380 11.580 52.300 11.660 ;
        RECT 60.190 11.550 62.120 11.660 ;
        RECT 95.010 11.630 96.170 11.660 ;
        RECT 1.930 8.330 2.430 8.440 ;
        RECT 70.900 8.360 71.290 8.370 ;
        RECT 70.890 8.330 71.290 8.360 ;
        RECT 1.930 8.050 71.290 8.330 ;
        RECT 1.930 7.970 2.430 8.050 ;
        RECT 70.890 8.030 71.290 8.050 ;
        RECT 70.900 8.020 71.290 8.030 ;
      LAYER via2 ;
        RECT 77.300 55.240 77.620 55.560 ;
        RECT 78.330 55.230 78.650 55.550 ;
    END
  END GENERALGATE01   
  PIN OUTPUTTA1    
    ANTENNADIFFAREA 4.694300 ;
    PORT
      LAYER nwell ;
        RECT 11.670 65.390 13.280 66.180 ;
        RECT 13.780 65.390 14.290 65.560 ;
        RECT 14.330 65.390 15.480 65.560 ;
        RECT 11.670 64.210 15.670 65.390 ;
        RECT 11.670 64.200 12.460 64.210 ;
        RECT 13.780 64.200 15.670 64.210 ;
        RECT 13.780 64.000 14.290 64.200 ;
        RECT 14.330 64.010 15.480 64.200 ;
        RECT 113.440 47.790 114.720 53.470 ;
      LAYER met2 ;
        RECT 0.770 66.200 1.450 67.080 ;
        RECT 0.770 65.880 4.130 66.200 ;
        RECT 0.770 65.730 1.450 65.880 ;
        RECT 0.000 65.520 12.010 65.730 ;
        RECT 0.770 64.760 1.450 65.520 ;
        RECT 3.460 65.490 4.040 65.520 ;
        RECT 3.460 65.460 3.780 65.490 ;
        RECT 11.430 65.070 11.670 65.520 ;
        RECT 11.410 64.740 11.720 65.070 ;
        RECT 112.870 63.180 113.640 63.330 ;
        RECT 3.380 62.760 113.640 63.180 ;
        RECT 112.870 62.620 113.640 62.760 ;
        RECT 112.680 43.420 113.460 43.570 ;
        RECT 115.420 43.420 116.320 44.340 ;
        RECT 112.680 42.950 116.320 43.420 ;
        RECT 112.680 42.800 113.460 42.950 ;
        RECT 115.420 42.250 116.320 42.950 ;
    END
  END OUTPUTTA1    
  PIN DRAINOUT
    ANTENNADIFFAREA 3.068100 ;
    PORT
      LAYER met2 ;
        RECT 83.360 56.770 83.680 56.780 ;
        RECT 83.120 56.760 83.680 56.770 ;
        RECT 80.950 56.580 92.470 56.760 ;
        RECT 115.460 56.580 116.320 58.560 ;
        RECT 83.120 56.440 83.430 56.580 ;
        RECT 87.110 56.460 116.320 56.580 ;
        RECT 87.110 56.210 116.210 56.460 ;
        RECT 87.110 56.180 87.520 56.210 ;
        RECT 49.450 34.320 49.760 34.340 ;
        RECT 87.090 34.320 87.540 34.350 ;
        RECT 49.450 33.910 87.540 34.320 ;
        RECT 49.450 33.890 49.760 33.910 ;
        RECT 54.980 33.780 55.290 33.910 ;
        RECT 87.090 33.890 87.540 33.910 ;
        RECT 52.820 33.600 62.890 33.780 ;
        RECT 54.980 33.580 55.290 33.600 ;
    END
  END DRAINOUT
  PIN COLUMN2
    ANTENNAGATEAREA 1.870000 ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met2 ;
        RECT 85.450 66.360 85.890 66.380 ;
        RECT 115.490 66.360 116.350 67.040 ;
        RECT 85.450 65.990 116.350 66.360 ;
        RECT 85.450 65.970 85.890 65.990 ;
        RECT 115.490 64.940 116.350 65.990 ;
        RECT 85.430 41.800 85.860 41.880 ;
        RECT 74.170 41.540 85.860 41.800 ;
        RECT 74.170 41.530 74.490 41.540 ;
        RECT 85.430 41.470 85.860 41.540 ;
    END
  END COLUMN2
  PIN COLUMN1
    ANTENNAGATEAREA 3.120400 ;
    ANTENNADIFFAREA 11.364100 ;
    PORT
      LAYER met2 ;
        RECT 84.620 69.820 85.080 69.840 ;
        RECT 115.490 69.820 116.350 71.170 ;
        RECT 84.620 69.450 116.350 69.820 ;
        RECT 84.620 69.430 85.080 69.450 ;
        RECT 115.490 69.070 116.350 69.450 ;
        RECT 54.260 48.540 54.580 48.660 ;
        RECT 76.460 48.540 76.780 48.660 ;
        RECT 54.260 48.360 76.780 48.540 ;
        RECT 75.590 45.850 75.910 46.110 ;
        RECT 75.630 45.830 76.810 45.850 ;
        RECT 75.630 45.570 76.850 45.830 ;
        RECT 75.630 45.510 76.810 45.570 ;
        RECT 75.590 45.500 76.810 45.510 ;
        RECT 75.590 45.250 75.910 45.500 ;
        RECT 56.830 42.400 57.150 42.410 ;
        RECT 84.640 42.400 85.100 42.470 ;
        RECT 56.830 42.120 85.100 42.400 ;
        RECT 56.830 42.070 57.150 42.120 ;
        RECT 84.640 42.060 85.100 42.120 ;
        RECT 55.630 40.910 75.370 41.090 ;
        RECT 55.630 40.770 56.050 40.910 ;
        RECT 75.030 40.780 75.370 40.910 ;
        RECT 58.220 31.280 58.540 31.300 ;
        RECT 56.010 31.060 56.330 31.120 ;
        RECT 58.220 31.090 66.140 31.280 ;
        RECT 66.300 31.090 66.610 31.130 ;
        RECT 58.220 31.070 66.610 31.090 ;
        RECT 58.220 31.060 58.540 31.070 ;
        RECT 60.030 31.060 60.360 31.070 ;
        RECT 56.010 30.890 60.360 31.060 ;
        RECT 56.010 30.840 56.330 30.890 ;
        RECT 60.030 30.830 60.360 30.890 ;
        RECT 65.930 30.880 66.610 31.070 ;
        RECT 66.300 30.800 66.610 30.880 ;
        RECT 55.260 30.660 62.890 30.670 ;
        RECT 54.950 30.640 62.890 30.660 ;
        RECT 53.930 30.530 62.890 30.640 ;
        RECT 52.820 30.500 62.890 30.530 ;
        RECT 52.820 30.350 55.380 30.500 ;
        RECT 53.870 30.160 54.150 30.350 ;
        RECT 54.950 30.330 55.290 30.350 ;
        RECT 54.950 30.240 55.100 30.330 ;
        RECT 58.200 30.240 58.520 30.250 ;
        RECT 54.950 30.100 58.520 30.240 ;
        RECT 52.820 30.090 58.520 30.100 ;
        RECT 52.820 29.920 55.290 30.090 ;
        RECT 58.080 29.990 58.520 30.090 ;
        RECT 54.980 29.780 55.290 29.920 ;
        RECT 47.270 25.270 47.590 25.320 ;
        RECT 53.880 25.270 54.200 25.370 ;
        RECT 47.270 25.110 54.200 25.270 ;
        RECT 47.270 25.060 47.590 25.110 ;
        RECT 53.880 25.090 54.200 25.110 ;
        RECT 47.030 23.780 50.090 23.790 ;
        RECT 46.940 23.450 50.090 23.780 ;
        RECT 46.940 22.770 47.260 23.450 ;
        RECT 49.760 23.440 50.070 23.450 ;
        RECT 46.790 22.390 47.260 22.770 ;
        RECT 46.940 21.000 47.260 22.390 ;
        RECT 46.940 20.670 50.100 21.000 ;
        RECT 46.940 19.630 47.260 20.670 ;
        RECT 46.940 19.310 50.100 19.630 ;
        RECT 47.560 19.300 47.870 19.310 ;
        RECT 48.660 19.300 48.970 19.310 ;
        RECT 49.760 19.300 50.070 19.310 ;
    END
  END COLUMN1
  PIN GATE2
    PORT
      LAYER met2 ;
        RECT 69.480 58.060 69.760 58.080 ;
        RECT 69.460 58.030 69.780 58.060 ;
        RECT 101.600 58.030 102.940 58.570 ;
        RECT 69.460 57.820 102.940 58.030 ;
        RECT 69.460 57.800 69.780 57.820 ;
        RECT 69.480 57.780 69.760 57.800 ;
        RECT 101.600 57.290 102.940 57.820 ;
    END
  END GATE2
  PIN DRAININJECT
    PORT
      LAYER met2 ;
        RECT 45.000 67.930 45.450 67.950 ;
        RECT 44.990 67.870 45.470 67.930 ;
        RECT 22.600 67.570 45.470 67.870 ;
        RECT 44.990 67.510 45.470 67.570 ;
        RECT 45.000 67.490 45.450 67.510 ;
    END
  END DRAININJECT
  PIN VTUN
    PORT
      LAYER met2 ;
        RECT 41.150 67.170 41.600 67.190 ;
        RECT 41.140 67.160 41.620 67.170 ;
        RECT 64.760 67.160 66.180 67.200 ;
        RECT 41.140 66.760 66.230 67.160 ;
        RECT 41.140 66.750 41.620 66.760 ;
        RECT 41.150 66.730 41.600 66.750 ;
        RECT 64.760 66.720 66.180 66.760 ;
    END
  END VTUN
  PIN LARGECAPACITOR
    ANTENNADIFFAREA 3.550400 ;
    PORT
      LAYER met2 ;
        RECT 0.320 61.940 1.000 62.610 ;
        RECT 9.240 61.940 9.710 61.960 ;
        RECT 0.320 61.360 9.710 61.940 ;
        RECT 0.320 61.290 1.040 61.360 ;
        RECT 9.240 61.340 9.710 61.360 ;
        RECT 10.690 61.290 11.000 61.410 ;
        RECT 20.550 61.290 20.860 61.430 ;
        RECT 0.000 61.100 20.860 61.290 ;
        RECT 0.000 61.080 20.830 61.100 ;
        RECT 0.320 60.290 1.000 61.080 ;
    END
  END LARGECAPACITOR
  PIN DRAIN6N
    PORT
      LAYER met2 ;
        RECT 11.610 17.530 11.980 17.540 ;
        RECT 0.720 16.710 1.990 17.410 ;
        RECT 10.290 17.150 12.900 17.530 ;
        RECT 10.290 16.710 10.670 17.150 ;
        RECT 11.610 17.130 11.980 17.150 ;
        RECT 0.720 16.330 10.670 16.710 ;
        RECT 0.720 15.530 1.990 16.330 ;
    END
  END DRAIN6N
  PIN DRAIN6P
    ANTENNADIFFAREA 4.317200 ;
    PORT
      LAYER met2 ;
        RECT 14.480 14.100 14.790 14.110 ;
        RECT 15.570 14.100 15.880 14.110 ;
        RECT 13.160 14.090 15.880 14.100 ;
        RECT 12.930 13.780 15.880 14.090 ;
        RECT 12.930 13.770 15.870 13.780 ;
        RECT 0.720 11.480 1.990 12.390 ;
        RECT 0.720 11.100 10.690 11.480 ;
        RECT 0.720 10.510 1.990 11.100 ;
        RECT 10.310 10.250 10.690 11.100 ;
        RECT 12.930 11.330 13.280 13.770 ;
        RECT 12.930 11.000 15.880 11.330 ;
        RECT 11.610 10.250 11.980 10.260 ;
        RECT 12.930 10.250 13.280 11.000 ;
        RECT 10.310 10.130 13.280 10.250 ;
        RECT 10.310 10.000 13.310 10.130 ;
        RECT 10.310 9.960 13.680 10.000 ;
        RECT 14.480 9.960 14.790 9.980 ;
        RECT 10.310 9.870 15.880 9.960 ;
        RECT 11.610 9.850 11.980 9.870 ;
        RECT 12.930 9.660 15.880 9.870 ;
        RECT 14.480 9.650 14.790 9.660 ;
        RECT 15.570 9.630 15.880 9.660 ;
    END
  END DRAIN6P
  PIN DRAIN5P
    PORT
      LAYER met2 ;
        RECT 9.880 27.160 10.290 27.180 ;
        RECT 11.650 27.160 13.640 27.180 ;
        RECT 9.880 27.120 13.640 27.160 ;
        RECT 9.880 26.900 14.970 27.120 ;
        RECT 9.880 26.790 12.030 26.900 ;
        RECT 9.880 26.770 10.290 26.790 ;
        RECT 11.650 26.770 12.020 26.790 ;
        RECT 0.660 20.920 1.930 21.700 ;
        RECT 9.890 20.920 10.300 20.940 ;
        RECT 0.660 20.550 10.300 20.920 ;
        RECT 0.660 19.820 1.930 20.550 ;
        RECT 9.890 20.530 10.300 20.550 ;
    END
  END DRAIN5P
  PIN DARIN4P
    PORT
      LAYER met2 ;
        RECT 0.720 30.170 1.990 30.940 ;
        RECT 0.720 29.800 6.710 30.170 ;
        RECT 0.720 29.060 1.990 29.800 ;
        RECT 6.340 28.140 6.710 29.800 ;
        RECT 6.340 27.960 12.290 28.140 ;
        RECT 6.340 27.890 12.360 27.960 ;
        RECT 13.750 27.890 14.970 27.900 ;
        RECT 6.340 27.770 14.970 27.890 ;
        RECT 11.650 27.730 14.970 27.770 ;
        RECT 12.010 27.680 14.970 27.730 ;
    END
  END DARIN4P
  PIN DRAIN5N
    PORT
      LAYER met2 ;
        RECT 4.650 31.820 5.420 32.010 ;
        RECT 11.650 31.820 12.040 31.840 ;
        RECT 4.650 31.780 12.040 31.820 ;
        RECT 4.650 31.570 14.960 31.780 ;
        RECT 4.650 31.450 12.030 31.570 ;
        RECT 4.650 31.270 5.420 31.450 ;
        RECT 11.650 31.430 12.020 31.450 ;
        RECT 0.720 26.030 1.990 26.850 ;
        RECT 4.650 26.030 5.450 26.170 ;
        RECT 0.720 25.530 5.450 26.030 ;
        RECT 0.720 24.970 1.990 25.530 ;
        RECT 4.650 25.400 5.450 25.530 ;
    END
  END DRAIN5N
  PIN DRAIN4N
    PORT
      LAYER met2 ;
        RECT 0.660 34.200 1.930 35.040 ;
        RECT 0.660 33.830 10.360 34.200 ;
        RECT 0.660 33.160 1.930 33.830 ;
        RECT 9.990 32.480 10.360 33.830 ;
        RECT 9.990 32.470 12.020 32.480 ;
        RECT 9.990 32.290 12.240 32.470 ;
        RECT 9.990 32.230 13.640 32.290 ;
        RECT 9.990 32.110 14.970 32.230 ;
        RECT 11.650 32.070 14.970 32.110 ;
        RECT 12.020 32.010 14.970 32.070 ;
    END
  END DRAIN4N
  PIN DRAIN3P
    PORT
      LAYER met2 ;
        RECT 11.650 49.720 17.300 49.910 ;
        RECT 0.720 38.350 1.990 39.260 ;
        RECT 11.650 38.350 12.020 49.720 ;
        RECT 0.720 37.980 12.020 38.350 ;
        RECT 0.720 37.380 1.990 37.980 ;
    END
  END DRAIN3P
  PIN DRAIN2P
    PORT
      LAYER met2 ;
        RECT 10.810 51.810 17.300 51.830 ;
        RECT 10.520 51.640 17.300 51.810 ;
        RECT 10.520 51.460 12.020 51.640 ;
        RECT 10.520 50.870 11.180 51.460 ;
        RECT 11.650 51.420 12.020 51.460 ;
        RECT 10.520 50.680 17.300 50.870 ;
        RECT 10.520 50.500 12.020 50.680 ;
        RECT 10.520 50.490 11.190 50.500 ;
        RECT 10.520 50.450 11.180 50.490 ;
        RECT 11.650 50.460 12.020 50.500 ;
        RECT 0.660 43.190 1.930 44.080 ;
        RECT 10.520 43.190 10.890 50.450 ;
        RECT 0.660 42.820 10.890 43.190 ;
        RECT 0.660 42.200 1.930 42.820 ;
    END
  END DRAIN2P
  PIN DRAIN3N
    ANTENNADIFFAREA 0.390600 ;
    PORT
      LAYER met2 ;
        RECT 11.650 54.900 12.020 54.910 ;
        RECT 9.860 54.670 12.020 54.900 ;
        RECT 17.700 54.770 18.010 54.860 ;
        RECT 17.110 54.670 18.010 54.770 ;
        RECT 9.860 54.600 18.010 54.670 ;
        RECT 9.860 54.540 17.280 54.600 ;
        RECT 9.860 53.840 10.480 54.540 ;
        RECT 11.650 54.500 17.280 54.540 ;
        RECT 17.700 54.530 18.010 54.600 ;
        RECT 11.650 53.840 12.020 53.880 ;
        RECT 9.330 53.750 12.020 53.840 ;
        RECT 17.710 53.780 18.020 53.870 ;
        RECT 17.180 53.750 18.020 53.780 ;
        RECT 9.330 53.610 18.020 53.750 ;
        RECT 9.330 53.580 17.280 53.610 ;
        RECT 9.330 53.470 12.020 53.580 ;
        RECT 17.710 53.540 18.020 53.610 ;
        RECT 9.330 53.360 10.480 53.470 ;
        RECT 9.330 52.910 10.440 53.360 ;
        RECT 11.650 52.910 12.020 52.950 ;
        RECT 9.330 52.830 12.020 52.910 ;
        RECT 9.330 52.800 17.280 52.830 ;
        RECT 9.330 52.790 17.320 52.800 ;
        RECT 17.710 52.790 18.020 52.880 ;
        RECT 9.330 52.660 18.020 52.790 ;
        RECT 9.330 52.540 12.020 52.660 ;
        RECT 17.180 52.620 18.020 52.660 ;
        RECT 17.710 52.550 18.020 52.620 ;
        RECT 9.330 52.500 10.230 52.540 ;
        RECT 0.720 47.950 1.990 48.830 ;
        RECT 9.330 47.950 9.700 52.500 ;
        RECT 0.720 47.580 9.700 47.950 ;
        RECT 0.720 46.950 1.990 47.580 ;
    END
  END DRAIN3N
  PIN SOURCEP
    ANTENNAGATEAREA 0.652600 ;
    ANTENNADIFFAREA 5.759000 ;
    PORT
      LAYER met2 ;
        RECT 0.000 56.790 1.270 58.250 ;
        RECT 11.350 56.790 11.650 56.800 ;
        RECT 20.940 56.790 21.230 56.810 ;
        RECT 0.000 56.400 21.260 56.790 ;
        RECT 0.000 56.370 1.270 56.400 ;
        RECT 20.940 56.380 21.230 56.400 ;
        RECT 20.920 51.770 21.240 51.800 ;
        RECT 19.110 51.570 21.340 51.770 ;
        RECT 20.920 51.540 21.240 51.570 ;
        RECT 20.930 50.810 21.250 50.840 ;
        RECT 19.110 50.610 21.340 50.810 ;
        RECT 20.930 50.580 21.250 50.610 ;
        RECT 20.920 49.850 21.240 49.880 ;
        RECT 19.100 49.650 21.340 49.850 ;
        RECT 20.920 49.620 21.240 49.650 ;
        RECT 21.090 30.770 21.400 30.840 ;
        RECT 21.090 30.560 22.080 30.770 ;
        RECT 21.090 30.510 21.400 30.560 ;
        RECT 18.550 28.000 21.530 28.020 ;
        RECT 18.550 27.860 21.850 28.000 ;
        RECT 18.070 27.810 21.850 27.860 ;
        RECT 18.070 27.650 21.240 27.810 ;
        RECT 21.530 27.680 21.850 27.810 ;
        RECT 18.070 26.830 18.280 27.650 ;
        RECT 20.920 27.630 21.240 27.650 ;
        RECT 20.930 27.610 21.220 27.630 ;
        RECT 21.130 25.610 21.440 25.680 ;
        RECT 21.130 25.400 22.080 25.610 ;
        RECT 21.130 25.350 21.440 25.400 ;
        RECT 13.930 13.420 14.240 13.430 ;
        RECT 15.030 13.420 15.340 13.430 ;
        RECT 16.130 13.420 16.440 13.430 ;
        RECT 13.900 13.100 17.060 13.420 ;
        RECT 16.740 12.060 17.060 13.100 ;
        RECT 13.900 11.730 17.060 12.060 ;
        RECT 13.930 9.280 14.240 9.290 ;
        RECT 16.740 9.280 17.060 11.730 ;
        RECT 20.860 9.280 21.170 9.300 ;
        RECT 13.910 8.940 21.170 9.280 ;
        RECT 20.860 8.920 21.170 8.940 ;
    END
  END SOURCEP
  PIN GATE1
    PORT
      LAYER met2 ;
        RECT 57.060 58.640 57.380 58.680 ;
        RECT 72.710 58.640 73.990 58.740 ;
        RECT 57.060 58.430 73.990 58.640 ;
        RECT 57.060 58.400 57.380 58.430 ;
    END
  END GATE1
  PIN VINJ
    PORT
      LAYER met2 ;
        RECT 0.620 68.190 3.100 68.200 ;
        RECT 0.620 67.800 4.570 68.190 ;
        RECT 2.890 67.430 4.570 67.800 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.320 59.790 0.830 59.910 ;
        RECT 0.320 59.500 3.420 59.790 ;
        RECT 0.830 59.490 3.420 59.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.200 65.070 54.930 71.940 ;
        RECT 54.360 54.680 54.530 65.070 ;
      LAYER via ;
        RECT 54.230 65.110 54.670 65.550 ;
    END
  END VINJ
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 2.770 64.390 4.300 64.550 ;
        RECT 0.960 64.060 4.300 64.390 ;
        RECT 0.960 63.990 3.230 64.060 ;
        RECT 0.960 63.790 1.360 63.990 ;
        RECT 0.610 63.390 1.360 63.790 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.350 71.790 60.330 71.940 ;
        RECT 59.360 64.540 60.330 71.790 ;
        RECT 59.340 64.070 60.350 64.540 ;
      LAYER via ;
        RECT 59.370 64.110 60.320 64.520 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 50.840 24.100 51.100 24.170 ;
        RECT 51.580 24.100 51.840 24.170 ;
        RECT 50.840 23.070 51.840 24.100 ;
        RECT 50.600 23.060 51.100 23.070 ;
        RECT 50.320 22.750 51.100 23.060 ;
        RECT 50.320 22.740 50.640 22.750 ;
        RECT 50.840 21.730 51.100 22.750 ;
        RECT 50.600 21.720 51.100 21.730 ;
        RECT 50.310 21.410 51.100 21.720 ;
        RECT 50.310 21.400 50.630 21.410 ;
        RECT 50.840 18.960 51.100 21.410 ;
        RECT 50.600 18.950 51.100 18.960 ;
        RECT 50.310 18.640 51.100 18.950 ;
        RECT 50.310 18.630 50.630 18.640 ;
        RECT 50.840 17.980 51.100 18.640 ;
        RECT 51.580 23.060 52.080 23.070 ;
        RECT 51.580 22.750 52.360 23.060 ;
        RECT 51.580 21.720 51.840 22.750 ;
        RECT 52.040 22.740 52.360 22.750 ;
        RECT 51.580 21.400 52.370 21.720 ;
        RECT 51.580 18.950 51.840 21.400 ;
        RECT 51.580 18.630 52.370 18.950 ;
        RECT 51.580 18.000 51.840 18.630 ;
        RECT 50.830 17.640 51.110 17.980 ;
        RECT 51.570 17.660 51.850 18.000 ;
        RECT 50.840 16.230 51.100 17.640 ;
        RECT 51.580 16.230 51.840 17.660 ;
        RECT 50.840 12.800 51.840 16.230 ;
        RECT 50.360 12.760 52.290 12.800 ;
        RECT 49.820 11.570 52.290 12.760 ;
        RECT 49.820 0.080 50.760 11.570 ;
      LAYER via ;
        RECT 50.350 22.770 50.610 23.030 ;
        RECT 50.340 21.430 50.600 21.690 ;
        RECT 50.340 18.660 50.600 18.920 ;
        RECT 52.070 22.770 52.330 23.030 ;
        RECT 52.080 21.430 52.340 21.690 ;
        RECT 52.080 18.660 52.340 18.920 ;
        RECT 50.830 17.670 51.110 17.950 ;
        RECT 51.570 17.690 51.850 17.970 ;
        RECT 51.150 12.720 52.270 12.740 ;
        RECT 50.410 11.620 52.270 12.720 ;
        RECT 50.410 11.600 51.530 11.620 ;
    END
    PORT
      LAYER met1 ;
        RECT 60.650 24.020 60.910 24.200 ;
        RECT 61.390 24.020 61.650 24.200 ;
        RECT 60.650 23.090 61.650 24.020 ;
        RECT 60.130 22.770 60.910 23.090 ;
        RECT 60.650 21.750 60.910 22.770 ;
        RECT 60.120 21.430 60.910 21.750 ;
        RECT 60.650 18.980 60.910 21.430 ;
        RECT 60.120 18.660 60.910 18.980 ;
        RECT 60.650 17.980 60.910 18.660 ;
        RECT 61.390 22.770 62.170 23.090 ;
        RECT 61.390 21.740 61.650 22.770 ;
        RECT 61.860 21.740 62.180 21.750 ;
        RECT 61.390 21.430 62.180 21.740 ;
        RECT 61.390 21.420 61.890 21.430 ;
        RECT 61.390 18.980 61.650 21.420 ;
        RECT 61.390 18.660 62.180 18.980 ;
        RECT 60.640 17.640 60.920 17.980 ;
        RECT 60.650 16.460 60.910 17.640 ;
        RECT 61.390 16.460 61.650 18.660 ;
        RECT 60.650 12.860 61.650 16.460 ;
        RECT 60.650 12.820 62.670 12.860 ;
        RECT 60.170 11.540 62.670 12.820 ;
        RECT 61.780 1.540 62.670 11.540 ;
        RECT 61.780 0.810 62.700 1.540 ;
        RECT 61.750 0.080 62.670 0.810 ;
      LAYER via ;
        RECT 60.160 22.800 60.420 23.060 ;
        RECT 60.150 21.460 60.410 21.720 ;
        RECT 60.150 18.690 60.410 18.950 ;
        RECT 61.880 22.800 62.140 23.060 ;
        RECT 61.890 21.460 62.150 21.720 ;
        RECT 61.890 18.690 62.150 18.950 ;
        RECT 60.640 17.670 60.920 17.950 ;
        RECT 60.220 11.570 62.080 12.760 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 0.000 69.190 4.530 75.180 ;
        RECT 6.460 65.900 10.460 67.540 ;
        RECT 17.230 67.000 19.940 67.040 ;
        RECT 17.220 65.350 19.940 67.000 ;
        RECT 22.420 65.300 24.640 66.990 ;
        RECT 6.460 61.550 10.460 64.740 ;
        RECT 12.460 64.010 12.730 64.190 ;
        RECT 17.230 64.010 19.940 64.050 ;
        RECT 17.220 61.350 19.940 64.010 ;
        RECT 76.230 59.360 77.960 61.260 ;
        RECT 76.230 55.220 77.960 57.120 ;
        RECT 110.860 55.490 112.590 57.390 ;
        RECT 85.100 53.070 85.420 53.370 ;
        RECT 59.840 48.260 61.570 51.830 ;
        RECT 91.710 51.220 92.130 51.290 ;
        RECT 63.790 49.230 63.800 50.420 ;
        RECT 63.790 49.180 63.840 49.230 ;
        RECT 63.790 49.080 63.850 49.180 ;
        RECT 60.440 47.930 61.000 48.260 ;
        RECT 63.800 47.960 63.850 49.080 ;
        RECT 96.360 49.070 98.090 52.640 ;
        RECT 80.830 48.570 82.110 48.710 ;
        RECT 79.970 48.530 82.110 48.570 ;
        RECT 65.470 44.390 67.200 47.960 ;
        RECT 69.220 46.320 71.940 47.970 ;
        RECT 79.970 46.670 81.700 48.530 ;
        RECT 69.220 46.280 71.930 46.320 ;
        RECT 78.310 45.770 78.760 46.000 ;
        RECT 69.220 44.950 71.930 44.990 ;
        RECT 66.040 44.060 66.600 44.390 ;
        RECT 54.020 43.160 54.100 43.340 ;
        RECT 69.220 43.300 71.940 44.950 ;
        RECT 79.990 44.260 81.720 45.180 ;
        RECT 79.990 41.270 82.460 44.260 ;
        RECT 82.550 43.110 83.830 48.790 ;
        RECT 96.930 48.740 97.490 49.070 ;
        RECT 108.370 47.140 111.130 48.750 ;
        RECT 111.490 45.950 113.350 48.940 ;
        RECT 111.490 42.900 113.350 45.890 ;
        RECT 79.990 41.210 81.720 41.270 ;
        RECT 59.520 34.690 61.750 41.180 ;
        RECT 65.430 39.850 65.550 40.030 ;
        RECT 64.340 39.500 64.930 39.610 ;
        RECT 66.050 39.500 66.640 39.610 ;
        RECT 63.770 37.260 67.210 39.100 ;
        RECT 64.340 36.220 64.930 36.410 ;
        RECT 66.050 36.220 66.640 36.410 ;
        RECT 69.230 34.690 71.460 41.180 ;
        RECT 79.990 38.690 82.460 41.210 ;
        RECT 80.600 38.220 82.460 38.690 ;
        RECT 61.730 34.130 62.320 34.290 ;
        RECT 61.160 31.890 62.890 33.730 ;
        RECT 60.750 31.490 61.130 31.590 ;
        RECT 64.780 31.450 65.180 31.590 ;
        RECT 61.730 30.890 62.320 31.040 ;
        RECT 19.150 27.760 21.520 27.960 ;
        RECT 19.150 25.790 22.080 27.760 ;
        RECT 19.150 25.090 21.520 25.790 ;
        RECT 102.210 16.300 103.060 17.910 ;
        RECT 102.210 1.810 103.060 3.420 ;
      LAYER li1 ;
        RECT 6.800 66.230 10.110 67.210 ;
        RECT 12.050 65.590 12.220 65.920 ;
        RECT 12.730 65.590 12.900 65.920 ;
        RECT 19.410 65.870 19.640 66.560 ;
        RECT 24.110 65.820 24.340 66.510 ;
        RECT 12.120 65.030 12.290 65.380 ;
        RECT 12.750 65.070 13.070 65.110 ;
        RECT 11.390 64.990 12.290 65.030 ;
        RECT 11.380 64.800 12.290 64.990 ;
        RECT 12.740 64.880 13.070 65.070 ;
        RECT 13.440 65.060 13.760 65.100 ;
        RECT 12.750 64.850 13.070 64.880 ;
        RECT 13.430 64.870 13.760 65.060 ;
        RECT 13.440 64.840 13.760 64.870 ;
        RECT 11.390 64.770 12.290 64.800 ;
        RECT 20.620 64.790 20.790 64.810 ;
        RECT 6.800 63.430 10.110 64.410 ;
        RECT 6.800 61.880 10.110 62.860 ;
        RECT 10.750 61.910 10.920 64.560 ;
        RECT 12.120 64.370 12.290 64.770 ;
        RECT 17.730 64.620 20.790 64.790 ;
        RECT 20.620 63.970 20.790 64.620 ;
        RECT 20.620 63.800 21.890 63.970 ;
        RECT 19.410 62.880 19.640 63.570 ;
        RECT 10.750 61.370 10.930 61.910 ;
        RECT 19.410 61.870 19.640 62.560 ;
        RECT 20.620 61.390 20.790 63.800 ;
        RECT 23.360 62.150 23.530 63.040 ;
        RECT 10.670 61.330 10.990 61.370 ;
        RECT 20.530 61.350 20.850 61.390 ;
        RECT 10.660 61.140 10.990 61.330 ;
        RECT 20.520 61.160 20.850 61.350 ;
        RECT 10.670 61.110 10.990 61.140 ;
        RECT 20.530 61.130 20.850 61.160 ;
        RECT 19.820 60.140 21.340 60.150 ;
        RECT 19.820 59.350 21.370 60.140 ;
        RECT 40.910 58.090 41.260 58.190 ;
        RECT 44.670 58.180 44.960 58.200 ;
        RECT 44.500 58.140 44.960 58.180 ;
        RECT 43.520 58.120 44.960 58.140 ;
        RECT 42.570 58.090 43.030 58.120 ;
        RECT 39.500 57.920 40.260 58.090 ;
        RECT 40.510 57.920 41.680 58.090 ;
        RECT 41.920 57.950 43.030 58.090 ;
        RECT 43.480 57.960 44.960 58.120 ;
        RECT 43.480 57.950 44.670 57.960 ;
        RECT 41.920 57.920 42.740 57.950 ;
        RECT 39.500 57.910 39.730 57.920 ;
        RECT 39.460 57.470 39.730 57.910 ;
        RECT 42.480 57.780 42.740 57.920 ;
        RECT 40.940 57.470 41.270 57.730 ;
        RECT 42.480 57.610 43.660 57.780 ;
        RECT 42.480 57.470 42.740 57.610 ;
        RECT 38.910 57.330 39.080 57.390 ;
        RECT 38.880 57.110 39.100 57.330 ;
        RECT 39.430 57.290 39.760 57.470 ;
        RECT 40.010 57.300 42.170 57.470 ;
        RECT 42.410 57.300 42.740 57.470 ;
        RECT 42.570 57.250 42.740 57.300 ;
        RECT 43.030 57.110 43.240 57.440 ;
        RECT 43.480 57.170 43.660 57.610 ;
        RECT 45.290 57.510 45.460 58.270 ;
        RECT 45.660 58.120 46.110 58.270 ;
        RECT 45.660 57.950 46.260 58.120 ;
        RECT 46.720 57.940 47.050 58.110 ;
        RECT 45.080 57.500 45.460 57.510 ;
        RECT 45.080 57.440 45.550 57.500 ;
        RECT 46.800 57.480 46.980 57.940 ;
        RECT 44.210 57.330 45.550 57.440 ;
        RECT 44.210 57.270 45.470 57.330 ;
        RECT 46.020 57.310 46.980 57.480 ;
        RECT 45.080 57.220 45.470 57.270 ;
        RECT 38.910 57.060 39.080 57.110 ;
        RECT 40.910 56.340 41.260 56.440 ;
        RECT 44.670 56.430 44.960 56.450 ;
        RECT 44.500 56.390 44.960 56.430 ;
        RECT 43.520 56.370 44.960 56.390 ;
        RECT 42.570 56.340 43.030 56.370 ;
        RECT 39.500 56.170 40.260 56.340 ;
        RECT 40.510 56.170 41.680 56.340 ;
        RECT 41.920 56.200 43.030 56.340 ;
        RECT 43.480 56.210 44.960 56.370 ;
        RECT 43.480 56.200 44.670 56.210 ;
        RECT 41.920 56.170 42.740 56.200 ;
        RECT 39.500 56.160 39.730 56.170 ;
        RECT 39.460 55.720 39.730 56.160 ;
        RECT 42.480 56.030 42.740 56.170 ;
        RECT 40.940 55.720 41.270 55.980 ;
        RECT 42.480 55.860 43.660 56.030 ;
        RECT 42.480 55.720 42.740 55.860 ;
        RECT 38.910 55.580 39.080 55.640 ;
        RECT 38.880 55.360 39.100 55.580 ;
        RECT 39.430 55.540 39.760 55.720 ;
        RECT 40.010 55.550 42.170 55.720 ;
        RECT 42.410 55.550 42.740 55.720 ;
        RECT 42.570 55.500 42.740 55.550 ;
        RECT 43.030 55.360 43.240 55.690 ;
        RECT 43.480 55.420 43.660 55.860 ;
        RECT 45.290 55.760 45.460 56.520 ;
        RECT 45.660 56.370 46.110 56.520 ;
        RECT 45.660 56.200 46.260 56.370 ;
        RECT 46.720 56.190 47.050 56.360 ;
        RECT 67.790 56.190 68.460 57.060 ;
        RECT 80.070 56.300 82.170 57.060 ;
        RECT 82.830 56.680 83.360 56.850 ;
        RECT 83.500 56.710 83.690 56.940 ;
        RECT 83.780 56.660 84.660 56.830 ;
        RECT 80.070 56.210 82.280 56.300 ;
        RECT 45.080 55.750 45.460 55.760 ;
        RECT 45.080 55.690 45.550 55.750 ;
        RECT 46.800 55.730 46.980 56.190 ;
        RECT 81.340 55.970 81.560 56.210 ;
        RECT 81.340 55.960 81.550 55.970 ;
        RECT 81.720 55.790 81.910 55.800 ;
        RECT 44.210 55.580 45.550 55.690 ;
        RECT 44.210 55.520 45.470 55.580 ;
        RECT 46.020 55.560 46.980 55.730 ;
        RECT 45.080 55.470 45.470 55.520 ;
        RECT 81.710 55.500 81.910 55.790 ;
        RECT 38.910 55.310 39.080 55.360 ;
        RECT 81.650 55.170 81.920 55.500 ;
        RECT 18.020 54.820 18.220 54.860 ;
        RECT 17.710 54.560 18.220 54.820 ;
        RECT 18.020 54.530 18.220 54.560 ;
        RECT 18.610 54.830 18.810 54.860 ;
        RECT 18.610 54.790 19.120 54.830 ;
        RECT 18.610 54.600 19.130 54.790 ;
        RECT 18.610 54.570 19.120 54.600 ;
        RECT 40.910 54.590 41.260 54.690 ;
        RECT 44.670 54.680 44.960 54.700 ;
        RECT 44.500 54.640 44.960 54.680 ;
        RECT 43.520 54.620 44.960 54.640 ;
        RECT 42.570 54.590 43.030 54.620 ;
        RECT 18.610 54.530 18.810 54.570 ;
        RECT 39.500 54.420 40.260 54.590 ;
        RECT 40.510 54.420 41.680 54.590 ;
        RECT 41.920 54.450 43.030 54.590 ;
        RECT 43.480 54.460 44.960 54.620 ;
        RECT 43.480 54.450 44.670 54.460 ;
        RECT 41.920 54.420 42.740 54.450 ;
        RECT 39.500 54.410 39.730 54.420 ;
        RECT 17.440 54.320 17.800 54.390 ;
        RECT 17.280 54.220 17.800 54.320 ;
        RECT 19.310 54.280 19.480 54.330 ;
        RECT 19.300 54.250 19.480 54.280 ;
        RECT 17.280 54.140 17.650 54.220 ;
        RECT 17.280 54.090 17.610 54.140 ;
        RECT 17.280 54.060 17.600 54.090 ;
        RECT 19.300 54.000 19.730 54.250 ;
        RECT 19.800 54.090 19.990 54.320 ;
        RECT 19.300 53.970 19.490 54.000 ;
        RECT 39.460 53.970 39.730 54.410 ;
        RECT 42.480 54.280 42.740 54.420 ;
        RECT 40.940 53.970 41.270 54.230 ;
        RECT 42.480 54.110 43.660 54.280 ;
        RECT 42.480 53.970 42.740 54.110 ;
        RECT 19.310 53.940 19.490 53.970 ;
        RECT 18.030 53.830 18.230 53.870 ;
        RECT 17.720 53.570 18.230 53.830 ;
        RECT 18.030 53.540 18.230 53.570 ;
        RECT 18.620 53.840 18.820 53.870 ;
        RECT 18.620 53.800 19.130 53.840 ;
        RECT 38.910 53.830 39.080 53.890 ;
        RECT 18.620 53.610 19.140 53.800 ;
        RECT 38.880 53.610 39.100 53.830 ;
        RECT 39.430 53.790 39.760 53.970 ;
        RECT 40.010 53.800 42.170 53.970 ;
        RECT 42.410 53.800 42.740 53.970 ;
        RECT 42.570 53.750 42.740 53.800 ;
        RECT 43.030 53.610 43.240 53.940 ;
        RECT 43.480 53.670 43.660 54.110 ;
        RECT 45.290 54.010 45.460 54.770 ;
        RECT 45.660 54.620 46.110 54.770 ;
        RECT 82.110 54.690 82.280 56.210 ;
        RECT 82.940 55.200 83.110 56.290 ;
        RECT 83.970 56.270 84.160 56.380 ;
        RECT 83.530 56.150 84.160 56.270 ;
        RECT 84.490 56.270 84.660 56.660 ;
        RECT 83.530 56.100 84.080 56.150 ;
        RECT 84.490 56.100 85.230 56.270 ;
        RECT 86.290 55.480 86.520 56.000 ;
        RECT 83.530 55.310 86.520 55.480 ;
        RECT 82.710 55.160 83.110 55.200 ;
        RECT 82.700 54.970 83.110 55.160 ;
        RECT 91.490 55.120 92.040 55.550 ;
        RECT 82.710 54.940 83.110 54.970 ;
        RECT 45.660 54.450 46.260 54.620 ;
        RECT 46.720 54.440 47.050 54.610 ;
        RECT 82.100 54.500 82.280 54.690 ;
        RECT 82.940 54.600 83.110 54.940 ;
        RECT 83.500 54.720 83.690 54.950 ;
        RECT 83.530 54.520 83.880 54.690 ;
        RECT 45.080 54.000 45.460 54.010 ;
        RECT 45.080 53.940 45.550 54.000 ;
        RECT 46.800 53.980 46.980 54.440 ;
        RECT 84.360 54.370 84.570 54.800 ;
        RECT 84.880 54.520 85.220 54.690 ;
        RECT 84.380 54.350 84.550 54.370 ;
        RECT 44.210 53.830 45.550 53.940 ;
        RECT 44.210 53.770 45.470 53.830 ;
        RECT 46.020 53.810 46.980 53.980 ;
        RECT 82.100 53.780 82.280 53.970 ;
        RECT 83.530 53.880 83.880 53.950 ;
        RECT 45.080 53.720 45.470 53.770 ;
        RECT 18.620 53.580 19.130 53.610 ;
        RECT 18.620 53.540 18.820 53.580 ;
        RECT 38.910 53.560 39.080 53.610 ;
        RECT 17.260 53.230 17.810 53.400 ;
        RECT 17.260 53.170 17.590 53.230 ;
        RECT 17.260 53.140 17.580 53.170 ;
        RECT 18.030 52.840 18.230 52.880 ;
        RECT 17.720 52.580 18.230 52.840 ;
        RECT 18.030 52.550 18.230 52.580 ;
        RECT 18.620 52.850 18.820 52.880 ;
        RECT 18.620 52.810 19.130 52.850 ;
        RECT 40.910 52.840 41.260 52.940 ;
        RECT 44.670 52.930 44.960 52.950 ;
        RECT 44.500 52.890 44.960 52.930 ;
        RECT 43.520 52.870 44.960 52.890 ;
        RECT 42.570 52.840 43.030 52.870 ;
        RECT 18.620 52.620 19.140 52.810 ;
        RECT 39.500 52.670 40.260 52.840 ;
        RECT 40.510 52.670 41.680 52.840 ;
        RECT 41.920 52.700 43.030 52.840 ;
        RECT 43.480 52.710 44.960 52.870 ;
        RECT 43.480 52.700 44.670 52.710 ;
        RECT 41.920 52.670 42.740 52.700 ;
        RECT 39.500 52.660 39.730 52.670 ;
        RECT 18.620 52.590 19.130 52.620 ;
        RECT 18.620 52.550 18.820 52.590 ;
        RECT 18.740 52.420 19.060 52.460 ;
        RECT 17.240 52.240 17.810 52.410 ;
        RECT 18.740 52.400 19.070 52.420 ;
        RECT 17.240 52.180 17.570 52.240 ;
        RECT 18.740 52.200 19.360 52.400 ;
        RECT 17.240 52.150 17.560 52.180 ;
        RECT 19.190 52.070 19.360 52.200 ;
        RECT 19.870 52.360 20.040 52.400 ;
        RECT 19.870 52.320 20.360 52.360 ;
        RECT 19.870 52.130 20.370 52.320 ;
        RECT 39.460 52.220 39.730 52.660 ;
        RECT 42.480 52.530 42.740 52.670 ;
        RECT 40.940 52.220 41.270 52.480 ;
        RECT 42.480 52.360 43.660 52.530 ;
        RECT 42.480 52.220 42.740 52.360 ;
        RECT 19.870 52.100 20.360 52.130 ;
        RECT 19.870 52.070 20.040 52.100 ;
        RECT 38.910 52.080 39.080 52.140 ;
        RECT 18.550 51.960 18.980 51.980 ;
        RECT 18.530 51.790 18.980 51.960 ;
        RECT 38.880 51.860 39.100 52.080 ;
        RECT 39.430 52.040 39.760 52.220 ;
        RECT 40.010 52.050 42.170 52.220 ;
        RECT 42.410 52.050 42.740 52.220 ;
        RECT 42.570 52.000 42.740 52.050 ;
        RECT 43.030 51.860 43.240 52.190 ;
        RECT 43.480 51.920 43.660 52.360 ;
        RECT 45.290 52.260 45.460 53.020 ;
        RECT 45.660 52.870 46.110 53.020 ;
        RECT 81.650 52.970 81.920 53.300 ;
        RECT 45.660 52.700 46.260 52.870 ;
        RECT 46.720 52.690 47.050 52.860 ;
        RECT 45.080 52.250 45.460 52.260 ;
        RECT 45.080 52.190 45.550 52.250 ;
        RECT 46.800 52.230 46.980 52.690 ;
        RECT 81.710 52.680 81.910 52.970 ;
        RECT 81.720 52.670 81.910 52.680 ;
        RECT 81.340 52.500 81.550 52.510 ;
        RECT 44.210 52.080 45.550 52.190 ;
        RECT 44.210 52.020 45.470 52.080 ;
        RECT 46.020 52.060 46.980 52.230 ;
        RECT 45.080 51.970 45.470 52.020 ;
        RECT 50.460 51.900 50.660 52.250 ;
        RECT 51.940 52.000 52.470 52.170 ;
        RECT 50.450 51.870 50.660 51.900 ;
        RECT 38.910 51.810 39.080 51.860 ;
        RECT 18.550 51.770 18.980 51.790 ;
        RECT 18.740 51.430 19.060 51.470 ;
        RECT 18.740 51.410 19.070 51.430 ;
        RECT 18.740 51.210 19.360 51.410 ;
        RECT 19.190 51.080 19.360 51.210 ;
        RECT 19.870 51.370 20.040 51.410 ;
        RECT 19.870 51.330 20.360 51.370 ;
        RECT 19.870 51.140 20.370 51.330 ;
        RECT 38.910 51.290 39.080 51.340 ;
        RECT 19.870 51.110 20.360 51.140 ;
        RECT 19.870 51.080 20.040 51.110 ;
        RECT 38.880 51.070 39.100 51.290 ;
        RECT 38.910 51.010 39.080 51.070 ;
        RECT 18.550 50.970 18.980 50.990 ;
        RECT 18.530 50.800 18.980 50.970 ;
        RECT 39.430 50.930 39.760 51.110 ;
        RECT 42.570 51.100 42.740 51.150 ;
        RECT 40.010 50.930 42.170 51.100 ;
        RECT 42.410 50.930 42.740 51.100 ;
        RECT 43.030 50.960 43.240 51.290 ;
        RECT 18.550 50.780 18.980 50.800 ;
        RECT 39.460 50.490 39.730 50.930 ;
        RECT 40.940 50.670 41.270 50.930 ;
        RECT 42.480 50.790 42.740 50.930 ;
        RECT 43.480 50.790 43.660 51.230 ;
        RECT 45.080 51.130 45.470 51.180 ;
        RECT 44.210 51.070 45.470 51.130 ;
        RECT 44.210 50.960 45.550 51.070 ;
        RECT 45.080 50.900 45.550 50.960 ;
        RECT 46.020 50.920 46.980 51.090 ;
        RECT 45.080 50.890 45.460 50.900 ;
        RECT 39.500 50.480 39.730 50.490 ;
        RECT 42.480 50.620 43.660 50.790 ;
        RECT 42.480 50.480 42.740 50.620 ;
        RECT 18.740 50.440 19.060 50.480 ;
        RECT 18.740 50.420 19.070 50.440 ;
        RECT 18.740 50.290 19.360 50.420 ;
        RECT 19.870 50.380 20.040 50.420 ;
        RECT 19.870 50.340 20.360 50.380 ;
        RECT 18.740 50.220 19.520 50.290 ;
        RECT 19.190 50.200 19.520 50.220 ;
        RECT 19.190 50.090 19.580 50.200 ;
        RECT 19.870 50.150 20.370 50.340 ;
        RECT 39.500 50.310 40.260 50.480 ;
        RECT 40.510 50.310 41.680 50.480 ;
        RECT 41.920 50.450 42.740 50.480 ;
        RECT 41.920 50.310 43.030 50.450 ;
        RECT 40.910 50.210 41.260 50.310 ;
        RECT 42.570 50.280 43.030 50.310 ;
        RECT 43.480 50.440 44.670 50.450 ;
        RECT 43.480 50.280 44.960 50.440 ;
        RECT 43.520 50.260 44.960 50.280 ;
        RECT 44.500 50.220 44.960 50.260 ;
        RECT 44.670 50.200 44.960 50.220 ;
        RECT 19.870 50.120 20.360 50.150 ;
        RECT 45.290 50.130 45.460 50.890 ;
        RECT 46.800 50.460 46.980 50.920 ;
        RECT 47.970 50.910 48.140 51.330 ;
        RECT 50.450 51.290 50.670 51.870 ;
        RECT 50.450 51.280 50.660 51.290 ;
        RECT 48.780 51.210 49.020 51.240 ;
        RECT 51.220 51.210 51.390 51.620 ;
        RECT 48.450 51.040 49.020 51.210 ;
        RECT 49.260 51.040 50.600 51.210 ;
        RECT 50.830 51.110 51.020 51.120 ;
        RECT 48.780 51.000 49.020 51.040 ;
        RECT 50.820 50.820 51.020 51.110 ;
        RECT 51.050 51.040 52.010 51.210 ;
        RECT 52.050 51.090 52.220 51.610 ;
        RECT 54.660 51.570 59.720 52.400 ;
        RECT 81.340 51.920 81.560 52.500 ;
        RECT 82.110 52.170 82.280 53.780 ;
        RECT 82.940 53.510 83.110 53.870 ;
        RECT 83.510 53.780 83.880 53.880 ;
        RECT 83.970 53.830 84.160 54.060 ;
        RECT 84.970 53.950 85.140 54.520 ;
        RECT 89.250 54.370 89.440 54.690 ;
        RECT 89.250 54.280 89.530 54.370 ;
        RECT 85.890 54.140 89.530 54.280 ;
        RECT 85.890 54.100 89.440 54.140 ;
        RECT 84.250 53.920 84.300 53.930 ;
        RECT 84.880 53.920 85.220 53.950 ;
        RECT 84.250 53.840 85.220 53.920 ;
        RECT 84.210 53.780 85.220 53.840 ;
        RECT 83.510 53.650 83.700 53.780 ;
        RECT 84.210 53.720 85.050 53.780 ;
        RECT 89.250 53.680 89.440 54.100 ;
        RECT 82.700 53.470 83.110 53.510 ;
        RECT 82.690 53.280 83.110 53.470 ;
        RECT 91.490 53.390 92.040 53.820 ;
        RECT 108.580 53.750 108.790 54.180 ;
        RECT 108.600 53.730 108.770 53.750 ;
        RECT 109.100 53.610 109.290 53.720 ;
        RECT 109.100 53.490 109.520 53.610 ;
        RECT 109.000 53.440 109.520 53.490 ;
        RECT 109.870 53.440 111.770 53.620 ;
        RECT 112.150 53.450 112.500 53.620 ;
        RECT 112.600 53.610 112.790 53.720 ;
        RECT 112.600 53.490 112.930 53.610 ;
        RECT 109.000 53.390 109.190 53.440 ;
        RECT 82.700 53.250 83.110 53.280 ;
        RECT 108.850 53.340 109.190 53.390 ;
        RECT 108.850 53.270 109.410 53.340 ;
        RECT 110.360 53.320 110.690 53.440 ;
        RECT 112.680 53.410 112.930 53.490 ;
        RECT 112.760 53.390 112.930 53.410 ;
        RECT 112.040 53.350 112.240 53.390 ;
        RECT 82.940 52.180 83.110 53.250 ;
        RECT 108.720 53.240 109.410 53.270 ;
        RECT 83.530 53.060 86.460 53.160 ;
        RECT 108.680 53.080 109.410 53.240 ;
        RECT 108.680 53.060 109.020 53.080 ;
        RECT 83.530 52.990 86.520 53.060 ;
        RECT 85.550 52.670 85.720 52.730 ;
        RECT 83.960 52.370 84.150 52.480 ;
        RECT 85.530 52.460 85.740 52.670 ;
        RECT 85.550 52.390 85.720 52.460 ;
        RECT 86.290 52.370 86.520 52.990 ;
        RECT 105.460 52.810 105.990 52.980 ;
        RECT 107.270 52.710 107.470 53.060 ;
        RECT 108.680 53.020 108.890 53.060 ;
        RECT 108.680 52.740 108.850 53.020 ;
        RECT 110.030 52.910 110.200 53.070 ;
        RECT 111.010 53.000 111.200 53.110 ;
        RECT 111.810 53.100 112.240 53.350 ;
        RECT 111.810 53.090 112.330 53.100 ;
        RECT 110.890 52.990 111.200 53.000 ;
        RECT 109.900 52.870 110.220 52.910 ;
        RECT 110.640 52.880 111.200 52.990 ;
        RECT 111.530 52.910 111.700 53.070 ;
        RECT 112.040 53.060 112.330 53.090 ;
        RECT 112.140 52.990 112.330 53.060 ;
        RECT 107.270 52.680 107.480 52.710 ;
        RECT 83.530 52.250 84.150 52.370 ;
        RECT 83.530 52.200 84.070 52.250 ;
        RECT 84.420 52.200 85.230 52.370 ;
        RECT 81.340 51.890 81.550 51.920 ;
        RECT 59.170 51.490 59.650 51.570 ;
        RECT 81.350 51.540 81.550 51.890 ;
        RECT 83.530 51.860 83.720 51.970 ;
        RECT 84.420 51.860 84.610 52.200 ;
        RECT 82.830 51.620 83.360 51.790 ;
        RECT 83.530 51.740 84.610 51.860 ;
        RECT 83.650 51.680 84.610 51.740 ;
        RECT 47.900 50.690 48.070 50.730 ;
        RECT 47.840 50.520 48.070 50.690 ;
        RECT 50.740 50.590 51.030 50.820 ;
        RECT 51.220 50.770 51.390 51.040 ;
        RECT 51.560 51.030 51.730 51.040 ;
        RECT 52.050 50.830 52.380 51.090 ;
        RECT 51.190 50.590 51.530 50.770 ;
        RECT 45.660 50.280 46.260 50.450 ;
        RECT 46.720 50.290 47.050 50.460 ;
        RECT 45.660 50.130 46.110 50.280 ;
        RECT 47.900 50.170 48.070 50.520 ;
        RECT 48.140 50.300 48.330 50.530 ;
        RECT 48.430 50.420 48.800 50.590 ;
        RECT 49.260 50.420 52.010 50.590 ;
        RECT 19.870 50.090 20.040 50.120 ;
        RECT 19.350 50.010 19.580 50.090 ;
        RECT 51.220 50.010 51.390 50.420 ;
        RECT 18.550 49.980 18.980 50.000 ;
        RECT 18.530 49.810 18.980 49.980 ;
        RECT 51.210 49.820 51.390 50.010 ;
        RECT 52.050 49.920 52.220 50.830 ;
        RECT 52.540 50.350 52.710 51.280 ;
        RECT 52.940 50.440 53.110 51.330 ;
        RECT 57.290 50.630 57.520 51.320 ;
        RECT 59.170 51.240 59.640 51.490 ;
        RECT 96.780 51.250 97.330 51.680 ;
        RECT 100.410 51.440 100.640 52.130 ;
        RECT 105.710 51.900 105.880 52.420 ;
        RECT 105.550 51.640 105.880 51.900 ;
        RECT 60.600 50.440 61.150 50.870 ;
        RECT 99.380 50.500 99.570 50.820 ;
        RECT 105.710 50.730 105.880 51.640 ;
        RECT 106.540 50.820 106.710 52.430 ;
        RECT 107.260 52.100 107.480 52.680 ;
        RECT 109.900 52.680 110.230 52.870 ;
        RECT 110.640 52.820 111.020 52.880 ;
        RECT 111.470 52.870 111.790 52.910 ;
        RECT 112.140 52.870 112.480 52.990 ;
        RECT 111.470 52.700 111.800 52.870 ;
        RECT 112.190 52.820 112.480 52.870 ;
        RECT 112.040 52.700 112.240 52.730 ;
        RECT 109.900 52.650 110.220 52.680 ;
        RECT 111.470 52.650 112.240 52.700 ;
        RECT 109.250 52.510 109.330 52.650 ;
        RECT 109.240 52.470 109.560 52.510 ;
        RECT 109.230 52.280 109.560 52.470 ;
        RECT 111.630 52.440 112.240 52.650 ;
        RECT 111.630 52.410 111.800 52.440 ;
        RECT 112.040 52.400 112.240 52.440 ;
        RECT 112.630 52.400 113.180 53.390 ;
        RECT 114.000 53.240 114.630 53.410 ;
        RECT 114.000 53.140 114.390 53.240 ;
        RECT 114.000 53.110 114.380 53.140 ;
        RECT 114.000 52.960 114.360 53.110 ;
        RECT 113.650 52.790 114.360 52.960 ;
        RECT 109.240 52.250 109.560 52.280 ;
        RECT 113.650 52.120 114.350 52.350 ;
        RECT 107.270 52.090 107.480 52.100 ;
        RECT 108.150 51.950 108.470 51.980 ;
        RECT 106.910 51.920 107.100 51.930 ;
        RECT 106.910 51.630 107.110 51.920 ;
        RECT 108.150 51.760 108.480 51.950 ;
        RECT 113.600 51.890 114.350 52.120 ;
        RECT 111.630 51.850 111.800 51.880 ;
        RECT 112.040 51.850 112.240 51.890 ;
        RECT 111.630 51.760 112.240 51.850 ;
        RECT 108.150 51.720 108.470 51.760 ;
        RECT 109.900 51.730 110.220 51.760 ;
        RECT 106.900 51.300 107.190 51.630 ;
        RECT 108.680 51.390 108.850 51.670 ;
        RECT 109.900 51.540 110.230 51.730 ;
        RECT 111.470 51.590 112.240 51.760 ;
        RECT 109.900 51.500 110.220 51.540 ;
        RECT 110.640 51.530 111.020 51.590 ;
        RECT 111.470 51.540 111.800 51.590 ;
        RECT 112.040 51.560 112.480 51.590 ;
        RECT 112.190 51.540 112.480 51.560 ;
        RECT 108.680 51.350 108.890 51.390 ;
        RECT 108.680 51.330 108.910 51.350 ;
        RECT 110.030 51.340 110.200 51.500 ;
        RECT 110.640 51.420 111.200 51.530 ;
        RECT 111.470 51.500 111.790 51.540 ;
        RECT 110.890 51.410 111.200 51.420 ;
        RECT 108.680 51.310 108.940 51.330 ;
        RECT 108.680 51.260 109.020 51.310 ;
        RECT 111.010 51.300 111.200 51.410 ;
        RECT 111.530 51.340 111.700 51.500 ;
        RECT 112.140 51.420 112.480 51.540 ;
        RECT 112.140 51.310 112.330 51.420 ;
        RECT 108.680 51.200 109.170 51.260 ;
        RECT 112.040 51.200 112.240 51.230 ;
        RECT 108.680 51.170 109.190 51.200 ;
        RECT 108.720 51.140 109.190 51.170 ;
        RECT 108.850 51.090 109.190 51.140 ;
        RECT 108.970 51.080 109.190 51.090 ;
        RECT 108.980 51.050 109.190 51.080 ;
        RECT 106.540 50.630 106.720 50.820 ;
        RECT 99.290 50.410 99.570 50.500 ;
        RECT 99.290 50.270 102.930 50.410 ;
        RECT 99.380 50.230 102.930 50.270 ;
        RECT 18.550 49.790 18.980 49.810 ;
        RECT 38.910 49.540 39.080 49.590 ;
        RECT 38.880 49.320 39.100 49.540 ;
        RECT 38.910 49.260 39.080 49.320 ;
        RECT 39.430 49.180 39.760 49.360 ;
        RECT 42.570 49.350 42.740 49.400 ;
        RECT 40.010 49.180 42.170 49.350 ;
        RECT 42.410 49.180 42.740 49.350 ;
        RECT 43.030 49.210 43.240 49.540 ;
        RECT 39.460 48.740 39.730 49.180 ;
        RECT 40.940 48.920 41.270 49.180 ;
        RECT 42.480 49.040 42.740 49.180 ;
        RECT 43.480 49.040 43.660 49.480 ;
        RECT 45.080 49.380 45.470 49.430 ;
        RECT 47.900 49.410 48.070 49.760 ;
        RECT 58.360 49.690 58.550 50.010 ;
        RECT 44.210 49.320 45.470 49.380 ;
        RECT 44.210 49.210 45.550 49.320 ;
        RECT 45.080 49.150 45.550 49.210 ;
        RECT 46.020 49.170 46.980 49.340 ;
        RECT 47.840 49.240 48.070 49.410 ;
        RECT 48.140 49.400 48.330 49.630 ;
        RECT 58.360 49.600 58.640 49.690 ;
        RECT 48.430 49.340 48.800 49.510 ;
        RECT 49.260 49.340 52.010 49.510 ;
        RECT 47.900 49.200 48.070 49.240 ;
        RECT 45.080 49.140 45.460 49.150 ;
        RECT 39.500 48.730 39.730 48.740 ;
        RECT 42.480 48.870 43.660 49.040 ;
        RECT 42.480 48.730 42.740 48.870 ;
        RECT 39.500 48.560 40.260 48.730 ;
        RECT 40.510 48.560 41.680 48.730 ;
        RECT 41.920 48.700 42.740 48.730 ;
        RECT 41.920 48.560 43.030 48.700 ;
        RECT 40.910 48.460 41.260 48.560 ;
        RECT 42.570 48.530 43.030 48.560 ;
        RECT 43.480 48.690 44.670 48.700 ;
        RECT 43.480 48.530 44.960 48.690 ;
        RECT 43.520 48.510 44.960 48.530 ;
        RECT 44.500 48.470 44.960 48.510 ;
        RECT 44.670 48.450 44.960 48.470 ;
        RECT 45.290 48.380 45.460 49.140 ;
        RECT 46.800 48.710 46.980 49.170 ;
        RECT 51.190 49.160 51.530 49.340 ;
        RECT 51.210 49.100 51.390 49.160 ;
        RECT 45.660 48.530 46.260 48.700 ;
        RECT 46.720 48.540 47.050 48.710 ;
        RECT 47.970 48.600 48.140 49.020 ;
        RECT 48.780 48.890 49.020 48.930 ;
        RECT 51.220 48.890 51.390 49.100 ;
        RECT 51.560 48.890 51.730 48.900 ;
        RECT 48.450 48.720 49.020 48.890 ;
        RECT 49.260 48.720 50.600 48.890 ;
        RECT 51.050 48.720 52.010 48.890 ;
        RECT 48.780 48.690 49.020 48.720 ;
        RECT 45.660 48.380 46.110 48.530 ;
        RECT 50.740 48.290 51.030 48.620 ;
        RECT 38.910 47.790 39.080 47.840 ;
        RECT 38.880 47.570 39.100 47.790 ;
        RECT 38.910 47.510 39.080 47.570 ;
        RECT 39.430 47.430 39.760 47.610 ;
        RECT 42.570 47.600 42.740 47.650 ;
        RECT 40.010 47.430 42.170 47.600 ;
        RECT 42.410 47.430 42.740 47.600 ;
        RECT 43.030 47.460 43.240 47.790 ;
        RECT 39.460 46.990 39.730 47.430 ;
        RECT 40.940 47.170 41.270 47.430 ;
        RECT 42.480 47.290 42.740 47.430 ;
        RECT 43.480 47.290 43.660 47.730 ;
        RECT 47.970 47.710 48.140 48.130 ;
        RECT 48.780 48.010 49.020 48.040 ;
        RECT 48.450 47.840 49.020 48.010 ;
        RECT 49.260 47.840 50.600 48.010 ;
        RECT 50.820 48.000 51.020 48.290 ;
        RECT 51.220 48.010 51.390 48.720 ;
        RECT 52.050 48.330 52.220 49.190 ;
        RECT 52.540 48.650 52.710 49.580 ;
        RECT 52.940 48.600 53.110 49.490 ;
        RECT 55.000 49.460 58.640 49.600 ;
        RECT 96.780 49.520 97.330 49.950 ;
        RECT 99.380 49.810 99.570 50.230 ;
        RECT 55.000 49.420 58.550 49.460 ;
        RECT 58.360 49.000 58.550 49.420 ;
        RECT 60.600 48.710 61.150 49.140 ;
        RECT 77.960 48.660 78.130 48.710 ;
        RECT 81.150 48.670 81.350 48.710 ;
        RECT 52.050 48.070 52.380 48.330 ;
        RECT 50.830 47.990 51.020 48.000 ;
        RECT 51.050 47.840 52.010 48.010 ;
        RECT 48.780 47.800 49.020 47.840 ;
        RECT 50.450 47.820 50.660 47.830 ;
        RECT 45.080 47.630 45.470 47.680 ;
        RECT 44.210 47.570 45.470 47.630 ;
        RECT 44.210 47.460 45.550 47.570 ;
        RECT 45.080 47.400 45.550 47.460 ;
        RECT 46.020 47.420 46.980 47.590 ;
        RECT 47.900 47.490 48.070 47.530 ;
        RECT 45.080 47.390 45.460 47.400 ;
        RECT 39.500 46.980 39.730 46.990 ;
        RECT 42.480 47.120 43.660 47.290 ;
        RECT 42.480 46.980 42.740 47.120 ;
        RECT 39.500 46.810 40.260 46.980 ;
        RECT 40.510 46.810 41.680 46.980 ;
        RECT 41.920 46.950 42.740 46.980 ;
        RECT 41.920 46.810 43.030 46.950 ;
        RECT 40.910 46.710 41.260 46.810 ;
        RECT 42.570 46.780 43.030 46.810 ;
        RECT 43.480 46.940 44.670 46.950 ;
        RECT 43.480 46.780 44.960 46.940 ;
        RECT 43.520 46.760 44.960 46.780 ;
        RECT 44.500 46.720 44.960 46.760 ;
        RECT 44.670 46.700 44.960 46.720 ;
        RECT 45.290 46.630 45.460 47.390 ;
        RECT 46.800 46.960 46.980 47.420 ;
        RECT 47.840 47.320 48.070 47.490 ;
        RECT 50.450 47.390 50.670 47.820 ;
        RECT 51.220 47.570 51.390 47.840 ;
        RECT 51.560 47.830 51.730 47.840 ;
        RECT 51.190 47.390 51.530 47.570 ;
        RECT 52.050 47.500 52.220 48.070 ;
        RECT 47.900 46.970 48.070 47.320 ;
        RECT 48.140 47.100 48.330 47.330 ;
        RECT 48.430 47.220 48.800 47.390 ;
        RECT 49.260 47.220 52.010 47.390 ;
        RECT 50.450 47.210 50.660 47.220 ;
        RECT 45.660 46.780 46.260 46.950 ;
        RECT 46.720 46.790 47.050 46.960 ;
        RECT 50.460 46.860 50.660 47.210 ;
        RECT 52.540 47.150 52.710 48.080 ;
        RECT 52.940 47.240 53.110 48.130 ;
        RECT 57.290 47.690 57.520 48.420 ;
        RECT 77.960 48.400 78.520 48.660 ;
        RECT 80.920 48.410 81.350 48.670 ;
        RECT 77.960 48.380 78.130 48.400 ;
        RECT 81.150 48.380 81.350 48.410 ;
        RECT 74.570 48.130 75.100 48.300 ;
        RECT 76.380 48.030 76.580 48.380 ;
        RECT 76.380 48.000 76.590 48.030 ;
        RECT 59.330 47.560 59.670 47.810 ;
        RECT 59.330 47.480 59.680 47.560 ;
        RECT 51.940 46.940 52.470 47.110 ;
        RECT 45.660 46.630 46.110 46.780 ;
        RECT 54.630 46.630 59.680 47.480 ;
        RECT 65.890 46.570 66.440 47.000 ;
        RECT 69.520 46.760 69.750 47.450 ;
        RECT 74.820 47.220 74.990 47.740 ;
        RECT 74.660 46.960 74.990 47.220 ;
        RECT 47.900 46.210 48.070 46.560 ;
        RECT 38.910 46.040 39.080 46.090 ;
        RECT 47.840 46.040 48.070 46.210 ;
        RECT 48.140 46.200 48.330 46.430 ;
        RECT 48.430 46.140 48.800 46.310 ;
        RECT 49.260 46.140 52.010 46.310 ;
        RECT 38.880 45.820 39.100 46.040 ;
        RECT 38.910 45.760 39.080 45.820 ;
        RECT 39.430 45.680 39.760 45.860 ;
        RECT 42.570 45.850 42.740 45.900 ;
        RECT 40.010 45.680 42.170 45.850 ;
        RECT 42.410 45.680 42.740 45.850 ;
        RECT 43.030 45.710 43.240 46.040 ;
        RECT 47.900 46.000 48.070 46.040 ;
        RECT 39.460 45.240 39.730 45.680 ;
        RECT 40.940 45.420 41.270 45.680 ;
        RECT 42.480 45.540 42.740 45.680 ;
        RECT 43.480 45.540 43.660 45.980 ;
        RECT 51.190 45.960 51.530 46.140 ;
        RECT 45.080 45.880 45.470 45.930 ;
        RECT 44.210 45.820 45.470 45.880 ;
        RECT 44.210 45.710 45.550 45.820 ;
        RECT 45.080 45.650 45.550 45.710 ;
        RECT 46.020 45.670 46.980 45.840 ;
        RECT 45.080 45.640 45.460 45.650 ;
        RECT 39.500 45.230 39.730 45.240 ;
        RECT 42.480 45.370 43.660 45.540 ;
        RECT 42.480 45.230 42.740 45.370 ;
        RECT 39.500 45.060 40.260 45.230 ;
        RECT 40.510 45.060 41.680 45.230 ;
        RECT 41.920 45.200 42.740 45.230 ;
        RECT 41.920 45.060 43.030 45.200 ;
        RECT 40.910 44.960 41.260 45.060 ;
        RECT 42.570 45.030 43.030 45.060 ;
        RECT 43.480 45.190 44.670 45.200 ;
        RECT 43.480 45.030 44.960 45.190 ;
        RECT 43.520 45.010 44.960 45.030 ;
        RECT 44.500 44.970 44.960 45.010 ;
        RECT 44.670 44.950 44.960 44.970 ;
        RECT 45.290 44.880 45.460 45.640 ;
        RECT 46.800 45.210 46.980 45.670 ;
        RECT 47.970 45.400 48.140 45.820 ;
        RECT 48.780 45.690 49.020 45.730 ;
        RECT 51.560 45.690 51.730 45.700 ;
        RECT 48.450 45.520 49.020 45.690 ;
        RECT 49.260 45.520 50.600 45.690 ;
        RECT 51.050 45.520 52.010 45.690 ;
        RECT 48.780 45.490 49.020 45.520 ;
        RECT 52.540 45.450 52.710 46.380 ;
        RECT 52.940 45.400 53.110 46.290 ;
        RECT 45.660 45.030 46.260 45.200 ;
        RECT 46.720 45.040 47.050 45.210 ;
        RECT 62.510 45.130 62.710 46.140 ;
        RECT 68.260 45.730 68.680 46.140 ;
        RECT 74.820 46.050 74.990 46.960 ;
        RECT 75.650 46.140 75.820 47.750 ;
        RECT 76.370 47.420 76.590 48.000 ;
        RECT 80.740 48.020 80.910 48.060 ;
        RECT 81.150 48.020 81.350 48.050 ;
        RECT 78.360 47.830 78.440 47.970 ;
        RECT 78.350 47.790 78.670 47.830 ;
        RECT 78.340 47.600 78.670 47.790 ;
        RECT 80.740 47.760 81.350 48.020 ;
        RECT 80.740 47.730 80.910 47.760 ;
        RECT 81.150 47.720 81.350 47.760 ;
        RECT 81.740 47.720 82.290 48.710 ;
        RECT 83.110 48.560 83.740 48.730 ;
        RECT 83.110 48.460 83.500 48.560 ;
        RECT 100.410 48.500 100.640 49.230 ;
        RECT 105.710 49.140 105.880 50.000 ;
        RECT 105.550 48.880 105.880 49.140 ;
        RECT 83.110 48.430 83.490 48.460 ;
        RECT 83.110 48.280 83.470 48.430 ;
        RECT 105.710 48.310 105.880 48.880 ;
        RECT 106.540 49.910 106.720 50.100 ;
        RECT 106.540 48.300 106.710 49.910 ;
        RECT 108.270 49.850 108.450 50.910 ;
        RECT 108.580 50.230 108.790 50.980 ;
        RECT 109.000 50.970 109.190 51.050 ;
        RECT 110.360 50.970 110.690 51.090 ;
        RECT 109.000 50.920 109.520 50.970 ;
        RECT 109.100 50.800 109.520 50.920 ;
        RECT 109.100 50.700 109.290 50.800 ;
        RECT 109.870 50.790 111.770 50.970 ;
        RECT 111.810 50.960 112.240 51.200 ;
        RECT 111.810 50.940 112.500 50.960 ;
        RECT 112.040 50.900 112.500 50.940 ;
        RECT 112.630 50.920 113.180 51.890 ;
        RECT 113.650 51.470 114.350 51.890 ;
        RECT 114.110 51.110 114.430 51.150 ;
        RECT 114.110 51.050 114.440 51.110 ;
        RECT 112.150 50.790 112.500 50.900 ;
        RECT 112.600 50.900 113.180 50.920 ;
        RECT 113.640 50.920 114.440 51.050 ;
        RECT 112.600 50.800 112.930 50.900 ;
        RECT 113.640 50.890 114.430 50.920 ;
        RECT 113.640 50.870 114.340 50.890 ;
        RECT 108.880 50.690 109.290 50.700 ;
        RECT 112.600 50.690 112.790 50.800 ;
        RECT 108.880 50.670 109.200 50.690 ;
        RECT 108.880 50.520 109.210 50.670 ;
        RECT 108.880 50.440 109.290 50.520 ;
        RECT 108.880 50.360 109.050 50.440 ;
        RECT 108.830 50.290 109.050 50.360 ;
        RECT 109.100 50.410 109.290 50.440 ;
        RECT 109.100 50.290 109.520 50.410 ;
        RECT 108.830 50.240 109.520 50.290 ;
        RECT 109.870 50.240 111.770 50.420 ;
        RECT 112.150 50.390 112.500 50.420 ;
        RECT 112.040 50.350 112.500 50.390 ;
        RECT 111.810 50.250 112.500 50.350 ;
        RECT 112.600 50.410 112.790 50.520 ;
        RECT 112.600 50.390 112.930 50.410 ;
        RECT 114.100 50.390 114.420 50.430 ;
        RECT 112.600 50.290 113.180 50.390 ;
        RECT 108.830 50.070 109.190 50.240 ;
        RECT 110.360 50.120 110.690 50.240 ;
        RECT 111.810 50.090 112.240 50.250 ;
        RECT 108.720 50.040 109.190 50.070 ;
        RECT 112.040 50.060 112.240 50.090 ;
        RECT 108.680 50.010 109.190 50.040 ;
        RECT 108.680 49.950 109.170 50.010 ;
        RECT 108.680 49.900 109.020 49.950 ;
        RECT 108.680 49.880 108.940 49.900 ;
        RECT 108.680 49.860 108.910 49.880 ;
        RECT 108.680 49.820 108.890 49.860 ;
        RECT 108.680 49.540 108.850 49.820 ;
        RECT 109.320 49.690 109.400 49.770 ;
        RECT 109.460 49.690 109.650 49.810 ;
        RECT 110.030 49.710 110.200 49.870 ;
        RECT 111.010 49.800 111.200 49.910 ;
        RECT 110.890 49.790 111.200 49.800 ;
        RECT 109.320 49.600 109.650 49.690 ;
        RECT 109.460 49.580 109.650 49.600 ;
        RECT 109.900 49.670 110.220 49.710 ;
        RECT 110.640 49.680 111.200 49.790 ;
        RECT 111.530 49.740 111.700 49.870 ;
        RECT 112.140 49.790 112.330 49.900 ;
        RECT 111.530 49.710 111.800 49.740 ;
        RECT 112.140 49.730 112.480 49.790 ;
        RECT 111.470 49.700 111.800 49.710 ;
        RECT 112.040 49.700 112.480 49.730 ;
        RECT 109.900 49.480 110.230 49.670 ;
        RECT 110.640 49.620 111.020 49.680 ;
        RECT 111.470 49.620 112.480 49.700 ;
        RECT 109.900 49.450 110.220 49.480 ;
        RECT 111.470 49.450 112.240 49.620 ;
        RECT 111.630 49.440 112.240 49.450 ;
        RECT 106.900 49.100 107.190 49.430 ;
        RECT 111.630 49.410 111.800 49.440 ;
        RECT 112.040 49.400 112.240 49.440 ;
        RECT 112.630 49.400 113.180 50.290 ;
        RECT 113.640 50.210 114.430 50.390 ;
        RECT 114.100 50.200 114.430 50.210 ;
        RECT 114.100 50.170 114.420 50.200 ;
        RECT 113.650 49.530 114.350 49.790 ;
        RECT 113.600 49.300 114.350 49.530 ;
        RECT 106.910 48.810 107.110 49.100 ;
        RECT 113.650 48.910 114.350 49.300 ;
        RECT 111.630 48.850 111.800 48.880 ;
        RECT 112.040 48.850 112.240 48.890 ;
        RECT 106.910 48.800 107.100 48.810 ;
        RECT 107.270 48.630 107.480 48.640 ;
        RECT 82.760 48.110 83.470 48.280 ;
        RECT 107.260 48.050 107.480 48.630 ;
        RECT 111.630 48.590 112.240 48.850 ;
        RECT 111.630 48.560 111.800 48.590 ;
        RECT 112.040 48.560 112.240 48.590 ;
        RECT 109.900 48.530 110.220 48.560 ;
        RECT 111.470 48.550 111.800 48.560 ;
        RECT 111.470 48.530 111.790 48.550 ;
        RECT 107.270 48.020 107.480 48.050 ;
        RECT 108.680 48.190 108.850 48.470 ;
        RECT 109.900 48.340 110.230 48.530 ;
        RECT 109.900 48.300 110.220 48.340 ;
        RECT 110.640 48.330 111.020 48.390 ;
        RECT 111.470 48.340 111.800 48.530 ;
        RECT 108.680 48.150 108.890 48.190 ;
        RECT 108.680 48.130 108.910 48.150 ;
        RECT 110.030 48.140 110.200 48.300 ;
        RECT 110.640 48.220 111.200 48.330 ;
        RECT 111.470 48.300 111.790 48.340 ;
        RECT 110.890 48.210 111.200 48.220 ;
        RECT 108.680 48.110 108.940 48.130 ;
        RECT 108.680 48.060 109.020 48.110 ;
        RECT 111.010 48.100 111.200 48.210 ;
        RECT 111.530 48.140 111.700 48.300 ;
        RECT 111.900 48.230 112.080 48.470 ;
        RECT 112.190 48.340 112.480 48.390 ;
        RECT 112.140 48.230 112.480 48.340 ;
        RECT 111.900 48.220 112.480 48.230 ;
        RECT 111.900 48.200 112.330 48.220 ;
        RECT 111.810 48.110 112.330 48.200 ;
        RECT 105.460 47.750 105.990 47.920 ;
        RECT 107.270 47.670 107.470 48.020 ;
        RECT 108.680 48.000 109.170 48.060 ;
        RECT 108.680 47.970 109.190 48.000 ;
        RECT 108.720 47.940 109.190 47.970 ;
        RECT 111.810 47.940 112.240 48.110 ;
        RECT 108.850 47.890 109.190 47.940 ;
        RECT 111.900 47.900 112.240 47.940 ;
        RECT 112.630 47.900 113.180 48.890 ;
        RECT 113.650 48.300 114.360 48.470 ;
        RECT 114.000 48.020 114.360 48.300 ;
        RECT 108.970 47.880 109.190 47.890 ;
        RECT 108.980 47.850 109.190 47.880 ;
        RECT 109.000 47.770 109.190 47.850 ;
        RECT 110.360 47.770 110.690 47.890 ;
        RECT 109.000 47.720 109.520 47.770 ;
        RECT 78.350 47.570 78.670 47.600 ;
        RECT 82.760 47.440 83.460 47.670 ;
        RECT 109.100 47.600 109.520 47.720 ;
        RECT 109.100 47.490 109.290 47.600 ;
        RECT 109.870 47.590 111.770 47.770 ;
        RECT 108.600 47.460 108.770 47.480 ;
        RECT 76.380 47.410 76.590 47.420 ;
        RECT 77.260 47.270 77.580 47.300 ;
        RECT 76.020 47.240 76.210 47.250 ;
        RECT 76.020 46.950 76.220 47.240 ;
        RECT 77.260 47.080 77.590 47.270 ;
        RECT 82.710 47.210 83.460 47.440 ;
        RECT 80.740 47.170 80.910 47.200 ;
        RECT 81.150 47.170 81.350 47.210 ;
        RECT 77.260 47.040 77.580 47.080 ;
        RECT 76.010 46.620 76.300 46.950 ;
        RECT 80.740 46.910 81.350 47.170 ;
        RECT 80.740 46.870 80.910 46.910 ;
        RECT 81.150 46.880 81.350 46.910 ;
        RECT 81.150 46.520 81.350 46.550 ;
        RECT 80.920 46.260 81.350 46.520 ;
        RECT 75.650 45.950 75.830 46.140 ;
        RECT 68.260 45.550 72.040 45.730 ;
        RECT 45.660 44.880 46.110 45.030 ;
        RECT 65.890 44.840 66.440 45.270 ;
        RECT 68.260 45.130 68.680 45.550 ;
        RECT 69.520 43.820 69.750 44.550 ;
        RECT 74.820 44.460 74.990 45.320 ;
        RECT 74.660 44.200 74.990 44.460 ;
        RECT 74.820 43.630 74.990 44.200 ;
        RECT 75.650 45.230 75.830 45.420 ;
        RECT 75.650 43.620 75.820 45.230 ;
        RECT 77.380 45.170 77.560 46.230 ;
        RECT 81.150 46.220 81.350 46.260 ;
        RECT 81.740 46.220 82.290 47.210 ;
        RECT 82.760 46.790 83.460 47.210 ;
        RECT 108.580 47.030 108.790 47.460 ;
        RECT 83.220 46.430 83.540 46.470 ;
        RECT 83.220 46.370 83.550 46.430 ;
        RECT 111.900 46.420 112.080 47.900 ;
        RECT 112.710 47.800 112.930 47.900 ;
        RECT 114.000 47.850 114.630 48.020 ;
        RECT 112.150 47.590 112.500 47.760 ;
        RECT 112.680 47.720 112.930 47.800 ;
        RECT 112.600 47.600 112.930 47.720 ;
        RECT 112.600 47.490 112.880 47.600 ;
        RECT 112.710 46.430 112.880 47.490 ;
        RECT 82.750 46.240 83.550 46.370 ;
        RECT 82.750 46.210 83.540 46.240 ;
        RECT 82.750 46.190 83.450 46.210 ;
        RECT 77.990 45.990 78.310 46.020 ;
        RECT 77.990 45.800 78.320 45.990 ;
        RECT 77.990 45.760 78.310 45.800 ;
        RECT 77.990 45.680 78.160 45.760 ;
        RECT 83.210 45.710 83.530 45.750 ;
        RECT 77.940 45.510 78.160 45.680 ;
        RECT 81.150 45.670 81.350 45.710 ;
        RECT 77.940 45.350 78.110 45.510 ;
        RECT 80.920 45.410 81.350 45.670 ;
        RECT 81.150 45.380 81.350 45.410 ;
        RECT 78.430 45.010 78.510 45.090 ;
        RECT 78.570 45.010 78.760 45.130 ;
        RECT 78.430 44.920 78.760 45.010 ;
        RECT 78.570 44.900 78.760 44.920 ;
        RECT 80.740 45.020 80.910 45.060 ;
        RECT 81.150 45.020 81.350 45.050 ;
        RECT 80.740 44.760 81.350 45.020 ;
        RECT 76.010 44.420 76.300 44.750 ;
        RECT 80.740 44.730 80.910 44.760 ;
        RECT 81.150 44.720 81.350 44.760 ;
        RECT 81.740 44.720 82.290 45.710 ;
        RECT 82.750 45.530 83.540 45.710 ;
        RECT 83.210 45.520 83.540 45.530 ;
        RECT 83.210 45.490 83.530 45.520 ;
        RECT 82.760 44.850 83.460 45.110 ;
        RECT 82.710 44.620 83.460 44.850 ;
        RECT 76.020 44.130 76.220 44.420 ;
        RECT 82.760 44.230 83.460 44.620 ;
        RECT 80.740 44.170 80.910 44.200 ;
        RECT 81.150 44.170 81.350 44.210 ;
        RECT 76.020 44.120 76.210 44.130 ;
        RECT 76.380 43.950 76.590 43.960 ;
        RECT 76.370 43.370 76.590 43.950 ;
        RECT 80.740 43.910 81.350 44.170 ;
        RECT 80.740 43.870 80.910 43.910 ;
        RECT 81.150 43.880 81.350 43.910 ;
        RECT 81.010 43.550 81.190 43.790 ;
        RECT 81.010 43.520 81.350 43.550 ;
        RECT 76.380 43.340 76.590 43.370 ;
        RECT 74.570 43.070 75.100 43.240 ;
        RECT 76.380 42.990 76.580 43.340 ;
        RECT 80.920 43.260 81.350 43.520 ;
        RECT 81.010 43.220 81.350 43.260 ;
        RECT 81.740 43.220 82.290 44.210 ;
        RECT 82.760 43.620 83.470 43.790 ;
        RECT 83.110 43.340 83.470 43.620 ;
        RECT 111.900 43.370 112.080 45.420 ;
        RECT 112.630 45.160 112.960 45.330 ;
        RECT 112.710 43.380 112.880 45.160 ;
        RECT 81.010 41.740 81.190 43.220 ;
        RECT 81.820 41.750 81.990 43.220 ;
        RECT 83.110 43.170 83.740 43.340 ;
        RECT 38.910 41.160 39.080 41.210 ;
        RECT 38.880 40.940 39.100 41.160 ;
        RECT 38.910 40.880 39.080 40.940 ;
        RECT 39.430 40.800 39.760 40.980 ;
        RECT 42.570 40.970 42.740 41.020 ;
        RECT 40.010 40.800 42.170 40.970 ;
        RECT 42.410 40.800 42.740 40.970 ;
        RECT 43.030 40.830 43.240 41.160 ;
        RECT 39.460 40.360 39.730 40.800 ;
        RECT 40.940 40.540 41.270 40.800 ;
        RECT 42.480 40.660 42.740 40.800 ;
        RECT 43.480 40.660 43.660 41.100 ;
        RECT 45.080 41.000 45.470 41.050 ;
        RECT 44.210 40.940 45.470 41.000 ;
        RECT 44.210 40.830 45.550 40.940 ;
        RECT 45.080 40.770 45.550 40.830 ;
        RECT 46.020 40.790 46.980 40.960 ;
        RECT 45.080 40.760 45.460 40.770 ;
        RECT 39.500 40.350 39.730 40.360 ;
        RECT 42.480 40.490 43.660 40.660 ;
        RECT 42.480 40.350 42.740 40.490 ;
        RECT 39.500 40.180 40.260 40.350 ;
        RECT 40.510 40.180 41.680 40.350 ;
        RECT 41.920 40.320 42.740 40.350 ;
        RECT 41.920 40.180 43.030 40.320 ;
        RECT 40.910 40.080 41.260 40.180 ;
        RECT 42.570 40.150 43.030 40.180 ;
        RECT 43.480 40.310 44.670 40.320 ;
        RECT 43.480 40.150 44.960 40.310 ;
        RECT 43.520 40.130 44.960 40.150 ;
        RECT 44.500 40.090 44.960 40.130 ;
        RECT 44.670 40.070 44.960 40.090 ;
        RECT 45.290 40.000 45.460 40.760 ;
        RECT 46.800 40.330 46.980 40.790 ;
        RECT 47.950 40.440 48.120 40.860 ;
        RECT 48.760 40.740 49.000 40.770 ;
        RECT 48.430 40.570 49.000 40.740 ;
        RECT 49.240 40.570 50.580 40.740 ;
        RECT 51.030 40.570 51.990 40.740 ;
        RECT 48.760 40.530 49.000 40.570 ;
        RECT 51.540 40.560 51.710 40.570 ;
        RECT 45.660 40.150 46.260 40.320 ;
        RECT 46.720 40.160 47.050 40.330 ;
        RECT 47.880 40.220 48.050 40.260 ;
        RECT 45.660 40.000 46.110 40.150 ;
        RECT 47.820 40.050 48.050 40.220 ;
        RECT 51.170 40.120 51.510 40.300 ;
        RECT 47.880 39.700 48.050 40.050 ;
        RECT 48.120 39.830 48.310 40.060 ;
        RECT 48.410 39.950 48.780 40.120 ;
        RECT 49.240 39.950 51.990 40.120 ;
        RECT 52.520 39.880 52.690 40.810 ;
        RECT 52.920 39.970 53.090 40.860 ;
        RECT 55.830 40.450 56.030 40.800 ;
        RECT 57.570 40.720 57.890 40.730 ;
        RECT 57.310 40.550 57.890 40.720 ;
        RECT 57.560 40.500 57.890 40.550 ;
        RECT 57.570 40.470 57.890 40.500 ;
        RECT 73.090 40.720 73.410 40.730 ;
        RECT 73.090 40.550 73.670 40.720 ;
        RECT 73.090 40.500 73.420 40.550 ;
        RECT 73.090 40.470 73.410 40.500 ;
        RECT 55.820 40.420 56.030 40.450 ;
        RECT 74.950 40.450 75.150 40.800 ;
        RECT 55.820 39.830 56.040 40.420 ;
        RECT 56.560 39.830 56.760 40.430 ;
        RECT 57.570 40.140 57.890 40.180 ;
        RECT 57.560 40.100 57.890 40.140 ;
        RECT 57.310 39.930 57.890 40.100 ;
        RECT 57.570 39.920 57.890 39.930 ;
        RECT 73.090 40.140 73.410 40.180 ;
        RECT 73.090 40.100 73.420 40.140 ;
        RECT 73.090 39.930 73.670 40.100 ;
        RECT 73.090 39.920 73.410 39.930 ;
        RECT 74.220 39.830 74.420 40.430 ;
        RECT 74.950 40.420 75.160 40.450 ;
        RECT 74.940 39.830 75.160 40.420 ;
        RECT 38.910 39.410 39.080 39.460 ;
        RECT 38.880 39.190 39.100 39.410 ;
        RECT 38.910 39.130 39.080 39.190 ;
        RECT 39.430 39.050 39.760 39.230 ;
        RECT 42.570 39.220 42.740 39.270 ;
        RECT 40.010 39.050 42.170 39.220 ;
        RECT 42.410 39.050 42.740 39.220 ;
        RECT 43.030 39.080 43.240 39.410 ;
        RECT 39.460 38.610 39.730 39.050 ;
        RECT 40.940 38.790 41.270 39.050 ;
        RECT 42.480 38.910 42.740 39.050 ;
        RECT 43.480 38.910 43.660 39.350 ;
        RECT 45.080 39.250 45.470 39.300 ;
        RECT 44.210 39.190 45.470 39.250 ;
        RECT 44.210 39.080 45.550 39.190 ;
        RECT 45.080 39.020 45.550 39.080 ;
        RECT 46.020 39.040 46.980 39.210 ;
        RECT 45.080 39.010 45.460 39.020 ;
        RECT 39.500 38.600 39.730 38.610 ;
        RECT 42.480 38.740 43.660 38.910 ;
        RECT 42.480 38.600 42.740 38.740 ;
        RECT 39.500 38.430 40.260 38.600 ;
        RECT 40.510 38.430 41.680 38.600 ;
        RECT 41.920 38.570 42.740 38.600 ;
        RECT 41.920 38.430 43.030 38.570 ;
        RECT 40.910 38.330 41.260 38.430 ;
        RECT 42.570 38.400 43.030 38.430 ;
        RECT 43.480 38.560 44.670 38.570 ;
        RECT 43.480 38.400 44.960 38.560 ;
        RECT 43.520 38.380 44.960 38.400 ;
        RECT 44.500 38.340 44.960 38.380 ;
        RECT 44.670 38.320 44.960 38.340 ;
        RECT 45.290 38.250 45.460 39.010 ;
        RECT 46.800 38.580 46.980 39.040 ;
        RECT 47.880 38.940 48.050 39.290 ;
        RECT 47.820 38.770 48.050 38.940 ;
        RECT 48.120 38.930 48.310 39.160 ;
        RECT 48.410 38.870 48.780 39.040 ;
        RECT 49.240 38.870 51.990 39.040 ;
        RECT 47.880 38.730 48.050 38.770 ;
        RECT 51.170 38.690 51.510 38.870 ;
        RECT 45.660 38.400 46.260 38.570 ;
        RECT 46.720 38.410 47.050 38.580 ;
        RECT 45.660 38.250 46.110 38.400 ;
        RECT 47.950 38.130 48.120 38.550 ;
        RECT 48.760 38.420 49.000 38.460 ;
        RECT 51.540 38.420 51.710 38.430 ;
        RECT 48.430 38.250 49.000 38.420 ;
        RECT 49.240 38.250 50.580 38.420 ;
        RECT 51.030 38.250 51.990 38.420 ;
        RECT 48.760 38.220 49.000 38.250 ;
        RECT 52.520 38.180 52.690 39.110 ;
        RECT 52.920 38.130 53.090 39.020 ;
        RECT 55.820 38.690 56.040 39.280 ;
        RECT 55.820 38.660 56.030 38.690 ;
        RECT 56.560 38.680 56.760 39.280 ;
        RECT 58.570 39.200 58.740 39.730 ;
        RECT 62.510 39.210 62.680 39.740 ;
        RECT 68.300 39.210 68.470 39.740 ;
        RECT 72.240 39.200 72.410 39.730 ;
        RECT 57.570 39.180 57.890 39.190 ;
        RECT 57.310 39.010 57.890 39.180 ;
        RECT 57.560 38.970 57.890 39.010 ;
        RECT 57.570 38.930 57.890 38.970 ;
        RECT 73.090 39.180 73.410 39.190 ;
        RECT 73.090 39.010 73.670 39.180 ;
        RECT 73.090 38.970 73.420 39.010 ;
        RECT 73.090 38.930 73.410 38.970 ;
        RECT 74.220 38.680 74.420 39.280 ;
        RECT 74.940 38.690 75.160 39.280 ;
        RECT 81.010 38.690 81.190 40.740 ;
        RECT 81.740 40.480 82.070 40.650 ;
        RECT 81.820 38.700 81.990 40.480 ;
        RECT 55.830 38.310 56.030 38.660 ;
        RECT 74.950 38.660 75.160 38.690 ;
        RECT 57.570 38.610 57.890 38.640 ;
        RECT 57.560 38.560 57.890 38.610 ;
        RECT 57.310 38.390 57.890 38.560 ;
        RECT 73.090 38.610 73.410 38.640 ;
        RECT 73.090 38.560 73.420 38.610 ;
        RECT 57.570 38.380 57.890 38.390 ;
        RECT 56.200 37.850 56.640 38.020 ;
        RECT 38.910 37.660 39.080 37.710 ;
        RECT 38.880 37.440 39.100 37.660 ;
        RECT 38.910 37.380 39.080 37.440 ;
        RECT 39.430 37.300 39.760 37.480 ;
        RECT 42.570 37.470 42.740 37.520 ;
        RECT 40.010 37.300 42.170 37.470 ;
        RECT 42.410 37.300 42.740 37.470 ;
        RECT 43.030 37.330 43.240 37.660 ;
        RECT 39.460 36.860 39.730 37.300 ;
        RECT 40.940 37.040 41.270 37.300 ;
        RECT 42.480 37.160 42.740 37.300 ;
        RECT 43.480 37.160 43.660 37.600 ;
        RECT 45.080 37.500 45.470 37.550 ;
        RECT 44.210 37.440 45.470 37.500 ;
        RECT 44.210 37.330 45.550 37.440 ;
        RECT 45.080 37.270 45.550 37.330 ;
        RECT 46.020 37.290 46.980 37.460 ;
        RECT 45.080 37.260 45.460 37.270 ;
        RECT 39.500 36.850 39.730 36.860 ;
        RECT 42.480 36.990 43.660 37.160 ;
        RECT 42.480 36.850 42.740 36.990 ;
        RECT 39.500 36.680 40.260 36.850 ;
        RECT 40.510 36.680 41.680 36.850 ;
        RECT 41.920 36.820 42.740 36.850 ;
        RECT 41.920 36.680 43.030 36.820 ;
        RECT 40.910 36.580 41.260 36.680 ;
        RECT 42.570 36.650 43.030 36.680 ;
        RECT 43.480 36.810 44.670 36.820 ;
        RECT 43.480 36.650 44.960 36.810 ;
        RECT 43.520 36.630 44.960 36.650 ;
        RECT 44.500 36.590 44.960 36.630 ;
        RECT 44.670 36.570 44.960 36.590 ;
        RECT 45.290 36.500 45.460 37.260 ;
        RECT 46.800 36.830 46.980 37.290 ;
        RECT 47.950 37.240 48.120 37.660 ;
        RECT 48.760 37.540 49.000 37.570 ;
        RECT 48.430 37.370 49.000 37.540 ;
        RECT 49.240 37.370 50.580 37.540 ;
        RECT 51.030 37.370 51.990 37.540 ;
        RECT 48.760 37.330 49.000 37.370 ;
        RECT 51.540 37.360 51.710 37.370 ;
        RECT 47.880 37.020 48.050 37.060 ;
        RECT 47.820 36.850 48.050 37.020 ;
        RECT 51.170 36.920 51.510 37.100 ;
        RECT 45.660 36.650 46.260 36.820 ;
        RECT 46.720 36.660 47.050 36.830 ;
        RECT 45.660 36.500 46.110 36.650 ;
        RECT 47.880 36.500 48.050 36.850 ;
        RECT 48.120 36.630 48.310 36.860 ;
        RECT 48.410 36.750 48.780 36.920 ;
        RECT 49.240 36.750 51.990 36.920 ;
        RECT 52.520 36.680 52.690 37.610 ;
        RECT 52.920 36.770 53.090 37.660 ;
        RECT 55.830 37.210 56.030 37.560 ;
        RECT 57.570 37.480 57.890 37.490 ;
        RECT 57.310 37.310 57.890 37.480 ;
        RECT 58.570 37.360 58.740 38.370 ;
        RECT 60.500 37.640 61.050 38.070 ;
        RECT 62.500 37.500 62.670 38.510 ;
        RECT 64.530 37.710 65.080 38.140 ;
        RECT 65.900 37.710 66.450 38.140 ;
        RECT 68.310 37.500 68.480 38.510 ;
        RECT 73.090 38.390 73.670 38.560 ;
        RECT 73.090 38.380 73.410 38.390 ;
        RECT 69.930 37.640 70.480 38.070 ;
        RECT 72.240 37.360 72.410 38.370 ;
        RECT 74.950 38.310 75.150 38.660 ;
        RECT 74.340 37.850 74.780 38.020 ;
        RECT 73.090 37.480 73.410 37.490 ;
        RECT 57.560 37.260 57.890 37.310 ;
        RECT 57.570 37.230 57.890 37.260 ;
        RECT 73.090 37.310 73.670 37.480 ;
        RECT 73.090 37.260 73.420 37.310 ;
        RECT 73.090 37.230 73.410 37.260 ;
        RECT 55.820 37.180 56.030 37.210 ;
        RECT 74.950 37.210 75.150 37.560 ;
        RECT 55.820 36.590 56.040 37.180 ;
        RECT 56.560 36.590 56.760 37.190 ;
        RECT 57.570 36.900 57.890 36.940 ;
        RECT 57.560 36.860 57.890 36.900 ;
        RECT 57.310 36.690 57.890 36.860 ;
        RECT 57.570 36.680 57.890 36.690 ;
        RECT 73.090 36.900 73.410 36.940 ;
        RECT 73.090 36.860 73.420 36.900 ;
        RECT 73.090 36.690 73.670 36.860 ;
        RECT 73.090 36.680 73.410 36.690 ;
        RECT 74.220 36.590 74.420 37.190 ;
        RECT 74.950 37.180 75.160 37.210 ;
        RECT 74.940 36.590 75.160 37.180 ;
        RECT 38.910 35.910 39.080 35.960 ;
        RECT 38.880 35.690 39.100 35.910 ;
        RECT 38.910 35.630 39.080 35.690 ;
        RECT 39.430 35.550 39.760 35.730 ;
        RECT 42.570 35.720 42.740 35.770 ;
        RECT 40.010 35.550 42.170 35.720 ;
        RECT 42.410 35.550 42.740 35.720 ;
        RECT 43.030 35.580 43.240 35.910 ;
        RECT 39.460 35.110 39.730 35.550 ;
        RECT 40.940 35.290 41.270 35.550 ;
        RECT 42.480 35.410 42.740 35.550 ;
        RECT 43.480 35.410 43.660 35.850 ;
        RECT 45.080 35.750 45.470 35.800 ;
        RECT 44.210 35.690 45.470 35.750 ;
        RECT 47.880 35.740 48.050 36.090 ;
        RECT 44.210 35.580 45.550 35.690 ;
        RECT 45.080 35.520 45.550 35.580 ;
        RECT 46.020 35.540 46.980 35.710 ;
        RECT 47.820 35.570 48.050 35.740 ;
        RECT 48.120 35.730 48.310 35.960 ;
        RECT 48.410 35.670 48.780 35.840 ;
        RECT 49.240 35.670 51.990 35.840 ;
        RECT 45.080 35.510 45.460 35.520 ;
        RECT 39.500 35.100 39.730 35.110 ;
        RECT 42.480 35.240 43.660 35.410 ;
        RECT 42.480 35.100 42.740 35.240 ;
        RECT 39.500 34.930 40.260 35.100 ;
        RECT 40.510 34.930 41.680 35.100 ;
        RECT 41.920 35.070 42.740 35.100 ;
        RECT 41.920 34.930 43.030 35.070 ;
        RECT 40.910 34.830 41.260 34.930 ;
        RECT 42.570 34.900 43.030 34.930 ;
        RECT 43.480 35.060 44.670 35.070 ;
        RECT 43.480 34.900 44.960 35.060 ;
        RECT 43.520 34.880 44.960 34.900 ;
        RECT 44.500 34.840 44.960 34.880 ;
        RECT 44.670 34.820 44.960 34.840 ;
        RECT 45.290 34.750 45.460 35.510 ;
        RECT 46.800 35.080 46.980 35.540 ;
        RECT 47.880 35.530 48.050 35.570 ;
        RECT 51.170 35.490 51.510 35.670 ;
        RECT 45.660 34.900 46.260 35.070 ;
        RECT 46.720 34.910 47.050 35.080 ;
        RECT 47.950 34.930 48.120 35.350 ;
        RECT 48.760 35.220 49.000 35.260 ;
        RECT 51.540 35.220 51.710 35.230 ;
        RECT 48.430 35.050 49.000 35.220 ;
        RECT 49.240 35.050 50.580 35.220 ;
        RECT 51.030 35.050 51.990 35.220 ;
        RECT 48.760 35.020 49.000 35.050 ;
        RECT 52.520 34.980 52.690 35.910 ;
        RECT 52.920 34.930 53.090 35.820 ;
        RECT 53.220 35.120 53.420 35.470 ;
        RECT 55.820 35.460 56.040 36.050 ;
        RECT 55.820 35.430 56.030 35.460 ;
        RECT 56.560 35.450 56.760 36.050 ;
        RECT 57.570 35.950 57.890 35.960 ;
        RECT 57.310 35.780 57.890 35.950 ;
        RECT 57.560 35.740 57.890 35.780 ;
        RECT 57.570 35.700 57.890 35.740 ;
        RECT 73.090 35.950 73.410 35.960 ;
        RECT 73.090 35.780 73.670 35.950 ;
        RECT 73.090 35.740 73.420 35.780 ;
        RECT 73.090 35.700 73.410 35.740 ;
        RECT 74.220 35.450 74.420 36.050 ;
        RECT 74.940 35.460 75.160 36.050 ;
        RECT 54.960 35.390 55.280 35.400 ;
        RECT 54.700 35.220 55.280 35.390 ;
        RECT 54.950 35.170 55.280 35.220 ;
        RECT 54.960 35.140 55.280 35.170 ;
        RECT 53.210 35.090 53.420 35.120 ;
        RECT 45.660 34.750 46.110 34.900 ;
        RECT 53.210 34.500 53.430 35.090 ;
        RECT 53.950 34.500 54.150 35.100 ;
        RECT 55.830 35.080 56.030 35.430 ;
        RECT 74.950 35.430 75.160 35.460 ;
        RECT 57.570 35.380 57.890 35.410 ;
        RECT 57.560 35.330 57.890 35.380 ;
        RECT 57.310 35.160 57.890 35.330 ;
        RECT 57.570 35.150 57.890 35.160 ;
        RECT 73.090 35.380 73.410 35.410 ;
        RECT 73.090 35.330 73.420 35.380 ;
        RECT 73.090 35.160 73.670 35.330 ;
        RECT 73.090 35.150 73.410 35.160 ;
        RECT 74.950 35.080 75.150 35.430 ;
        RECT 54.960 34.810 55.280 34.850 ;
        RECT 54.950 34.770 55.280 34.810 ;
        RECT 54.700 34.600 55.280 34.770 ;
        RECT 54.960 34.590 55.280 34.600 ;
        RECT 53.210 33.380 53.430 33.970 ;
        RECT 53.210 33.350 53.420 33.380 ;
        RECT 53.950 33.370 54.150 33.970 ;
        RECT 54.960 33.870 55.280 33.880 ;
        RECT 54.700 33.700 55.280 33.870 ;
        RECT 56.090 33.810 56.260 34.340 ;
        RECT 60.110 33.840 60.280 34.370 ;
        RECT 54.950 33.660 55.280 33.700 ;
        RECT 54.960 33.620 55.280 33.660 ;
        RECT 53.220 33.000 53.420 33.350 ;
        RECT 54.960 33.300 55.280 33.330 ;
        RECT 54.950 33.250 55.280 33.300 ;
        RECT 54.700 33.080 55.280 33.250 ;
        RECT 54.960 33.070 55.280 33.080 ;
        RECT 53.590 32.540 54.030 32.710 ;
        RECT 38.870 32.100 39.040 32.150 ;
        RECT 38.840 31.880 39.060 32.100 ;
        RECT 38.870 31.820 39.040 31.880 ;
        RECT 39.390 31.740 39.720 31.920 ;
        RECT 42.530 31.910 42.700 31.960 ;
        RECT 39.970 31.740 42.130 31.910 ;
        RECT 42.370 31.740 42.700 31.910 ;
        RECT 42.990 31.770 43.200 32.100 ;
        RECT 39.420 31.300 39.690 31.740 ;
        RECT 40.900 31.480 41.230 31.740 ;
        RECT 42.440 31.600 42.700 31.740 ;
        RECT 43.440 31.600 43.620 32.040 ;
        RECT 45.040 31.940 45.430 31.990 ;
        RECT 44.170 31.880 45.430 31.940 ;
        RECT 44.170 31.770 45.510 31.880 ;
        RECT 45.040 31.710 45.510 31.770 ;
        RECT 45.980 31.730 46.940 31.900 ;
        RECT 53.220 31.880 53.420 32.230 ;
        RECT 54.960 32.150 55.280 32.160 ;
        RECT 54.700 31.980 55.280 32.150 ;
        RECT 54.950 31.930 55.280 31.980 ;
        RECT 56.080 31.950 56.250 33.140 ;
        RECT 57.890 32.270 58.440 32.700 ;
        RECT 54.960 31.900 55.280 31.930 ;
        RECT 60.100 31.910 60.270 33.080 ;
        RECT 61.920 32.340 62.470 32.770 ;
        RECT 45.040 31.700 45.420 31.710 ;
        RECT 39.460 31.290 39.690 31.300 ;
        RECT 42.440 31.430 43.620 31.600 ;
        RECT 42.440 31.290 42.700 31.430 ;
        RECT 39.460 31.120 40.220 31.290 ;
        RECT 40.470 31.120 41.640 31.290 ;
        RECT 41.880 31.260 42.700 31.290 ;
        RECT 41.880 31.120 42.990 31.260 ;
        RECT 40.870 31.020 41.220 31.120 ;
        RECT 42.530 31.090 42.990 31.120 ;
        RECT 43.440 31.250 44.630 31.260 ;
        RECT 43.440 31.090 44.920 31.250 ;
        RECT 43.480 31.070 44.920 31.090 ;
        RECT 44.460 31.030 44.920 31.070 ;
        RECT 44.630 31.010 44.920 31.030 ;
        RECT 45.250 30.940 45.420 31.700 ;
        RECT 46.760 31.270 46.940 31.730 ;
        RECT 53.210 31.850 53.420 31.880 ;
        RECT 45.620 31.090 46.220 31.260 ;
        RECT 46.680 31.100 47.010 31.270 ;
        RECT 47.980 31.170 48.150 31.590 ;
        RECT 48.790 31.470 49.030 31.500 ;
        RECT 48.460 31.300 49.030 31.470 ;
        RECT 49.270 31.300 50.610 31.470 ;
        RECT 51.060 31.300 52.020 31.470 ;
        RECT 48.790 31.260 49.030 31.300 ;
        RECT 51.570 31.290 51.740 31.300 ;
        RECT 45.620 30.940 46.070 31.090 ;
        RECT 47.910 30.950 48.080 30.990 ;
        RECT 19.380 30.370 19.550 30.860 ;
        RECT 19.230 30.340 19.550 30.370 ;
        RECT 19.930 30.370 20.100 30.860 ;
        RECT 20.570 30.810 20.740 30.860 ;
        RECT 21.120 30.810 21.290 30.860 ;
        RECT 20.450 30.780 20.770 30.810 ;
        RECT 21.100 30.780 21.420 30.810 ;
        RECT 47.850 30.780 48.080 30.950 ;
        RECT 51.200 30.850 51.540 31.030 ;
        RECT 20.450 30.590 20.780 30.780 ;
        RECT 21.100 30.590 21.430 30.780 ;
        RECT 20.450 30.550 20.770 30.590 ;
        RECT 21.100 30.550 21.420 30.590 ;
        RECT 19.930 30.340 20.250 30.370 ;
        RECT 19.230 30.150 19.560 30.340 ;
        RECT 19.930 30.150 20.260 30.340 ;
        RECT 19.230 30.110 19.550 30.150 ;
        RECT 19.380 28.460 19.550 30.110 ;
        RECT 19.930 30.110 20.250 30.150 ;
        RECT 19.930 28.460 20.100 30.110 ;
        RECT 20.570 28.460 20.740 30.550 ;
        RECT 21.120 28.460 21.290 30.550 ;
        RECT 47.910 30.430 48.080 30.780 ;
        RECT 48.150 30.560 48.340 30.790 ;
        RECT 48.440 30.680 48.810 30.850 ;
        RECT 49.270 30.680 52.020 30.850 ;
        RECT 52.550 30.610 52.720 31.540 ;
        RECT 52.950 30.700 53.120 31.590 ;
        RECT 53.210 31.260 53.430 31.850 ;
        RECT 53.950 31.260 54.150 31.860 ;
        RECT 54.960 31.570 55.280 31.610 ;
        RECT 54.950 31.530 55.280 31.570 ;
        RECT 54.700 31.360 55.280 31.530 ;
        RECT 54.960 31.350 55.280 31.360 ;
        RECT 66.310 31.070 66.630 31.100 ;
        RECT 66.310 30.900 68.100 31.070 ;
        RECT 66.310 30.880 66.640 30.900 ;
        RECT 66.310 30.840 66.630 30.880 ;
        RECT 38.870 30.350 39.040 30.400 ;
        RECT 38.840 30.130 39.060 30.350 ;
        RECT 38.870 30.070 39.040 30.130 ;
        RECT 39.390 29.990 39.720 30.170 ;
        RECT 42.530 30.160 42.700 30.210 ;
        RECT 39.970 29.990 42.130 30.160 ;
        RECT 42.370 29.990 42.700 30.160 ;
        RECT 42.990 30.020 43.200 30.350 ;
        RECT 21.670 29.100 21.840 29.950 ;
        RECT 39.420 29.550 39.690 29.990 ;
        RECT 40.900 29.730 41.230 29.990 ;
        RECT 42.440 29.850 42.700 29.990 ;
        RECT 43.440 29.850 43.620 30.290 ;
        RECT 45.040 30.190 45.430 30.240 ;
        RECT 44.170 30.130 45.430 30.190 ;
        RECT 44.170 30.020 45.510 30.130 ;
        RECT 45.040 29.960 45.510 30.020 ;
        RECT 45.980 29.980 46.940 30.150 ;
        RECT 53.210 30.130 53.430 30.720 ;
        RECT 53.210 30.100 53.420 30.130 ;
        RECT 53.950 30.120 54.150 30.720 ;
        RECT 67.930 30.670 68.100 30.900 ;
        RECT 54.960 30.620 55.280 30.630 ;
        RECT 54.700 30.450 55.280 30.620 ;
        RECT 54.950 30.410 55.280 30.450 ;
        RECT 66.780 30.420 67.120 30.670 ;
        RECT 67.290 30.500 67.620 30.670 ;
        RECT 67.840 30.500 68.180 30.670 ;
        RECT 54.960 30.370 55.280 30.410 ;
        RECT 66.460 30.160 67.120 30.420 ;
        RECT 67.370 30.330 67.540 30.500 ;
        RECT 67.930 30.330 68.100 30.500 ;
        RECT 67.290 30.160 67.620 30.330 ;
        RECT 67.840 30.160 68.180 30.330 ;
        RECT 45.040 29.950 45.420 29.960 ;
        RECT 39.460 29.540 39.690 29.550 ;
        RECT 42.440 29.680 43.620 29.850 ;
        RECT 42.440 29.540 42.700 29.680 ;
        RECT 39.460 29.370 40.220 29.540 ;
        RECT 40.470 29.370 41.640 29.540 ;
        RECT 41.880 29.510 42.700 29.540 ;
        RECT 41.880 29.370 42.990 29.510 ;
        RECT 40.870 29.270 41.220 29.370 ;
        RECT 42.530 29.340 42.990 29.370 ;
        RECT 43.440 29.500 44.630 29.510 ;
        RECT 43.440 29.340 44.920 29.500 ;
        RECT 43.480 29.320 44.920 29.340 ;
        RECT 44.460 29.280 44.920 29.320 ;
        RECT 44.630 29.260 44.920 29.280 ;
        RECT 45.250 29.190 45.420 29.950 ;
        RECT 46.760 29.520 46.940 29.980 ;
        RECT 47.910 29.670 48.080 30.020 ;
        RECT 45.620 29.340 46.220 29.510 ;
        RECT 46.680 29.350 47.010 29.520 ;
        RECT 47.850 29.500 48.080 29.670 ;
        RECT 48.150 29.660 48.340 29.890 ;
        RECT 48.440 29.600 48.810 29.770 ;
        RECT 49.270 29.600 52.020 29.770 ;
        RECT 47.910 29.460 48.080 29.500 ;
        RECT 51.200 29.420 51.540 29.600 ;
        RECT 45.620 29.190 46.070 29.340 ;
        RECT 47.980 28.860 48.150 29.280 ;
        RECT 48.790 29.150 49.030 29.190 ;
        RECT 51.570 29.150 51.740 29.160 ;
        RECT 48.460 28.980 49.030 29.150 ;
        RECT 49.270 28.980 50.610 29.150 ;
        RECT 51.060 28.980 52.020 29.150 ;
        RECT 48.790 28.950 49.030 28.980 ;
        RECT 52.550 28.910 52.720 29.840 ;
        RECT 53.220 29.750 53.420 30.100 ;
        RECT 54.960 30.050 55.280 30.080 ;
        RECT 54.950 30.000 55.280 30.050 ;
        RECT 54.700 29.830 55.280 30.000 ;
        RECT 54.960 29.820 55.280 29.830 ;
        RECT 67.370 29.930 67.620 30.160 ;
        RECT 68.500 30.080 69.010 30.750 ;
        RECT 67.370 29.760 68.040 29.930 ;
        RECT 52.950 28.860 53.120 29.750 ;
        RECT 67.370 29.530 67.620 29.760 ;
        RECT 66.460 29.270 67.120 29.530 ;
        RECT 67.290 29.360 67.620 29.530 ;
        RECT 67.840 29.360 68.180 29.530 ;
        RECT 66.780 29.020 67.120 29.270 ;
        RECT 67.370 29.190 67.540 29.360 ;
        RECT 67.930 29.190 68.100 29.360 ;
        RECT 67.290 29.020 67.620 29.190 ;
        RECT 67.840 29.020 68.180 29.190 ;
        RECT 66.310 28.810 66.630 28.850 ;
        RECT 66.310 28.790 66.640 28.810 ;
        RECT 67.930 28.790 68.100 29.020 ;
        RECT 68.500 28.940 69.010 29.610 ;
        RECT 38.870 28.600 39.040 28.650 ;
        RECT 66.310 28.620 68.100 28.790 ;
        RECT 21.560 28.470 21.990 28.490 ;
        RECT 18.750 28.390 18.920 28.410 ;
        RECT 18.730 28.270 18.940 28.390 ;
        RECT 21.560 28.300 22.010 28.470 ;
        RECT 38.840 28.380 39.060 28.600 ;
        RECT 38.870 28.320 39.040 28.380 ;
        RECT 21.560 28.280 21.990 28.300 ;
        RECT 18.730 27.960 19.130 28.270 ;
        RECT 39.390 28.240 39.720 28.420 ;
        RECT 42.530 28.410 42.700 28.460 ;
        RECT 39.970 28.240 42.130 28.410 ;
        RECT 42.370 28.240 42.700 28.410 ;
        RECT 42.990 28.270 43.200 28.600 ;
        RECT 66.310 28.590 66.630 28.620 ;
        RECT 18.920 27.840 19.130 27.960 ;
        RECT 21.570 27.930 22.000 27.950 ;
        RECT 18.940 27.820 19.110 27.840 ;
        RECT 19.390 26.490 19.560 27.810 ;
        RECT 19.260 26.460 19.580 26.490 ;
        RECT 19.940 26.480 20.110 27.820 ;
        RECT 13.960 25.790 14.280 25.820 ;
        RECT 15.060 25.800 15.380 25.830 ;
        RECT 16.150 25.800 16.470 25.830 ;
        RECT 13.950 25.600 14.280 25.790 ;
        RECT 15.050 25.610 15.380 25.800 ;
        RECT 16.140 25.610 16.470 25.800 ;
        RECT 12.380 23.180 12.550 25.580 ;
        RECT 12.930 23.180 13.100 25.580 ;
        RECT 13.480 23.180 13.650 25.580 ;
        RECT 13.960 25.560 14.280 25.600 ;
        RECT 14.030 23.110 14.200 25.560 ;
        RECT 14.580 25.150 14.750 25.580 ;
        RECT 15.060 25.570 15.380 25.610 ;
        RECT 16.150 25.570 16.470 25.610 ;
        RECT 17.190 25.610 17.700 26.290 ;
        RECT 19.260 26.270 19.590 26.460 ;
        RECT 19.940 26.450 20.270 26.480 ;
        RECT 19.260 26.230 19.580 26.270 ;
        RECT 19.940 26.260 20.280 26.450 ;
        RECT 14.510 25.120 14.830 25.150 ;
        RECT 14.500 24.930 14.830 25.120 ;
        RECT 14.510 24.890 14.830 24.930 ;
        RECT 14.580 23.780 14.750 24.890 ;
        RECT 14.510 23.750 14.830 23.780 ;
        RECT 14.500 23.560 14.830 23.750 ;
        RECT 14.510 23.520 14.830 23.560 ;
        RECT 14.580 23.110 14.750 23.520 ;
        RECT 15.130 23.110 15.300 25.570 ;
        RECT 17.190 25.540 17.710 25.610 ;
        RECT 17.200 25.280 17.710 25.540 ;
        RECT 19.390 25.320 19.560 26.230 ;
        RECT 19.940 26.220 20.270 26.260 ;
        RECT 19.940 25.320 20.110 26.220 ;
        RECT 20.570 25.710 20.740 27.810 ;
        RECT 20.430 25.680 20.750 25.710 ;
        RECT 20.430 25.490 20.760 25.680 ;
        RECT 21.120 25.650 21.290 27.820 ;
        RECT 21.570 27.760 22.020 27.930 ;
        RECT 39.420 27.800 39.690 28.240 ;
        RECT 40.900 27.980 41.230 28.240 ;
        RECT 42.440 28.100 42.700 28.240 ;
        RECT 43.440 28.100 43.620 28.540 ;
        RECT 45.040 28.440 45.430 28.490 ;
        RECT 44.170 28.380 45.430 28.440 ;
        RECT 44.170 28.270 45.510 28.380 ;
        RECT 45.040 28.210 45.510 28.270 ;
        RECT 45.980 28.230 46.940 28.400 ;
        RECT 45.040 28.200 45.420 28.210 ;
        RECT 39.460 27.790 39.690 27.800 ;
        RECT 42.440 27.930 43.620 28.100 ;
        RECT 42.440 27.790 42.700 27.930 ;
        RECT 21.570 27.740 22.000 27.760 ;
        RECT 39.460 27.620 40.220 27.790 ;
        RECT 40.470 27.620 41.640 27.790 ;
        RECT 41.880 27.760 42.700 27.790 ;
        RECT 41.880 27.620 42.990 27.760 ;
        RECT 40.870 27.520 41.220 27.620 ;
        RECT 42.530 27.590 42.990 27.620 ;
        RECT 43.440 27.750 44.630 27.760 ;
        RECT 43.440 27.590 44.920 27.750 ;
        RECT 43.480 27.570 44.920 27.590 ;
        RECT 44.460 27.530 44.920 27.570 ;
        RECT 44.630 27.510 44.920 27.530 ;
        RECT 45.250 27.440 45.420 28.200 ;
        RECT 46.760 27.770 46.940 28.230 ;
        RECT 47.980 27.970 48.150 28.390 ;
        RECT 48.790 28.270 49.030 28.300 ;
        RECT 48.460 28.100 49.030 28.270 ;
        RECT 49.270 28.100 50.610 28.270 ;
        RECT 51.060 28.100 52.020 28.270 ;
        RECT 48.790 28.060 49.030 28.100 ;
        RECT 51.570 28.090 51.740 28.100 ;
        RECT 45.620 27.590 46.220 27.760 ;
        RECT 46.680 27.600 47.010 27.770 ;
        RECT 47.910 27.750 48.080 27.790 ;
        RECT 45.620 27.440 46.070 27.590 ;
        RECT 47.850 27.580 48.080 27.750 ;
        RECT 51.200 27.650 51.540 27.830 ;
        RECT 47.910 27.230 48.080 27.580 ;
        RECT 48.150 27.360 48.340 27.590 ;
        RECT 48.440 27.480 48.810 27.650 ;
        RECT 49.270 27.480 52.020 27.650 ;
        RECT 52.550 27.410 52.720 28.340 ;
        RECT 52.950 27.500 53.120 28.390 ;
        RECT 66.310 28.300 66.630 28.330 ;
        RECT 66.310 28.130 68.100 28.300 ;
        RECT 66.310 28.110 66.640 28.130 ;
        RECT 66.310 28.070 66.630 28.110 ;
        RECT 67.930 27.900 68.100 28.130 ;
        RECT 66.780 27.650 67.120 27.900 ;
        RECT 67.290 27.730 67.620 27.900 ;
        RECT 67.840 27.730 68.180 27.900 ;
        RECT 66.460 27.390 67.120 27.650 ;
        RECT 67.370 27.560 67.540 27.730 ;
        RECT 67.930 27.560 68.100 27.730 ;
        RECT 67.290 27.390 67.620 27.560 ;
        RECT 67.840 27.390 68.180 27.560 ;
        RECT 21.660 26.550 21.830 27.220 ;
        RECT 67.370 27.160 67.620 27.390 ;
        RECT 68.500 27.310 69.010 27.980 ;
        RECT 67.370 26.990 68.040 27.160 ;
        RECT 38.870 26.850 39.040 26.900 ;
        RECT 38.840 26.630 39.060 26.850 ;
        RECT 38.870 26.570 39.040 26.630 ;
        RECT 39.390 26.490 39.720 26.670 ;
        RECT 42.530 26.660 42.700 26.710 ;
        RECT 39.970 26.490 42.130 26.660 ;
        RECT 42.370 26.490 42.700 26.660 ;
        RECT 42.990 26.520 43.200 26.850 ;
        RECT 39.420 26.050 39.690 26.490 ;
        RECT 40.900 26.230 41.230 26.490 ;
        RECT 42.440 26.350 42.700 26.490 ;
        RECT 43.440 26.350 43.620 26.790 ;
        RECT 45.040 26.690 45.430 26.740 ;
        RECT 44.170 26.630 45.430 26.690 ;
        RECT 44.170 26.520 45.510 26.630 ;
        RECT 45.040 26.460 45.510 26.520 ;
        RECT 45.980 26.480 46.940 26.650 ;
        RECT 45.040 26.450 45.420 26.460 ;
        RECT 39.460 26.040 39.690 26.050 ;
        RECT 42.440 26.180 43.620 26.350 ;
        RECT 42.440 26.040 42.700 26.180 ;
        RECT 39.460 25.870 40.220 26.040 ;
        RECT 40.470 25.870 41.640 26.040 ;
        RECT 41.880 26.010 42.700 26.040 ;
        RECT 41.880 25.870 42.990 26.010 ;
        RECT 40.870 25.770 41.220 25.870 ;
        RECT 42.530 25.840 42.990 25.870 ;
        RECT 43.440 26.000 44.630 26.010 ;
        RECT 43.440 25.840 44.920 26.000 ;
        RECT 43.480 25.820 44.920 25.840 ;
        RECT 44.460 25.780 44.920 25.820 ;
        RECT 44.630 25.760 44.920 25.780 ;
        RECT 45.250 25.690 45.420 26.450 ;
        RECT 46.760 26.020 46.940 26.480 ;
        RECT 47.910 26.470 48.080 26.820 ;
        RECT 67.370 26.760 67.620 26.990 ;
        RECT 47.850 26.300 48.080 26.470 ;
        RECT 48.150 26.460 48.340 26.690 ;
        RECT 54.870 26.660 55.190 26.700 ;
        RECT 48.440 26.400 48.810 26.570 ;
        RECT 49.270 26.400 52.020 26.570 ;
        RECT 47.910 26.260 48.080 26.300 ;
        RECT 51.200 26.220 51.540 26.400 ;
        RECT 45.620 25.840 46.220 26.010 ;
        RECT 46.680 25.850 47.010 26.020 ;
        RECT 45.620 25.690 46.070 25.840 ;
        RECT 47.980 25.660 48.150 26.080 ;
        RECT 48.790 25.950 49.030 25.990 ;
        RECT 51.570 25.950 51.740 25.960 ;
        RECT 48.460 25.780 49.030 25.950 ;
        RECT 49.270 25.780 50.610 25.950 ;
        RECT 51.060 25.780 52.020 25.950 ;
        RECT 48.790 25.750 49.030 25.780 ;
        RECT 52.550 25.710 52.720 26.640 ;
        RECT 52.950 25.660 53.120 26.550 ;
        RECT 54.870 26.470 55.200 26.660 ;
        RECT 66.460 26.500 67.120 26.760 ;
        RECT 67.290 26.590 67.620 26.760 ;
        RECT 67.840 26.590 68.180 26.760 ;
        RECT 54.870 26.440 55.190 26.470 ;
        RECT 54.920 25.740 55.100 26.440 ;
        RECT 66.780 26.250 67.120 26.500 ;
        RECT 67.370 26.420 67.540 26.590 ;
        RECT 67.930 26.420 68.100 26.590 ;
        RECT 67.290 26.250 67.620 26.420 ;
        RECT 67.840 26.250 68.180 26.420 ;
        RECT 66.310 26.040 66.630 26.080 ;
        RECT 66.310 26.020 66.640 26.040 ;
        RECT 67.930 26.020 68.100 26.250 ;
        RECT 68.500 26.170 69.010 26.840 ;
        RECT 66.310 25.850 68.100 26.020 ;
        RECT 66.310 25.820 66.630 25.850 ;
        RECT 54.920 25.700 55.240 25.740 ;
        RECT 21.120 25.620 21.460 25.650 ;
        RECT 20.430 25.450 20.750 25.490 ;
        RECT 20.570 25.320 20.740 25.450 ;
        RECT 21.120 25.430 21.470 25.620 ;
        RECT 54.920 25.510 55.250 25.700 ;
        RECT 54.920 25.480 55.240 25.510 ;
        RECT 21.120 25.390 21.460 25.430 ;
        RECT 21.120 25.320 21.290 25.390 ;
        RECT 15.610 25.120 15.930 25.150 ;
        RECT 16.710 25.120 17.030 25.150 ;
        RECT 15.600 24.930 15.930 25.120 ;
        RECT 16.700 24.930 17.030 25.120 ;
        RECT 15.610 24.890 15.930 24.930 ;
        RECT 16.710 24.890 17.030 24.930 ;
        RECT 17.490 23.870 17.660 25.090 ;
        RECT 15.610 23.750 15.930 23.780 ;
        RECT 16.710 23.750 17.030 23.780 ;
        RECT 15.600 23.560 15.930 23.750 ;
        RECT 16.700 23.560 17.030 23.750 ;
        RECT 47.660 23.740 47.830 23.830 ;
        RECT 15.610 23.520 15.930 23.560 ;
        RECT 16.710 23.520 17.030 23.560 ;
        RECT 47.580 23.700 47.900 23.740 ;
        RECT 47.580 23.510 47.910 23.700 ;
        RECT 15.680 23.110 15.850 23.490 ;
        RECT 16.230 23.110 16.400 23.490 ;
        RECT 16.780 23.110 16.950 23.490 ;
        RECT 47.580 23.480 47.900 23.510 ;
        RECT 13.960 23.020 14.280 23.050 ;
        RECT 15.060 23.020 15.380 23.050 ;
        RECT 16.150 23.020 16.470 23.050 ;
        RECT 13.950 22.830 14.280 23.020 ;
        RECT 15.050 22.830 15.380 23.020 ;
        RECT 16.140 22.830 16.470 23.020 ;
        RECT 12.380 20.400 12.550 22.800 ;
        RECT 12.930 20.400 13.100 22.800 ;
        RECT 13.480 20.400 13.650 22.800 ;
        RECT 13.960 22.790 14.280 22.830 ;
        RECT 14.030 21.710 14.200 22.790 ;
        RECT 13.950 21.680 14.270 21.710 ;
        RECT 13.940 21.490 14.270 21.680 ;
        RECT 13.950 21.450 14.270 21.490 ;
        RECT 14.030 20.400 14.200 21.450 ;
        RECT 14.580 21.010 14.750 22.800 ;
        RECT 15.060 22.790 15.380 22.830 ;
        RECT 16.150 22.790 16.470 22.830 ;
        RECT 15.130 21.700 15.300 22.790 ;
        RECT 15.060 21.670 15.380 21.700 ;
        RECT 15.050 21.480 15.380 21.670 ;
        RECT 16.150 21.650 16.470 21.680 ;
        RECT 15.060 21.440 15.380 21.480 ;
        RECT 16.140 21.460 16.470 21.650 ;
        RECT 23.820 21.590 24.580 22.010 ;
        RECT 14.510 20.980 14.830 21.010 ;
        RECT 14.500 20.790 14.830 20.980 ;
        RECT 14.510 20.750 14.830 20.790 ;
        RECT 14.580 20.400 14.750 20.750 ;
        RECT 15.130 20.400 15.300 21.440 ;
        RECT 16.150 21.420 16.470 21.460 ;
        RECT 15.610 20.970 15.930 21.000 ;
        RECT 16.700 20.970 17.020 21.000 ;
        RECT 15.600 20.780 15.930 20.970 ;
        RECT 16.690 20.780 17.020 20.970 ;
        RECT 23.840 20.800 24.580 21.590 ;
        RECT 47.660 20.960 47.830 23.480 ;
        RECT 48.210 23.060 48.380 23.830 ;
        RECT 48.760 23.740 48.930 23.830 ;
        RECT 48.670 23.700 48.990 23.740 ;
        RECT 48.670 23.510 49.000 23.700 ;
        RECT 48.670 23.480 48.990 23.510 ;
        RECT 48.130 23.020 48.450 23.060 ;
        RECT 48.130 22.830 48.460 23.020 ;
        RECT 48.130 22.800 48.450 22.830 ;
        RECT 48.210 21.690 48.380 22.800 ;
        RECT 48.130 21.650 48.450 21.690 ;
        RECT 48.130 21.460 48.460 21.650 ;
        RECT 48.130 21.430 48.450 21.460 ;
        RECT 47.570 20.920 47.890 20.960 ;
        RECT 15.610 20.740 15.930 20.780 ;
        RECT 16.700 20.740 17.020 20.780 ;
        RECT 47.570 20.730 47.900 20.920 ;
        RECT 47.570 20.700 47.890 20.730 ;
        RECT 47.660 19.590 47.830 20.700 ;
        RECT 47.570 19.550 47.890 19.590 ;
        RECT 47.570 19.360 47.900 19.550 ;
        RECT 47.570 19.330 47.890 19.360 ;
        RECT 46.890 19.120 47.400 19.200 ;
        RECT 46.890 18.870 47.410 19.120 ;
        RECT 46.900 18.190 47.410 18.870 ;
        RECT 47.660 18.510 47.830 19.330 ;
        RECT 48.210 18.910 48.380 21.430 ;
        RECT 48.760 20.960 48.930 23.480 ;
        RECT 49.310 23.040 49.480 23.830 ;
        RECT 49.860 23.730 50.030 23.830 ;
        RECT 49.770 23.690 50.090 23.730 ;
        RECT 49.770 23.500 50.100 23.690 ;
        RECT 49.770 23.470 50.090 23.500 ;
        RECT 49.220 23.000 49.540 23.040 ;
        RECT 49.220 22.810 49.550 23.000 ;
        RECT 49.220 22.780 49.540 22.810 ;
        RECT 49.310 21.690 49.480 22.780 ;
        RECT 49.220 21.650 49.540 21.690 ;
        RECT 49.220 21.460 49.550 21.650 ;
        RECT 49.220 21.430 49.540 21.460 ;
        RECT 48.670 20.920 48.990 20.960 ;
        RECT 48.670 20.730 49.000 20.920 ;
        RECT 48.670 20.700 48.990 20.730 ;
        RECT 48.760 19.590 48.930 20.700 ;
        RECT 48.670 19.550 48.990 19.590 ;
        RECT 48.670 19.360 49.000 19.550 ;
        RECT 48.670 19.330 48.990 19.360 ;
        RECT 48.130 18.870 48.450 18.910 ;
        RECT 48.130 18.680 48.460 18.870 ;
        RECT 48.130 18.650 48.450 18.680 ;
        RECT 48.210 18.500 48.380 18.650 ;
        RECT 48.760 18.500 48.930 19.330 ;
        RECT 49.310 18.910 49.480 21.430 ;
        RECT 49.860 20.960 50.030 23.470 ;
        RECT 50.410 23.030 50.580 23.830 ;
        RECT 50.950 23.100 51.120 23.860 ;
        RECT 51.560 23.100 51.730 23.860 ;
        RECT 52.100 23.030 52.270 23.830 ;
        RECT 52.650 23.730 52.820 23.830 ;
        RECT 52.590 23.690 52.910 23.730 ;
        RECT 52.580 23.500 52.910 23.690 ;
        RECT 52.590 23.470 52.910 23.500 ;
        RECT 50.330 22.990 50.650 23.030 ;
        RECT 52.030 22.990 52.350 23.030 ;
        RECT 50.330 22.800 50.660 22.990 ;
        RECT 52.020 22.800 52.350 22.990 ;
        RECT 50.330 22.770 50.650 22.800 ;
        RECT 52.030 22.770 52.350 22.800 ;
        RECT 50.410 21.690 50.580 22.770 ;
        RECT 52.100 21.690 52.270 22.770 ;
        RECT 50.320 21.650 50.640 21.690 ;
        RECT 52.040 21.650 52.360 21.690 ;
        RECT 50.320 21.460 50.650 21.650 ;
        RECT 52.030 21.460 52.360 21.650 ;
        RECT 50.320 21.430 50.640 21.460 ;
        RECT 52.040 21.430 52.360 21.460 ;
        RECT 49.770 20.920 50.090 20.960 ;
        RECT 49.770 20.730 50.100 20.920 ;
        RECT 49.770 20.700 50.090 20.730 ;
        RECT 49.860 19.590 50.030 20.700 ;
        RECT 49.770 19.550 50.090 19.590 ;
        RECT 49.770 19.360 50.100 19.550 ;
        RECT 49.770 19.330 50.090 19.360 ;
        RECT 49.220 18.870 49.540 18.910 ;
        RECT 49.220 18.680 49.550 18.870 ;
        RECT 49.220 18.650 49.540 18.680 ;
        RECT 49.310 18.500 49.480 18.650 ;
        RECT 49.860 18.500 50.030 19.330 ;
        RECT 50.410 18.920 50.580 21.430 ;
        RECT 52.100 18.920 52.270 21.430 ;
        RECT 52.650 20.960 52.820 23.470 ;
        RECT 53.200 23.040 53.370 23.830 ;
        RECT 53.750 23.740 53.920 23.830 ;
        RECT 53.690 23.700 54.010 23.740 ;
        RECT 53.680 23.510 54.010 23.700 ;
        RECT 53.690 23.480 54.010 23.510 ;
        RECT 53.140 23.000 53.460 23.040 ;
        RECT 53.130 22.810 53.460 23.000 ;
        RECT 53.140 22.780 53.460 22.810 ;
        RECT 53.200 21.690 53.370 22.780 ;
        RECT 53.140 21.650 53.460 21.690 ;
        RECT 53.130 21.460 53.460 21.650 ;
        RECT 53.140 21.430 53.460 21.460 ;
        RECT 52.590 20.920 52.910 20.960 ;
        RECT 52.580 20.730 52.910 20.920 ;
        RECT 52.590 20.700 52.910 20.730 ;
        RECT 52.650 19.590 52.820 20.700 ;
        RECT 52.590 19.550 52.910 19.590 ;
        RECT 52.580 19.360 52.910 19.550 ;
        RECT 52.590 19.330 52.910 19.360 ;
        RECT 50.320 18.880 50.640 18.920 ;
        RECT 52.040 18.880 52.360 18.920 ;
        RECT 50.320 18.690 50.650 18.880 ;
        RECT 52.030 18.690 52.360 18.880 ;
        RECT 50.320 18.660 50.640 18.690 ;
        RECT 52.040 18.660 52.360 18.690 ;
        RECT 50.410 18.500 50.580 18.660 ;
        RECT 52.100 18.500 52.270 18.660 ;
        RECT 52.650 18.500 52.820 19.330 ;
        RECT 53.200 18.910 53.370 21.430 ;
        RECT 53.750 20.960 53.920 23.480 ;
        RECT 54.300 23.060 54.470 23.830 ;
        RECT 54.850 23.740 55.020 23.830 ;
        RECT 57.470 23.770 57.640 23.860 ;
        RECT 54.780 23.700 55.100 23.740 ;
        RECT 54.770 23.510 55.100 23.700 ;
        RECT 57.390 23.730 57.710 23.770 ;
        RECT 57.390 23.540 57.720 23.730 ;
        RECT 57.390 23.510 57.710 23.540 ;
        RECT 54.780 23.480 55.100 23.510 ;
        RECT 54.230 23.020 54.550 23.060 ;
        RECT 54.220 22.830 54.550 23.020 ;
        RECT 54.230 22.800 54.550 22.830 ;
        RECT 54.300 21.690 54.470 22.800 ;
        RECT 54.230 21.650 54.550 21.690 ;
        RECT 54.220 21.460 54.550 21.650 ;
        RECT 54.230 21.430 54.550 21.460 ;
        RECT 53.690 20.920 54.010 20.960 ;
        RECT 53.680 20.730 54.010 20.920 ;
        RECT 53.690 20.700 54.010 20.730 ;
        RECT 53.750 19.590 53.920 20.700 ;
        RECT 53.690 19.550 54.010 19.590 ;
        RECT 53.680 19.360 54.010 19.550 ;
        RECT 53.690 19.330 54.010 19.360 ;
        RECT 53.140 18.870 53.460 18.910 ;
        RECT 53.130 18.680 53.460 18.870 ;
        RECT 53.140 18.650 53.460 18.680 ;
        RECT 53.200 18.500 53.370 18.650 ;
        RECT 53.750 18.500 53.920 19.330 ;
        RECT 54.300 18.910 54.470 21.430 ;
        RECT 54.850 20.960 55.020 23.480 ;
        RECT 57.470 20.990 57.640 23.510 ;
        RECT 58.020 23.090 58.190 23.860 ;
        RECT 58.570 23.770 58.740 23.860 ;
        RECT 58.480 23.730 58.800 23.770 ;
        RECT 58.480 23.540 58.810 23.730 ;
        RECT 58.480 23.510 58.800 23.540 ;
        RECT 57.940 23.050 58.260 23.090 ;
        RECT 57.940 22.860 58.270 23.050 ;
        RECT 57.940 22.830 58.260 22.860 ;
        RECT 58.020 21.720 58.190 22.830 ;
        RECT 57.940 21.680 58.260 21.720 ;
        RECT 57.940 21.490 58.270 21.680 ;
        RECT 57.940 21.460 58.260 21.490 ;
        RECT 54.790 20.920 55.110 20.960 ;
        RECT 54.780 20.730 55.110 20.920 ;
        RECT 57.380 20.950 57.700 20.990 ;
        RECT 57.380 20.760 57.710 20.950 ;
        RECT 57.380 20.730 57.700 20.760 ;
        RECT 54.790 20.700 55.110 20.730 ;
        RECT 54.850 19.590 55.020 20.700 ;
        RECT 57.470 19.620 57.640 20.730 ;
        RECT 54.790 19.550 55.110 19.590 ;
        RECT 54.780 19.360 55.110 19.550 ;
        RECT 57.380 19.580 57.700 19.620 ;
        RECT 57.380 19.390 57.710 19.580 ;
        RECT 57.380 19.360 57.700 19.390 ;
        RECT 54.790 19.330 55.110 19.360 ;
        RECT 54.230 18.870 54.550 18.910 ;
        RECT 54.220 18.680 54.550 18.870 ;
        RECT 54.230 18.650 54.550 18.680 ;
        RECT 54.300 18.500 54.470 18.650 ;
        RECT 54.850 18.510 55.020 19.330 ;
        RECT 55.280 19.120 55.790 19.200 ;
        RECT 55.270 18.870 55.790 19.120 ;
        RECT 56.700 19.150 57.210 19.230 ;
        RECT 56.700 18.900 57.220 19.150 ;
        RECT 55.270 18.190 55.780 18.870 ;
        RECT 56.710 18.220 57.220 18.900 ;
        RECT 57.470 18.540 57.640 19.360 ;
        RECT 58.020 18.940 58.190 21.460 ;
        RECT 58.570 20.990 58.740 23.510 ;
        RECT 59.120 23.070 59.290 23.860 ;
        RECT 59.670 23.760 59.840 23.860 ;
        RECT 59.580 23.720 59.900 23.760 ;
        RECT 59.580 23.530 59.910 23.720 ;
        RECT 59.580 23.500 59.900 23.530 ;
        RECT 59.030 23.030 59.350 23.070 ;
        RECT 59.030 22.840 59.360 23.030 ;
        RECT 59.030 22.810 59.350 22.840 ;
        RECT 59.120 21.720 59.290 22.810 ;
        RECT 59.030 21.680 59.350 21.720 ;
        RECT 59.030 21.490 59.360 21.680 ;
        RECT 59.030 21.460 59.350 21.490 ;
        RECT 58.480 20.950 58.800 20.990 ;
        RECT 58.480 20.760 58.810 20.950 ;
        RECT 58.480 20.730 58.800 20.760 ;
        RECT 58.570 19.620 58.740 20.730 ;
        RECT 58.480 19.580 58.800 19.620 ;
        RECT 58.480 19.390 58.810 19.580 ;
        RECT 58.480 19.360 58.800 19.390 ;
        RECT 57.940 18.900 58.260 18.940 ;
        RECT 57.940 18.710 58.270 18.900 ;
        RECT 57.940 18.680 58.260 18.710 ;
        RECT 58.020 18.530 58.190 18.680 ;
        RECT 58.570 18.530 58.740 19.360 ;
        RECT 59.120 18.940 59.290 21.460 ;
        RECT 59.670 20.990 59.840 23.500 ;
        RECT 60.220 23.060 60.390 23.860 ;
        RECT 60.760 23.130 60.930 23.890 ;
        RECT 61.370 23.130 61.540 23.890 ;
        RECT 61.910 23.060 62.080 23.860 ;
        RECT 62.460 23.760 62.630 23.860 ;
        RECT 62.400 23.720 62.720 23.760 ;
        RECT 62.390 23.530 62.720 23.720 ;
        RECT 62.400 23.500 62.720 23.530 ;
        RECT 60.140 23.020 60.460 23.060 ;
        RECT 61.840 23.020 62.160 23.060 ;
        RECT 60.140 22.830 60.470 23.020 ;
        RECT 61.830 22.830 62.160 23.020 ;
        RECT 60.140 22.800 60.460 22.830 ;
        RECT 61.840 22.800 62.160 22.830 ;
        RECT 60.220 21.720 60.390 22.800 ;
        RECT 61.910 21.720 62.080 22.800 ;
        RECT 60.130 21.680 60.450 21.720 ;
        RECT 61.850 21.680 62.170 21.720 ;
        RECT 60.130 21.490 60.460 21.680 ;
        RECT 61.840 21.490 62.170 21.680 ;
        RECT 60.130 21.460 60.450 21.490 ;
        RECT 61.850 21.460 62.170 21.490 ;
        RECT 59.580 20.950 59.900 20.990 ;
        RECT 59.580 20.760 59.910 20.950 ;
        RECT 59.580 20.730 59.900 20.760 ;
        RECT 59.670 19.620 59.840 20.730 ;
        RECT 59.580 19.580 59.900 19.620 ;
        RECT 59.580 19.390 59.910 19.580 ;
        RECT 59.580 19.360 59.900 19.390 ;
        RECT 59.030 18.900 59.350 18.940 ;
        RECT 59.030 18.710 59.360 18.900 ;
        RECT 59.030 18.680 59.350 18.710 ;
        RECT 59.120 18.530 59.290 18.680 ;
        RECT 59.670 18.530 59.840 19.360 ;
        RECT 60.220 18.950 60.390 21.460 ;
        RECT 61.910 18.950 62.080 21.460 ;
        RECT 62.460 20.990 62.630 23.500 ;
        RECT 63.010 23.070 63.180 23.860 ;
        RECT 63.560 23.770 63.730 23.860 ;
        RECT 63.500 23.730 63.820 23.770 ;
        RECT 63.490 23.540 63.820 23.730 ;
        RECT 63.500 23.510 63.820 23.540 ;
        RECT 62.950 23.030 63.270 23.070 ;
        RECT 62.940 22.840 63.270 23.030 ;
        RECT 62.950 22.810 63.270 22.840 ;
        RECT 63.010 21.720 63.180 22.810 ;
        RECT 62.950 21.680 63.270 21.720 ;
        RECT 62.940 21.490 63.270 21.680 ;
        RECT 62.950 21.460 63.270 21.490 ;
        RECT 62.400 20.950 62.720 20.990 ;
        RECT 62.390 20.760 62.720 20.950 ;
        RECT 62.400 20.730 62.720 20.760 ;
        RECT 62.460 19.620 62.630 20.730 ;
        RECT 62.400 19.580 62.720 19.620 ;
        RECT 62.390 19.390 62.720 19.580 ;
        RECT 62.400 19.360 62.720 19.390 ;
        RECT 60.130 18.910 60.450 18.950 ;
        RECT 61.850 18.910 62.170 18.950 ;
        RECT 60.130 18.720 60.460 18.910 ;
        RECT 61.840 18.720 62.170 18.910 ;
        RECT 60.130 18.690 60.450 18.720 ;
        RECT 61.850 18.690 62.170 18.720 ;
        RECT 60.220 18.530 60.390 18.690 ;
        RECT 61.910 18.530 62.080 18.690 ;
        RECT 62.460 18.530 62.630 19.360 ;
        RECT 63.010 18.940 63.180 21.460 ;
        RECT 63.560 20.990 63.730 23.510 ;
        RECT 64.110 23.090 64.280 23.860 ;
        RECT 64.660 23.770 64.830 23.860 ;
        RECT 64.590 23.730 64.910 23.770 ;
        RECT 64.580 23.540 64.910 23.730 ;
        RECT 64.590 23.510 64.910 23.540 ;
        RECT 64.040 23.050 64.360 23.090 ;
        RECT 64.030 22.860 64.360 23.050 ;
        RECT 64.040 22.830 64.360 22.860 ;
        RECT 64.110 21.720 64.280 22.830 ;
        RECT 64.040 21.680 64.360 21.720 ;
        RECT 64.030 21.490 64.360 21.680 ;
        RECT 64.040 21.460 64.360 21.490 ;
        RECT 63.500 20.950 63.820 20.990 ;
        RECT 63.490 20.760 63.820 20.950 ;
        RECT 63.500 20.730 63.820 20.760 ;
        RECT 63.560 19.620 63.730 20.730 ;
        RECT 63.500 19.580 63.820 19.620 ;
        RECT 63.490 19.390 63.820 19.580 ;
        RECT 63.500 19.360 63.820 19.390 ;
        RECT 62.950 18.900 63.270 18.940 ;
        RECT 62.940 18.710 63.270 18.900 ;
        RECT 62.950 18.680 63.270 18.710 ;
        RECT 63.010 18.530 63.180 18.680 ;
        RECT 63.560 18.530 63.730 19.360 ;
        RECT 64.110 18.940 64.280 21.460 ;
        RECT 64.660 20.990 64.830 23.510 ;
        RECT 64.600 20.950 64.920 20.990 ;
        RECT 64.590 20.760 64.920 20.950 ;
        RECT 64.600 20.730 64.920 20.760 ;
        RECT 64.660 19.620 64.830 20.730 ;
        RECT 64.600 19.580 64.920 19.620 ;
        RECT 64.590 19.390 64.920 19.580 ;
        RECT 64.600 19.360 64.920 19.390 ;
        RECT 64.040 18.900 64.360 18.940 ;
        RECT 64.030 18.710 64.360 18.900 ;
        RECT 64.040 18.680 64.360 18.710 ;
        RECT 64.110 18.530 64.280 18.680 ;
        RECT 64.660 18.540 64.830 19.360 ;
        RECT 65.090 19.150 65.600 19.230 ;
        RECT 65.080 18.900 65.600 19.150 ;
        RECT 65.080 18.220 65.590 18.900 ;
        RECT 66.650 17.500 66.820 19.900 ;
        RECT 67.200 17.500 67.370 19.900 ;
        RECT 67.750 17.500 67.920 19.900 ;
        RECT 68.300 18.850 68.470 19.900 ;
        RECT 68.850 19.550 69.020 19.900 ;
        RECT 68.780 19.510 69.100 19.550 ;
        RECT 68.770 19.320 69.100 19.510 ;
        RECT 68.780 19.290 69.100 19.320 ;
        RECT 68.220 18.810 68.540 18.850 ;
        RECT 68.210 18.620 68.540 18.810 ;
        RECT 68.220 18.590 68.540 18.620 ;
        RECT 68.300 17.510 68.470 18.590 ;
        RECT 68.230 17.470 68.550 17.510 ;
        RECT 68.850 17.500 69.020 19.290 ;
        RECT 69.400 18.860 69.570 19.900 ;
        RECT 69.880 19.520 70.200 19.560 ;
        RECT 70.970 19.520 71.290 19.560 ;
        RECT 69.870 19.330 70.200 19.520 ;
        RECT 70.960 19.330 71.290 19.520 ;
        RECT 69.880 19.300 70.200 19.330 ;
        RECT 70.970 19.300 71.290 19.330 ;
        RECT 69.330 18.820 69.650 18.860 ;
        RECT 70.420 18.840 70.740 18.880 ;
        RECT 69.320 18.630 69.650 18.820 ;
        RECT 70.410 18.650 70.740 18.840 ;
        RECT 69.330 18.600 69.650 18.630 ;
        RECT 70.420 18.620 70.740 18.650 ;
        RECT 69.400 17.510 69.570 18.600 ;
        RECT 69.330 17.470 69.650 17.510 ;
        RECT 70.420 17.470 70.740 17.510 ;
        RECT 68.220 17.280 68.550 17.470 ;
        RECT 69.320 17.280 69.650 17.470 ;
        RECT 70.410 17.280 70.740 17.470 ;
        RECT 68.230 17.250 68.550 17.280 ;
        RECT 69.330 17.250 69.650 17.280 ;
        RECT 70.420 17.250 70.740 17.280 ;
        RECT 66.650 14.720 66.820 17.120 ;
        RECT 67.200 14.720 67.370 17.120 ;
        RECT 67.750 14.720 67.920 17.120 ;
        RECT 68.300 14.740 68.470 17.190 ;
        RECT 68.850 16.780 69.020 17.190 ;
        RECT 68.780 16.740 69.100 16.780 ;
        RECT 68.770 16.550 69.100 16.740 ;
        RECT 68.780 16.520 69.100 16.550 ;
        RECT 68.850 15.410 69.020 16.520 ;
        RECT 68.780 15.370 69.100 15.410 ;
        RECT 68.770 15.180 69.100 15.370 ;
        RECT 68.780 15.150 69.100 15.180 ;
        RECT 68.230 14.700 68.550 14.740 ;
        RECT 68.850 14.720 69.020 15.150 ;
        RECT 69.400 14.730 69.570 17.190 ;
        RECT 69.950 16.810 70.120 17.190 ;
        RECT 70.500 16.810 70.670 17.190 ;
        RECT 71.050 16.810 71.220 17.190 ;
        RECT 69.880 16.740 70.200 16.780 ;
        RECT 70.980 16.740 71.300 16.780 ;
        RECT 69.870 16.550 70.200 16.740 ;
        RECT 70.970 16.550 71.300 16.740 ;
        RECT 69.880 16.520 70.200 16.550 ;
        RECT 70.980 16.520 71.300 16.550 ;
        RECT 69.880 15.370 70.200 15.410 ;
        RECT 70.980 15.370 71.300 15.410 ;
        RECT 69.870 15.180 70.200 15.370 ;
        RECT 70.970 15.180 71.300 15.370 ;
        RECT 71.760 15.210 71.930 16.430 ;
        RECT 102.290 15.920 102.520 16.030 ;
        RECT 102.190 15.750 106.850 15.920 ;
        RECT 105.170 15.470 105.500 15.640 ;
        RECT 106.130 15.470 106.460 15.640 ;
        RECT 107.090 15.470 107.420 15.640 ;
        RECT 108.050 15.470 108.380 15.640 ;
        RECT 107.750 15.270 107.940 15.280 ;
        RECT 103.410 15.230 107.210 15.240 ;
        RECT 107.720 15.230 107.980 15.270 ;
        RECT 69.880 15.150 70.200 15.180 ;
        RECT 70.980 15.150 71.300 15.180 ;
        RECT 103.410 15.070 107.980 15.230 ;
        RECT 106.980 15.060 107.980 15.070 ;
        RECT 71.470 14.760 71.980 15.020 ;
        RECT 106.980 14.960 107.210 15.060 ;
        RECT 105.170 14.790 105.500 14.960 ;
        RECT 106.130 14.790 106.460 14.960 ;
        RECT 106.980 14.790 107.420 14.960 ;
        RECT 107.720 14.950 107.980 15.060 ;
        RECT 108.050 14.790 108.380 14.960 ;
        RECT 13.420 14.070 13.590 14.230 ;
        RECT 13.360 14.040 13.680 14.070 ;
        RECT 13.350 13.850 13.680 14.040 ;
        RECT 13.360 13.810 13.680 13.850 ;
        RECT 13.420 11.300 13.590 13.810 ;
        RECT 13.970 13.400 14.140 14.230 ;
        RECT 14.520 14.080 14.690 14.230 ;
        RECT 14.460 14.050 14.780 14.080 ;
        RECT 14.450 13.860 14.780 14.050 ;
        RECT 14.460 13.820 14.780 13.860 ;
        RECT 13.910 13.370 14.230 13.400 ;
        RECT 13.900 13.180 14.230 13.370 ;
        RECT 13.910 13.140 14.230 13.180 ;
        RECT 13.970 12.030 14.140 13.140 ;
        RECT 13.910 12.000 14.230 12.030 ;
        RECT 13.900 11.810 14.230 12.000 ;
        RECT 13.910 11.770 14.230 11.810 ;
        RECT 13.360 11.270 13.680 11.300 ;
        RECT 13.350 11.080 13.680 11.270 ;
        RECT 13.360 11.040 13.680 11.080 ;
        RECT 13.420 9.960 13.590 11.040 ;
        RECT 13.350 9.930 13.670 9.960 ;
        RECT 13.340 9.740 13.670 9.930 ;
        RECT 13.350 9.700 13.670 9.740 ;
        RECT 12.880 8.870 13.050 9.630 ;
        RECT 13.420 8.900 13.590 9.700 ;
        RECT 13.970 9.260 14.140 11.770 ;
        RECT 14.520 11.300 14.690 13.820 ;
        RECT 15.070 13.400 15.240 14.230 ;
        RECT 15.620 14.080 15.790 14.230 ;
        RECT 15.550 14.050 15.870 14.080 ;
        RECT 15.540 13.860 15.870 14.050 ;
        RECT 15.550 13.820 15.870 13.860 ;
        RECT 15.010 13.370 15.330 13.400 ;
        RECT 15.000 13.180 15.330 13.370 ;
        RECT 15.010 13.140 15.330 13.180 ;
        RECT 15.070 12.030 15.240 13.140 ;
        RECT 15.010 12.000 15.330 12.030 ;
        RECT 15.000 11.810 15.330 12.000 ;
        RECT 15.010 11.770 15.330 11.810 ;
        RECT 14.460 11.270 14.780 11.300 ;
        RECT 14.450 11.080 14.780 11.270 ;
        RECT 14.460 11.040 14.780 11.080 ;
        RECT 14.520 9.950 14.690 11.040 ;
        RECT 14.460 9.920 14.780 9.950 ;
        RECT 14.450 9.730 14.780 9.920 ;
        RECT 14.460 9.690 14.780 9.730 ;
        RECT 13.910 9.230 14.230 9.260 ;
        RECT 13.900 9.040 14.230 9.230 ;
        RECT 13.910 9.000 14.230 9.040 ;
        RECT 13.970 8.900 14.140 9.000 ;
        RECT 14.520 8.900 14.690 9.690 ;
        RECT 15.070 9.250 15.240 11.770 ;
        RECT 15.620 11.300 15.790 13.820 ;
        RECT 16.170 13.400 16.340 14.220 ;
        RECT 16.590 13.860 17.100 14.540 ;
        RECT 68.220 14.510 68.550 14.700 ;
        RECT 69.330 14.690 69.650 14.730 ;
        RECT 70.420 14.690 70.740 14.730 ;
        RECT 68.230 14.480 68.550 14.510 ;
        RECT 69.320 14.500 69.650 14.690 ;
        RECT 70.410 14.500 70.740 14.690 ;
        RECT 69.330 14.470 69.650 14.500 ;
        RECT 70.420 14.470 70.740 14.500 ;
        RECT 71.460 14.690 71.980 14.760 ;
        RECT 71.460 14.010 71.970 14.690 ;
        RECT 106.980 14.600 107.210 14.790 ;
        RECT 107.750 14.600 107.940 14.610 ;
        RECT 102.290 14.310 102.520 14.420 ;
        RECT 106.980 14.390 107.990 14.600 ;
        RECT 102.190 14.140 106.670 14.310 ;
        RECT 106.980 14.030 107.210 14.390 ;
        RECT 107.720 14.280 107.980 14.390 ;
        RECT 105.170 13.860 105.500 14.030 ;
        RECT 106.130 13.860 106.460 14.030 ;
        RECT 106.980 13.860 107.420 14.030 ;
        RECT 108.050 13.860 108.380 14.030 ;
        RECT 16.590 13.610 17.110 13.860 ;
        RECT 106.980 13.630 107.210 13.860 ;
        RECT 16.600 13.530 17.110 13.610 ;
        RECT 103.440 13.460 107.210 13.630 ;
        RECT 16.110 13.370 16.430 13.400 ;
        RECT 16.100 13.180 16.430 13.370 ;
        RECT 106.980 13.350 107.210 13.460 ;
        RECT 16.110 13.140 16.430 13.180 ;
        RECT 16.170 12.030 16.340 13.140 ;
        RECT 18.170 12.900 20.560 13.270 ;
        RECT 105.170 13.180 105.500 13.350 ;
        RECT 106.130 13.180 106.460 13.350 ;
        RECT 106.980 13.180 107.420 13.350 ;
        RECT 108.050 13.290 108.380 13.350 ;
        RECT 107.700 13.270 108.380 13.290 ;
        RECT 107.680 13.180 108.380 13.270 ;
        RECT 16.110 12.000 16.430 12.030 ;
        RECT 16.100 11.810 16.430 12.000 ;
        RECT 16.110 11.770 16.430 11.810 ;
        RECT 15.550 11.270 15.870 11.300 ;
        RECT 15.540 11.080 15.870 11.270 ;
        RECT 15.550 11.040 15.870 11.080 ;
        RECT 15.620 9.930 15.790 11.040 ;
        RECT 15.550 9.900 15.870 9.930 ;
        RECT 15.540 9.710 15.870 9.900 ;
        RECT 15.550 9.670 15.870 9.710 ;
        RECT 15.010 9.220 15.330 9.250 ;
        RECT 15.000 9.030 15.330 9.220 ;
        RECT 15.010 8.990 15.330 9.030 ;
        RECT 15.070 8.900 15.240 8.990 ;
        RECT 15.620 8.900 15.790 9.670 ;
        RECT 16.170 9.250 16.340 11.770 ;
        RECT 18.220 9.640 20.560 12.900 ;
        RECT 102.290 12.710 102.520 12.820 ;
        RECT 102.190 12.540 106.690 12.710 ;
        RECT 106.980 12.420 107.210 13.180 ;
        RECT 107.680 13.100 108.130 13.180 ;
        RECT 107.700 13.080 108.130 13.100 ;
        RECT 105.170 12.250 105.500 12.420 ;
        RECT 106.130 12.250 106.460 12.420 ;
        RECT 106.980 12.250 107.420 12.420 ;
        RECT 108.050 12.250 108.380 12.420 ;
        RECT 106.980 12.020 107.210 12.250 ;
        RECT 103.450 11.850 107.210 12.020 ;
        RECT 106.980 11.740 107.210 11.850 ;
        RECT 103.750 11.660 104.180 11.680 ;
        RECT 103.730 11.490 104.180 11.660 ;
        RECT 105.170 11.570 105.500 11.740 ;
        RECT 106.130 11.570 106.460 11.740 ;
        RECT 106.980 11.570 107.420 11.740 ;
        RECT 108.050 11.680 108.380 11.740 ;
        RECT 107.700 11.660 108.380 11.680 ;
        RECT 107.680 11.570 108.380 11.660 ;
        RECT 103.750 11.470 104.180 11.490 ;
        RECT 102.290 11.090 102.520 11.200 ;
        RECT 102.190 10.920 106.690 11.090 ;
        RECT 106.980 10.420 107.210 11.570 ;
        RECT 107.680 11.490 108.130 11.570 ;
        RECT 107.700 11.470 108.130 11.490 ;
        RECT 103.440 10.410 107.210 10.420 ;
        RECT 103.430 10.250 107.210 10.410 ;
        RECT 103.430 10.240 103.760 10.250 ;
        RECT 105.350 10.240 105.680 10.250 ;
        RECT 106.310 10.240 106.640 10.250 ;
        RECT 104.230 10.020 104.660 10.040 ;
        RECT 104.230 9.850 104.680 10.020 ;
        RECT 104.230 9.830 104.660 9.850 ;
        RECT 18.220 9.630 20.550 9.640 ;
        RECT 102.290 9.490 102.520 9.600 ;
        RECT 102.190 9.320 106.640 9.490 ;
        RECT 103.430 9.310 103.760 9.320 ;
        RECT 104.390 9.310 104.720 9.320 ;
        RECT 105.350 9.310 105.680 9.320 ;
        RECT 106.310 9.310 106.640 9.320 ;
        RECT 16.100 9.220 16.420 9.250 ;
        RECT 16.090 9.030 16.420 9.220 ;
        RECT 16.100 8.990 16.420 9.030 ;
        RECT 16.170 8.900 16.340 8.990 ;
        RECT 106.980 8.800 107.210 10.250 ;
        RECT 107.690 10.050 108.120 10.070 ;
        RECT 107.670 9.880 108.120 10.050 ;
        RECT 107.690 9.860 108.120 9.880 ;
        RECT 103.420 8.630 107.210 8.800 ;
        RECT 105.660 8.440 106.090 8.460 ;
        RECT 105.640 8.270 106.090 8.440 ;
        RECT 105.660 8.250 106.090 8.270 ;
        RECT 102.290 7.870 102.520 7.980 ;
        RECT 102.190 7.700 106.690 7.870 ;
        RECT 106.980 7.590 107.210 8.630 ;
        RECT 107.700 8.430 108.130 8.450 ;
        RECT 107.680 8.260 108.130 8.430 ;
        RECT 107.700 8.240 108.130 8.260 ;
        RECT 105.170 7.420 105.500 7.590 ;
        RECT 106.130 7.420 106.460 7.590 ;
        RECT 106.980 7.420 107.420 7.590 ;
        RECT 108.050 7.420 108.380 7.590 ;
        RECT 106.980 7.180 107.210 7.420 ;
        RECT 103.420 7.010 107.210 7.180 ;
        RECT 106.980 6.910 107.210 7.010 ;
        RECT 105.170 6.740 105.500 6.910 ;
        RECT 106.130 6.740 106.460 6.910 ;
        RECT 106.980 6.740 107.420 6.910 ;
        RECT 108.050 6.840 108.380 6.910 ;
        RECT 107.690 6.820 108.380 6.840 ;
        RECT 107.670 6.740 108.380 6.820 ;
        RECT 102.290 6.270 102.520 6.380 ;
        RECT 102.190 6.100 106.610 6.270 ;
        RECT 106.980 5.980 107.210 6.740 ;
        RECT 107.670 6.650 108.120 6.740 ;
        RECT 107.690 6.630 108.120 6.650 ;
        RECT 105.170 5.810 105.500 5.980 ;
        RECT 106.130 5.810 106.460 5.980 ;
        RECT 106.980 5.810 107.420 5.980 ;
        RECT 108.050 5.810 108.380 5.980 ;
        RECT 106.980 5.590 107.210 5.810 ;
        RECT 103.420 5.420 107.220 5.590 ;
        RECT 106.980 5.300 107.210 5.420 ;
        RECT 105.170 5.130 105.500 5.300 ;
        RECT 106.130 5.130 106.460 5.300 ;
        RECT 106.980 5.130 107.420 5.300 ;
        RECT 102.290 4.640 102.520 4.760 ;
        RECT 102.190 4.470 106.650 4.640 ;
        RECT 106.980 4.370 107.210 5.130 ;
        RECT 107.490 4.780 107.700 5.210 ;
        RECT 108.050 5.130 108.380 5.300 ;
        RECT 107.510 4.760 107.680 4.780 ;
        RECT 105.170 4.200 105.500 4.370 ;
        RECT 106.130 4.200 106.460 4.370 ;
        RECT 106.980 4.200 107.420 4.370 ;
        RECT 108.050 4.200 108.380 4.370 ;
        RECT 106.980 3.980 107.210 4.200 ;
        RECT 103.420 3.810 107.210 3.980 ;
        RECT 105.170 3.520 105.500 3.690 ;
        RECT 106.130 3.520 106.460 3.690 ;
        RECT 107.090 3.520 107.420 3.690 ;
        RECT 108.050 3.640 108.380 3.690 ;
        RECT 107.690 3.620 108.380 3.640 ;
        RECT 107.670 3.520 108.380 3.620 ;
        RECT 107.670 3.450 108.120 3.520 ;
        RECT 107.690 3.430 108.120 3.450 ;
        RECT 108.400 2.640 108.770 17.510 ;
        RECT 108.400 2.390 108.780 2.640 ;
        RECT 104.450 1.910 104.880 1.930 ;
        RECT 105.390 1.910 105.820 1.930 ;
        RECT 107.650 1.910 108.080 1.930 ;
        RECT 104.430 1.740 104.880 1.910 ;
        RECT 105.370 1.740 105.820 1.910 ;
        RECT 106.340 1.890 106.770 1.910 ;
        RECT 104.450 1.720 104.880 1.740 ;
        RECT 105.390 1.720 105.820 1.740 ;
        RECT 106.320 1.720 106.770 1.890 ;
        RECT 107.630 1.740 108.080 1.910 ;
        RECT 107.650 1.720 108.080 1.740 ;
        RECT 106.340 1.700 106.770 1.720 ;
      LAYER mcon ;
        RECT 8.370 66.980 8.540 67.150 ;
        RECT 8.370 66.290 8.540 66.460 ;
        RECT 19.440 66.350 19.610 66.520 ;
        RECT 19.440 65.900 19.610 66.070 ;
        RECT 24.140 66.300 24.310 66.470 ;
        RECT 24.140 65.850 24.310 66.020 ;
        RECT 11.480 64.810 11.650 64.980 ;
        RECT 12.840 64.890 13.010 65.060 ;
        RECT 13.530 64.880 13.700 65.050 ;
        RECT 8.370 64.180 8.540 64.350 ;
        RECT 8.370 63.490 8.540 63.660 ;
        RECT 8.370 62.630 8.540 62.800 ;
        RECT 8.370 61.940 8.540 62.110 ;
        RECT 19.440 63.360 19.610 63.530 ;
        RECT 19.440 62.910 19.610 63.080 ;
        RECT 19.440 62.350 19.610 62.520 ;
        RECT 19.440 61.900 19.610 62.070 ;
        RECT 23.360 62.840 23.530 63.010 ;
        RECT 10.760 61.150 10.930 61.320 ;
        RECT 20.620 61.170 20.790 61.340 ;
        RECT 19.890 59.380 20.320 60.120 ;
        RECT 40.990 57.960 41.200 58.170 ;
        RECT 44.730 57.980 44.900 58.150 ;
        RECT 39.520 57.590 39.690 57.760 ;
        RECT 45.770 58.020 45.940 58.190 ;
        RECT 46.810 57.680 46.980 57.850 ;
        RECT 46.810 57.320 46.980 57.490 ;
        RECT 40.990 56.210 41.200 56.420 ;
        RECT 44.730 56.230 44.900 56.400 ;
        RECT 39.520 55.840 39.690 56.010 ;
        RECT 45.770 56.270 45.940 56.440 ;
        RECT 68.180 56.220 68.440 57.040 ;
        RECT 80.130 56.250 80.450 57.040 ;
        RECT 83.180 56.680 83.360 56.850 ;
        RECT 83.510 56.740 83.680 56.910 ;
        RECT 81.370 56.380 81.540 56.550 ;
        RECT 46.810 55.930 46.980 56.100 ;
        RECT 46.810 55.570 46.980 55.740 ;
        RECT 81.720 55.540 81.900 55.730 ;
        RECT 17.770 54.600 17.940 54.770 ;
        RECT 18.860 54.610 19.030 54.780 ;
        RECT 40.990 54.460 41.200 54.670 ;
        RECT 44.730 54.480 44.900 54.650 ;
        RECT 17.340 54.100 17.510 54.270 ;
        RECT 19.810 54.120 19.980 54.290 ;
        RECT 39.520 54.090 39.690 54.260 ;
        RECT 17.780 53.610 17.950 53.780 ;
        RECT 18.870 53.620 19.040 53.790 ;
        RECT 83.980 56.180 84.150 56.350 ;
        RECT 86.320 55.800 86.490 55.970 ;
        RECT 86.320 55.350 86.490 55.520 ;
        RECT 82.800 54.980 82.970 55.150 ;
        RECT 91.770 55.200 92.040 55.470 ;
        RECT 45.770 54.520 45.940 54.690 ;
        RECT 83.510 54.750 83.680 54.920 ;
        RECT 46.810 54.180 46.980 54.350 ;
        RECT 46.810 53.820 46.980 53.990 ;
        RECT 17.320 53.180 17.490 53.350 ;
        RECT 17.780 52.620 17.950 52.790 ;
        RECT 18.870 52.630 19.040 52.800 ;
        RECT 40.990 52.710 41.200 52.920 ;
        RECT 44.730 52.730 44.900 52.900 ;
        RECT 17.300 52.190 17.470 52.360 ;
        RECT 18.800 52.240 18.970 52.410 ;
        RECT 39.520 52.340 39.690 52.510 ;
        RECT 20.100 52.140 20.270 52.310 ;
        RECT 45.770 52.770 45.940 52.940 ;
        RECT 81.720 52.740 81.900 52.930 ;
        RECT 46.810 52.430 46.980 52.600 ;
        RECT 46.810 52.070 46.980 52.240 ;
        RECT 52.290 52.000 52.470 52.170 ;
        RECT 50.480 51.700 50.650 51.870 ;
        RECT 18.800 51.250 18.970 51.420 ;
        RECT 20.100 51.150 20.270 51.320 ;
        RECT 39.520 50.640 39.690 50.810 ;
        RECT 47.970 51.160 48.140 51.330 ;
        RECT 46.810 50.910 46.980 51.080 ;
        RECT 48.810 51.040 48.980 51.210 ;
        RECT 49.560 51.040 49.730 51.210 ;
        RECT 18.800 50.260 18.970 50.430 ;
        RECT 19.380 50.020 19.550 50.190 ;
        RECT 20.100 50.160 20.270 50.330 ;
        RECT 40.990 50.230 41.200 50.440 ;
        RECT 44.730 50.250 44.900 50.420 ;
        RECT 50.830 50.860 51.010 51.050 ;
        RECT 46.810 50.550 46.980 50.720 ;
        RECT 83.520 53.680 83.690 53.850 ;
        RECT 83.980 53.860 84.150 54.030 ;
        RECT 89.350 54.170 89.520 54.340 ;
        RECT 82.790 53.290 82.960 53.460 ;
        RECT 91.770 53.470 92.040 53.740 ;
        RECT 109.110 53.520 109.280 53.690 ;
        RECT 112.610 53.520 112.780 53.690 ;
        RECT 109.180 53.120 109.350 53.290 ;
        RECT 111.870 53.130 112.040 53.300 ;
        RECT 86.320 52.850 86.490 53.020 ;
        RECT 111.020 52.910 111.190 53.080 ;
        RECT 83.970 52.280 84.140 52.450 ;
        RECT 86.320 52.400 86.490 52.570 ;
        RECT 107.280 52.510 107.450 52.680 ;
        RECT 109.960 52.690 110.130 52.860 ;
        RECT 112.150 52.900 112.320 53.070 ;
        RECT 111.530 52.690 111.700 52.860 ;
        RECT 112.950 52.890 113.120 53.060 ;
        RECT 114.120 53.150 114.290 53.320 ;
        RECT 81.370 51.920 81.540 52.090 ;
        RECT 83.180 51.620 83.360 51.790 ;
        RECT 83.540 51.770 83.710 51.940 ;
        RECT 100.440 51.930 100.610 52.100 ;
        RECT 52.150 50.870 52.320 51.040 ;
        RECT 45.770 50.210 45.940 50.380 ;
        RECT 48.150 50.330 48.320 50.500 ;
        RECT 52.540 50.710 52.710 50.880 ;
        RECT 52.940 51.160 53.110 51.330 ;
        RECT 52.940 50.800 53.110 50.970 ;
        RECT 57.320 51.120 57.490 51.290 ;
        RECT 59.410 51.280 59.580 51.450 ;
        RECT 96.780 51.330 97.050 51.600 ;
        RECT 100.440 51.480 100.610 51.650 ;
        RECT 105.610 51.680 105.780 51.850 ;
        RECT 57.320 50.670 57.490 50.840 ;
        RECT 60.880 50.520 61.150 50.790 ;
        RECT 109.330 52.290 109.500 52.460 ;
        RECT 111.820 52.480 111.990 52.650 ;
        RECT 106.920 51.670 107.100 51.860 ;
        RECT 108.210 51.770 108.380 51.940 ;
        RECT 113.610 51.920 113.780 52.090 ;
        RECT 109.960 51.550 110.130 51.720 ;
        RECT 111.530 51.550 111.700 51.720 ;
        RECT 111.820 51.640 111.990 51.810 ;
        RECT 111.020 51.330 111.190 51.500 ;
        RECT 112.150 51.340 112.320 51.510 ;
        RECT 112.950 51.230 113.120 51.400 ;
        RECT 99.300 50.300 99.470 50.470 ;
        RECT 39.520 48.890 39.690 49.060 ;
        RECT 46.810 49.160 46.980 49.330 ;
        RECT 48.150 49.430 48.320 49.600 ;
        RECT 40.990 48.480 41.200 48.690 ;
        RECT 44.730 48.500 44.900 48.670 ;
        RECT 58.460 49.490 58.630 49.660 ;
        RECT 96.780 49.600 97.050 49.870 ;
        RECT 46.810 48.800 46.980 48.970 ;
        RECT 45.770 48.460 45.940 48.630 ;
        RECT 48.810 48.720 48.980 48.890 ;
        RECT 49.560 48.720 49.730 48.890 ;
        RECT 51.560 48.730 51.730 48.900 ;
        RECT 47.970 47.960 48.140 48.130 ;
        RECT 50.830 48.060 51.010 48.250 ;
        RECT 39.520 47.140 39.690 47.310 ;
        RECT 48.810 47.840 48.980 48.010 ;
        RECT 49.560 47.840 49.730 48.010 ;
        RECT 52.540 49.050 52.710 49.220 ;
        RECT 52.940 49.320 53.110 49.490 ;
        RECT 52.940 48.960 53.110 49.130 ;
        RECT 60.880 48.790 61.150 49.060 ;
        RECT 100.440 48.980 100.610 49.150 ;
        RECT 78.290 48.440 78.460 48.610 ;
        RECT 80.980 48.450 81.150 48.620 ;
        RECT 52.150 48.110 52.320 48.280 ;
        RECT 57.320 48.170 57.490 48.340 ;
        RECT 46.810 47.410 46.980 47.580 ;
        RECT 40.990 46.730 41.200 46.940 ;
        RECT 44.730 46.750 44.900 46.920 ;
        RECT 46.810 47.050 46.980 47.220 ;
        RECT 48.150 47.130 48.320 47.300 ;
        RECT 50.480 47.240 50.650 47.410 ;
        RECT 52.540 47.510 52.710 47.680 ;
        RECT 45.770 46.710 45.940 46.880 ;
        RECT 52.940 47.960 53.110 48.130 ;
        RECT 52.940 47.600 53.110 47.770 ;
        RECT 82.060 48.210 82.230 48.380 ;
        RECT 83.230 48.470 83.400 48.640 ;
        RECT 105.610 48.920 105.780 49.090 ;
        RECT 100.440 48.530 100.610 48.700 ;
        RECT 111.870 50.990 112.040 51.160 ;
        RECT 109.110 50.720 109.280 50.890 ;
        RECT 114.170 50.930 114.340 51.100 ;
        RECT 108.600 50.510 108.770 50.700 ;
        RECT 112.610 50.720 112.780 50.890 ;
        RECT 108.940 50.490 109.110 50.660 ;
        RECT 109.110 50.320 109.280 50.490 ;
        RECT 111.870 50.130 112.040 50.300 ;
        RECT 112.610 50.320 112.780 50.490 ;
        RECT 114.160 50.210 114.330 50.380 ;
        RECT 109.470 49.610 109.640 49.780 ;
        RECT 111.020 49.710 111.190 49.880 ;
        RECT 112.150 49.700 112.320 49.870 ;
        RECT 112.950 49.890 113.120 50.060 ;
        RECT 109.960 49.490 110.130 49.660 ;
        RECT 111.530 49.490 111.700 49.660 ;
        RECT 111.820 49.480 111.990 49.650 ;
        RECT 113.610 49.330 113.780 49.500 ;
        RECT 106.920 48.870 107.100 49.060 ;
        RECT 111.820 48.640 111.990 48.810 ;
        RECT 57.320 47.720 57.490 47.890 ;
        RECT 76.390 47.830 76.560 48.000 ;
        RECT 59.440 47.590 59.610 47.760 ;
        RECT 52.290 46.940 52.470 47.110 ;
        RECT 69.550 47.250 69.720 47.420 ;
        RECT 65.890 46.650 66.160 46.920 ;
        RECT 69.550 46.800 69.720 46.970 ;
        RECT 74.720 47.000 74.890 47.170 ;
        RECT 48.150 46.230 48.320 46.400 ;
        RECT 39.520 45.390 39.690 45.560 ;
        RECT 52.540 45.850 52.710 46.020 ;
        RECT 46.810 45.660 46.980 45.830 ;
        RECT 40.990 44.980 41.200 45.190 ;
        RECT 44.730 45.000 44.900 45.170 ;
        RECT 46.810 45.300 46.980 45.470 ;
        RECT 48.810 45.520 48.980 45.690 ;
        RECT 49.560 45.520 49.730 45.690 ;
        RECT 51.560 45.530 51.730 45.700 ;
        RECT 52.940 46.120 53.110 46.290 ;
        RECT 52.940 45.760 53.110 45.930 ;
        RECT 62.520 45.900 62.690 46.070 ;
        RECT 45.770 44.960 45.940 45.130 ;
        RECT 62.530 45.180 62.700 45.350 ;
        RECT 68.310 45.900 68.480 46.070 ;
        RECT 78.440 47.610 78.610 47.780 ;
        RECT 80.930 47.800 81.100 47.970 ;
        RECT 107.280 48.050 107.450 48.220 ;
        RECT 109.960 48.350 110.130 48.520 ;
        RECT 111.530 48.350 111.700 48.520 ;
        RECT 111.020 48.130 111.190 48.300 ;
        RECT 111.870 47.990 112.040 48.160 ;
        RECT 112.150 48.140 112.320 48.310 ;
        RECT 112.950 48.230 113.120 48.400 ;
        RECT 114.080 47.960 114.250 48.130 ;
        RECT 109.110 47.520 109.280 47.690 ;
        RECT 76.030 46.990 76.210 47.180 ;
        RECT 77.320 47.090 77.490 47.260 ;
        RECT 82.720 47.240 82.890 47.410 ;
        RECT 80.930 46.960 81.100 47.130 ;
        RECT 108.600 47.310 108.770 47.480 ;
        RECT 82.060 46.550 82.230 46.720 ;
        RECT 80.980 46.310 81.150 46.480 ;
        RECT 68.410 45.620 68.580 45.790 ;
        RECT 65.890 44.920 66.160 45.190 ;
        RECT 68.310 45.180 68.480 45.350 ;
        RECT 69.550 44.300 69.720 44.470 ;
        RECT 74.720 44.240 74.890 44.410 ;
        RECT 69.550 43.850 69.720 44.020 ;
        RECT 112.610 47.520 112.780 47.690 ;
        RECT 83.280 46.250 83.450 46.420 ;
        RECT 78.050 45.810 78.220 45.980 ;
        RECT 80.980 45.450 81.150 45.620 ;
        RECT 83.270 45.530 83.440 45.700 ;
        RECT 82.060 45.210 82.230 45.380 ;
        RECT 78.580 44.930 78.750 45.100 ;
        RECT 80.930 44.800 81.100 44.970 ;
        RECT 82.720 44.650 82.890 44.820 ;
        RECT 76.030 44.190 76.210 44.380 ;
        RECT 80.930 43.960 81.100 44.130 ;
        RECT 76.390 43.370 76.560 43.540 ;
        RECT 82.060 43.550 82.230 43.720 ;
        RECT 80.980 43.310 81.150 43.480 ;
        RECT 83.190 43.280 83.360 43.450 ;
        RECT 39.520 40.510 39.690 40.680 ;
        RECT 46.810 40.780 46.980 40.950 ;
        RECT 40.990 40.100 41.200 40.310 ;
        RECT 44.730 40.120 44.900 40.290 ;
        RECT 46.810 40.420 46.980 40.590 ;
        RECT 47.950 40.690 48.120 40.860 ;
        RECT 48.790 40.570 48.960 40.740 ;
        RECT 49.540 40.570 49.710 40.740 ;
        RECT 45.770 40.080 45.940 40.250 ;
        RECT 52.520 40.240 52.690 40.410 ;
        RECT 48.130 39.860 48.300 40.030 ;
        RECT 52.920 40.690 53.090 40.860 ;
        RECT 52.920 40.330 53.090 40.500 ;
        RECT 57.660 40.510 57.830 40.680 ;
        RECT 73.150 40.510 73.320 40.680 ;
        RECT 55.850 40.250 56.020 40.420 ;
        RECT 56.580 40.220 56.750 40.390 ;
        RECT 74.230 40.220 74.400 40.390 ;
        RECT 57.660 39.960 57.830 40.130 ;
        RECT 73.150 39.960 73.320 40.130 ;
        RECT 74.960 40.250 75.130 40.420 ;
        RECT 58.570 39.560 58.740 39.730 ;
        RECT 39.520 38.760 39.690 38.930 ;
        RECT 46.810 39.030 46.980 39.200 ;
        RECT 40.990 38.350 41.200 38.560 ;
        RECT 44.730 38.370 44.900 38.540 ;
        RECT 46.810 38.670 46.980 38.840 ;
        RECT 48.130 38.960 48.300 39.130 ;
        RECT 52.520 38.580 52.690 38.750 ;
        RECT 45.770 38.330 45.940 38.500 ;
        RECT 48.790 38.250 48.960 38.420 ;
        RECT 49.540 38.250 49.710 38.420 ;
        RECT 51.540 38.260 51.710 38.430 ;
        RECT 52.920 38.850 53.090 39.020 ;
        RECT 55.850 38.690 56.020 38.860 ;
        RECT 62.510 39.570 62.680 39.740 ;
        RECT 68.300 39.570 68.470 39.740 ;
        RECT 72.240 39.560 72.410 39.730 ;
        RECT 57.660 38.980 57.830 39.150 ;
        RECT 73.150 38.980 73.320 39.150 ;
        RECT 56.580 38.720 56.750 38.890 ;
        RECT 74.230 38.720 74.400 38.890 ;
        RECT 74.960 38.690 75.130 38.860 ;
        RECT 52.920 38.490 53.090 38.660 ;
        RECT 57.660 38.430 57.830 38.600 ;
        RECT 58.570 37.970 58.740 38.140 ;
        RECT 62.500 38.110 62.670 38.280 ;
        RECT 73.150 38.430 73.320 38.600 ;
        RECT 39.520 37.010 39.690 37.180 ;
        RECT 47.950 37.490 48.120 37.660 ;
        RECT 46.810 37.280 46.980 37.450 ;
        RECT 40.990 36.600 41.200 36.810 ;
        RECT 44.730 36.620 44.900 36.790 ;
        RECT 48.790 37.370 48.960 37.540 ;
        RECT 49.540 37.370 49.710 37.540 ;
        RECT 46.810 36.920 46.980 37.090 ;
        RECT 52.520 37.040 52.690 37.210 ;
        RECT 45.770 36.580 45.940 36.750 ;
        RECT 48.130 36.660 48.300 36.830 ;
        RECT 52.920 37.490 53.090 37.660 ;
        RECT 58.570 37.610 58.740 37.780 ;
        RECT 60.780 37.720 61.050 37.990 ;
        RECT 62.500 37.750 62.670 37.920 ;
        RECT 52.920 37.130 53.090 37.300 ;
        RECT 57.660 37.270 57.830 37.440 ;
        RECT 64.810 37.790 65.080 38.060 ;
        RECT 65.900 37.790 66.170 38.060 ;
        RECT 68.310 38.110 68.480 38.280 ;
        RECT 68.310 37.750 68.480 37.920 ;
        RECT 69.930 37.720 70.200 37.990 ;
        RECT 72.240 37.970 72.410 38.140 ;
        RECT 74.600 37.850 74.780 38.020 ;
        RECT 72.240 37.610 72.410 37.780 ;
        RECT 73.150 37.270 73.320 37.440 ;
        RECT 55.850 37.010 56.020 37.180 ;
        RECT 56.580 36.980 56.750 37.150 ;
        RECT 74.230 36.980 74.400 37.150 ;
        RECT 57.660 36.720 57.830 36.890 ;
        RECT 73.150 36.720 73.320 36.890 ;
        RECT 74.960 37.010 75.130 37.180 ;
        RECT 39.520 35.260 39.690 35.430 ;
        RECT 46.810 35.530 46.980 35.700 ;
        RECT 48.130 35.760 48.300 35.930 ;
        RECT 40.990 34.850 41.200 35.060 ;
        RECT 44.730 34.870 44.900 35.040 ;
        RECT 52.520 35.380 52.690 35.550 ;
        RECT 46.810 35.170 46.980 35.340 ;
        RECT 45.770 34.830 45.940 35.000 ;
        RECT 48.790 35.050 48.960 35.220 ;
        RECT 49.540 35.050 49.710 35.220 ;
        RECT 51.540 35.060 51.710 35.230 ;
        RECT 52.920 35.650 53.090 35.820 ;
        RECT 52.920 35.290 53.090 35.460 ;
        RECT 55.850 35.460 56.020 35.630 ;
        RECT 57.660 35.750 57.830 35.920 ;
        RECT 73.150 35.750 73.320 35.920 ;
        RECT 56.580 35.490 56.750 35.660 ;
        RECT 74.230 35.490 74.400 35.660 ;
        RECT 74.960 35.460 75.130 35.630 ;
        RECT 55.050 35.180 55.220 35.350 ;
        RECT 53.240 34.920 53.410 35.090 ;
        RECT 57.660 35.200 57.830 35.370 ;
        RECT 73.150 35.200 73.320 35.370 ;
        RECT 53.970 34.890 54.140 35.060 ;
        RECT 55.050 34.630 55.220 34.800 ;
        RECT 56.090 34.170 56.260 34.340 ;
        RECT 53.240 33.380 53.410 33.550 ;
        RECT 55.050 33.670 55.220 33.840 ;
        RECT 60.110 34.200 60.280 34.370 ;
        RECT 53.970 33.410 54.140 33.580 ;
        RECT 55.050 33.120 55.220 33.290 ;
        RECT 56.080 32.970 56.250 33.140 ;
        RECT 60.100 32.910 60.270 33.080 ;
        RECT 56.080 32.310 56.250 32.480 ;
        RECT 39.480 31.450 39.650 31.620 ;
        RECT 46.770 31.720 46.940 31.890 ;
        RECT 55.050 31.940 55.220 32.110 ;
        RECT 58.170 32.350 58.440 32.620 ;
        RECT 60.100 32.270 60.270 32.440 ;
        RECT 62.200 32.420 62.470 32.690 ;
        RECT 40.950 31.040 41.160 31.250 ;
        RECT 44.690 31.060 44.860 31.230 ;
        RECT 53.240 31.680 53.410 31.850 ;
        RECT 46.770 31.360 46.940 31.530 ;
        RECT 47.980 31.420 48.150 31.590 ;
        RECT 45.730 31.020 45.900 31.190 ;
        RECT 48.820 31.300 48.990 31.470 ;
        RECT 49.570 31.300 49.740 31.470 ;
        RECT 52.550 30.970 52.720 31.140 ;
        RECT 20.510 30.600 20.680 30.770 ;
        RECT 21.160 30.600 21.330 30.770 ;
        RECT 19.290 30.160 19.460 30.330 ;
        RECT 19.990 30.160 20.160 30.330 ;
        RECT 48.160 30.590 48.330 30.760 ;
        RECT 52.950 31.420 53.120 31.590 ;
        RECT 53.970 31.650 54.140 31.820 ;
        RECT 55.050 31.390 55.220 31.560 ;
        RECT 52.950 31.060 53.120 31.230 ;
        RECT 66.370 30.890 66.540 31.060 ;
        RECT 21.670 29.780 21.840 29.950 ;
        RECT 39.480 29.700 39.650 29.870 ;
        RECT 46.770 29.970 46.940 30.140 ;
        RECT 53.240 30.130 53.410 30.300 ;
        RECT 55.050 30.420 55.220 30.590 ;
        RECT 53.970 30.160 54.140 30.330 ;
        RECT 66.520 30.210 66.690 30.380 ;
        RECT 68.670 30.330 68.840 30.500 ;
        RECT 40.950 29.290 41.160 29.500 ;
        RECT 44.690 29.310 44.860 29.480 ;
        RECT 46.770 29.610 46.940 29.780 ;
        RECT 45.730 29.270 45.900 29.440 ;
        RECT 48.160 29.690 48.330 29.860 ;
        RECT 55.050 29.870 55.220 30.040 ;
        RECT 67.410 29.760 67.580 29.930 ;
        RECT 52.550 29.310 52.720 29.480 ;
        RECT 48.820 28.980 48.990 29.150 ;
        RECT 49.570 28.980 49.740 29.150 ;
        RECT 51.570 28.990 51.740 29.160 ;
        RECT 52.950 29.580 53.120 29.750 ;
        RECT 52.950 29.220 53.120 29.390 ;
        RECT 66.520 29.310 66.690 29.480 ;
        RECT 68.670 29.190 68.840 29.360 ;
        RECT 66.370 28.630 66.540 28.800 ;
        RECT 18.750 28.240 18.920 28.410 ;
        RECT 21.840 28.300 22.010 28.470 ;
        RECT 39.480 27.950 39.650 28.120 ;
        RECT 46.770 28.220 46.940 28.390 ;
        RECT 19.320 26.280 19.490 26.450 ;
        RECT 20.010 26.270 20.180 26.440 ;
        RECT 17.360 26.050 17.530 26.220 ;
        RECT 14.050 25.610 14.220 25.780 ;
        RECT 15.150 25.620 15.320 25.790 ;
        RECT 16.240 25.620 16.410 25.790 ;
        RECT 17.370 25.580 17.540 25.750 ;
        RECT 14.600 24.940 14.770 25.110 ;
        RECT 14.600 23.570 14.770 23.740 ;
        RECT 20.490 25.500 20.660 25.670 ;
        RECT 21.850 27.760 22.020 27.930 ;
        RECT 40.950 27.540 41.160 27.750 ;
        RECT 44.690 27.560 44.860 27.730 ;
        RECT 46.770 27.860 46.940 28.030 ;
        RECT 47.980 28.220 48.150 28.390 ;
        RECT 48.820 28.100 48.990 28.270 ;
        RECT 49.570 28.100 49.740 28.270 ;
        RECT 45.730 27.520 45.900 27.690 ;
        RECT 52.550 27.770 52.720 27.940 ;
        RECT 48.160 27.390 48.330 27.560 ;
        RECT 52.950 28.220 53.120 28.390 ;
        RECT 66.370 28.120 66.540 28.290 ;
        RECT 52.950 27.860 53.120 28.030 ;
        RECT 66.520 27.440 66.690 27.610 ;
        RECT 68.670 27.560 68.840 27.730 ;
        RECT 21.660 26.800 21.830 26.970 ;
        RECT 67.410 26.990 67.580 27.160 ;
        RECT 39.480 26.200 39.650 26.370 ;
        RECT 46.770 26.470 46.940 26.640 ;
        RECT 40.950 25.790 41.160 26.000 ;
        RECT 44.690 25.810 44.860 25.980 ;
        RECT 48.160 26.490 48.330 26.660 ;
        RECT 46.770 26.110 46.940 26.280 ;
        RECT 52.550 26.110 52.720 26.280 ;
        RECT 45.730 25.770 45.900 25.940 ;
        RECT 48.820 25.780 48.990 25.950 ;
        RECT 49.570 25.780 49.740 25.950 ;
        RECT 51.570 25.790 51.740 25.960 ;
        RECT 52.950 26.380 53.120 26.550 ;
        RECT 54.930 26.480 55.100 26.650 ;
        RECT 66.520 26.540 66.690 26.710 ;
        RECT 52.950 26.020 53.120 26.190 ;
        RECT 68.670 26.420 68.840 26.590 ;
        RECT 66.370 25.860 66.540 26.030 ;
        RECT 21.200 25.440 21.370 25.610 ;
        RECT 54.980 25.520 55.150 25.690 ;
        RECT 15.700 24.940 15.870 25.110 ;
        RECT 16.800 24.940 16.970 25.110 ;
        RECT 17.490 24.920 17.660 25.090 ;
        RECT 17.490 24.230 17.660 24.400 ;
        RECT 15.700 23.570 15.870 23.740 ;
        RECT 16.800 23.570 16.970 23.740 ;
        RECT 47.640 23.520 47.810 23.690 ;
        RECT 14.050 22.840 14.220 23.010 ;
        RECT 15.150 22.840 15.320 23.010 ;
        RECT 16.240 22.840 16.410 23.010 ;
        RECT 14.040 21.500 14.210 21.670 ;
        RECT 15.150 21.490 15.320 21.660 ;
        RECT 16.240 21.470 16.410 21.640 ;
        RECT 24.040 21.670 24.210 22.010 ;
        RECT 24.410 21.670 24.580 22.010 ;
        RECT 14.600 20.800 14.770 20.970 ;
        RECT 15.700 20.790 15.870 20.960 ;
        RECT 16.790 20.790 16.960 20.960 ;
        RECT 48.730 23.520 48.900 23.690 ;
        RECT 48.190 22.840 48.360 23.010 ;
        RECT 48.190 21.470 48.360 21.640 ;
        RECT 47.630 20.740 47.800 20.910 ;
        RECT 47.630 19.370 47.800 19.540 ;
        RECT 47.060 18.730 47.230 18.900 ;
        RECT 49.830 23.510 50.000 23.680 ;
        RECT 49.280 22.820 49.450 22.990 ;
        RECT 49.280 21.470 49.450 21.640 ;
        RECT 48.730 20.740 48.900 20.910 ;
        RECT 48.730 19.370 48.900 19.540 ;
        RECT 48.190 18.690 48.360 18.860 ;
        RECT 50.950 23.690 51.120 23.860 ;
        RECT 50.950 23.330 51.120 23.500 ;
        RECT 51.560 23.690 51.730 23.860 ;
        RECT 51.560 23.330 51.730 23.500 ;
        RECT 52.680 23.510 52.850 23.680 ;
        RECT 50.390 22.810 50.560 22.980 ;
        RECT 52.120 22.810 52.290 22.980 ;
        RECT 50.380 21.470 50.550 21.640 ;
        RECT 52.130 21.470 52.300 21.640 ;
        RECT 49.830 20.740 50.000 20.910 ;
        RECT 49.830 19.370 50.000 19.540 ;
        RECT 49.280 18.690 49.450 18.860 ;
        RECT 53.780 23.520 53.950 23.690 ;
        RECT 53.230 22.820 53.400 22.990 ;
        RECT 53.230 21.470 53.400 21.640 ;
        RECT 52.680 20.740 52.850 20.910 ;
        RECT 52.680 19.370 52.850 19.540 ;
        RECT 50.380 18.700 50.550 18.870 ;
        RECT 52.130 18.700 52.300 18.870 ;
        RECT 54.870 23.520 55.040 23.690 ;
        RECT 57.450 23.550 57.620 23.720 ;
        RECT 54.320 22.840 54.490 23.010 ;
        RECT 54.320 21.470 54.490 21.640 ;
        RECT 53.780 20.740 53.950 20.910 ;
        RECT 53.780 19.370 53.950 19.540 ;
        RECT 53.230 18.690 53.400 18.860 ;
        RECT 58.540 23.550 58.710 23.720 ;
        RECT 58.000 22.870 58.170 23.040 ;
        RECT 58.000 21.500 58.170 21.670 ;
        RECT 54.880 20.740 55.050 20.910 ;
        RECT 57.440 20.770 57.610 20.940 ;
        RECT 54.880 19.370 55.050 19.540 ;
        RECT 57.440 19.400 57.610 19.570 ;
        RECT 54.320 18.690 54.490 18.860 ;
        RECT 55.450 18.730 55.620 18.900 ;
        RECT 47.070 18.260 47.240 18.430 ;
        RECT 55.440 18.260 55.610 18.430 ;
        RECT 56.870 18.760 57.040 18.930 ;
        RECT 59.640 23.540 59.810 23.710 ;
        RECT 59.090 22.850 59.260 23.020 ;
        RECT 59.090 21.500 59.260 21.670 ;
        RECT 58.540 20.770 58.710 20.940 ;
        RECT 58.540 19.400 58.710 19.570 ;
        RECT 58.000 18.720 58.170 18.890 ;
        RECT 60.760 23.720 60.930 23.890 ;
        RECT 60.760 23.360 60.930 23.530 ;
        RECT 61.370 23.720 61.540 23.890 ;
        RECT 61.370 23.360 61.540 23.530 ;
        RECT 62.490 23.540 62.660 23.710 ;
        RECT 60.200 22.840 60.370 23.010 ;
        RECT 61.930 22.840 62.100 23.010 ;
        RECT 60.190 21.500 60.360 21.670 ;
        RECT 61.940 21.500 62.110 21.670 ;
        RECT 59.640 20.770 59.810 20.940 ;
        RECT 59.640 19.400 59.810 19.570 ;
        RECT 59.090 18.720 59.260 18.890 ;
        RECT 63.590 23.550 63.760 23.720 ;
        RECT 63.040 22.850 63.210 23.020 ;
        RECT 63.040 21.500 63.210 21.670 ;
        RECT 62.490 20.770 62.660 20.940 ;
        RECT 62.490 19.400 62.660 19.570 ;
        RECT 60.190 18.730 60.360 18.900 ;
        RECT 61.940 18.730 62.110 18.900 ;
        RECT 64.680 23.550 64.850 23.720 ;
        RECT 64.130 22.870 64.300 23.040 ;
        RECT 64.130 21.500 64.300 21.670 ;
        RECT 63.590 20.770 63.760 20.940 ;
        RECT 63.590 19.400 63.760 19.570 ;
        RECT 63.040 18.720 63.210 18.890 ;
        RECT 64.690 20.770 64.860 20.940 ;
        RECT 64.690 19.400 64.860 19.570 ;
        RECT 64.130 18.720 64.300 18.890 ;
        RECT 65.260 18.760 65.430 18.930 ;
        RECT 56.880 18.290 57.050 18.460 ;
        RECT 65.250 18.290 65.420 18.460 ;
        RECT 68.870 19.330 69.040 19.500 ;
        RECT 68.310 18.630 68.480 18.800 ;
        RECT 69.970 19.340 70.140 19.510 ;
        RECT 71.060 19.340 71.230 19.510 ;
        RECT 69.420 18.640 69.590 18.810 ;
        RECT 70.510 18.660 70.680 18.830 ;
        RECT 68.320 17.290 68.490 17.460 ;
        RECT 69.420 17.290 69.590 17.460 ;
        RECT 70.510 17.290 70.680 17.460 ;
        RECT 68.870 16.560 69.040 16.730 ;
        RECT 68.870 15.190 69.040 15.360 ;
        RECT 69.970 16.560 70.140 16.730 ;
        RECT 71.070 16.560 71.240 16.730 ;
        RECT 71.760 16.260 71.930 16.430 ;
        RECT 71.760 15.900 71.930 16.070 ;
        RECT 69.970 15.190 70.140 15.360 ;
        RECT 71.070 15.190 71.240 15.360 ;
        RECT 102.320 15.850 102.490 16.020 ;
        RECT 107.760 15.010 107.930 15.180 ;
        RECT 68.320 14.520 68.490 14.690 ;
        RECT 69.420 14.510 69.590 14.680 ;
        RECT 70.510 14.510 70.680 14.680 ;
        RECT 71.640 14.550 71.810 14.720 ;
        RECT 16.760 14.300 16.930 14.470 ;
        RECT 13.450 13.860 13.620 14.030 ;
        RECT 14.550 13.870 14.720 14.040 ;
        RECT 14.000 13.190 14.170 13.360 ;
        RECT 14.000 11.820 14.170 11.990 ;
        RECT 13.450 11.090 13.620 11.260 ;
        RECT 13.440 9.750 13.610 9.920 ;
        RECT 12.880 9.230 13.050 9.400 ;
        RECT 15.640 13.870 15.810 14.040 ;
        RECT 15.100 13.190 15.270 13.360 ;
        RECT 15.100 11.820 15.270 11.990 ;
        RECT 14.550 11.090 14.720 11.260 ;
        RECT 14.550 9.740 14.720 9.910 ;
        RECT 14.000 9.050 14.170 9.220 ;
        RECT 71.630 14.080 71.800 14.250 ;
        RECT 102.320 14.240 102.490 14.410 ;
        RECT 107.760 14.340 107.930 14.510 ;
        RECT 16.770 13.830 16.940 14.000 ;
        RECT 16.200 13.190 16.370 13.360 ;
        RECT 16.200 11.820 16.370 11.990 ;
        RECT 15.640 11.090 15.810 11.260 ;
        RECT 15.640 9.720 15.810 9.890 ;
        RECT 15.100 9.040 15.270 9.210 ;
        RECT 18.230 9.700 18.400 13.220 ;
        RECT 18.590 9.700 18.760 13.220 ;
        RECT 18.950 9.700 19.120 13.220 ;
        RECT 19.640 9.700 19.810 13.220 ;
        RECT 20.000 9.700 20.170 13.220 ;
        RECT 20.360 9.700 20.530 13.220 ;
        RECT 102.320 12.640 102.490 12.810 ;
        RECT 102.320 11.020 102.490 11.190 ;
        RECT 104.510 9.850 104.680 10.020 ;
        RECT 102.320 9.420 102.490 9.590 ;
        RECT 16.190 9.040 16.360 9.210 ;
        RECT 102.320 7.800 102.490 7.970 ;
        RECT 102.320 6.200 102.490 6.370 ;
        RECT 102.320 4.580 102.490 4.750 ;
        RECT 108.600 2.490 108.770 17.440 ;
      LAYER met1 ;
        RECT 80.150 74.040 80.490 74.180 ;
        RECT 88.030 74.040 88.750 75.780 ;
        RECT 80.150 73.320 88.750 74.040 ;
        RECT 28.080 70.870 29.420 71.320 ;
        RECT 1.980 70.030 2.480 70.510 ;
        RECT 28.080 70.450 41.600 70.870 ;
        RECT 43.390 70.780 46.580 71.900 ;
        RECT 28.080 70.310 29.420 70.450 ;
        RECT 2.080 67.070 2.470 70.030 ;
        RECT 22.670 69.710 25.440 69.950 ;
        RECT 22.670 69.300 22.910 69.710 ;
        RECT 2.080 66.580 2.550 67.070 ;
        RECT 2.080 66.570 2.530 66.580 ;
        RECT 8.340 66.570 8.580 67.210 ;
        RECT 13.550 66.650 13.790 67.060 ;
        RECT 0.180 61.010 0.470 62.070 ;
        RECT 2.080 8.460 2.470 66.570 ;
        RECT 8.340 66.310 8.570 66.570 ;
        RECT 8.330 66.090 8.570 66.310 ;
        RECT 19.390 65.810 19.660 67.060 ;
        RECT 24.100 65.770 24.360 67.060 ;
        RECT 3.490 65.430 3.750 65.750 ;
        RECT 3.500 63.210 3.740 65.430 ;
        RECT 11.400 64.740 11.720 65.060 ;
        RECT 12.760 64.820 13.080 65.140 ;
        RECT 13.450 64.810 13.770 65.130 ;
        RECT 8.340 63.770 8.580 64.410 ;
        RECT 8.340 63.510 8.570 63.770 ;
        RECT 8.330 63.290 8.570 63.510 ;
        RECT 3.410 62.730 3.830 63.210 ;
        RECT 8.340 62.220 8.580 62.860 ;
        RECT 8.340 61.960 8.570 62.220 ;
        RECT 9.300 61.970 9.590 63.890 ;
        RECT 19.400 63.600 19.660 63.620 ;
        RECT 8.330 61.740 8.570 61.960 ;
        RECT 9.280 61.300 9.690 61.970 ;
        RECT 10.680 61.080 11.000 61.400 ;
        RECT 13.540 61.010 13.780 62.890 ;
        RECT 19.360 61.010 19.670 63.600 ;
        RECT 20.540 61.100 20.860 61.420 ;
        RECT 22.660 60.610 22.900 63.840 ;
        RECT 23.330 63.060 23.560 63.230 ;
        RECT 23.320 61.190 23.570 63.060 ;
        RECT 23.320 61.010 23.580 61.190 ;
        RECT 22.610 60.270 22.950 60.610 ;
        RECT 19.860 60.170 20.350 60.180 ;
        RECT 15.930 51.480 16.160 54.960 ;
        RECT 16.600 54.340 16.820 54.960 ;
        RECT 17.700 54.530 18.020 54.850 ;
        RECT 18.790 54.540 19.110 54.860 ;
        RECT 16.570 54.020 16.830 54.340 ;
        RECT 17.270 54.030 17.590 54.350 ;
        RECT 16.600 53.420 16.820 54.020 ;
        RECT 17.710 53.540 18.030 53.860 ;
        RECT 18.800 53.550 19.120 53.870 ;
        RECT 16.540 53.100 16.820 53.420 ;
        RECT 17.250 53.110 17.570 53.430 ;
        RECT 16.600 52.500 16.820 53.100 ;
        RECT 17.710 52.550 18.030 52.870 ;
        RECT 18.800 52.560 19.120 52.880 ;
        RECT 16.550 52.180 16.820 52.500 ;
        RECT 15.900 51.160 16.160 51.480 ;
        RECT 15.930 50.520 16.160 51.160 ;
        RECT 15.860 50.200 16.160 50.520 ;
        RECT 15.930 49.560 16.160 50.200 ;
        RECT 15.900 49.240 16.160 49.560 ;
        RECT 15.930 34.490 16.160 49.240 ;
        RECT 16.600 34.490 16.820 52.180 ;
        RECT 17.230 52.120 17.550 52.440 ;
        RECT 18.730 52.170 19.050 52.490 ;
        RECT 18.700 51.990 19.020 52.030 ;
        RECT 18.470 51.760 19.020 51.990 ;
        RECT 18.700 51.710 19.020 51.760 ;
        RECT 18.730 51.180 19.050 51.500 ;
        RECT 18.700 51.000 19.020 51.040 ;
        RECT 18.470 50.770 19.020 51.000 ;
        RECT 18.700 50.720 19.020 50.770 ;
        RECT 18.730 50.190 19.050 50.510 ;
        RECT 19.290 50.290 19.510 59.230 ;
        RECT 19.850 59.020 20.360 60.170 ;
        RECT 25.200 59.240 25.440 69.710 ;
        RECT 28.510 69.380 31.540 69.650 ;
        RECT 33.220 69.390 33.480 70.450 ;
        RECT 28.480 60.210 28.790 63.910 ;
        RECT 28.400 59.840 28.790 60.210 ;
        RECT 31.270 59.700 31.540 69.380 ;
        RECT 41.180 67.200 41.600 70.450 ;
        RECT 44.990 67.960 45.410 70.780 ;
        RECT 71.980 70.770 75.170 71.890 ;
        RECT 44.990 67.480 45.460 67.960 ;
        RECT 41.140 66.720 41.620 67.200 ;
        RECT 64.750 66.700 66.220 67.230 ;
        RECT 46.690 65.110 47.130 65.610 ;
        RECT 52.410 65.110 52.850 65.610 ;
        RECT 42.270 64.090 42.710 64.590 ;
        RECT 32.440 60.700 32.690 63.850 ;
        RECT 39.480 61.350 39.800 61.400 ;
        RECT 39.390 61.060 39.800 61.350 ;
        RECT 32.400 60.340 32.730 60.700 ;
        RECT 31.230 59.390 31.570 59.700 ;
        RECT 19.800 58.920 20.360 59.020 ;
        RECT 25.150 58.920 25.490 59.240 ;
        RECT 19.270 50.220 19.510 50.290 ;
        RECT 19.690 58.520 20.360 58.920 ;
        RECT 39.390 58.630 39.630 61.060 ;
        RECT 42.330 58.630 42.640 64.090 ;
        RECT 19.690 58.490 20.350 58.520 ;
        RECT 19.690 54.350 19.910 58.490 ;
        RECT 39.390 57.560 39.730 58.630 ;
        RECT 40.910 57.920 41.260 58.210 ;
        RECT 40.910 57.900 41.110 57.920 ;
        RECT 38.750 57.060 39.160 57.390 ;
        RECT 20.910 56.370 21.260 56.830 ;
        RECT 37.340 56.390 37.710 56.700 ;
        RECT 20.310 56.010 20.560 56.130 ;
        RECT 20.280 55.550 20.600 56.010 ;
        RECT 20.310 54.760 20.560 55.550 ;
        RECT 20.310 54.440 20.600 54.760 ;
        RECT 19.690 54.060 20.010 54.350 ;
        RECT 19.270 50.120 19.610 50.220 ;
        RECT 18.700 50.010 19.020 50.050 ;
        RECT 18.470 49.780 19.020 50.010 ;
        RECT 18.700 49.730 19.020 49.780 ;
        RECT 19.290 49.990 19.610 50.120 ;
        RECT 15.820 33.960 16.160 34.490 ;
        RECT 16.480 33.960 16.820 34.490 ;
        RECT 14.510 33.220 14.740 33.290 ;
        RECT 14.470 32.960 14.790 33.220 ;
        RECT 14.020 32.850 14.250 32.890 ;
        RECT 13.980 32.530 14.250 32.850 ;
        RECT 4.670 31.290 5.390 31.990 ;
        RECT 4.680 26.140 5.340 31.290 ;
        RECT 14.020 29.010 14.250 32.530 ;
        RECT 14.510 30.490 14.740 32.960 ;
        RECT 15.930 32.870 16.160 33.960 ;
        RECT 16.600 33.230 16.820 33.960 ;
        RECT 18.360 33.250 18.630 33.290 ;
        RECT 16.580 32.910 16.840 33.230 ;
        RECT 18.340 32.920 18.630 33.250 ;
        RECT 15.920 32.550 16.180 32.870 ;
        RECT 17.810 31.380 18.100 31.410 ;
        RECT 14.510 30.120 15.240 30.490 ;
        RECT 14.020 28.940 14.280 29.010 ;
        RECT 14.000 28.930 14.280 28.940 ;
        RECT 13.970 28.620 14.290 28.930 ;
        RECT 9.870 26.760 10.300 27.190 ;
        RECT 4.680 25.420 5.420 26.140 ;
        RECT 9.920 20.950 10.290 26.760 ;
        RECT 13.970 25.530 14.290 25.850 ;
        RECT 14.510 25.180 14.740 30.120 ;
        RECT 18.360 29.950 18.630 32.920 ;
        RECT 18.240 29.700 18.630 29.950 ;
        RECT 18.840 32.850 19.080 32.890 ;
        RECT 18.840 32.530 19.100 32.850 ;
        RECT 18.840 29.390 19.080 32.530 ;
        RECT 19.290 30.400 19.510 49.990 ;
        RECT 19.690 31.100 19.910 54.060 ;
        RECT 20.310 53.840 20.560 54.440 ;
        RECT 20.310 53.520 20.600 53.840 ;
        RECT 20.310 52.920 20.560 53.520 ;
        RECT 20.310 52.600 20.570 52.920 ;
        RECT 20.310 52.390 20.560 52.600 ;
        RECT 20.030 52.070 20.560 52.390 ;
        RECT 20.310 51.400 20.560 52.070 ;
        RECT 20.030 51.080 20.560 51.400 ;
        RECT 20.310 50.410 20.560 51.080 ;
        RECT 20.030 50.090 20.560 50.410 ;
        RECT 20.310 32.250 20.560 50.090 ;
        RECT 20.930 51.830 21.190 56.370 ;
        RECT 36.700 54.670 37.090 55.040 ;
        RECT 36.120 53.180 36.510 53.570 ;
        RECT 20.930 51.510 21.210 51.830 ;
        RECT 35.480 51.590 35.870 51.970 ;
        RECT 35.510 51.580 35.850 51.590 ;
        RECT 20.930 50.870 21.190 51.510 ;
        RECT 34.870 51.390 35.210 51.400 ;
        RECT 34.860 51.000 35.220 51.390 ;
        RECT 20.930 50.550 21.220 50.870 ;
        RECT 20.930 49.910 21.190 50.550 ;
        RECT 20.930 49.590 21.210 49.910 ;
        RECT 20.310 32.230 20.570 32.250 ;
        RECT 20.300 31.950 20.580 32.230 ;
        RECT 20.310 31.930 20.570 31.950 ;
        RECT 19.650 30.780 19.970 31.100 ;
        RECT 20.310 30.840 20.560 31.930 ;
        RECT 20.930 30.840 21.190 49.590 ;
        RECT 34.250 49.440 34.610 49.830 ;
        RECT 33.600 47.900 34.010 48.300 ;
        RECT 33.070 46.340 33.430 46.730 ;
        RECT 32.490 41.280 32.820 41.300 ;
        RECT 32.430 40.860 32.820 41.280 ;
        RECT 31.860 39.670 32.190 39.690 ;
        RECT 31.810 39.280 32.200 39.670 ;
        RECT 31.240 38.120 31.570 38.130 ;
        RECT 31.210 37.730 31.570 38.120 ;
        RECT 30.590 36.250 30.980 36.650 ;
        RECT 29.920 31.080 30.350 31.480 ;
        RECT 19.220 30.080 19.540 30.400 ;
        RECT 18.240 29.160 19.080 29.390 ;
        RECT 18.840 29.050 19.080 29.160 ;
        RECT 18.800 28.730 19.080 29.050 ;
        RECT 18.840 28.470 19.080 28.730 ;
        RECT 19.290 28.490 19.510 30.080 ;
        RECT 18.720 28.270 19.080 28.470 ;
        RECT 18.720 27.960 19.140 28.270 ;
        RECT 19.250 28.170 19.530 28.490 ;
        RECT 18.840 27.760 19.140 27.960 ;
        RECT 18.840 27.500 19.080 27.760 ;
        RECT 18.800 27.180 19.080 27.500 ;
        RECT 17.280 25.970 17.600 26.290 ;
        RECT 15.070 25.540 15.390 25.860 ;
        RECT 16.160 25.540 16.480 25.860 ;
        RECT 17.290 25.500 17.610 25.820 ;
        RECT 14.510 24.860 14.840 25.180 ;
        RECT 15.620 24.860 15.940 25.180 ;
        RECT 16.720 24.860 17.040 25.180 ;
        RECT 14.510 23.810 14.740 24.860 ;
        RECT 17.430 24.690 17.720 25.120 ;
        RECT 17.430 24.670 17.900 24.690 ;
        RECT 17.440 24.370 17.900 24.670 ;
        RECT 17.440 23.840 17.720 24.370 ;
        RECT 17.450 23.810 17.720 23.840 ;
        RECT 14.510 23.490 14.840 23.810 ;
        RECT 15.620 23.490 15.940 23.810 ;
        RECT 16.720 23.490 17.040 23.810 ;
        RECT 13.970 22.760 14.290 23.080 ;
        RECT 14.510 22.620 14.740 23.490 ;
        RECT 15.070 22.760 15.390 23.080 ;
        RECT 16.160 22.760 16.480 23.080 ;
        RECT 14.510 22.390 16.960 22.620 ;
        RECT 16.640 22.060 16.960 22.390 ;
        RECT 13.960 21.420 14.280 21.740 ;
        RECT 15.070 21.410 15.390 21.730 ;
        RECT 16.160 21.390 16.480 21.710 ;
        RECT 9.880 20.520 10.310 20.950 ;
        RECT 14.520 20.720 14.840 21.040 ;
        RECT 15.620 20.710 15.940 21.030 ;
        RECT 16.710 20.710 17.030 21.030 ;
        RECT 17.400 20.490 17.730 20.520 ;
        RECT 17.260 20.410 17.730 20.490 ;
        RECT 17.020 20.170 17.730 20.410 ;
        RECT 17.400 20.100 17.730 20.170 ;
        RECT 12.890 14.860 13.180 15.210 ;
        RECT 12.900 9.570 13.160 14.860 ;
        RECT 16.680 14.220 17.000 14.540 ;
        RECT 18.840 14.500 19.080 27.180 ;
        RECT 19.290 26.520 19.510 28.170 ;
        RECT 19.250 26.200 19.570 26.520 ;
        RECT 19.290 15.200 19.510 26.200 ;
        RECT 19.690 22.960 19.910 30.780 ;
        RECT 20.310 30.520 20.760 30.840 ;
        RECT 20.930 30.520 21.410 30.840 ;
        RECT 19.920 30.080 20.240 30.400 ;
        RECT 19.940 26.190 20.260 26.510 ;
        RECT 20.310 25.740 20.560 30.520 ;
        RECT 20.930 27.920 21.190 30.520 ;
        RECT 21.610 29.070 21.900 29.980 ;
        RECT 29.260 29.510 29.670 29.910 ;
        RECT 21.520 28.500 21.840 28.540 ;
        RECT 21.520 28.270 22.080 28.500 ;
        RECT 21.520 28.220 21.840 28.270 ;
        RECT 21.530 27.960 21.850 28.000 ;
        RECT 20.920 27.600 21.230 27.920 ;
        RECT 21.530 27.730 22.080 27.960 ;
        RECT 28.650 27.870 29.040 28.270 ;
        RECT 21.530 27.680 21.850 27.730 ;
        RECT 20.310 25.420 20.740 25.740 ;
        RECT 20.930 25.680 21.190 27.600 ;
        RECT 21.600 27.050 21.870 27.230 ;
        RECT 21.580 26.730 21.900 27.050 ;
        RECT 21.600 26.560 21.870 26.730 ;
        RECT 27.960 26.430 28.370 26.820 ;
        RECT 19.690 22.480 19.980 22.960 ;
        RECT 19.690 20.520 19.910 22.480 ;
        RECT 19.670 20.100 19.930 20.520 ;
        RECT 19.690 15.480 19.910 20.100 ;
        RECT 20.310 16.860 20.560 25.420 ;
        RECT 20.930 25.360 21.450 25.680 ;
        RECT 20.270 16.460 20.570 16.860 ;
        RECT 19.690 15.340 19.930 15.480 ;
        RECT 19.250 14.850 19.560 15.200 ;
        RECT 19.700 14.710 19.930 15.340 ;
        RECT 13.370 13.780 13.690 14.100 ;
        RECT 14.470 13.790 14.790 14.110 ;
        RECT 15.560 13.790 15.880 14.110 ;
        RECT 16.690 13.750 17.010 14.070 ;
        RECT 18.050 13.940 19.080 14.500 ;
        RECT 19.690 14.680 19.930 14.710 ;
        RECT 18.050 13.830 18.840 13.940 ;
        RECT 13.920 13.110 14.240 13.430 ;
        RECT 15.020 13.110 15.340 13.430 ;
        RECT 16.120 13.110 16.440 13.430 ;
        RECT 19.690 13.290 19.910 14.680 ;
        RECT 13.920 11.740 14.240 12.060 ;
        RECT 15.020 11.740 15.340 12.060 ;
        RECT 16.120 11.740 16.440 12.060 ;
        RECT 13.370 11.010 13.690 11.330 ;
        RECT 14.470 11.010 14.790 11.330 ;
        RECT 15.560 11.010 15.880 11.330 ;
        RECT 13.360 9.670 13.680 9.990 ;
        RECT 14.470 9.660 14.790 9.980 ;
        RECT 15.560 9.640 15.880 9.960 ;
        RECT 18.160 9.610 20.580 13.290 ;
        RECT 12.850 8.760 13.160 9.570 ;
        RECT 20.930 9.320 21.190 25.360 ;
        RECT 23.750 21.280 24.680 22.930 ;
        RECT 23.840 20.800 24.580 21.280 ;
        RECT 13.920 8.970 14.240 9.290 ;
        RECT 15.020 8.960 15.340 9.280 ;
        RECT 16.110 8.960 16.430 9.280 ;
        RECT 20.840 8.910 21.190 9.320 ;
        RECT 12.900 8.560 13.160 8.760 ;
        RECT 1.910 7.940 2.470 8.460 ;
        RECT 28.020 3.090 28.350 26.430 ;
        RECT 27.970 3.080 28.400 3.090 ;
        RECT 27.940 2.620 28.430 3.080 ;
        RECT 27.970 2.600 28.400 2.620 ;
        RECT 28.670 2.300 29.000 27.870 ;
        RECT 28.580 1.810 29.070 2.300 ;
        RECT 29.320 1.590 29.650 29.510 ;
        RECT 29.290 1.130 29.690 1.590 ;
        RECT 29.080 0.640 29.660 0.750 ;
        RECT 29.990 0.640 30.320 31.080 ;
        RECT 30.630 5.220 30.960 36.250 ;
        RECT 30.630 0.760 30.950 5.220 ;
        RECT 31.240 1.370 31.570 37.730 ;
        RECT 31.860 1.620 32.190 39.280 ;
        RECT 32.490 2.650 32.820 40.860 ;
        RECT 33.090 2.950 33.420 46.340 ;
        RECT 33.670 3.520 34.000 47.900 ;
        RECT 34.280 4.550 34.610 49.440 ;
        RECT 34.870 5.160 35.200 51.000 ;
        RECT 35.510 5.830 35.840 51.580 ;
        RECT 36.130 6.480 36.460 53.180 ;
        RECT 36.730 7.110 37.060 54.670 ;
        RECT 37.360 7.720 37.690 56.390 ;
        RECT 38.750 55.310 39.160 55.640 ;
        RECT 38.750 53.560 39.160 53.890 ;
        RECT 38.750 51.810 39.160 52.140 ;
        RECT 38.750 51.010 39.160 51.340 ;
        RECT 38.750 49.260 39.160 49.590 ;
        RECT 38.750 47.510 39.160 47.840 ;
        RECT 38.750 45.760 39.160 46.090 ;
        RECT 39.490 45.480 39.730 57.560 ;
        RECT 42.330 57.490 42.740 58.630 ;
        RECT 44.650 58.200 44.960 58.210 ;
        RECT 44.650 57.930 44.970 58.200 ;
        RECT 45.690 57.970 46.010 58.270 ;
        RECT 44.670 57.920 44.960 57.930 ;
        RECT 40.910 56.170 41.260 56.460 ;
        RECT 40.910 56.150 41.110 56.170 ;
        RECT 40.910 54.420 41.260 54.710 ;
        RECT 40.910 54.400 41.110 54.420 ;
        RECT 40.910 52.670 41.260 52.960 ;
        RECT 40.910 52.650 41.110 52.670 ;
        RECT 40.910 50.480 41.110 50.500 ;
        RECT 40.910 50.190 41.260 50.480 ;
        RECT 40.910 48.730 41.110 48.750 ;
        RECT 40.910 48.440 41.260 48.730 ;
        RECT 40.910 46.980 41.110 47.000 ;
        RECT 40.910 46.690 41.260 46.980 ;
        RECT 42.430 45.550 42.740 57.490 ;
        RECT 42.990 57.170 43.270 57.500 ;
        RECT 44.650 56.450 44.960 56.460 ;
        RECT 44.650 56.180 44.970 56.450 ;
        RECT 45.690 56.220 46.010 56.520 ;
        RECT 44.670 56.170 44.960 56.180 ;
        RECT 42.990 55.420 43.270 55.750 ;
        RECT 44.650 54.700 44.960 54.710 ;
        RECT 44.650 54.430 44.970 54.700 ;
        RECT 45.690 54.470 46.010 54.770 ;
        RECT 44.670 54.420 44.960 54.430 ;
        RECT 42.990 53.670 43.270 54.000 ;
        RECT 44.650 52.950 44.960 52.960 ;
        RECT 44.650 52.680 44.970 52.950 ;
        RECT 45.690 52.720 46.010 53.020 ;
        RECT 44.670 52.670 44.960 52.680 ;
        RECT 42.990 51.920 43.270 52.250 ;
        RECT 42.990 50.900 43.270 51.230 ;
        RECT 44.670 50.470 44.960 50.480 ;
        RECT 44.650 50.200 44.970 50.470 ;
        RECT 44.650 50.190 44.960 50.200 ;
        RECT 45.690 50.130 46.010 50.430 ;
        RECT 42.990 49.150 43.270 49.480 ;
        RECT 44.670 48.720 44.960 48.730 ;
        RECT 44.650 48.450 44.970 48.720 ;
        RECT 44.650 48.440 44.960 48.450 ;
        RECT 45.690 48.380 46.010 48.680 ;
        RECT 42.990 47.400 43.270 47.730 ;
        RECT 44.670 46.970 44.960 46.980 ;
        RECT 44.650 46.700 44.970 46.970 ;
        RECT 44.650 46.690 44.960 46.700 ;
        RECT 45.690 46.630 46.010 46.930 ;
        RECT 42.990 45.650 43.270 45.980 ;
        RECT 39.390 44.520 39.730 45.480 ;
        RECT 40.910 45.230 41.110 45.250 ;
        RECT 40.910 44.940 41.260 45.230 ;
        RECT 42.330 44.520 42.740 45.550 ;
        RECT 44.670 45.220 44.960 45.230 ;
        RECT 44.650 44.950 44.970 45.220 ;
        RECT 44.650 44.940 44.960 44.950 ;
        RECT 45.690 44.880 46.010 45.180 ;
        RECT 39.390 41.390 39.630 44.520 ;
        RECT 42.330 41.390 42.640 44.520 ;
        RECT 38.750 40.880 39.160 41.210 ;
        RECT 39.390 41.110 39.730 41.390 ;
        RECT 38.750 39.130 39.160 39.460 ;
        RECT 38.750 37.380 39.160 37.710 ;
        RECT 38.750 35.630 39.160 35.960 ;
        RECT 39.490 35.350 39.730 41.110 ;
        RECT 42.330 41.040 42.740 41.390 ;
        RECT 40.910 40.350 41.110 40.370 ;
        RECT 40.910 40.060 41.260 40.350 ;
        RECT 40.910 38.600 41.110 38.620 ;
        RECT 40.910 38.310 41.260 38.600 ;
        RECT 40.910 36.850 41.110 36.870 ;
        RECT 40.910 36.560 41.260 36.850 ;
        RECT 42.430 35.420 42.740 41.040 ;
        RECT 42.990 40.770 43.270 41.100 ;
        RECT 44.670 40.340 44.960 40.350 ;
        RECT 44.650 40.070 44.970 40.340 ;
        RECT 44.650 40.060 44.960 40.070 ;
        RECT 45.690 40.000 46.010 40.300 ;
        RECT 42.990 39.020 43.270 39.350 ;
        RECT 44.670 38.590 44.960 38.600 ;
        RECT 44.650 38.320 44.970 38.590 ;
        RECT 44.650 38.310 44.960 38.320 ;
        RECT 45.690 38.250 46.010 38.550 ;
        RECT 42.990 37.270 43.270 37.600 ;
        RECT 44.670 36.840 44.960 36.850 ;
        RECT 44.650 36.570 44.970 36.840 ;
        RECT 44.650 36.560 44.960 36.570 ;
        RECT 45.690 36.500 46.010 36.800 ;
        RECT 42.990 35.520 43.270 35.850 ;
        RECT 38.710 31.820 39.120 32.150 ;
        RECT 39.390 31.580 39.730 35.350 ;
        RECT 40.910 35.100 41.110 35.120 ;
        RECT 40.910 34.810 41.260 35.100 ;
        RECT 42.330 31.580 42.740 35.420 ;
        RECT 44.670 35.090 44.960 35.100 ;
        RECT 44.650 34.820 44.970 35.090 ;
        RECT 44.650 34.810 44.960 34.820 ;
        RECT 45.690 34.750 46.010 35.050 ;
        RECT 46.760 32.330 47.050 65.110 ;
        RECT 47.950 64.120 48.450 64.560 ;
        RECT 48.220 51.390 48.410 64.120 ;
        RECT 50.300 51.930 50.580 52.580 ;
        RECT 47.940 50.900 48.410 51.390 ;
        RECT 48.800 51.250 49.170 51.270 ;
        RECT 48.750 50.990 49.170 51.250 ;
        RECT 48.800 50.980 49.170 50.990 ;
        RECT 47.760 50.460 48.080 50.740 ;
        RECT 48.220 50.560 48.410 50.900 ;
        RECT 48.120 50.270 48.410 50.560 ;
        RECT 48.220 49.660 48.410 50.270 ;
        RECT 47.760 49.190 48.080 49.470 ;
        RECT 48.120 49.370 48.410 49.660 ;
        RECT 48.220 49.030 48.410 49.370 ;
        RECT 47.940 48.540 48.410 49.030 ;
        RECT 48.800 48.940 49.170 48.950 ;
        RECT 48.750 48.680 49.170 48.940 ;
        RECT 48.800 48.660 49.170 48.680 ;
        RECT 48.220 48.190 48.410 48.540 ;
        RECT 47.940 47.700 48.410 48.190 ;
        RECT 48.800 48.050 49.170 48.070 ;
        RECT 48.750 47.790 49.170 48.050 ;
        RECT 48.800 47.780 49.170 47.790 ;
        RECT 47.760 47.260 48.080 47.540 ;
        RECT 48.220 47.360 48.410 47.700 ;
        RECT 48.120 47.070 48.410 47.360 ;
        RECT 48.220 46.460 48.410 47.070 ;
        RECT 47.760 45.990 48.080 46.270 ;
        RECT 48.120 46.170 48.410 46.460 ;
        RECT 48.220 45.830 48.410 46.170 ;
        RECT 47.940 45.340 48.410 45.830 ;
        RECT 48.800 45.740 49.170 45.750 ;
        RECT 48.750 45.480 49.170 45.740 ;
        RECT 48.800 45.460 49.170 45.480 ;
        RECT 48.220 41.570 48.410 45.340 ;
        RECT 49.530 41.670 49.760 51.610 ;
        RECT 50.300 51.330 50.690 51.930 ;
        RECT 50.300 47.780 50.580 51.330 ;
        RECT 50.830 51.120 51.020 52.580 ;
        RECT 52.500 52.200 52.750 65.110 ;
        RECT 62.380 64.090 62.820 64.590 ;
        RECT 56.580 60.340 56.920 60.630 ;
        RECT 56.630 60.310 56.890 60.340 ;
        RECT 54.750 56.780 55.010 57.100 ;
        RECT 54.780 54.550 54.970 56.780 ;
        RECT 56.650 54.530 56.860 60.310 ;
        RECT 60.220 59.710 60.480 59.720 ;
        RECT 60.200 59.410 60.500 59.710 ;
        RECT 60.220 59.400 60.480 59.410 ;
        RECT 57.050 58.380 57.390 58.700 ;
        RECT 57.120 54.550 57.310 58.380 ;
        RECT 57.490 56.290 57.780 56.610 ;
        RECT 57.530 54.530 57.740 56.290 ;
        RECT 58.530 55.810 58.870 56.130 ;
        RECT 58.610 54.560 58.790 55.810 ;
        RECT 52.230 51.760 52.750 52.200 ;
        RECT 52.500 51.390 52.750 51.760 ;
        RECT 51.260 51.230 51.600 51.280 ;
        RECT 51.260 51.210 51.820 51.230 ;
        RECT 50.800 51.090 51.020 51.120 ;
        RECT 50.790 50.820 51.040 51.090 ;
        RECT 51.140 51.040 51.820 51.210 ;
        RECT 51.260 51.000 51.820 51.040 ;
        RECT 51.260 50.960 51.600 51.000 ;
        RECT 50.790 50.810 51.030 50.820 ;
        RECT 50.800 50.570 51.030 50.810 ;
        RECT 52.070 50.800 52.390 51.120 ;
        RECT 50.830 48.540 50.990 50.570 ;
        RECT 52.500 50.320 53.140 51.390 ;
        RECT 57.310 51.370 57.540 52.580 ;
        RECT 58.530 51.610 58.760 52.580 ;
        RECT 57.280 50.580 57.540 51.370 ;
        RECT 58.520 51.360 58.760 51.610 ;
        RECT 51.180 50.010 51.420 50.140 ;
        RECT 51.160 49.690 51.420 50.010 ;
        RECT 52.500 49.610 52.750 50.320 ;
        RECT 51.160 49.090 51.420 49.410 ;
        RECT 51.180 48.970 51.420 49.090 ;
        RECT 51.260 48.930 51.600 48.970 ;
        RECT 51.260 48.890 51.820 48.930 ;
        RECT 51.140 48.720 51.820 48.890 ;
        RECT 51.260 48.700 51.820 48.720 ;
        RECT 51.260 48.650 51.600 48.700 ;
        RECT 52.500 48.540 53.140 49.610 ;
        RECT 54.260 48.660 54.540 48.710 ;
        RECT 50.800 48.300 51.030 48.540 ;
        RECT 50.790 48.290 51.030 48.300 ;
        RECT 50.790 48.020 51.040 48.290 ;
        RECT 51.260 48.030 51.600 48.080 ;
        RECT 52.070 48.040 52.390 48.360 ;
        RECT 52.500 48.190 52.750 48.540 ;
        RECT 54.260 48.380 54.580 48.660 ;
        RECT 54.790 48.650 54.980 48.710 ;
        RECT 57.310 48.430 57.540 50.580 ;
        RECT 58.530 49.720 58.760 51.360 ;
        RECT 59.330 51.210 59.650 51.530 ;
        RECT 58.430 49.430 58.760 49.720 ;
        RECT 50.800 47.990 51.020 48.020 ;
        RECT 51.260 48.010 51.820 48.030 ;
        RECT 50.300 47.180 50.690 47.780 ;
        RECT 50.300 46.530 50.580 47.180 ;
        RECT 50.830 46.530 51.020 47.990 ;
        RECT 51.140 47.840 51.820 48.010 ;
        RECT 51.260 47.800 51.820 47.840 ;
        RECT 51.260 47.760 51.600 47.800 ;
        RECT 52.500 47.350 53.140 48.190 ;
        RECT 57.280 47.640 57.540 48.430 ;
        RECT 52.230 47.120 53.140 47.350 ;
        RECT 52.230 46.910 52.750 47.120 ;
        RECT 52.500 46.410 52.750 46.910 ;
        RECT 57.310 46.530 57.540 47.640 ;
        RECT 58.530 46.530 58.760 49.430 ;
        RECT 60.250 49.170 60.450 59.400 ;
        RECT 62.480 54.510 62.710 64.090 ;
        RECT 63.380 60.320 63.660 60.640 ;
        RECT 62.940 59.410 63.220 59.730 ;
        RECT 60.230 49.040 60.450 49.170 ;
        RECT 60.180 48.710 60.510 49.040 ;
        RECT 59.360 47.520 59.680 47.840 ;
        RECT 60.820 46.540 61.240 52.580 ;
        RECT 62.710 48.700 62.720 48.760 ;
        RECT 61.270 48.620 61.500 48.700 ;
        RECT 62.490 48.620 62.720 48.700 ;
        RECT 62.710 48.600 62.720 48.620 ;
        RECT 62.970 47.870 63.190 59.410 ;
        RECT 62.960 47.800 63.190 47.870 ;
        RECT 62.950 47.200 63.150 47.800 ;
        RECT 63.400 47.350 63.630 60.320 ;
        RECT 64.770 54.320 65.190 66.700 ;
        RECT 65.800 54.320 66.220 66.700 ;
        RECT 68.180 64.050 68.620 64.550 ;
        RECT 68.280 57.070 68.510 64.050 ;
        RECT 72.700 58.800 73.980 70.770 ;
        RECT 76.460 65.580 76.740 65.700 ;
        RECT 76.460 65.080 76.790 65.580 ;
        RECT 72.700 58.720 74.000 58.800 ;
        RECT 72.690 58.420 74.000 58.720 ;
        RECT 69.470 57.770 69.770 58.090 ;
        RECT 68.150 57.060 68.510 57.070 ;
        RECT 68.120 56.170 68.510 57.060 ;
        RECT 68.280 54.510 68.510 56.170 ;
        RECT 69.500 54.510 69.730 57.770 ;
        RECT 75.780 57.220 76.210 57.560 ;
        RECT 76.020 54.550 76.210 57.220 ;
        RECT 76.460 54.460 76.740 65.080 ;
        RECT 78.160 60.320 78.420 60.640 ;
        RECT 77.270 59.450 77.530 59.770 ;
        RECT 77.300 55.730 77.490 59.450 ;
        RECT 78.180 55.730 78.400 60.320 ;
        RECT 80.150 57.100 80.490 73.320 ;
        RECT 100.550 70.800 103.740 71.920 ;
        RECT 84.650 69.860 85.020 69.870 ;
        RECT 84.600 69.410 85.100 69.860 ;
        RECT 80.800 61.000 81.120 61.370 ;
        RECT 80.100 57.020 80.490 57.100 ;
        RECT 80.090 56.250 80.490 57.020 ;
        RECT 80.100 56.180 80.490 56.250 ;
        RECT 77.130 55.040 77.810 55.730 ;
        RECT 78.170 55.040 78.850 55.730 ;
        RECT 80.150 54.400 80.490 56.180 ;
        RECT 80.820 55.620 81.090 61.000 ;
        RECT 84.650 57.260 85.020 69.410 ;
        RECT 85.440 65.960 85.900 66.390 ;
        RECT 81.310 56.610 81.470 57.260 ;
        RECT 81.310 56.060 81.580 56.610 ;
        RECT 81.300 56.010 81.580 56.060 ;
        RECT 81.300 55.920 81.470 56.010 ;
        RECT 81.310 55.620 81.470 55.920 ;
        RECT 81.720 55.800 81.910 57.260 ;
        RECT 83.590 56.970 83.800 57.260 ;
        RECT 83.120 56.440 83.430 56.880 ;
        RECT 83.480 56.680 83.800 56.970 ;
        RECT 81.690 55.770 81.910 55.800 ;
        RECT 80.820 55.120 81.500 55.620 ;
        RECT 81.680 55.500 81.930 55.770 ;
        RECT 81.680 55.490 81.920 55.500 ;
        RECT 81.690 55.250 81.920 55.490 ;
        RECT 80.820 54.470 81.090 55.120 ;
        RECT 81.310 52.550 81.470 55.120 ;
        RECT 81.720 53.220 81.880 55.250 ;
        RECT 82.720 54.910 83.040 55.230 ;
        RECT 83.590 54.980 83.800 56.680 ;
        RECT 84.060 56.410 84.250 57.260 ;
        RECT 83.950 56.120 84.250 56.410 ;
        RECT 82.070 54.400 82.310 54.820 ;
        RECT 83.480 54.690 83.800 54.980 ;
        RECT 83.590 54.470 83.800 54.690 ;
        RECT 82.040 54.080 82.310 54.400 ;
        RECT 84.060 54.090 84.250 56.120 ;
        RECT 84.470 54.800 85.020 57.260 ;
        RECT 84.350 54.290 85.020 54.800 ;
        RECT 82.070 53.650 82.310 54.080 ;
        RECT 83.610 53.910 83.800 53.960 ;
        RECT 83.490 53.620 83.800 53.910 ;
        RECT 83.950 53.800 84.250 54.090 ;
        RECT 82.710 53.220 83.030 53.540 ;
        RECT 81.690 52.980 81.920 53.220 ;
        RECT 81.680 52.970 81.920 52.980 ;
        RECT 81.680 52.700 81.930 52.970 ;
        RECT 81.690 52.670 81.910 52.700 ;
        RECT 81.300 52.460 81.470 52.550 ;
        RECT 81.300 52.410 81.580 52.460 ;
        RECT 81.310 51.860 81.580 52.410 ;
        RECT 81.310 51.210 81.470 51.860 ;
        RECT 81.720 51.210 81.910 52.670 ;
        RECT 83.120 51.590 83.430 52.030 ;
        RECT 83.610 52.000 83.800 53.620 ;
        RECT 84.060 52.510 84.250 53.800 ;
        RECT 83.940 52.220 84.250 52.510 ;
        RECT 83.510 51.710 83.800 52.000 ;
        RECT 83.600 51.210 83.830 51.710 ;
        RECT 84.060 51.210 84.250 52.220 ;
        RECT 84.470 51.210 85.020 54.290 ;
        RECT 85.460 53.390 85.830 65.960 ;
        RECT 86.210 61.250 86.660 61.680 ;
        RECT 85.260 53.370 85.420 53.390 ;
        RECT 85.100 53.070 85.420 53.370 ;
        RECT 85.460 53.330 85.860 53.390 ;
        RECT 64.780 48.550 66.220 48.710 ;
        RECT 62.960 47.170 63.190 47.200 ;
        RECT 51.260 45.730 51.600 45.770 ;
        RECT 51.260 45.690 51.820 45.730 ;
        RECT 51.140 45.520 51.820 45.690 ;
        RECT 51.260 45.500 51.820 45.520 ;
        RECT 51.260 45.450 51.600 45.500 ;
        RECT 52.500 45.340 53.140 46.410 ;
        RECT 62.520 45.890 62.690 46.070 ;
        RECT 52.500 41.680 52.750 45.340 ;
        RECT 62.500 45.300 62.820 45.600 ;
        RECT 62.500 45.190 62.740 45.300 ;
        RECT 62.530 45.180 62.700 45.190 ;
        RECT 62.720 45.130 62.740 45.190 ;
        RECT 62.970 43.970 63.190 47.170 ;
        RECT 62.970 43.880 63.320 43.970 ;
        RECT 62.970 43.660 63.480 43.880 ;
        RECT 48.200 41.070 48.410 41.570 ;
        RECT 49.510 41.260 49.760 41.670 ;
        RECT 52.480 41.260 52.750 41.680 ;
        RECT 54.260 41.830 54.540 42.940 ;
        RECT 54.790 42.250 54.980 42.850 ;
        RECT 56.790 42.410 57.180 42.430 ;
        RECT 56.780 42.320 57.180 42.410 ;
        RECT 56.630 42.310 57.180 42.320 ;
        RECT 54.790 42.060 56.390 42.250 ;
        RECT 54.260 41.550 55.980 41.830 ;
        RECT 55.780 41.320 55.980 41.550 ;
        RECT 48.200 40.920 48.390 41.070 ;
        RECT 47.920 40.430 48.390 40.920 ;
        RECT 48.780 40.780 49.150 40.800 ;
        RECT 48.730 40.520 49.150 40.780 ;
        RECT 48.780 40.510 49.150 40.520 ;
        RECT 47.740 39.990 48.060 40.270 ;
        RECT 48.200 40.090 48.390 40.430 ;
        RECT 48.100 39.800 48.390 40.090 ;
        RECT 48.200 39.190 48.390 39.800 ;
        RECT 47.740 38.720 48.060 39.000 ;
        RECT 48.100 38.900 48.390 39.190 ;
        RECT 48.200 38.560 48.390 38.900 ;
        RECT 47.920 38.070 48.390 38.560 ;
        RECT 48.780 38.470 49.150 38.480 ;
        RECT 48.730 38.210 49.150 38.470 ;
        RECT 48.780 38.190 49.150 38.210 ;
        RECT 48.200 37.720 48.390 38.070 ;
        RECT 47.920 37.230 48.390 37.720 ;
        RECT 48.780 37.580 49.150 37.600 ;
        RECT 48.730 37.320 49.150 37.580 ;
        RECT 48.780 37.310 49.150 37.320 ;
        RECT 47.740 36.790 48.060 37.070 ;
        RECT 48.200 36.890 48.390 37.230 ;
        RECT 48.100 36.600 48.390 36.890 ;
        RECT 48.200 35.990 48.390 36.600 ;
        RECT 47.740 35.520 48.060 35.800 ;
        RECT 48.100 35.700 48.390 35.990 ;
        RECT 48.200 35.400 48.390 35.700 ;
        RECT 49.510 35.440 49.740 41.260 ;
        RECT 52.480 40.920 52.730 41.260 ;
        RECT 55.790 41.060 55.950 41.320 ;
        RECT 55.640 40.920 55.950 41.060 ;
        RECT 51.240 40.760 51.580 40.810 ;
        RECT 51.240 40.740 51.800 40.760 ;
        RECT 51.120 40.570 51.800 40.740 ;
        RECT 51.240 40.530 51.800 40.570 ;
        RECT 51.240 40.490 51.580 40.530 ;
        RECT 52.480 39.850 53.120 40.920 ;
        RECT 55.630 40.770 55.950 40.920 ;
        RECT 55.790 40.480 55.950 40.770 ;
        RECT 55.790 39.930 56.060 40.480 ;
        RECT 55.780 39.880 56.060 39.930 ;
        RECT 56.200 40.140 56.390 42.060 ;
        RECT 56.600 42.070 57.180 42.310 ;
        RECT 56.600 42.050 57.170 42.070 ;
        RECT 56.600 42.040 56.790 42.050 ;
        RECT 56.600 41.200 56.770 42.040 ;
        RECT 61.270 41.980 61.500 42.890 ;
        RECT 62.490 42.010 62.720 42.890 ;
        RECT 60.750 41.910 61.500 41.980 ;
        RECT 60.720 41.750 61.500 41.910 ;
        RECT 62.470 41.950 62.720 42.010 ;
        RECT 65.800 42.080 66.220 48.550 ;
        RECT 68.280 45.850 68.510 48.710 ;
        RECT 69.500 47.500 69.730 48.710 ;
        RECT 74.500 47.890 74.810 48.330 ;
        RECT 69.500 46.710 69.760 47.500 ;
        RECT 76.020 47.250 76.210 48.710 ;
        RECT 76.460 48.660 76.740 48.710 ;
        RECT 76.460 48.360 76.780 48.660 ;
        RECT 78.210 48.370 78.530 48.690 ;
        RECT 80.150 48.570 80.490 48.710 ;
        RECT 80.810 48.700 81.090 48.710 ;
        RECT 80.810 48.560 81.230 48.700 ;
        RECT 80.910 48.380 81.230 48.560 ;
        RECT 81.870 48.440 82.210 48.830 ;
        RECT 76.460 48.060 76.740 48.360 ;
        RECT 76.350 47.460 76.740 48.060 ;
        RECT 81.870 48.150 82.260 48.440 ;
        RECT 78.360 47.540 78.680 47.860 ;
        RECT 80.860 47.730 81.180 48.050 ;
        RECT 74.650 46.930 74.970 47.250 ;
        RECT 76.020 47.220 76.240 47.250 ;
        RECT 76.000 46.950 76.250 47.220 ;
        RECT 76.010 46.940 76.250 46.950 ;
        RECT 68.280 45.560 68.610 45.850 ;
        RECT 68.280 45.550 68.510 45.560 ;
        RECT 68.200 45.230 68.520 45.550 ;
        RECT 68.280 43.020 68.510 45.230 ;
        RECT 69.500 44.560 69.730 46.710 ;
        RECT 76.010 46.700 76.240 46.940 ;
        RECT 75.620 46.140 75.860 46.270 ;
        RECT 75.620 45.820 75.880 46.140 ;
        RECT 75.620 45.220 75.880 45.540 ;
        RECT 75.620 45.100 75.860 45.220 ;
        RECT 76.050 44.670 76.210 46.700 ;
        RECT 76.460 45.860 76.740 47.460 ;
        RECT 77.250 47.010 77.570 47.330 ;
        RECT 78.470 46.850 78.680 46.960 ;
        RECT 80.860 46.880 81.180 47.200 ;
        RECT 78.450 46.530 78.710 46.850 ;
        RECT 81.870 46.780 82.210 48.150 ;
        RECT 82.540 47.470 82.810 48.820 ;
        RECT 83.160 48.400 83.480 48.720 ;
        RECT 82.540 47.180 82.920 47.470 ;
        RECT 76.460 45.540 76.820 45.860 ;
        RECT 77.980 45.730 78.300 46.050 ;
        RECT 69.500 43.770 69.760 44.560 ;
        RECT 74.650 44.170 74.970 44.490 ;
        RECT 76.010 44.430 76.240 44.670 ;
        RECT 76.010 44.420 76.250 44.430 ;
        RECT 76.000 44.150 76.250 44.420 ;
        RECT 76.020 44.120 76.240 44.150 ;
        RECT 68.200 42.720 68.520 43.020 ;
        RECT 60.720 41.300 61.130 41.750 ;
        RECT 56.600 40.450 56.760 41.200 ;
        RECT 56.560 40.430 56.760 40.450 ;
        RECT 57.580 40.440 57.900 40.760 ;
        RECT 56.550 40.190 56.780 40.430 ;
        RECT 56.550 40.140 56.760 40.190 ;
        RECT 56.200 40.020 56.370 40.140 ;
        RECT 52.480 39.140 52.730 39.850 ;
        RECT 55.780 39.790 55.950 39.880 ;
        RECT 55.790 39.320 55.950 39.790 ;
        RECT 55.780 39.230 55.950 39.320 ;
        RECT 55.780 39.180 56.060 39.230 ;
        RECT 51.240 38.460 51.580 38.500 ;
        RECT 51.240 38.420 51.800 38.460 ;
        RECT 51.120 38.250 51.800 38.420 ;
        RECT 51.240 38.230 51.800 38.250 ;
        RECT 51.240 38.180 51.580 38.230 ;
        RECT 52.480 38.070 53.120 39.140 ;
        RECT 55.790 38.630 56.060 39.180 ;
        RECT 56.200 39.090 56.360 40.020 ;
        RECT 56.200 38.970 56.370 39.090 ;
        RECT 56.600 38.970 56.760 40.140 ;
        RECT 57.580 39.890 57.900 40.210 ;
        RECT 58.540 39.800 58.780 41.190 ;
        RECT 52.480 37.720 52.730 38.070 ;
        RECT 51.240 37.560 51.580 37.610 ;
        RECT 51.240 37.540 51.800 37.560 ;
        RECT 51.120 37.370 51.800 37.540 ;
        RECT 51.240 37.330 51.800 37.370 ;
        RECT 51.240 37.290 51.580 37.330 ;
        RECT 52.480 36.650 53.120 37.720 ;
        RECT 55.790 37.240 55.950 38.630 ;
        RECT 56.200 38.050 56.390 38.970 ;
        RECT 56.550 38.920 56.760 38.970 ;
        RECT 56.550 38.680 56.780 38.920 ;
        RECT 57.580 38.900 57.900 39.220 ;
        RECT 58.530 39.140 58.800 39.800 ;
        RECT 56.560 38.660 56.760 38.680 ;
        RECT 56.170 38.030 56.410 38.050 ;
        RECT 56.600 38.030 56.760 38.660 ;
        RECT 57.580 38.350 57.900 38.670 ;
        RECT 56.170 37.840 56.760 38.030 ;
        RECT 56.170 37.820 56.410 37.840 ;
        RECT 55.790 36.690 56.060 37.240 ;
        RECT 52.480 35.940 52.730 36.650 ;
        RECT 55.780 36.640 56.060 36.690 ;
        RECT 56.200 36.900 56.390 37.820 ;
        RECT 56.600 37.210 56.760 37.840 ;
        RECT 56.560 37.190 56.760 37.210 ;
        RECT 57.580 37.200 57.900 37.520 ;
        RECT 56.550 36.950 56.780 37.190 ;
        RECT 56.550 36.900 56.760 36.950 ;
        RECT 56.200 36.780 56.370 36.900 ;
        RECT 55.780 36.550 55.950 36.640 ;
        RECT 55.790 36.090 55.950 36.550 ;
        RECT 55.780 36.000 55.950 36.090 ;
        RECT 55.780 35.950 56.060 36.000 ;
        RECT 48.200 35.360 48.410 35.400 ;
        RECT 47.920 34.870 48.410 35.360 ;
        RECT 48.780 35.270 49.150 35.280 ;
        RECT 48.730 35.010 49.150 35.270 ;
        RECT 48.780 34.990 49.150 35.010 ;
        RECT 48.200 34.650 48.410 34.870 ;
        RECT 49.510 34.650 49.760 35.440 ;
        RECT 51.240 35.260 51.580 35.300 ;
        RECT 51.240 35.220 51.800 35.260 ;
        RECT 51.120 35.050 51.800 35.220 ;
        RECT 51.240 35.030 51.800 35.050 ;
        RECT 51.240 34.980 51.580 35.030 ;
        RECT 52.480 34.870 53.120 35.940 ;
        RECT 55.790 35.860 56.060 35.950 ;
        RECT 56.200 35.860 56.360 36.780 ;
        RECT 53.180 35.150 53.340 35.850 ;
        RECT 52.480 34.650 52.750 34.870 ;
        RECT 42.950 31.710 43.230 32.040 ;
        RECT 39.450 31.340 39.730 31.580 ;
        RECT 38.710 30.070 39.120 30.400 ;
        RECT 38.710 28.320 39.120 28.650 ;
        RECT 38.710 26.570 39.120 26.900 ;
        RECT 39.450 25.580 39.690 31.340 ;
        RECT 42.390 31.310 42.740 31.580 ;
        RECT 46.720 31.580 47.050 32.330 ;
        RECT 48.220 31.870 48.410 34.650 ;
        RECT 49.530 34.360 49.760 34.650 ;
        RECT 49.440 33.880 49.770 34.360 ;
        RECT 49.530 31.870 49.760 33.880 ;
        RECT 52.500 31.870 52.750 34.650 ;
        RECT 53.180 34.600 53.450 35.150 ;
        RECT 53.170 34.550 53.450 34.600 ;
        RECT 53.590 34.810 53.780 35.800 ;
        RECT 53.990 35.120 54.150 35.850 ;
        RECT 55.790 35.740 56.370 35.860 ;
        RECT 56.600 35.740 56.760 36.900 ;
        RECT 57.580 36.650 57.900 36.970 ;
        RECT 58.540 36.550 58.780 39.140 ;
        RECT 60.720 39.040 61.100 41.300 ;
        RECT 62.470 39.780 62.710 41.950 ;
        RECT 65.800 41.900 66.230 42.080 ;
        RECT 65.800 41.510 66.240 41.900 ;
        RECT 68.280 41.690 68.510 42.720 ;
        RECT 65.830 41.300 66.240 41.510 ;
        RECT 64.750 40.820 65.150 41.190 ;
        RECT 65.830 40.820 66.230 41.300 ;
        RECT 64.750 40.600 66.230 40.820 ;
        RECT 62.460 39.120 62.720 39.780 ;
        RECT 60.720 37.180 61.110 39.040 ;
        RECT 58.530 36.230 58.790 36.550 ;
        RECT 53.950 35.100 54.150 35.120 ;
        RECT 54.970 35.110 55.290 35.430 ;
        RECT 55.790 35.400 56.390 35.740 ;
        RECT 56.550 35.690 56.760 35.740 ;
        RECT 56.550 35.450 56.780 35.690 ;
        RECT 57.580 35.670 57.900 35.990 ;
        RECT 56.560 35.430 56.760 35.450 ;
        RECT 53.940 34.860 54.170 35.100 ;
        RECT 53.940 34.810 54.150 34.860 ;
        RECT 53.590 34.690 53.760 34.810 ;
        RECT 53.170 34.460 53.340 34.550 ;
        RECT 53.180 34.010 53.340 34.460 ;
        RECT 53.170 33.920 53.340 34.010 ;
        RECT 53.170 33.870 53.450 33.920 ;
        RECT 53.180 33.320 53.450 33.870 ;
        RECT 53.590 33.780 53.750 34.690 ;
        RECT 53.590 33.660 53.760 33.780 ;
        RECT 53.990 33.660 54.150 34.810 ;
        RECT 54.970 34.560 55.290 34.880 ;
        RECT 55.790 34.700 55.980 35.400 ;
        RECT 53.180 31.910 53.340 33.320 ;
        RECT 53.590 32.740 53.780 33.660 ;
        RECT 53.940 33.610 54.150 33.660 ;
        RECT 53.940 33.370 54.170 33.610 ;
        RECT 54.970 33.590 55.290 33.910 ;
        RECT 53.950 33.350 54.150 33.370 ;
        RECT 53.560 32.710 53.800 32.740 ;
        RECT 53.990 32.710 54.150 33.350 ;
        RECT 54.970 33.040 55.290 33.360 ;
        RECT 53.560 32.540 54.150 32.710 ;
        RECT 53.560 32.510 53.800 32.540 ;
        RECT 48.220 31.650 48.420 31.870 ;
        RECT 40.870 31.290 41.070 31.310 ;
        RECT 40.870 31.000 41.220 31.290 ;
        RECT 40.870 29.540 41.070 29.560 ;
        RECT 40.870 29.250 41.220 29.540 ;
        RECT 40.870 27.790 41.070 27.810 ;
        RECT 40.870 27.500 41.220 27.790 ;
        RECT 40.870 26.040 41.070 26.060 ;
        RECT 40.870 25.750 41.220 26.040 ;
        RECT 42.390 25.650 42.700 31.310 ;
        RECT 44.630 31.280 44.920 31.290 ;
        RECT 44.610 31.010 44.930 31.280 ;
        RECT 44.610 31.000 44.920 31.010 ;
        RECT 45.650 30.940 45.970 31.240 ;
        RECT 42.950 29.960 43.230 30.290 ;
        RECT 44.630 29.530 44.920 29.540 ;
        RECT 44.610 29.260 44.930 29.530 ;
        RECT 44.610 29.250 44.920 29.260 ;
        RECT 45.650 29.190 45.970 29.490 ;
        RECT 42.950 28.210 43.230 28.540 ;
        RECT 44.630 27.780 44.920 27.790 ;
        RECT 44.610 27.510 44.930 27.780 ;
        RECT 44.610 27.500 44.920 27.510 ;
        RECT 45.650 27.440 45.970 27.740 ;
        RECT 42.950 26.460 43.230 26.790 ;
        RECT 44.630 26.030 44.920 26.040 ;
        RECT 44.610 25.760 44.930 26.030 ;
        RECT 44.610 25.750 44.920 25.760 ;
        RECT 45.650 25.690 45.970 25.990 ;
        RECT 39.390 25.330 39.690 25.580 ;
        RECT 42.330 25.330 42.700 25.650 ;
        RECT 46.720 25.630 47.010 31.580 ;
        RECT 47.950 31.160 48.420 31.650 ;
        RECT 48.810 31.510 49.180 31.530 ;
        RECT 48.760 31.250 49.180 31.510 ;
        RECT 49.530 31.270 49.770 31.870 ;
        RECT 52.500 31.650 52.760 31.870 ;
        RECT 51.270 31.490 51.610 31.540 ;
        RECT 51.270 31.470 51.830 31.490 ;
        RECT 52.500 31.480 53.150 31.650 ;
        RECT 51.150 31.300 51.830 31.470 ;
        RECT 48.810 31.240 49.180 31.250 ;
        RECT 47.770 30.720 48.090 31.000 ;
        RECT 48.230 30.820 48.420 31.160 ;
        RECT 48.130 30.530 48.420 30.820 ;
        RECT 48.230 29.920 48.420 30.530 ;
        RECT 47.770 29.450 48.090 29.730 ;
        RECT 48.130 29.630 48.420 29.920 ;
        RECT 48.230 29.290 48.420 29.630 ;
        RECT 47.950 28.800 48.420 29.290 ;
        RECT 48.810 29.200 49.180 29.210 ;
        RECT 48.760 28.940 49.180 29.200 ;
        RECT 48.810 28.920 49.180 28.940 ;
        RECT 48.230 28.450 48.420 28.800 ;
        RECT 47.950 27.960 48.420 28.450 ;
        RECT 48.810 28.310 49.180 28.330 ;
        RECT 48.760 28.050 49.180 28.310 ;
        RECT 48.810 28.040 49.180 28.050 ;
        RECT 47.770 27.520 48.090 27.800 ;
        RECT 48.230 27.620 48.420 27.960 ;
        RECT 48.130 27.330 48.420 27.620 ;
        RECT 48.230 26.720 48.420 27.330 ;
        RECT 47.770 26.250 48.090 26.530 ;
        RECT 48.130 26.430 48.420 26.720 ;
        RECT 48.230 26.090 48.420 26.430 ;
        RECT 46.720 25.330 47.050 25.630 ;
        RECT 47.950 25.600 48.420 26.090 ;
        RECT 48.810 26.000 49.180 26.010 ;
        RECT 48.760 25.740 49.180 26.000 ;
        RECT 48.810 25.720 49.180 25.740 ;
        RECT 48.220 25.380 48.420 25.600 ;
        RECT 49.540 25.380 49.770 31.270 ;
        RECT 51.270 31.260 51.830 31.300 ;
        RECT 51.270 31.220 51.610 31.260 ;
        RECT 52.510 30.580 53.150 31.480 ;
        RECT 53.180 31.360 53.450 31.910 ;
        RECT 53.170 31.310 53.450 31.360 ;
        RECT 53.590 31.570 53.780 32.510 ;
        RECT 53.990 31.880 54.150 32.540 ;
        RECT 53.950 31.860 54.150 31.880 ;
        RECT 54.970 31.870 55.290 32.190 ;
        RECT 53.940 31.620 54.170 31.860 ;
        RECT 53.940 31.570 54.150 31.620 ;
        RECT 53.590 31.450 53.760 31.570 ;
        RECT 53.170 31.220 53.340 31.310 ;
        RECT 53.180 30.760 53.340 31.220 ;
        RECT 53.170 30.670 53.340 30.760 ;
        RECT 53.170 30.620 53.450 30.670 ;
        RECT 52.510 29.870 52.760 30.580 ;
        RECT 53.180 30.070 53.450 30.620 ;
        RECT 53.590 30.530 53.750 31.450 ;
        RECT 53.590 30.410 53.760 30.530 ;
        RECT 53.990 30.490 54.150 31.570 ;
        RECT 54.970 31.320 55.290 31.640 ;
        RECT 55.820 31.420 55.980 34.700 ;
        RECT 56.050 34.750 56.390 35.400 ;
        RECT 56.050 31.590 56.300 34.750 ;
        RECT 56.600 34.700 56.760 35.430 ;
        RECT 57.580 35.120 57.900 35.440 ;
        RECT 58.110 33.670 58.490 35.860 ;
        RECT 58.540 35.550 58.780 36.230 ;
        RECT 58.540 34.690 58.810 35.550 ;
        RECT 58.110 31.810 58.500 33.670 ;
        RECT 58.570 31.830 58.810 34.690 ;
        RECT 56.050 31.520 56.420 31.590 ;
        RECT 56.630 31.520 56.790 31.590 ;
        RECT 56.050 31.150 56.300 31.520 ;
        RECT 58.110 31.330 58.490 31.810 ;
        RECT 58.550 31.580 58.940 31.830 ;
        RECT 58.690 31.330 58.940 31.580 ;
        RECT 56.030 31.120 56.310 31.150 ;
        RECT 56.020 30.840 56.320 31.120 ;
        RECT 58.110 31.010 58.510 31.330 ;
        RECT 60.060 31.120 60.330 35.860 ;
        RECT 60.720 35.690 61.100 37.180 ;
        RECT 62.470 36.510 62.710 39.120 ;
        RECT 62.460 36.190 62.720 36.510 ;
        RECT 62.470 35.860 62.710 36.190 ;
        RECT 60.720 34.690 61.130 35.690 ;
        RECT 60.750 31.200 61.130 34.690 ;
        RECT 62.140 35.550 62.710 35.860 ;
        RECT 64.750 35.710 65.150 40.600 ;
        RECT 62.140 31.810 62.740 35.550 ;
        RECT 64.750 34.690 65.180 35.710 ;
        RECT 65.830 34.690 66.230 40.600 ;
        RECT 68.270 39.780 68.510 41.690 ;
        RECT 69.500 42.000 69.730 43.770 ;
        RECT 74.500 43.040 74.810 43.480 ;
        RECT 69.500 41.620 70.260 42.000 ;
        RECT 76.020 41.870 76.210 44.120 ;
        RECT 76.460 43.910 76.740 45.540 ;
        RECT 78.470 45.190 78.680 46.530 ;
        RECT 80.910 46.230 81.230 46.550 ;
        RECT 81.870 46.490 82.260 46.780 ;
        RECT 80.910 45.380 81.230 45.700 ;
        RECT 81.870 45.440 82.210 46.490 ;
        RECT 78.550 44.870 78.780 45.160 ;
        RECT 81.870 45.150 82.260 45.440 ;
        RECT 80.860 44.730 81.180 45.050 ;
        RECT 76.350 43.310 76.740 43.910 ;
        RECT 80.860 43.880 81.180 44.200 ;
        RECT 81.870 43.780 82.210 45.150 ;
        RECT 82.540 44.880 82.810 47.180 ;
        RECT 83.210 46.180 83.530 46.500 ;
        RECT 83.200 45.460 83.520 45.780 ;
        RECT 82.540 44.590 82.920 44.880 ;
        RECT 68.260 39.120 68.520 39.780 ;
        RECT 68.270 36.510 68.510 39.120 ;
        RECT 69.880 39.040 70.260 41.620 ;
        RECT 74.190 41.500 74.470 41.820 ;
        RECT 74.620 41.680 76.210 41.870 ;
        RECT 72.200 39.800 72.440 41.190 ;
        RECT 73.080 40.440 73.400 40.760 ;
        RECT 74.220 40.450 74.380 41.500 ;
        RECT 74.620 41.350 74.810 41.680 ;
        RECT 76.460 41.490 76.740 43.310 ;
        RECT 80.910 43.230 81.230 43.550 ;
        RECT 81.870 43.490 82.260 43.780 ;
        RECT 78.640 42.860 78.970 43.150 ;
        RECT 81.870 43.110 82.210 43.490 ;
        RECT 82.540 43.120 82.810 44.590 ;
        RECT 83.120 43.210 83.440 43.530 ;
        RECT 78.630 42.830 79.050 42.860 ;
        RECT 79.650 42.850 80.150 42.860 ;
        RECT 79.650 42.830 80.490 42.850 ;
        RECT 78.630 42.720 80.490 42.830 ;
        RECT 78.910 42.690 79.810 42.720 ;
        RECT 80.150 42.660 80.490 42.720 ;
        RECT 80.820 42.660 81.090 42.870 ;
        RECT 84.650 42.500 85.020 51.210 ;
        RECT 84.620 42.040 85.070 42.500 ;
        RECT 84.650 42.000 85.020 42.040 ;
        RECT 85.460 41.910 85.830 53.330 ;
        RECT 75.070 41.480 76.740 41.490 ;
        RECT 74.590 41.240 74.810 41.350 ;
        RECT 74.220 40.430 74.420 40.450 ;
        RECT 73.080 39.890 73.400 40.210 ;
        RECT 74.200 40.190 74.430 40.430 ;
        RECT 74.220 40.140 74.430 40.190 ;
        RECT 74.590 40.140 74.780 41.240 ;
        RECT 75.030 41.210 76.740 41.480 ;
        RECT 85.430 41.450 85.870 41.910 ;
        RECT 85.460 41.400 85.830 41.450 ;
        RECT 75.030 41.070 75.190 41.210 ;
        RECT 75.030 40.790 75.360 41.070 ;
        RECT 75.030 40.480 75.190 40.790 ;
        RECT 72.180 39.140 72.450 39.800 ;
        RECT 69.870 37.180 70.260 39.040 ;
        RECT 68.260 36.190 68.520 36.510 ;
        RECT 68.270 35.550 68.510 36.190 ;
        RECT 68.270 34.690 68.540 35.550 ;
        RECT 69.880 34.690 70.260 37.180 ;
        RECT 72.200 36.550 72.440 39.140 ;
        RECT 73.080 38.900 73.400 39.220 ;
        RECT 74.220 38.970 74.380 40.140 ;
        RECT 74.610 40.020 74.780 40.140 ;
        RECT 74.620 39.090 74.780 40.020 ;
        RECT 74.920 39.930 75.190 40.480 ;
        RECT 74.920 39.880 75.200 39.930 ;
        RECT 75.030 39.790 75.200 39.880 ;
        RECT 75.030 39.320 75.190 39.790 ;
        RECT 86.230 39.560 86.600 61.250 ;
        RECT 92.780 60.200 93.360 60.760 ;
        RECT 89.570 58.630 90.130 59.280 ;
        RECT 90.520 59.120 91.080 59.700 ;
        RECT 91.600 59.580 92.160 60.170 ;
        RECT 89.590 57.260 90.090 58.630 ;
        RECT 87.100 56.170 87.530 56.610 ;
        RECT 86.200 39.550 86.600 39.560 ;
        RECT 75.030 39.230 75.200 39.320 ;
        RECT 74.610 38.970 74.780 39.090 ;
        RECT 74.220 38.920 74.430 38.970 ;
        RECT 74.200 38.680 74.430 38.920 ;
        RECT 73.080 38.350 73.400 38.670 ;
        RECT 74.220 38.660 74.420 38.680 ;
        RECT 74.220 38.030 74.380 38.660 ;
        RECT 74.590 38.050 74.780 38.970 ;
        RECT 74.920 39.180 75.200 39.230 ;
        RECT 74.920 38.630 75.190 39.180 ;
        RECT 86.190 39.130 86.610 39.550 ;
        RECT 86.230 39.120 86.600 39.130 ;
        RECT 74.570 38.030 74.810 38.050 ;
        RECT 74.220 37.840 74.810 38.030 ;
        RECT 73.080 37.200 73.400 37.520 ;
        RECT 74.220 37.210 74.380 37.840 ;
        RECT 74.570 37.820 74.810 37.840 ;
        RECT 74.220 37.190 74.420 37.210 ;
        RECT 73.080 36.650 73.400 36.970 ;
        RECT 74.200 36.950 74.430 37.190 ;
        RECT 74.220 36.900 74.430 36.950 ;
        RECT 74.590 36.900 74.780 37.820 ;
        RECT 75.030 37.240 75.190 38.630 ;
        RECT 72.190 36.230 72.450 36.550 ;
        RECT 72.200 34.690 72.440 36.230 ;
        RECT 73.080 35.670 73.400 35.990 ;
        RECT 74.220 35.740 74.380 36.900 ;
        RECT 74.610 36.780 74.780 36.900 ;
        RECT 74.620 35.860 74.780 36.780 ;
        RECT 74.920 36.690 75.190 37.240 ;
        RECT 74.920 36.640 75.200 36.690 ;
        RECT 75.030 36.550 75.200 36.640 ;
        RECT 75.030 36.090 75.190 36.550 ;
        RECT 75.030 36.000 75.200 36.090 ;
        RECT 74.610 35.740 74.780 35.860 ;
        RECT 74.220 35.690 74.430 35.740 ;
        RECT 74.200 35.450 74.430 35.690 ;
        RECT 73.080 35.120 73.400 35.440 ;
        RECT 74.220 35.430 74.420 35.450 ;
        RECT 74.220 34.700 74.380 35.430 ;
        RECT 74.590 34.750 74.780 35.740 ;
        RECT 74.920 35.950 75.200 36.000 ;
        RECT 74.920 35.400 75.190 35.950 ;
        RECT 75.030 34.700 75.190 35.400 ;
        RECT 62.140 31.540 62.970 31.810 ;
        RECT 56.030 30.820 56.310 30.840 ;
        RECT 51.270 29.190 51.610 29.230 ;
        RECT 51.270 29.150 51.830 29.190 ;
        RECT 51.150 28.980 51.830 29.150 ;
        RECT 51.270 28.960 51.830 28.980 ;
        RECT 51.270 28.910 51.610 28.960 ;
        RECT 52.510 28.800 53.150 29.870 ;
        RECT 53.180 29.370 53.340 30.070 ;
        RECT 53.590 29.420 53.780 30.410 ;
        RECT 53.850 30.150 54.170 30.490 ;
        RECT 54.970 30.340 55.290 30.660 ;
        RECT 53.930 30.120 54.170 30.150 ;
        RECT 53.930 29.370 54.150 30.120 ;
        RECT 54.970 29.790 55.290 30.110 ;
        RECT 54.960 29.660 55.220 29.780 ;
        RECT 54.950 29.460 55.220 29.660 ;
        RECT 52.510 28.450 52.760 28.800 ;
        RECT 51.270 28.290 51.610 28.340 ;
        RECT 51.270 28.270 51.830 28.290 ;
        RECT 51.150 28.100 51.830 28.270 ;
        RECT 51.270 28.060 51.830 28.100 ;
        RECT 51.270 28.020 51.610 28.060 ;
        RECT 52.510 27.380 53.150 28.450 ;
        RECT 52.510 26.670 52.760 27.380 ;
        RECT 51.270 25.990 51.610 26.030 ;
        RECT 51.270 25.950 51.830 25.990 ;
        RECT 51.150 25.780 51.830 25.950 ;
        RECT 51.270 25.760 51.830 25.780 ;
        RECT 51.270 25.710 51.610 25.760 ;
        RECT 52.510 25.700 53.150 26.670 ;
        RECT 52.500 25.600 53.150 25.700 ;
        RECT 52.500 25.380 52.760 25.600 ;
        RECT 53.930 25.390 54.140 29.370 ;
        RECT 54.950 28.770 55.160 29.460 ;
        RECT 56.050 29.360 56.300 30.820 ;
        RECT 58.110 29.360 58.490 31.010 ;
        RECT 60.040 30.810 60.350 31.120 ;
        RECT 60.060 29.360 60.330 30.810 ;
        RECT 62.140 29.360 62.540 31.540 ;
        RECT 62.700 31.310 62.970 31.540 ;
        RECT 64.780 31.180 65.180 34.690 ;
        RECT 68.300 33.040 68.540 34.690 ;
        RECT 87.110 34.380 87.480 56.170 ;
        RECT 89.420 54.400 90.090 57.260 ;
        RECT 89.320 54.110 90.090 54.400 ;
        RECT 87.540 53.280 87.750 53.390 ;
        RECT 88.010 53.310 88.200 53.390 ;
        RECT 88.420 53.330 88.630 53.390 ;
        RECT 89.420 51.210 90.090 54.110 ;
        RECT 87.550 47.350 87.780 47.470 ;
        RECT 87.070 33.870 87.560 34.380 ;
        RECT 87.110 33.840 87.480 33.870 ;
        RECT 68.300 32.800 68.880 33.040 ;
        RECT 66.300 30.810 66.620 31.130 ;
        RECT 66.450 30.130 66.770 30.450 ;
        RECT 66.450 29.240 66.770 29.560 ;
        RECT 54.940 28.710 55.200 28.770 ;
        RECT 54.940 28.460 55.580 28.710 ;
        RECT 66.300 28.560 66.620 28.880 ;
        RECT 54.940 28.450 55.200 28.460 ;
        RECT 54.470 27.360 54.810 27.700 ;
        RECT 54.510 27.340 54.730 27.360 ;
        RECT 39.390 12.950 39.630 25.330 ;
        RECT 42.330 24.500 42.640 25.330 ;
        RECT 46.760 25.010 47.050 25.330 ;
        RECT 47.260 25.030 47.600 25.350 ;
        RECT 46.730 24.660 47.080 25.010 ;
        RECT 42.290 24.170 42.660 24.500 ;
        RECT 46.760 24.200 47.050 24.660 ;
        RECT 47.260 24.420 47.510 25.030 ;
        RECT 48.220 24.440 48.410 25.380 ;
        RECT 52.500 24.970 52.750 25.380 ;
        RECT 53.900 25.070 54.180 25.390 ;
        RECT 54.510 25.060 54.710 27.340 ;
        RECT 54.860 26.410 55.180 26.730 ;
        RECT 54.970 25.770 55.160 25.880 ;
        RECT 54.910 25.450 55.230 25.770 ;
        RECT 52.470 24.680 52.810 24.970 ;
        RECT 54.470 24.740 54.750 25.060 ;
        RECT 54.930 25.050 55.210 25.450 ;
        RECT 42.330 22.960 42.640 24.170 ;
        RECT 46.190 23.920 47.050 24.200 ;
        RECT 46.110 23.910 47.050 23.920 ;
        RECT 47.210 24.310 47.510 24.420 ;
        RECT 46.110 23.440 46.570 23.910 ;
        RECT 42.280 22.480 42.700 22.960 ;
        RECT 47.210 22.800 47.400 24.310 ;
        RECT 48.160 24.120 48.480 24.440 ;
        RECT 55.400 23.830 55.580 28.460 ;
        RECT 58.230 28.080 58.490 28.400 ;
        RECT 58.230 27.220 58.390 28.080 ;
        RECT 66.300 28.040 66.620 28.360 ;
        RECT 66.450 27.360 66.770 27.680 ;
        RECT 58.100 26.900 58.390 27.220 ;
        RECT 66.450 26.470 66.770 26.790 ;
        RECT 56.720 24.990 56.980 25.020 ;
        RECT 56.700 24.690 57.000 24.990 ;
        RECT 56.720 24.680 56.980 24.690 ;
        RECT 47.570 23.450 47.890 23.770 ;
        RECT 48.660 23.450 48.980 23.770 ;
        RECT 49.760 23.440 50.080 23.760 ;
        RECT 52.600 23.440 52.920 23.760 ;
        RECT 53.700 23.450 54.020 23.770 ;
        RECT 54.790 23.450 55.110 23.770 ;
        RECT 55.400 23.530 55.880 23.830 ;
        RECT 56.730 23.760 56.950 24.680 ;
        RECT 58.690 24.550 58.940 25.780 ;
        RECT 60.750 25.540 61.130 25.640 ;
        RECT 62.700 24.570 62.970 25.800 ;
        RECT 66.300 25.790 66.620 26.110 ;
        RECT 67.380 25.540 67.610 31.590 ;
        RECT 68.640 31.460 68.880 32.800 ;
        RECT 68.640 27.240 68.870 31.460 ;
        RECT 73.760 30.400 74.020 30.460 ;
        RECT 73.750 30.140 74.020 30.400 ;
        RECT 73.240 29.210 73.500 29.530 ;
        RECT 72.770 27.370 73.030 27.690 ;
        RECT 68.600 27.230 68.880 27.240 ;
        RECT 68.600 26.910 68.900 27.230 ;
        RECT 65.520 25.000 65.950 25.400 ;
        RECT 58.680 24.290 59.000 24.550 ;
        RECT 62.700 24.260 63.050 24.570 ;
        RECT 55.480 23.420 55.880 23.530 ;
        RECT 56.670 23.360 57.010 23.760 ;
        RECT 57.380 23.480 57.700 23.800 ;
        RECT 58.470 23.480 58.790 23.800 ;
        RECT 59.570 23.470 59.890 23.790 ;
        RECT 62.410 23.470 62.730 23.790 ;
        RECT 63.510 23.480 63.830 23.800 ;
        RECT 64.600 23.480 64.920 23.800 ;
        RECT 56.730 23.280 56.950 23.360 ;
        RECT 65.560 23.210 65.910 25.000 ;
        RECT 67.380 24.440 67.600 25.540 ;
        RECT 68.640 25.040 68.870 26.910 ;
        RECT 72.270 26.440 72.530 26.760 ;
        RECT 68.640 24.810 71.850 25.040 ;
        RECT 68.640 24.800 68.870 24.810 ;
        RECT 67.090 24.200 67.600 24.440 ;
        RECT 46.770 22.480 47.400 22.800 ;
        RECT 48.120 22.770 48.440 23.090 ;
        RECT 49.210 22.750 49.530 23.070 ;
        RECT 53.150 22.750 53.470 23.070 ;
        RECT 54.240 22.770 54.560 23.090 ;
        RECT 57.930 22.800 58.250 23.120 ;
        RECT 59.020 22.780 59.340 23.100 ;
        RECT 62.960 22.780 63.280 23.100 ;
        RECT 64.050 22.800 64.370 23.120 ;
        RECT 67.090 22.950 67.320 24.200 ;
        RECT 71.620 23.840 71.850 24.810 ;
        RECT 71.570 23.440 71.880 23.840 ;
        RECT 66.980 22.510 67.440 22.950 ;
        RECT 46.770 22.380 47.210 22.480 ;
        RECT 48.120 21.400 48.440 21.720 ;
        RECT 49.210 21.400 49.530 21.720 ;
        RECT 53.150 21.400 53.470 21.720 ;
        RECT 54.240 21.400 54.560 21.720 ;
        RECT 57.930 21.430 58.250 21.750 ;
        RECT 59.020 21.430 59.340 21.750 ;
        RECT 62.960 21.430 63.280 21.750 ;
        RECT 64.050 21.430 64.370 21.750 ;
        RECT 47.560 20.670 47.880 20.990 ;
        RECT 48.660 20.670 48.980 20.990 ;
        RECT 49.760 20.670 50.080 20.990 ;
        RECT 52.600 20.670 52.920 20.990 ;
        RECT 53.700 20.670 54.020 20.990 ;
        RECT 54.800 20.670 55.120 20.990 ;
        RECT 57.370 20.700 57.690 21.020 ;
        RECT 58.470 20.700 58.790 21.020 ;
        RECT 59.570 20.700 59.890 21.020 ;
        RECT 62.410 20.700 62.730 21.020 ;
        RECT 63.510 20.700 63.830 21.020 ;
        RECT 64.610 20.700 64.930 21.020 ;
        RECT 71.620 20.270 71.850 23.440 ;
        RECT 71.490 20.050 71.850 20.270 ;
        RECT 71.290 19.820 71.850 20.050 ;
        RECT 71.290 19.810 71.830 19.820 ;
        RECT 47.560 19.300 47.880 19.620 ;
        RECT 48.660 19.300 48.980 19.620 ;
        RECT 49.760 19.300 50.080 19.620 ;
        RECT 52.600 19.300 52.920 19.620 ;
        RECT 53.700 19.300 54.020 19.620 ;
        RECT 54.800 19.300 55.120 19.620 ;
        RECT 57.370 19.330 57.690 19.650 ;
        RECT 58.470 19.330 58.790 19.650 ;
        RECT 59.570 19.330 59.890 19.650 ;
        RECT 62.410 19.330 62.730 19.650 ;
        RECT 63.510 19.330 63.830 19.650 ;
        RECT 64.610 19.330 64.930 19.650 ;
        RECT 68.790 19.260 69.110 19.580 ;
        RECT 69.890 19.270 70.210 19.590 ;
        RECT 70.980 19.270 71.300 19.590 ;
        RECT 46.990 18.950 47.310 18.980 ;
        RECT 55.370 18.970 55.690 18.980 ;
        RECT 46.980 18.660 47.310 18.950 ;
        RECT 46.980 18.510 47.300 18.660 ;
        RECT 48.120 18.620 48.440 18.940 ;
        RECT 49.210 18.620 49.530 18.940 ;
        RECT 53.150 18.620 53.470 18.940 ;
        RECT 54.240 18.620 54.560 18.940 ;
        RECT 46.980 18.190 47.320 18.510 ;
        RECT 46.980 17.200 47.300 18.190 ;
        RECT 46.860 16.600 47.400 17.200 ;
        RECT 55.350 16.180 55.690 18.970 ;
        RECT 56.800 18.960 57.120 19.010 ;
        RECT 56.780 18.540 57.120 18.960 ;
        RECT 57.930 18.650 58.250 18.970 ;
        RECT 59.020 18.650 59.340 18.970 ;
        RECT 62.960 18.650 63.280 18.970 ;
        RECT 64.050 18.650 64.370 18.970 ;
        RECT 65.180 18.690 65.500 19.010 ;
        RECT 65.200 18.540 65.470 18.690 ;
        RECT 68.230 18.560 68.550 18.880 ;
        RECT 69.340 18.570 69.660 18.890 ;
        RECT 70.430 18.590 70.750 18.910 ;
        RECT 72.270 18.600 72.520 26.440 ;
        RECT 72.770 19.500 73.020 27.370 ;
        RECT 73.250 20.410 73.500 29.210 ;
        RECT 73.750 21.300 74.000 30.140 ;
        RECT 89.590 22.800 90.090 51.210 ;
        RECT 90.520 28.080 91.020 59.120 ;
        RECT 91.650 33.310 92.150 59.580 ;
        RECT 92.780 38.480 93.280 60.200 ;
        RECT 101.640 58.600 102.920 70.800 ;
        RECT 101.630 57.260 102.920 58.600 ;
        RECT 101.640 56.770 102.920 57.260 ;
        RECT 106.000 55.590 106.200 55.620 ;
        RECT 105.910 55.090 106.220 55.590 ;
        RECT 102.090 53.820 102.440 54.300 ;
        RECT 95.660 53.240 96.080 53.390 ;
        RECT 96.690 53.240 97.110 53.390 ;
        RECT 95.660 53.100 97.110 53.240 ;
        RECT 93.320 47.390 93.640 47.690 ;
        RECT 96.690 47.340 97.110 53.100 ;
        RECT 98.100 50.620 98.570 51.110 ;
        RECT 92.730 37.920 93.280 38.480 ;
        RECT 91.640 32.750 92.160 33.310 ;
        RECT 90.510 27.560 91.030 28.080 ;
        RECT 89.430 22.230 90.090 22.800 ;
        RECT 73.700 20.720 74.070 21.300 ;
        RECT 73.170 19.830 73.540 20.410 ;
        RECT 72.680 18.920 73.050 19.500 ;
        RECT 56.780 18.220 57.130 18.540 ;
        RECT 65.170 18.220 65.490 18.540 ;
        RECT 55.290 15.660 55.750 16.180 ;
        RECT 56.780 15.290 57.120 18.220 ;
        RECT 56.690 14.770 57.210 15.290 ;
        RECT 65.200 14.410 65.470 18.220 ;
        RECT 68.240 17.220 68.560 17.540 ;
        RECT 69.340 17.220 69.660 17.540 ;
        RECT 70.430 17.220 70.750 17.540 ;
        RECT 70.940 16.810 71.270 18.380 ;
        RECT 72.210 18.030 72.560 18.600 ;
        RECT 68.790 16.490 69.110 16.810 ;
        RECT 69.890 16.490 70.210 16.810 ;
        RECT 70.940 16.490 71.310 16.810 ;
        RECT 70.940 15.440 71.270 16.490 ;
        RECT 71.720 16.460 71.990 16.490 ;
        RECT 71.710 15.930 71.990 16.460 ;
        RECT 71.710 15.630 72.170 15.930 ;
        RECT 71.700 15.610 72.170 15.630 ;
        RECT 68.790 15.120 69.110 15.440 ;
        RECT 69.890 15.120 70.210 15.440 ;
        RECT 70.940 15.120 71.310 15.440 ;
        RECT 71.700 15.180 71.990 15.610 ;
        RECT 68.240 14.450 68.560 14.770 ;
        RECT 69.340 14.440 69.660 14.760 ;
        RECT 70.430 14.440 70.750 14.760 ;
        RECT 65.090 13.850 65.580 14.410 ;
        RECT 38.990 11.630 39.640 12.950 ;
        RECT 70.940 8.390 71.270 15.120 ;
        RECT 71.560 14.480 71.880 14.800 ;
        RECT 71.550 14.010 71.870 14.330 ;
        RECT 89.590 13.920 90.090 22.230 ;
        RECT 90.520 14.830 91.020 27.560 ;
        RECT 91.650 15.700 92.150 32.750 ;
        RECT 92.780 17.210 93.280 37.920 ;
        RECT 95.670 24.770 96.250 25.330 ;
        RECT 95.700 24.760 96.210 24.770 ;
        RECT 92.780 16.650 93.340 17.210 ;
        RECT 92.780 16.520 93.280 16.650 ;
        RECT 95.700 12.890 96.200 24.760 ;
        RECT 95.070 11.610 96.200 12.890 ;
        RECT 70.880 8.000 71.310 8.390 ;
        RECT 37.340 7.340 37.710 7.720 ;
        RECT 98.150 7.270 98.550 50.620 ;
        RECT 99.170 50.530 99.400 53.390 ;
        RECT 100.390 52.180 100.620 53.390 ;
        RECT 100.390 51.390 100.650 52.180 ;
        RECT 99.170 50.370 99.500 50.530 ;
        RECT 99.070 50.240 99.500 50.370 ;
        RECT 99.070 50.010 99.490 50.240 ;
        RECT 36.690 6.720 37.080 7.110 ;
        RECT 98.140 6.810 98.610 7.270 ;
        RECT 36.090 6.090 36.470 6.480 ;
        RECT 99.080 6.470 99.470 50.010 ;
        RECT 100.390 49.240 100.620 51.390 ;
        RECT 100.390 48.450 100.650 49.240 ;
        RECT 100.390 48.050 100.620 48.450 ;
        RECT 99.990 47.620 100.620 48.050 ;
        RECT 100.010 47.340 100.620 47.620 ;
        RECT 100.850 47.360 101.230 47.370 ;
        RECT 99.050 6.000 99.510 6.470 ;
        RECT 35.500 5.460 35.850 5.830 ;
        RECT 100.010 5.650 100.400 47.340 ;
        RECT 100.830 47.060 101.250 47.360 ;
        RECT 99.990 5.190 100.460 5.650 ;
        RECT 34.860 4.780 35.220 5.160 ;
        RECT 100.850 4.850 101.230 47.060 ;
        RECT 102.190 23.830 102.420 53.820 ;
        RECT 105.390 52.570 105.700 53.010 ;
        RECT 105.540 51.610 105.860 51.930 ;
        RECT 106.000 51.840 106.200 55.090 ;
        RECT 108.580 53.960 108.800 54.180 ;
        RECT 108.570 53.920 108.800 53.960 ;
        RECT 106.360 53.640 106.560 53.680 ;
        RECT 108.570 53.600 108.830 53.920 ;
        RECT 108.990 53.750 109.190 54.070 ;
        RECT 108.990 53.460 109.310 53.750 ;
        RECT 106.910 51.930 107.100 53.390 ;
        RECT 107.350 53.370 107.630 53.390 ;
        RECT 108.990 53.370 109.190 53.460 ;
        RECT 107.350 53.070 107.690 53.370 ;
        RECT 107.350 52.740 107.630 53.070 ;
        RECT 107.240 52.140 107.630 52.740 ;
        RECT 108.990 53.050 109.420 53.370 ;
        RECT 108.990 52.460 109.190 53.050 ;
        RECT 109.510 52.540 109.700 72.120 ;
        RECT 112.850 63.270 113.670 63.360 ;
        RECT 112.790 62.580 113.670 63.270 ;
        RECT 109.870 53.620 110.060 53.680 ;
        RECT 110.840 53.530 111.100 53.850 ;
        RECT 111.840 53.790 112.110 53.860 ;
        RECT 111.840 53.540 112.210 53.790 ;
        RECT 110.910 53.390 111.100 53.530 ;
        RECT 110.910 53.250 111.380 53.390 ;
        RECT 111.700 53.380 111.980 53.390 ;
        RECT 112.020 53.380 112.210 53.540 ;
        RECT 110.910 53.140 111.100 53.250 ;
        RECT 111.700 53.240 112.210 53.380 ;
        RECT 110.910 53.060 111.220 53.140 ;
        RECT 111.800 53.130 112.210 53.240 ;
        RECT 112.500 53.750 112.690 54.070 ;
        RECT 112.790 53.750 113.500 62.580 ;
        RECT 112.500 53.500 113.500 53.750 ;
        RECT 112.500 53.460 113.700 53.500 ;
        RECT 111.800 53.060 112.350 53.130 ;
        RECT 109.890 52.620 110.210 52.940 ;
        RECT 110.890 52.850 111.220 53.060 ;
        RECT 112.020 53.040 112.350 53.060 ;
        RECT 110.890 52.770 111.120 52.850 ;
        RECT 111.460 52.730 111.780 52.940 ;
        RECT 112.120 52.840 112.350 53.040 ;
        RECT 111.460 52.620 112.070 52.730 ;
        RECT 109.250 52.220 109.700 52.540 ;
        RECT 111.750 52.410 112.070 52.620 ;
        RECT 112.500 52.460 112.690 53.460 ;
        RECT 106.910 51.900 107.130 51.930 ;
        RECT 106.890 51.630 107.140 51.900 ;
        RECT 106.900 51.620 107.140 51.630 ;
        RECT 106.900 51.380 107.130 51.620 ;
        RECT 106.510 50.820 106.750 50.950 ;
        RECT 106.510 50.500 106.770 50.820 ;
        RECT 106.510 49.900 106.770 50.220 ;
        RECT 106.510 49.780 106.750 49.900 ;
        RECT 106.940 49.350 107.100 51.380 ;
        RECT 107.350 50.540 107.630 52.140 ;
        RECT 108.140 51.690 108.460 52.010 ;
        RECT 108.580 50.810 108.800 50.980 ;
        RECT 108.990 50.950 109.190 51.950 ;
        RECT 109.510 51.850 109.700 52.220 ;
        RECT 112.760 52.150 113.700 53.460 ;
        RECT 114.050 53.080 114.370 53.400 ;
        RECT 111.750 51.790 112.070 51.880 ;
        RECT 109.360 51.530 109.570 51.640 ;
        RECT 109.340 51.210 109.600 51.530 ;
        RECT 109.890 51.470 110.210 51.790 ;
        RECT 110.890 51.560 111.120 51.640 ;
        RECT 111.460 51.560 112.070 51.790 ;
        RECT 110.890 51.350 111.220 51.560 ;
        RECT 111.460 51.470 111.780 51.560 ;
        RECT 112.120 51.370 112.350 51.570 ;
        RECT 110.910 51.270 111.220 51.350 ;
        RECT 112.020 51.280 112.350 51.370 ;
        RECT 107.350 50.220 107.710 50.540 ;
        RECT 108.570 50.400 108.830 50.810 ;
        RECT 108.990 50.730 109.310 50.950 ;
        RECT 108.870 50.660 109.310 50.730 ;
        RECT 108.870 50.550 109.190 50.660 ;
        RECT 108.870 50.410 109.310 50.550 ;
        RECT 108.580 50.230 108.800 50.400 ;
        RECT 108.990 50.260 109.310 50.410 ;
        RECT 105.540 48.850 105.860 49.170 ;
        RECT 106.900 49.110 107.130 49.350 ;
        RECT 106.900 49.100 107.140 49.110 ;
        RECT 106.890 48.830 107.140 49.100 ;
        RECT 106.910 48.800 107.130 48.830 ;
        RECT 105.390 47.720 105.700 48.160 ;
        RECT 106.360 47.630 106.560 47.670 ;
        RECT 106.910 47.340 107.100 48.800 ;
        RECT 107.350 48.590 107.630 50.220 ;
        RECT 108.990 49.260 109.190 50.260 ;
        RECT 109.360 49.870 109.570 51.210 ;
        RECT 110.910 50.880 111.100 51.270 ;
        RECT 112.020 51.230 112.210 51.280 ;
        RECT 111.800 50.910 112.210 51.230 ;
        RECT 110.840 50.330 111.100 50.880 ;
        RECT 112.020 50.870 112.210 50.910 ;
        RECT 111.840 50.620 112.210 50.870 ;
        RECT 112.500 50.950 112.690 51.950 ;
        RECT 112.760 51.860 113.810 52.150 ;
        RECT 112.760 50.950 113.700 51.860 ;
        RECT 112.500 50.660 113.700 50.950 ;
        RECT 114.100 50.860 114.420 51.180 ;
        RECT 111.840 50.590 112.110 50.620 ;
        RECT 111.840 50.380 112.210 50.590 ;
        RECT 110.910 49.940 111.100 50.330 ;
        RECT 111.800 50.060 112.210 50.380 ;
        RECT 110.910 49.860 111.220 49.940 ;
        RECT 109.440 49.550 109.670 49.840 ;
        RECT 109.890 49.420 110.210 49.740 ;
        RECT 110.890 49.650 111.220 49.860 ;
        RECT 112.020 49.930 112.210 50.060 ;
        RECT 112.500 50.550 112.690 50.660 ;
        RECT 112.760 50.550 113.700 50.660 ;
        RECT 112.500 50.260 113.700 50.550 ;
        RECT 112.020 49.840 112.350 49.930 ;
        RECT 111.460 49.730 111.780 49.740 ;
        RECT 110.890 49.570 111.120 49.650 ;
        RECT 111.460 49.420 112.070 49.730 ;
        RECT 112.120 49.640 112.350 49.840 ;
        RECT 111.750 49.410 112.070 49.420 ;
        RECT 112.500 49.260 112.690 50.260 ;
        RECT 112.760 49.560 113.700 50.260 ;
        RECT 114.090 50.140 114.410 50.460 ;
        RECT 112.760 49.270 113.810 49.560 ;
        RECT 107.240 47.990 107.630 48.590 ;
        RECT 107.350 47.340 107.630 47.990 ;
        RECT 108.990 47.750 109.190 48.750 ;
        RECT 111.750 48.590 112.070 48.880 ;
        RECT 109.890 48.270 110.210 48.590 ;
        RECT 111.460 48.560 112.070 48.590 ;
        RECT 110.890 48.360 111.120 48.440 ;
        RECT 110.890 48.150 111.220 48.360 ;
        RECT 111.460 48.270 111.780 48.560 ;
        RECT 112.120 48.230 112.350 48.370 ;
        RECT 110.910 48.070 111.220 48.150 ;
        RECT 111.800 48.080 112.350 48.230 ;
        RECT 108.570 47.290 108.830 47.610 ;
        RECT 108.990 47.460 109.310 47.750 ;
        RECT 109.510 47.540 109.830 47.840 ;
        RECT 109.870 47.630 110.060 47.690 ;
        RECT 110.910 47.680 111.100 48.070 ;
        RECT 111.800 47.910 112.210 48.080 ;
        RECT 110.840 47.540 111.100 47.680 ;
        RECT 112.020 47.670 112.210 47.910 ;
        RECT 111.840 47.550 112.210 47.670 ;
        RECT 109.510 47.510 109.940 47.540 ;
        RECT 110.540 47.530 111.100 47.540 ;
        RECT 110.540 47.510 111.380 47.530 ;
        RECT 109.510 47.480 111.380 47.510 ;
        RECT 108.570 47.250 108.800 47.290 ;
        RECT 108.580 47.030 108.800 47.250 ;
        RECT 108.990 47.140 109.190 47.460 ;
        RECT 109.660 47.430 111.380 47.480 ;
        RECT 109.690 47.400 111.380 47.430 ;
        RECT 109.720 47.380 111.380 47.400 ;
        RECT 109.790 47.370 110.750 47.380 ;
        RECT 110.840 47.360 111.380 47.380 ;
        RECT 111.040 47.340 111.380 47.360 ;
        RECT 111.710 47.420 112.210 47.550 ;
        RECT 112.500 47.750 112.690 48.750 ;
        RECT 112.760 47.800 113.700 49.270 ;
        RECT 114.010 47.890 114.330 48.210 ;
        RECT 112.760 47.790 113.500 47.800 ;
        RECT 112.790 47.750 113.500 47.790 ;
        RECT 112.500 47.460 113.500 47.750 ;
        RECT 111.710 47.350 112.110 47.420 ;
        RECT 111.710 47.340 111.980 47.350 ;
        RECT 112.500 47.140 112.690 47.460 ;
        RECT 112.790 43.580 113.500 47.460 ;
        RECT 112.660 42.790 113.500 43.580 ;
        RECT 108.380 24.750 109.100 25.320 ;
        RECT 102.190 23.600 102.430 23.830 ;
        RECT 102.190 16.050 102.420 23.600 ;
        RECT 108.440 17.740 108.950 24.750 ;
        RECT 108.300 17.690 108.950 17.740 ;
        RECT 108.290 17.510 108.950 17.690 ;
        RECT 108.260 17.500 108.950 17.510 ;
        RECT 108.260 17.130 108.860 17.500 ;
        RECT 102.190 15.820 102.550 16.050 ;
        RECT 102.190 14.440 102.420 15.820 ;
        RECT 108.260 15.260 108.840 17.130 ;
        RECT 107.690 14.940 108.840 15.260 ;
        RECT 107.910 14.590 108.840 14.940 ;
        RECT 102.190 14.210 102.550 14.440 ;
        RECT 107.690 14.270 108.840 14.590 ;
        RECT 102.190 12.840 102.420 14.210 ;
        RECT 108.260 13.490 108.840 14.270 ;
        RECT 107.850 13.300 108.170 13.350 ;
        RECT 107.620 13.070 108.170 13.300 ;
        RECT 107.850 13.030 108.170 13.070 ;
        RECT 108.310 12.890 108.840 13.490 ;
        RECT 108.270 12.880 108.840 12.890 ;
        RECT 102.190 12.610 102.550 12.840 ;
        RECT 102.190 11.220 102.420 12.610 ;
        RECT 108.260 11.880 108.840 12.880 ;
        RECT 107.850 11.690 108.170 11.740 ;
        RECT 103.670 11.630 104.180 11.690 ;
        RECT 103.670 11.460 105.910 11.630 ;
        RECT 107.620 11.460 108.170 11.690 ;
        RECT 103.900 11.430 105.910 11.460 ;
        RECT 102.190 10.990 102.550 11.220 ;
        RECT 102.190 9.620 102.420 10.990 ;
        RECT 102.910 9.910 103.230 9.990 ;
        RECT 104.230 9.910 104.740 10.050 ;
        RECT 102.910 9.730 104.750 9.910 ;
        RECT 102.190 9.390 102.550 9.620 ;
        RECT 102.190 8.000 102.420 9.390 ;
        RECT 105.740 8.470 105.910 11.430 ;
        RECT 107.850 11.420 108.170 11.460 ;
        RECT 108.310 11.280 108.840 11.880 ;
        RECT 108.260 10.270 108.840 11.280 ;
        RECT 107.840 10.080 108.160 10.130 ;
        RECT 107.610 9.850 108.160 10.080 ;
        RECT 107.840 9.810 108.160 9.850 ;
        RECT 108.300 9.670 108.840 10.270 ;
        RECT 108.260 8.650 108.840 9.670 ;
        RECT 105.580 8.250 106.090 8.470 ;
        RECT 107.850 8.460 108.170 8.510 ;
        RECT 105.580 8.240 105.910 8.250 ;
        RECT 105.740 8.180 105.910 8.240 ;
        RECT 107.620 8.230 108.170 8.460 ;
        RECT 107.850 8.190 108.170 8.230 ;
        RECT 108.310 8.050 108.840 8.650 ;
        RECT 102.190 7.770 102.550 8.000 ;
        RECT 102.190 6.400 102.420 7.770 ;
        RECT 108.260 7.040 108.840 8.050 ;
        RECT 107.840 6.850 108.160 6.900 ;
        RECT 107.610 6.620 108.160 6.850 ;
        RECT 107.840 6.580 108.160 6.620 ;
        RECT 108.300 6.440 108.840 7.040 ;
        RECT 102.190 6.170 102.550 6.400 ;
        RECT 34.270 4.540 34.610 4.550 ;
        RECT 34.250 4.170 34.630 4.540 ;
        RECT 100.820 4.390 101.260 4.850 ;
        RECT 102.190 4.780 102.420 6.170 ;
        RECT 107.430 4.930 107.750 5.250 ;
        RECT 102.190 4.550 102.550 4.780 ;
        RECT 107.480 4.700 107.710 4.930 ;
        RECT 108.260 4.570 108.840 6.440 ;
        RECT 102.190 4.480 102.420 4.550 ;
        RECT 34.270 4.160 34.600 4.170 ;
        RECT 107.840 3.650 108.160 3.700 ;
        RECT 107.610 3.420 108.160 3.650 ;
        RECT 107.840 3.380 108.160 3.420 ;
        RECT 32.490 2.320 32.840 2.650 ;
        RECT 108.300 2.360 108.840 4.570 ;
        RECT 32.510 2.260 32.840 2.320 ;
        RECT 104.600 1.940 104.920 1.990 ;
        RECT 105.540 1.940 105.860 1.990 ;
        RECT 104.370 1.710 104.920 1.940 ;
        RECT 105.310 1.710 105.860 1.940 ;
        RECT 106.490 1.920 106.810 1.970 ;
        RECT 107.800 1.940 108.120 1.990 ;
        RECT 104.600 1.670 104.920 1.710 ;
        RECT 105.540 1.670 105.860 1.710 ;
        RECT 106.260 1.690 106.810 1.920 ;
        RECT 107.570 1.710 108.120 1.940 ;
        RECT 106.490 1.650 106.810 1.690 ;
        RECT 107.800 1.670 108.120 1.710 ;
        RECT 31.220 1.040 31.570 1.370 ;
        RECT 31.220 0.970 31.550 1.040 ;
        RECT 29.080 0.310 30.320 0.640 ;
        RECT 30.610 0.340 31.050 0.760 ;
        RECT 29.080 0.200 29.660 0.310 ;
      LAYER via ;
        RECT 2.030 70.080 2.420 70.470 ;
        RECT 2.110 66.630 2.500 67.020 ;
        RECT 3.490 65.460 3.750 65.720 ;
        RECT 11.430 64.770 11.690 65.030 ;
        RECT 12.790 64.850 13.050 65.110 ;
        RECT 13.480 64.840 13.740 65.100 ;
        RECT 3.410 62.760 3.830 63.180 ;
        RECT 9.360 61.360 9.650 61.940 ;
        RECT 10.710 61.110 10.970 61.370 ;
        RECT 20.570 61.130 20.830 61.390 ;
        RECT 22.650 60.300 22.910 60.560 ;
        RECT 17.730 54.560 17.990 54.820 ;
        RECT 18.820 54.570 19.080 54.830 ;
        RECT 16.570 54.050 16.830 54.310 ;
        RECT 17.300 54.060 17.560 54.320 ;
        RECT 17.740 53.570 18.000 53.830 ;
        RECT 18.830 53.580 19.090 53.840 ;
        RECT 16.540 53.130 16.800 53.390 ;
        RECT 17.280 53.140 17.540 53.400 ;
        RECT 17.740 52.580 18.000 52.840 ;
        RECT 18.830 52.590 19.090 52.850 ;
        RECT 16.550 52.210 16.810 52.470 ;
        RECT 15.900 51.190 16.160 51.450 ;
        RECT 15.860 50.230 16.120 50.490 ;
        RECT 15.900 49.270 16.160 49.530 ;
        RECT 17.260 52.150 17.520 52.410 ;
        RECT 18.760 52.200 19.020 52.460 ;
        RECT 18.730 51.740 18.990 52.000 ;
        RECT 18.760 51.210 19.020 51.470 ;
        RECT 18.730 50.750 18.990 51.010 ;
        RECT 18.760 50.220 19.020 50.480 ;
        RECT 28.440 59.870 28.750 60.180 ;
        RECT 45.020 67.510 45.440 67.930 ;
        RECT 41.170 66.750 41.590 67.170 ;
        RECT 64.790 66.750 66.140 67.170 ;
        RECT 46.690 65.140 47.130 65.580 ;
        RECT 52.410 65.140 52.850 65.580 ;
        RECT 42.270 64.120 42.710 64.560 ;
        RECT 39.510 61.100 39.770 61.360 ;
        RECT 32.440 60.410 32.700 60.670 ;
        RECT 31.270 59.420 31.540 59.680 ;
        RECT 19.940 58.640 20.290 58.990 ;
        RECT 25.190 58.950 25.450 59.210 ;
        RECT 40.960 57.930 41.220 58.190 ;
        RECT 38.860 57.090 39.120 57.350 ;
        RECT 20.960 56.400 21.220 56.790 ;
        RECT 37.360 56.410 37.690 56.670 ;
        RECT 20.320 55.580 20.580 55.980 ;
        RECT 20.340 54.470 20.600 54.730 ;
        RECT 18.730 49.760 18.990 50.020 ;
        RECT 15.860 33.990 16.120 34.460 ;
        RECT 16.500 33.990 16.760 34.460 ;
        RECT 14.500 32.960 14.760 33.220 ;
        RECT 13.980 32.560 14.240 32.820 ;
        RECT 4.700 31.310 5.360 31.970 ;
        RECT 16.580 32.940 16.840 33.200 ;
        RECT 18.340 32.950 18.610 33.220 ;
        RECT 15.920 32.580 16.180 32.840 ;
        RECT 14.000 28.650 14.260 28.910 ;
        RECT 9.910 26.790 10.280 27.160 ;
        RECT 4.740 25.450 5.400 26.110 ;
        RECT 14.000 25.560 14.260 25.820 ;
        RECT 18.840 32.560 19.100 32.820 ;
        RECT 20.340 53.550 20.600 53.810 ;
        RECT 20.310 52.630 20.570 52.890 ;
        RECT 20.060 52.100 20.320 52.360 ;
        RECT 20.060 51.110 20.320 51.370 ;
        RECT 20.060 50.120 20.320 50.380 ;
        RECT 36.730 54.690 37.060 55.020 ;
        RECT 36.160 53.210 36.490 53.540 ;
        RECT 20.950 51.540 21.210 51.800 ;
        RECT 35.520 51.610 35.850 51.940 ;
        RECT 34.880 51.040 35.210 51.370 ;
        RECT 20.960 50.580 21.220 50.840 ;
        RECT 20.950 49.620 21.210 49.880 ;
        RECT 20.310 31.960 20.570 32.220 ;
        RECT 19.690 30.810 19.950 31.070 ;
        RECT 34.270 49.470 34.600 49.800 ;
        RECT 33.640 47.940 33.970 48.270 ;
        RECT 33.080 46.370 33.410 46.700 ;
        RECT 32.460 40.900 32.790 41.230 ;
        RECT 31.830 39.310 32.160 39.640 ;
        RECT 31.210 37.760 31.540 38.090 ;
        RECT 30.610 36.280 30.940 36.610 ;
        RECT 29.970 31.110 30.300 31.440 ;
        RECT 19.250 30.110 19.510 30.370 ;
        RECT 18.800 28.760 19.060 29.020 ;
        RECT 19.270 28.200 19.530 28.460 ;
        RECT 18.800 27.210 19.060 27.470 ;
        RECT 17.310 26.000 17.570 26.260 ;
        RECT 15.100 25.570 15.360 25.830 ;
        RECT 16.190 25.570 16.450 25.830 ;
        RECT 17.320 25.530 17.580 25.790 ;
        RECT 14.550 24.890 14.810 25.150 ;
        RECT 15.650 24.890 15.910 25.150 ;
        RECT 16.750 24.890 17.010 25.150 ;
        RECT 14.550 23.520 14.810 23.780 ;
        RECT 15.650 23.520 15.910 23.780 ;
        RECT 16.750 23.520 17.010 23.780 ;
        RECT 14.000 22.790 14.260 23.050 ;
        RECT 15.100 22.790 15.360 23.050 ;
        RECT 16.190 22.790 16.450 23.050 ;
        RECT 13.990 21.450 14.250 21.710 ;
        RECT 15.100 21.440 15.360 21.700 ;
        RECT 16.190 21.420 16.450 21.680 ;
        RECT 9.900 20.550 10.270 20.920 ;
        RECT 14.550 20.750 14.810 21.010 ;
        RECT 15.650 20.740 15.910 21.000 ;
        RECT 16.740 20.740 17.000 21.000 ;
        RECT 17.440 20.130 17.700 20.490 ;
        RECT 12.890 14.890 13.180 15.180 ;
        RECT 16.710 14.250 16.970 14.510 ;
        RECT 19.280 26.230 19.540 26.490 ;
        RECT 20.470 30.550 20.730 30.810 ;
        RECT 21.120 30.550 21.380 30.810 ;
        RECT 19.950 30.110 20.210 30.370 ;
        RECT 19.970 26.220 20.230 26.480 ;
        RECT 21.630 29.380 21.890 29.640 ;
        RECT 29.300 29.540 29.630 29.870 ;
        RECT 21.550 28.250 21.810 28.510 ;
        RECT 20.950 27.630 21.210 27.890 ;
        RECT 21.560 27.710 21.820 27.970 ;
        RECT 28.680 27.900 29.010 28.230 ;
        RECT 20.450 25.450 20.710 25.710 ;
        RECT 21.610 26.760 21.870 27.020 ;
        RECT 28.000 26.460 28.330 26.790 ;
        RECT 19.710 22.510 19.970 22.930 ;
        RECT 19.670 20.130 19.930 20.490 ;
        RECT 21.160 25.390 21.420 25.650 ;
        RECT 20.290 16.500 20.550 16.830 ;
        RECT 19.260 14.880 19.550 15.170 ;
        RECT 13.400 13.810 13.660 14.070 ;
        RECT 14.500 13.820 14.760 14.080 ;
        RECT 15.590 13.820 15.850 14.080 ;
        RECT 16.720 13.780 16.980 14.040 ;
        RECT 18.100 13.870 18.700 14.470 ;
        RECT 13.950 13.140 14.210 13.400 ;
        RECT 15.050 13.140 15.310 13.400 ;
        RECT 16.150 13.140 16.410 13.400 ;
        RECT 13.950 11.770 14.210 12.030 ;
        RECT 15.050 11.770 15.310 12.030 ;
        RECT 16.150 11.770 16.410 12.030 ;
        RECT 13.400 11.040 13.660 11.300 ;
        RECT 14.500 11.040 14.760 11.300 ;
        RECT 15.590 11.040 15.850 11.300 ;
        RECT 13.390 9.700 13.650 9.960 ;
        RECT 14.500 9.690 14.760 9.950 ;
        RECT 15.590 9.670 15.850 9.930 ;
        RECT 23.960 22.100 24.540 22.810 ;
        RECT 13.950 9.000 14.210 9.260 ;
        RECT 15.050 8.990 15.310 9.250 ;
        RECT 16.140 8.990 16.400 9.250 ;
        RECT 20.880 8.940 21.140 9.280 ;
        RECT 1.970 8.000 2.360 8.390 ;
        RECT 27.970 2.630 28.400 3.060 ;
        RECT 28.620 1.840 29.050 2.270 ;
        RECT 29.290 1.160 29.690 1.560 ;
        RECT 29.120 0.220 29.630 0.730 ;
        RECT 38.860 55.340 39.120 55.600 ;
        RECT 38.860 53.590 39.120 53.850 ;
        RECT 38.860 51.840 39.120 52.100 ;
        RECT 38.860 51.050 39.120 51.310 ;
        RECT 38.860 49.300 39.120 49.560 ;
        RECT 38.860 47.550 39.120 47.810 ;
        RECT 38.860 45.800 39.120 46.060 ;
        RECT 44.680 57.940 44.940 58.200 ;
        RECT 45.720 57.980 45.980 58.240 ;
        RECT 40.960 56.180 41.220 56.440 ;
        RECT 40.960 54.430 41.220 54.690 ;
        RECT 40.960 52.680 41.220 52.940 ;
        RECT 40.960 50.210 41.220 50.470 ;
        RECT 40.960 48.460 41.220 48.720 ;
        RECT 40.960 46.710 41.220 46.970 ;
        RECT 43.000 57.210 43.260 57.470 ;
        RECT 44.680 56.190 44.940 56.450 ;
        RECT 45.720 56.230 45.980 56.490 ;
        RECT 43.000 55.460 43.260 55.720 ;
        RECT 44.680 54.440 44.940 54.700 ;
        RECT 45.720 54.480 45.980 54.740 ;
        RECT 43.000 53.710 43.260 53.970 ;
        RECT 44.680 52.690 44.940 52.950 ;
        RECT 45.720 52.730 45.980 52.990 ;
        RECT 43.000 51.960 43.260 52.220 ;
        RECT 43.000 50.930 43.260 51.190 ;
        RECT 44.680 50.200 44.940 50.460 ;
        RECT 45.720 50.160 45.980 50.420 ;
        RECT 43.000 49.180 43.260 49.440 ;
        RECT 44.680 48.450 44.940 48.710 ;
        RECT 45.720 48.410 45.980 48.670 ;
        RECT 43.000 47.430 43.260 47.690 ;
        RECT 44.680 46.700 44.940 46.960 ;
        RECT 45.720 46.660 45.980 46.920 ;
        RECT 43.000 45.680 43.260 45.940 ;
        RECT 40.960 44.960 41.220 45.220 ;
        RECT 44.680 44.950 44.940 45.210 ;
        RECT 45.720 44.910 45.980 45.170 ;
        RECT 38.860 40.920 39.120 41.180 ;
        RECT 38.860 39.170 39.120 39.430 ;
        RECT 38.860 37.420 39.120 37.680 ;
        RECT 38.860 35.670 39.120 35.930 ;
        RECT 40.960 40.080 41.220 40.340 ;
        RECT 40.960 38.330 41.220 38.590 ;
        RECT 40.960 36.580 41.220 36.840 ;
        RECT 43.000 40.800 43.260 41.060 ;
        RECT 44.680 40.070 44.940 40.330 ;
        RECT 45.720 40.030 45.980 40.290 ;
        RECT 43.000 39.050 43.260 39.310 ;
        RECT 44.680 38.320 44.940 38.580 ;
        RECT 45.720 38.280 45.980 38.540 ;
        RECT 43.000 37.300 43.260 37.560 ;
        RECT 44.680 36.570 44.940 36.830 ;
        RECT 45.720 36.530 45.980 36.790 ;
        RECT 43.000 35.550 43.260 35.810 ;
        RECT 38.820 31.860 39.080 32.120 ;
        RECT 40.960 34.830 41.220 35.090 ;
        RECT 44.680 34.820 44.940 35.080 ;
        RECT 45.720 34.780 45.980 35.040 ;
        RECT 47.980 64.120 48.420 64.560 ;
        RECT 48.880 50.990 49.140 51.250 ;
        RECT 47.790 50.470 48.050 50.730 ;
        RECT 47.790 49.200 48.050 49.460 ;
        RECT 48.880 48.680 49.140 48.940 ;
        RECT 48.880 47.790 49.140 48.050 ;
        RECT 47.790 47.270 48.050 47.530 ;
        RECT 47.790 46.000 48.050 46.260 ;
        RECT 48.880 45.480 49.140 45.740 ;
        RECT 62.380 64.120 62.820 64.560 ;
        RECT 56.630 60.340 56.890 60.600 ;
        RECT 54.750 56.810 55.010 57.070 ;
        RECT 60.220 59.430 60.480 59.690 ;
        RECT 57.090 58.410 57.350 58.670 ;
        RECT 57.510 56.320 57.770 56.580 ;
        RECT 58.570 55.840 58.830 56.100 ;
        RECT 52.250 51.790 52.510 52.050 ;
        RECT 51.290 50.990 51.550 51.250 ;
        RECT 52.100 50.830 52.360 51.090 ;
        RECT 51.160 49.720 51.420 49.980 ;
        RECT 51.160 49.120 51.420 49.380 ;
        RECT 51.290 48.680 51.550 48.940 ;
        RECT 51.290 47.790 51.550 48.050 ;
        RECT 52.100 48.070 52.360 48.330 ;
        RECT 54.290 48.390 54.550 48.650 ;
        RECT 59.360 51.240 59.620 51.500 ;
        RECT 52.250 47.060 52.510 47.320 ;
        RECT 63.390 60.350 63.650 60.610 ;
        RECT 62.950 59.440 63.210 59.700 ;
        RECT 60.210 48.740 60.480 49.010 ;
        RECT 59.390 47.550 59.650 47.810 ;
        RECT 68.180 64.080 68.620 64.520 ;
        RECT 76.510 65.110 76.790 65.550 ;
        RECT 72.730 58.450 73.950 58.710 ;
        RECT 69.490 57.800 69.750 58.060 ;
        RECT 75.820 57.260 76.080 57.520 ;
        RECT 78.160 60.350 78.420 60.610 ;
        RECT 77.270 59.480 77.530 59.740 ;
        RECT 84.680 69.450 85.050 69.820 ;
        RECT 80.830 61.060 81.090 61.330 ;
        RECT 77.270 55.270 77.530 55.530 ;
        RECT 78.290 55.280 78.550 55.540 ;
        RECT 85.500 65.990 85.870 66.360 ;
        RECT 83.140 56.470 83.400 56.730 ;
        RECT 81.040 55.160 81.470 55.590 ;
        RECT 82.750 54.940 83.010 55.200 ;
        RECT 82.040 54.110 82.300 54.370 ;
        RECT 82.740 53.250 83.000 53.510 ;
        RECT 83.140 51.740 83.400 52.000 ;
        RECT 86.270 61.280 86.640 61.650 ;
        RECT 85.130 53.090 85.390 53.350 ;
        RECT 51.290 45.480 51.550 45.740 ;
        RECT 62.530 45.320 62.790 45.580 ;
        RECT 48.860 40.520 49.120 40.780 ;
        RECT 47.770 40.000 48.030 40.260 ;
        RECT 47.770 38.730 48.030 38.990 ;
        RECT 48.860 38.210 49.120 38.470 ;
        RECT 48.860 37.320 49.120 37.580 ;
        RECT 47.770 36.800 48.030 37.060 ;
        RECT 47.770 35.530 48.030 35.790 ;
        RECT 51.270 40.520 51.530 40.780 ;
        RECT 55.670 40.790 55.930 41.050 ;
        RECT 56.850 42.100 57.130 42.380 ;
        RECT 74.530 47.920 74.790 48.180 ;
        RECT 76.490 48.380 76.750 48.640 ;
        RECT 78.240 48.400 78.500 48.660 ;
        RECT 80.940 48.410 81.200 48.670 ;
        RECT 78.390 47.570 78.650 47.830 ;
        RECT 80.890 47.760 81.150 48.020 ;
        RECT 74.680 46.960 74.940 47.220 ;
        RECT 68.230 45.260 68.490 45.520 ;
        RECT 75.620 45.850 75.880 46.110 ;
        RECT 75.620 45.250 75.880 45.510 ;
        RECT 77.280 47.040 77.540 47.300 ;
        RECT 80.890 46.910 81.150 47.170 ;
        RECT 78.450 46.560 78.710 46.820 ;
        RECT 83.190 48.430 83.450 48.690 ;
        RECT 76.560 45.570 76.820 45.830 ;
        RECT 78.010 45.760 78.270 46.020 ;
        RECT 74.680 44.200 74.940 44.460 ;
        RECT 68.230 42.740 68.490 43.000 ;
        RECT 57.610 40.470 57.870 40.730 ;
        RECT 51.270 38.210 51.530 38.470 ;
        RECT 57.610 39.920 57.870 40.180 ;
        RECT 51.270 37.320 51.530 37.580 ;
        RECT 57.610 38.930 57.870 39.190 ;
        RECT 57.610 38.380 57.870 38.640 ;
        RECT 57.610 37.230 57.870 37.490 ;
        RECT 48.860 35.010 49.120 35.270 ;
        RECT 51.270 35.010 51.530 35.270 ;
        RECT 42.960 31.740 43.220 32.000 ;
        RECT 38.820 30.110 39.080 30.370 ;
        RECT 38.820 28.360 39.080 28.620 ;
        RECT 38.820 26.610 39.080 26.870 ;
        RECT 49.480 33.910 49.740 34.320 ;
        RECT 57.610 36.680 57.870 36.940 ;
        RECT 58.530 36.260 58.790 36.520 ;
        RECT 55.000 35.140 55.260 35.400 ;
        RECT 57.610 35.700 57.870 35.960 ;
        RECT 55.000 34.590 55.260 34.850 ;
        RECT 55.000 33.620 55.260 33.880 ;
        RECT 55.000 33.070 55.260 33.330 ;
        RECT 40.920 31.020 41.180 31.280 ;
        RECT 40.920 29.270 41.180 29.530 ;
        RECT 40.920 27.520 41.180 27.780 ;
        RECT 40.920 25.770 41.180 26.030 ;
        RECT 44.640 31.010 44.900 31.270 ;
        RECT 45.680 30.970 45.940 31.230 ;
        RECT 42.960 29.990 43.220 30.250 ;
        RECT 44.640 29.260 44.900 29.520 ;
        RECT 45.680 29.220 45.940 29.480 ;
        RECT 42.960 28.240 43.220 28.500 ;
        RECT 44.640 27.510 44.900 27.770 ;
        RECT 45.680 27.470 45.940 27.730 ;
        RECT 42.960 26.490 43.220 26.750 ;
        RECT 44.640 25.760 44.900 26.020 ;
        RECT 45.680 25.720 45.940 25.980 ;
        RECT 48.890 31.250 49.150 31.510 ;
        RECT 47.800 30.730 48.060 30.990 ;
        RECT 47.800 29.460 48.060 29.720 ;
        RECT 48.890 28.940 49.150 29.200 ;
        RECT 48.890 28.050 49.150 28.310 ;
        RECT 47.800 27.530 48.060 27.790 ;
        RECT 47.800 26.260 48.060 26.520 ;
        RECT 48.890 25.740 49.150 26.000 ;
        RECT 51.300 31.250 51.560 31.510 ;
        RECT 55.000 31.900 55.260 32.160 ;
        RECT 55.000 31.350 55.260 31.610 ;
        RECT 57.610 35.150 57.870 35.410 ;
        RECT 56.040 30.850 56.300 31.110 ;
        RECT 58.250 31.040 58.510 31.300 ;
        RECT 62.460 36.220 62.720 36.480 ;
        RECT 74.530 43.190 74.790 43.450 ;
        RECT 80.940 46.260 81.200 46.520 ;
        RECT 80.940 45.410 81.200 45.670 ;
        RECT 80.890 44.760 81.150 45.020 ;
        RECT 80.890 43.910 81.150 44.170 ;
        RECT 83.240 46.210 83.500 46.470 ;
        RECT 83.230 45.490 83.490 45.750 ;
        RECT 74.200 41.530 74.460 41.790 ;
        RECT 73.110 40.470 73.370 40.730 ;
        RECT 80.940 43.260 81.200 43.520 ;
        RECT 78.670 42.870 78.940 43.130 ;
        RECT 83.150 43.240 83.410 43.500 ;
        RECT 84.690 42.080 85.060 42.450 ;
        RECT 73.110 39.920 73.370 40.180 ;
        RECT 85.460 41.490 85.830 41.860 ;
        RECT 75.070 40.800 75.330 41.060 ;
        RECT 68.260 36.220 68.520 36.480 ;
        RECT 73.110 38.930 73.370 39.190 ;
        RECT 92.820 60.230 93.320 60.730 ;
        RECT 89.600 58.670 90.100 59.170 ;
        RECT 90.550 59.160 91.050 59.660 ;
        RECT 91.630 59.630 92.130 60.130 ;
        RECT 87.150 56.210 87.520 56.580 ;
        RECT 73.110 38.380 73.370 38.640 ;
        RECT 86.200 39.160 86.570 39.530 ;
        RECT 73.110 37.230 73.370 37.490 ;
        RECT 73.110 36.680 73.370 36.940 ;
        RECT 72.190 36.260 72.450 36.520 ;
        RECT 73.110 35.700 73.370 35.960 ;
        RECT 73.110 35.150 73.370 35.410 ;
        RECT 51.300 28.940 51.560 29.200 ;
        RECT 53.880 30.190 54.140 30.450 ;
        RECT 55.000 30.370 55.260 30.630 ;
        RECT 55.000 29.820 55.260 30.080 ;
        RECT 54.960 29.490 55.220 29.750 ;
        RECT 51.300 28.050 51.560 28.310 ;
        RECT 51.300 25.740 51.560 26.000 ;
        RECT 60.060 30.830 60.330 31.090 ;
        RECT 58.230 29.990 58.490 30.250 ;
        RECT 87.130 33.910 87.500 34.320 ;
        RECT 66.330 30.840 66.590 31.100 ;
        RECT 66.480 30.160 66.740 30.420 ;
        RECT 66.480 29.270 66.740 29.530 ;
        RECT 54.940 28.480 55.200 28.740 ;
        RECT 66.330 28.590 66.590 28.850 ;
        RECT 54.510 27.410 54.770 27.670 ;
        RECT 47.300 25.060 47.560 25.320 ;
        RECT 46.760 24.690 47.050 24.980 ;
        RECT 42.320 24.180 42.630 24.490 ;
        RECT 53.910 25.100 54.170 25.360 ;
        RECT 54.890 26.440 55.150 26.700 ;
        RECT 54.940 25.480 55.200 25.740 ;
        RECT 54.940 25.090 55.200 25.350 ;
        RECT 52.510 24.690 52.770 24.950 ;
        RECT 54.480 24.770 54.740 25.030 ;
        RECT 46.130 23.470 46.550 23.890 ;
        RECT 42.280 22.510 42.700 22.930 ;
        RECT 48.190 24.150 48.450 24.410 ;
        RECT 58.230 28.110 58.490 28.370 ;
        RECT 66.330 28.070 66.590 28.330 ;
        RECT 66.480 27.390 66.740 27.650 ;
        RECT 58.100 26.930 58.360 27.190 ;
        RECT 66.480 26.500 66.740 26.760 ;
        RECT 66.330 25.820 66.590 26.080 ;
        RECT 56.720 24.710 56.980 24.970 ;
        RECT 47.600 23.480 47.860 23.740 ;
        RECT 48.690 23.480 48.950 23.740 ;
        RECT 49.790 23.470 50.050 23.730 ;
        RECT 52.630 23.470 52.890 23.730 ;
        RECT 53.730 23.480 53.990 23.740 ;
        RECT 54.820 23.480 55.080 23.740 ;
        RECT 55.520 23.460 55.850 23.790 ;
        RECT 73.760 30.170 74.020 30.430 ;
        RECT 73.240 29.240 73.500 29.500 ;
        RECT 72.770 27.400 73.030 27.660 ;
        RECT 68.610 26.940 68.880 27.210 ;
        RECT 65.560 25.020 65.910 25.370 ;
        RECT 58.710 24.290 58.970 24.550 ;
        RECT 62.750 24.260 63.020 24.530 ;
        RECT 56.670 23.390 57.010 23.730 ;
        RECT 57.410 23.510 57.670 23.770 ;
        RECT 58.500 23.510 58.760 23.770 ;
        RECT 59.600 23.500 59.860 23.760 ;
        RECT 62.440 23.500 62.700 23.760 ;
        RECT 63.540 23.510 63.800 23.770 ;
        RECT 64.630 23.510 64.890 23.770 ;
        RECT 72.270 26.470 72.530 26.730 ;
        RECT 65.600 23.250 65.860 23.570 ;
        RECT 48.150 22.800 48.410 23.060 ;
        RECT 49.240 22.780 49.500 23.040 ;
        RECT 53.180 22.780 53.440 23.040 ;
        RECT 54.270 22.800 54.530 23.060 ;
        RECT 57.960 22.830 58.220 23.090 ;
        RECT 59.050 22.810 59.310 23.070 ;
        RECT 62.990 22.810 63.250 23.070 ;
        RECT 64.080 22.830 64.340 23.090 ;
        RECT 71.590 23.470 71.850 23.810 ;
        RECT 46.810 22.420 47.130 22.740 ;
        RECT 67.020 22.540 67.400 22.920 ;
        RECT 48.150 21.430 48.410 21.690 ;
        RECT 49.240 21.430 49.500 21.690 ;
        RECT 53.180 21.430 53.440 21.690 ;
        RECT 54.270 21.430 54.530 21.690 ;
        RECT 57.960 21.460 58.220 21.720 ;
        RECT 59.050 21.460 59.310 21.720 ;
        RECT 62.990 21.460 63.250 21.720 ;
        RECT 64.080 21.460 64.340 21.720 ;
        RECT 47.590 20.700 47.850 20.960 ;
        RECT 48.690 20.700 48.950 20.960 ;
        RECT 49.790 20.700 50.050 20.960 ;
        RECT 52.630 20.700 52.890 20.960 ;
        RECT 53.730 20.700 53.990 20.960 ;
        RECT 54.830 20.700 55.090 20.960 ;
        RECT 57.400 20.730 57.660 20.990 ;
        RECT 58.500 20.730 58.760 20.990 ;
        RECT 59.600 20.730 59.860 20.990 ;
        RECT 62.440 20.730 62.700 20.990 ;
        RECT 63.540 20.730 63.800 20.990 ;
        RECT 64.640 20.730 64.900 20.990 ;
        RECT 47.590 19.330 47.850 19.590 ;
        RECT 48.690 19.330 48.950 19.590 ;
        RECT 49.790 19.330 50.050 19.590 ;
        RECT 52.630 19.330 52.890 19.590 ;
        RECT 53.730 19.330 53.990 19.590 ;
        RECT 54.830 19.330 55.090 19.590 ;
        RECT 57.400 19.360 57.660 19.620 ;
        RECT 58.500 19.360 58.760 19.620 ;
        RECT 59.600 19.360 59.860 19.620 ;
        RECT 62.440 19.360 62.700 19.620 ;
        RECT 63.540 19.360 63.800 19.620 ;
        RECT 64.640 19.360 64.900 19.620 ;
        RECT 68.820 19.290 69.080 19.550 ;
        RECT 69.920 19.300 70.180 19.560 ;
        RECT 71.010 19.300 71.270 19.560 ;
        RECT 47.020 18.690 47.280 18.950 ;
        RECT 48.150 18.650 48.410 18.910 ;
        RECT 49.240 18.650 49.500 18.910 ;
        RECT 53.180 18.650 53.440 18.910 ;
        RECT 54.270 18.650 54.530 18.910 ;
        RECT 55.400 18.690 55.660 18.950 ;
        RECT 47.030 18.220 47.290 18.480 ;
        RECT 55.390 18.220 55.650 18.480 ;
        RECT 46.910 16.640 47.370 17.100 ;
        RECT 56.830 18.720 57.090 18.980 ;
        RECT 57.960 18.680 58.220 18.940 ;
        RECT 59.050 18.680 59.310 18.940 ;
        RECT 62.990 18.680 63.250 18.940 ;
        RECT 64.080 18.680 64.340 18.940 ;
        RECT 65.210 18.720 65.470 18.980 ;
        RECT 68.260 18.590 68.520 18.850 ;
        RECT 69.370 18.600 69.630 18.860 ;
        RECT 70.460 18.620 70.720 18.880 ;
        RECT 101.630 57.290 102.910 58.570 ;
        RECT 105.950 55.130 106.210 55.560 ;
        RECT 102.120 53.850 102.380 54.270 ;
        RECT 93.350 47.410 93.610 47.670 ;
        RECT 98.120 50.650 98.520 51.050 ;
        RECT 92.730 37.950 93.230 38.450 ;
        RECT 91.650 32.760 92.150 33.230 ;
        RECT 90.520 27.570 91.020 28.070 ;
        RECT 89.470 22.270 89.970 22.770 ;
        RECT 73.740 20.760 74.000 21.260 ;
        RECT 73.200 19.860 73.460 20.360 ;
        RECT 72.730 18.960 72.990 19.460 ;
        RECT 56.840 18.250 57.100 18.510 ;
        RECT 65.200 18.250 65.460 18.510 ;
        RECT 55.290 15.690 55.750 16.150 ;
        RECT 56.720 14.800 57.180 15.260 ;
        RECT 68.270 17.250 68.530 17.510 ;
        RECT 69.370 17.250 69.630 17.510 ;
        RECT 70.460 17.250 70.720 17.510 ;
        RECT 72.250 18.060 72.510 18.560 ;
        RECT 68.820 16.520 69.080 16.780 ;
        RECT 69.920 16.520 70.180 16.780 ;
        RECT 71.020 16.520 71.280 16.780 ;
        RECT 68.820 15.150 69.080 15.410 ;
        RECT 69.920 15.150 70.180 15.410 ;
        RECT 71.020 15.150 71.280 15.410 ;
        RECT 68.270 14.480 68.530 14.740 ;
        RECT 69.370 14.470 69.630 14.730 ;
        RECT 70.460 14.470 70.720 14.730 ;
        RECT 65.110 13.890 65.570 14.350 ;
        RECT 39.040 11.660 39.300 12.780 ;
        RECT 71.590 14.510 71.850 14.770 ;
        RECT 95.710 24.790 96.210 25.290 ;
        RECT 92.840 16.680 93.340 17.180 ;
        RECT 91.650 15.730 92.150 16.190 ;
        RECT 90.520 14.860 91.020 15.320 ;
        RECT 71.580 14.040 71.840 14.300 ;
        RECT 89.590 13.950 90.090 14.410 ;
        RECT 95.130 11.660 96.070 12.780 ;
        RECT 70.920 8.030 71.250 8.360 ;
        RECT 37.360 7.370 37.690 7.700 ;
        RECT 99.100 50.010 99.460 50.370 ;
        RECT 99.150 47.410 99.410 47.670 ;
        RECT 100.020 47.640 100.410 48.030 ;
        RECT 36.740 6.750 37.070 7.080 ;
        RECT 98.180 6.840 98.580 7.240 ;
        RECT 36.110 6.120 36.440 6.450 ;
        RECT 99.090 6.040 99.480 6.430 ;
        RECT 35.510 5.490 35.840 5.820 ;
        RECT 100.850 47.080 101.230 47.340 ;
        RECT 100.020 5.220 100.410 5.610 ;
        RECT 34.870 4.810 35.200 5.140 ;
        RECT 105.420 52.600 105.680 52.860 ;
        RECT 105.570 51.640 105.830 51.900 ;
        RECT 108.570 53.630 108.830 53.890 ;
        RECT 107.400 53.090 107.660 53.350 ;
        RECT 109.130 53.080 109.390 53.340 ;
        RECT 112.900 62.620 113.610 63.330 ;
        RECT 110.840 53.560 111.100 53.820 ;
        RECT 111.850 53.570 112.110 53.830 ;
        RECT 111.830 53.090 112.090 53.350 ;
        RECT 109.920 52.650 110.180 52.910 ;
        RECT 111.490 52.650 111.750 52.910 ;
        RECT 109.280 52.250 109.540 52.510 ;
        RECT 111.780 52.440 112.040 52.700 ;
        RECT 106.510 50.530 106.770 50.790 ;
        RECT 106.510 49.930 106.770 50.190 ;
        RECT 108.170 51.720 108.430 51.980 ;
        RECT 114.080 53.110 114.340 53.370 ;
        RECT 109.340 51.240 109.600 51.500 ;
        RECT 109.920 51.500 110.180 51.760 ;
        RECT 111.490 51.500 111.750 51.760 ;
        RECT 111.780 51.590 112.040 51.850 ;
        RECT 107.450 50.250 107.710 50.510 ;
        RECT 108.570 50.430 108.830 50.780 ;
        RECT 108.900 50.440 109.160 50.700 ;
        RECT 105.570 48.880 105.830 49.140 ;
        RECT 105.420 47.870 105.680 48.130 ;
        RECT 111.830 50.940 112.090 51.200 ;
        RECT 110.840 50.360 111.100 50.850 ;
        RECT 111.850 50.370 112.110 50.840 ;
        RECT 114.130 50.890 114.390 51.150 ;
        RECT 111.830 50.090 112.090 50.350 ;
        RECT 109.920 49.450 110.180 49.710 ;
        RECT 111.490 49.450 111.750 49.710 ;
        RECT 111.780 49.440 112.040 49.700 ;
        RECT 114.120 50.170 114.380 50.430 ;
        RECT 111.780 48.590 112.040 48.850 ;
        RECT 109.920 48.300 110.180 48.560 ;
        RECT 111.490 48.300 111.750 48.560 ;
        RECT 108.570 47.320 108.830 47.580 ;
        RECT 109.540 47.560 109.800 47.820 ;
        RECT 111.830 47.940 112.090 48.200 ;
        RECT 110.840 47.390 111.100 47.650 ;
        RECT 111.850 47.380 112.110 47.640 ;
        RECT 114.040 47.920 114.300 48.180 ;
        RECT 112.710 42.830 113.420 43.540 ;
        RECT 108.510 24.780 109.020 25.290 ;
        RECT 107.720 14.970 107.980 15.230 ;
        RECT 107.720 14.300 107.980 14.560 ;
        RECT 107.880 13.060 108.140 13.320 ;
        RECT 102.940 9.730 103.200 9.990 ;
        RECT 107.880 11.450 108.140 11.710 ;
        RECT 107.870 9.840 108.130 10.100 ;
        RECT 107.880 8.220 108.140 8.480 ;
        RECT 107.870 6.610 108.130 6.870 ;
        RECT 34.270 4.190 34.600 4.520 ;
        RECT 100.840 4.430 101.220 4.810 ;
        RECT 107.460 4.960 107.720 5.220 ;
        RECT 33.670 3.550 34.000 3.880 ;
        RECT 107.870 3.410 108.130 3.670 ;
        RECT 33.090 2.980 33.420 3.310 ;
        RECT 32.510 2.290 32.840 2.620 ;
        RECT 31.860 1.650 32.190 1.980 ;
        RECT 104.630 1.700 104.890 1.960 ;
        RECT 105.570 1.700 105.830 1.960 ;
        RECT 106.520 1.680 106.780 1.940 ;
        RECT 107.830 1.700 108.090 1.960 ;
        RECT 31.220 1.000 31.550 1.340 ;
        RECT 30.640 0.360 31.010 0.730 ;
      LAYER met2 ;
        RECT 20.550 68.100 21.300 68.110 ;
        RECT 20.550 67.800 22.170 68.100 ;
        RECT 20.550 67.630 20.790 67.800 ;
        RECT 21.870 67.580 22.170 67.800 ;
        RECT 12.750 65.150 13.050 65.290 ;
        RECT 12.750 64.830 13.080 65.150 ;
        RECT 13.480 65.140 13.780 65.280 ;
        RECT 12.770 64.820 13.080 64.830 ;
        RECT 13.460 64.820 13.780 65.140 ;
        RECT 13.460 64.810 13.770 64.820 ;
        RECT 40.960 57.420 41.220 58.220 ;
        RECT 44.660 58.200 44.980 58.210 ;
        RECT 44.650 58.190 44.980 58.200 ;
        RECT 45.690 58.190 46.010 58.240 ;
        RECT 44.650 57.990 49.970 58.190 ;
        RECT 44.650 57.940 44.980 57.990 ;
        RECT 45.690 57.980 46.010 57.990 ;
        RECT 44.660 57.920 44.980 57.940 ;
        RECT 49.770 57.490 49.970 57.990 ;
        RECT 75.790 57.490 76.100 57.550 ;
        RECT 42.960 57.420 43.300 57.480 ;
        RECT 40.860 57.200 43.300 57.420 ;
        RECT 49.770 57.290 76.100 57.490 ;
        RECT 75.790 57.230 76.100 57.290 ;
        RECT 54.720 57.020 55.040 57.070 ;
        RECT 49.720 56.820 55.090 57.020 ;
        RECT 40.960 55.670 41.220 56.470 ;
        RECT 44.660 56.450 44.980 56.460 ;
        RECT 44.650 56.440 44.980 56.450 ;
        RECT 45.690 56.440 46.010 56.490 ;
        RECT 49.720 56.440 49.920 56.820 ;
        RECT 54.720 56.810 55.040 56.820 ;
        RECT 57.480 56.580 57.790 56.590 ;
        RECT 57.480 56.550 57.800 56.580 ;
        RECT 44.650 56.240 49.920 56.440 ;
        RECT 50.230 56.350 57.800 56.550 ;
        RECT 44.650 56.190 44.980 56.240 ;
        RECT 45.690 56.230 46.010 56.240 ;
        RECT 44.660 56.170 44.980 56.190 ;
        RECT 42.960 55.670 43.300 55.730 ;
        RECT 40.860 55.450 43.300 55.670 ;
        RECT 40.960 53.920 41.220 54.720 ;
        RECT 44.660 54.700 44.980 54.710 ;
        RECT 44.650 54.690 44.980 54.700 ;
        RECT 45.690 54.690 46.010 54.740 ;
        RECT 50.230 54.690 50.430 56.350 ;
        RECT 57.480 56.320 57.800 56.350 ;
        RECT 57.480 56.310 57.790 56.320 ;
        RECT 58.540 56.070 58.860 56.110 ;
        RECT 44.650 54.490 50.430 54.690 ;
        RECT 50.780 55.870 58.940 56.070 ;
        RECT 44.650 54.440 44.980 54.490 ;
        RECT 45.690 54.480 46.010 54.490 ;
        RECT 44.660 54.420 44.980 54.440 ;
        RECT 42.960 53.920 43.300 53.980 ;
        RECT 40.860 53.700 43.300 53.920 ;
        RECT 18.730 52.390 19.040 52.500 ;
        RECT 18.390 52.200 19.040 52.390 ;
        RECT 18.730 52.170 19.040 52.200 ;
        RECT 40.960 52.170 41.220 52.970 ;
        RECT 44.660 52.950 44.980 52.960 ;
        RECT 44.650 52.940 44.980 52.950 ;
        RECT 45.690 52.940 46.010 52.990 ;
        RECT 50.780 52.940 50.980 55.870 ;
        RECT 58.540 55.830 58.860 55.870 ;
        RECT 105.620 53.450 105.670 53.650 ;
        RECT 109.110 53.370 109.420 53.380 ;
        RECT 108.540 53.360 109.420 53.370 ;
        RECT 108.470 53.120 109.420 53.360 ;
        RECT 109.110 53.050 109.420 53.120 ;
        RECT 44.650 52.740 50.980 52.940 ;
        RECT 105.390 52.890 105.700 52.900 ;
        RECT 44.650 52.690 44.980 52.740 ;
        RECT 45.690 52.730 46.010 52.740 ;
        RECT 84.900 52.710 84.980 52.890 ;
        RECT 96.340 52.710 107.870 52.890 ;
        RECT 44.660 52.670 44.980 52.690 ;
        RECT 105.390 52.570 105.700 52.710 ;
        RECT 105.620 52.470 105.680 52.570 ;
        RECT 109.260 52.510 109.570 52.550 ;
        RECT 109.080 52.260 109.800 52.510 ;
        RECT 42.960 52.170 43.300 52.230 ;
        RECT 18.700 51.970 19.020 52.030 ;
        RECT 18.390 51.780 19.020 51.970 ;
        RECT 40.860 51.950 43.300 52.170 ;
        RECT 18.700 51.710 19.020 51.780 ;
        RECT 78.280 51.640 78.880 52.200 ;
        RECT 87.480 52.030 96.630 52.260 ;
        RECT 109.260 52.220 109.800 52.260 ;
        RECT 109.530 52.150 109.800 52.220 ;
        RECT 96.340 51.930 96.630 52.030 ;
        RECT 104.320 51.930 105.460 52.010 ;
        RECT 96.340 51.810 105.460 51.930 ;
        RECT 96.340 51.730 104.670 51.810 ;
        RECT 96.340 51.720 96.630 51.730 ;
        RECT 18.730 51.400 19.040 51.510 ;
        RECT 18.390 51.210 19.040 51.400 ;
        RECT 59.340 51.490 59.650 51.540 ;
        RECT 59.340 51.480 59.800 51.490 ;
        RECT 59.340 51.300 61.590 51.480 ;
        RECT 59.340 51.210 59.650 51.300 ;
        RECT 81.890 51.210 87.110 51.430 ;
        RECT 18.730 51.180 19.040 51.210 ;
        RECT 18.700 50.980 19.020 51.040 ;
        RECT 40.860 50.980 43.300 51.200 ;
        RECT 18.390 50.790 19.020 50.980 ;
        RECT 18.700 50.720 19.020 50.790 ;
        RECT 40.960 50.180 41.220 50.980 ;
        RECT 42.960 50.920 43.300 50.980 ;
        RECT 105.620 50.760 105.670 50.960 ;
        RECT 105.620 50.250 105.670 50.450 ;
        RECT 18.700 49.990 19.020 50.050 ;
        RECT 18.390 49.800 19.020 49.990 ;
        RECT 112.890 49.860 113.000 50.080 ;
        RECT 18.700 49.730 19.020 49.800 ;
        RECT 40.860 49.230 43.300 49.450 ;
        RECT 105.620 49.270 105.680 49.470 ;
        RECT 40.960 48.430 41.220 49.230 ;
        RECT 42.960 49.170 43.300 49.230 ;
        RECT 77.220 48.690 77.780 48.710 ;
        RECT 78.220 48.690 78.530 48.700 ;
        RECT 77.220 48.440 78.530 48.690 ;
        RECT 74.500 48.210 74.810 48.220 ;
        RECT 65.450 48.030 76.980 48.210 ;
        RECT 77.220 48.170 77.780 48.440 ;
        RECT 78.220 48.370 78.530 48.440 ;
        RECT 74.500 47.890 74.810 48.030 ;
        RECT 80.860 47.980 81.170 48.060 ;
        RECT 59.370 47.770 59.680 47.850 ;
        RECT 78.370 47.830 78.680 47.870 ;
        RECT 40.860 47.480 43.300 47.700 ;
        RECT 59.370 47.560 61.590 47.770 ;
        RECT 59.370 47.520 59.680 47.560 ;
        RECT 40.960 46.680 41.220 47.480 ;
        RECT 42.960 47.420 43.300 47.480 ;
        RECT 62.920 47.430 63.760 47.630 ;
        RECT 78.190 47.580 78.910 47.830 ;
        RECT 80.560 47.770 81.170 47.980 ;
        RECT 84.900 47.840 84.980 48.020 ;
        RECT 80.860 47.730 81.170 47.770 ;
        RECT 78.370 47.540 78.910 47.580 ;
        RECT 78.640 47.470 78.910 47.540 ;
        RECT 74.650 47.190 74.960 47.260 ;
        RECT 77.250 47.190 77.560 47.330 ;
        RECT 63.370 46.960 73.510 47.180 ;
        RECT 47.750 46.210 48.090 46.280 ;
        RECT 47.610 46.160 48.090 46.210 ;
        RECT 47.410 45.980 48.090 46.160 ;
        RECT 63.320 45.990 72.330 46.210 ;
        RECT 40.860 45.730 43.300 45.950 ;
        RECT 40.960 44.930 41.220 45.730 ;
        RECT 42.960 45.670 43.300 45.730 ;
        RECT 44.660 45.210 44.980 45.230 ;
        RECT 44.650 45.160 44.980 45.210 ;
        RECT 45.690 45.160 46.010 45.170 ;
        RECT 47.410 45.160 47.590 45.980 ;
        RECT 48.850 45.690 49.170 45.770 ;
        RECT 51.260 45.710 51.580 45.740 ;
        RECT 51.260 45.690 53.870 45.710 ;
        RECT 48.850 45.530 53.870 45.690 ;
        RECT 48.850 45.500 51.580 45.530 ;
        RECT 48.850 45.450 49.170 45.500 ;
        RECT 51.260 45.480 51.580 45.500 ;
        RECT 44.650 44.960 47.600 45.160 ;
        RECT 44.650 44.950 44.980 44.960 ;
        RECT 44.660 44.940 44.980 44.950 ;
        RECT 45.690 44.910 46.010 44.960 ;
        RECT 53.690 43.340 53.870 45.530 ;
        RECT 62.500 45.550 62.820 45.600 ;
        RECT 62.500 45.300 68.520 45.550 ;
        RECT 68.200 45.230 68.520 45.300 ;
        RECT 63.370 44.210 69.030 44.430 ;
        RECT 62.870 43.910 63.350 43.920 ;
        RECT 62.870 43.670 63.760 43.910 ;
        RECT 68.810 43.880 69.030 44.210 ;
        RECT 72.110 44.380 72.330 45.990 ;
        RECT 73.290 45.760 73.510 46.960 ;
        RECT 74.650 47.000 77.560 47.190 ;
        RECT 80.860 47.160 81.170 47.200 ;
        RECT 74.650 46.970 77.250 47.000 ;
        RECT 74.650 46.930 74.960 46.970 ;
        RECT 80.560 46.950 81.170 47.160 ;
        RECT 78.710 46.900 78.910 46.910 ;
        RECT 78.710 46.820 78.930 46.900 ;
        RECT 80.860 46.870 81.170 46.950 ;
        RECT 78.420 46.800 78.930 46.820 ;
        RECT 78.370 46.560 78.930 46.800 ;
        RECT 78.370 46.550 78.840 46.560 ;
        RECT 78.260 46.050 78.880 46.150 ;
        RECT 87.480 46.120 104.670 46.300 ;
        RECT 87.480 46.100 105.460 46.120 ;
        RECT 77.980 46.010 78.880 46.050 ;
        RECT 77.660 45.770 78.880 46.010 ;
        RECT 104.410 45.920 105.460 46.100 ;
        RECT 73.260 45.720 73.510 45.760 ;
        RECT 77.980 45.720 78.880 45.770 ;
        RECT 73.260 45.080 73.520 45.720 ;
        RECT 78.260 45.620 78.880 45.720 ;
        RECT 73.260 44.870 77.390 45.080 ;
        RECT 80.860 44.980 81.170 45.060 ;
        RECT 77.180 44.730 77.390 44.870 ;
        RECT 80.560 44.770 81.170 44.980 ;
        RECT 80.860 44.730 81.170 44.770 ;
        RECT 77.180 44.520 79.200 44.730 ;
        RECT 74.650 44.430 74.960 44.500 ;
        RECT 74.650 44.380 76.980 44.430 ;
        RECT 72.110 44.220 76.980 44.380 ;
        RECT 72.110 44.160 74.960 44.220 ;
        RECT 80.860 44.160 81.170 44.200 ;
        RECT 80.560 43.950 81.170 44.160 ;
        RECT 73.180 43.880 79.200 43.930 ;
        RECT 68.810 43.720 79.200 43.880 ;
        RECT 80.860 43.870 81.170 43.950 ;
        RECT 68.810 43.660 73.570 43.720 ;
        RECT 74.500 43.340 74.810 43.480 ;
        RECT 53.690 43.160 54.230 43.340 ;
        RECT 74.500 43.330 76.980 43.340 ;
        RECT 65.450 43.180 76.980 43.330 ;
        RECT 74.500 43.160 76.980 43.180 ;
        RECT 74.500 43.150 74.810 43.160 ;
        RECT 68.200 43.010 68.520 43.020 ;
        RECT 78.640 43.010 78.970 43.150 ;
        RECT 68.200 42.850 78.970 43.010 ;
        RECT 68.200 42.840 68.890 42.850 ;
        RECT 68.200 42.720 68.520 42.840 ;
        RECT 40.860 40.850 43.300 41.070 ;
        RECT 40.960 40.050 41.220 40.850 ;
        RECT 42.960 40.790 43.300 40.850 ;
        RECT 48.830 40.760 49.150 40.810 ;
        RECT 51.240 40.760 51.560 40.780 ;
        RECT 48.830 40.740 53.310 40.760 ;
        RECT 53.610 40.740 53.790 40.750 ;
        RECT 48.830 40.630 53.790 40.740 ;
        RECT 57.590 40.630 57.900 40.770 ;
        RECT 73.080 40.630 73.390 40.770 ;
        RECT 48.830 40.590 75.550 40.630 ;
        RECT 48.830 40.570 51.560 40.590 ;
        RECT 48.830 40.490 49.150 40.570 ;
        RECT 51.240 40.520 51.560 40.570 ;
        RECT 53.270 40.560 75.550 40.590 ;
        RECT 53.610 40.450 75.550 40.560 ;
        RECT 57.590 40.440 57.900 40.450 ;
        RECT 73.080 40.440 73.390 40.450 ;
        RECT 44.660 40.330 44.980 40.350 ;
        RECT 44.650 40.280 44.980 40.330 ;
        RECT 45.690 40.280 46.010 40.290 ;
        RECT 44.650 40.080 48.070 40.280 ;
        RECT 57.590 40.200 57.900 40.220 ;
        RECT 73.080 40.200 73.390 40.220 ;
        RECT 44.650 40.070 44.980 40.080 ;
        RECT 44.660 40.060 44.980 40.070 ;
        RECT 45.690 40.030 46.010 40.080 ;
        RECT 47.590 40.050 48.070 40.080 ;
        RECT 47.730 39.980 48.070 40.050 ;
        RECT 55.430 40.190 57.990 40.200 ;
        RECT 72.990 40.190 75.550 40.200 ;
        RECT 55.430 40.020 75.550 40.190 ;
        RECT 57.590 40.010 73.390 40.020 ;
        RECT 57.590 39.890 57.900 40.010 ;
        RECT 73.080 39.890 73.390 40.010 ;
        RECT 40.860 39.100 43.300 39.320 ;
        RECT 40.960 38.300 41.220 39.100 ;
        RECT 42.960 39.040 43.300 39.100 ;
        RECT 47.730 38.940 48.070 39.010 ;
        RECT 47.590 38.890 48.070 38.940 ;
        RECT 47.390 38.880 48.070 38.890 ;
        RECT 47.370 38.710 48.070 38.880 ;
        RECT 44.660 38.580 44.980 38.600 ;
        RECT 44.650 38.530 44.980 38.580 ;
        RECT 45.690 38.530 46.010 38.540 ;
        RECT 47.370 38.530 47.570 38.710 ;
        RECT 57.590 38.660 57.900 38.670 ;
        RECT 73.080 38.660 73.390 38.670 ;
        RECT 44.650 38.330 47.570 38.530 ;
        RECT 53.350 38.500 75.550 38.660 ;
        RECT 48.830 38.420 49.150 38.500 ;
        RECT 51.310 38.480 75.550 38.500 ;
        RECT 51.310 38.470 53.530 38.480 ;
        RECT 51.240 38.420 53.530 38.470 ;
        RECT 48.830 38.340 53.530 38.420 ;
        RECT 57.590 38.340 57.900 38.480 ;
        RECT 73.080 38.340 73.390 38.480 ;
        RECT 44.650 38.320 44.980 38.330 ;
        RECT 44.660 38.310 44.980 38.320 ;
        RECT 45.690 38.280 46.010 38.330 ;
        RECT 48.830 38.230 51.560 38.340 ;
        RECT 52.040 38.330 53.530 38.340 ;
        RECT 52.740 38.320 53.530 38.330 ;
        RECT 48.830 38.180 49.150 38.230 ;
        RECT 51.240 38.210 51.560 38.230 ;
        RECT 40.860 37.350 43.300 37.570 ;
        RECT 40.960 36.550 41.220 37.350 ;
        RECT 42.960 37.290 43.300 37.350 ;
        RECT 48.830 37.560 49.150 37.610 ;
        RECT 51.240 37.560 51.560 37.580 ;
        RECT 48.830 37.540 51.560 37.560 ;
        RECT 48.830 37.530 53.550 37.540 ;
        RECT 48.830 37.390 53.560 37.530 ;
        RECT 57.590 37.390 57.900 37.530 ;
        RECT 73.080 37.390 73.390 37.530 ;
        RECT 48.830 37.380 75.550 37.390 ;
        RECT 48.830 37.370 51.560 37.380 ;
        RECT 48.830 37.290 49.150 37.370 ;
        RECT 51.240 37.320 51.560 37.370 ;
        RECT 53.380 37.210 75.550 37.380 ;
        RECT 57.590 37.200 57.900 37.210 ;
        RECT 73.080 37.200 73.390 37.210 ;
        RECT 47.590 37.060 48.070 37.080 ;
        RECT 44.660 36.830 44.980 36.850 ;
        RECT 44.650 36.780 44.980 36.830 ;
        RECT 45.690 36.780 46.010 36.790 ;
        RECT 47.320 36.780 48.070 37.060 ;
        RECT 57.590 36.960 57.900 36.980 ;
        RECT 73.080 36.960 73.390 36.980 ;
        RECT 55.430 36.780 75.550 36.960 ;
        RECT 44.650 36.730 47.810 36.780 ;
        RECT 44.650 36.580 47.670 36.730 ;
        RECT 57.590 36.650 57.900 36.780 ;
        RECT 73.080 36.650 73.390 36.780 ;
        RECT 44.650 36.570 44.980 36.580 ;
        RECT 44.660 36.560 44.980 36.570 ;
        RECT 45.690 36.530 46.010 36.580 ;
        RECT 58.500 36.470 58.820 36.530 ;
        RECT 62.430 36.470 62.750 36.480 ;
        RECT 68.230 36.470 68.550 36.480 ;
        RECT 72.160 36.470 72.480 36.530 ;
        RECT 58.500 36.290 72.480 36.470 ;
        RECT 58.500 36.240 58.820 36.290 ;
        RECT 62.430 36.220 62.750 36.290 ;
        RECT 68.230 36.220 68.550 36.290 ;
        RECT 72.160 36.240 72.480 36.290 ;
        RECT 57.590 35.860 57.900 35.990 ;
        RECT 73.080 35.860 73.390 35.990 ;
        RECT 40.860 35.600 43.300 35.820 ;
        RECT 47.730 35.740 48.070 35.810 ;
        RECT 40.960 34.800 41.220 35.600 ;
        RECT 42.960 35.540 43.300 35.600 ;
        RECT 47.360 35.510 48.070 35.740 ;
        RECT 55.430 35.680 75.550 35.860 ;
        RECT 57.590 35.660 57.900 35.680 ;
        RECT 73.080 35.660 73.390 35.680 ;
        RECT 44.660 35.080 44.980 35.100 ;
        RECT 44.650 35.030 44.980 35.080 ;
        RECT 45.690 35.030 46.010 35.040 ;
        RECT 47.360 35.030 47.560 35.510 ;
        RECT 54.980 35.430 55.290 35.440 ;
        RECT 57.590 35.430 57.900 35.440 ;
        RECT 73.080 35.430 73.390 35.440 ;
        RECT 53.340 35.300 75.550 35.430 ;
        RECT 44.650 34.830 47.560 35.030 ;
        RECT 48.830 35.220 49.150 35.300 ;
        RECT 51.240 35.240 51.560 35.270 ;
        RECT 52.820 35.260 75.550 35.300 ;
        RECT 52.820 35.250 57.900 35.260 ;
        RECT 52.820 35.240 55.290 35.250 ;
        RECT 51.240 35.220 55.290 35.240 ;
        RECT 48.830 35.120 55.290 35.220 ;
        RECT 48.830 35.060 53.540 35.120 ;
        RECT 54.980 35.110 55.290 35.120 ;
        RECT 57.590 35.110 57.900 35.250 ;
        RECT 73.080 35.250 75.550 35.260 ;
        RECT 73.080 35.110 73.390 35.250 ;
        RECT 48.830 35.030 51.560 35.060 ;
        RECT 48.830 34.980 49.150 35.030 ;
        RECT 51.240 35.010 51.560 35.030 ;
        RECT 54.980 34.870 55.290 34.890 ;
        RECT 44.650 34.820 44.980 34.830 ;
        RECT 44.660 34.810 44.980 34.820 ;
        RECT 45.690 34.780 46.010 34.830 ;
        RECT 52.820 34.690 62.890 34.870 ;
        RECT 54.980 34.680 62.890 34.690 ;
        RECT 54.980 34.560 55.290 34.680 ;
        RECT 54.980 32.070 55.290 32.200 ;
        RECT 54.980 32.060 55.410 32.070 ;
        RECT 40.820 31.790 43.260 32.010 ;
        RECT 52.820 31.900 55.410 32.060 ;
        RECT 52.820 31.880 55.290 31.900 ;
        RECT 54.980 31.870 55.290 31.880 ;
        RECT 40.920 30.990 41.180 31.790 ;
        RECT 42.920 31.730 43.260 31.790 ;
        RECT 54.980 31.630 55.290 31.650 ;
        RECT 48.860 31.490 49.180 31.540 ;
        RECT 51.270 31.490 51.590 31.510 ;
        RECT 52.820 31.490 62.120 31.630 ;
        RECT 48.860 31.460 62.120 31.490 ;
        RECT 62.420 31.490 62.890 31.650 ;
        RECT 62.420 31.480 62.880 31.490 ;
        RECT 48.860 31.450 55.380 31.460 ;
        RECT 48.860 31.320 53.470 31.450 ;
        RECT 54.980 31.320 55.290 31.450 ;
        RECT 48.860 31.300 51.590 31.320 ;
        RECT 53.160 31.300 53.470 31.320 ;
        RECT 44.620 31.270 44.940 31.290 ;
        RECT 44.610 31.220 44.940 31.270 ;
        RECT 45.650 31.220 45.970 31.230 ;
        RECT 48.860 31.220 49.180 31.300 ;
        RECT 51.270 31.250 51.590 31.300 ;
        RECT 44.610 31.020 47.690 31.220 ;
        RECT 53.290 31.120 55.640 31.300 ;
        RECT 44.610 31.010 44.940 31.020 ;
        RECT 44.620 31.000 44.940 31.010 ;
        RECT 45.650 30.970 45.970 31.020 ;
        RECT 47.490 31.010 47.690 31.020 ;
        RECT 47.490 30.780 48.100 31.010 ;
        RECT 47.760 30.710 48.100 30.780 ;
        RECT 19.920 30.330 20.230 30.400 ;
        RECT 19.920 30.110 22.080 30.330 ;
        RECT 19.920 30.070 20.230 30.110 ;
        RECT 40.820 30.040 43.260 30.260 ;
        RECT 21.600 29.610 21.920 29.670 ;
        RECT 21.600 29.400 22.080 29.610 ;
        RECT 21.600 29.350 21.920 29.400 ;
        RECT 40.920 29.240 41.180 30.040 ;
        RECT 42.920 29.980 43.260 30.040 ;
        RECT 47.760 29.670 48.100 29.740 ;
        RECT 47.620 29.630 48.100 29.670 ;
        RECT 44.620 29.520 44.940 29.540 ;
        RECT 44.610 29.470 44.940 29.520 ;
        RECT 45.650 29.470 45.970 29.480 ;
        RECT 47.480 29.470 48.100 29.630 ;
        RECT 54.930 29.490 55.250 29.760 ;
        RECT 44.610 29.440 48.100 29.470 ;
        RECT 44.610 29.270 47.800 29.440 ;
        RECT 44.610 29.260 44.940 29.270 ;
        RECT 44.620 29.250 44.940 29.260 ;
        RECT 45.650 29.220 45.970 29.270 ;
        RECT 53.270 29.230 55.460 29.350 ;
        RECT 48.860 29.150 49.180 29.230 ;
        RECT 51.340 29.200 55.460 29.230 ;
        RECT 51.270 29.170 55.460 29.200 ;
        RECT 51.270 29.150 53.450 29.170 ;
        RECT 48.860 29.070 53.450 29.150 ;
        RECT 48.860 28.960 51.590 29.070 ;
        RECT 52.070 29.060 53.450 29.070 ;
        RECT 52.770 29.050 53.450 29.060 ;
        RECT 48.860 28.910 49.180 28.960 ;
        RECT 51.270 28.940 51.590 28.960 ;
        RECT 53.130 29.020 53.450 29.050 ;
        RECT 53.130 28.940 53.310 29.020 ;
        RECT 58.160 29.010 58.390 29.020 ;
        RECT 58.160 28.980 65.730 29.010 ;
        RECT 58.160 28.810 65.790 28.980 ;
        RECT 66.300 28.810 66.610 28.890 ;
        RECT 54.910 28.710 55.230 28.740 ;
        RECT 58.160 28.710 58.400 28.810 ;
        RECT 54.910 28.530 58.400 28.710 ;
        RECT 65.600 28.610 66.610 28.810 ;
        RECT 66.200 28.600 66.610 28.610 ;
        RECT 66.300 28.560 66.610 28.600 ;
        RECT 54.910 28.510 58.320 28.530 ;
        RECT 40.820 28.290 43.260 28.510 ;
        RECT 54.910 28.480 55.230 28.510 ;
        RECT 40.920 27.490 41.180 28.290 ;
        RECT 42.920 28.230 43.260 28.290 ;
        RECT 48.860 28.290 49.180 28.340 ;
        RECT 58.200 28.330 58.520 28.370 ;
        RECT 58.200 28.310 65.750 28.330 ;
        RECT 66.300 28.320 66.610 28.360 ;
        RECT 66.200 28.310 66.610 28.320 ;
        RECT 51.270 28.290 51.590 28.310 ;
        RECT 48.860 28.270 51.590 28.290 ;
        RECT 48.860 28.110 53.380 28.270 ;
        RECT 58.200 28.110 66.610 28.310 ;
        RECT 48.860 28.100 51.590 28.110 ;
        RECT 48.860 28.020 49.180 28.100 ;
        RECT 51.270 28.050 51.590 28.100 ;
        RECT 53.200 28.060 53.380 28.110 ;
        RECT 58.300 28.100 58.620 28.110 ;
        RECT 53.200 27.880 55.460 28.060 ;
        RECT 66.300 28.030 66.610 28.110 ;
        RECT 44.620 27.770 44.940 27.790 ;
        RECT 44.610 27.720 44.940 27.770 ;
        RECT 45.650 27.720 45.970 27.730 ;
        RECT 47.620 27.720 48.100 27.810 ;
        RECT 44.610 27.520 48.100 27.720 ;
        RECT 44.610 27.510 44.940 27.520 ;
        RECT 44.620 27.500 44.940 27.510 ;
        RECT 45.650 27.470 45.970 27.520 ;
        RECT 47.560 27.510 48.100 27.520 ;
        RECT 54.480 27.650 54.800 27.690 ;
        RECT 47.560 27.430 47.850 27.510 ;
        RECT 54.480 27.370 55.090 27.650 ;
        RECT 54.890 27.150 55.090 27.370 ;
        RECT 58.070 27.150 58.390 27.190 ;
        RECT 21.580 27.000 21.900 27.050 ;
        RECT 21.580 26.790 22.080 27.000 ;
        RECT 54.890 26.950 58.440 27.150 ;
        RECT 68.580 27.130 68.910 27.220 ;
        RECT 62.230 26.960 68.910 27.130 ;
        RECT 58.070 26.930 58.390 26.950 ;
        RECT 68.580 26.930 68.910 26.960 ;
        RECT 21.580 26.730 21.900 26.790 ;
        RECT 40.820 26.540 43.260 26.760 ;
        RECT 47.540 26.550 47.840 26.590 ;
        RECT 19.940 26.440 20.250 26.510 ;
        RECT 17.290 25.960 17.900 26.290 ;
        RECT 19.940 26.230 22.080 26.440 ;
        RECT 19.940 26.180 20.250 26.230 ;
        RECT 17.300 25.470 17.900 25.960 ;
        RECT 40.920 25.740 41.180 26.540 ;
        RECT 42.920 26.480 43.260 26.540 ;
        RECT 47.530 26.540 47.840 26.550 ;
        RECT 47.530 26.240 48.100 26.540 ;
        RECT 54.860 26.410 55.170 26.740 ;
        RECT 44.620 26.020 44.940 26.040 ;
        RECT 44.610 25.970 44.940 26.020 ;
        RECT 45.650 25.970 45.970 25.980 ;
        RECT 47.530 25.970 47.730 26.240 ;
        RECT 44.610 25.770 47.730 25.970 ;
        RECT 48.860 25.950 49.180 26.030 ;
        RECT 51.270 25.970 51.590 26.000 ;
        RECT 53.440 25.970 55.460 26.100 ;
        RECT 66.300 26.060 66.610 26.120 ;
        RECT 65.750 26.050 66.610 26.060 ;
        RECT 51.270 25.950 55.460 25.970 ;
        RECT 48.860 25.920 55.460 25.950 ;
        RECT 48.860 25.790 53.620 25.920 ;
        RECT 58.170 25.830 66.610 26.050 ;
        RECT 58.170 25.820 65.760 25.830 ;
        RECT 58.170 25.810 58.940 25.820 ;
        RECT 44.610 25.760 44.940 25.770 ;
        RECT 44.620 25.750 44.940 25.760 ;
        RECT 45.650 25.720 45.970 25.770 ;
        RECT 48.860 25.760 51.590 25.790 ;
        RECT 48.860 25.710 49.180 25.760 ;
        RECT 51.270 25.740 51.590 25.760 ;
        RECT 54.910 25.770 55.220 25.780 ;
        RECT 54.910 25.640 55.270 25.770 ;
        RECT 58.170 25.640 58.410 25.810 ;
        RECT 66.300 25.790 66.610 25.830 ;
        RECT 54.910 25.400 58.410 25.640 ;
        RECT 54.910 25.250 55.230 25.400 ;
        RECT 65.530 25.270 65.940 25.380 ;
        RECT 58.560 25.250 65.940 25.270 ;
        RECT 54.910 25.110 65.940 25.250 ;
        RECT 54.910 25.080 55.230 25.110 ;
        RECT 58.480 25.040 65.940 25.110 ;
        RECT 54.470 25.030 54.750 25.040 ;
        RECT 54.450 24.940 54.770 25.030 ;
        RECT 65.530 25.010 65.940 25.040 ;
        RECT 56.690 24.940 57.010 24.970 ;
        RECT 54.420 24.780 57.010 24.940 ;
        RECT 54.450 24.770 54.770 24.780 ;
        RECT 54.470 24.760 54.750 24.770 ;
        RECT 56.690 24.710 57.010 24.780 ;
        RECT 56.710 24.700 56.990 24.710 ;
        RECT 55.490 23.790 55.870 23.820 ;
        RECT 56.840 23.810 59.900 23.820 ;
        RECT 52.590 23.450 55.870 23.790 ;
        RECT 56.750 23.730 59.900 23.810 ;
        RECT 52.610 23.440 52.920 23.450 ;
        RECT 55.420 23.430 55.870 23.450 ;
        RECT 56.640 23.480 59.900 23.730 ;
        RECT 62.400 23.810 65.460 23.820 ;
        RECT 71.570 23.810 71.870 23.830 ;
        RECT 62.400 23.590 65.550 23.810 ;
        RECT 62.400 23.480 65.890 23.590 ;
        RECT 55.420 21.000 55.740 23.430 ;
        RECT 56.640 23.390 57.070 23.480 ;
        RECT 59.570 23.470 59.880 23.480 ;
        RECT 62.420 23.470 62.730 23.480 ;
        RECT 52.580 20.670 55.740 21.000 ;
        RECT 55.420 19.630 55.740 20.670 ;
        RECT 52.580 19.310 55.740 19.630 ;
        RECT 56.750 21.030 57.070 23.390 ;
        RECT 65.230 23.230 65.890 23.480 ;
        RECT 70.860 23.470 71.880 23.810 ;
        RECT 71.570 23.450 71.880 23.470 ;
        RECT 65.230 21.030 65.550 23.230 ;
        RECT 66.980 22.510 67.430 22.940 ;
        RECT 56.750 20.700 59.910 21.030 ;
        RECT 62.390 20.700 65.550 21.030 ;
        RECT 56.750 19.660 57.070 20.700 ;
        RECT 65.230 19.660 65.550 20.700 ;
        RECT 56.750 19.340 59.910 19.660 ;
        RECT 62.390 19.340 65.550 19.660 ;
        RECT 57.370 19.330 57.680 19.340 ;
        RECT 58.470 19.330 58.780 19.340 ;
        RECT 59.570 19.330 59.880 19.340 ;
        RECT 62.420 19.330 62.730 19.340 ;
        RECT 63.520 19.330 63.830 19.340 ;
        RECT 64.620 19.330 64.930 19.340 ;
        RECT 52.610 19.300 52.920 19.310 ;
        RECT 53.710 19.300 54.020 19.310 ;
        RECT 54.810 19.300 55.120 19.310 ;
        RECT 0.590 4.970 1.860 6.850 ;
        RECT 0.660 0.220 1.930 2.100 ;
        RECT 104.600 1.670 104.920 1.990 ;
        RECT 105.540 1.670 105.860 1.990 ;
      LAYER via2 ;
        RECT 78.410 51.750 78.750 52.090 ;
        RECT 77.340 48.270 77.670 48.620 ;
        RECT 78.430 45.700 78.770 46.060 ;
  END
END sky130_hilas_TopLevelTextStructure

MACRO sky130_hilas_pFETLarge
  CLASS CORE ;
  FOREIGN sky130_hilas_pFETLarge ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.640 BY 5.990 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA 5.476200 ;
    ANTENNADIFFAREA 1.032200 ;
    PORT
      LAYER met2 ;
        RECT 0.430 0.830 0.740 0.960 ;
        RECT 0.000 0.630 0.740 0.830 ;
        RECT 0.000 0.490 0.600 0.630 ;
        RECT 0.000 0.160 0.750 0.490 ;
        RECT 0.000 0.010 0.600 0.160 ;
    END
  END GATE
  PIN SOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 2.622000 ;
    PORT
      LAYER met2 ;
        RECT 1.010 5.610 1.320 5.750 ;
        RECT 2.100 5.610 2.410 5.750 ;
        RECT 3.200 5.610 3.510 5.740 ;
        RECT 0.330 5.600 3.510 5.610 ;
        RECT 0.240 5.410 3.510 5.600 ;
        RECT 0.240 5.270 3.390 5.410 ;
        RECT 0.240 2.820 0.560 5.270 ;
        RECT 1.000 2.820 1.310 2.970 ;
        RECT 2.100 2.820 2.410 2.970 ;
        RECT 3.200 2.820 3.510 2.970 ;
        RECT 0.240 2.640 3.510 2.820 ;
        RECT 0.240 2.490 3.400 2.640 ;
        RECT 0.240 1.450 0.560 2.490 ;
        RECT 1.000 1.450 1.310 1.600 ;
        RECT 2.100 1.450 2.410 1.600 ;
        RECT 3.200 1.450 3.510 1.600 ;
        RECT 0.240 1.270 3.510 1.450 ;
        RECT 0.240 1.130 3.400 1.270 ;
    END
  END SOURCE
  PIN DRAIN
    USE ANALOG ;
    ANTENNADIFFAREA 1.334000 ;
    PORT
      LAYER met2 ;
        RECT 1.560 4.890 1.870 5.070 ;
        RECT 2.650 4.890 2.960 5.050 ;
        RECT 3.760 4.890 4.070 5.040 ;
        RECT 1.430 4.590 4.370 4.890 ;
        RECT 3.620 4.550 4.370 4.590 ;
        RECT 3.990 4.420 4.370 4.550 ;
        RECT 4.020 3.700 4.370 4.420 ;
        RECT 1.560 3.550 1.870 3.700 ;
        RECT 2.650 3.550 2.960 3.700 ;
        RECT 3.750 3.550 4.370 3.700 ;
        RECT 1.420 3.220 4.370 3.550 ;
        RECT 4.020 0.930 4.370 3.220 ;
        RECT 1.560 0.780 1.870 0.920 ;
        RECT 2.650 0.780 2.960 0.920 ;
        RECT 3.750 0.780 4.370 0.930 ;
        RECT 1.430 0.460 4.370 0.780 ;
        RECT 1.430 0.450 4.140 0.460 ;
    END
  END DRAIN
  PIN WELL
    USE ANALOG ;
    ANTENNADIFFAREA 0.213200 ;
    PORT
      LAYER nwell ;
        RECT 4.020 0.180 4.640 5.880 ;
      LAYER met1 ;
        RECT 4.140 5.790 4.400 5.990 ;
        RECT 4.140 4.980 4.450 5.790 ;
        RECT 4.140 0.000 4.400 4.980 ;
    END
  END WELL
  OBS
      LAYER nwell ;
        RECT 0.000 0.490 2.700 5.990 ;
        RECT 3.640 3.060 3.650 3.100 ;
      LAYER li1 ;
        RECT 0.100 3.460 0.270 5.960 ;
        RECT 0.650 3.460 0.820 5.960 ;
        RECT 1.200 5.710 1.370 5.960 ;
        RECT 1.020 5.450 1.370 5.710 ;
        RECT 1.200 3.460 1.370 5.450 ;
        RECT 1.750 5.030 1.920 5.960 ;
        RECT 2.300 5.710 2.470 5.960 ;
        RECT 2.110 5.450 2.470 5.710 ;
        RECT 1.570 4.770 1.920 5.030 ;
        RECT 1.750 3.660 1.920 4.770 ;
        RECT 1.570 3.460 1.920 3.660 ;
        RECT 2.300 3.460 2.470 5.450 ;
        RECT 3.210 5.660 3.530 5.700 ;
        RECT 3.210 5.470 3.540 5.660 ;
        RECT 3.210 5.440 3.530 5.470 ;
        RECT 2.660 4.970 2.980 5.010 ;
        RECT 2.660 4.780 2.990 4.970 ;
        RECT 3.770 4.960 4.090 5.000 ;
        RECT 2.660 4.750 2.980 4.780 ;
        RECT 3.770 4.770 4.100 4.960 ;
        RECT 4.250 4.920 4.420 5.680 ;
        RECT 3.770 4.740 4.090 4.770 ;
        RECT 2.660 3.620 2.980 3.660 ;
        RECT 3.760 3.620 4.080 3.660 ;
        RECT 1.570 3.430 1.900 3.460 ;
        RECT 2.660 3.430 2.990 3.620 ;
        RECT 3.760 3.430 4.090 3.620 ;
        RECT 1.570 3.400 1.890 3.430 ;
        RECT 2.660 3.400 2.980 3.430 ;
        RECT 3.760 3.400 4.080 3.430 ;
        RECT 0.960 3.160 1.120 3.190 ;
        RECT 0.100 1.020 0.270 3.130 ;
        RECT 0.650 1.020 0.820 3.130 ;
        RECT 0.960 2.930 1.130 3.160 ;
        RECT 1.510 3.150 1.670 3.190 ;
        RECT 1.200 2.930 1.370 3.130 ;
        RECT 0.960 2.810 1.370 2.930 ;
        RECT 1.510 2.820 1.680 3.150 ;
        RECT 1.510 2.810 1.670 2.820 ;
        RECT 1.010 2.670 1.370 2.810 ;
        RECT 1.200 1.560 1.370 2.670 ;
        RECT 1.010 1.300 1.370 1.560 ;
        RECT 0.100 0.630 0.820 1.020 ;
        RECT 1.200 0.630 1.370 1.300 ;
        RECT 1.750 0.880 1.920 3.130 ;
        RECT 2.060 2.930 2.230 3.220 ;
        RECT 2.610 3.150 2.770 3.190 ;
        RECT 3.160 3.150 3.320 3.190 ;
        RECT 3.710 3.170 3.870 3.190 ;
        RECT 2.300 2.930 2.470 3.130 ;
        RECT 2.060 2.810 2.470 2.930 ;
        RECT 2.610 2.820 2.780 3.150 ;
        RECT 3.160 2.930 3.330 3.150 ;
        RECT 3.160 2.890 3.530 2.930 ;
        RECT 2.610 2.810 2.770 2.820 ;
        RECT 3.160 2.810 3.540 2.890 ;
        RECT 3.710 2.820 3.880 3.170 ;
        RECT 3.710 2.810 3.870 2.820 ;
        RECT 2.110 2.670 2.470 2.810 ;
        RECT 3.210 2.700 3.540 2.810 ;
        RECT 3.210 2.670 3.530 2.700 ;
        RECT 2.300 1.560 2.470 2.670 ;
        RECT 2.110 1.300 2.470 1.560 ;
        RECT 3.210 1.520 3.530 1.560 ;
        RECT 3.210 1.330 3.540 1.520 ;
        RECT 3.210 1.300 3.530 1.330 ;
        RECT 1.570 0.630 1.920 0.880 ;
        RECT 2.300 0.630 2.470 1.300 ;
        RECT 2.660 0.840 2.980 0.880 ;
        RECT 3.760 0.850 4.080 0.890 ;
        RECT 2.660 0.650 2.990 0.840 ;
        RECT 3.760 0.660 4.090 0.850 ;
        RECT 0.200 0.450 0.710 0.630 ;
        RECT 1.570 0.620 1.890 0.630 ;
        RECT 2.660 0.620 2.980 0.650 ;
        RECT 3.760 0.630 4.080 0.660 ;
        RECT 0.200 0.410 0.770 0.450 ;
        RECT 0.200 0.220 0.780 0.410 ;
        RECT 0.200 0.190 0.770 0.220 ;
        RECT 0.200 0.010 0.710 0.190 ;
      LAYER mcon ;
        RECT 1.080 5.490 1.250 5.660 ;
        RECT 2.170 5.490 2.340 5.660 ;
        RECT 1.630 4.810 1.800 4.980 ;
        RECT 1.630 3.440 1.800 3.610 ;
        RECT 3.270 5.480 3.440 5.650 ;
        RECT 4.250 5.510 4.420 5.680 ;
        RECT 4.250 5.150 4.420 5.320 ;
        RECT 2.720 4.790 2.890 4.960 ;
        RECT 3.830 4.780 4.000 4.950 ;
        RECT 2.720 3.440 2.890 3.610 ;
        RECT 3.820 3.440 3.990 3.610 ;
        RECT 1.070 2.710 1.240 2.880 ;
        RECT 1.070 1.340 1.240 1.510 ;
        RECT 0.500 0.700 0.670 0.870 ;
        RECT 2.170 2.710 2.340 2.880 ;
        RECT 3.270 2.710 3.440 2.880 ;
        RECT 2.170 1.340 2.340 1.510 ;
        RECT 3.270 1.340 3.440 1.510 ;
        RECT 1.630 0.660 1.800 0.830 ;
        RECT 2.720 0.660 2.890 0.830 ;
        RECT 3.820 0.670 3.990 0.840 ;
        RECT 0.510 0.230 0.680 0.400 ;
      LAYER met1 ;
        RECT 1.010 5.420 1.330 5.740 ;
        RECT 2.100 5.420 2.420 5.740 ;
        RECT 3.200 5.410 3.520 5.730 ;
        RECT 1.560 4.740 1.880 5.060 ;
        RECT 2.650 4.720 2.970 5.040 ;
        RECT 3.760 4.710 4.080 5.030 ;
        RECT 1.560 3.370 1.880 3.690 ;
        RECT 2.650 3.370 2.970 3.690 ;
        RECT 3.750 3.370 4.070 3.690 ;
        RECT 1.000 2.640 1.320 2.960 ;
        RECT 2.100 2.640 2.420 2.960 ;
        RECT 3.200 2.640 3.520 2.960 ;
        RECT 1.000 1.270 1.320 1.590 ;
        RECT 2.100 1.270 2.420 1.590 ;
        RECT 3.200 1.270 3.520 1.590 ;
        RECT 0.430 0.630 0.750 0.950 ;
        RECT 1.560 0.590 1.880 0.910 ;
        RECT 2.650 0.590 2.970 0.910 ;
        RECT 3.750 0.600 4.070 0.920 ;
        RECT 0.440 0.160 0.760 0.480 ;
      LAYER via ;
        RECT 1.040 5.450 1.300 5.710 ;
        RECT 2.130 5.450 2.390 5.710 ;
        RECT 3.230 5.440 3.490 5.700 ;
        RECT 1.590 4.770 1.850 5.030 ;
        RECT 2.680 4.750 2.940 5.010 ;
        RECT 3.790 4.740 4.050 5.000 ;
        RECT 1.590 3.400 1.850 3.660 ;
        RECT 2.680 3.400 2.940 3.660 ;
        RECT 3.780 3.400 4.040 3.660 ;
        RECT 1.030 2.670 1.290 2.930 ;
        RECT 2.130 2.670 2.390 2.930 ;
        RECT 3.230 2.670 3.490 2.930 ;
        RECT 1.030 1.300 1.290 1.560 ;
        RECT 2.130 1.300 2.390 1.560 ;
        RECT 3.230 1.300 3.490 1.560 ;
        RECT 0.460 0.660 0.720 0.920 ;
        RECT 1.590 0.620 1.850 0.880 ;
        RECT 2.680 0.620 2.940 0.880 ;
        RECT 3.780 0.630 4.040 0.890 ;
        RECT 0.470 0.190 0.730 0.450 ;
  END
END sky130_hilas_pFETLarge

MACRO sky130_hilas_VinjInv2
  CLASS CORE ;
  FOREIGN sky130_hilas_VinjInv2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.610 BY 1.640 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 0.000 0.000 1.980 1.640 ;
      LAYER li1 ;
        RECT 0.620 1.210 0.790 1.350 ;
        RECT 0.620 1.040 0.810 1.210 ;
        RECT 0.620 0.940 0.790 1.040 ;
        RECT 0.190 0.560 0.360 0.660 ;
        RECT 0.170 0.390 0.360 0.560 ;
        RECT 0.190 0.330 0.360 0.390 ;
        RECT 0.610 0.600 0.780 0.660 ;
        RECT 0.610 0.330 0.860 0.600 ;
        RECT 1.350 0.580 1.600 0.660 ;
        RECT 1.350 0.410 2.650 0.580 ;
        RECT 3.210 0.570 3.380 1.200 ;
        RECT 0.620 0.310 0.860 0.330 ;
        RECT 1.430 0.320 1.600 0.410 ;
        RECT 3.130 0.400 3.460 0.570 ;
      LAYER mcon ;
        RECT 0.640 1.040 0.810 1.210 ;
        RECT 3.210 0.680 3.380 0.850 ;
        RECT 0.650 0.360 0.820 0.530 ;
        RECT 1.990 0.410 2.160 0.580 ;
      LAYER met1 ;
        RECT 0.610 1.260 0.830 1.600 ;
        RECT 0.610 1.000 0.840 1.260 ;
        RECT 0.080 0.320 0.390 0.670 ;
        RECT 0.610 0.600 0.830 1.000 ;
        RECT 0.610 0.290 0.860 0.600 ;
        RECT 1.910 0.360 2.230 0.620 ;
        RECT 0.610 0.090 0.830 0.290 ;
        RECT 3.180 0.090 3.410 1.600 ;
      LAYER via ;
        RECT 0.110 0.350 0.370 0.610 ;
        RECT 1.940 0.360 2.200 0.620 ;
      LAYER met2 ;
        RECT 0.000 1.030 3.610 1.210 ;
        RECT 0.080 0.510 0.400 0.610 ;
        RECT 0.070 0.350 0.400 0.510 ;
        RECT 1.910 0.540 2.230 0.620 ;
        RECT 1.910 0.360 3.610 0.540 ;
  END
END sky130_hilas_VinjInv2

MACRO sky130_hilas_capacitorSize03
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize03 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.020 BY 5.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.420 2.830 5.790 3.110 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.020 2.790 0.290 3.070 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 0.000 5.270 5.780 5.450 ;
        RECT 0.000 4.840 5.780 5.020 ;
        RECT 0.030 3.840 5.780 4.020 ;
        RECT 0.030 3.530 5.780 3.590 ;
        RECT 0.030 3.410 5.820 3.530 ;
        RECT 0.600 3.090 0.970 3.410 ;
        RECT 5.450 3.130 5.820 3.410 ;
        RECT 0.030 2.260 5.780 2.430 ;
        RECT 0.030 1.840 5.780 2.010 ;
        RECT 0.030 0.860 5.780 1.030 ;
        RECT 0.030 0.420 5.780 0.590 ;
      LAYER via2 ;
        RECT 0.650 3.150 0.930 3.430 ;
        RECT 5.500 3.190 5.780 3.470 ;
      LAYER met3 ;
        RECT 0.380 2.890 1.170 3.640 ;
        RECT 1.450 3.320 4.290 5.870 ;
        RECT 5.230 3.320 6.020 3.680 ;
        RECT 1.450 2.930 6.020 3.320 ;
        RECT 1.450 2.570 5.590 2.930 ;
        RECT 1.450 0.000 4.290 2.570 ;
      LAYER via3 ;
        RECT 0.570 3.040 1.000 3.520 ;
        RECT 5.420 3.080 5.850 3.560 ;
      LAYER met4 ;
        RECT 2.570 4.530 3.020 4.540 ;
        RECT 2.550 4.040 3.070 4.530 ;
        RECT 0.470 3.190 1.130 3.610 ;
        RECT 2.580 3.200 3.020 4.040 ;
        RECT 1.160 3.190 2.170 3.200 ;
        RECT 2.570 3.190 3.030 3.200 ;
        RECT 0.450 2.690 3.030 3.190 ;
        RECT 5.320 2.990 5.980 3.650 ;
        RECT 0.450 2.680 1.520 2.690 ;
        RECT 2.570 2.030 3.030 2.690 ;
        RECT 2.570 1.520 3.050 2.030 ;
        RECT 2.550 1.030 3.070 1.520 ;
  END
END sky130_hilas_capacitorSize03

MACRO sky130_hilas_swc4x1BiasCell
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x1BiasCell ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 10.500 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN ROW1
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 7.610 5.510 7.920 5.530 ;
        RECT 0.010 5.330 10.080 5.510 ;
        RECT 0.010 5.320 7.920 5.330 ;
        RECT 7.610 5.200 7.920 5.320 ;
    END
  END ROW1
  PIN ROW2
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 7.610 4.420 7.920 4.550 ;
        RECT 0.010 4.240 10.080 4.420 ;
        RECT 7.610 4.220 7.920 4.240 ;
    END
  END ROW2
  PIN ROW3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.010 2.130 0.480 2.290 ;
        RECT 0.020 2.120 0.480 2.130 ;
    END
    PORT
      LAYER met2 ;
        RECT 7.610 2.270 7.920 2.290 ;
        RECT 0.780 2.100 10.080 2.270 ;
        RECT 7.520 2.090 10.080 2.100 ;
        RECT 7.610 1.960 7.920 2.090 ;
    END
  END ROW3
  PIN ROW4
    USE ANALOG ;
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 0.010 1.300 7.640 1.310 ;
        RECT 0.010 1.170 7.920 1.300 ;
        RECT 0.010 1.140 10.080 1.170 ;
        RECT 7.520 0.990 10.080 1.140 ;
        RECT 7.610 0.970 7.920 0.990 ;
    END
  END ROW4
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 0.436600 ;
    PORT
      LAYER nwell ;
        RECT 0.010 2.530 1.740 4.370 ;
      LAYER met1 ;
        RECT 0.360 0.000 0.760 6.500 ;
    END
  END VTUN
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 3.253900 ;
    PORT
      LAYER nwell ;
        RECT 3.760 0.000 5.990 6.490 ;
      LAYER met1 ;
        RECT 4.410 4.310 4.790 6.500 ;
        RECT 4.400 2.450 4.790 4.310 ;
        RECT 4.410 0.000 4.790 2.450 ;
    END
  END GATE1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 7.520 0.000 10.080 6.500 ;
      LAYER met1 ;
        RECT 9.560 5.790 9.720 6.490 ;
        RECT 9.450 5.240 9.720 5.790 ;
        RECT 9.450 5.190 9.730 5.240 ;
        RECT 9.560 5.100 9.730 5.190 ;
        RECT 9.560 4.650 9.720 5.100 ;
        RECT 9.560 4.560 9.730 4.650 ;
        RECT 9.450 4.510 9.730 4.560 ;
        RECT 9.450 3.960 9.720 4.510 ;
        RECT 9.560 2.550 9.720 3.960 ;
        RECT 9.450 2.000 9.720 2.550 ;
        RECT 9.450 1.950 9.730 2.000 ;
        RECT 9.560 1.860 9.730 1.950 ;
        RECT 9.560 1.400 9.720 1.860 ;
        RECT 9.560 1.310 9.730 1.400 ;
        RECT 9.450 1.260 9.730 1.310 ;
        RECT 9.450 0.710 9.720 1.260 ;
        RECT 9.560 0.010 9.720 0.710 ;
    END
  END VINJ
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 8.750 5.760 8.910 6.490 ;
        RECT 8.750 5.740 8.950 5.760 ;
        RECT 8.730 5.500 8.960 5.740 ;
        RECT 8.750 5.450 8.960 5.500 ;
        RECT 9.120 5.450 9.310 6.440 ;
        RECT 8.750 4.300 8.910 5.450 ;
        RECT 9.140 5.330 9.310 5.450 ;
        RECT 9.150 4.420 9.310 5.330 ;
        RECT 9.140 4.300 9.310 4.420 ;
        RECT 8.750 4.250 8.960 4.300 ;
        RECT 8.730 4.010 8.960 4.250 ;
        RECT 8.750 3.990 8.950 4.010 ;
        RECT 8.750 3.350 8.910 3.990 ;
        RECT 9.120 3.380 9.310 4.300 ;
        RECT 9.100 3.350 9.340 3.380 ;
        RECT 8.750 3.180 9.340 3.350 ;
        RECT 8.750 2.520 8.910 3.180 ;
        RECT 9.100 3.150 9.340 3.180 ;
        RECT 8.750 2.500 8.950 2.520 ;
        RECT 8.730 2.260 8.960 2.500 ;
        RECT 8.750 2.210 8.960 2.260 ;
        RECT 9.120 2.210 9.310 3.150 ;
        RECT 8.750 1.050 8.910 2.210 ;
        RECT 9.140 2.090 9.310 2.210 ;
        RECT 9.150 1.170 9.310 2.090 ;
        RECT 9.140 1.050 9.310 1.170 ;
        RECT 8.750 1.000 8.960 1.050 ;
        RECT 8.730 0.760 8.960 1.000 ;
        RECT 8.750 0.740 8.950 0.760 ;
        RECT 8.750 0.010 8.910 0.740 ;
        RECT 9.120 0.060 9.310 1.050 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 2.540 1.700 2.870 1.730 ;
        RECT 6.570 1.700 6.890 1.760 ;
        RECT 2.540 1.530 6.890 1.700 ;
        RECT 2.540 1.470 2.870 1.530 ;
        RECT 6.570 1.480 6.890 1.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.600 1.790 6.850 6.500 ;
        RECT 6.590 1.760 6.870 1.790 ;
        RECT 6.580 1.480 6.880 1.760 ;
        RECT 6.590 1.460 6.870 1.480 ;
        RECT 6.600 0.000 6.850 1.460 ;
      LAYER via ;
        RECT 6.600 1.490 6.860 1.750 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.570 1.760 2.840 6.500 ;
        RECT 2.550 1.450 2.860 1.760 ;
        RECT 2.570 0.000 2.840 1.450 ;
      LAYER via ;
        RECT 2.570 1.470 2.840 1.730 ;
    END
  END VGND
  PIN DRAIN3
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 7.610 2.710 7.920 2.840 ;
        RECT 7.490 2.700 7.920 2.710 ;
        RECT 7.490 2.540 10.080 2.700 ;
        RECT 7.610 2.520 10.080 2.540 ;
        RECT 7.610 2.510 7.920 2.520 ;
    END
  END DRAIN3
  PIN DRAIN4
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 7.610 0.740 7.920 0.750 ;
        RECT 7.610 0.560 10.080 0.740 ;
        RECT 7.610 0.420 7.920 0.560 ;
    END
  END DRAIN4
  PIN DRAIN1
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 7.610 5.940 7.920 6.080 ;
        RECT 7.610 5.760 10.080 5.940 ;
        RECT 7.610 5.750 7.920 5.760 ;
    END
  END DRAIN1
  PIN DRAIN2
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 7.610 3.990 7.920 4.000 ;
        RECT 7.610 3.830 10.080 3.990 ;
        RECT 7.520 3.810 10.080 3.830 ;
        RECT 7.520 3.690 7.920 3.810 ;
        RECT 7.610 3.670 7.920 3.690 ;
    END
  END DRAIN2
  OBS
      LAYER nwell ;
        RECT 0.580 4.770 1.170 4.930 ;
        RECT 14.520 4.000 16.250 10.500 ;
        RECT 0.580 1.530 1.170 1.680 ;
      LAYER li1 ;
        RECT 7.620 6.030 7.940 6.040 ;
        RECT 7.620 5.860 8.200 6.030 ;
        RECT 7.620 5.810 7.950 5.860 ;
        RECT 7.620 5.780 7.940 5.810 ;
        RECT 9.480 5.760 9.680 6.110 ;
        RECT 7.620 5.450 7.940 5.490 ;
        RECT 7.620 5.410 7.950 5.450 ;
        RECT 7.620 5.240 8.200 5.410 ;
        RECT 7.620 5.230 7.940 5.240 ;
        RECT 8.750 5.140 8.950 5.740 ;
        RECT 9.480 5.730 9.690 5.760 ;
        RECT 9.470 5.140 9.690 5.730 ;
        RECT 2.620 4.480 2.790 5.010 ;
        RECT 6.640 4.450 6.810 4.980 ;
        RECT 7.620 4.510 7.940 4.520 ;
        RECT 7.620 4.340 8.200 4.510 ;
        RECT 7.620 4.300 7.950 4.340 ;
        RECT 7.620 4.260 7.940 4.300 ;
        RECT 8.750 4.010 8.950 4.610 ;
        RECT 9.470 4.020 9.690 4.610 ;
        RECT 9.480 3.990 9.690 4.020 ;
        RECT 7.620 3.940 7.940 3.970 ;
        RECT 7.620 3.890 7.950 3.940 ;
        RECT 0.430 2.980 0.980 3.410 ;
        RECT 2.630 2.550 2.800 3.720 ;
        RECT 4.460 2.910 5.010 3.340 ;
        RECT 6.650 2.590 6.820 3.780 ;
        RECT 7.620 3.720 8.200 3.890 ;
        RECT 7.620 3.710 7.940 3.720 ;
        RECT 9.480 3.640 9.680 3.990 ;
        RECT 8.870 3.180 9.310 3.350 ;
        RECT 7.620 2.790 7.940 2.800 ;
        RECT 7.620 2.620 8.200 2.790 ;
        RECT 7.620 2.570 7.950 2.620 ;
        RECT 7.620 2.540 7.940 2.570 ;
        RECT 9.480 2.520 9.680 2.870 ;
        RECT 7.620 2.210 7.940 2.250 ;
        RECT 7.620 2.170 7.950 2.210 ;
        RECT 7.620 2.000 8.200 2.170 ;
        RECT 7.620 1.990 7.940 2.000 ;
        RECT 8.750 1.900 8.950 2.500 ;
        RECT 9.480 2.490 9.690 2.520 ;
        RECT 9.470 1.900 9.690 2.490 ;
        RECT 7.620 1.260 7.940 1.270 ;
        RECT 7.620 1.090 8.200 1.260 ;
        RECT 7.620 1.050 7.950 1.090 ;
        RECT 7.620 1.010 7.940 1.050 ;
        RECT 8.750 0.760 8.950 1.360 ;
        RECT 9.470 0.770 9.690 1.360 ;
        RECT 9.480 0.740 9.690 0.770 ;
        RECT 7.620 0.690 7.940 0.720 ;
        RECT 7.620 0.640 7.950 0.690 ;
        RECT 7.620 0.470 8.200 0.640 ;
        RECT 7.620 0.460 7.940 0.470 ;
        RECT 9.480 0.390 9.680 0.740 ;
      LAYER mcon ;
        RECT 7.680 5.820 7.850 5.990 ;
        RECT 8.760 5.530 8.930 5.700 ;
        RECT 7.680 5.270 7.850 5.440 ;
        RECT 9.490 5.560 9.660 5.730 ;
        RECT 2.620 4.840 2.790 5.010 ;
        RECT 6.640 4.810 6.810 4.980 ;
        RECT 7.680 4.310 7.850 4.480 ;
        RECT 8.760 4.050 8.930 4.220 ;
        RECT 9.490 4.020 9.660 4.190 ;
        RECT 2.630 3.550 2.800 3.720 ;
        RECT 0.430 3.060 0.700 3.330 ;
        RECT 6.650 3.610 6.820 3.780 ;
        RECT 7.680 3.760 7.850 3.930 ;
        RECT 2.630 2.910 2.800 3.080 ;
        RECT 4.460 2.990 4.730 3.260 ;
        RECT 9.130 3.180 9.310 3.350 ;
        RECT 6.650 2.950 6.820 3.120 ;
        RECT 7.680 2.580 7.850 2.750 ;
        RECT 8.760 2.290 8.930 2.460 ;
        RECT 7.680 2.030 7.850 2.200 ;
        RECT 9.490 2.320 9.660 2.490 ;
        RECT 7.680 1.060 7.850 1.230 ;
        RECT 8.760 0.800 8.930 0.970 ;
        RECT 9.490 0.770 9.660 0.940 ;
        RECT 7.680 0.510 7.850 0.680 ;
      LAYER met1 ;
        RECT 7.610 5.750 7.930 6.070 ;
        RECT 7.610 5.200 7.930 5.520 ;
        RECT 7.610 4.230 7.930 4.550 ;
        RECT 7.610 3.680 7.930 4.000 ;
        RECT 7.610 2.510 7.930 2.830 ;
        RECT 7.610 1.960 7.930 2.280 ;
        RECT 7.610 0.980 7.930 1.300 ;
        RECT 7.610 0.430 7.930 0.750 ;
      LAYER via ;
        RECT 7.640 5.780 7.900 6.040 ;
        RECT 7.640 5.230 7.900 5.490 ;
        RECT 7.640 4.260 7.900 4.520 ;
        RECT 7.640 3.710 7.900 3.970 ;
        RECT 7.640 2.540 7.900 2.800 ;
        RECT 7.640 1.990 7.900 2.250 ;
        RECT 7.640 1.010 7.900 1.270 ;
        RECT 7.640 0.460 7.900 0.720 ;
  END
END sky130_hilas_swc4x1BiasCell

MACRO sky130_hilas_FGtrans2x1cell
  CLASS CORE ;
  FOREIGN sky130_hilas_FGtrans2x1cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.240 BY 10.100 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN COLSEL1
    USE ANALOG ;
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT 10.560 4.640 10.750 6.100 ;
        RECT 10.560 4.610 10.780 4.640 ;
        RECT 10.540 4.340 10.790 4.610 ;
        RECT 10.550 4.330 10.790 4.340 ;
        RECT 10.550 4.090 10.780 4.330 ;
        RECT 10.590 2.060 10.750 4.090 ;
        RECT 10.550 1.820 10.780 2.060 ;
        RECT 10.550 1.810 10.790 1.820 ;
        RECT 10.540 1.540 10.790 1.810 ;
        RECT 10.560 1.510 10.780 1.540 ;
        RECT 10.560 0.050 10.750 1.510 ;
    END
  END COLSEL1
  PIN VINJ
    USE ANALOG ;
    ANTENNADIFFAREA 0.544000 ;
    PORT
      LAYER nwell ;
        RECT 8.210 0.000 11.520 6.150 ;
      LAYER met1 ;
        RECT 11.000 5.450 11.160 6.100 ;
        RECT 10.890 4.900 11.160 5.450 ;
        RECT 10.890 4.850 11.170 4.900 ;
        RECT 11.000 4.760 11.170 4.850 ;
        RECT 11.000 1.390 11.160 4.760 ;
        RECT 11.000 1.300 11.170 1.390 ;
        RECT 10.890 1.250 11.170 1.300 ;
        RECT 10.890 0.700 11.160 1.250 ;
        RECT 11.000 0.050 11.160 0.700 ;
    END
  END VINJ
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 8.790 5.610 9.110 5.620 ;
        RECT 8.790 5.600 9.350 5.610 ;
        RECT 0.000 5.420 11.520 5.600 ;
        RECT 9.040 5.280 9.350 5.420 ;
    END
  END DRAIN1
  PIN DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 9.040 0.730 9.350 0.870 ;
        RECT 9.040 0.720 11.520 0.730 ;
        RECT 0.000 0.570 11.520 0.720 ;
        RECT 9.040 0.550 11.520 0.570 ;
        RECT 9.040 0.540 9.350 0.550 ;
    END
  END DRAIN2
  PIN PROG
    USE ANALOG ;
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER met1 ;
        RECT 7.790 3.380 8.000 6.100 ;
        RECT 7.790 2.870 8.030 3.380 ;
        RECT 7.790 0.050 8.000 2.870 ;
    END
  END PROG
  PIN RUN
    USE ANALOG ;
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER met1 ;
        RECT 6.740 1.570 6.920 6.100 ;
        RECT 6.690 1.230 6.980 1.570 ;
        RECT 6.740 0.050 6.920 1.230 ;
    END
  END RUN
  PIN VIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.217200 ;
    PORT
      LAYER met1 ;
        RECT 8.670 2.670 8.860 2.800 ;
        RECT 8.650 2.380 8.880 2.670 ;
        RECT 8.670 0.760 8.860 2.380 ;
        RECT 8.630 0.550 8.860 0.760 ;
        RECT 8.630 0.470 8.870 0.550 ;
        RECT 8.640 0.050 8.870 0.470 ;
    END
  END VIN2
  PIN VIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.217200 ;
    PORT
      LAYER met1 ;
        RECT 8.670 5.730 8.880 6.100 ;
        RECT 8.660 5.440 8.890 5.730 ;
        RECT 8.670 3.740 8.880 5.440 ;
        RECT 8.660 3.450 8.890 3.740 ;
        RECT 8.670 3.310 8.880 3.450 ;
    END
  END VIN1
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 0.434600 ;
    PORT
      LAYER met1 ;
        RECT 8.220 5.170 8.410 6.100 ;
        RECT 8.190 4.880 8.420 5.170 ;
        RECT 8.220 2.850 8.410 4.880 ;
        RECT 8.190 2.560 8.420 2.850 ;
        RECT 8.220 1.270 8.410 2.560 ;
        RECT 8.200 0.980 8.430 1.270 ;
        RECT 8.220 0.050 8.410 0.980 ;
    END
  END GATE1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2.820 0.050 3.050 6.100 ;
    END
  END VGND
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 1.808400 ;
    PORT
      LAYER nwell ;
        RECT 0.010 1.780 1.740 5.350 ;
        RECT 0.580 1.450 1.140 1.780 ;
      LAYER met1 ;
        RECT 0.340 0.050 0.760 6.100 ;
    END
  END VTUN
  PIN COL1
    ANTENNADIFFAREA 1.030400 ;
    PORT
      LAYER met2 ;
        RECT 10.140 3.180 10.460 3.210 ;
        RECT 0.000 2.950 10.460 3.180 ;
    END
  END COL1
  PIN ROW1
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 9.430 4.060 9.740 4.080 ;
        RECT 0.000 3.870 9.740 4.060 ;
        RECT 9.430 3.750 9.740 3.870 ;
    END
  END ROW1
  PIN ROW2
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 9.440 2.200 9.750 2.390 ;
        RECT 0.000 2.060 9.750 2.200 ;
        RECT 0.000 2.010 9.720 2.060 ;
    END
  END ROW2
  OBS
      LAYER nwell ;
        RECT 14.510 8.200 16.240 10.100 ;
        RECT 3.760 3.710 6.480 5.360 ;
        RECT 14.510 4.060 16.240 5.960 ;
        RECT 3.770 3.670 6.480 3.710 ;
        RECT 3.770 2.340 6.480 2.380 ;
        RECT 3.760 0.690 6.480 2.340 ;
        RECT 0.340 0.060 0.760 0.130 ;
      LAYER li1 ;
        RECT 8.680 5.670 8.870 5.700 ;
        RECT 7.810 5.500 8.870 5.670 ;
        RECT 9.110 5.520 9.640 5.690 ;
        RECT 7.810 5.110 7.980 5.500 ;
        RECT 8.680 5.470 8.870 5.500 ;
        RECT 10.920 5.420 11.120 5.770 ;
        RECT 10.920 5.390 11.130 5.420 ;
        RECT 7.240 4.940 7.980 5.110 ;
        RECT 8.210 5.110 8.400 5.140 ;
        RECT 8.210 4.940 8.940 5.110 ;
        RECT 8.210 4.910 8.400 4.940 ;
        RECT 0.430 3.960 0.980 4.390 ;
        RECT 5.950 4.320 6.180 4.840 ;
        RECT 5.950 4.150 8.940 4.320 ;
        RECT 9.360 4.040 9.530 5.130 ;
        RECT 9.360 4.000 9.760 4.040 ;
        RECT 9.360 3.810 9.770 4.000 ;
        RECT 9.360 3.780 9.760 3.810 ;
        RECT 8.680 3.530 8.870 3.710 ;
        RECT 3.030 3.130 3.220 3.530 ;
        RECT 7.250 3.360 7.590 3.530 ;
        RECT 2.840 3.120 3.220 3.130 ;
        RECT 2.840 2.940 6.580 3.120 ;
        RECT 2.840 2.900 3.220 2.940 ;
        RECT 0.430 2.230 0.980 2.660 ;
        RECT 3.030 2.520 3.220 2.900 ;
        RECT 7.330 2.790 7.500 3.360 ;
        RECT 7.810 2.950 8.020 3.380 ;
        RECT 8.590 3.360 8.940 3.530 ;
        RECT 9.360 3.440 9.530 3.780 ;
        RECT 10.190 3.530 10.360 5.140 ;
        RECT 10.910 4.810 11.130 5.390 ;
        RECT 10.920 4.800 11.130 4.810 ;
        RECT 10.560 4.630 10.750 4.640 ;
        RECT 10.560 4.340 10.760 4.630 ;
        RECT 10.550 4.010 10.820 4.340 ;
        RECT 10.190 3.340 10.370 3.530 ;
        RECT 7.830 2.930 8.000 2.950 ;
        RECT 7.250 2.760 7.590 2.790 ;
        RECT 8.210 2.770 8.400 2.820 ;
        RECT 8.170 2.760 8.400 2.770 ;
        RECT 7.250 2.620 8.400 2.760 ;
        RECT 8.590 2.620 8.940 2.790 ;
        RECT 7.420 2.590 8.400 2.620 ;
        RECT 7.420 2.560 8.260 2.590 ;
        RECT 8.670 2.410 8.860 2.620 ;
        RECT 9.360 2.350 9.530 2.710 ;
        RECT 10.190 2.620 10.370 2.810 ;
        RECT 9.360 2.310 9.770 2.350 ;
        RECT 9.360 2.120 9.780 2.310 ;
        RECT 9.360 2.090 9.770 2.120 ;
        RECT 6.010 1.900 8.940 2.000 ;
        RECT 5.950 1.830 8.940 1.900 ;
        RECT 5.950 1.210 6.180 1.830 ;
        RECT 6.750 1.510 6.920 1.570 ;
        RECT 6.730 1.300 6.940 1.510 ;
        RECT 6.750 1.230 6.920 1.300 ;
        RECT 8.220 1.210 8.410 1.240 ;
        RECT 7.240 1.040 8.050 1.210 ;
        RECT 7.860 0.700 8.050 1.040 ;
        RECT 8.220 1.040 8.940 1.210 ;
        RECT 8.220 1.010 8.410 1.040 ;
        RECT 9.360 1.020 9.530 2.090 ;
        RECT 10.190 1.010 10.360 2.620 ;
        RECT 10.550 1.810 10.820 2.140 ;
        RECT 10.560 1.520 10.760 1.810 ;
        RECT 10.560 1.510 10.750 1.520 ;
        RECT 10.920 1.340 11.130 1.350 ;
        RECT 10.910 0.760 11.130 1.340 ;
        RECT 10.920 0.730 11.130 0.760 ;
        RECT 8.650 0.700 8.840 0.730 ;
        RECT 7.860 0.520 8.840 0.700 ;
        RECT 8.650 0.500 8.840 0.520 ;
        RECT 9.110 0.460 9.640 0.630 ;
        RECT 10.920 0.380 11.120 0.730 ;
      LAYER mcon ;
        RECT 8.690 5.500 8.860 5.670 ;
        RECT 10.930 5.220 11.100 5.390 ;
        RECT 8.220 4.940 8.390 5.110 ;
        RECT 5.980 4.640 6.150 4.810 ;
        RECT 0.430 4.040 0.700 4.310 ;
        RECT 5.980 4.190 6.150 4.360 ;
        RECT 9.500 3.820 9.670 3.990 ;
        RECT 8.690 3.510 8.860 3.680 ;
        RECT 2.850 2.930 3.020 3.100 ;
        RECT 0.430 2.310 0.700 2.580 ;
        RECT 10.570 4.380 10.750 4.570 ;
        RECT 8.220 2.620 8.390 2.790 ;
        RECT 8.680 2.440 8.850 2.610 ;
        RECT 9.510 2.130 9.680 2.300 ;
        RECT 5.980 1.690 6.150 1.860 ;
        RECT 5.980 1.240 6.150 1.410 ;
        RECT 8.230 1.040 8.400 1.210 ;
        RECT 10.570 1.580 10.750 1.770 ;
        RECT 10.930 0.760 11.100 0.930 ;
        RECT 8.660 0.530 8.830 0.700 ;
      LAYER met1 ;
        RECT 9.040 5.280 9.350 5.720 ;
        RECT 5.940 4.100 6.200 4.890 ;
        RECT 9.430 3.750 9.750 4.070 ;
        RECT 10.160 3.240 10.400 3.660 ;
        RECT 10.160 2.920 10.430 3.240 ;
        RECT 10.160 2.490 10.400 2.920 ;
        RECT 9.440 2.060 9.760 2.380 ;
        RECT 5.940 1.160 6.200 1.950 ;
        RECT 9.040 0.430 9.350 0.870 ;
      LAYER via ;
        RECT 9.070 5.310 9.330 5.570 ;
        RECT 9.460 3.780 9.720 4.040 ;
        RECT 10.170 2.950 10.430 3.210 ;
        RECT 9.470 2.090 9.730 2.350 ;
        RECT 9.070 0.580 9.330 0.840 ;
  END
END sky130_hilas_FGtrans2x1cell

MACRO sky130_hilas_capacitorSize01
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.090 BY 7.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 10.060 2.380 10.420 2.660 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.020 2.370 0.290 2.650 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 0.000 4.850 10.420 5.030 ;
        RECT 0.000 4.420 10.420 4.600 ;
        RECT 0.030 3.420 10.420 3.600 ;
        RECT 8.510 3.170 10.420 3.180 ;
        RECT 0.030 3.080 10.420 3.170 ;
        RECT 0.030 2.990 10.460 3.080 ;
        RECT 0.600 2.670 0.970 2.990 ;
        RECT 10.090 2.680 10.460 2.990 ;
        RECT 0.030 1.840 10.420 2.010 ;
        RECT 0.030 1.420 10.420 1.590 ;
        RECT 0.030 0.440 10.420 0.610 ;
        RECT 0.030 0.000 10.420 0.170 ;
      LAYER via2 ;
        RECT 0.650 2.730 0.930 3.010 ;
        RECT 10.140 2.740 10.420 3.020 ;
      LAYER met3 ;
        RECT 5.890 7.840 8.710 7.870 ;
        RECT 0.380 2.470 1.170 3.220 ;
        RECT 5.890 2.060 13.090 7.840 ;
        RECT 8.680 2.040 13.090 2.060 ;
      LAYER via3 ;
        RECT 0.570 2.620 1.000 3.100 ;
        RECT 10.060 2.630 10.490 3.110 ;
      LAYER met4 ;
        RECT 0.470 2.770 1.130 3.190 ;
        RECT 6.780 3.140 9.820 3.610 ;
        RECT 1.160 2.770 2.170 2.780 ;
        RECT 0.450 2.270 3.800 2.770 ;
        RECT 9.960 2.540 10.620 3.200 ;
        RECT 0.450 2.260 1.520 2.270 ;
        RECT 3.160 1.150 3.790 2.270 ;
        RECT 3.160 0.850 5.310 1.150 ;
        RECT 3.490 0.840 5.310 0.850 ;
  END
END sky130_hilas_capacitorSize01

MACRO sky130_hilas_Tgate4Double01
  CLASS CORE ;
  FOREIGN sky130_hilas_Tgate4Double01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.080 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER nwell ;
        RECT 0.120 0.000 3.590 6.050 ;
      LAYER met1 ;
        RECT 0.740 5.100 0.940 6.050 ;
        RECT 0.740 4.810 1.060 5.100 ;
        RECT 0.740 4.260 0.940 4.810 ;
        RECT 0.740 3.970 1.060 4.260 ;
        RECT 0.740 2.080 0.940 3.970 ;
        RECT 0.740 1.790 1.060 2.080 ;
        RECT 0.740 1.240 0.940 1.790 ;
        RECT 0.740 0.950 1.060 1.240 ;
        RECT 0.740 0.000 0.940 0.950 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.570 5.100 6.760 6.050 ;
        RECT 6.570 4.810 6.880 5.100 ;
        RECT 6.570 4.260 6.760 4.810 ;
        RECT 6.570 3.970 6.880 4.260 ;
        RECT 6.570 2.080 6.760 3.970 ;
        RECT 6.570 1.790 6.880 2.080 ;
        RECT 6.570 1.240 6.760 1.790 ;
        RECT 6.570 0.950 6.880 1.240 ;
        RECT 6.570 0.000 6.760 0.950 ;
    END
  END VGND
  PIN INPUT1_1
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.450 5.940 2.760 5.950 ;
        RECT 0.000 5.740 5.840 5.940 ;
        RECT 2.450 5.620 2.760 5.740 ;
        RECT 5.530 5.610 5.840 5.740 ;
    END
  END INPUT1_1
  PIN SELECT1
    ANTENNAGATEAREA 0.992000 ;
    PORT
      LAYER met2 ;
        RECT 0.000 4.760 0.610 4.960 ;
        RECT 0.290 4.670 0.610 4.760 ;
        RECT 0.290 4.310 0.610 4.400 ;
        RECT 0.000 4.110 0.610 4.310 ;
    END
  END SELECT1
  PIN INPUT2_2
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 1.100 3.810 1.410 3.820 ;
        RECT 4.020 3.810 4.330 3.820 ;
        RECT 0.000 3.610 4.370 3.810 ;
        RECT 1.100 3.490 1.410 3.610 ;
        RECT 4.020 3.490 4.330 3.610 ;
    END
  END INPUT2_2
  PIN INPUT1_2
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.450 3.330 2.760 3.450 ;
        RECT 5.530 3.330 5.840 3.460 ;
        RECT 0.000 3.130 5.840 3.330 ;
        RECT 2.450 3.120 2.760 3.130 ;
    END
  END INPUT1_2
  PIN SELECT3
    ANTENNAGATEAREA 0.992000 ;
    PORT
      LAYER met2 ;
        RECT 0.000 1.740 0.610 1.940 ;
        RECT 0.290 1.650 0.610 1.740 ;
        RECT 0.290 1.290 0.610 1.380 ;
        RECT 0.000 1.090 0.610 1.290 ;
    END
  END SELECT3
  PIN INPUT2_3
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 1.100 2.440 1.410 2.560 ;
        RECT 4.020 2.440 4.330 2.560 ;
        RECT 0.000 2.240 4.370 2.440 ;
        RECT 1.100 2.230 1.410 2.240 ;
        RECT 4.020 2.230 4.330 2.240 ;
    END
  END INPUT2_3
  PIN INPUT2_4
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 1.100 0.790 1.410 0.800 ;
        RECT 4.020 0.790 4.330 0.800 ;
        RECT 0.000 0.590 4.370 0.790 ;
        RECT 1.100 0.470 1.410 0.590 ;
        RECT 4.020 0.470 4.330 0.590 ;
    END
  END INPUT2_4
  PIN INPUT1_4
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.450 0.310 2.760 0.430 ;
        RECT 5.530 0.310 5.840 0.440 ;
        RECT 0.000 0.110 5.840 0.310 ;
        RECT 2.450 0.100 2.760 0.110 ;
    END
  END INPUT1_4
  PIN OUTPUT4
    ANTENNADIFFAREA 0.275900 ;
    PORT
      LAYER met2 ;
        RECT 1.680 1.290 2.000 1.300 ;
        RECT 3.100 1.290 3.420 1.310 ;
        RECT 4.850 1.290 5.170 1.330 ;
        RECT 5.890 1.290 6.210 1.320 ;
        RECT 1.680 1.090 7.080 1.290 ;
        RECT 1.680 1.040 2.000 1.090 ;
        RECT 3.100 1.050 3.420 1.090 ;
        RECT 4.850 1.070 5.170 1.090 ;
        RECT 5.890 1.060 6.210 1.090 ;
    END
  END OUTPUT4
  PIN OUTPUT3
    ANTENNADIFFAREA 0.275900 ;
    PORT
      LAYER met2 ;
        RECT 1.680 1.940 2.000 1.990 ;
        RECT 3.100 1.940 3.420 1.980 ;
        RECT 4.850 1.940 5.170 1.960 ;
        RECT 5.890 1.940 6.210 1.970 ;
        RECT 1.680 1.740 7.080 1.940 ;
        RECT 1.680 1.730 2.000 1.740 ;
        RECT 3.100 1.720 3.420 1.740 ;
        RECT 4.850 1.700 5.170 1.740 ;
        RECT 5.890 1.710 6.210 1.740 ;
    END
  END OUTPUT3
  PIN OUTPUT2
    ANTENNADIFFAREA 0.275900 ;
    PORT
      LAYER met2 ;
        RECT 1.680 4.310 2.000 4.320 ;
        RECT 3.100 4.310 3.420 4.330 ;
        RECT 4.850 4.310 5.170 4.350 ;
        RECT 5.890 4.310 6.210 4.340 ;
        RECT 1.680 4.110 7.080 4.310 ;
        RECT 1.680 4.060 2.000 4.110 ;
        RECT 3.100 4.070 3.420 4.110 ;
        RECT 4.850 4.090 5.170 4.110 ;
        RECT 5.890 4.080 6.210 4.110 ;
    END
  END OUTPUT2
  PIN OUTPUT1
    ANTENNADIFFAREA 0.275900 ;
    PORT
      LAYER met2 ;
        RECT 1.680 4.960 2.000 5.010 ;
        RECT 3.100 4.960 3.420 5.000 ;
        RECT 4.850 4.960 5.170 4.980 ;
        RECT 5.890 4.960 6.210 4.990 ;
        RECT 1.680 4.760 7.080 4.960 ;
        RECT 1.680 4.750 2.000 4.760 ;
        RECT 3.100 4.740 3.420 4.760 ;
        RECT 4.850 4.720 5.170 4.760 ;
        RECT 5.890 4.730 6.210 4.760 ;
    END
  END OUTPUT1
  PIN INPUT2_1
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 1.100 5.460 1.410 5.580 ;
        RECT 4.020 5.460 4.330 5.580 ;
        RECT 0.000 5.260 4.370 5.460 ;
        RECT 1.100 5.250 1.410 5.260 ;
        RECT 4.020 5.250 4.330 5.260 ;
    END
  END INPUT2_1
  PIN INPUT1_3
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.450 2.920 2.760 2.930 ;
        RECT 0.000 2.720 5.840 2.920 ;
        RECT 2.450 2.600 2.760 2.720 ;
        RECT 5.530 2.590 5.840 2.720 ;
    END
  END INPUT1_3
  OBS
      LAYER li1 ;
        RECT 2.460 5.890 2.780 5.920 ;
        RECT 0.430 5.540 0.600 5.820 ;
        RECT 0.940 5.580 1.290 5.750 ;
        RECT 1.110 5.550 1.290 5.580 ;
        RECT 0.430 5.500 0.640 5.540 ;
        RECT 1.110 5.520 1.430 5.550 ;
        RECT 0.430 5.480 0.660 5.500 ;
        RECT 0.430 5.460 0.690 5.480 ;
        RECT 0.430 5.410 0.770 5.460 ;
        RECT 0.430 5.350 0.920 5.410 ;
        RECT 0.430 5.320 0.940 5.350 ;
        RECT 0.470 5.290 0.940 5.320 ;
        RECT 1.110 5.330 1.440 5.520 ;
        RECT 1.710 5.480 1.880 5.830 ;
        RECT 2.460 5.700 2.790 5.890 ;
        RECT 5.540 5.880 5.860 5.910 ;
        RECT 2.460 5.660 2.780 5.700 ;
        RECT 2.490 5.490 2.660 5.660 ;
        RECT 3.180 5.480 3.350 5.830 ;
        RECT 4.140 5.550 4.310 5.830 ;
        RECT 4.030 5.520 4.350 5.550 ;
        RECT 1.710 5.340 2.010 5.480 ;
        RECT 1.110 5.290 1.430 5.330 ;
        RECT 0.600 5.240 0.940 5.290 ;
        RECT 1.820 5.250 2.010 5.340 ;
        RECT 0.720 5.230 0.940 5.240 ;
        RECT 0.730 5.200 0.940 5.230 ;
        RECT 0.750 5.120 0.940 5.200 ;
        RECT 2.110 5.120 2.440 5.240 ;
        RECT 3.270 5.230 3.460 5.460 ;
        RECT 4.030 5.330 4.360 5.520 ;
        RECT 4.880 5.470 5.050 5.840 ;
        RECT 5.540 5.690 5.870 5.880 ;
        RECT 6.260 5.690 6.550 5.740 ;
        RECT 5.540 5.650 5.860 5.690 ;
        RECT 5.600 5.490 5.770 5.650 ;
        RECT 6.210 5.570 6.550 5.690 ;
        RECT 4.880 5.460 5.170 5.470 ;
        RECT 6.210 5.460 6.400 5.570 ;
        RECT 4.030 5.290 4.350 5.330 ;
        RECT 4.980 5.240 5.170 5.460 ;
        RECT 6.830 5.150 7.000 5.830 ;
        RECT 0.750 5.070 1.270 5.120 ;
        RECT 0.850 4.950 1.270 5.070 ;
        RECT 0.850 4.840 1.040 4.950 ;
        RECT 1.620 4.940 5.840 5.120 ;
        RECT 6.220 4.940 6.570 5.110 ;
        RECT 6.750 5.070 7.000 5.150 ;
        RECT 6.670 4.950 7.000 5.070 ;
        RECT 6.670 4.840 6.860 4.950 ;
        RECT 0.350 4.810 0.520 4.830 ;
        RECT 0.330 4.260 0.540 4.810 ;
        RECT 0.350 4.240 0.520 4.260 ;
        RECT 0.850 4.120 1.040 4.230 ;
        RECT 0.850 4.000 1.270 4.120 ;
        RECT 0.750 3.950 1.270 4.000 ;
        RECT 1.620 3.950 5.840 4.130 ;
        RECT 6.220 3.960 6.570 4.130 ;
        RECT 6.670 4.120 6.860 4.230 ;
        RECT 6.670 4.000 7.000 4.120 ;
        RECT 0.750 3.870 0.940 3.950 ;
        RECT 0.730 3.840 0.940 3.870 ;
        RECT 0.720 3.830 0.940 3.840 ;
        RECT 2.110 3.830 2.440 3.950 ;
        RECT 6.750 3.920 7.000 4.000 ;
        RECT 0.600 3.780 0.940 3.830 ;
        RECT 0.470 3.750 0.940 3.780 ;
        RECT 0.430 3.720 0.940 3.750 ;
        RECT 1.110 3.740 1.430 3.780 ;
        RECT 0.430 3.660 0.920 3.720 ;
        RECT 0.430 3.610 0.770 3.660 ;
        RECT 0.430 3.590 0.690 3.610 ;
        RECT 0.430 3.570 0.660 3.590 ;
        RECT 0.430 3.530 0.640 3.570 ;
        RECT 1.110 3.550 1.440 3.740 ;
        RECT 1.820 3.730 2.010 3.820 ;
        RECT 1.710 3.590 2.010 3.730 ;
        RECT 3.270 3.610 3.460 3.840 ;
        RECT 4.030 3.740 4.350 3.780 ;
        RECT 0.430 3.250 0.600 3.530 ;
        RECT 1.110 3.520 1.430 3.550 ;
        RECT 1.110 3.490 1.290 3.520 ;
        RECT 0.940 3.320 1.290 3.490 ;
        RECT 1.710 3.240 1.880 3.590 ;
        RECT 2.490 3.410 2.660 3.580 ;
        RECT 2.460 3.370 2.780 3.410 ;
        RECT 2.460 3.180 2.790 3.370 ;
        RECT 3.180 3.240 3.350 3.590 ;
        RECT 4.030 3.550 4.360 3.740 ;
        RECT 4.980 3.610 5.170 3.830 ;
        RECT 4.880 3.600 5.170 3.610 ;
        RECT 4.030 3.520 4.350 3.550 ;
        RECT 4.140 3.240 4.310 3.520 ;
        RECT 4.880 3.230 5.050 3.600 ;
        RECT 5.600 3.420 5.770 3.580 ;
        RECT 6.210 3.500 6.400 3.610 ;
        RECT 5.540 3.380 5.860 3.420 ;
        RECT 6.210 3.380 6.550 3.500 ;
        RECT 5.540 3.190 5.870 3.380 ;
        RECT 6.260 3.330 6.550 3.380 ;
        RECT 6.830 3.240 7.000 3.920 ;
        RECT 2.460 3.150 2.780 3.180 ;
        RECT 5.540 3.160 5.860 3.190 ;
        RECT 2.460 2.870 2.780 2.900 ;
        RECT 0.430 2.520 0.600 2.800 ;
        RECT 0.940 2.560 1.290 2.730 ;
        RECT 1.110 2.530 1.290 2.560 ;
        RECT 0.430 2.480 0.640 2.520 ;
        RECT 1.110 2.500 1.430 2.530 ;
        RECT 0.430 2.460 0.660 2.480 ;
        RECT 0.430 2.440 0.690 2.460 ;
        RECT 0.430 2.390 0.770 2.440 ;
        RECT 0.430 2.330 0.920 2.390 ;
        RECT 0.430 2.300 0.940 2.330 ;
        RECT 0.470 2.270 0.940 2.300 ;
        RECT 1.110 2.310 1.440 2.500 ;
        RECT 1.710 2.460 1.880 2.810 ;
        RECT 2.460 2.680 2.790 2.870 ;
        RECT 5.540 2.860 5.860 2.890 ;
        RECT 2.460 2.640 2.780 2.680 ;
        RECT 2.490 2.470 2.660 2.640 ;
        RECT 3.180 2.460 3.350 2.810 ;
        RECT 4.140 2.530 4.310 2.810 ;
        RECT 4.030 2.500 4.350 2.530 ;
        RECT 1.710 2.320 2.010 2.460 ;
        RECT 1.110 2.270 1.430 2.310 ;
        RECT 0.600 2.220 0.940 2.270 ;
        RECT 1.820 2.230 2.010 2.320 ;
        RECT 0.720 2.210 0.940 2.220 ;
        RECT 0.730 2.180 0.940 2.210 ;
        RECT 0.750 2.100 0.940 2.180 ;
        RECT 2.110 2.100 2.440 2.220 ;
        RECT 3.270 2.210 3.460 2.440 ;
        RECT 4.030 2.310 4.360 2.500 ;
        RECT 4.880 2.450 5.050 2.820 ;
        RECT 5.540 2.670 5.870 2.860 ;
        RECT 6.260 2.670 6.550 2.720 ;
        RECT 5.540 2.630 5.860 2.670 ;
        RECT 5.600 2.470 5.770 2.630 ;
        RECT 6.210 2.550 6.550 2.670 ;
        RECT 4.880 2.440 5.170 2.450 ;
        RECT 6.210 2.440 6.400 2.550 ;
        RECT 4.030 2.270 4.350 2.310 ;
        RECT 4.980 2.220 5.170 2.440 ;
        RECT 6.830 2.130 7.000 2.810 ;
        RECT 0.750 2.050 1.270 2.100 ;
        RECT 0.850 1.930 1.270 2.050 ;
        RECT 0.850 1.820 1.040 1.930 ;
        RECT 1.620 1.920 5.840 2.100 ;
        RECT 6.220 1.920 6.570 2.090 ;
        RECT 6.750 2.050 7.000 2.130 ;
        RECT 6.670 1.930 7.000 2.050 ;
        RECT 6.670 1.820 6.860 1.930 ;
        RECT 0.350 1.790 0.520 1.810 ;
        RECT 0.330 1.240 0.540 1.790 ;
        RECT 0.350 1.220 0.520 1.240 ;
        RECT 0.850 1.100 1.040 1.210 ;
        RECT 0.850 0.980 1.270 1.100 ;
        RECT 0.750 0.930 1.270 0.980 ;
        RECT 1.620 0.930 5.840 1.110 ;
        RECT 6.220 0.940 6.570 1.110 ;
        RECT 6.670 1.100 6.860 1.210 ;
        RECT 6.670 0.980 7.000 1.100 ;
        RECT 0.750 0.850 0.940 0.930 ;
        RECT 0.730 0.820 0.940 0.850 ;
        RECT 0.720 0.810 0.940 0.820 ;
        RECT 2.110 0.810 2.440 0.930 ;
        RECT 6.750 0.900 7.000 0.980 ;
        RECT 0.600 0.760 0.940 0.810 ;
        RECT 0.470 0.730 0.940 0.760 ;
        RECT 0.430 0.700 0.940 0.730 ;
        RECT 1.110 0.720 1.430 0.760 ;
        RECT 0.430 0.640 0.920 0.700 ;
        RECT 0.430 0.590 0.770 0.640 ;
        RECT 0.430 0.570 0.690 0.590 ;
        RECT 0.430 0.550 0.660 0.570 ;
        RECT 0.430 0.510 0.640 0.550 ;
        RECT 1.110 0.530 1.440 0.720 ;
        RECT 1.820 0.710 2.010 0.800 ;
        RECT 1.710 0.570 2.010 0.710 ;
        RECT 3.270 0.590 3.460 0.820 ;
        RECT 4.030 0.720 4.350 0.760 ;
        RECT 0.430 0.230 0.600 0.510 ;
        RECT 1.110 0.500 1.430 0.530 ;
        RECT 1.110 0.470 1.290 0.500 ;
        RECT 0.940 0.300 1.290 0.470 ;
        RECT 1.710 0.220 1.880 0.570 ;
        RECT 2.490 0.390 2.660 0.560 ;
        RECT 2.460 0.350 2.780 0.390 ;
        RECT 2.460 0.160 2.790 0.350 ;
        RECT 3.180 0.220 3.350 0.570 ;
        RECT 4.030 0.530 4.360 0.720 ;
        RECT 4.980 0.590 5.170 0.810 ;
        RECT 4.880 0.580 5.170 0.590 ;
        RECT 4.030 0.500 4.350 0.530 ;
        RECT 4.140 0.220 4.310 0.500 ;
        RECT 4.880 0.210 5.050 0.580 ;
        RECT 5.600 0.400 5.770 0.560 ;
        RECT 6.210 0.480 6.400 0.590 ;
        RECT 5.540 0.360 5.860 0.400 ;
        RECT 6.210 0.360 6.550 0.480 ;
        RECT 5.540 0.170 5.870 0.360 ;
        RECT 6.260 0.310 6.550 0.360 ;
        RECT 6.830 0.220 7.000 0.900 ;
        RECT 2.460 0.130 2.780 0.160 ;
        RECT 5.540 0.140 5.860 0.170 ;
      LAYER mcon ;
        RECT 1.170 5.340 1.340 5.510 ;
        RECT 2.520 5.710 2.690 5.880 ;
        RECT 1.830 5.280 2.000 5.450 ;
        RECT 3.280 5.260 3.450 5.430 ;
        RECT 4.090 5.340 4.260 5.510 ;
        RECT 5.600 5.700 5.770 5.870 ;
        RECT 6.220 5.490 6.390 5.660 ;
        RECT 4.990 5.270 5.160 5.440 ;
        RECT 0.860 4.870 1.030 5.040 ;
        RECT 6.680 4.870 6.850 5.040 ;
        RECT 0.350 4.660 0.520 4.830 ;
        RECT 0.860 4.030 1.030 4.200 ;
        RECT 6.680 4.030 6.850 4.200 ;
        RECT 1.170 3.560 1.340 3.730 ;
        RECT 1.830 3.620 2.000 3.790 ;
        RECT 3.280 3.640 3.450 3.810 ;
        RECT 2.520 3.190 2.690 3.360 ;
        RECT 4.090 3.560 4.260 3.730 ;
        RECT 4.990 3.630 5.160 3.800 ;
        RECT 6.220 3.410 6.390 3.580 ;
        RECT 5.600 3.200 5.770 3.370 ;
        RECT 1.170 2.320 1.340 2.490 ;
        RECT 2.520 2.690 2.690 2.860 ;
        RECT 1.830 2.260 2.000 2.430 ;
        RECT 3.280 2.240 3.450 2.410 ;
        RECT 4.090 2.320 4.260 2.490 ;
        RECT 5.600 2.680 5.770 2.850 ;
        RECT 6.220 2.470 6.390 2.640 ;
        RECT 4.990 2.250 5.160 2.420 ;
        RECT 0.860 1.850 1.030 2.020 ;
        RECT 6.680 1.850 6.850 2.020 ;
        RECT 0.350 1.640 0.520 1.810 ;
        RECT 0.860 1.010 1.030 1.180 ;
        RECT 6.680 1.010 6.850 1.180 ;
        RECT 1.170 0.540 1.340 0.710 ;
        RECT 1.830 0.600 2.000 0.770 ;
        RECT 3.280 0.620 3.450 0.790 ;
        RECT 2.520 0.170 2.690 0.340 ;
        RECT 4.090 0.540 4.260 0.710 ;
        RECT 4.990 0.610 5.160 0.780 ;
        RECT 6.220 0.390 6.390 0.560 ;
        RECT 5.600 0.180 5.770 0.350 ;
      LAYER met1 ;
        RECT 2.450 5.630 2.770 5.950 ;
        RECT 5.530 5.620 5.850 5.940 ;
        RECT 1.100 5.260 1.420 5.580 ;
        RECT 1.800 5.310 2.030 5.510 ;
        RECT 1.720 5.220 2.030 5.310 ;
        RECT 3.250 5.290 3.480 5.490 ;
        RECT 1.720 5.040 1.890 5.220 ;
        RECT 3.170 5.200 3.480 5.290 ;
        RECT 4.020 5.260 4.340 5.580 ;
        RECT 6.190 5.520 6.420 5.720 ;
        RECT 4.960 5.320 5.190 5.500 ;
        RECT 4.890 5.210 5.190 5.320 ;
        RECT 6.090 5.430 6.420 5.520 ;
        RECT 0.320 4.640 0.580 4.960 ;
        RECT 1.710 4.720 1.970 5.040 ;
        RECT 3.170 5.030 3.340 5.200 ;
        RECT 3.130 4.710 3.390 5.030 ;
        RECT 4.890 5.010 5.060 5.210 ;
        RECT 6.090 5.020 6.280 5.430 ;
        RECT 4.880 4.690 5.140 5.010 ;
        RECT 5.920 4.770 6.280 5.020 ;
        RECT 5.920 4.700 6.180 4.770 ;
        RECT 0.320 4.600 0.550 4.640 ;
        RECT 0.330 4.470 0.550 4.600 ;
        RECT 0.320 4.430 0.550 4.470 ;
        RECT 0.320 4.110 0.580 4.430 ;
        RECT 1.710 4.030 1.970 4.350 ;
        RECT 3.130 4.040 3.390 4.360 ;
        RECT 4.880 4.060 5.140 4.380 ;
        RECT 5.920 4.300 6.180 4.370 ;
        RECT 1.720 3.850 1.890 4.030 ;
        RECT 3.170 3.870 3.340 4.040 ;
        RECT 1.100 3.490 1.420 3.810 ;
        RECT 1.720 3.760 2.030 3.850 ;
        RECT 3.170 3.780 3.480 3.870 ;
        RECT 4.890 3.860 5.060 4.060 ;
        RECT 5.920 4.050 6.280 4.300 ;
        RECT 1.800 3.560 2.030 3.760 ;
        RECT 3.250 3.580 3.480 3.780 ;
        RECT 4.020 3.490 4.340 3.810 ;
        RECT 4.890 3.750 5.190 3.860 ;
        RECT 4.960 3.570 5.190 3.750 ;
        RECT 6.090 3.640 6.280 4.050 ;
        RECT 6.090 3.550 6.420 3.640 ;
        RECT 2.450 3.120 2.770 3.440 ;
        RECT 5.530 3.130 5.850 3.450 ;
        RECT 6.190 3.350 6.420 3.550 ;
        RECT 2.450 2.610 2.770 2.930 ;
        RECT 5.530 2.600 5.850 2.920 ;
        RECT 1.100 2.240 1.420 2.560 ;
        RECT 1.800 2.290 2.030 2.490 ;
        RECT 1.720 2.200 2.030 2.290 ;
        RECT 3.250 2.270 3.480 2.470 ;
        RECT 1.720 2.020 1.890 2.200 ;
        RECT 3.170 2.180 3.480 2.270 ;
        RECT 4.020 2.240 4.340 2.560 ;
        RECT 6.190 2.500 6.420 2.700 ;
        RECT 4.960 2.300 5.190 2.480 ;
        RECT 4.890 2.190 5.190 2.300 ;
        RECT 6.090 2.410 6.420 2.500 ;
        RECT 0.320 1.620 0.580 1.940 ;
        RECT 1.710 1.700 1.970 2.020 ;
        RECT 3.170 2.010 3.340 2.180 ;
        RECT 3.130 1.690 3.390 2.010 ;
        RECT 4.890 1.990 5.060 2.190 ;
        RECT 6.090 2.000 6.280 2.410 ;
        RECT 4.880 1.670 5.140 1.990 ;
        RECT 5.920 1.750 6.280 2.000 ;
        RECT 5.920 1.680 6.180 1.750 ;
        RECT 0.320 1.580 0.550 1.620 ;
        RECT 0.330 1.450 0.550 1.580 ;
        RECT 0.320 1.410 0.550 1.450 ;
        RECT 0.320 1.090 0.580 1.410 ;
        RECT 1.710 1.010 1.970 1.330 ;
        RECT 3.130 1.020 3.390 1.340 ;
        RECT 4.880 1.040 5.140 1.360 ;
        RECT 5.920 1.280 6.180 1.350 ;
        RECT 1.720 0.830 1.890 1.010 ;
        RECT 3.170 0.850 3.340 1.020 ;
        RECT 1.100 0.470 1.420 0.790 ;
        RECT 1.720 0.740 2.030 0.830 ;
        RECT 3.170 0.760 3.480 0.850 ;
        RECT 4.890 0.840 5.060 1.040 ;
        RECT 5.920 1.030 6.280 1.280 ;
        RECT 1.800 0.540 2.030 0.740 ;
        RECT 3.250 0.560 3.480 0.760 ;
        RECT 4.020 0.470 4.340 0.790 ;
        RECT 4.890 0.730 5.190 0.840 ;
        RECT 4.960 0.550 5.190 0.730 ;
        RECT 6.090 0.620 6.280 1.030 ;
        RECT 6.090 0.530 6.420 0.620 ;
        RECT 2.450 0.100 2.770 0.420 ;
        RECT 5.530 0.110 5.850 0.430 ;
        RECT 6.190 0.330 6.420 0.530 ;
      LAYER via ;
        RECT 2.480 5.660 2.740 5.920 ;
        RECT 5.560 5.650 5.820 5.910 ;
        RECT 1.130 5.290 1.390 5.550 ;
        RECT 4.050 5.290 4.310 5.550 ;
        RECT 0.320 4.670 0.580 4.930 ;
        RECT 1.710 4.750 1.970 5.010 ;
        RECT 3.130 4.740 3.390 5.000 ;
        RECT 4.880 4.720 5.140 4.980 ;
        RECT 5.920 4.730 6.180 4.990 ;
        RECT 0.320 4.140 0.580 4.400 ;
        RECT 1.710 4.060 1.970 4.320 ;
        RECT 3.130 4.070 3.390 4.330 ;
        RECT 4.880 4.090 5.140 4.350 ;
        RECT 5.920 4.080 6.180 4.340 ;
        RECT 1.130 3.520 1.390 3.780 ;
        RECT 4.050 3.520 4.310 3.780 ;
        RECT 2.480 3.150 2.740 3.410 ;
        RECT 5.560 3.160 5.820 3.420 ;
        RECT 2.480 2.640 2.740 2.900 ;
        RECT 5.560 2.630 5.820 2.890 ;
        RECT 1.130 2.270 1.390 2.530 ;
        RECT 4.050 2.270 4.310 2.530 ;
        RECT 0.320 1.650 0.580 1.910 ;
        RECT 1.710 1.730 1.970 1.990 ;
        RECT 3.130 1.720 3.390 1.980 ;
        RECT 4.880 1.700 5.140 1.960 ;
        RECT 5.920 1.710 6.180 1.970 ;
        RECT 0.320 1.120 0.580 1.380 ;
        RECT 1.710 1.040 1.970 1.300 ;
        RECT 3.130 1.050 3.390 1.310 ;
        RECT 4.880 1.070 5.140 1.330 ;
        RECT 5.920 1.060 6.180 1.320 ;
        RECT 1.130 0.500 1.390 0.760 ;
        RECT 4.050 0.500 4.310 0.760 ;
        RECT 2.480 0.130 2.740 0.390 ;
        RECT 5.560 0.140 5.820 0.400 ;
  END
END sky130_hilas_Tgate4Double01

MACRO sky130_hilas_cellAttempt01
  CLASS CORE ;
  FOREIGN sky130_hilas_cellAttempt01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.240 BY 10.490 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 0.350 0.000 0.750 6.500 ;
    END
  END VTUN
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 9.550 6.220 9.710 6.270 ;
    END
  END VINJ
  PIN COLSEL1
    PORT
      LAYER met1 ;
        RECT 9.110 6.220 9.300 6.270 ;
    END
  END COLSEL1
  PIN COL1
    PORT
      LAYER met1 ;
        RECT 8.740 6.230 8.900 6.270 ;
    END
  END COL1
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT 4.400 6.170 4.780 6.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.400 0.000 4.780 0.600 ;
    END
  END GATE1
  PIN ROW4
    PORT
      LAYER met2 ;
        RECT 0.000 0.990 7.620 1.170 ;
    END
  END ROW4
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 2.750 1.780 3.070 1.790 ;
        RECT 6.680 1.780 7.000 1.840 ;
        RECT 2.750 1.600 7.000 1.780 ;
        RECT 2.750 1.530 3.070 1.600 ;
        RECT 6.680 1.550 7.000 1.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.720 5.110 6.960 6.500 ;
        RECT 6.700 4.450 6.970 5.110 ;
        RECT 6.720 1.860 6.960 4.450 ;
        RECT 6.710 1.540 6.970 1.860 ;
        RECT 6.720 0.000 6.960 1.540 ;
      LAYER via ;
        RECT 6.710 1.570 6.970 1.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.790 5.090 3.030 6.500 ;
        RECT 2.780 4.430 3.040 5.090 ;
        RECT 2.790 1.820 3.030 4.430 ;
        RECT 2.780 1.500 3.040 1.820 ;
        RECT 2.790 0.000 3.030 1.500 ;
      LAYER via ;
        RECT 2.780 1.530 3.040 1.790 ;
    END
  END VGND
  PIN DRAIN4
    PORT
      LAYER met2 ;
        RECT 0.000 0.570 7.600 0.740 ;
    END
  END DRAIN4
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 0.000 5.760 7.630 5.940 ;
    END
  END DRAIN1
  PIN ROW1
    PORT
      LAYER met2 ;
        RECT 0.000 5.320 7.630 5.500 ;
    END
  END ROW1
  PIN ROW3
    PORT
      LAYER met2 ;
        RECT 0.000 2.090 7.630 2.270 ;
    END
  END ROW3
  PIN DRAIN3
    PORT
      LAYER met2 ;
        RECT 0.000 2.520 7.620 2.700 ;
    END
  END DRAIN3
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 0.000 3.790 7.630 3.970 ;
    END
  END DRAIN2
  PIN ROW2
    PORT
      LAYER met2 ;
        RECT 0.000 4.220 7.630 4.400 ;
    END
  END ROW2
  OBS
      LAYER nwell ;
        RECT 14.510 10.440 16.240 10.490 ;
        RECT 0.000 5.160 0.070 5.340 ;
        RECT 10.400 5.000 12.960 6.910 ;
        RECT 0.570 4.810 1.160 4.920 ;
        RECT 4.310 4.750 5.420 4.980 ;
        RECT 8.950 3.320 9.300 3.330 ;
        RECT 8.950 3.160 9.120 3.320 ;
        RECT 9.290 3.160 9.300 3.320 ;
        RECT 0.570 1.530 1.160 1.720 ;
        RECT 4.310 1.510 5.420 1.780 ;
        RECT 10.400 1.760 12.960 4.730 ;
        RECT 13.320 4.000 16.240 10.440 ;
        RECT 13.320 3.950 15.550 4.000 ;
        RECT 10.400 0.000 12.960 1.500 ;
      LAYER li1 ;
        RECT 14.900 7.430 15.450 7.860 ;
        RECT 10.640 6.560 10.960 6.600 ;
        RECT 10.640 6.440 10.970 6.560 ;
        RECT 10.640 6.340 11.080 6.440 ;
        RECT 10.740 6.270 11.080 6.340 ;
        RECT 12.360 6.170 12.560 6.520 ;
        RECT 10.640 6.010 10.960 6.050 ;
        RECT 10.640 5.820 10.970 6.010 ;
        RECT 10.640 5.790 11.080 5.820 ;
        RECT 10.740 5.650 11.080 5.790 ;
        RECT 11.630 5.550 11.830 6.150 ;
        RECT 12.360 6.140 12.570 6.170 ;
        RECT 12.350 5.550 12.570 6.140 ;
        RECT 2.820 4.520 2.990 5.050 ;
        RECT 6.760 4.510 6.930 5.040 ;
        RECT 10.740 3.940 11.080 4.080 ;
        RECT 10.640 3.910 11.080 3.940 ;
        RECT 2.830 2.810 3.000 3.820 ;
        RECT 10.640 3.720 10.970 3.910 ;
        RECT 10.640 3.680 10.960 3.720 ;
        RECT 6.760 2.670 6.930 3.680 ;
        RECT 11.630 3.580 11.830 4.180 ;
        RECT 12.350 3.590 12.570 4.180 ;
        RECT 12.360 3.560 12.570 3.590 ;
        RECT 10.740 3.390 11.080 3.460 ;
        RECT 8.860 3.160 9.300 3.330 ;
        RECT 10.640 3.290 11.080 3.390 ;
        RECT 10.640 3.200 10.970 3.290 ;
        RECT 10.640 3.100 11.080 3.200 ;
        RECT 10.740 3.030 11.080 3.100 ;
        RECT 12.360 2.930 12.560 3.560 ;
        RECT 10.640 2.770 10.960 2.810 ;
        RECT 10.640 2.580 10.970 2.770 ;
        RECT 10.640 2.550 11.080 2.580 ;
        RECT 10.740 2.410 11.080 2.550 ;
        RECT 11.630 2.310 11.830 2.910 ;
        RECT 12.360 2.900 12.570 2.930 ;
        RECT 12.350 2.310 12.570 2.900 ;
        RECT 10.740 0.710 11.080 0.850 ;
        RECT 10.640 0.680 11.080 0.710 ;
        RECT 10.640 0.490 10.970 0.680 ;
        RECT 10.640 0.450 10.960 0.490 ;
        RECT 11.630 0.350 11.830 0.950 ;
        RECT 12.350 0.360 12.570 0.950 ;
        RECT 12.360 0.330 12.570 0.360 ;
        RECT 10.740 0.160 11.080 0.230 ;
        RECT 10.640 0.060 11.080 0.160 ;
        RECT 10.640 0.000 10.970 0.060 ;
        RECT 12.360 0.000 12.560 0.330 ;
      LAYER mcon ;
        RECT 14.900 7.510 15.170 7.780 ;
        RECT 10.700 6.380 10.870 6.550 ;
        RECT 10.700 5.830 10.870 6.000 ;
        RECT 11.640 5.940 11.810 6.110 ;
        RECT 12.370 5.970 12.540 6.140 ;
        RECT 2.820 4.880 2.990 5.050 ;
        RECT 6.760 4.870 6.930 5.040 ;
        RECT 10.700 3.730 10.870 3.900 ;
        RECT 2.830 3.420 3.000 3.590 ;
        RECT 2.830 3.060 3.000 3.230 ;
        RECT 11.640 3.620 11.810 3.790 ;
        RECT 12.370 3.590 12.540 3.760 ;
        RECT 6.760 3.280 6.930 3.450 ;
        RECT 9.120 3.160 9.300 3.330 ;
        RECT 10.700 3.140 10.870 3.350 ;
        RECT 6.760 2.920 6.930 3.090 ;
        RECT 10.700 2.590 10.870 2.760 ;
        RECT 11.640 2.700 11.810 2.870 ;
        RECT 12.370 2.730 12.540 2.900 ;
        RECT 10.700 0.500 10.870 0.670 ;
        RECT 11.640 0.390 11.810 0.560 ;
        RECT 12.370 0.360 12.540 0.530 ;
        RECT 10.700 0.000 10.870 0.120 ;
      LAYER met1 ;
        RECT 10.630 6.310 10.950 6.630 ;
        RECT 11.630 6.170 11.790 6.900 ;
        RECT 11.630 6.150 11.830 6.170 ;
        RECT 10.630 5.760 10.950 6.080 ;
        RECT 11.610 5.910 11.840 6.150 ;
        RECT 11.630 5.860 11.840 5.910 ;
        RECT 12.000 5.860 12.190 6.850 ;
        RECT 12.440 6.200 12.600 6.900 ;
        RECT 11.630 5.000 11.790 5.860 ;
        RECT 12.020 5.740 12.190 5.860 ;
        RECT 12.030 5.000 12.190 5.740 ;
        RECT 12.330 5.650 12.600 6.200 ;
        RECT 12.330 5.600 12.610 5.650 ;
        RECT 12.440 5.510 12.610 5.600 ;
        RECT 12.440 5.000 12.600 5.510 ;
        RECT 10.630 3.650 10.950 3.970 ;
        RECT 11.630 3.870 11.790 4.730 ;
        RECT 12.030 3.990 12.190 4.730 ;
        RECT 12.440 4.220 12.600 4.730 ;
        RECT 12.440 4.130 12.610 4.220 ;
        RECT 12.020 3.870 12.190 3.990 ;
        RECT 11.630 3.820 11.840 3.870 ;
        RECT 11.610 3.580 11.840 3.820 ;
        RECT 11.630 3.560 11.830 3.580 ;
        RECT 9.170 3.360 9.300 3.380 ;
        RECT 9.090 3.340 9.330 3.360 ;
        RECT 8.890 3.150 9.330 3.340 ;
        RECT 9.090 3.130 9.330 3.150 ;
        RECT 9.190 3.090 9.300 3.130 ;
        RECT 10.630 3.070 10.950 3.420 ;
        RECT 11.630 2.930 11.790 3.560 ;
        RECT 11.630 2.910 11.830 2.930 ;
        RECT 10.630 2.520 10.950 2.840 ;
        RECT 11.610 2.670 11.840 2.910 ;
        RECT 11.630 2.620 11.840 2.670 ;
        RECT 12.000 2.620 12.190 3.870 ;
        RECT 12.330 4.080 12.610 4.130 ;
        RECT 12.330 3.530 12.600 4.080 ;
        RECT 13.970 3.950 14.350 10.450 ;
        RECT 14.840 6.970 15.230 8.830 ;
        RECT 12.440 2.960 12.600 3.530 ;
        RECT 11.630 1.760 11.790 2.620 ;
        RECT 12.020 2.500 12.190 2.620 ;
        RECT 12.030 1.760 12.190 2.500 ;
        RECT 12.330 2.410 12.600 2.960 ;
        RECT 12.330 2.360 12.610 2.410 ;
        RECT 12.440 2.270 12.610 2.360 ;
        RECT 12.440 1.760 12.600 2.270 ;
        RECT 10.630 0.420 10.950 0.740 ;
        RECT 11.630 0.640 11.790 1.500 ;
        RECT 12.030 0.760 12.190 1.500 ;
        RECT 12.440 0.990 12.600 1.500 ;
        RECT 12.440 0.900 12.610 0.990 ;
        RECT 12.020 0.640 12.190 0.760 ;
        RECT 11.630 0.590 11.840 0.640 ;
        RECT 11.610 0.350 11.840 0.590 ;
        RECT 11.630 0.330 11.830 0.350 ;
        RECT 10.630 0.000 10.950 0.190 ;
        RECT 11.630 0.000 11.790 0.330 ;
        RECT 12.000 0.000 12.190 0.640 ;
        RECT 12.330 0.850 12.610 0.900 ;
        RECT 12.330 0.300 12.600 0.850 ;
        RECT 12.440 0.000 12.600 0.300 ;
      LAYER via ;
        RECT 10.660 6.340 10.920 6.600 ;
        RECT 10.660 5.790 10.920 6.050 ;
        RECT 10.660 3.680 10.920 3.940 ;
        RECT 10.660 3.100 10.920 3.390 ;
        RECT 10.660 2.550 10.920 2.810 ;
        RECT 10.660 0.450 10.920 0.710 ;
        RECT 10.660 0.000 10.920 0.160 ;
      LAYER met2 ;
        RECT 10.630 6.350 10.940 6.640 ;
        RECT 10.630 6.310 12.960 6.350 ;
        RECT 10.780 6.170 12.960 6.310 ;
        RECT 10.630 5.920 10.940 6.090 ;
        RECT 10.400 5.740 10.490 5.920 ;
        RECT 10.630 5.760 12.960 5.920 ;
        RECT 10.790 5.740 12.960 5.760 ;
        RECT 10.400 3.810 10.490 3.990 ;
        RECT 10.790 3.970 12.960 3.990 ;
        RECT 10.630 3.810 12.960 3.970 ;
        RECT 10.630 3.640 10.940 3.810 ;
        RECT 10.780 3.420 12.960 3.560 ;
        RECT 10.630 3.380 12.960 3.420 ;
        RECT 10.630 3.110 10.940 3.380 ;
        RECT 10.630 3.070 12.960 3.110 ;
        RECT 10.780 2.930 12.960 3.070 ;
        RECT 10.630 2.680 10.940 2.850 ;
        RECT 10.400 2.500 10.490 2.680 ;
        RECT 10.630 2.520 12.960 2.680 ;
        RECT 10.790 2.500 12.960 2.520 ;
        RECT 10.400 0.580 10.490 0.760 ;
        RECT 10.790 0.740 12.960 0.760 ;
        RECT 10.630 0.580 12.960 0.740 ;
        RECT 10.630 0.410 10.940 0.580 ;
        RECT 10.780 0.190 12.960 0.330 ;
        RECT 10.630 0.150 12.960 0.190 ;
        RECT 10.630 0.000 10.940 0.150 ;
  END
END sky130_hilas_cellAttempt01

MACRO sky130_hilas_StepUpDigital
  CLASS CORE ;
  FOREIGN sky130_hilas_StepUpDigital ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.700 BY 1.750 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 0.000 0.000 2.500 1.750 ;
        RECT 3.590 0.580 5.360 1.750 ;
        RECT 6.370 1.680 8.140 1.750 ;
        RECT 6.370 0.000 8.140 0.090 ;
      LAYER li1 ;
        RECT 0.000 1.730 1.090 1.750 ;
        RECT 0.000 1.560 1.130 1.730 ;
        RECT 1.580 1.700 2.040 1.730 ;
        RECT 3.350 1.700 3.700 1.750 ;
        RECT 1.580 1.560 2.690 1.700 ;
        RECT 1.870 1.530 2.690 1.560 ;
        RECT 2.930 1.530 4.100 1.700 ;
        RECT 4.350 1.530 5.110 1.700 ;
        RECT 1.870 1.390 2.130 1.530 ;
        RECT 0.340 1.060 0.670 1.230 ;
        RECT 0.950 1.220 2.130 1.390 ;
        RECT 4.880 1.520 5.110 1.530 ;
        RECT 0.950 1.070 1.730 1.220 ;
        RECT 1.870 1.080 2.130 1.220 ;
        RECT 2.430 1.290 2.720 1.320 ;
        RECT 2.430 1.120 2.760 1.290 ;
        RECT 2.430 1.080 2.720 1.120 ;
        RECT 3.340 1.080 3.670 1.340 ;
        RECT 4.880 1.080 5.150 1.520 ;
        RECT 0.000 0.880 0.400 1.050 ;
        RECT 0.410 0.600 0.590 1.060 ;
        RECT 0.950 0.780 1.130 1.070 ;
        RECT 1.370 0.720 1.580 1.050 ;
        RECT 1.870 0.910 2.200 1.080 ;
        RECT 2.440 0.910 4.600 1.080 ;
        RECT 1.870 0.860 2.100 0.910 ;
        RECT 4.850 0.900 5.180 1.080 ;
        RECT 5.530 0.940 5.700 1.000 ;
        RECT 1.930 0.630 2.100 0.860 ;
        RECT 5.510 0.720 5.730 0.940 ;
        RECT 5.530 0.670 5.700 0.720 ;
        RECT 1.930 0.620 2.310 0.630 ;
        RECT 0.410 0.430 1.370 0.600 ;
        RECT 1.840 0.560 2.310 0.620 ;
        RECT 1.840 0.510 2.650 0.560 ;
        RECT 1.840 0.450 2.660 0.510 ;
        RECT 1.920 0.390 2.660 0.450 ;
        RECT 1.920 0.340 2.310 0.390 ;
      LAYER mcon ;
        RECT 3.410 1.570 3.620 1.750 ;
        RECT 1.450 1.140 1.620 1.310 ;
        RECT 2.490 1.100 2.660 1.270 ;
        RECT 4.920 1.200 5.090 1.370 ;
        RECT 0.410 0.800 0.580 0.970 ;
        RECT 0.410 0.440 0.580 0.610 ;
      LAYER met1 ;
        RECT 0.340 0.000 0.630 1.750 ;
        RECT 1.380 1.110 1.700 1.390 ;
        RECT 1.340 1.090 1.700 1.110 ;
        RECT 1.340 0.780 1.620 1.090 ;
        RECT 1.870 0.490 2.180 1.750 ;
        RECT 3.350 1.530 3.700 1.750 ;
        RECT 4.650 1.690 5.120 1.750 ;
        RECT 3.500 1.510 3.700 1.530 ;
        RECT 2.430 1.320 2.740 1.330 ;
        RECT 2.420 1.050 2.740 1.320 ;
        RECT 2.430 1.040 2.720 1.050 ;
        RECT 4.880 0.490 5.120 1.690 ;
        RECT 7.660 1.680 7.900 1.750 ;
        RECT 5.450 0.670 5.860 1.000 ;
      LAYER via ;
        RECT 1.410 1.100 1.670 1.360 ;
        RECT 1.350 0.820 1.610 1.080 ;
        RECT 3.390 1.540 3.650 1.750 ;
        RECT 2.450 1.060 2.710 1.320 ;
        RECT 5.490 0.700 5.750 0.960 ;
      LAYER met2 ;
        RECT 1.380 1.310 1.700 1.360 ;
        RECT 2.410 1.320 2.730 1.330 ;
        RECT 2.410 1.310 2.740 1.320 ;
        RECT 0.070 1.110 2.740 1.310 ;
        RECT 1.380 1.100 1.700 1.110 ;
        RECT 1.310 1.030 1.650 1.090 ;
        RECT 2.410 1.060 2.740 1.110 ;
        RECT 2.410 1.040 2.730 1.060 ;
        RECT 3.390 1.030 3.650 1.750 ;
        RECT 1.310 0.810 3.750 1.030 ;
        RECT 5.460 0.670 5.920 0.990 ;
  END
END sky130_hilas_StepUpDigital

MACRO sky130_hilas_VinjNOR3
  CLASS CORE ;
  FOREIGN sky130_hilas_VinjNOR3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.880 BY 1.640 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 0.010 0.000 3.450 1.640 ;
      LAYER li1 ;
        RECT 0.630 1.210 0.800 1.350 ;
        RECT 1.360 1.230 1.530 1.310 ;
        RECT 2.170 1.230 2.340 1.310 ;
        RECT 3.710 1.270 3.880 1.390 ;
        RECT 0.630 1.040 0.820 1.210 ;
        RECT 0.630 0.940 0.800 1.040 ;
        RECT 1.360 0.660 1.570 1.230 ;
        RECT 2.130 0.980 2.340 1.230 ;
        RECT 2.730 1.050 2.900 1.150 ;
        RECT 3.670 1.100 3.880 1.270 ;
        RECT 5.600 1.200 5.860 1.270 ;
        RECT 6.400 1.200 6.580 1.330 ;
        RECT 3.710 1.060 3.880 1.100 ;
        RECT 2.130 0.660 2.300 0.980 ;
        RECT 2.700 0.880 2.900 1.050 ;
        RECT 2.730 0.780 2.900 0.880 ;
        RECT 4.270 1.020 5.140 1.190 ;
        RECT 5.600 1.020 6.580 1.200 ;
        RECT 0.200 0.560 0.370 0.660 ;
        RECT 0.180 0.390 0.370 0.560 ;
        RECT 0.200 0.330 0.370 0.390 ;
        RECT 0.620 0.600 0.790 0.660 ;
        RECT 0.620 0.330 0.870 0.600 ;
        RECT 1.360 0.410 1.610 0.660 ;
        RECT 0.630 0.310 0.870 0.330 ;
        RECT 1.440 0.320 1.610 0.410 ;
        RECT 2.090 0.410 2.300 0.660 ;
        RECT 4.270 0.580 4.440 1.020 ;
        RECT 5.600 0.580 5.860 1.020 ;
        RECT 6.400 0.910 6.580 1.020 ;
        RECT 2.810 0.410 4.440 0.580 ;
        RECT 4.890 0.410 5.860 0.580 ;
        RECT 6.310 0.410 6.650 0.580 ;
        RECT 2.090 0.330 2.260 0.410 ;
        RECT 3.580 0.370 3.750 0.410 ;
      LAYER mcon ;
        RECT 0.650 1.040 0.820 1.210 ;
        RECT 0.660 0.360 0.830 0.530 ;
        RECT 5.630 0.700 5.810 0.880 ;
      LAYER met1 ;
        RECT 0.620 1.260 0.840 1.600 ;
        RECT 0.620 1.000 0.850 1.260 ;
        RECT 0.090 0.320 0.400 0.670 ;
        RECT 0.620 0.600 0.840 1.000 ;
        RECT 2.640 0.840 2.970 1.100 ;
        RECT 3.610 1.060 4.040 1.350 ;
        RECT 0.620 0.290 0.870 0.600 ;
        RECT 3.480 0.310 3.870 0.580 ;
        RECT 0.620 0.090 0.840 0.290 ;
        RECT 5.590 0.090 5.860 1.610 ;
        RECT 6.410 0.320 6.720 0.640 ;
      LAYER via ;
        RECT 0.120 0.350 0.380 0.610 ;
        RECT 2.680 0.840 2.940 1.100 ;
        RECT 3.670 1.090 3.930 1.350 ;
        RECT 3.540 0.310 3.800 0.570 ;
        RECT 6.440 0.350 6.700 0.610 ;
      LAYER met2 ;
        RECT 0.000 1.290 4.040 1.450 ;
        RECT 2.640 1.020 2.970 1.100 ;
        RECT 3.620 1.060 4.040 1.290 ;
        RECT 2.370 1.000 2.970 1.020 ;
        RECT 0.010 0.840 2.970 1.000 ;
        RECT 0.090 0.510 0.410 0.610 ;
        RECT 0.010 0.350 0.410 0.510 ;
        RECT 3.500 0.490 3.870 0.570 ;
        RECT 3.500 0.480 4.530 0.490 ;
        RECT 6.410 0.480 6.720 0.640 ;
        RECT 3.500 0.310 6.880 0.480 ;
  END
END sky130_hilas_VinjNOR3

MACRO sky130_hilas_VinjDiodeProtect01
  CLASS CORE ;
  FOREIGN sky130_hilas_VinjDiodeProtect01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.590 BY 10.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN OUTPUT 
    ANTENNADIFFAREA 58.900799 ;
    PORT
      LAYER met1 ;
        RECT 14.350 10.250 14.700 10.410 ;
        RECT 14.340 9.300 14.710 10.250 ;
        RECT 13.990 8.930 16.460 9.300 ;
        RECT 12.550 7.470 16.460 8.930 ;
        RECT 2.840 7.460 16.460 7.470 ;
        RECT 2.170 6.900 16.460 7.460 ;
        RECT 2.170 2.600 25.520 6.900 ;
        RECT 2.170 2.320 16.460 2.600 ;
        RECT 12.550 0.770 16.460 2.320 ;
        RECT 12.530 0.000 16.480 0.770 ;
    END
  END OUTPUT 
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.000 7.380 28.590 8.780 ;
        RECT 0.470 7.370 1.400 7.380 ;
        RECT 0.720 6.260 0.890 7.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.440 8.130 2.810 8.760 ;
        RECT 23.780 8.280 27.910 8.680 ;
        RECT 23.780 8.190 27.920 8.280 ;
        RECT 0.470 6.170 1.420 8.130 ;
        RECT 2.170 8.110 2.750 8.130 ;
        RECT 27.390 7.290 27.920 8.190 ;
        RECT 0.700 0.500 1.420 6.170 ;
      LAYER via ;
        RECT 0.660 8.280 2.690 8.610 ;
        RECT 24.050 8.280 27.040 8.630 ;
        RECT 0.600 7.420 1.300 8.040 ;
        RECT 27.480 7.480 27.830 8.240 ;
    END
  END VGND
  PIN VINJ
    ANTENNADIFFAREA 9.088799 ;
    PORT
      LAYER nwell ;
        RECT 14.870 1.910 26.920 7.850 ;
      LAYER met2 ;
        RECT 26.340 2.480 26.980 5.490 ;
        RECT 0.000 1.080 28.590 2.480 ;
        RECT 25.440 0.950 28.070 1.080 ;
        RECT 25.440 0.440 27.990 0.950 ;
        RECT 25.440 0.370 26.060 0.440 ;
    END
  END VINJ
  PIN INPUT
    PORT
      LAYER met1 ;
        RECT 7.710 10.280 11.610 10.870 ;
        RECT 7.710 8.930 8.000 10.280 ;
    END
  END INPUT
  OBS
      LAYER li1 ;
        RECT 7.730 8.930 7.980 10.390 ;
        RECT 7.770 8.920 7.940 8.930 ;
        RECT 14.410 8.900 14.660 10.380 ;
        RECT 0.550 8.180 27.930 8.690 ;
        RECT 0.550 6.250 1.350 8.180 ;
        RECT 1.930 7.730 2.100 7.810 ;
        RECT 13.170 7.730 13.400 7.820 ;
        RECT 1.930 7.720 13.400 7.730 ;
        RECT 0.550 1.670 1.060 6.250 ;
        RECT 1.920 2.250 13.400 7.720 ;
        RECT 1.850 2.080 13.400 2.250 ;
        RECT 1.920 2.020 2.110 2.080 ;
        RECT 13.170 1.840 13.400 2.080 ;
        RECT 1.800 1.670 3.600 1.680 ;
        RECT 13.960 1.670 14.470 8.180 ;
        RECT 15.230 7.290 26.480 7.460 ;
        RECT 15.230 2.420 15.400 7.290 ;
        RECT 15.790 6.960 25.900 6.980 ;
        RECT 15.790 6.920 25.920 6.960 ;
        RECT 15.740 6.750 25.920 6.920 ;
        RECT 15.790 2.730 25.920 6.750 ;
        RECT 26.310 5.530 26.480 7.290 ;
        RECT 15.790 2.650 25.900 2.730 ;
        RECT 15.220 2.350 15.400 2.420 ;
        RECT 26.310 2.350 26.920 5.530 ;
        RECT 15.220 2.180 26.920 2.350 ;
        RECT 26.380 2.070 26.920 2.180 ;
        RECT 27.380 1.830 27.930 8.180 ;
        RECT 27.370 1.670 27.930 1.830 ;
        RECT 0.550 1.330 27.930 1.670 ;
        RECT 0.580 1.160 27.930 1.330 ;
        RECT 0.580 1.140 1.270 1.160 ;
        RECT 1.780 1.150 3.580 1.160 ;
      LAYER mcon ;
        RECT 7.770 9.870 7.940 10.040 ;
        RECT 7.770 9.510 7.940 9.680 ;
        RECT 7.770 9.140 7.940 9.310 ;
        RECT 14.450 10.190 14.620 10.360 ;
        RECT 14.450 9.830 14.620 10.000 ;
        RECT 14.450 9.470 14.620 9.640 ;
        RECT 14.450 9.110 14.620 9.280 ;
        RECT 0.630 8.520 2.490 8.530 ;
        RECT 0.630 8.350 2.500 8.520 ;
        RECT 23.990 8.340 27.150 8.520 ;
        RECT 0.670 6.260 0.850 8.160 ;
        RECT 1.070 6.250 1.250 8.160 ;
        RECT 2.260 7.220 13.240 7.390 ;
        RECT 2.260 6.600 13.240 6.770 ;
        RECT 2.270 5.980 13.250 6.150 ;
        RECT 2.290 5.400 13.270 5.570 ;
        RECT 2.300 4.810 13.280 4.980 ;
        RECT 2.300 4.210 13.280 4.380 ;
        RECT 2.250 3.610 13.230 3.780 ;
        RECT 2.260 3.000 13.240 3.170 ;
        RECT 2.250 2.400 13.230 2.570 ;
        RECT 15.990 6.460 25.440 6.630 ;
        RECT 15.980 5.710 25.370 5.880 ;
        RECT 16.010 4.990 25.410 5.160 ;
        RECT 16.020 4.330 25.390 4.500 ;
        RECT 16.010 3.680 25.460 3.850 ;
        RECT 16.020 3.040 25.410 3.210 ;
        RECT 27.560 7.360 27.760 8.290 ;
        RECT 26.490 2.120 26.840 5.420 ;
      LAYER met1 ;
        RECT 26.290 5.480 26.860 5.490 ;
        RECT 26.290 2.060 26.910 5.480 ;
        RECT 26.290 2.050 26.860 2.060 ;
        RECT 25.460 0.420 26.020 0.920 ;
        RECT 25.470 0.200 26.020 0.420 ;
      LAYER via ;
        RECT 26.450 2.190 26.870 5.360 ;
        RECT 25.480 0.370 26.000 0.890 ;
  END
END sky130_hilas_VinjDiodeProtect01

MACRO sky130_hilas_LevelShift4InputUp
  CLASS CORE ;
  FOREIGN sky130_hilas_LevelShift4InputUp ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.700 BY 7.000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 7.660 6.950 7.900 7.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 7.660 0.000 7.900 0.050 ;
    END
  END VPWR
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 0.340 0.000 0.630 0.120 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.000 0.440 2.310 7.000 ;
      LAYER met1 ;
        RECT 0.150 6.910 0.630 7.000 ;
        RECT 0.150 0.440 0.440 6.910 ;
    END
  END VINJ
  PIN OUTPUT1
    PORT
      LAYER met2 ;
        RECT 0.000 6.360 0.160 6.560 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    PORT
      LAYER met2 ;
        RECT 0.000 4.610 0.170 4.810 ;
    END
  END OUTPUT2
  PIN OUTPUT3
    PORT
      LAYER met2 ;
        RECT 0.000 2.860 0.190 3.060 ;
    END
  END OUTPUT3
  PIN OUTPUT4
    PORT
      LAYER met2 ;
        RECT 0.000 1.110 0.160 1.310 ;
    END
  END OUTPUT4
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 4.650 0.000 4.960 0.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.650 6.940 4.960 7.000 ;
        RECT 4.690 6.180 4.930 6.940 ;
    END
  END VGND
  PIN INPUT1
    PORT
      LAYER met2 ;
        RECT 8.600 5.430 8.700 5.750 ;
    END
  END INPUT1
  PIN INPUT2
    PORT
      LAYER met2 ;
        RECT 8.600 3.680 8.700 4.000 ;
    END
  END INPUT2
  PIN INPUT3
    PORT
      LAYER met2 ;
        RECT 8.600 1.930 8.700 2.250 ;
    END
  END INPUT3
  PIN INPUT4
    PORT
      LAYER met2 ;
        RECT 8.600 0.180 8.700 0.500 ;
    END
  END INPUT4
  OBS
      LAYER nwell ;
        RECT 3.400 6.270 5.170 7.000 ;
        RECT 3.400 4.520 5.170 6.110 ;
        RECT 6.180 5.620 7.950 5.780 ;
        RECT 3.400 2.770 5.170 4.360 ;
        RECT 6.180 3.870 7.950 4.030 ;
        RECT 3.400 1.020 5.170 2.610 ;
        RECT 6.180 2.120 7.950 2.280 ;
        RECT 6.180 0.440 7.950 0.530 ;
      LAYER li1 ;
        RECT 0.150 6.750 0.480 6.920 ;
        RECT 0.760 6.910 1.940 7.000 ;
        RECT 0.760 6.760 1.540 6.910 ;
        RECT 1.680 6.770 1.940 6.910 ;
        RECT 2.240 6.980 2.530 7.000 ;
        RECT 2.240 6.810 2.570 6.980 ;
        RECT 2.240 6.770 2.530 6.810 ;
        RECT 3.150 6.770 3.480 7.000 ;
        RECT 4.690 6.770 4.960 7.000 ;
        RECT 0.000 6.570 0.210 6.740 ;
        RECT 0.220 6.290 0.400 6.750 ;
        RECT 0.760 6.470 0.940 6.760 ;
        RECT 1.180 6.410 1.390 6.740 ;
        RECT 1.680 6.600 2.010 6.770 ;
        RECT 2.250 6.600 4.410 6.770 ;
        RECT 1.680 6.550 1.910 6.600 ;
        RECT 4.660 6.590 4.990 6.770 ;
        RECT 5.340 6.630 5.510 6.690 ;
        RECT 1.740 6.320 1.910 6.550 ;
        RECT 5.320 6.410 5.540 6.630 ;
        RECT 5.340 6.360 5.510 6.410 ;
        RECT 1.740 6.310 2.120 6.320 ;
        RECT 0.220 6.120 1.180 6.290 ;
        RECT 1.650 6.250 2.120 6.310 ;
        RECT 1.650 6.200 2.460 6.250 ;
        RECT 1.650 6.140 2.470 6.200 ;
        RECT 1.730 6.080 2.470 6.140 ;
        RECT 1.730 6.030 2.120 6.080 ;
        RECT 0.000 5.670 0.900 5.690 ;
        RECT 0.000 5.500 0.940 5.670 ;
        RECT 1.390 5.640 1.850 5.670 ;
        RECT 3.160 5.640 3.510 5.740 ;
        RECT 1.390 5.500 2.500 5.640 ;
        RECT 1.680 5.470 2.500 5.500 ;
        RECT 2.740 5.470 3.910 5.640 ;
        RECT 4.160 5.470 4.920 5.640 ;
        RECT 1.680 5.330 1.940 5.470 ;
        RECT 0.150 5.000 0.480 5.170 ;
        RECT 0.760 5.160 1.940 5.330 ;
        RECT 4.690 5.460 4.920 5.470 ;
        RECT 0.760 5.010 1.540 5.160 ;
        RECT 1.680 5.020 1.940 5.160 ;
        RECT 2.240 5.230 2.530 5.260 ;
        RECT 2.240 5.060 2.570 5.230 ;
        RECT 2.240 5.020 2.530 5.060 ;
        RECT 3.150 5.020 3.480 5.280 ;
        RECT 4.690 5.020 4.960 5.460 ;
        RECT 0.000 4.820 0.210 4.990 ;
        RECT 0.220 4.540 0.400 5.000 ;
        RECT 0.760 4.720 0.940 5.010 ;
        RECT 1.180 4.660 1.390 4.990 ;
        RECT 1.680 4.850 2.010 5.020 ;
        RECT 2.250 4.850 4.410 5.020 ;
        RECT 1.680 4.800 1.910 4.850 ;
        RECT 4.660 4.840 4.990 5.020 ;
        RECT 5.340 4.880 5.510 4.940 ;
        RECT 1.740 4.570 1.910 4.800 ;
        RECT 5.320 4.660 5.540 4.880 ;
        RECT 5.340 4.610 5.510 4.660 ;
        RECT 1.740 4.560 2.120 4.570 ;
        RECT 0.220 4.370 1.180 4.540 ;
        RECT 1.650 4.500 2.120 4.560 ;
        RECT 1.650 4.450 2.460 4.500 ;
        RECT 1.650 4.390 2.470 4.450 ;
        RECT 1.730 4.330 2.470 4.390 ;
        RECT 1.730 4.280 2.120 4.330 ;
        RECT 0.000 3.920 0.900 3.940 ;
        RECT 0.000 3.750 0.940 3.920 ;
        RECT 1.390 3.890 1.850 3.920 ;
        RECT 3.160 3.890 3.510 3.990 ;
        RECT 1.390 3.750 2.500 3.890 ;
        RECT 1.680 3.720 2.500 3.750 ;
        RECT 2.740 3.720 3.910 3.890 ;
        RECT 4.160 3.720 4.920 3.890 ;
        RECT 1.680 3.580 1.940 3.720 ;
        RECT 0.150 3.250 0.480 3.420 ;
        RECT 0.760 3.410 1.940 3.580 ;
        RECT 4.690 3.710 4.920 3.720 ;
        RECT 0.760 3.260 1.540 3.410 ;
        RECT 1.680 3.270 1.940 3.410 ;
        RECT 2.240 3.480 2.530 3.510 ;
        RECT 2.240 3.310 2.570 3.480 ;
        RECT 2.240 3.270 2.530 3.310 ;
        RECT 3.150 3.270 3.480 3.530 ;
        RECT 4.690 3.270 4.960 3.710 ;
        RECT 0.000 3.070 0.210 3.240 ;
        RECT 0.220 2.790 0.400 3.250 ;
        RECT 0.760 2.970 0.940 3.260 ;
        RECT 1.180 2.910 1.390 3.240 ;
        RECT 1.680 3.100 2.010 3.270 ;
        RECT 2.250 3.100 4.410 3.270 ;
        RECT 1.680 3.050 1.910 3.100 ;
        RECT 4.660 3.090 4.990 3.270 ;
        RECT 5.340 3.130 5.510 3.190 ;
        RECT 1.740 2.820 1.910 3.050 ;
        RECT 5.320 2.910 5.540 3.130 ;
        RECT 5.340 2.860 5.510 2.910 ;
        RECT 1.740 2.810 2.120 2.820 ;
        RECT 0.220 2.620 1.180 2.790 ;
        RECT 1.650 2.750 2.120 2.810 ;
        RECT 1.650 2.700 2.460 2.750 ;
        RECT 1.650 2.640 2.470 2.700 ;
        RECT 1.730 2.580 2.470 2.640 ;
        RECT 1.730 2.530 2.120 2.580 ;
        RECT 0.000 2.170 0.900 2.190 ;
        RECT 0.000 2.000 0.940 2.170 ;
        RECT 1.390 2.140 1.850 2.170 ;
        RECT 3.160 2.140 3.510 2.240 ;
        RECT 1.390 2.000 2.500 2.140 ;
        RECT 1.680 1.970 2.500 2.000 ;
        RECT 2.740 1.970 3.910 2.140 ;
        RECT 4.160 1.970 4.920 2.140 ;
        RECT 1.680 1.830 1.940 1.970 ;
        RECT 0.150 1.500 0.480 1.670 ;
        RECT 0.760 1.660 1.940 1.830 ;
        RECT 4.690 1.960 4.920 1.970 ;
        RECT 0.760 1.510 1.540 1.660 ;
        RECT 1.680 1.520 1.940 1.660 ;
        RECT 2.240 1.730 2.530 1.760 ;
        RECT 2.240 1.560 2.570 1.730 ;
        RECT 2.240 1.520 2.530 1.560 ;
        RECT 3.150 1.520 3.480 1.780 ;
        RECT 4.690 1.520 4.960 1.960 ;
        RECT 0.000 1.320 0.210 1.490 ;
        RECT 0.220 1.040 0.400 1.500 ;
        RECT 0.760 1.220 0.940 1.510 ;
        RECT 1.180 1.160 1.390 1.490 ;
        RECT 1.680 1.350 2.010 1.520 ;
        RECT 2.250 1.350 4.410 1.520 ;
        RECT 1.680 1.300 1.910 1.350 ;
        RECT 4.660 1.340 4.990 1.520 ;
        RECT 5.340 1.380 5.510 1.440 ;
        RECT 1.740 1.070 1.910 1.300 ;
        RECT 5.320 1.160 5.540 1.380 ;
        RECT 5.340 1.110 5.510 1.160 ;
        RECT 1.740 1.060 2.120 1.070 ;
        RECT 0.220 0.870 1.180 1.040 ;
        RECT 1.650 1.000 2.120 1.060 ;
        RECT 1.650 0.950 2.460 1.000 ;
        RECT 1.650 0.890 2.470 0.950 ;
        RECT 1.730 0.830 2.470 0.890 ;
        RECT 1.730 0.780 2.120 0.830 ;
      LAYER mcon ;
        RECT 1.260 6.830 1.430 7.000 ;
        RECT 2.300 6.790 2.470 6.960 ;
        RECT 4.730 6.890 4.900 7.000 ;
        RECT 0.220 6.490 0.390 6.660 ;
        RECT 0.220 6.130 0.390 6.300 ;
        RECT 3.220 5.510 3.430 5.720 ;
        RECT 1.260 5.080 1.430 5.250 ;
        RECT 2.300 5.040 2.470 5.210 ;
        RECT 4.730 5.140 4.900 5.310 ;
        RECT 0.220 4.740 0.390 4.910 ;
        RECT 0.220 4.380 0.390 4.550 ;
        RECT 3.220 3.760 3.430 3.970 ;
        RECT 1.260 3.330 1.430 3.500 ;
        RECT 2.300 3.290 2.470 3.460 ;
        RECT 4.730 3.390 4.900 3.560 ;
        RECT 0.220 2.990 0.390 3.160 ;
        RECT 0.220 2.630 0.390 2.800 ;
        RECT 3.220 2.010 3.430 2.220 ;
        RECT 1.260 1.580 1.430 1.750 ;
        RECT 2.300 1.540 2.470 1.710 ;
        RECT 4.730 1.640 4.900 1.810 ;
        RECT 0.220 1.240 0.390 1.410 ;
        RECT 0.220 0.880 0.390 1.050 ;
      LAYER met1 ;
        RECT 1.190 6.800 1.510 7.000 ;
        RECT 1.150 6.780 1.510 6.800 ;
        RECT 1.150 6.470 1.430 6.780 ;
        RECT 1.680 6.180 1.990 7.000 ;
        RECT 2.230 6.740 2.550 7.000 ;
        RECT 2.240 6.730 2.530 6.740 ;
        RECT 5.260 6.360 5.670 6.690 ;
        RECT 1.190 5.050 1.510 5.330 ;
        RECT 1.150 5.030 1.510 5.050 ;
        RECT 1.150 4.720 1.430 5.030 ;
        RECT 1.680 4.430 1.990 6.120 ;
        RECT 3.160 5.470 3.510 5.760 ;
        RECT 4.690 5.690 4.930 6.110 ;
        RECT 4.460 5.630 4.930 5.690 ;
        RECT 3.310 5.450 3.510 5.470 ;
        RECT 2.240 5.260 2.550 5.270 ;
        RECT 2.230 4.990 2.550 5.260 ;
        RECT 2.240 4.980 2.530 4.990 ;
        RECT 4.690 4.430 4.930 5.630 ;
        RECT 7.470 5.620 7.710 5.690 ;
        RECT 5.260 4.610 5.670 4.940 ;
        RECT 1.190 3.300 1.510 3.580 ;
        RECT 1.150 3.280 1.510 3.300 ;
        RECT 1.150 2.970 1.430 3.280 ;
        RECT 1.680 2.680 1.990 4.370 ;
        RECT 3.160 3.720 3.510 4.010 ;
        RECT 4.690 3.940 4.930 4.360 ;
        RECT 4.460 3.880 4.930 3.940 ;
        RECT 3.310 3.700 3.510 3.720 ;
        RECT 2.240 3.510 2.550 3.520 ;
        RECT 2.230 3.240 2.550 3.510 ;
        RECT 2.240 3.230 2.530 3.240 ;
        RECT 4.690 2.680 4.930 3.880 ;
        RECT 7.470 3.870 7.710 3.940 ;
        RECT 5.260 2.860 5.670 3.190 ;
        RECT 1.190 1.550 1.510 1.830 ;
        RECT 1.150 1.530 1.510 1.550 ;
        RECT 1.150 1.220 1.430 1.530 ;
        RECT 1.680 0.930 1.990 2.620 ;
        RECT 3.160 1.970 3.510 2.260 ;
        RECT 4.690 2.190 4.930 2.610 ;
        RECT 4.460 2.130 4.930 2.190 ;
        RECT 3.310 1.950 3.510 1.970 ;
        RECT 2.240 1.760 2.550 1.770 ;
        RECT 2.230 1.490 2.550 1.760 ;
        RECT 2.240 1.480 2.530 1.490 ;
        RECT 4.690 0.930 4.930 2.130 ;
        RECT 7.470 2.120 7.710 2.190 ;
        RECT 5.260 1.110 5.670 1.440 ;
      LAYER via ;
        RECT 1.220 6.790 1.480 7.000 ;
        RECT 1.160 6.510 1.420 6.770 ;
        RECT 2.260 6.750 2.520 7.000 ;
        RECT 5.300 6.390 5.560 6.650 ;
        RECT 1.220 5.040 1.480 5.300 ;
        RECT 1.160 4.760 1.420 5.020 ;
        RECT 3.200 5.480 3.460 5.740 ;
        RECT 2.260 5.000 2.520 5.260 ;
        RECT 5.300 4.640 5.560 4.900 ;
        RECT 1.220 3.290 1.480 3.550 ;
        RECT 1.160 3.010 1.420 3.270 ;
        RECT 3.200 3.730 3.460 3.990 ;
        RECT 2.260 3.250 2.520 3.510 ;
        RECT 5.300 2.890 5.560 3.150 ;
        RECT 1.220 1.540 1.480 1.800 ;
        RECT 1.160 1.260 1.420 1.520 ;
        RECT 3.200 1.980 3.460 2.240 ;
        RECT 2.260 1.500 2.520 1.760 ;
        RECT 5.300 1.140 5.560 1.400 ;
      LAYER met2 ;
        RECT 0.000 6.800 2.550 7.000 ;
        RECT 1.190 6.790 1.510 6.800 ;
        RECT 1.120 6.720 1.460 6.780 ;
        RECT 2.220 6.750 2.550 6.800 ;
        RECT 2.220 6.730 2.540 6.750 ;
        RECT 3.200 6.720 3.460 7.000 ;
        RECT 1.120 6.500 3.560 6.720 ;
        RECT 5.270 6.360 5.730 6.680 ;
        RECT 1.190 5.250 1.510 5.300 ;
        RECT 2.220 5.260 2.540 5.270 ;
        RECT 2.220 5.250 2.550 5.260 ;
        RECT 0.000 5.050 2.550 5.250 ;
        RECT 1.190 5.040 1.510 5.050 ;
        RECT 1.120 4.970 1.460 5.030 ;
        RECT 2.220 5.000 2.550 5.050 ;
        RECT 2.220 4.980 2.540 5.000 ;
        RECT 3.200 4.970 3.460 5.770 ;
        RECT 1.120 4.750 3.560 4.970 ;
        RECT 5.270 4.610 5.730 4.930 ;
        RECT 1.190 3.500 1.510 3.550 ;
        RECT 2.220 3.510 2.540 3.520 ;
        RECT 2.220 3.500 2.550 3.510 ;
        RECT 0.000 3.300 2.550 3.500 ;
        RECT 1.190 3.290 1.510 3.300 ;
        RECT 1.120 3.220 1.460 3.280 ;
        RECT 2.220 3.250 2.550 3.300 ;
        RECT 2.220 3.230 2.540 3.250 ;
        RECT 3.200 3.220 3.460 4.020 ;
        RECT 1.120 3.000 3.560 3.220 ;
        RECT 5.270 2.860 5.730 3.180 ;
        RECT 1.190 1.750 1.510 1.800 ;
        RECT 2.220 1.760 2.540 1.770 ;
        RECT 2.220 1.750 2.550 1.760 ;
        RECT 0.000 1.550 2.550 1.750 ;
        RECT 1.190 1.540 1.510 1.550 ;
        RECT 1.120 1.470 1.460 1.530 ;
        RECT 2.220 1.500 2.550 1.550 ;
        RECT 2.220 1.480 2.540 1.500 ;
        RECT 3.200 1.470 3.460 2.270 ;
        RECT 1.120 1.250 3.560 1.470 ;
        RECT 5.270 1.110 5.730 1.430 ;
  END
END sky130_hilas_LevelShift4InputUp

MACRO sky130_hilas_WTA4Stage01
  CLASS CORE ;
  FOREIGN sky130_hilas_WTA4Stage01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.740 BY 10.500 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 19.290 1.770 19.620 1.860 ;
        RECT 12.940 1.600 19.620 1.770 ;
        RECT 19.290 1.570 19.620 1.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.350 1.880 19.580 6.230 ;
        RECT 19.310 1.870 19.590 1.880 ;
        RECT 19.310 1.550 19.610 1.870 ;
        RECT 19.350 0.180 19.580 1.550 ;
      LAYER via ;
        RECT 19.320 1.580 19.590 1.850 ;
    END
  END VGND
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 17.450 4.940 19.740 5.030 ;
        RECT 17.300 4.870 19.740 4.940 ;
        RECT 17.300 4.610 17.610 4.870 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 16.240 4.360 17.440 4.420 ;
        RECT 16.240 4.320 17.610 4.360 ;
        RECT 16.230 4.240 17.610 4.320 ;
        RECT 17.160 4.120 17.610 4.240 ;
        RECT 17.160 4.100 17.190 4.120 ;
        RECT 17.300 4.100 17.610 4.120 ;
        RECT 17.300 4.030 19.740 4.100 ;
        RECT 17.450 3.940 19.740 4.030 ;
    END
  END OUTPUT2
  PIN OUTPUT3
    USE ANALOG ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 17.450 2.170 19.740 2.260 ;
        RECT 17.300 2.100 19.740 2.170 ;
        RECT 17.300 1.840 17.610 2.100 ;
    END
  END OUTPUT3
  PIN OUTPUT4
    USE ANALOG ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 17.300 1.330 17.610 1.590 ;
        RECT 17.300 1.260 19.740 1.330 ;
        RECT 17.450 1.170 19.740 1.260 ;
    END
  END OUTPUT4
  PIN INPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 1.267500 ;
    PORT
      LAYER met2 ;
        RECT 8.930 5.920 9.250 5.940 ;
        RECT 6.720 5.700 7.040 5.760 ;
        RECT 8.930 5.730 16.850 5.920 ;
        RECT 8.930 5.710 17.030 5.730 ;
        RECT 8.930 5.700 9.250 5.710 ;
        RECT 10.740 5.700 11.070 5.710 ;
        RECT 6.720 5.530 11.070 5.700 ;
        RECT 6.720 5.480 7.040 5.530 ;
        RECT 10.740 5.470 11.070 5.530 ;
        RECT 16.640 5.520 17.030 5.710 ;
        RECT 5.660 5.170 5.810 5.300 ;
        RECT 3.530 5.150 5.810 5.170 ;
        RECT 3.530 4.990 5.860 5.150 ;
        RECT 5.550 4.880 5.860 4.990 ;
        RECT 8.910 4.880 9.230 4.890 ;
        RECT 5.550 4.820 9.230 4.880 ;
        RECT 5.660 4.740 9.230 4.820 ;
        RECT 3.530 4.730 9.230 4.740 ;
        RECT 3.530 4.600 5.710 4.730 ;
        RECT 8.790 4.630 9.230 4.730 ;
        RECT 3.530 4.560 5.860 4.600 ;
        RECT 5.550 4.400 5.860 4.560 ;
        RECT 5.550 4.270 5.960 4.400 ;
        RECT 5.640 4.130 5.960 4.270 ;
        RECT 8.870 3.650 9.100 3.660 ;
        RECT 8.870 3.620 16.440 3.650 ;
        RECT 8.870 3.450 16.500 3.620 ;
        RECT 5.620 3.350 5.940 3.380 ;
        RECT 8.870 3.350 9.110 3.450 ;
        RECT 5.620 3.170 9.110 3.350 ;
        RECT 16.310 3.250 17.030 3.450 ;
        RECT 16.910 3.240 17.030 3.250 ;
        RECT 5.620 3.150 9.030 3.170 ;
        RECT 5.620 3.120 5.940 3.150 ;
    END
  END INPUT1
  PIN INPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met1 ;
        RECT 5.540 4.420 5.860 4.600 ;
        RECT 5.540 4.280 5.930 4.420 ;
        RECT 5.660 4.100 5.930 4.280 ;
        RECT 5.660 3.410 5.870 4.100 ;
        RECT 5.650 3.090 5.910 3.410 ;
      LAYER via ;
        RECT 5.570 4.390 5.830 4.570 ;
        RECT 5.570 4.310 5.930 4.390 ;
        RECT 5.670 4.130 5.930 4.310 ;
        RECT 5.650 3.120 5.910 3.380 ;
    END
  END INPUT2
  PIN INPUT3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 8.910 2.970 9.230 3.010 ;
        RECT 8.910 2.950 16.460 2.970 ;
        RECT 16.910 2.950 17.030 2.960 ;
        RECT 8.910 2.750 17.030 2.950 ;
        RECT 9.010 2.740 9.330 2.750 ;
        RECT 5.600 1.790 5.800 2.290 ;
        RECT 8.780 1.790 9.100 1.830 ;
        RECT 5.600 1.590 9.150 1.790 ;
        RECT 8.780 1.570 9.100 1.590 ;
    END
  END INPUT3
  PIN INPUT4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.710 1.350 6.020 1.530 ;
        RECT 5.590 1.200 6.020 1.350 ;
        RECT 5.590 1.080 5.870 1.200 ;
        RECT 5.600 0.560 6.170 0.740 ;
        RECT 16.460 0.690 17.010 0.700 ;
        RECT 8.880 0.680 17.010 0.690 ;
        RECT 5.760 0.410 6.070 0.560 ;
        RECT 5.640 0.280 6.070 0.410 ;
        RECT 8.880 0.470 17.030 0.680 ;
        RECT 8.880 0.460 16.470 0.470 ;
        RECT 8.880 0.450 9.650 0.460 ;
        RECT 8.880 0.280 9.120 0.450 ;
        RECT 5.640 0.200 9.120 0.280 ;
        RECT 5.750 0.040 9.120 0.200 ;
    END
  END INPUT4
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 5.620 5.760 6.350 5.940 ;
    END
  END DRAIN1
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT 11.460 6.130 11.840 6.230 ;
    END
  END GATE1
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 15.490 5.950 15.890 6.230 ;
    END
  END VTUN
  PIN WTAMIDDLENODE
    ANTENNAGATEAREA 0.472000 ;
    ANTENNADIFFAREA 0.708000 ;
    PORT
      LAYER met1 ;
        RECT 18.090 0.180 18.320 6.230 ;
    END
  END WTAMIDDLENODE
  PIN COLSEL1
    ANTENNADIFFAREA 0.512300 ;
    PORT
      LAYER met1 ;
        RECT 6.760 6.230 7.010 10.500 ;
        RECT 6.760 6.160 7.130 6.230 ;
        RECT 6.760 5.790 7.010 6.160 ;
        RECT 6.740 5.760 7.020 5.790 ;
        RECT 6.730 5.480 7.030 5.760 ;
        RECT 6.740 5.460 7.020 5.480 ;
        RECT 6.760 4.000 7.010 5.460 ;
      LAYER via ;
        RECT 6.750 5.490 7.010 5.750 ;
    END
  END COLSEL1
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 7.340 6.160 7.500 6.230 ;
    END
  END VPWR
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 6.530 6.160 6.690 6.230 ;
    END
  END VINJ
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 5.590 3.810 6.170 3.990 ;
    END
  END DRAIN2
  PIN DRAIN3
    PORT
      LAYER met2 ;
        RECT 5.620 2.520 6.170 2.700 ;
    END
  END DRAIN3
  OBS
      LAYER nwell ;
        RECT 3.530 6.230 6.090 10.500 ;
        RECT 7.620 6.230 9.850 10.490 ;
        RECT 12.440 8.770 13.030 8.930 ;
        RECT 3.530 6.220 9.850 6.230 ;
        RECT 3.530 6.070 6.180 6.220 ;
        RECT 3.530 6.060 6.360 6.070 ;
        RECT 3.530 4.000 6.180 6.060 ;
        RECT 7.620 4.000 9.850 6.220 ;
        RECT 11.460 6.130 11.840 6.230 ;
        RECT 15.490 6.090 15.890 6.230 ;
        RECT 12.440 5.530 13.030 5.680 ;
        RECT 5.660 3.880 6.180 4.000 ;
        RECT 5.660 3.680 6.170 3.880 ;
        RECT 5.660 3.150 6.180 3.680 ;
        RECT 5.770 0.190 6.180 3.150 ;
      LAYER li1 ;
        RECT 5.530 10.150 5.850 10.190 ;
        RECT 3.930 9.760 4.130 10.110 ;
        RECT 5.520 10.030 5.850 10.150 ;
        RECT 5.410 9.930 5.850 10.030 ;
        RECT 5.410 9.860 5.750 9.930 ;
        RECT 3.920 9.730 4.130 9.760 ;
        RECT 3.920 9.140 4.140 9.730 ;
        RECT 4.660 9.140 4.860 9.740 ;
        RECT 5.530 9.600 5.850 9.640 ;
        RECT 5.520 9.410 5.850 9.600 ;
        RECT 5.410 9.380 5.850 9.410 ;
        RECT 5.410 9.240 5.750 9.380 ;
        RECT 3.920 8.020 4.140 8.610 ;
        RECT 3.920 7.990 4.130 8.020 ;
        RECT 4.660 8.010 4.860 8.610 ;
        RECT 5.410 8.370 5.750 8.510 ;
        RECT 6.800 8.450 6.970 8.980 ;
        RECT 10.820 8.480 10.990 9.010 ;
        RECT 5.410 8.340 5.850 8.370 ;
        RECT 5.520 8.150 5.850 8.340 ;
        RECT 5.530 8.110 5.850 8.150 ;
        RECT 3.930 7.640 4.130 7.990 ;
        RECT 5.410 7.820 5.750 7.890 ;
        RECT 5.410 7.720 5.850 7.820 ;
        RECT 5.520 7.600 5.850 7.720 ;
        RECT 5.530 7.560 5.850 7.600 ;
        RECT 4.300 7.180 4.740 7.350 ;
        RECT 5.530 6.910 5.850 6.950 ;
        RECT 3.930 6.520 4.130 6.870 ;
        RECT 5.520 6.790 5.850 6.910 ;
        RECT 5.410 6.690 5.850 6.790 ;
        RECT 5.410 6.620 5.750 6.690 ;
        RECT 6.790 6.590 6.960 7.780 ;
        RECT 10.810 6.550 10.980 7.720 ;
        RECT 3.920 6.490 4.130 6.520 ;
        RECT 3.920 5.900 4.140 6.490 ;
        RECT 4.660 5.900 4.860 6.500 ;
        RECT 5.530 6.360 5.850 6.400 ;
        RECT 5.520 6.170 5.850 6.360 ;
        RECT 5.410 6.140 5.850 6.170 ;
        RECT 5.410 6.000 5.750 6.140 ;
        RECT 17.350 5.590 18.810 5.710 ;
        RECT 17.160 5.540 18.810 5.590 ;
        RECT 17.160 5.370 17.490 5.540 ;
        RECT 3.920 4.770 4.140 5.360 ;
        RECT 3.920 4.740 4.130 4.770 ;
        RECT 4.660 4.760 4.860 5.360 ;
        RECT 17.160 5.330 17.480 5.370 ;
        RECT 18.640 5.310 18.810 5.540 ;
        RECT 5.410 5.120 5.750 5.260 ;
        RECT 5.410 5.090 5.850 5.120 ;
        RECT 5.520 4.900 5.850 5.090 ;
        RECT 17.490 4.910 17.830 5.310 ;
        RECT 18.000 5.140 18.330 5.310 ;
        RECT 18.550 5.140 18.890 5.310 ;
        RECT 18.080 4.970 18.250 5.140 ;
        RECT 18.640 4.970 18.810 5.140 ;
        RECT 5.530 4.860 5.850 4.900 ;
        RECT 17.310 4.800 17.830 4.910 ;
        RECT 18.000 4.800 18.330 4.970 ;
        RECT 18.550 4.800 18.890 4.970 ;
        RECT 3.930 4.390 4.130 4.740 ;
        RECT 17.310 4.690 17.640 4.800 ;
        RECT 17.310 4.650 17.630 4.690 ;
        RECT 5.410 4.570 5.750 4.640 ;
        RECT 18.080 4.570 18.330 4.800 ;
        RECT 19.210 4.720 19.720 5.390 ;
        RECT 5.410 4.470 5.850 4.570 ;
        RECT 5.520 4.350 5.850 4.470 ;
        RECT 5.530 4.310 5.850 4.350 ;
        RECT 18.080 4.400 18.750 4.570 ;
        RECT 17.310 4.280 17.630 4.320 ;
        RECT 17.310 4.170 17.640 4.280 ;
        RECT 18.080 4.170 18.330 4.400 ;
        RECT 17.310 4.060 17.830 4.170 ;
        RECT 17.490 3.660 17.830 4.060 ;
        RECT 18.000 4.000 18.330 4.170 ;
        RECT 18.550 4.000 18.890 4.170 ;
        RECT 18.080 3.830 18.250 4.000 ;
        RECT 18.640 3.830 18.810 4.000 ;
        RECT 18.000 3.660 18.330 3.830 ;
        RECT 18.550 3.660 18.890 3.830 ;
        RECT 17.160 3.600 17.480 3.640 ;
        RECT 17.160 3.430 17.490 3.600 ;
        RECT 18.640 3.430 18.810 3.660 ;
        RECT 19.210 3.580 19.720 4.250 ;
        RECT 17.160 3.380 18.810 3.430 ;
        RECT 17.350 3.260 18.810 3.380 ;
        RECT 17.350 2.820 18.810 2.940 ;
        RECT 17.160 2.770 18.810 2.820 ;
        RECT 17.160 2.600 17.490 2.770 ;
        RECT 17.160 2.560 17.480 2.600 ;
        RECT 18.640 2.540 18.810 2.770 ;
        RECT 17.490 2.140 17.830 2.540 ;
        RECT 18.000 2.370 18.330 2.540 ;
        RECT 18.550 2.370 18.890 2.540 ;
        RECT 18.080 2.200 18.250 2.370 ;
        RECT 18.640 2.200 18.810 2.370 ;
        RECT 17.310 2.030 17.830 2.140 ;
        RECT 18.000 2.030 18.330 2.200 ;
        RECT 18.550 2.030 18.890 2.200 ;
        RECT 17.310 1.920 17.640 2.030 ;
        RECT 17.310 1.880 17.630 1.920 ;
        RECT 18.080 1.800 18.330 2.030 ;
        RECT 19.210 1.950 19.720 2.620 ;
        RECT 18.080 1.630 18.750 1.800 ;
        RECT 17.310 1.510 17.630 1.550 ;
        RECT 5.720 1.450 6.040 1.490 ;
        RECT 5.720 1.280 6.050 1.450 ;
        RECT 17.310 1.400 17.640 1.510 ;
        RECT 18.080 1.400 18.330 1.630 ;
        RECT 17.310 1.290 17.830 1.400 ;
        RECT 5.630 1.260 6.050 1.280 ;
        RECT 5.630 1.230 6.040 1.260 ;
        RECT 5.630 0.530 5.810 1.230 ;
        RECT 17.490 0.890 17.830 1.290 ;
        RECT 18.000 1.230 18.330 1.400 ;
        RECT 18.550 1.230 18.890 1.400 ;
        RECT 18.080 1.060 18.250 1.230 ;
        RECT 18.640 1.060 18.810 1.230 ;
        RECT 18.000 0.890 18.330 1.060 ;
        RECT 18.550 0.890 18.890 1.060 ;
        RECT 17.160 0.830 17.480 0.870 ;
        RECT 17.160 0.660 17.490 0.830 ;
        RECT 18.640 0.660 18.810 0.890 ;
        RECT 19.210 0.810 19.720 1.480 ;
        RECT 17.160 0.610 18.810 0.660 ;
        RECT 5.630 0.490 6.090 0.530 ;
        RECT 17.350 0.490 18.810 0.610 ;
        RECT 5.630 0.360 6.100 0.490 ;
        RECT 5.770 0.300 6.100 0.360 ;
        RECT 5.770 0.270 6.090 0.300 ;
      LAYER mcon ;
        RECT 5.620 9.970 5.790 10.140 ;
        RECT 3.950 9.560 4.120 9.730 ;
        RECT 4.680 9.530 4.850 9.700 ;
        RECT 5.620 9.420 5.790 9.590 ;
        RECT 6.800 8.810 6.970 8.980 ;
        RECT 3.950 8.020 4.120 8.190 ;
        RECT 10.820 8.840 10.990 9.010 ;
        RECT 4.680 8.050 4.850 8.220 ;
        RECT 5.620 8.160 5.790 8.330 ;
        RECT 5.620 7.610 5.790 7.780 ;
        RECT 6.790 7.610 6.960 7.780 ;
        RECT 6.790 6.950 6.960 7.120 ;
        RECT 5.620 6.730 5.790 6.900 ;
        RECT 10.810 7.550 10.980 7.720 ;
        RECT 10.810 6.910 10.980 7.080 ;
        RECT 3.950 6.320 4.120 6.490 ;
        RECT 4.680 6.290 4.850 6.460 ;
        RECT 5.620 6.180 5.790 6.350 ;
        RECT 17.220 5.380 17.390 5.550 ;
        RECT 3.950 4.770 4.120 4.940 ;
        RECT 4.680 4.800 4.850 4.970 ;
        RECT 5.620 4.910 5.790 5.080 ;
        RECT 19.380 4.970 19.550 5.140 ;
        RECT 17.370 4.700 17.540 4.870 ;
        RECT 5.620 4.360 5.790 4.530 ;
        RECT 18.120 4.400 18.290 4.570 ;
        RECT 17.370 4.100 17.540 4.270 ;
        RECT 19.380 3.830 19.550 4.000 ;
        RECT 17.220 3.420 17.390 3.590 ;
        RECT 17.220 2.610 17.390 2.780 ;
        RECT 19.380 2.200 19.550 2.370 ;
        RECT 17.370 1.930 17.540 2.100 ;
        RECT 18.120 1.630 18.290 1.800 ;
        RECT 5.780 1.270 5.950 1.440 ;
        RECT 17.370 1.330 17.540 1.500 ;
        RECT 19.380 1.060 19.550 1.230 ;
        RECT 17.220 0.650 17.390 0.820 ;
        RECT 5.830 0.310 6.000 0.480 ;
      LAYER met1 ;
        RECT 3.890 9.790 4.050 10.490 ;
        RECT 3.890 9.240 4.160 9.790 ;
        RECT 3.880 9.190 4.160 9.240 ;
        RECT 4.300 9.450 4.490 10.440 ;
        RECT 4.700 9.760 4.860 10.490 ;
        RECT 5.540 9.900 5.860 10.220 ;
        RECT 4.660 9.740 4.860 9.760 ;
        RECT 4.650 9.500 4.880 9.740 ;
        RECT 4.650 9.450 4.860 9.500 ;
        RECT 4.300 9.330 4.470 9.450 ;
        RECT 3.880 9.100 4.050 9.190 ;
        RECT 3.890 8.650 4.050 9.100 ;
        RECT 3.880 8.560 4.050 8.650 ;
        RECT 3.880 8.510 4.160 8.560 ;
        RECT 3.890 7.960 4.160 8.510 ;
        RECT 4.300 8.420 4.460 9.330 ;
        RECT 4.300 8.300 4.470 8.420 ;
        RECT 4.700 8.300 4.860 9.450 ;
        RECT 5.540 9.350 5.860 9.670 ;
        RECT 3.890 6.550 4.050 7.960 ;
        RECT 4.300 7.380 4.490 8.300 ;
        RECT 4.650 8.250 4.860 8.300 ;
        RECT 4.650 8.010 4.880 8.250 ;
        RECT 5.540 8.080 5.860 8.400 ;
        RECT 4.660 7.990 4.860 8.010 ;
        RECT 4.270 7.350 4.510 7.380 ;
        RECT 4.700 7.350 4.860 7.990 ;
        RECT 5.540 7.530 5.860 7.850 ;
        RECT 4.270 7.180 4.860 7.350 ;
        RECT 4.270 7.150 4.510 7.180 ;
        RECT 3.890 6.000 4.160 6.550 ;
        RECT 3.880 5.950 4.160 6.000 ;
        RECT 4.300 6.210 4.490 7.150 ;
        RECT 4.700 6.520 4.860 7.180 ;
        RECT 5.540 6.660 5.860 6.980 ;
        RECT 4.660 6.500 4.860 6.520 ;
        RECT 4.650 6.260 4.880 6.500 ;
        RECT 4.650 6.210 4.860 6.260 ;
        RECT 4.300 6.090 4.470 6.210 ;
        RECT 3.880 5.860 4.050 5.950 ;
        RECT 3.890 5.400 4.050 5.860 ;
        RECT 3.880 5.310 4.050 5.400 ;
        RECT 3.880 5.260 4.160 5.310 ;
        RECT 3.890 4.710 4.160 5.260 ;
        RECT 4.300 5.170 4.460 6.090 ;
        RECT 4.300 5.050 4.470 5.170 ;
        RECT 4.700 5.050 4.860 6.210 ;
        RECT 5.540 6.110 5.860 6.430 ;
        RECT 8.820 5.970 9.200 10.500 ;
        RECT 8.820 5.650 9.220 5.970 ;
        RECT 10.770 5.760 11.040 10.500 ;
        RECT 3.890 4.010 4.050 4.710 ;
        RECT 4.300 4.060 4.490 5.050 ;
        RECT 4.650 5.000 4.860 5.050 ;
        RECT 4.650 4.760 4.880 5.000 ;
        RECT 5.540 4.830 5.860 5.150 ;
        RECT 4.660 4.740 4.860 4.760 ;
        RECT 4.700 4.010 4.860 4.740 ;
        RECT 8.820 4.000 9.200 5.650 ;
        RECT 10.750 5.450 11.060 5.760 ;
        RECT 10.770 4.000 11.040 5.450 ;
        RECT 12.850 4.000 13.250 10.500 ;
        RECT 17.150 5.300 17.470 5.620 ;
        RECT 17.300 4.620 17.620 4.940 ;
        RECT 17.300 4.030 17.620 4.350 ;
        RECT 17.150 3.350 17.470 3.670 ;
        RECT 8.940 2.720 9.200 3.040 ;
        RECT 8.940 1.860 9.100 2.720 ;
        RECT 17.150 2.530 17.470 2.850 ;
        RECT 8.810 1.540 9.100 1.860 ;
        RECT 17.300 1.850 17.620 2.170 ;
        RECT 5.710 1.200 6.030 1.520 ;
        RECT 17.300 1.260 17.620 1.580 ;
        RECT 17.150 0.580 17.470 0.900 ;
        RECT 5.760 0.240 6.080 0.560 ;
        RECT 11.460 0.180 11.840 0.280 ;
      LAYER via ;
        RECT 5.570 9.930 5.830 10.190 ;
        RECT 5.570 9.380 5.830 9.640 ;
        RECT 5.570 8.110 5.830 8.370 ;
        RECT 5.570 7.560 5.830 7.820 ;
        RECT 5.570 6.690 5.830 6.950 ;
        RECT 5.570 6.140 5.830 6.400 ;
        RECT 8.960 5.680 9.220 5.940 ;
        RECT 5.570 4.860 5.830 5.120 ;
        RECT 10.770 5.470 11.040 5.730 ;
        RECT 8.940 4.630 9.200 4.890 ;
        RECT 17.180 5.330 17.440 5.590 ;
        RECT 17.330 4.650 17.590 4.910 ;
        RECT 17.330 4.060 17.590 4.320 ;
        RECT 17.180 3.380 17.440 3.640 ;
        RECT 8.940 2.750 9.200 3.010 ;
        RECT 17.180 2.560 17.440 2.820 ;
        RECT 17.330 1.880 17.590 2.140 ;
        RECT 8.810 1.570 9.070 1.830 ;
        RECT 5.740 1.230 6.000 1.490 ;
        RECT 17.330 1.290 17.590 1.550 ;
        RECT 17.180 0.610 17.440 0.870 ;
        RECT 5.790 0.270 6.050 0.530 ;
      LAYER met2 ;
        RECT 5.550 9.940 5.860 10.230 ;
        RECT 3.530 9.900 5.860 9.940 ;
        RECT 3.530 9.760 5.710 9.900 ;
        RECT 5.550 9.510 5.860 9.680 ;
        RECT 3.530 9.350 5.860 9.510 ;
        RECT 3.530 9.330 5.700 9.350 ;
        RECT 5.990 9.320 13.600 9.510 ;
        RECT 3.530 8.400 5.700 8.420 ;
        RECT 3.530 8.240 5.860 8.400 ;
        RECT 5.970 8.240 13.600 8.420 ;
        RECT 5.550 8.070 5.860 8.240 ;
        RECT 3.530 7.850 5.710 7.990 ;
        RECT 3.530 7.810 5.860 7.850 ;
        RECT 5.550 7.520 5.860 7.810 ;
        RECT 6.000 7.800 6.090 7.830 ;
        RECT 5.970 7.690 6.090 7.800 ;
        RECT 5.550 6.700 5.860 6.990 ;
        RECT 3.530 6.660 5.860 6.700 ;
        RECT 3.530 6.520 5.710 6.660 ;
        RECT 5.970 6.540 6.120 6.710 ;
        RECT 5.550 6.270 5.860 6.440 ;
        RECT 3.530 6.110 5.860 6.270 ;
        RECT 3.530 6.090 5.700 6.110 ;
        RECT 5.970 6.100 12.830 6.270 ;
        RECT 13.130 6.130 13.600 6.290 ;
        RECT 13.130 6.120 13.590 6.130 ;
        RECT 6.000 6.090 6.090 6.100 ;
        RECT 16.130 5.510 16.270 5.520 ;
        RECT 5.970 5.140 13.600 5.310 ;
        RECT 16.130 5.180 16.280 5.510 ;
        RECT 17.150 5.290 17.460 5.620 ;
        RECT 6.000 4.990 6.090 5.140 ;
        RECT 16.130 4.980 17.340 5.180 ;
        RECT 17.150 3.350 17.460 3.680 ;
        RECT 17.150 2.520 17.460 2.850 ;
        RECT 16.220 2.130 17.220 2.290 ;
        RECT 16.230 1.150 17.230 1.320 ;
        RECT 16.230 1.140 17.170 1.150 ;
        RECT 17.150 0.580 17.460 0.910 ;
  END
END sky130_hilas_WTA4Stage01

MACRO sky130_hilas_Trans4small
  CLASS CORE ;
  FOREIGN sky130_hilas_Trans4small ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.400 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN NFET_SOURCE1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 5.710 0.070 5.750 ;
        RECT 0.000 5.480 0.140 5.710 ;
    END
  END NFET_SOURCE1
  PIN NFET_GATE1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 5.070 0.160 5.240 ;
    END
  END NFET_GATE1
  PIN NFET_SOURCE2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 4.560 0.140 4.730 ;
    END
  END NFET_SOURCE2
  PIN NFET_GATE2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 4.150 0.170 4.320 ;
    END
  END NFET_GATE2
  PIN NFET_SOURCE3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 3.780 0.140 3.810 ;
        RECT 0.000 3.640 0.210 3.780 ;
    END
  END NFET_SOURCE3
  PIN NFET_GATE3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 3.230 0.160 3.400 ;
    END
  END NFET_GATE3
  PIN PFET_SOURCE1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 2.620 0.140 2.810 ;
    END
  END PFET_SOURCE1
  PIN PFET_GATE1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 2.200 0.140 2.390 ;
    END
  END PFET_GATE1
  PIN PFET_SOURCE2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 1.830 0.140 1.850 ;
        RECT 0.000 1.660 0.070 1.830 ;
    END
  END PFET_SOURCE2
  PIN PFET_GATE2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 1.410 0.140 1.430 ;
        RECT 0.000 1.240 0.070 1.410 ;
    END
  END PFET_GATE2
  PIN PFET_SOURCE3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 0.840 0.140 0.890 ;
        RECT 0.000 0.700 0.070 0.840 ;
    END
  END PFET_SOURCE3
  PIN PFET_GATE3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 0.450 0.140 0.470 ;
        RECT 0.000 0.280 0.150 0.450 ;
    END
  END PFET_GATE3
  PIN WELL
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 1.280 0.680 3.310 3.650 ;
        RECT 2.100 0.630 2.640 0.680 ;
        RECT 1.920 0.180 2.640 0.630 ;
        RECT 0.070 0.000 2.640 0.180 ;
      LAYER met2 ;
        RECT 1.850 1.790 2.170 1.930 ;
        RECT 1.850 1.650 2.800 1.790 ;
        RECT 1.760 1.590 2.800 1.650 ;
        RECT 1.760 1.320 2.070 1.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.850 1.890 2.170 1.930 ;
        RECT 1.620 1.660 2.170 1.890 ;
        RECT 1.850 1.640 2.170 1.660 ;
        RECT 1.760 1.610 2.170 1.640 ;
        RECT 1.760 1.320 2.080 1.610 ;
        RECT 2.180 1.270 2.400 5.880 ;
        RECT 2.160 1.200 2.400 1.270 ;
        RECT 2.160 1.100 2.500 1.200 ;
        RECT 2.180 0.970 2.500 1.100 ;
        RECT 2.180 0.000 2.400 0.970 ;
      LAYER via ;
        RECT 1.880 1.640 2.140 1.900 ;
        RECT 1.790 1.350 2.050 1.610 ;
    END
  END WELL
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 1.850 5.080 2.160 5.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.850 5.080 2.170 5.400 ;
        RECT 2.580 5.330 2.800 5.880 ;
        RECT 2.580 5.040 2.900 5.330 ;
        RECT 2.580 0.000 2.800 5.040 ;
      LAYER via ;
        RECT 1.880 5.110 2.140 5.370 ;
    END
  END VGND
  PIN PFET_DRAIN3
    USE ANALOG ;
    ANTENNAGATEAREA 0.163800 ;
    PORT
      LAYER met2 ;
        RECT 1.850 0.830 2.170 0.940 ;
        RECT 1.850 0.630 2.800 0.830 ;
        RECT 1.850 0.620 2.170 0.630 ;
    END
  END PFET_DRAIN3
  PIN PFET_DRAIN1
    USE ANALOG ;
    ANTENNAGATEAREA 0.163800 ;
    ANTENNADIFFAREA 0.117600 ;
    PORT
      LAYER met2 ;
        RECT 1.850 2.750 2.170 2.920 ;
        RECT 1.850 2.640 2.800 2.750 ;
        RECT 1.760 2.550 2.800 2.640 ;
        RECT 1.760 2.310 2.070 2.550 ;
    END
  END PFET_DRAIN1
  PIN NFET_DRAIN3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.980 3.650 2.800 3.820 ;
    END
  END NFET_DRAIN3
  PIN NFET_DRAIN2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.980 4.570 2.800 4.740 ;
    END
  END NFET_DRAIN2
  PIN NFET_DRAIN1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.980 5.490 2.800 5.660 ;
    END
  END NFET_DRAIN1
  OBS
      LAYER li1 ;
        RECT 2.020 5.920 2.220 6.050 ;
        RECT 2.610 5.920 2.810 6.050 ;
        RECT 1.470 5.610 1.800 5.780 ;
        RECT 0.310 5.410 0.630 5.450 ;
        RECT 0.310 5.220 0.640 5.410 ;
        RECT 1.860 5.330 2.180 5.370 ;
        RECT 2.950 5.340 3.270 5.380 ;
        RECT 1.860 5.260 2.190 5.330 ;
        RECT 2.200 5.260 2.370 5.310 ;
        RECT 2.690 5.260 2.880 5.300 ;
        RECT 1.860 5.230 2.370 5.260 ;
        RECT 2.620 5.230 2.880 5.260 ;
        RECT 0.310 5.190 0.630 5.220 ;
        RECT 0.330 5.120 0.540 5.190 ;
        RECT 1.860 5.110 2.880 5.230 ;
        RECT 2.950 5.150 3.280 5.340 ;
        RECT 2.950 5.120 3.270 5.150 ;
        RECT 2.030 5.070 2.880 5.110 ;
        RECT 2.030 4.980 2.820 5.070 ;
        RECT 2.030 4.930 2.380 4.980 ;
        RECT 2.620 4.930 2.820 4.980 ;
        RECT 2.200 4.920 2.380 4.930 ;
        RECT 1.480 4.620 1.810 4.790 ;
        RECT 0.290 4.490 0.610 4.530 ;
        RECT 0.290 4.300 0.620 4.490 ;
        RECT 1.860 4.340 2.180 4.380 ;
        RECT 2.950 4.350 3.270 4.390 ;
        RECT 0.290 4.270 0.610 4.300 ;
        RECT 1.860 4.270 2.190 4.340 ;
        RECT 1.860 4.120 2.230 4.270 ;
        RECT 2.030 3.940 2.230 4.120 ;
        RECT 2.620 3.940 2.820 4.270 ;
        RECT 2.950 4.160 3.280 4.350 ;
        RECT 2.950 4.130 3.270 4.160 ;
        RECT 1.480 3.630 1.810 3.800 ;
        RECT 1.770 3.550 2.090 3.590 ;
        RECT 0.270 3.500 0.590 3.540 ;
        RECT 0.270 3.310 0.600 3.500 ;
        RECT 1.770 3.380 2.100 3.550 ;
        RECT 3.070 3.450 3.390 3.490 ;
        RECT 1.770 3.330 2.250 3.380 ;
        RECT 0.270 3.280 0.590 3.310 ;
        RECT 1.940 3.200 2.250 3.330 ;
        RECT 1.920 3.180 2.250 3.200 ;
        RECT 2.080 3.050 2.250 3.180 ;
        RECT 2.760 3.050 2.930 3.380 ;
        RECT 3.070 3.260 3.400 3.450 ;
        RECT 3.070 3.230 3.390 3.260 ;
        RECT 1.700 2.850 2.130 2.870 ;
        RECT 1.680 2.680 2.130 2.850 ;
        RECT 1.700 2.660 2.130 2.680 ;
        RECT 1.770 2.560 2.090 2.600 ;
        RECT 1.770 2.390 2.100 2.560 ;
        RECT 3.070 2.460 3.390 2.500 ;
        RECT 1.770 2.340 2.250 2.390 ;
        RECT 1.940 2.210 2.250 2.340 ;
        RECT 1.920 2.190 2.250 2.210 ;
        RECT 2.080 2.060 2.250 2.190 ;
        RECT 2.760 2.060 2.930 2.390 ;
        RECT 3.070 2.270 3.400 2.460 ;
        RECT 3.070 2.240 3.390 2.270 ;
        RECT 1.700 1.860 2.130 1.880 ;
        RECT 1.680 1.690 2.130 1.860 ;
        RECT 1.700 1.670 2.130 1.690 ;
        RECT 1.770 1.570 2.090 1.610 ;
        RECT 1.770 1.400 2.100 1.570 ;
        RECT 3.070 1.470 3.390 1.510 ;
        RECT 1.770 1.350 2.250 1.400 ;
        RECT 1.940 1.270 2.250 1.350 ;
        RECT 1.940 1.220 2.410 1.270 ;
        RECT 1.920 1.200 2.410 1.220 ;
        RECT 2.080 1.180 2.410 1.200 ;
        RECT 2.080 1.070 2.470 1.180 ;
        RECT 2.760 1.070 2.930 1.400 ;
        RECT 3.070 1.280 3.400 1.470 ;
        RECT 3.070 1.250 3.390 1.280 ;
        RECT 2.240 0.990 2.470 1.070 ;
        RECT 1.700 0.870 2.130 0.890 ;
        RECT 1.680 0.700 2.130 0.870 ;
        RECT 1.700 0.680 2.130 0.700 ;
      LAYER mcon ;
        RECT 0.370 5.230 0.540 5.400 ;
        RECT 1.920 5.150 2.090 5.320 ;
        RECT 2.700 5.100 2.870 5.270 ;
        RECT 3.010 5.160 3.180 5.330 ;
        RECT 0.350 4.310 0.520 4.480 ;
        RECT 1.920 4.160 2.090 4.330 ;
        RECT 3.010 4.170 3.180 4.340 ;
        RECT 0.330 3.320 0.500 3.490 ;
        RECT 1.830 3.370 2.000 3.540 ;
        RECT 3.130 3.270 3.300 3.440 ;
        RECT 1.830 2.380 2.000 2.550 ;
        RECT 3.130 2.280 3.300 2.450 ;
        RECT 1.830 1.390 2.000 1.560 ;
        RECT 2.270 1.000 2.440 1.170 ;
        RECT 3.130 1.290 3.300 1.460 ;
      LAYER met1 ;
        RECT 0.300 5.160 0.620 5.480 ;
        RECT 2.940 5.090 3.260 5.410 ;
        RECT 0.280 4.240 0.600 4.560 ;
        RECT 1.850 4.090 2.170 4.410 ;
        RECT 2.940 4.100 3.260 4.420 ;
        RECT 0.260 3.250 0.580 3.570 ;
        RECT 1.760 3.300 2.080 3.620 ;
        RECT 3.060 3.200 3.380 3.520 ;
        RECT 1.850 2.880 2.170 2.920 ;
        RECT 1.620 2.650 2.170 2.880 ;
        RECT 1.850 2.630 2.170 2.650 ;
        RECT 1.760 2.600 2.170 2.630 ;
        RECT 1.760 2.310 2.080 2.600 ;
        RECT 3.060 2.210 3.380 2.530 ;
        RECT 3.060 1.220 3.380 1.540 ;
        RECT 1.850 0.900 2.170 0.940 ;
        RECT 1.620 0.670 2.170 0.900 ;
        RECT 1.850 0.620 2.170 0.670 ;
      LAYER via ;
        RECT 0.330 5.190 0.590 5.450 ;
        RECT 2.970 5.120 3.230 5.380 ;
        RECT 0.310 4.270 0.570 4.530 ;
        RECT 1.880 4.120 2.140 4.380 ;
        RECT 2.970 4.130 3.230 4.390 ;
        RECT 0.290 3.280 0.550 3.540 ;
        RECT 1.790 3.330 2.050 3.590 ;
        RECT 3.090 3.230 3.350 3.490 ;
        RECT 1.880 2.630 2.140 2.890 ;
        RECT 1.790 2.340 2.050 2.600 ;
        RECT 3.090 2.240 3.350 2.500 ;
        RECT 3.090 1.250 3.350 1.510 ;
        RECT 1.880 0.650 2.140 0.910 ;
      LAYER met2 ;
        RECT 1.170 5.990 1.770 6.050 ;
        RECT 3.030 6.000 3.250 6.050 ;
        RECT 0.300 5.160 0.610 5.490 ;
        RECT 2.940 5.180 3.250 5.420 ;
        RECT 1.180 5.000 1.780 5.170 ;
        RECT 2.940 5.090 3.260 5.180 ;
        RECT 3.040 5.010 3.260 5.090 ;
        RECT 0.280 4.240 0.590 4.570 ;
        RECT 1.180 4.010 1.780 4.180 ;
        RECT 1.850 4.090 2.160 4.420 ;
        RECT 2.940 4.190 3.250 4.430 ;
        RECT 2.940 4.100 3.260 4.190 ;
        RECT 3.040 4.020 3.260 4.100 ;
        RECT 0.260 3.250 0.570 3.580 ;
        RECT 1.280 3.180 1.650 3.370 ;
        RECT 1.760 3.300 2.070 3.630 ;
        RECT 3.060 3.200 3.370 3.530 ;
        RECT 1.280 2.760 1.660 2.950 ;
        RECT 1.280 2.190 1.650 2.380 ;
        RECT 3.060 2.210 3.370 2.540 ;
        RECT 1.280 1.770 1.660 1.960 ;
        RECT 1.280 1.200 1.650 1.390 ;
        RECT 3.060 1.220 3.370 1.550 ;
        RECT 1.280 0.780 1.660 0.970 ;
  END
END sky130_hilas_Trans4small

MACRO sky130_hilas_FGBiasWeakGate2x1cell
  CLASS CORE ;
  FOREIGN sky130_hilas_FGBiasWeakGate2x1cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 10.100 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 9.050 5.600 9.360 5.610 ;
        RECT 0.000 5.420 11.530 5.600 ;
        RECT 9.050 5.280 9.360 5.420 ;
    END
  END DRAIN1
  PIN VIN11
    PORT
      LAYER met2 ;
        RECT 1.940 5.010 2.250 5.060 ;
        RECT 1.790 5.000 2.250 5.010 ;
        RECT 0.000 4.820 2.250 5.000 ;
        RECT 1.940 4.730 2.250 4.820 ;
    END
  END VIN11
  PIN ROW1
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 9.200 4.580 9.510 4.650 ;
        RECT 9.200 4.570 11.530 4.580 ;
        RECT 0.000 4.360 11.530 4.570 ;
        RECT 0.000 4.350 10.220 4.360 ;
        RECT 9.200 4.320 9.510 4.350 ;
    END
  END ROW1
  PIN ROW2
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 9.200 1.820 9.510 1.890 ;
        RECT 0.000 1.610 11.530 1.820 ;
        RECT 0.000 1.600 10.220 1.610 ;
        RECT 9.200 1.560 9.510 1.600 ;
    END
  END ROW2
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 8.220 0.000 11.530 6.150 ;
      LAYER met1 ;
        RECT 11.010 5.450 11.290 6.100 ;
        RECT 10.900 4.850 11.290 5.450 ;
        RECT 11.010 1.300 11.290 4.850 ;
        RECT 10.900 0.700 11.290 1.300 ;
        RECT 11.010 0.050 11.290 0.700 ;
    END
  END VINJ
  PIN COLSEL1
    USE ANALOG ;
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT 10.570 4.640 10.760 6.100 ;
        RECT 10.570 4.610 10.790 4.640 ;
        RECT 10.550 4.340 10.800 4.610 ;
        RECT 10.560 4.330 10.800 4.340 ;
        RECT 10.560 4.090 10.790 4.330 ;
        RECT 10.600 2.060 10.760 4.090 ;
        RECT 10.560 1.820 10.790 2.060 ;
        RECT 10.560 1.810 10.800 1.820 ;
        RECT 10.550 1.540 10.800 1.810 ;
        RECT 10.570 1.510 10.790 1.540 ;
        RECT 10.570 0.050 10.760 1.510 ;
    END
  END COLSEL1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2.830 5.130 3.060 6.100 ;
        RECT 2.830 4.880 3.070 5.130 ;
        RECT 2.830 0.050 3.060 4.880 ;
    END
  END VGND
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT 3.770 3.710 6.490 5.360 ;
        RECT 3.770 3.670 6.480 3.710 ;
        RECT 3.770 2.340 6.480 2.380 ;
        RECT 3.770 0.690 6.490 2.340 ;
      LAYER met1 ;
        RECT 4.050 4.890 4.280 6.100 ;
        RECT 4.050 4.100 4.310 4.890 ;
        RECT 4.050 1.950 4.280 4.100 ;
        RECT 4.050 1.160 4.310 1.950 ;
        RECT 4.050 0.050 4.280 1.160 ;
    END
  END GATE1
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 1.808400 ;
    PORT
      LAYER nwell ;
        RECT 0.020 1.780 1.750 5.350 ;
        RECT 0.590 1.450 1.150 1.780 ;
      LAYER met1 ;
        RECT 0.350 0.060 0.770 6.100 ;
    END
  END VTUN
  PIN DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 9.050 0.730 9.360 0.870 ;
        RECT 9.050 0.720 11.530 0.730 ;
        RECT 0.000 0.570 11.530 0.720 ;
        RECT 9.050 0.550 11.530 0.570 ;
        RECT 9.050 0.540 9.360 0.550 ;
    END
  END DRAIN2
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 1.290 2.220 1.370 ;
        RECT 0.000 1.080 2.220 1.290 ;
        RECT 1.910 1.040 2.220 1.080 ;
    END
  END VIN12
  PIN COMMONSOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 1.030400 ;
    PORT
      LAYER met2 ;
        RECT 0.000 3.380 10.460 3.600 ;
        RECT 10.140 3.240 10.460 3.380 ;
        RECT 10.180 2.900 10.440 3.240 ;
        RECT 10.140 2.640 10.460 2.900 ;
    END
  END COMMONSOURCE
  OBS
      LAYER nwell ;
        RECT 14.520 8.200 16.250 10.100 ;
        RECT 14.520 4.060 16.250 5.960 ;
      LAYER li1 ;
        RECT 1.870 5.090 6.930 5.920 ;
        RECT 9.120 5.520 9.650 5.690 ;
        RECT 10.930 5.420 11.130 5.770 ;
        RECT 10.930 5.390 11.140 5.420 ;
        RECT 1.940 5.010 2.420 5.090 ;
        RECT 1.950 4.760 2.420 5.010 ;
        RECT 0.440 3.960 0.990 4.390 ;
        RECT 4.070 4.150 4.300 4.840 ;
        RECT 9.370 4.610 9.540 5.130 ;
        RECT 9.210 4.350 9.540 4.610 ;
        RECT 3.040 3.130 3.230 3.530 ;
        RECT 9.370 3.440 9.540 4.350 ;
        RECT 10.200 3.530 10.370 5.140 ;
        RECT 10.920 4.810 11.140 5.390 ;
        RECT 10.930 4.800 11.140 4.810 ;
        RECT 10.570 4.630 10.760 4.640 ;
        RECT 10.570 4.340 10.770 4.630 ;
        RECT 10.560 4.010 10.850 4.340 ;
        RECT 10.200 3.340 10.380 3.530 ;
        RECT 2.850 3.120 3.230 3.130 ;
        RECT 2.850 2.940 6.590 3.120 ;
        RECT 2.850 2.900 3.230 2.940 ;
        RECT 0.440 2.230 0.990 2.660 ;
        RECT 3.040 2.520 3.230 2.900 ;
        RECT 1.920 1.080 2.260 1.330 ;
        RECT 4.070 1.210 4.300 1.940 ;
        RECT 9.370 1.850 9.540 2.710 ;
        RECT 9.210 1.590 9.540 1.850 ;
        RECT 1.910 1.000 2.260 1.080 ;
        RECT 9.370 1.020 9.540 1.590 ;
        RECT 10.200 2.620 10.380 2.810 ;
        RECT 10.200 1.010 10.370 2.620 ;
        RECT 10.560 1.810 10.850 2.140 ;
        RECT 10.570 1.520 10.770 1.810 ;
        RECT 10.570 1.510 10.760 1.520 ;
        RECT 10.930 1.340 11.140 1.350 ;
        RECT 1.910 0.150 6.960 1.000 ;
        RECT 10.920 0.760 11.140 1.340 ;
        RECT 10.930 0.730 11.140 0.760 ;
        RECT 9.120 0.460 9.650 0.630 ;
        RECT 10.930 0.380 11.130 0.730 ;
      LAYER mcon ;
        RECT 10.940 5.220 11.110 5.390 ;
        RECT 2.010 4.800 2.180 4.970 ;
        RECT 4.100 4.640 4.270 4.810 ;
        RECT 0.440 4.040 0.710 4.310 ;
        RECT 4.100 4.190 4.270 4.360 ;
        RECT 9.270 4.390 9.440 4.560 ;
        RECT 10.580 4.380 10.760 4.570 ;
        RECT 2.860 2.930 3.030 3.100 ;
        RECT 0.440 2.310 0.710 2.580 ;
        RECT 4.100 1.690 4.270 1.860 ;
        RECT 9.270 1.630 9.440 1.800 ;
        RECT 1.980 1.110 2.150 1.280 ;
        RECT 4.100 1.240 4.270 1.410 ;
        RECT 10.580 1.580 10.760 1.770 ;
        RECT 10.940 0.760 11.110 0.930 ;
      LAYER met1 ;
        RECT 9.050 5.280 9.360 5.720 ;
        RECT 1.940 4.730 2.260 5.050 ;
        RECT 9.200 4.320 9.520 4.640 ;
        RECT 10.170 3.530 10.410 3.660 ;
        RECT 10.170 3.210 10.430 3.530 ;
        RECT 10.170 2.610 10.430 2.930 ;
        RECT 10.170 2.490 10.410 2.610 ;
        RECT 9.200 1.560 9.520 1.880 ;
        RECT 1.910 1.040 2.230 1.360 ;
        RECT 9.050 0.430 9.360 0.870 ;
      LAYER via ;
        RECT 9.080 5.310 9.340 5.570 ;
        RECT 1.970 4.760 2.230 5.020 ;
        RECT 9.230 4.350 9.490 4.610 ;
        RECT 10.170 3.240 10.430 3.500 ;
        RECT 10.170 2.640 10.430 2.900 ;
        RECT 9.230 1.590 9.490 1.850 ;
        RECT 1.940 1.070 2.200 1.330 ;
        RECT 9.080 0.580 9.340 0.840 ;
  END
END sky130_hilas_FGBiasWeakGate2x1cell

MACRO sky130_hilas_swc4x2cell
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x2cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 32.460 BY 10.490 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 20.620 0.000 21.000 6.500 ;
    END
  END GATE2
  PIN VTUN
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 15.490 6.130 15.890 6.500 ;
        RECT 16.570 6.130 16.970 6.500 ;
        RECT 15.490 5.910 16.970 6.130 ;
        RECT 15.490 0.000 15.890 5.910 ;
        RECT 16.570 0.000 16.970 5.910 ;
    END
  END VTUN
  PIN GATE1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 11.460 0.000 11.840 6.500 ;
    END
  END GATE1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 6.170 0.000 8.730 6.500 ;
        RECT 23.730 0.000 26.290 6.500 ;
      LAYER met2 ;
        RECT 6.370 6.220 26.110 6.400 ;
        RECT 6.370 6.080 6.790 6.220 ;
        RECT 8.190 5.940 8.500 6.220 ;
        RECT 6.170 5.900 8.500 5.940 ;
        RECT 23.960 5.940 24.270 6.220 ;
        RECT 25.770 6.090 26.110 6.220 ;
        RECT 23.960 5.900 26.290 5.940 ;
        RECT 6.170 5.760 8.350 5.900 ;
        RECT 24.110 5.760 26.290 5.900 ;
    END
  END VINJ
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 25.770 6.380 25.930 6.490 ;
        RECT 25.770 6.100 26.100 6.380 ;
        RECT 25.770 5.790 25.930 6.100 ;
        RECT 25.660 5.240 25.930 5.790 ;
        RECT 25.660 5.190 25.940 5.240 ;
        RECT 25.770 5.100 25.940 5.190 ;
        RECT 25.770 4.630 25.930 5.100 ;
        RECT 25.770 4.540 25.940 4.630 ;
        RECT 25.660 4.490 25.940 4.540 ;
        RECT 25.660 3.940 25.930 4.490 ;
        RECT 25.770 2.550 25.930 3.940 ;
        RECT 25.660 2.000 25.930 2.550 ;
        RECT 25.660 1.950 25.940 2.000 ;
        RECT 25.770 1.860 25.940 1.950 ;
        RECT 25.770 1.400 25.930 1.860 ;
        RECT 25.770 1.310 25.940 1.400 ;
        RECT 25.660 1.260 25.940 1.310 ;
        RECT 25.660 0.710 25.930 1.260 ;
        RECT 25.770 0.010 25.930 0.710 ;
      LAYER via ;
        RECT 25.810 6.110 26.070 6.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.530 6.370 6.690 6.490 ;
        RECT 6.380 6.230 6.690 6.370 ;
        RECT 6.370 6.080 6.690 6.230 ;
        RECT 6.530 5.790 6.690 6.080 ;
        RECT 6.530 5.240 6.800 5.790 ;
        RECT 6.520 5.190 6.800 5.240 ;
        RECT 6.520 5.100 6.690 5.190 ;
        RECT 6.530 4.630 6.690 5.100 ;
        RECT 6.520 4.540 6.690 4.630 ;
        RECT 6.520 4.490 6.800 4.540 ;
        RECT 6.530 3.940 6.800 4.490 ;
        RECT 6.530 2.550 6.690 3.940 ;
        RECT 6.530 2.000 6.800 2.550 ;
        RECT 6.520 1.950 6.800 2.000 ;
        RECT 6.520 1.860 6.690 1.950 ;
        RECT 6.530 1.400 6.690 1.860 ;
        RECT 6.520 1.310 6.690 1.400 ;
        RECT 6.520 1.260 6.800 1.310 ;
        RECT 6.530 0.710 6.800 1.260 ;
        RECT 6.530 0.010 6.690 0.710 ;
      LAYER via ;
        RECT 6.410 6.100 6.670 6.360 ;
    END
  END VINJ
  PIN GATESELECT1
    USE ANALOG ;
    ANTENNAGATEAREA 0.720000 ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met1 ;
        RECT 6.940 5.450 7.130 6.440 ;
        RECT 7.340 5.760 7.500 6.490 ;
        RECT 7.300 5.740 7.500 5.760 ;
        RECT 7.290 5.500 7.520 5.740 ;
        RECT 7.290 5.450 7.500 5.500 ;
        RECT 6.940 5.330 7.110 5.450 ;
        RECT 6.940 4.400 7.100 5.330 ;
        RECT 6.940 4.280 7.110 4.400 ;
        RECT 7.340 4.280 7.500 5.450 ;
        RECT 6.940 3.360 7.130 4.280 ;
        RECT 7.290 4.230 7.500 4.280 ;
        RECT 7.290 3.990 7.520 4.230 ;
        RECT 7.300 3.970 7.500 3.990 ;
        RECT 6.910 3.340 7.150 3.360 ;
        RECT 7.340 3.340 7.500 3.970 ;
        RECT 6.910 3.150 7.500 3.340 ;
        RECT 6.910 3.130 7.150 3.150 ;
        RECT 6.940 2.210 7.130 3.130 ;
        RECT 7.340 2.520 7.500 3.150 ;
        RECT 7.300 2.500 7.500 2.520 ;
        RECT 7.290 2.260 7.520 2.500 ;
        RECT 7.290 2.210 7.500 2.260 ;
        RECT 6.940 2.090 7.110 2.210 ;
        RECT 6.940 1.170 7.100 2.090 ;
        RECT 6.940 1.050 7.110 1.170 ;
        RECT 7.340 1.050 7.500 2.210 ;
        RECT 6.940 0.060 7.130 1.050 ;
        RECT 7.290 1.000 7.500 1.050 ;
        RECT 7.290 0.760 7.520 1.000 ;
        RECT 7.300 0.740 7.500 0.760 ;
        RECT 7.340 0.010 7.500 0.740 ;
    END
  END GATESELECT1
  PIN GATESELECT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.720000 ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met1 ;
        RECT 24.960 5.760 25.120 6.490 ;
        RECT 24.960 5.740 25.160 5.760 ;
        RECT 24.940 5.500 25.170 5.740 ;
        RECT 24.960 5.450 25.170 5.500 ;
        RECT 25.330 5.450 25.520 6.440 ;
        RECT 24.960 4.280 25.120 5.450 ;
        RECT 25.350 5.330 25.520 5.450 ;
        RECT 25.360 4.400 25.520 5.330 ;
        RECT 25.350 4.280 25.520 4.400 ;
        RECT 24.960 4.230 25.170 4.280 ;
        RECT 24.940 3.990 25.170 4.230 ;
        RECT 24.960 3.970 25.160 3.990 ;
        RECT 24.960 3.340 25.120 3.970 ;
        RECT 25.330 3.360 25.520 4.280 ;
        RECT 25.310 3.340 25.550 3.360 ;
        RECT 24.960 3.150 25.550 3.340 ;
        RECT 24.960 2.520 25.120 3.150 ;
        RECT 25.310 3.130 25.550 3.150 ;
        RECT 24.960 2.500 25.160 2.520 ;
        RECT 24.940 2.260 25.170 2.500 ;
        RECT 24.960 2.210 25.170 2.260 ;
        RECT 25.330 2.210 25.520 3.130 ;
        RECT 24.960 1.050 25.120 2.210 ;
        RECT 25.350 2.090 25.520 2.210 ;
        RECT 25.360 1.170 25.520 2.090 ;
        RECT 25.350 1.050 25.520 1.170 ;
        RECT 24.960 1.000 25.170 1.050 ;
        RECT 24.940 0.760 25.170 1.000 ;
        RECT 24.960 0.740 25.160 0.760 ;
        RECT 24.960 0.010 25.120 0.740 ;
        RECT 25.330 0.060 25.520 1.050 ;
    END
  END GATESELECT2
  PIN ROW1
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 8.190 5.510 8.500 5.680 ;
        RECT 6.170 5.350 8.500 5.510 ;
        RECT 6.170 5.330 8.340 5.350 ;
    END
    PORT
      LAYER met2 ;
        RECT 23.960 5.510 24.270 5.680 ;
        RECT 23.960 5.350 26.290 5.510 ;
        RECT 24.120 5.330 26.290 5.350 ;
    END
  END ROW1
  PIN ROW2
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 6.170 4.380 8.340 4.400 ;
        RECT 6.170 4.220 8.500 4.380 ;
        RECT 8.190 4.050 8.500 4.220 ;
    END
    PORT
      LAYER met2 ;
        RECT 24.120 4.380 26.290 4.400 ;
        RECT 23.960 4.220 26.290 4.380 ;
        RECT 23.960 4.050 24.270 4.220 ;
    END
  END ROW2
  PIN DRAIN2
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 6.170 3.830 8.350 3.970 ;
        RECT 6.170 3.790 8.500 3.830 ;
        RECT 8.190 3.500 8.500 3.790 ;
    END
    PORT
      LAYER met2 ;
        RECT 24.110 3.830 26.290 3.970 ;
        RECT 23.960 3.790 26.290 3.830 ;
        RECT 23.960 3.500 24.270 3.790 ;
    END
  END DRAIN2
  PIN DRAIN3
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 8.190 2.700 8.500 2.990 ;
        RECT 6.170 2.660 8.500 2.700 ;
        RECT 6.170 2.520 8.350 2.660 ;
    END
    PORT
      LAYER met2 ;
        RECT 23.960 2.700 24.270 2.990 ;
        RECT 23.960 2.660 26.290 2.700 ;
        RECT 24.110 2.520 26.290 2.660 ;
    END
  END DRAIN3
  PIN ROW3
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 8.190 2.270 8.500 2.440 ;
        RECT 6.170 2.110 8.500 2.270 ;
        RECT 6.170 2.090 8.340 2.110 ;
    END
    PORT
      LAYER met2 ;
        RECT 23.960 2.270 24.270 2.440 ;
        RECT 23.960 2.110 26.290 2.270 ;
        RECT 24.120 2.090 26.290 2.110 ;
    END
  END ROW3
  PIN ROW4
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 6.170 1.150 8.340 1.170 ;
        RECT 6.170 0.990 8.500 1.150 ;
        RECT 8.190 0.820 8.500 0.990 ;
    END
    PORT
      LAYER met2 ;
        RECT 24.120 1.150 26.290 1.170 ;
        RECT 23.960 0.990 26.290 1.150 ;
        RECT 23.960 0.820 24.270 0.990 ;
    END
  END ROW4
  PIN DRAIN4
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 6.170 0.600 8.350 0.740 ;
        RECT 6.170 0.560 8.500 0.600 ;
        RECT 8.190 0.270 8.500 0.560 ;
    END
    PORT
      LAYER met2 ;
        RECT 24.110 0.600 26.290 0.740 ;
        RECT 23.960 0.560 26.290 0.600 ;
        RECT 23.960 0.270 24.270 0.560 ;
    END
  END DRAIN4
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 9.240 1.780 9.560 1.840 ;
        RECT 13.170 1.780 13.490 1.790 ;
        RECT 18.970 1.780 19.290 1.790 ;
        RECT 22.900 1.780 23.220 1.840 ;
        RECT 9.240 1.600 23.220 1.780 ;
        RECT 9.240 1.550 9.560 1.600 ;
        RECT 13.170 1.530 13.490 1.600 ;
        RECT 18.970 1.530 19.290 1.600 ;
        RECT 22.900 1.550 23.220 1.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 9.280 5.110 9.520 6.500 ;
        RECT 9.270 4.450 9.540 5.110 ;
        RECT 9.280 1.860 9.520 4.450 ;
        RECT 9.270 1.540 9.530 1.860 ;
        RECT 9.280 0.000 9.520 1.540 ;
      LAYER via ;
        RECT 9.270 1.570 9.530 1.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.210 5.090 13.450 6.500 ;
        RECT 13.200 4.430 13.460 5.090 ;
        RECT 13.210 1.820 13.450 4.430 ;
        RECT 13.200 1.500 13.460 1.820 ;
        RECT 13.210 0.000 13.450 1.500 ;
      LAYER via ;
        RECT 13.200 1.530 13.460 1.790 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.010 5.090 19.250 6.500 ;
        RECT 19.000 4.430 19.260 5.090 ;
        RECT 19.010 1.820 19.250 4.430 ;
        RECT 19.000 1.500 19.260 1.820 ;
        RECT 19.010 0.000 19.250 1.500 ;
      LAYER via ;
        RECT 19.000 1.530 19.260 1.790 ;
    END
    PORT
      LAYER met1 ;
        RECT 22.940 5.110 23.180 6.500 ;
        RECT 22.920 4.450 23.190 5.110 ;
        RECT 22.940 1.860 23.180 4.450 ;
        RECT 22.930 1.540 23.190 1.860 ;
        RECT 22.940 0.000 23.180 1.540 ;
      LAYER via ;
        RECT 22.930 1.570 23.190 1.830 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 0.000 8.820 1.730 10.490 ;
        RECT 30.730 8.820 32.460 10.490 ;
        RECT 0.000 6.980 1.760 8.820 ;
        RECT 30.700 6.980 32.460 8.820 ;
        RECT 0.000 4.000 1.730 6.980 ;
        RECT 10.260 0.000 12.490 6.490 ;
        RECT 16.170 5.160 16.290 5.340 ;
        RECT 15.080 4.810 15.670 4.920 ;
        RECT 16.790 4.810 17.380 4.920 ;
        RECT 15.080 1.530 15.670 1.720 ;
        RECT 16.790 1.530 17.380 1.720 ;
        RECT 19.970 0.000 22.200 6.490 ;
        RECT 30.730 4.000 32.460 6.980 ;
      LAYER li1 ;
        RECT 0.790 7.430 1.340 7.860 ;
        RECT 31.120 7.430 31.670 7.860 ;
        RECT 8.170 6.150 8.490 6.190 ;
        RECT 6.570 5.760 6.770 6.110 ;
        RECT 8.160 6.030 8.490 6.150 ;
        RECT 8.050 5.930 8.490 6.030 ;
        RECT 23.970 6.150 24.290 6.190 ;
        RECT 23.970 6.030 24.300 6.150 ;
        RECT 23.970 5.930 24.410 6.030 ;
        RECT 8.050 5.860 8.390 5.930 ;
        RECT 24.070 5.860 24.410 5.930 ;
        RECT 6.560 5.730 6.770 5.760 ;
        RECT 25.690 5.760 25.890 6.110 ;
        RECT 6.560 5.140 6.780 5.730 ;
        RECT 7.300 5.140 7.500 5.740 ;
        RECT 8.170 5.600 8.490 5.640 ;
        RECT 8.160 5.410 8.490 5.600 ;
        RECT 8.050 5.380 8.490 5.410 ;
        RECT 23.970 5.600 24.290 5.640 ;
        RECT 23.970 5.410 24.300 5.600 ;
        RECT 23.970 5.380 24.410 5.410 ;
        RECT 8.050 5.240 8.390 5.380 ;
        RECT 24.070 5.240 24.410 5.380 ;
        RECT 24.960 5.140 25.160 5.740 ;
        RECT 25.690 5.730 25.900 5.760 ;
        RECT 25.680 5.140 25.900 5.730 ;
        RECT 6.560 4.000 6.780 4.590 ;
        RECT 6.560 3.970 6.770 4.000 ;
        RECT 7.300 3.990 7.500 4.590 ;
        RECT 9.310 4.510 9.480 5.040 ;
        RECT 13.250 4.520 13.420 5.050 ;
        RECT 19.040 4.520 19.210 5.050 ;
        RECT 22.980 4.510 23.150 5.040 ;
        RECT 8.050 4.350 8.390 4.490 ;
        RECT 24.070 4.350 24.410 4.490 ;
        RECT 8.050 4.320 8.490 4.350 ;
        RECT 8.160 4.130 8.490 4.320 ;
        RECT 8.170 4.090 8.490 4.130 ;
        RECT 23.970 4.320 24.410 4.350 ;
        RECT 23.970 4.130 24.300 4.320 ;
        RECT 23.970 4.090 24.290 4.130 ;
        RECT 24.960 3.990 25.160 4.590 ;
        RECT 25.680 4.000 25.900 4.590 ;
        RECT 6.570 3.620 6.770 3.970 ;
        RECT 25.690 3.970 25.900 4.000 ;
        RECT 8.050 3.800 8.390 3.870 ;
        RECT 8.050 3.700 8.490 3.800 ;
        RECT 8.160 3.580 8.490 3.700 ;
        RECT 8.170 3.540 8.490 3.580 ;
        RECT 6.940 3.160 7.380 3.330 ;
        RECT 8.170 2.910 8.490 2.950 ;
        RECT 6.570 2.520 6.770 2.870 ;
        RECT 8.160 2.790 8.490 2.910 ;
        RECT 8.050 2.690 8.490 2.790 ;
        RECT 8.050 2.620 8.390 2.690 ;
        RECT 9.310 2.670 9.480 3.680 ;
        RECT 13.240 2.810 13.410 3.820 ;
        RECT 19.050 2.810 19.220 3.820 ;
        RECT 24.070 3.800 24.410 3.870 ;
        RECT 23.970 3.700 24.410 3.800 ;
        RECT 22.980 2.670 23.150 3.680 ;
        RECT 23.970 3.580 24.300 3.700 ;
        RECT 25.690 3.620 25.890 3.970 ;
        RECT 23.970 3.540 24.290 3.580 ;
        RECT 25.080 3.160 25.520 3.330 ;
        RECT 23.970 2.910 24.290 2.950 ;
        RECT 23.970 2.790 24.300 2.910 ;
        RECT 23.970 2.690 24.410 2.790 ;
        RECT 24.070 2.620 24.410 2.690 ;
        RECT 6.560 2.490 6.770 2.520 ;
        RECT 25.690 2.520 25.890 2.870 ;
        RECT 6.560 1.900 6.780 2.490 ;
        RECT 7.300 1.900 7.500 2.500 ;
        RECT 8.170 2.360 8.490 2.400 ;
        RECT 8.160 2.170 8.490 2.360 ;
        RECT 8.050 2.140 8.490 2.170 ;
        RECT 23.970 2.360 24.290 2.400 ;
        RECT 23.970 2.170 24.300 2.360 ;
        RECT 23.970 2.140 24.410 2.170 ;
        RECT 8.050 2.000 8.390 2.140 ;
        RECT 24.070 2.000 24.410 2.140 ;
        RECT 24.960 1.900 25.160 2.500 ;
        RECT 25.690 2.490 25.900 2.520 ;
        RECT 25.680 1.900 25.900 2.490 ;
        RECT 6.560 0.770 6.780 1.360 ;
        RECT 6.560 0.740 6.770 0.770 ;
        RECT 7.300 0.760 7.500 1.360 ;
        RECT 8.050 1.120 8.390 1.260 ;
        RECT 24.070 1.120 24.410 1.260 ;
        RECT 8.050 1.090 8.490 1.120 ;
        RECT 8.160 0.900 8.490 1.090 ;
        RECT 8.170 0.860 8.490 0.900 ;
        RECT 23.970 1.090 24.410 1.120 ;
        RECT 23.970 0.900 24.300 1.090 ;
        RECT 23.970 0.860 24.290 0.900 ;
        RECT 24.960 0.760 25.160 1.360 ;
        RECT 25.680 0.770 25.900 1.360 ;
        RECT 6.570 0.390 6.770 0.740 ;
        RECT 25.690 0.740 25.900 0.770 ;
        RECT 8.050 0.570 8.390 0.640 ;
        RECT 24.070 0.570 24.410 0.640 ;
        RECT 8.050 0.470 8.490 0.570 ;
        RECT 8.160 0.350 8.490 0.470 ;
        RECT 8.170 0.310 8.490 0.350 ;
        RECT 23.970 0.470 24.410 0.570 ;
        RECT 23.970 0.350 24.300 0.470 ;
        RECT 25.690 0.390 25.890 0.740 ;
        RECT 23.970 0.310 24.290 0.350 ;
      LAYER mcon ;
        RECT 1.070 7.510 1.340 7.780 ;
        RECT 31.120 7.510 31.390 7.780 ;
        RECT 8.260 5.970 8.430 6.140 ;
        RECT 24.030 5.970 24.200 6.140 ;
        RECT 6.590 5.560 6.760 5.730 ;
        RECT 7.320 5.530 7.490 5.700 ;
        RECT 8.260 5.420 8.430 5.590 ;
        RECT 24.030 5.420 24.200 5.590 ;
        RECT 24.970 5.530 25.140 5.700 ;
        RECT 25.700 5.560 25.870 5.730 ;
        RECT 9.310 4.870 9.480 5.040 ;
        RECT 6.590 4.000 6.760 4.170 ;
        RECT 13.250 4.880 13.420 5.050 ;
        RECT 19.040 4.880 19.210 5.050 ;
        RECT 22.980 4.870 23.150 5.040 ;
        RECT 7.320 4.030 7.490 4.200 ;
        RECT 8.260 4.140 8.430 4.310 ;
        RECT 24.030 4.140 24.200 4.310 ;
        RECT 24.970 4.030 25.140 4.200 ;
        RECT 25.700 4.000 25.870 4.170 ;
        RECT 8.260 3.590 8.430 3.760 ;
        RECT 9.310 3.280 9.480 3.450 ;
        RECT 8.260 2.730 8.430 2.900 ;
        RECT 9.310 2.920 9.480 3.090 ;
        RECT 13.240 3.420 13.410 3.590 ;
        RECT 13.240 3.060 13.410 3.230 ;
        RECT 19.050 3.420 19.220 3.590 ;
        RECT 19.050 3.060 19.220 3.230 ;
        RECT 24.030 3.590 24.200 3.760 ;
        RECT 22.980 3.280 23.150 3.450 ;
        RECT 25.340 3.160 25.520 3.330 ;
        RECT 22.980 2.920 23.150 3.090 ;
        RECT 24.030 2.730 24.200 2.900 ;
        RECT 6.590 2.320 6.760 2.490 ;
        RECT 7.320 2.290 7.490 2.460 ;
        RECT 8.260 2.180 8.430 2.350 ;
        RECT 24.030 2.180 24.200 2.350 ;
        RECT 24.970 2.290 25.140 2.460 ;
        RECT 25.700 2.320 25.870 2.490 ;
        RECT 6.590 0.770 6.760 0.940 ;
        RECT 7.320 0.800 7.490 0.970 ;
        RECT 8.260 0.910 8.430 1.080 ;
        RECT 24.030 0.910 24.200 1.080 ;
        RECT 24.970 0.800 25.140 0.970 ;
        RECT 25.700 0.770 25.870 0.940 ;
        RECT 8.260 0.360 8.430 0.530 ;
        RECT 24.030 0.360 24.200 0.530 ;
      LAYER met1 ;
        RECT 1.010 6.970 1.400 8.830 ;
        RECT 31.060 6.970 31.450 8.830 ;
        RECT 8.180 5.900 8.500 6.220 ;
        RECT 23.960 5.900 24.280 6.220 ;
        RECT 8.180 5.350 8.500 5.670 ;
        RECT 23.960 5.350 24.280 5.670 ;
        RECT 8.180 4.060 8.500 4.380 ;
        RECT 23.960 4.060 24.280 4.380 ;
        RECT 8.180 3.510 8.500 3.830 ;
        RECT 23.960 3.510 24.280 3.830 ;
        RECT 8.180 2.660 8.500 2.980 ;
        RECT 23.960 2.660 24.280 2.980 ;
        RECT 8.180 2.110 8.500 2.430 ;
        RECT 23.960 2.110 24.280 2.430 ;
        RECT 8.180 0.830 8.500 1.150 ;
        RECT 23.960 0.830 24.280 1.150 ;
        RECT 8.180 0.280 8.500 0.600 ;
        RECT 23.960 0.280 24.280 0.600 ;
      LAYER via ;
        RECT 8.210 5.930 8.470 6.190 ;
        RECT 23.990 5.930 24.250 6.190 ;
        RECT 8.210 5.380 8.470 5.640 ;
        RECT 23.990 5.380 24.250 5.640 ;
        RECT 8.210 4.090 8.470 4.350 ;
        RECT 23.990 4.090 24.250 4.350 ;
        RECT 8.210 3.540 8.470 3.800 ;
        RECT 23.990 3.540 24.250 3.800 ;
        RECT 8.210 2.690 8.470 2.950 ;
        RECT 23.990 2.690 24.250 2.950 ;
        RECT 8.210 2.140 8.470 2.400 ;
        RECT 23.990 2.140 24.250 2.400 ;
        RECT 8.210 0.860 8.470 1.120 ;
        RECT 23.990 0.860 24.250 1.120 ;
        RECT 8.210 0.310 8.470 0.570 ;
        RECT 23.990 0.310 24.250 0.570 ;
      LAYER met2 ;
        RECT 8.610 5.760 23.850 5.940 ;
        RECT 8.640 5.500 8.730 5.510 ;
        RECT 23.730 5.500 23.820 5.510 ;
        RECT 8.610 5.320 23.850 5.500 ;
        RECT 8.610 4.220 23.850 4.400 ;
        RECT 8.610 3.790 23.850 3.970 ;
        RECT 8.620 2.520 23.840 2.700 ;
        RECT 8.610 2.090 23.850 2.270 ;
        RECT 8.620 0.990 23.840 1.170 ;
        RECT 8.640 0.570 23.820 0.740 ;
  END
END sky130_hilas_swc4x2cell

MACRO sky130_hilas_polyresistorGND
  CLASS CORE ;
  FOREIGN sky130_hilas_polyresistorGND ;
  ORIGIN 0.000 0.000 ;
  SIZE 55.470 BY 10.890 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN INPUT
    PORT
      LAYER met1 ;
        RECT 21.060 10.250 23.470 10.890 ;
        RECT 21.080 8.900 21.490 10.250 ;
    END
  END INPUT
  PIN OUTPUT
    ANTENNADIFFAREA 16.452000 ;
    PORT
      LAYER met2 ;
        RECT 0.000 7.380 55.470 8.770 ;
    END
  END OUTPUT
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 27.810 9.590 28.220 10.360 ;
        RECT 27.540 9.320 28.220 9.590 ;
        RECT 27.540 8.890 29.230 9.320 ;
        RECT 0.330 8.710 24.700 8.730 ;
        RECT 0.270 8.320 24.700 8.710 ;
        RECT 0.270 0.070 0.680 8.320 ;
        RECT 26.870 0.820 29.230 8.890 ;
        RECT 33.500 8.720 54.860 8.730 ;
        RECT 33.440 8.330 54.860 8.720 ;
        RECT 33.440 8.320 54.700 8.330 ;
        RECT 26.750 0.000 29.230 0.820 ;
      LAYER via ;
        RECT 0.820 8.410 24.620 8.670 ;
        RECT 33.500 8.410 54.360 8.670 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 21.140 9.120 21.360 10.240 ;
        RECT 21.090 8.930 21.420 9.120 ;
        RECT 27.880 8.930 28.120 10.280 ;
        RECT 0.380 8.460 55.120 8.730 ;
        RECT 0.380 8.330 24.720 8.460 ;
        RECT 33.410 8.330 55.120 8.460 ;
        RECT 0.380 0.730 0.550 8.330 ;
        RECT 54.950 1.250 55.120 8.330 ;
        RECT 26.820 0.390 29.180 0.560 ;
      LAYER mcon ;
        RECT 21.170 10.040 21.340 10.210 ;
        RECT 21.170 9.680 21.340 9.850 ;
        RECT 21.170 9.320 21.340 9.490 ;
        RECT 21.170 8.960 21.340 9.130 ;
        RECT 27.920 9.870 28.090 10.040 ;
        RECT 27.920 9.510 28.090 9.680 ;
        RECT 27.920 9.150 28.090 9.320 ;
        RECT 0.720 8.350 24.620 8.520 ;
        RECT 33.500 8.350 54.670 8.520 ;
        RECT 27.190 0.390 27.360 0.560 ;
        RECT 27.560 0.390 27.730 0.560 ;
        RECT 27.920 0.390 28.090 0.560 ;
        RECT 28.280 0.390 28.450 0.560 ;
        RECT 28.640 0.390 28.820 0.560 ;
        RECT 29.010 0.390 29.180 0.560 ;
      LAYER met2 ;
        RECT 0.000 1.080 55.470 2.480 ;
  END
END sky130_hilas_polyresistorGND

MACRO sky130_hilas_swc4x2cellOverlap
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x2cellOverlap ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.980 BY 6.160 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VERT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met1 ;
        RECT 1.170 5.420 1.330 6.150 ;
        RECT 1.130 5.400 1.330 5.420 ;
        RECT 1.120 5.160 1.350 5.400 ;
        RECT 1.120 5.110 1.330 5.160 ;
        RECT 1.170 4.050 1.330 5.110 ;
        RECT 1.120 4.000 1.330 4.050 ;
        RECT 1.120 3.760 1.350 4.000 ;
        RECT 1.130 3.740 1.330 3.760 ;
        RECT 1.170 2.410 1.330 3.740 ;
        RECT 1.130 2.390 1.330 2.410 ;
        RECT 1.120 2.150 1.350 2.390 ;
        RECT 1.120 2.100 1.330 2.150 ;
        RECT 1.170 1.050 1.330 2.100 ;
        RECT 1.120 1.000 1.330 1.050 ;
        RECT 1.120 0.760 1.350 1.000 ;
        RECT 1.130 0.740 1.330 0.760 ;
        RECT 1.170 0.010 1.330 0.740 ;
    END
  END VERT1
  PIN HORIZ1
    USE ANALOG ;
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT 2.160 5.170 2.470 5.190 ;
        RECT 15.500 5.170 15.810 5.190 ;
        RECT 0.000 4.990 17.980 5.170 ;
        RECT 2.160 4.860 2.470 4.990 ;
        RECT 15.500 4.860 15.810 4.990 ;
    END
  END HORIZ1
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT 2.160 5.600 2.470 5.740 ;
        RECT 15.500 5.600 15.810 5.740 ;
        RECT 0.000 5.420 17.970 5.600 ;
        RECT 2.160 5.410 2.470 5.420 ;
        RECT 15.500 5.410 15.810 5.420 ;
    END
  END DRAIN1
  PIN HORIZ2
    USE ANALOG ;
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT 2.160 4.170 2.470 4.300 ;
        RECT 15.500 4.170 15.810 4.300 ;
        RECT 0.000 3.990 17.980 4.170 ;
        RECT 2.160 3.970 2.470 3.990 ;
        RECT 15.500 3.970 15.810 3.990 ;
    END
  END HORIZ2
  PIN DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT 2.160 3.740 2.470 3.750 ;
        RECT 15.500 3.740 15.810 3.750 ;
        RECT 0.000 3.560 17.980 3.740 ;
        RECT 2.160 3.420 2.470 3.560 ;
        RECT 15.500 3.420 15.810 3.560 ;
    END
  END DRAIN2
  PIN DRAIN3
    USE ANALOG ;
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT 2.160 2.590 2.470 2.730 ;
        RECT 0.000 2.580 2.470 2.590 ;
        RECT 15.500 2.590 15.810 2.730 ;
        RECT 15.500 2.580 17.970 2.590 ;
        RECT 0.000 2.410 17.970 2.580 ;
        RECT 2.160 2.400 2.470 2.410 ;
        RECT 15.500 2.400 15.810 2.410 ;
    END
  END DRAIN3
  PIN HORIZ3
    USE ANALOG ;
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT 2.160 2.160 2.470 2.180 ;
        RECT 15.500 2.160 15.810 2.180 ;
        RECT 0.000 1.990 17.970 2.160 ;
        RECT 0.000 1.980 2.560 1.990 ;
        RECT 15.410 1.980 17.970 1.990 ;
        RECT 2.160 1.850 2.470 1.980 ;
        RECT 15.500 1.850 15.810 1.980 ;
    END
  END HORIZ3
  PIN HORIZ4
    USE ANALOG ;
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT 2.160 1.180 2.470 1.300 ;
        RECT 15.500 1.180 15.810 1.300 ;
        RECT 2.160 1.170 15.810 1.180 ;
        RECT 0.000 1.010 17.970 1.170 ;
        RECT 0.000 0.990 2.560 1.010 ;
        RECT 15.410 0.990 17.970 1.010 ;
        RECT 2.160 0.970 2.470 0.990 ;
        RECT 15.500 0.970 15.810 0.990 ;
    END
  END HORIZ4
  PIN DRAIN4
    USE ANALOG ;
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT 2.160 0.740 2.470 0.750 ;
        RECT 15.500 0.740 15.810 0.750 ;
        RECT 0.000 0.570 17.970 0.740 ;
        RECT 0.000 0.560 2.470 0.570 ;
        RECT 2.160 0.420 2.470 0.560 ;
        RECT 15.500 0.560 17.970 0.570 ;
        RECT 15.500 0.420 15.810 0.560 ;
    END
  END DRAIN4
  PIN VINJ
    ANTENNADIFFAREA 1.088000 ;
    PORT
      LAYER nwell ;
        RECT 0.000 6.100 2.560 6.160 ;
        RECT 0.000 0.050 6.560 6.100 ;
        RECT 0.000 0.000 2.560 0.050 ;
      LAYER met1 ;
        RECT 0.360 5.450 0.520 6.150 ;
        RECT 0.360 4.900 0.630 5.450 ;
        RECT 0.350 4.850 0.630 4.900 ;
        RECT 0.350 4.760 0.520 4.850 ;
        RECT 0.360 4.400 0.520 4.760 ;
        RECT 0.350 4.310 0.520 4.400 ;
        RECT 0.350 4.260 0.630 4.310 ;
        RECT 0.360 3.710 0.630 4.260 ;
        RECT 0.360 2.440 0.520 3.710 ;
        RECT 0.360 1.890 0.630 2.440 ;
        RECT 0.350 1.840 0.630 1.890 ;
        RECT 0.350 1.750 0.520 1.840 ;
        RECT 0.360 1.400 0.520 1.750 ;
        RECT 0.350 1.310 0.520 1.400 ;
        RECT 0.350 1.260 0.630 1.310 ;
        RECT 0.360 0.710 0.630 1.260 ;
        RECT 0.360 0.010 0.520 0.710 ;
    END
    PORT
      LAYER nwell ;
        RECT 15.410 6.100 17.970 6.160 ;
        RECT 11.410 0.050 17.970 6.100 ;
        RECT 15.410 0.000 17.970 0.050 ;
      LAYER met1 ;
        RECT 17.450 5.450 17.610 6.150 ;
        RECT 17.340 4.900 17.610 5.450 ;
        RECT 17.340 4.850 17.620 4.900 ;
        RECT 17.450 4.760 17.620 4.850 ;
        RECT 17.450 4.400 17.610 4.760 ;
        RECT 17.450 4.310 17.620 4.400 ;
        RECT 17.340 4.260 17.620 4.310 ;
        RECT 17.340 3.710 17.610 4.260 ;
        RECT 17.450 2.440 17.610 3.710 ;
        RECT 17.340 1.890 17.610 2.440 ;
        RECT 17.340 1.840 17.620 1.890 ;
        RECT 17.450 1.750 17.620 1.840 ;
        RECT 17.450 1.400 17.610 1.750 ;
        RECT 17.450 1.310 17.620 1.400 ;
        RECT 17.340 1.260 17.620 1.310 ;
        RECT 17.340 0.710 17.610 1.260 ;
        RECT 17.450 0.010 17.610 0.710 ;
    END
  END VINJ
  PIN GATESELECT1
    USE ANALOG ;
    ANTENNAGATEAREA 0.720000 ;
    PORT
      LAYER met1 ;
        RECT 0.770 5.110 0.960 6.100 ;
        RECT 0.770 4.990 0.940 5.110 ;
        RECT 0.770 4.170 0.930 4.990 ;
        RECT 0.770 4.050 0.940 4.170 ;
        RECT 0.770 3.190 0.960 4.050 ;
        RECT 0.740 2.960 0.980 3.190 ;
        RECT 0.770 2.100 0.960 2.960 ;
        RECT 0.770 1.980 0.940 2.100 ;
        RECT 0.770 1.170 0.930 1.980 ;
        RECT 0.770 1.050 0.940 1.170 ;
        RECT 0.770 0.060 0.960 1.050 ;
    END
  END GATESELECT1
  PIN VERT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met1 ;
        RECT 16.640 5.420 16.800 6.150 ;
        RECT 16.640 5.400 16.840 5.420 ;
        RECT 16.620 5.160 16.850 5.400 ;
        RECT 16.640 5.110 16.850 5.160 ;
        RECT 16.640 4.050 16.800 5.110 ;
        RECT 16.640 4.000 16.850 4.050 ;
        RECT 16.620 3.760 16.850 4.000 ;
        RECT 16.640 3.740 16.840 3.760 ;
        RECT 16.640 2.410 16.800 3.740 ;
        RECT 16.640 2.390 16.840 2.410 ;
        RECT 16.620 2.150 16.850 2.390 ;
        RECT 16.640 2.100 16.850 2.150 ;
        RECT 16.640 1.050 16.800 2.100 ;
        RECT 16.640 1.000 16.850 1.050 ;
        RECT 16.620 0.760 16.850 1.000 ;
        RECT 16.640 0.740 16.840 0.760 ;
        RECT 16.640 0.010 16.800 0.740 ;
    END
  END VERT2
  PIN GATESELECT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.720000 ;
    PORT
      LAYER met1 ;
        RECT 17.010 5.110 17.200 6.100 ;
        RECT 17.030 4.990 17.200 5.110 ;
        RECT 17.040 4.170 17.200 4.990 ;
        RECT 17.030 4.050 17.200 4.170 ;
        RECT 17.010 3.190 17.200 4.050 ;
        RECT 16.990 2.960 17.230 3.190 ;
        RECT 17.010 2.100 17.200 2.960 ;
        RECT 17.030 1.980 17.200 2.100 ;
        RECT 17.040 1.170 17.200 1.980 ;
        RECT 17.030 1.050 17.200 1.170 ;
        RECT 17.010 0.060 17.200 1.050 ;
    END
  END GATESELECT2
  PIN GATE2
    USE ANALOG ;
    ANTENNADIFFAREA 1.345600 ;
    PORT
      LAYER met1 ;
        RECT 13.290 4.870 13.530 6.100 ;
        RECT 13.290 4.650 13.540 4.870 ;
        RECT 13.290 3.400 13.530 4.650 ;
        RECT 13.290 3.180 13.540 3.400 ;
        RECT 13.290 1.930 13.530 3.180 ;
        RECT 13.290 1.710 13.540 1.930 ;
        RECT 13.290 0.460 13.530 1.710 ;
        RECT 13.290 0.240 13.540 0.460 ;
        RECT 13.290 0.050 13.530 0.240 ;
    END
  END GATE2
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 1.345600 ;
    PORT
      LAYER met1 ;
        RECT 4.440 4.870 4.690 6.100 ;
        RECT 4.430 4.650 4.690 4.870 ;
        RECT 4.440 3.400 4.690 4.650 ;
        RECT 4.430 3.180 4.690 3.400 ;
        RECT 4.440 1.930 4.690 3.180 ;
        RECT 4.430 1.710 4.690 1.930 ;
        RECT 4.440 0.460 4.690 1.710 ;
        RECT 4.430 0.240 4.690 0.460 ;
        RECT 4.440 0.050 4.690 0.240 ;
    END
  END GATE1
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 0.336400 ;
    PORT
      LAYER met1 ;
        RECT 8.050 0.050 8.350 6.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 9.630 0.050 9.930 6.100 ;
    END
  END VTUN
  OBS
      LAYER li1 ;
        RECT 0.400 5.420 0.600 5.770 ;
        RECT 2.140 5.690 2.460 5.700 ;
        RECT 1.880 5.520 2.460 5.690 ;
        RECT 2.130 5.470 2.460 5.520 ;
        RECT 2.140 5.440 2.460 5.470 ;
        RECT 0.390 5.390 0.600 5.420 ;
        RECT 0.390 4.800 0.610 5.390 ;
        RECT 1.130 4.800 1.330 5.400 ;
        RECT 2.140 5.110 2.460 5.150 ;
        RECT 2.130 5.070 2.460 5.110 ;
        RECT 1.880 4.900 2.460 5.070 ;
        RECT 2.140 4.890 2.460 4.900 ;
        RECT 2.900 4.790 6.210 5.770 ;
        RECT 8.120 4.890 8.290 5.780 ;
        RECT 9.680 4.890 9.850 5.780 ;
        RECT 11.760 4.790 15.070 5.770 ;
        RECT 15.510 5.690 15.830 5.700 ;
        RECT 15.510 5.520 16.090 5.690 ;
        RECT 15.510 5.470 15.840 5.520 ;
        RECT 15.510 5.440 15.830 5.470 ;
        RECT 17.370 5.420 17.570 5.770 ;
        RECT 15.510 5.110 15.830 5.150 ;
        RECT 15.510 5.070 15.840 5.110 ;
        RECT 15.510 4.900 16.090 5.070 ;
        RECT 15.510 4.890 15.830 4.900 ;
        RECT 16.640 4.800 16.840 5.400 ;
        RECT 17.370 5.390 17.580 5.420 ;
        RECT 17.360 4.800 17.580 5.390 ;
        RECT 0.390 3.770 0.610 4.360 ;
        RECT 0.390 3.740 0.600 3.770 ;
        RECT 1.130 3.760 1.330 4.360 ;
        RECT 2.140 4.260 2.460 4.270 ;
        RECT 1.880 4.090 2.460 4.260 ;
        RECT 2.130 4.050 2.460 4.090 ;
        RECT 2.140 4.010 2.460 4.050 ;
        RECT 0.400 3.390 0.600 3.740 ;
        RECT 2.140 3.690 2.460 3.720 ;
        RECT 2.130 3.640 2.460 3.690 ;
        RECT 1.880 3.470 2.460 3.640 ;
        RECT 2.140 3.460 2.460 3.470 ;
        RECT 2.900 3.320 6.210 4.300 ;
        RECT 8.120 3.370 8.290 4.260 ;
        RECT 9.680 3.370 9.850 4.260 ;
        RECT 11.760 3.320 15.070 4.300 ;
        RECT 15.510 4.260 15.830 4.270 ;
        RECT 15.510 4.090 16.090 4.260 ;
        RECT 15.510 4.050 15.840 4.090 ;
        RECT 15.510 4.010 15.830 4.050 ;
        RECT 16.640 3.760 16.840 4.360 ;
        RECT 17.360 3.770 17.580 4.360 ;
        RECT 17.370 3.740 17.580 3.770 ;
        RECT 15.510 3.690 15.830 3.720 ;
        RECT 15.510 3.640 15.840 3.690 ;
        RECT 15.510 3.470 16.090 3.640 ;
        RECT 15.510 3.460 15.830 3.470 ;
        RECT 17.370 3.390 17.570 3.740 ;
        RECT 0.770 2.990 1.210 3.160 ;
        RECT 16.760 2.990 17.200 3.160 ;
        RECT 0.400 2.410 0.600 2.760 ;
        RECT 2.140 2.680 2.460 2.690 ;
        RECT 1.880 2.510 2.460 2.680 ;
        RECT 2.130 2.460 2.460 2.510 ;
        RECT 2.140 2.430 2.460 2.460 ;
        RECT 0.390 2.380 0.600 2.410 ;
        RECT 0.390 1.790 0.610 2.380 ;
        RECT 1.130 1.790 1.330 2.390 ;
        RECT 2.140 2.100 2.460 2.140 ;
        RECT 2.130 2.060 2.460 2.100 ;
        RECT 1.880 1.890 2.460 2.060 ;
        RECT 2.140 1.880 2.460 1.890 ;
        RECT 2.900 1.850 6.210 2.830 ;
        RECT 8.120 1.920 8.290 2.810 ;
        RECT 9.680 1.920 9.850 2.810 ;
        RECT 11.760 1.850 15.070 2.830 ;
        RECT 15.510 2.680 15.830 2.690 ;
        RECT 15.510 2.510 16.090 2.680 ;
        RECT 15.510 2.460 15.840 2.510 ;
        RECT 15.510 2.430 15.830 2.460 ;
        RECT 17.370 2.410 17.570 2.760 ;
        RECT 15.510 2.100 15.830 2.140 ;
        RECT 15.510 2.060 15.840 2.100 ;
        RECT 15.510 1.890 16.090 2.060 ;
        RECT 15.510 1.880 15.830 1.890 ;
        RECT 16.640 1.790 16.840 2.390 ;
        RECT 17.370 2.380 17.580 2.410 ;
        RECT 17.360 1.790 17.580 2.380 ;
        RECT 0.390 0.770 0.610 1.360 ;
        RECT 0.390 0.740 0.600 0.770 ;
        RECT 1.130 0.760 1.330 1.360 ;
        RECT 2.140 1.260 2.460 1.270 ;
        RECT 1.880 1.090 2.460 1.260 ;
        RECT 2.130 1.050 2.460 1.090 ;
        RECT 2.140 1.010 2.460 1.050 ;
        RECT 0.400 0.390 0.600 0.740 ;
        RECT 2.140 0.690 2.460 0.720 ;
        RECT 2.130 0.640 2.460 0.690 ;
        RECT 1.880 0.470 2.460 0.640 ;
        RECT 2.140 0.460 2.460 0.470 ;
        RECT 2.900 0.380 6.210 1.360 ;
        RECT 8.120 0.380 8.290 1.270 ;
        RECT 9.680 0.380 9.850 1.270 ;
        RECT 11.760 0.380 15.070 1.360 ;
        RECT 15.510 1.260 15.830 1.270 ;
        RECT 15.510 1.090 16.090 1.260 ;
        RECT 15.510 1.050 15.840 1.090 ;
        RECT 15.510 1.010 15.830 1.050 ;
        RECT 16.640 0.760 16.840 1.360 ;
        RECT 17.360 0.770 17.580 1.360 ;
        RECT 17.370 0.740 17.580 0.770 ;
        RECT 15.510 0.690 15.830 0.720 ;
        RECT 15.510 0.640 15.840 0.690 ;
        RECT 15.510 0.470 16.090 0.640 ;
        RECT 15.510 0.460 15.830 0.470 ;
        RECT 17.370 0.390 17.570 0.740 ;
      LAYER mcon ;
        RECT 2.230 5.480 2.400 5.650 ;
        RECT 4.470 5.540 4.640 5.710 ;
        RECT 0.420 5.220 0.590 5.390 ;
        RECT 1.150 5.190 1.320 5.360 ;
        RECT 2.230 4.930 2.400 5.100 ;
        RECT 4.470 4.850 4.640 5.020 ;
        RECT 8.120 5.580 8.290 5.750 ;
        RECT 9.680 5.580 9.850 5.750 ;
        RECT 13.330 5.540 13.500 5.710 ;
        RECT 15.570 5.480 15.740 5.650 ;
        RECT 16.650 5.190 16.820 5.360 ;
        RECT 13.330 4.850 13.500 5.020 ;
        RECT 15.570 4.930 15.740 5.100 ;
        RECT 17.380 5.220 17.550 5.390 ;
        RECT 0.420 3.770 0.590 3.940 ;
        RECT 2.230 4.060 2.400 4.230 ;
        RECT 4.470 4.070 4.640 4.240 ;
        RECT 1.150 3.800 1.320 3.970 ;
        RECT 2.230 3.510 2.400 3.680 ;
        RECT 4.470 3.380 4.640 3.550 ;
        RECT 8.120 4.060 8.290 4.230 ;
        RECT 9.680 4.060 9.850 4.230 ;
        RECT 13.330 4.070 13.500 4.240 ;
        RECT 15.570 4.060 15.740 4.230 ;
        RECT 16.650 3.800 16.820 3.970 ;
        RECT 17.380 3.770 17.550 3.940 ;
        RECT 13.330 3.380 13.500 3.550 ;
        RECT 15.570 3.510 15.740 3.680 ;
        RECT 17.020 2.990 17.200 3.160 ;
        RECT 2.230 2.470 2.400 2.640 ;
        RECT 4.470 2.600 4.640 2.770 ;
        RECT 0.420 2.210 0.590 2.380 ;
        RECT 1.150 2.180 1.320 2.350 ;
        RECT 2.230 1.920 2.400 2.090 ;
        RECT 4.470 1.910 4.640 2.080 ;
        RECT 8.120 2.610 8.290 2.780 ;
        RECT 9.680 2.610 9.850 2.780 ;
        RECT 13.330 2.600 13.500 2.770 ;
        RECT 15.570 2.470 15.740 2.640 ;
        RECT 16.650 2.180 16.820 2.350 ;
        RECT 13.330 1.910 13.500 2.080 ;
        RECT 15.570 1.920 15.740 2.090 ;
        RECT 17.380 2.210 17.550 2.380 ;
        RECT 0.420 0.770 0.590 0.940 ;
        RECT 2.230 1.060 2.400 1.230 ;
        RECT 4.470 1.130 4.640 1.300 ;
        RECT 1.150 0.800 1.320 0.970 ;
        RECT 2.230 0.510 2.400 0.680 ;
        RECT 4.470 0.440 4.640 0.610 ;
        RECT 8.120 1.070 8.290 1.240 ;
        RECT 9.680 1.070 9.850 1.240 ;
        RECT 13.330 1.130 13.500 1.300 ;
        RECT 15.570 1.060 15.740 1.230 ;
        RECT 16.650 0.800 16.820 0.970 ;
        RECT 17.380 0.770 17.550 0.940 ;
        RECT 13.330 0.440 13.500 0.610 ;
        RECT 15.570 0.510 15.740 0.680 ;
      LAYER met1 ;
        RECT 2.150 5.410 2.470 5.730 ;
        RECT 15.500 5.410 15.820 5.730 ;
        RECT 2.150 4.860 2.470 5.180 ;
        RECT 15.500 4.860 15.820 5.180 ;
        RECT 2.150 3.980 2.470 4.300 ;
        RECT 15.500 3.980 15.820 4.300 ;
        RECT 2.150 3.430 2.470 3.750 ;
        RECT 15.500 3.430 15.820 3.750 ;
        RECT 2.150 2.400 2.470 2.720 ;
        RECT 15.500 2.400 15.820 2.720 ;
        RECT 2.150 1.850 2.470 2.170 ;
        RECT 15.500 1.850 15.820 2.170 ;
        RECT 2.150 0.980 2.470 1.300 ;
        RECT 15.500 0.980 15.820 1.300 ;
        RECT 2.150 0.430 2.470 0.750 ;
        RECT 15.500 0.430 15.820 0.750 ;
      LAYER via ;
        RECT 2.180 5.440 2.440 5.700 ;
        RECT 15.530 5.440 15.790 5.700 ;
        RECT 2.180 4.890 2.440 5.150 ;
        RECT 15.530 4.890 15.790 5.150 ;
        RECT 2.180 4.010 2.440 4.270 ;
        RECT 15.530 4.010 15.790 4.270 ;
        RECT 2.180 3.460 2.440 3.720 ;
        RECT 15.530 3.460 15.790 3.720 ;
        RECT 2.180 2.430 2.440 2.690 ;
        RECT 15.530 2.430 15.790 2.690 ;
        RECT 2.180 1.880 2.440 2.140 ;
        RECT 15.530 1.880 15.790 2.140 ;
        RECT 2.180 1.010 2.440 1.270 ;
        RECT 15.530 1.010 15.790 1.270 ;
        RECT 2.180 0.460 2.440 0.720 ;
        RECT 15.530 0.460 15.790 0.720 ;
  END
END sky130_hilas_swc4x2cellOverlap

MACRO sky130_hilas_FGBias2x1cell
  CLASS CORE ;
  FOREIGN sky130_hilas_FGBias2x1cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 10.100 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VTUN
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 0.350 0.050 0.770 6.100 ;
    END
  END VTUN
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2.830 3.240 3.060 6.100 ;
        RECT 2.830 2.950 3.160 3.240 ;
        RECT 2.830 0.050 3.060 2.950 ;
    END
  END VGND
  PIN GATE_CONTROL
    USE ANALOG ;
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT 3.770 3.710 6.490 5.360 ;
        RECT 3.770 3.670 6.480 3.710 ;
        RECT 3.770 2.340 6.480 2.380 ;
        RECT 3.770 0.690 6.490 2.340 ;
      LAYER met1 ;
        RECT 4.050 4.890 4.280 6.100 ;
        RECT 4.050 4.100 4.310 4.890 ;
        RECT 4.050 1.950 4.280 4.100 ;
        RECT 4.050 1.160 4.310 1.950 ;
        RECT 4.050 0.050 4.280 1.160 ;
    END
  END GATE_CONTROL
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 9.050 5.600 9.360 5.610 ;
        RECT 0.000 5.420 11.530 5.600 ;
        RECT 9.050 5.280 9.360 5.420 ;
    END
  END DRAIN1
  PIN DRAIN4
    USE ANALOG ;
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 9.050 0.730 9.360 0.870 ;
        RECT 9.050 0.720 11.530 0.730 ;
        RECT 0.000 0.570 11.530 0.720 ;
        RECT 9.050 0.550 11.530 0.570 ;
        RECT 9.050 0.540 9.360 0.550 ;
    END
  END DRAIN4
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 8.220 0.000 11.530 6.150 ;
      LAYER met2 ;
        RECT 10.140 3.240 10.460 3.500 ;
        RECT 10.180 3.220 11.360 3.240 ;
        RECT 10.180 2.960 11.400 3.220 ;
        RECT 10.180 2.900 11.360 2.960 ;
        RECT 10.140 2.890 11.360 2.900 ;
        RECT 10.140 2.640 10.460 2.890 ;
    END
  END VINJ
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 9.340 4.580 9.650 4.800 ;
        RECT 9.340 4.470 11.530 4.580 ;
        RECT 9.500 4.360 11.530 4.470 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 9.340 1.820 9.650 2.040 ;
        RECT 9.340 1.710 11.530 1.820 ;
        RECT 9.490 1.610 11.530 1.710 ;
    END
  END OUTPUT2
  PIN GATECOL
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT 10.570 4.640 10.760 6.100 ;
        RECT 10.570 4.610 10.790 4.640 ;
        RECT 10.550 4.340 10.800 4.610 ;
        RECT 10.560 4.330 10.800 4.340 ;
        RECT 10.560 4.090 10.790 4.330 ;
        RECT 10.600 2.060 10.760 4.090 ;
        RECT 10.560 1.820 10.790 2.060 ;
        RECT 10.560 1.810 10.800 1.820 ;
        RECT 10.550 1.540 10.800 1.810 ;
        RECT 10.570 1.510 10.790 1.540 ;
        RECT 10.570 0.050 10.760 1.510 ;
    END
  END GATECOL
  PIN VINJ
    ANTENNADIFFAREA 0.544000 ;
    PORT
      LAYER met1 ;
        RECT 11.010 5.450 11.290 6.100 ;
        RECT 10.900 4.850 11.290 5.450 ;
        RECT 11.010 3.250 11.290 4.850 ;
        RECT 11.010 2.930 11.370 3.250 ;
        RECT 11.010 1.300 11.290 2.930 ;
        RECT 10.900 0.700 11.290 1.300 ;
        RECT 11.010 0.050 11.290 0.700 ;
      LAYER via ;
        RECT 11.110 2.960 11.370 3.220 ;
    END
  END VINJ
  OBS
      LAYER nwell ;
        RECT 14.520 9.760 16.250 10.100 ;
        RECT 14.500 8.200 16.250 9.760 ;
        RECT 14.500 6.190 16.230 8.200 ;
        RECT 14.520 4.060 16.250 5.960 ;
        RECT 0.590 1.450 1.150 3.870 ;
      LAYER li1 ;
        RECT 14.920 8.370 15.470 8.800 ;
        RECT 14.920 6.640 15.470 7.070 ;
        RECT 9.120 5.520 9.650 5.690 ;
        RECT 10.930 5.420 11.130 5.770 ;
        RECT 10.930 5.390 11.140 5.420 ;
        RECT 4.070 4.150 4.300 4.840 ;
        RECT 9.370 4.760 9.540 5.130 ;
        RECT 9.350 4.720 9.670 4.760 ;
        RECT 9.350 4.530 9.680 4.720 ;
        RECT 9.350 4.500 9.670 4.530 ;
        RECT 3.040 3.210 3.230 3.530 ;
        RECT 9.370 3.440 9.540 4.500 ;
        RECT 10.200 3.530 10.370 5.140 ;
        RECT 10.920 4.810 11.140 5.390 ;
        RECT 10.930 4.800 11.140 4.810 ;
        RECT 10.570 4.630 10.760 4.640 ;
        RECT 10.570 4.340 10.770 4.630 ;
        RECT 10.560 4.010 10.850 4.340 ;
        RECT 10.200 3.340 10.380 3.530 ;
        RECT 2.950 3.120 3.230 3.210 ;
        RECT 2.950 2.980 6.590 3.120 ;
        RECT 3.040 2.940 6.590 2.980 ;
        RECT 3.040 2.520 3.230 2.940 ;
        RECT 9.370 2.000 9.540 2.710 ;
        RECT 10.200 2.620 10.380 2.810 ;
        RECT 9.350 1.960 9.670 2.000 ;
        RECT 4.070 1.210 4.300 1.940 ;
        RECT 9.350 1.770 9.680 1.960 ;
        RECT 9.350 1.740 9.670 1.770 ;
        RECT 9.370 1.020 9.540 1.740 ;
        RECT 10.200 1.010 10.370 2.620 ;
        RECT 10.560 1.810 10.850 2.140 ;
        RECT 10.570 1.520 10.770 1.810 ;
        RECT 10.570 1.510 10.760 1.520 ;
        RECT 10.930 1.340 11.140 1.350 ;
        RECT 10.920 0.760 11.140 1.340 ;
        RECT 10.930 0.730 11.140 0.760 ;
        RECT 9.120 0.460 9.650 0.630 ;
        RECT 10.930 0.380 11.130 0.730 ;
      LAYER mcon ;
        RECT 14.920 8.450 15.190 8.720 ;
        RECT 14.920 6.720 15.190 6.990 ;
        RECT 10.940 5.220 11.110 5.390 ;
        RECT 4.100 4.640 4.270 4.810 ;
        RECT 9.410 4.540 9.580 4.710 ;
        RECT 4.100 4.190 4.270 4.360 ;
        RECT 10.580 4.380 10.760 4.570 ;
        RECT 2.960 3.010 3.130 3.180 ;
        RECT 4.100 1.690 4.270 1.860 ;
        RECT 9.410 1.780 9.580 1.950 ;
        RECT 4.100 1.240 4.270 1.410 ;
        RECT 10.580 1.580 10.760 1.770 ;
        RECT 10.940 0.760 11.110 0.930 ;
      LAYER met1 ;
        RECT 14.860 6.180 15.250 9.770 ;
        RECT 9.050 5.280 9.360 5.720 ;
        RECT 9.340 4.470 9.660 4.790 ;
        RECT 10.170 3.530 10.410 3.660 ;
        RECT 10.170 3.210 10.430 3.530 ;
        RECT 10.170 2.610 10.430 2.930 ;
        RECT 10.170 2.490 10.410 2.610 ;
        RECT 9.340 1.710 9.660 2.030 ;
        RECT 9.050 0.430 9.360 0.870 ;
      LAYER via ;
        RECT 9.080 5.310 9.340 5.570 ;
        RECT 9.370 4.500 9.630 4.760 ;
        RECT 10.170 3.240 10.430 3.500 ;
        RECT 10.170 2.640 10.430 2.900 ;
        RECT 9.370 1.740 9.630 2.000 ;
        RECT 9.080 0.580 9.340 0.840 ;
  END
END sky130_hilas_FGBias2x1cell

MACRO sky130_hilas_drainSelect01
  CLASS CORE ;
  FOREIGN sky130_hilas_drainSelect01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.720 BY 6.590 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DRAIN3
    ANTENNADIFFAREA 0.322600 ;
    PORT
      LAYER met2 ;
        RECT 1.750 2.960 2.070 2.980 ;
        RECT 4.160 2.960 4.480 3.010 ;
        RECT 0.000 2.860 0.570 2.870 ;
        RECT 0.000 2.850 1.270 2.860 ;
        RECT 1.750 2.850 4.480 2.960 ;
        RECT 0.000 2.770 4.480 2.850 ;
        RECT 0.000 2.720 2.070 2.770 ;
        RECT 0.000 2.690 2.000 2.720 ;
        RECT 4.160 2.690 4.480 2.770 ;
    END
  END DRAIN3
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.000 0.000 3.420 6.590 ;
      LAYER met1 ;
        RECT 0.580 6.320 0.830 6.540 ;
        RECT 0.190 5.250 0.830 6.320 ;
        RECT 0.580 4.540 0.830 5.250 ;
        RECT 0.190 3.470 0.830 4.540 ;
        RECT 0.580 3.120 0.830 3.470 ;
        RECT 0.190 2.050 0.830 3.120 ;
        RECT 0.580 1.340 0.830 2.050 ;
        RECT 0.190 0.270 0.830 1.340 ;
        RECT 0.580 0.050 0.830 0.270 ;
    END
  END VINJ
  PIN DRAIN_MUX
    USE ANALOG ;
    ANTENNADIFFAREA 0.846400 ;
    PORT
      LAYER met1 ;
        RECT 3.570 0.050 3.800 6.540 ;
    END
  END DRAIN_MUX
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 4.920 6.320 5.110 6.540 ;
        RECT 4.920 5.830 5.390 6.320 ;
        RECT 4.920 5.490 5.110 5.830 ;
        RECT 4.920 5.200 5.210 5.490 ;
        RECT 4.920 4.590 5.110 5.200 ;
        RECT 4.920 4.300 5.210 4.590 ;
        RECT 4.920 3.960 5.110 4.300 ;
        RECT 4.920 3.470 5.390 3.960 ;
        RECT 4.920 3.120 5.110 3.470 ;
        RECT 4.920 2.630 5.390 3.120 ;
        RECT 4.920 2.290 5.110 2.630 ;
        RECT 4.920 2.000 5.210 2.290 ;
        RECT 4.920 1.390 5.110 2.000 ;
        RECT 4.920 1.100 5.210 1.390 ;
        RECT 4.920 0.760 5.110 1.100 ;
        RECT 4.920 0.270 5.390 0.760 ;
        RECT 4.920 0.050 5.110 0.270 ;
    END
  END VGND
  PIN SELECT2
    ANTENNAGATEAREA 0.730000 ;
    PORT
      LAYER met2 ;
        RECT 5.240 4.350 5.580 4.410 ;
        RECT 5.240 4.110 5.720 4.350 ;
    END
  END SELECT2
  PIN SELECT1
    ANTENNAGATEAREA 0.730000 ;
    PORT
      LAYER met2 ;
        RECT 5.240 5.450 5.720 5.680 ;
        RECT 5.240 5.380 5.580 5.450 ;
    END
  END SELECT1
  PIN SELECT3
    ANTENNAGATEAREA 0.730000 ;
    PORT
      LAYER met2 ;
        RECT 5.240 2.250 5.720 2.480 ;
        RECT 5.240 2.180 5.580 2.250 ;
    END
  END SELECT3
  PIN SELECT4
    ANTENNAGATEAREA 0.730000 ;
    PORT
      LAYER met2 ;
        RECT 5.240 1.140 5.580 1.210 ;
        RECT 5.240 0.910 5.720 1.140 ;
    END
  END SELECT4
  OBS
      LAYER li1 ;
        RECT 0.220 5.370 0.390 6.260 ;
        RECT 0.620 5.280 0.790 6.210 ;
        RECT 4.310 6.140 4.550 6.170 ;
        RECT 1.320 5.970 2.280 6.140 ;
        RECT 2.730 5.970 4.070 6.140 ;
        RECT 4.310 5.970 4.880 6.140 ;
        RECT 1.600 5.960 1.770 5.970 ;
        RECT 4.310 5.930 4.550 5.970 ;
        RECT 5.190 5.840 5.360 6.260 ;
        RECT 1.800 5.520 2.140 5.700 ;
        RECT 5.260 5.620 5.430 5.660 ;
        RECT 1.320 5.350 4.070 5.520 ;
        RECT 4.530 5.350 4.900 5.520 ;
        RECT 5.000 5.230 5.190 5.460 ;
        RECT 5.260 5.450 5.490 5.620 ;
        RECT 5.260 5.100 5.430 5.450 ;
        RECT 0.220 3.530 0.390 4.420 ;
        RECT 0.620 3.580 0.790 4.510 ;
        RECT 1.320 4.270 4.070 4.440 ;
        RECT 4.530 4.270 4.900 4.440 ;
        RECT 5.000 4.330 5.190 4.560 ;
        RECT 5.260 4.340 5.430 4.690 ;
        RECT 1.800 4.090 2.140 4.270 ;
        RECT 5.260 4.170 5.490 4.340 ;
        RECT 5.260 4.130 5.430 4.170 ;
        RECT 1.600 3.820 1.770 3.830 ;
        RECT 4.310 3.820 4.550 3.860 ;
        RECT 1.320 3.650 2.280 3.820 ;
        RECT 2.730 3.650 4.070 3.820 ;
        RECT 4.310 3.650 4.880 3.820 ;
        RECT 4.310 3.620 4.550 3.650 ;
        RECT 5.190 3.530 5.360 3.950 ;
        RECT 0.220 2.170 0.390 3.060 ;
        RECT 0.620 2.080 0.790 3.010 ;
        RECT 4.310 2.940 4.550 2.970 ;
        RECT 1.320 2.770 2.280 2.940 ;
        RECT 2.730 2.770 4.070 2.940 ;
        RECT 4.310 2.770 4.880 2.940 ;
        RECT 1.600 2.760 1.770 2.770 ;
        RECT 4.310 2.730 4.550 2.770 ;
        RECT 5.190 2.640 5.360 3.060 ;
        RECT 1.800 2.320 2.140 2.500 ;
        RECT 5.260 2.420 5.430 2.460 ;
        RECT 1.320 2.150 4.070 2.320 ;
        RECT 4.530 2.150 4.900 2.320 ;
        RECT 5.000 2.030 5.190 2.260 ;
        RECT 5.260 2.250 5.490 2.420 ;
        RECT 5.260 1.900 5.430 2.250 ;
        RECT 0.220 0.330 0.390 1.220 ;
        RECT 0.620 0.380 0.790 1.310 ;
        RECT 1.320 1.070 4.070 1.240 ;
        RECT 4.530 1.070 4.900 1.240 ;
        RECT 5.000 1.130 5.190 1.360 ;
        RECT 5.260 1.140 5.430 1.490 ;
        RECT 1.800 0.890 2.140 1.070 ;
        RECT 5.260 0.970 5.490 1.140 ;
        RECT 5.260 0.930 5.430 0.970 ;
        RECT 1.600 0.620 1.770 0.630 ;
        RECT 4.310 0.620 4.550 0.660 ;
        RECT 1.320 0.450 2.280 0.620 ;
        RECT 2.730 0.450 4.070 0.620 ;
        RECT 4.310 0.450 4.880 0.620 ;
        RECT 4.310 0.420 4.550 0.450 ;
        RECT 5.190 0.330 5.360 0.750 ;
      LAYER mcon ;
        RECT 0.220 6.090 0.390 6.260 ;
        RECT 0.220 5.730 0.390 5.900 ;
        RECT 3.600 5.970 3.770 6.140 ;
        RECT 4.350 5.970 4.520 6.140 ;
        RECT 5.190 6.090 5.360 6.260 ;
        RECT 0.620 5.640 0.790 5.810 ;
        RECT 5.010 5.260 5.180 5.430 ;
        RECT 5.320 5.450 5.490 5.620 ;
        RECT 0.220 4.250 0.390 4.420 ;
        RECT 0.220 3.890 0.390 4.060 ;
        RECT 5.010 4.360 5.180 4.530 ;
        RECT 0.620 3.980 0.790 4.150 ;
        RECT 5.320 4.170 5.490 4.340 ;
        RECT 1.600 3.660 1.770 3.830 ;
        RECT 3.600 3.650 3.770 3.820 ;
        RECT 4.350 3.650 4.520 3.820 ;
        RECT 0.220 2.890 0.390 3.060 ;
        RECT 0.220 2.530 0.390 2.700 ;
        RECT 3.600 2.770 3.770 2.940 ;
        RECT 4.350 2.770 4.520 2.940 ;
        RECT 5.190 2.890 5.360 3.060 ;
        RECT 0.620 2.440 0.790 2.610 ;
        RECT 5.010 2.060 5.180 2.230 ;
        RECT 5.320 2.250 5.490 2.420 ;
        RECT 0.220 1.050 0.390 1.220 ;
        RECT 0.220 0.690 0.390 0.860 ;
        RECT 5.010 1.160 5.180 1.330 ;
        RECT 0.620 0.780 0.790 0.950 ;
        RECT 5.320 0.970 5.490 1.140 ;
        RECT 1.600 0.460 1.770 0.630 ;
        RECT 3.600 0.450 3.770 0.620 ;
        RECT 4.350 0.450 4.520 0.620 ;
      LAYER met1 ;
        RECT 1.730 6.160 2.070 6.210 ;
        RECT 1.510 6.140 2.070 6.160 ;
        RECT 4.160 6.180 4.530 6.200 ;
        RECT 1.510 5.970 2.190 6.140 ;
        RECT 1.510 5.930 2.070 5.970 ;
        RECT 1.730 5.890 2.070 5.930 ;
        RECT 4.160 5.920 4.580 6.180 ;
        RECT 4.160 5.910 4.530 5.920 ;
        RECT 5.250 5.390 5.570 5.670 ;
        RECT 5.250 4.120 5.570 4.400 ;
        RECT 1.730 3.860 2.070 3.900 ;
        RECT 1.510 3.820 2.070 3.860 ;
        RECT 4.160 3.870 4.530 3.880 ;
        RECT 1.510 3.650 2.190 3.820 ;
        RECT 1.510 3.630 2.070 3.650 ;
        RECT 1.730 3.580 2.070 3.630 ;
        RECT 4.160 3.610 4.580 3.870 ;
        RECT 4.160 3.590 4.530 3.610 ;
        RECT 1.730 2.960 2.070 3.010 ;
        RECT 1.510 2.940 2.070 2.960 ;
        RECT 4.160 2.980 4.530 3.000 ;
        RECT 1.510 2.770 2.190 2.940 ;
        RECT 1.510 2.730 2.070 2.770 ;
        RECT 1.730 2.690 2.070 2.730 ;
        RECT 4.160 2.720 4.580 2.980 ;
        RECT 4.160 2.710 4.530 2.720 ;
        RECT 5.250 2.190 5.570 2.470 ;
        RECT 5.250 0.920 5.570 1.200 ;
        RECT 1.730 0.660 2.070 0.700 ;
        RECT 1.510 0.620 2.070 0.660 ;
        RECT 4.160 0.670 4.530 0.680 ;
        RECT 1.510 0.450 2.190 0.620 ;
        RECT 1.510 0.430 2.070 0.450 ;
        RECT 1.730 0.380 2.070 0.430 ;
        RECT 4.160 0.410 4.580 0.670 ;
        RECT 4.160 0.390 4.530 0.410 ;
      LAYER via ;
        RECT 1.780 5.920 2.040 6.180 ;
        RECT 4.190 5.920 4.450 6.180 ;
        RECT 5.280 5.400 5.540 5.660 ;
        RECT 5.280 4.130 5.540 4.390 ;
        RECT 1.780 3.610 2.040 3.870 ;
        RECT 4.190 3.610 4.450 3.870 ;
        RECT 1.780 2.720 2.040 2.980 ;
        RECT 4.190 2.720 4.450 2.980 ;
        RECT 5.280 2.200 5.540 2.460 ;
        RECT 5.280 0.930 5.540 1.190 ;
        RECT 1.780 0.410 2.040 0.670 ;
        RECT 4.190 0.410 4.450 0.670 ;
      LAYER met2 ;
        RECT 1.750 6.160 2.070 6.180 ;
        RECT 4.160 6.160 4.480 6.210 ;
        RECT 1.750 6.130 4.480 6.160 ;
        RECT 0.000 5.970 4.480 6.130 ;
        RECT 0.000 5.950 2.070 5.970 ;
        RECT 1.750 5.920 2.070 5.950 ;
        RECT 4.160 5.890 4.480 5.970 ;
        RECT 1.750 3.820 2.070 3.870 ;
        RECT 4.160 3.820 4.480 3.900 ;
        RECT 1.750 3.810 4.480 3.820 ;
        RECT 0.000 3.650 4.480 3.810 ;
        RECT 1.750 3.630 4.480 3.650 ;
        RECT 1.750 3.610 2.070 3.630 ;
        RECT 4.160 3.580 4.480 3.630 ;
        RECT 1.750 0.620 2.070 0.670 ;
        RECT 4.160 0.620 4.480 0.700 ;
        RECT 1.750 0.600 4.480 0.620 ;
        RECT 0.000 0.430 4.480 0.600 ;
        RECT 1.750 0.410 2.070 0.430 ;
        RECT 4.160 0.380 4.480 0.430 ;
  END
END sky130_hilas_drainSelect01

MACRO sky130_hilas_DAC5bit01
  CLASS CORE ;
  FOREIGN sky130_hilas_DAC5bit01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.580 BY 7.410 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 8.350 0.980 8.670 1.110 ;
        RECT 0.000 0.850 8.670 0.980 ;
        RECT 0.000 0.780 8.540 0.850 ;
    END
  END A0
  PIN A1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 11.710 2.100 11.860 5.840 ;
        RECT 0.000 1.900 11.870 2.100 ;
        RECT 0.000 1.890 0.140 1.900 ;
    END
  END A1
  PIN A2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 10.110 3.080 10.310 5.680 ;
        RECT 0.000 2.870 10.310 3.080 ;
        RECT 0.320 2.670 0.640 2.870 ;
    END
  END A2
  PIN A3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 4.950 2.060 5.010 ;
        RECT 3.480 4.950 3.700 5.410 ;
        RECT 8.400 4.960 8.650 5.720 ;
        RECT 8.400 4.950 8.680 4.960 ;
        RECT 0.000 4.800 8.680 4.950 ;
        RECT 0.260 4.560 0.620 4.800 ;
        RECT 1.900 4.650 8.680 4.800 ;
    END
  END A3
  PIN A4
    USE ANALOG ;
    ANTENNAGATEAREA 2.933400 ;
    ANTENNADIFFAREA 1.649500 ;
    PORT
      LAYER met2 ;
        RECT 0.320 5.960 0.640 6.190 ;
        RECT 2.030 5.960 2.350 6.230 ;
        RECT 5.230 5.960 5.550 6.230 ;
        RECT 6.840 5.960 7.160 6.240 ;
        RECT 12.970 5.960 13.280 5.980 ;
        RECT 13.640 5.960 13.950 5.980 ;
        RECT 0.000 5.920 7.160 5.960 ;
        RECT 0.000 5.770 7.050 5.920 ;
        RECT 0.000 5.750 0.290 5.770 ;
        RECT 12.710 5.680 13.950 5.960 ;
        RECT 12.970 5.650 13.280 5.680 ;
        RECT 13.460 5.670 13.950 5.680 ;
        RECT 13.640 5.650 13.950 5.670 ;
        RECT 3.750 5.150 4.070 5.470 ;
    END
  END A4
  PIN VPWR
    USE ANALOG ;
    ANTENNAGATEAREA 2.529900 ;
    ANTENNADIFFAREA 1.583800 ;
    PORT
      LAYER met1 ;
        RECT 2.030 5.910 2.350 6.230 ;
        RECT 2.070 5.680 2.300 5.910 ;
        RECT 12.970 5.650 13.290 5.970 ;
        RECT 13.640 5.650 13.960 5.970 ;
        RECT 3.750 5.430 4.070 5.470 ;
        RECT 3.520 5.200 4.070 5.430 ;
        RECT 3.750 5.150 4.070 5.200 ;
      LAYER via ;
        RECT 2.060 5.940 2.320 6.200 ;
        RECT 13.000 5.680 13.260 5.940 ;
        RECT 13.670 5.680 13.930 5.940 ;
        RECT 3.780 5.180 4.040 5.440 ;
    END
  END VPWR
  PIN OUT
    USE ANALOG ;
    ANTENNADIFFAREA 0.365200 ;
    PORT
      LAYER met1 ;
        RECT 3.110 0.230 3.340 0.360 ;
        RECT 4.730 0.230 4.960 0.360 ;
        RECT 6.330 0.230 6.560 0.360 ;
        RECT 7.950 0.230 8.180 0.360 ;
        RECT 9.550 0.230 9.780 0.360 ;
        RECT 11.170 0.230 11.400 0.360 ;
        RECT 12.770 0.230 13.000 0.360 ;
        RECT 14.380 0.230 14.610 0.360 ;
        RECT 3.040 0.000 16.580 0.230 ;
    END
  END OUT
  OBS
      LAYER nwell ;
        RECT 0.890 6.980 7.330 7.410 ;
        RECT 7.390 6.980 9.000 7.410 ;
        RECT 10.550 6.980 16.580 7.410 ;
        RECT 0.890 6.450 2.500 6.980 ;
        RECT 0.890 5.020 6.530 6.450 ;
        RECT 6.590 5.020 8.200 6.450 ;
        RECT 9.220 5.240 14.580 6.450 ;
        RECT 9.750 5.020 14.580 5.240 ;
        RECT 0.890 4.950 14.580 5.020 ;
        RECT 0.890 3.140 6.530 4.950 ;
        RECT 1.700 2.610 6.530 3.140 ;
        RECT 0.090 1.760 6.530 2.610 ;
        RECT 6.590 1.760 8.200 4.950 ;
        RECT 9.750 4.710 14.580 4.950 ;
        RECT 8.420 2.610 14.580 4.710 ;
        RECT 15.380 3.140 16.580 6.980 ;
        RECT 8.420 2.540 16.190 2.610 ;
        RECT 9.210 2.480 16.190 2.540 ;
        RECT 9.750 1.830 16.190 2.480 ;
        RECT 8.420 1.760 16.190 1.830 ;
        RECT 8.420 0.020 10.030 1.760 ;
      LAYER li1 ;
        RECT 6.890 6.190 7.100 6.200 ;
        RECT 0.370 5.720 0.580 6.150 ;
        RECT 2.080 5.760 2.290 6.190 ;
        RECT 2.760 5.860 2.930 6.190 ;
        RECT 3.690 5.860 3.860 6.190 ;
        RECT 4.370 5.860 4.540 6.190 ;
        RECT 5.280 5.760 5.490 6.190 ;
        RECT 5.980 5.860 6.150 6.190 ;
        RECT 6.890 5.860 7.140 6.190 ;
        RECT 7.650 5.860 7.820 6.190 ;
        RECT 6.890 5.770 7.100 5.860 ;
        RECT 2.100 5.740 2.270 5.760 ;
        RECT 5.300 5.740 5.470 5.760 ;
        RECT 6.910 5.750 7.080 5.770 ;
        RECT 8.510 5.760 8.720 6.190 ;
        RECT 10.120 5.770 10.330 6.200 ;
        RECT 10.810 5.860 10.980 6.190 ;
        RECT 11.730 5.770 11.940 6.200 ;
        RECT 12.420 5.860 12.590 6.190 ;
        RECT 12.980 5.900 13.300 5.940 ;
        RECT 12.980 5.800 13.310 5.900 ;
        RECT 13.350 5.860 13.520 6.190 ;
        RECT 13.650 5.900 13.970 5.940 ;
        RECT 8.530 5.740 8.700 5.760 ;
        RECT 10.140 5.750 10.310 5.770 ;
        RECT 11.750 5.750 11.920 5.770 ;
        RECT 0.390 5.700 0.560 5.720 ;
        RECT 12.950 5.710 13.310 5.800 ;
        RECT 13.650 5.710 13.980 5.900 ;
        RECT 14.030 5.860 14.200 6.190 ;
        RECT 12.950 5.680 13.300 5.710 ;
        RECT 13.650 5.700 13.970 5.710 ;
        RECT 13.620 5.680 13.970 5.700 ;
        RECT 3.600 5.400 4.030 5.420 ;
        RECT 3.580 5.230 4.030 5.400 ;
        RECT 2.080 4.900 2.250 5.230 ;
        RECT 2.760 5.020 2.930 5.230 ;
        RECT 3.600 5.210 4.030 5.230 ;
        RECT 3.690 5.020 3.860 5.210 ;
        RECT 3.980 5.020 4.150 5.030 ;
        RECT 4.370 5.020 4.540 5.230 ;
        RECT 5.300 5.020 5.470 5.230 ;
        RECT 5.980 5.020 6.150 5.230 ;
        RECT 6.590 5.210 6.800 5.640 ;
        RECT 6.610 5.190 6.780 5.210 ;
        RECT 6.970 5.020 7.140 5.230 ;
        RECT 7.650 5.020 7.820 5.230 ;
        RECT 10.130 5.020 10.300 5.230 ;
        RECT 10.810 5.020 10.980 5.230 ;
        RECT 11.740 5.020 11.910 5.230 ;
        RECT 12.420 5.020 12.590 5.230 ;
        RECT 12.950 5.020 13.160 5.680 ;
        RECT 13.350 5.020 13.520 5.230 ;
        RECT 13.620 5.020 13.790 5.680 ;
        RECT 0.350 4.410 0.560 4.840 ;
        RECT 2.370 4.790 13.800 5.020 ;
        RECT 14.030 4.900 14.200 5.230 ;
        RECT 0.370 4.390 0.540 4.410 ;
        RECT 2.080 3.940 2.250 4.270 ;
        RECT 0.370 3.460 0.580 3.890 ;
        RECT 0.390 3.440 0.560 3.460 ;
        RECT 2.080 2.980 2.250 3.310 ;
        RECT 0.370 2.520 0.580 2.950 ;
        RECT 0.390 2.500 0.560 2.520 ;
        RECT 2.370 1.230 2.540 4.790 ;
        RECT 2.760 3.940 2.930 4.270 ;
        RECT 2.760 2.980 2.930 3.310 ;
        RECT 3.030 0.330 3.200 4.460 ;
        RECT 3.690 3.940 3.860 4.270 ;
        RECT 3.690 2.980 3.860 3.310 ;
        RECT 3.980 1.230 4.150 4.790 ;
        RECT 4.370 3.940 4.540 4.270 ;
        RECT 4.370 2.980 4.540 3.310 ;
        RECT 4.660 0.330 4.830 4.420 ;
        RECT 5.300 3.940 5.470 4.270 ;
        RECT 5.300 2.980 5.470 3.310 ;
        RECT 5.570 1.230 5.740 4.790 ;
        RECT 5.980 3.940 6.150 4.270 ;
        RECT 5.980 2.980 6.150 3.310 ;
        RECT 6.260 0.330 6.430 4.500 ;
        RECT 6.970 3.940 7.140 4.270 ;
        RECT 6.970 2.980 7.140 3.310 ;
        RECT 7.190 1.230 7.360 4.790 ;
        RECT 8.810 4.450 8.980 4.790 ;
        RECT 7.650 3.940 7.820 4.270 ;
        RECT 7.650 2.980 7.820 3.310 ;
        RECT 7.880 0.330 8.050 4.450 ;
        RECT 8.190 4.210 8.360 4.230 ;
        RECT 8.170 3.780 8.380 4.210 ;
        RECT 8.800 4.120 8.980 4.450 ;
        RECT 8.810 3.490 8.980 4.120 ;
        RECT 8.800 3.160 8.980 3.490 ;
        RECT 8.810 1.570 8.980 3.160 ;
        RECT 8.800 1.250 8.980 1.570 ;
        RECT 8.800 1.240 8.970 1.250 ;
        RECT 9.480 0.330 9.650 4.500 ;
        RECT 10.130 3.940 10.300 4.270 ;
        RECT 10.130 2.980 10.300 3.310 ;
        RECT 10.410 1.260 10.580 4.790 ;
        RECT 10.810 3.940 10.980 4.270 ;
        RECT 10.810 2.980 10.980 3.310 ;
        RECT 10.820 2.460 11.030 2.890 ;
        RECT 10.840 2.440 11.010 2.460 ;
        RECT 11.100 0.330 11.270 4.500 ;
        RECT 11.740 3.940 11.910 4.270 ;
        RECT 11.740 2.980 11.910 3.310 ;
        RECT 12.020 1.250 12.190 4.790 ;
        RECT 12.420 3.940 12.590 4.270 ;
        RECT 12.420 2.980 12.590 3.310 ;
        RECT 12.700 0.330 12.870 4.480 ;
        RECT 13.350 3.940 13.520 4.270 ;
        RECT 13.350 2.980 13.520 3.310 ;
        RECT 13.630 1.220 13.800 4.790 ;
        RECT 14.030 3.940 14.200 4.270 ;
        RECT 14.030 2.980 14.200 3.310 ;
        RECT 14.310 0.330 14.480 4.660 ;
        RECT 3.030 0.100 3.320 0.330 ;
        RECT 4.660 0.100 4.940 0.330 ;
        RECT 6.260 0.100 6.540 0.330 ;
        RECT 7.880 0.100 8.160 0.330 ;
        RECT 9.480 0.100 9.760 0.330 ;
        RECT 11.100 0.100 11.380 0.330 ;
        RECT 12.700 0.100 12.980 0.330 ;
        RECT 14.310 0.100 14.590 0.330 ;
        RECT 3.030 0.000 3.200 0.100 ;
        RECT 4.660 0.000 4.830 0.100 ;
        RECT 6.260 0.000 6.430 0.100 ;
        RECT 7.880 0.000 8.050 0.100 ;
        RECT 9.480 0.000 9.650 0.100 ;
        RECT 11.100 0.000 11.270 0.100 ;
        RECT 12.700 0.000 12.870 0.100 ;
        RECT 14.310 0.000 14.480 0.100 ;
      LAYER mcon ;
        RECT 13.040 5.720 13.210 5.890 ;
        RECT 13.710 5.720 13.880 5.890 ;
        RECT 8.190 4.060 8.360 4.230 ;
        RECT 3.140 0.130 3.310 0.300 ;
        RECT 4.760 0.130 4.930 0.300 ;
        RECT 6.360 0.130 6.530 0.300 ;
        RECT 7.980 0.130 8.150 0.300 ;
        RECT 9.580 0.130 9.750 0.300 ;
        RECT 11.200 0.130 11.370 0.300 ;
        RECT 12.800 0.130 12.970 0.300 ;
        RECT 14.410 0.130 14.580 0.300 ;
      LAYER met1 ;
        RECT 0.320 5.870 0.640 6.190 ;
        RECT 5.230 5.910 5.550 6.230 ;
        RECT 6.840 5.920 7.160 6.240 ;
        RECT 0.360 5.640 0.590 5.870 ;
        RECT 5.270 5.680 5.500 5.910 ;
        RECT 6.880 5.690 7.110 5.920 ;
        RECT 8.460 5.910 8.780 6.230 ;
        RECT 10.070 5.920 10.390 6.240 ;
        RECT 11.680 5.920 12.000 6.240 ;
        RECT 8.500 5.680 8.730 5.910 ;
        RECT 10.110 5.690 10.340 5.920 ;
        RECT 11.720 5.690 11.950 5.920 ;
        RECT 6.590 5.420 6.810 5.640 ;
        RECT 6.580 5.130 6.810 5.420 ;
        RECT 0.300 4.560 0.620 4.880 ;
        RECT 0.340 4.330 0.570 4.560 ;
        RECT 8.160 4.000 8.390 4.290 ;
        RECT 0.320 3.610 0.640 3.930 ;
        RECT 8.170 3.780 8.390 4.000 ;
        RECT 0.360 3.380 0.590 3.610 ;
        RECT 6.740 3.550 10.190 3.720 ;
        RECT 0.320 2.670 0.640 2.990 ;
        RECT 0.360 2.440 0.590 2.670 ;
        RECT 8.290 1.140 8.470 2.560 ;
        RECT 9.990 1.710 10.190 3.550 ;
        RECT 10.820 2.670 11.040 2.890 ;
        RECT 10.810 2.380 11.040 2.670 ;
        RECT 8.290 1.020 8.640 1.140 ;
        RECT 8.380 0.820 8.640 1.020 ;
      LAYER via ;
        RECT 0.350 5.900 0.610 6.160 ;
        RECT 5.260 5.940 5.520 6.200 ;
        RECT 6.870 5.950 7.130 6.210 ;
        RECT 8.490 5.940 8.750 6.200 ;
        RECT 10.100 5.950 10.360 6.210 ;
        RECT 11.710 5.950 11.970 6.210 ;
        RECT 0.330 4.590 0.590 4.850 ;
        RECT 0.350 3.640 0.610 3.900 ;
        RECT 0.350 2.700 0.610 2.960 ;
        RECT 8.380 0.850 8.640 1.110 ;
      LAYER met2 ;
        RECT 8.460 5.910 8.780 6.230 ;
        RECT 10.070 5.920 10.390 6.240 ;
        RECT 11.680 5.920 12.000 6.240 ;
        RECT 0.320 3.610 0.640 3.930 ;
  END
END sky130_hilas_DAC5bit01

MACRO sky130_hilas_capacitorSize04
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize04 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.170 BY 7.320 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAP1TERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 4.960 3.700 5.620 4.360 ;
    END
  END CAP1TERM02
  PIN CAP2TERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 4.960 0.700 5.620 1.360 ;
    END
  END CAP2TERM02
  PIN CAP2TERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 0.120 1.100 0.780 1.360 ;
        RECT 0.120 0.700 2.690 1.100 ;
        RECT 0.570 0.690 2.690 0.700 ;
    END
  END CAP2TERM01
  PIN CAP1TERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 0.090 4.110 0.750 4.360 ;
        RECT 0.090 3.700 3.050 4.110 ;
    END
  END CAP1TERM01
  OBS
      LAYER met2 ;
        RECT 0.020 4.850 5.770 5.030 ;
        RECT 0.020 4.420 5.770 4.600 ;
        RECT 0.220 4.180 0.590 4.240 ;
        RECT 0.020 3.900 0.590 4.180 ;
        RECT 0.220 3.840 0.590 3.900 ;
        RECT 5.090 4.180 5.460 4.240 ;
        RECT 5.090 3.900 5.770 4.180 ;
        RECT 5.090 3.840 5.460 3.900 ;
        RECT 0.020 3.420 5.770 3.600 ;
        RECT 0.020 2.990 5.770 3.170 ;
        RECT 0.020 1.840 5.770 2.010 ;
        RECT 0.020 1.420 5.770 1.590 ;
        RECT 0.250 1.180 0.620 1.240 ;
        RECT 0.020 0.900 0.620 1.180 ;
        RECT 0.250 0.840 0.620 0.900 ;
        RECT 5.090 1.180 5.460 1.240 ;
        RECT 5.090 0.900 5.780 1.180 ;
        RECT 5.090 0.840 5.460 0.900 ;
        RECT 0.020 0.440 5.770 0.610 ;
        RECT 0.020 0.000 5.770 0.170 ;
      LAYER via2 ;
        RECT 0.270 3.900 0.550 4.180 ;
        RECT 5.140 3.900 5.420 4.180 ;
        RECT 0.300 0.900 0.580 1.180 ;
        RECT 5.140 0.900 5.420 1.180 ;
      LAYER met3 ;
        RECT 5.870 5.040 8.170 7.320 ;
        RECT 0.000 3.640 0.790 4.390 ;
        RECT 3.860 3.640 5.660 4.390 ;
        RECT 5.870 2.030 8.170 4.310 ;
        RECT 0.030 0.640 0.820 1.390 ;
        RECT 4.870 1.380 5.660 1.390 ;
        RECT 3.850 0.650 5.660 1.380 ;
        RECT 4.870 0.640 5.660 0.650 ;
      LAYER via3 ;
        RECT 0.190 3.790 0.620 4.270 ;
        RECT 5.060 3.790 5.490 4.270 ;
        RECT 0.220 0.790 0.650 1.270 ;
        RECT 5.060 0.790 5.490 1.270 ;
      LAYER met4 ;
        RECT 6.720 6.270 7.170 6.280 ;
        RECT 6.700 5.780 7.220 6.270 ;
        RECT 6.720 3.260 7.170 3.270 ;
        RECT 6.700 2.770 7.220 3.260 ;
  END
END sky130_hilas_capacitorSize04

MACRO sky130_hilas_capacitorArray01
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorArray01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.700 BY 10.490 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM2
    USE ANALOG ;
    PORT
      LAYER met3 ;
        RECT 35.230 2.420 36.380 4.060 ;
        RECT 35.680 2.410 36.380 2.420 ;
    END
  END CAPTERM2
  PIN CAPTERM1
    USE ANALOG ;
    ANTENNAGATEAREA 0.720000 ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met3 ;
        RECT 11.250 5.960 11.630 6.250 ;
        RECT 11.170 4.710 11.710 5.960 ;
    END
  END CAPTERM1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 7.520 6.270 10.080 6.500 ;
        RECT 14.520 6.270 16.250 10.490 ;
        RECT 7.520 0.230 35.420 6.270 ;
        RECT 7.520 0.000 10.080 0.230 ;
        RECT 12.000 0.220 35.420 0.230 ;
      LAYER met1 ;
        RECT 9.560 5.790 9.720 6.490 ;
        RECT 9.450 5.240 9.720 5.790 ;
        RECT 9.450 5.190 9.730 5.240 ;
        RECT 9.560 5.100 9.730 5.190 ;
        RECT 9.560 4.630 9.720 5.100 ;
        RECT 9.560 4.540 9.730 4.630 ;
        RECT 9.450 4.490 9.730 4.540 ;
        RECT 9.450 3.940 9.720 4.490 ;
        RECT 9.560 2.550 9.720 3.940 ;
        RECT 9.450 2.000 9.720 2.550 ;
        RECT 9.450 1.950 9.730 2.000 ;
        RECT 9.560 1.860 9.730 1.950 ;
        RECT 9.560 1.400 9.720 1.860 ;
        RECT 9.560 1.310 9.730 1.400 ;
        RECT 9.450 1.260 9.730 1.310 ;
        RECT 9.450 0.710 9.720 1.260 ;
        RECT 9.560 0.010 9.720 0.710 ;
    END
  END VINJ
  PIN GATESELECT
    ANTENNAGATEAREA 0.720000 ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met2 ;
        RECT 10.740 6.240 11.250 6.270 ;
        RECT 8.670 6.150 8.990 6.220 ;
        RECT 10.740 6.150 11.670 6.240 ;
        RECT 8.670 5.960 11.670 6.150 ;
        RECT 11.170 5.940 11.670 5.960 ;
      LAYER via2 ;
        RECT 11.300 5.940 11.580 6.220 ;
    END
  END GATESELECT
  PIN VTUN
    ANTENNADIFFAREA 0.436600 ;
    PORT
      LAYER nwell ;
        RECT 0.010 3.910 1.740 4.410 ;
        RECT 0.000 3.730 1.740 3.910 ;
        RECT 0.010 2.570 1.740 3.730 ;
      LAYER met1 ;
        RECT 0.360 0.000 0.760 6.500 ;
    END
  END VTUN
  PIN GATE
    USE ANALOG ;
    ANTENNADIFFAREA 3.253900 ;
    PORT
      LAYER nwell ;
        RECT 3.760 0.000 5.990 6.490 ;
      LAYER met1 ;
        RECT 4.410 4.350 4.790 6.500 ;
        RECT 4.400 2.490 4.790 4.350 ;
        RECT 4.410 0.370 4.790 2.490 ;
        RECT 4.400 0.220 4.790 0.370 ;
        RECT 4.410 0.000 4.790 0.220 ;
    END
  END GATE
  PIN DRAIN2
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 7.610 3.970 7.920 3.980 ;
        RECT 0.010 3.910 10.080 3.970 ;
        RECT 35.690 3.910 36.700 3.920 ;
        RECT 0.000 3.790 36.700 3.910 ;
        RECT 0.000 3.730 0.120 3.790 ;
        RECT 7.610 3.650 7.920 3.790 ;
        RECT 8.940 3.730 36.700 3.790 ;
    END
  END DRAIN2
  PIN DRAIN1
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 7.610 5.940 7.920 6.080 ;
        RECT 0.010 5.770 10.080 5.940 ;
        RECT 0.010 5.760 36.700 5.770 ;
        RECT 0.010 5.590 0.120 5.760 ;
        RECT 7.610 5.750 7.920 5.760 ;
        RECT 8.980 5.590 36.700 5.760 ;
    END
  END DRAIN1
  PIN DRAIN4
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 0.020 0.740 0.120 0.910 ;
        RECT 7.610 0.740 7.920 0.750 ;
        RECT 8.810 0.740 36.700 0.910 ;
        RECT 0.010 0.570 10.080 0.740 ;
        RECT 7.610 0.560 10.080 0.570 ;
        RECT 7.610 0.420 7.920 0.560 ;
    END
  END DRAIN4
  PIN DRAIN3
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 0.020 2.700 0.120 2.750 ;
        RECT 7.610 2.700 7.920 2.840 ;
        RECT 8.770 2.700 36.700 2.750 ;
        RECT 0.010 2.580 36.700 2.700 ;
        RECT 0.010 2.520 10.080 2.580 ;
        RECT 7.610 2.510 7.920 2.520 ;
    END
  END DRAIN3
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 2.760 1.780 3.080 1.790 ;
        RECT 6.690 1.780 7.010 1.840 ;
        RECT 2.760 1.600 7.010 1.780 ;
        RECT 2.760 1.530 3.080 1.600 ;
        RECT 6.690 1.550 7.010 1.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.730 5.110 6.970 6.500 ;
        RECT 6.710 4.450 6.980 5.110 ;
        RECT 6.730 1.860 6.970 4.450 ;
        RECT 6.720 1.540 6.980 1.860 ;
        RECT 6.730 0.000 6.970 1.540 ;
      LAYER via ;
        RECT 6.720 1.570 6.980 1.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.800 5.090 3.040 6.500 ;
        RECT 2.790 4.430 3.050 5.090 ;
        RECT 2.800 1.820 3.040 4.430 ;
        RECT 2.790 1.500 3.050 1.820 ;
        RECT 2.800 0.000 3.040 1.500 ;
      LAYER via ;
        RECT 2.790 1.530 3.050 1.790 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 0.010 5.590 0.120 5.770 ;
        RECT 0.010 5.160 0.080 5.340 ;
        RECT 0.580 4.810 1.170 4.920 ;
        RECT 0.580 1.530 1.170 1.720 ;
        RECT 0.020 0.740 0.120 0.910 ;
      LAYER li1 ;
        RECT 7.620 6.030 7.940 6.040 ;
        RECT 7.620 5.860 8.200 6.030 ;
        RECT 7.620 5.810 7.950 5.860 ;
        RECT 7.620 5.780 7.940 5.810 ;
        RECT 9.480 5.760 9.680 6.110 ;
        RECT 7.620 5.450 7.940 5.490 ;
        RECT 7.620 5.410 7.950 5.450 ;
        RECT 7.620 5.240 8.200 5.410 ;
        RECT 7.620 5.230 7.940 5.240 ;
        RECT 8.750 5.140 8.950 5.740 ;
        RECT 9.480 5.730 9.690 5.760 ;
        RECT 9.470 5.140 9.690 5.730 ;
        RECT 2.830 4.520 3.000 5.050 ;
        RECT 6.770 4.510 6.940 5.040 ;
        RECT 7.620 4.490 7.940 4.500 ;
        RECT 7.620 4.320 8.200 4.490 ;
        RECT 7.620 4.280 7.950 4.320 ;
        RECT 7.620 4.240 7.940 4.280 ;
        RECT 8.750 3.990 8.950 4.590 ;
        RECT 9.470 4.000 9.690 4.590 ;
        RECT 9.480 3.970 9.690 4.000 ;
        RECT 7.620 3.920 7.940 3.950 ;
        RECT 7.620 3.870 7.950 3.920 ;
        RECT 0.430 3.020 0.980 3.450 ;
        RECT 2.840 2.810 3.010 3.820 ;
        RECT 7.620 3.700 8.200 3.870 ;
        RECT 7.620 3.690 7.940 3.700 ;
        RECT 4.460 2.950 5.010 3.380 ;
        RECT 6.770 2.670 6.940 3.680 ;
        RECT 9.480 3.620 9.680 3.970 ;
        RECT 8.870 3.160 9.310 3.330 ;
        RECT 7.620 2.790 7.940 2.800 ;
        RECT 7.620 2.620 8.200 2.790 ;
        RECT 7.620 2.570 7.950 2.620 ;
        RECT 7.620 2.540 7.940 2.570 ;
        RECT 9.480 2.520 9.680 2.870 ;
        RECT 7.620 2.210 7.940 2.250 ;
        RECT 7.620 2.170 7.950 2.210 ;
        RECT 7.620 2.000 8.200 2.170 ;
        RECT 7.620 1.990 7.940 2.000 ;
        RECT 8.750 1.900 8.950 2.500 ;
        RECT 9.480 2.490 9.690 2.520 ;
        RECT 9.470 1.900 9.690 2.490 ;
        RECT 7.620 1.260 7.940 1.270 ;
        RECT 7.620 1.090 8.200 1.260 ;
        RECT 7.620 1.050 7.950 1.090 ;
        RECT 7.620 1.010 7.940 1.050 ;
        RECT 8.750 0.760 8.950 1.360 ;
        RECT 9.470 0.770 9.690 1.360 ;
        RECT 9.480 0.740 9.690 0.770 ;
        RECT 7.620 0.690 7.940 0.720 ;
        RECT 7.620 0.640 7.950 0.690 ;
        RECT 7.620 0.470 8.200 0.640 ;
        RECT 7.620 0.460 7.940 0.470 ;
        RECT 9.480 0.390 9.680 0.740 ;
      LAYER mcon ;
        RECT 7.680 5.820 7.850 5.990 ;
        RECT 8.760 5.530 8.930 5.700 ;
        RECT 7.680 5.270 7.850 5.440 ;
        RECT 9.490 5.560 9.660 5.730 ;
        RECT 2.830 4.880 3.000 5.050 ;
        RECT 6.770 4.870 6.940 5.040 ;
        RECT 7.680 4.290 7.850 4.460 ;
        RECT 8.760 4.030 8.930 4.200 ;
        RECT 9.490 4.000 9.660 4.170 ;
        RECT 7.680 3.740 7.850 3.910 ;
        RECT 0.430 3.100 0.700 3.370 ;
        RECT 2.840 3.420 3.010 3.590 ;
        RECT 2.840 3.060 3.010 3.230 ;
        RECT 4.460 3.030 4.730 3.300 ;
        RECT 6.770 3.280 6.940 3.450 ;
        RECT 9.130 3.160 9.310 3.330 ;
        RECT 6.770 2.920 6.940 3.090 ;
        RECT 7.680 2.580 7.850 2.750 ;
        RECT 8.760 2.290 8.930 2.460 ;
        RECT 7.680 2.030 7.850 2.200 ;
        RECT 9.490 2.320 9.660 2.490 ;
        RECT 7.680 1.060 7.850 1.230 ;
        RECT 8.760 0.800 8.930 0.970 ;
        RECT 9.490 0.770 9.660 0.940 ;
        RECT 7.680 0.510 7.850 0.680 ;
      LAYER met1 ;
        RECT 8.750 6.250 8.910 6.490 ;
        RECT 7.610 5.750 7.930 6.070 ;
        RECT 8.700 5.930 8.960 6.250 ;
        RECT 8.750 5.760 8.910 5.930 ;
        RECT 8.750 5.740 8.950 5.760 ;
        RECT 7.610 5.200 7.930 5.520 ;
        RECT 8.730 5.500 8.960 5.740 ;
        RECT 8.750 5.450 8.960 5.500 ;
        RECT 9.120 5.450 9.310 6.440 ;
        RECT 7.610 4.210 7.930 4.530 ;
        RECT 8.750 4.280 8.910 5.450 ;
        RECT 9.140 5.330 9.310 5.450 ;
        RECT 9.150 4.400 9.310 5.330 ;
        RECT 9.140 4.280 9.310 4.400 ;
        RECT 8.750 4.230 8.960 4.280 ;
        RECT 8.730 3.990 8.960 4.230 ;
        RECT 7.610 3.660 7.930 3.980 ;
        RECT 8.750 3.970 8.950 3.990 ;
        RECT 8.750 3.340 8.910 3.970 ;
        RECT 9.120 3.360 9.310 4.280 ;
        RECT 9.100 3.340 9.340 3.360 ;
        RECT 8.750 3.150 9.340 3.340 ;
        RECT 7.610 2.510 7.930 2.830 ;
        RECT 8.750 2.520 8.910 3.150 ;
        RECT 9.100 3.130 9.340 3.150 ;
        RECT 8.750 2.500 8.950 2.520 ;
        RECT 7.610 1.960 7.930 2.280 ;
        RECT 8.730 2.260 8.960 2.500 ;
        RECT 8.750 2.210 8.960 2.260 ;
        RECT 9.120 2.210 9.310 3.130 ;
        RECT 7.610 0.980 7.930 1.300 ;
        RECT 8.750 1.050 8.910 2.210 ;
        RECT 9.140 2.090 9.310 2.210 ;
        RECT 9.150 1.170 9.310 2.090 ;
        RECT 9.140 1.050 9.310 1.170 ;
        RECT 8.750 1.000 8.960 1.050 ;
        RECT 8.730 0.760 8.960 1.000 ;
        RECT 7.610 0.430 7.930 0.750 ;
        RECT 8.750 0.740 8.950 0.760 ;
        RECT 8.750 0.010 8.910 0.740 ;
        RECT 9.120 0.060 9.310 1.050 ;
      LAYER via ;
        RECT 7.640 5.780 7.900 6.040 ;
        RECT 8.700 5.960 8.960 6.220 ;
        RECT 7.640 5.230 7.900 5.490 ;
        RECT 7.640 4.240 7.900 4.500 ;
        RECT 7.640 3.690 7.900 3.950 ;
        RECT 7.640 2.540 7.900 2.800 ;
        RECT 7.640 1.990 7.900 2.250 ;
        RECT 7.640 1.010 7.900 1.270 ;
        RECT 7.640 0.460 7.900 0.720 ;
      LAYER met2 ;
        RECT 7.610 5.510 7.920 5.530 ;
        RECT 7.520 5.500 10.080 5.510 ;
        RECT 0.010 5.340 10.080 5.500 ;
        RECT 0.010 5.330 36.700 5.340 ;
        RECT 0.010 5.320 7.920 5.330 ;
        RECT 7.610 5.200 7.920 5.320 ;
        RECT 8.920 5.160 36.700 5.330 ;
        RECT 7.610 4.400 7.920 4.530 ;
        RECT 9.880 4.400 10.250 4.510 ;
        RECT 0.010 4.340 10.250 4.400 ;
        RECT 0.010 4.220 36.700 4.340 ;
        RECT 7.610 4.200 7.920 4.220 ;
        RECT 8.980 4.160 36.700 4.220 ;
        RECT 9.880 4.110 10.250 4.160 ;
        RECT 36.010 3.010 36.700 3.420 ;
        RECT 9.840 2.330 10.210 2.420 ;
        RECT 7.610 2.270 7.920 2.290 ;
        RECT 8.870 2.270 36.700 2.330 ;
        RECT 0.010 2.160 36.700 2.270 ;
        RECT 0.010 2.090 10.210 2.160 ;
        RECT 7.610 1.960 7.920 2.090 ;
        RECT 9.840 2.020 10.210 2.090 ;
        RECT 10.930 1.350 11.300 1.550 ;
        RECT 7.610 1.170 7.920 1.300 ;
        RECT 8.850 1.180 36.700 1.350 ;
        RECT 0.010 0.990 10.080 1.170 ;
        RECT 10.930 1.150 11.300 1.180 ;
        RECT 7.610 0.970 7.920 0.990 ;
      LAYER via2 ;
        RECT 9.930 4.170 10.210 4.450 ;
        RECT 36.080 3.070 36.370 3.350 ;
        RECT 9.890 2.080 10.170 2.360 ;
        RECT 10.980 1.210 11.260 1.490 ;
      LAYER met3 ;
        RECT 9.660 3.910 10.450 4.660 ;
        RECT 9.620 2.520 10.410 2.570 ;
        RECT 9.620 2.220 10.550 2.520 ;
        RECT 9.620 1.820 10.410 2.220 ;
        RECT 10.710 1.310 11.500 1.700 ;
        RECT 10.710 1.010 11.640 1.310 ;
        RECT 10.710 0.950 11.500 1.010 ;
      LAYER via3 ;
        RECT 9.850 4.060 10.280 4.540 ;
        RECT 9.810 1.970 10.240 2.450 ;
        RECT 10.900 1.100 11.330 1.580 ;
      LAYER met4 ;
        RECT 12.790 5.600 16.890 5.900 ;
        RECT 11.100 4.990 13.800 5.100 ;
        RECT 11.100 4.690 14.010 4.990 ;
        RECT 9.750 4.270 10.410 4.630 ;
        RECT 13.500 4.350 14.010 4.690 ;
        RECT 16.510 4.400 16.890 5.600 ;
        RECT 19.350 4.430 22.630 4.730 ;
        RECT 9.750 3.970 11.770 4.270 ;
        RECT 11.470 3.410 11.770 3.970 ;
        RECT 19.350 3.410 19.650 4.430 ;
        RECT 22.330 3.410 22.630 4.430 ;
        RECT 11.470 3.110 22.630 3.410 ;
        RECT 25.030 4.410 33.920 4.710 ;
        RECT 9.710 2.520 10.370 2.540 ;
        RECT 13.710 2.520 16.900 2.550 ;
        RECT 19.350 2.520 19.650 2.550 ;
        RECT 9.710 2.220 22.570 2.520 ;
        RECT 9.710 1.880 10.370 2.220 ;
        RECT 13.710 1.850 14.010 2.220 ;
        RECT 16.600 1.880 16.900 2.220 ;
        RECT 19.350 1.880 19.650 2.220 ;
        RECT 16.600 1.850 19.650 1.880 ;
        RECT 22.270 1.850 22.570 2.220 ;
        RECT 10.800 1.310 11.460 1.670 ;
        RECT 13.710 1.550 22.570 1.850 ;
        RECT 25.030 1.890 25.330 4.410 ;
        RECT 27.860 4.380 30.970 4.410 ;
        RECT 27.860 1.890 28.160 4.380 ;
        RECT 30.670 1.890 30.970 4.380 ;
        RECT 33.620 1.890 33.920 4.410 ;
        RECT 25.030 1.590 33.980 1.890 ;
        RECT 30.670 1.580 33.980 1.590 ;
        RECT 10.800 1.010 11.850 1.310 ;
        RECT 11.550 0.770 11.850 1.010 ;
        RECT 33.680 0.770 33.980 1.580 ;
        RECT 11.550 0.470 33.980 0.770 ;
  END
END sky130_hilas_capacitorArray01

MACRO sky130_hilas_pFETmed
  CLASS CORE ;
  FOREIGN sky130_hilas_pFETmed ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.190 BY 2.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 0.000 0.000 1.190 2.870 ;
      LAYER li1 ;
        RECT 0.240 0.150 0.410 2.640 ;
        RECT 0.790 0.140 0.960 2.640 ;
  END
END sky130_hilas_pFETmed

MACRO sky130_hilas_swc4x1cellOverlap2
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x1cellOverlap2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.350 BY 6.160 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 6.790 0.000 9.350 6.160 ;
      LAYER li1 ;
        RECT 1.680 5.320 1.850 6.160 ;
        RECT 7.030 5.810 7.350 5.850 ;
        RECT 7.030 5.690 7.360 5.810 ;
        RECT 7.030 5.590 7.470 5.690 ;
        RECT 7.130 5.520 7.470 5.590 ;
        RECT 7.030 5.260 7.350 5.300 ;
        RECT 7.030 5.070 7.360 5.260 ;
        RECT 7.030 5.040 7.470 5.070 ;
        RECT 7.130 4.900 7.470 5.040 ;
        RECT 8.020 4.800 8.220 5.400 ;
        RECT 8.350 5.330 9.350 6.160 ;
        RECT 8.740 4.840 8.960 5.330 ;
        RECT 1.680 3.800 1.850 4.690 ;
        RECT 7.130 4.120 7.470 4.260 ;
        RECT 7.030 4.090 7.470 4.120 ;
        RECT 7.030 3.900 7.360 4.090 ;
        RECT 7.030 3.860 7.350 3.900 ;
        RECT 8.020 3.760 8.220 4.360 ;
        RECT 8.350 3.860 9.350 4.840 ;
        RECT 8.740 3.770 8.960 3.860 ;
        RECT 8.750 3.740 8.960 3.770 ;
        RECT 7.130 3.570 7.470 3.640 ;
        RECT 7.030 3.470 7.470 3.570 ;
        RECT 7.030 3.350 7.360 3.470 ;
        RECT 8.750 3.390 8.950 3.740 ;
        RECT 7.030 3.310 7.350 3.350 ;
        RECT 1.680 2.350 1.850 3.240 ;
        RECT 8.350 3.160 9.350 3.370 ;
        RECT 8.140 2.990 9.350 3.160 ;
        RECT 7.030 2.800 7.350 2.840 ;
        RECT 7.030 2.680 7.360 2.800 ;
        RECT 7.030 2.580 7.470 2.680 ;
        RECT 7.130 2.510 7.470 2.580 ;
        RECT 8.350 2.390 9.350 2.990 ;
        RECT 7.030 2.250 7.350 2.290 ;
        RECT 7.030 2.060 7.360 2.250 ;
        RECT 7.030 2.030 7.470 2.060 ;
        RECT 7.130 1.890 7.470 2.030 ;
        RECT 8.020 1.790 8.220 2.390 ;
        RECT 8.750 2.380 8.960 2.390 ;
        RECT 8.740 1.900 8.960 2.380 ;
        RECT 1.680 0.810 1.850 1.700 ;
        RECT 7.130 1.120 7.470 1.260 ;
        RECT 7.030 1.090 7.470 1.120 ;
        RECT 7.030 0.900 7.360 1.090 ;
        RECT 7.030 0.860 7.350 0.900 ;
        RECT 8.020 0.760 8.220 1.360 ;
        RECT 8.350 0.920 9.350 1.900 ;
        RECT 8.740 0.770 8.960 0.920 ;
        RECT 8.750 0.740 8.960 0.770 ;
        RECT 7.130 0.570 7.470 0.640 ;
        RECT 7.030 0.470 7.470 0.570 ;
        RECT 7.030 0.350 7.360 0.470 ;
        RECT 8.750 0.390 8.950 0.740 ;
        RECT 7.030 0.310 7.350 0.350 ;
      LAYER mcon ;
        RECT 1.680 6.010 1.850 6.160 ;
        RECT 7.090 5.630 7.260 5.800 ;
        RECT 7.090 5.080 7.260 5.250 ;
        RECT 8.030 5.190 8.200 5.360 ;
        RECT 8.760 5.220 8.930 5.390 ;
        RECT 1.680 4.490 1.850 4.660 ;
        RECT 7.090 3.910 7.260 4.080 ;
        RECT 8.030 3.800 8.200 3.970 ;
        RECT 8.760 3.770 8.930 3.940 ;
        RECT 7.090 3.360 7.260 3.530 ;
        RECT 1.680 3.040 1.850 3.210 ;
        RECT 8.400 2.990 8.580 3.160 ;
        RECT 7.090 2.620 7.260 2.790 ;
        RECT 7.090 2.070 7.260 2.240 ;
        RECT 8.030 2.180 8.200 2.350 ;
        RECT 8.760 2.210 8.930 2.380 ;
        RECT 1.680 1.500 1.850 1.670 ;
        RECT 7.090 0.910 7.260 1.080 ;
        RECT 8.030 0.800 8.200 0.970 ;
        RECT 8.760 0.770 8.930 0.940 ;
        RECT 7.090 0.360 7.260 0.530 ;
      LAYER met1 ;
        RECT 1.010 0.050 1.280 6.100 ;
        RECT 1.650 5.110 1.880 6.160 ;
        RECT 7.020 5.560 7.340 5.880 ;
        RECT 8.020 5.420 8.180 6.150 ;
        RECT 8.020 5.400 8.220 5.420 ;
        RECT 7.020 5.010 7.340 5.330 ;
        RECT 8.000 5.160 8.230 5.400 ;
        RECT 8.020 5.110 8.230 5.160 ;
        RECT 8.390 5.110 8.580 6.100 ;
        RECT 8.830 5.450 8.990 6.150 ;
        RECT 1.650 3.590 1.880 4.880 ;
        RECT 7.020 3.830 7.340 4.150 ;
        RECT 8.020 4.050 8.180 5.110 ;
        RECT 8.410 4.990 8.580 5.110 ;
        RECT 8.420 4.170 8.580 4.990 ;
        RECT 8.720 4.900 8.990 5.450 ;
        RECT 8.720 4.850 9.000 4.900 ;
        RECT 8.830 4.760 9.000 4.850 ;
        RECT 8.830 4.400 8.990 4.760 ;
        RECT 8.830 4.310 9.000 4.400 ;
        RECT 8.410 4.050 8.580 4.170 ;
        RECT 8.020 4.000 8.230 4.050 ;
        RECT 8.000 3.760 8.230 4.000 ;
        RECT 8.020 3.740 8.220 3.760 ;
        RECT 1.650 2.140 1.880 3.430 ;
        RECT 7.020 3.280 7.340 3.600 ;
        RECT 7.020 2.550 7.340 2.870 ;
        RECT 8.020 2.410 8.180 3.740 ;
        RECT 8.390 3.190 8.580 4.050 ;
        RECT 8.720 4.260 9.000 4.310 ;
        RECT 8.720 3.710 8.990 4.260 ;
        RECT 8.370 2.960 8.610 3.190 ;
        RECT 8.020 2.390 8.220 2.410 ;
        RECT 7.020 2.000 7.340 2.320 ;
        RECT 8.000 2.150 8.230 2.390 ;
        RECT 8.020 2.100 8.230 2.150 ;
        RECT 8.390 2.100 8.580 2.960 ;
        RECT 8.830 2.440 8.990 3.710 ;
        RECT 1.650 0.600 1.880 1.890 ;
        RECT 7.020 0.830 7.340 1.150 ;
        RECT 8.020 1.050 8.180 2.100 ;
        RECT 8.410 1.980 8.580 2.100 ;
        RECT 8.420 1.170 8.580 1.980 ;
        RECT 8.720 1.890 8.990 2.440 ;
        RECT 8.720 1.840 9.000 1.890 ;
        RECT 8.830 1.750 9.000 1.840 ;
        RECT 8.830 1.400 8.990 1.750 ;
        RECT 8.830 1.310 9.000 1.400 ;
        RECT 8.410 1.050 8.580 1.170 ;
        RECT 8.020 1.000 8.230 1.050 ;
        RECT 8.000 0.760 8.230 1.000 ;
        RECT 8.020 0.740 8.220 0.760 ;
        RECT 7.020 0.280 7.340 0.600 ;
        RECT 8.020 0.010 8.180 0.740 ;
        RECT 8.390 0.060 8.580 1.050 ;
        RECT 8.720 1.260 9.000 1.310 ;
        RECT 8.720 0.710 8.990 1.260 ;
        RECT 8.830 0.010 8.990 0.710 ;
      LAYER via ;
        RECT 7.050 5.590 7.310 5.850 ;
        RECT 7.050 5.040 7.310 5.300 ;
        RECT 7.050 3.860 7.310 4.120 ;
        RECT 7.050 3.310 7.310 3.570 ;
        RECT 7.050 2.580 7.310 2.840 ;
        RECT 7.050 2.030 7.310 2.290 ;
        RECT 7.050 0.860 7.310 1.120 ;
        RECT 7.050 0.310 7.310 0.570 ;
      LAYER met2 ;
        RECT 7.020 5.600 7.330 5.890 ;
        RECT 0.000 5.530 6.880 5.600 ;
        RECT 7.020 5.560 9.350 5.600 ;
        RECT 0.000 5.420 6.910 5.530 ;
        RECT 7.170 5.420 9.350 5.560 ;
        RECT 7.020 5.170 7.330 5.340 ;
        RECT 0.000 4.990 9.350 5.170 ;
        RECT 0.000 4.110 6.880 4.170 ;
        RECT 7.180 4.150 9.350 4.170 ;
        RECT 0.000 3.990 6.910 4.110 ;
        RECT 7.020 3.990 9.350 4.150 ;
        RECT 7.020 3.820 7.330 3.990 ;
        RECT 0.000 3.670 6.870 3.740 ;
        RECT 0.000 3.560 6.910 3.670 ;
        RECT 7.170 3.600 9.350 3.740 ;
        RECT 7.020 3.560 9.350 3.600 ;
        RECT 7.020 3.270 7.330 3.560 ;
        RECT 7.020 2.590 7.330 2.880 ;
        RECT 0.000 2.410 6.910 2.580 ;
        RECT 7.020 2.550 9.350 2.590 ;
        RECT 7.170 2.410 9.350 2.550 ;
        RECT 7.020 2.160 7.330 2.330 ;
        RECT 0.000 1.990 6.910 2.160 ;
        RECT 7.020 2.000 9.350 2.160 ;
        RECT 6.790 1.980 6.880 1.990 ;
        RECT 7.180 1.980 9.350 2.000 ;
        RECT 0.000 1.010 6.910 1.180 ;
        RECT 7.180 1.150 9.350 1.170 ;
        RECT 6.790 0.990 6.880 1.010 ;
        RECT 7.020 0.990 9.350 1.150 ;
        RECT 7.020 0.820 7.330 0.990 ;
        RECT 0.000 0.570 6.910 0.740 ;
        RECT 7.170 0.600 9.350 0.740 ;
        RECT 7.020 0.560 9.350 0.600 ;
        RECT 7.020 0.270 7.330 0.560 ;
  END
END sky130_hilas_swc4x1cellOverlap2

MACRO sky130_hilas_TA2SignalBiasCell
  CLASS CORE ;
  FOREIGN sky130_hilas_TA2SignalBiasCell ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.600 BY 6.360 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VOUT_AMP2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 8.730 3.480 8.880 3.700 ;
    END
  END VOUT_AMP2
  PIN VOUT_AMP1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 8.730 2.660 8.880 2.880 ;
    END
  END VOUT_AMP1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 6.920 0.140 7.260 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.920 6.050 7.260 6.190 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 7.590 0.140 7.860 0.350 ;
    END
    PORT
      LAYER met2 ;
        RECT 7.820 6.110 8.130 6.340 ;
        RECT 10.070 6.110 10.380 6.360 ;
        RECT 7.690 6.030 10.380 6.110 ;
        RECT 7.690 5.880 10.230 6.030 ;
    END
    PORT
      LAYER nwell ;
        RECT 4.060 6.190 7.670 6.360 ;
        RECT 0.000 6.180 1.910 6.190 ;
        RECT 4.060 6.180 8.880 6.190 ;
        RECT 0.000 6.010 8.880 6.180 ;
        RECT 0.000 4.590 7.670 6.010 ;
        RECT 0.000 0.580 5.600 4.590 ;
        RECT 0.000 0.400 0.430 0.580 ;
        RECT 0.000 0.170 0.710 0.400 ;
        RECT 0.000 0.150 0.430 0.170 ;
      LAYER met2 ;
        RECT 0.790 6.160 1.030 6.190 ;
        RECT 0.790 5.830 1.200 6.160 ;
        RECT 0.790 5.720 1.030 5.830 ;
        RECT 0.270 5.370 1.030 5.720 ;
        RECT 0.270 5.140 4.810 5.370 ;
        RECT 0.270 4.900 1.030 5.140 ;
        RECT 0.270 4.890 0.720 4.900 ;
        RECT 4.580 4.780 4.810 5.140 ;
        RECT 7.600 4.780 7.930 4.930 ;
        RECT 4.580 4.580 7.930 4.780 ;
        RECT 4.840 4.570 7.930 4.580 ;
        RECT 7.330 4.530 7.930 4.570 ;
        RECT 7.330 4.430 8.080 4.530 ;
        RECT 7.600 4.200 8.080 4.430 ;
        RECT 7.600 4.000 7.930 4.200 ;
        RECT 0.850 1.670 1.160 2.000 ;
    END
  END VPWR
  PIN VIN22
    USE ANALOG ;
    ANTENNAGATEAREA 0.626300 ;
    PORT
      LAYER met2 ;
        RECT 4.390 6.170 4.640 6.180 ;
        RECT 4.850 6.170 5.160 6.330 ;
        RECT 4.390 5.920 5.300 6.170 ;
    END
  END VIN22
  PIN VIN21
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.660 3.480 5.090 3.490 ;
        RECT 4.430 3.250 5.530 3.480 ;
        RECT 4.890 3.050 5.200 3.250 ;
    END
  END VIN21
  PIN VIN11
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 3.330 3.080 3.640 3.280 ;
        RECT 2.870 2.850 3.970 3.080 ;
        RECT 2.870 2.840 3.530 2.850 ;
    END
  END VIN11
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 2.830 0.160 3.740 0.410 ;
        RECT 3.290 0.000 3.600 0.160 ;
    END
  END VIN12
  PIN VBIAS2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.110 0.400 1.990 0.410 ;
        RECT 0.050 0.170 1.990 0.400 ;
        RECT 1.110 0.160 1.990 0.170 ;
        RECT 1.540 0.000 1.850 0.160 ;
    END
  END VBIAS2
  PIN VBIAS1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.580 3.080 1.890 3.280 ;
        RECT 0.010 2.850 2.220 3.080 ;
        RECT 0.010 2.840 1.780 2.850 ;
        RECT 0.010 2.830 0.650 2.840 ;
    END
  END VBIAS1
  OBS
      LAYER nwell ;
        RECT 7.370 0.000 9.230 1.740 ;
        RECT 9.320 0.590 10.600 6.270 ;
      LAYER li1 ;
        RECT 0.900 6.080 1.220 6.120 ;
        RECT 0.900 5.890 1.230 6.080 ;
        RECT 0.900 5.860 1.220 5.890 ;
        RECT 0.670 5.710 1.010 5.720 ;
        RECT 0.420 5.520 1.010 5.710 ;
        RECT 0.250 5.300 1.010 5.520 ;
        RECT 0.250 5.130 0.840 5.300 ;
        RECT 0.250 4.980 1.010 5.130 ;
        RECT 4.470 5.060 4.650 6.360 ;
        RECT 4.830 6.250 5.150 6.290 ;
        RECT 4.820 6.190 5.150 6.250 ;
        RECT 4.730 6.030 5.150 6.190 ;
        RECT 4.730 5.880 4.970 6.030 ;
        RECT 4.730 5.860 4.900 5.880 ;
        RECT 5.280 5.460 5.450 6.360 ;
        RECT 4.980 5.420 5.450 5.460 ;
        RECT 4.970 5.320 5.450 5.420 ;
        RECT 4.970 5.230 5.530 5.320 ;
        RECT 4.980 5.200 5.530 5.230 ;
        RECT 5.200 5.150 5.530 5.200 ;
        RECT 6.220 5.060 6.400 6.360 ;
        RECT 7.030 5.320 7.200 6.360 ;
        RECT 7.830 6.260 8.150 6.300 ;
        RECT 10.080 6.280 10.400 6.320 ;
        RECT 7.830 6.070 8.160 6.260 ;
        RECT 10.080 6.210 10.410 6.280 ;
        RECT 7.830 6.040 8.150 6.070 ;
        RECT 7.920 5.860 8.120 6.040 ;
        RECT 7.780 5.610 8.100 5.650 ;
        RECT 6.950 5.150 7.280 5.320 ;
        RECT 7.510 5.210 7.680 5.540 ;
        RECT 7.780 5.530 8.110 5.610 ;
        RECT 7.780 5.390 8.120 5.530 ;
        RECT 7.920 5.200 8.120 5.390 ;
        RECT 8.510 5.200 9.060 6.190 ;
        RECT 9.880 6.040 10.510 6.210 ;
        RECT 9.880 5.760 10.240 6.040 ;
        RECT 9.530 5.590 10.240 5.760 ;
        RECT 0.250 3.650 0.420 4.980 ;
        RECT 0.840 4.960 1.010 4.980 ;
        RECT 9.530 4.920 10.230 5.150 ;
        RECT 1.740 4.800 2.060 4.840 ;
        RECT 1.740 4.610 2.070 4.800 ;
        RECT 7.650 4.680 7.900 4.890 ;
        RECT 9.480 4.690 10.230 4.920 ;
        RECT 1.740 4.580 2.060 4.610 ;
        RECT 4.170 4.600 4.490 4.630 ;
        RECT 4.170 4.410 4.500 4.600 ;
        RECT 7.510 4.500 7.900 4.680 ;
        RECT 7.920 4.500 8.120 4.690 ;
        RECT 4.170 4.370 4.490 4.410 ;
        RECT 7.510 4.360 8.120 4.500 ;
        RECT 7.510 4.350 8.110 4.360 ;
        RECT 7.650 4.280 8.110 4.350 ;
        RECT 7.650 4.240 8.100 4.280 ;
        RECT 7.650 4.000 7.860 4.240 ;
        RECT 2.030 3.930 2.220 3.950 ;
        RECT 3.780 3.930 3.970 3.950 ;
        RECT 1.890 3.840 2.220 3.930 ;
        RECT 1.890 3.760 1.970 3.840 ;
        RECT 2.030 3.720 2.220 3.840 ;
        RECT 3.640 3.840 3.970 3.930 ;
        RECT 7.920 3.850 8.120 4.030 ;
        RECT 3.640 3.760 3.720 3.840 ;
        RECT 3.780 3.720 3.970 3.840 ;
        RECT 7.830 3.820 8.150 3.850 ;
        RECT 0.840 2.620 1.020 3.680 ;
        RECT 1.400 3.340 1.570 3.500 ;
        RECT 1.400 3.240 1.620 3.340 ;
        RECT 1.400 3.200 1.910 3.240 ;
        RECT 1.400 3.170 1.920 3.200 ;
        RECT 1.450 3.080 1.920 3.170 ;
        RECT 1.590 3.010 1.920 3.080 ;
        RECT 1.590 2.980 1.910 3.010 ;
        RECT 2.590 2.620 2.770 3.680 ;
        RECT 3.150 3.340 3.320 3.500 ;
        RECT 3.150 3.240 3.370 3.340 ;
        RECT 3.150 3.200 3.660 3.240 ;
        RECT 3.150 3.170 3.670 3.200 ;
        RECT 3.200 3.080 3.670 3.170 ;
        RECT 3.340 3.010 3.670 3.080 ;
        RECT 3.340 2.980 3.660 3.010 ;
        RECT 4.150 2.650 4.330 3.710 ;
        RECT 7.830 3.630 8.160 3.820 ;
        RECT 8.510 3.700 9.060 4.690 ;
        RECT 9.530 4.270 10.230 4.690 ;
        RECT 10.130 4.060 10.450 4.100 ;
        RECT 10.130 3.870 10.460 4.060 ;
        RECT 10.130 3.850 10.450 3.870 ;
        RECT 9.520 3.840 10.450 3.850 ;
        RECT 9.520 3.670 10.220 3.840 ;
        RECT 7.830 3.590 8.150 3.630 ;
        RECT 4.900 3.320 5.220 3.350 ;
        RECT 10.120 3.340 10.440 3.380 ;
        RECT 4.900 3.250 5.230 3.320 ;
        RECT 4.760 3.160 5.230 3.250 ;
        RECT 4.710 3.130 5.230 3.160 ;
        RECT 7.830 3.260 8.150 3.300 ;
        RECT 4.710 3.090 5.220 3.130 ;
        RECT 4.710 2.990 4.930 3.090 ;
        RECT 7.830 3.070 8.160 3.260 ;
        RECT 10.120 3.190 10.450 3.340 ;
        RECT 7.830 3.040 8.150 3.070 ;
        RECT 4.710 2.830 4.880 2.990 ;
        RECT 7.920 2.860 8.120 3.040 ;
        RECT 7.780 2.610 8.100 2.650 ;
        RECT 5.200 2.490 5.280 2.570 ;
        RECT 5.340 2.490 5.530 2.610 ;
        RECT 0.260 0.710 0.430 2.490 ;
        RECT 5.200 2.400 5.530 2.490 ;
        RECT 5.340 2.380 5.530 2.400 ;
        RECT 7.510 2.210 7.680 2.540 ;
        RECT 7.780 2.530 8.110 2.610 ;
        RECT 7.780 2.390 8.120 2.530 ;
        RECT 7.920 2.200 8.120 2.390 ;
        RECT 8.510 2.200 9.060 3.190 ;
        RECT 9.520 3.150 10.450 3.190 ;
        RECT 9.520 3.120 10.440 3.150 ;
        RECT 9.520 3.010 10.220 3.120 ;
        RECT 9.530 2.330 10.230 2.590 ;
        RECT 9.480 2.100 10.230 2.330 ;
        RECT 0.860 1.920 1.180 1.960 ;
        RECT 2.610 1.920 2.930 1.960 ;
        RECT 0.860 1.730 1.190 1.920 ;
        RECT 2.610 1.730 2.940 1.920 ;
        RECT 0.860 1.700 1.180 1.730 ;
        RECT 2.610 1.700 2.930 1.730 ;
        RECT 9.530 1.710 10.230 2.100 ;
        RECT 7.510 1.350 7.680 1.680 ;
        RECT 7.920 1.500 8.120 1.690 ;
        RECT 7.780 1.360 8.120 1.500 ;
        RECT 7.780 1.280 8.110 1.360 ;
        RECT 7.780 1.240 8.100 1.280 ;
        RECT 1.670 1.100 1.990 1.130 ;
        RECT 3.420 1.100 3.740 1.130 ;
        RECT 1.660 0.910 1.990 1.100 ;
        RECT 3.410 0.910 3.740 1.100 ;
        RECT 1.670 0.870 1.990 0.910 ;
        RECT 3.420 0.870 3.740 0.910 ;
        RECT 7.780 1.030 7.960 1.240 ;
        RECT 7.780 0.850 8.120 1.030 ;
        RECT 7.780 0.820 8.150 0.850 ;
        RECT 7.780 0.630 8.160 0.820 ;
        RECT 8.510 0.700 9.060 1.690 ;
        RECT 9.530 1.130 10.240 1.270 ;
        RECT 9.530 1.100 10.360 1.130 ;
        RECT 9.880 1.090 10.360 1.100 ;
        RECT 9.880 0.900 10.370 1.090 ;
        RECT 9.880 0.870 10.360 0.900 ;
        RECT 9.880 0.820 10.240 0.870 ;
        RECT 7.780 0.590 8.150 0.630 ;
        RECT 1.420 0.450 1.590 0.470 ;
        RECT 3.170 0.450 3.340 0.470 ;
        RECT 1.420 0.300 1.660 0.450 ;
        RECT 3.170 0.300 3.410 0.450 ;
        RECT 1.420 0.140 1.840 0.300 ;
        RECT 3.170 0.140 3.590 0.300 ;
        RECT 1.510 0.080 1.840 0.140 ;
        RECT 3.260 0.080 3.590 0.140 ;
        RECT 1.520 0.040 1.840 0.080 ;
        RECT 3.270 0.040 3.590 0.080 ;
        RECT 7.780 0.000 7.960 0.590 ;
        RECT 8.590 0.000 8.760 0.700 ;
        RECT 9.880 0.650 10.510 0.820 ;
      LAYER mcon ;
        RECT 0.960 5.900 1.130 6.070 ;
        RECT 0.250 5.350 0.420 5.520 ;
        RECT 0.840 5.300 1.010 5.470 ;
        RECT 0.250 5.010 0.420 5.180 ;
        RECT 4.920 6.070 5.090 6.240 ;
        RECT 5.070 5.240 5.240 5.410 ;
        RECT 7.890 6.080 8.060 6.250 ;
        RECT 8.830 5.690 9.000 5.860 ;
        RECT 10.140 6.100 10.310 6.270 ;
        RECT 7.840 5.430 8.010 5.600 ;
        RECT 0.250 4.670 0.420 4.840 ;
        RECT 1.800 4.620 1.970 4.790 ;
        RECT 7.670 4.720 7.840 4.890 ;
        RECT 9.490 4.720 9.660 4.890 ;
        RECT 0.250 4.330 0.420 4.500 ;
        RECT 4.230 4.420 4.400 4.590 ;
        RECT 0.250 3.990 0.420 4.160 ;
        RECT 7.840 4.290 8.010 4.460 ;
        RECT 7.670 4.020 7.840 4.190 ;
        RECT 8.830 4.030 9.000 4.200 ;
        RECT 2.040 3.750 2.210 3.920 ;
        RECT 3.790 3.750 3.960 3.920 ;
        RECT 1.650 3.020 1.820 3.190 ;
        RECT 3.400 3.020 3.570 3.190 ;
        RECT 7.890 3.640 8.060 3.810 ;
        RECT 10.190 3.880 10.360 4.050 ;
        RECT 4.960 3.140 5.130 3.310 ;
        RECT 7.890 3.080 8.060 3.250 ;
        RECT 10.180 3.160 10.350 3.330 ;
        RECT 8.830 2.690 9.000 2.860 ;
        RECT 0.260 2.320 0.430 2.490 ;
        RECT 5.350 2.410 5.520 2.580 ;
        RECT 7.840 2.430 8.010 2.600 ;
        RECT 0.260 1.980 0.430 2.150 ;
        RECT 9.490 2.130 9.660 2.300 ;
        RECT 0.260 1.640 0.430 1.810 ;
        RECT 0.920 1.740 1.090 1.910 ;
        RECT 2.670 1.740 2.840 1.910 ;
        RECT 0.260 1.300 0.430 1.470 ;
        RECT 7.840 1.290 8.010 1.460 ;
        RECT 0.260 0.960 0.430 1.130 ;
        RECT 1.760 0.920 1.930 1.090 ;
        RECT 3.510 0.920 3.680 1.090 ;
        RECT 8.830 1.030 9.000 1.200 ;
        RECT 7.890 0.640 8.060 0.810 ;
        RECT 10.100 0.910 10.270 1.080 ;
        RECT 1.610 0.090 1.780 0.260 ;
        RECT 3.360 0.090 3.530 0.260 ;
      LAYER met1 ;
        RECT 0.890 5.830 1.210 6.150 ;
        RECT 4.840 6.000 5.160 6.320 ;
        RECT 7.820 6.190 8.140 6.330 ;
        RECT 7.590 6.040 8.140 6.190 ;
        RECT 7.820 6.010 8.140 6.040 ;
        RECT 8.640 5.920 8.980 6.310 ;
        RECT 0.220 5.720 0.750 5.730 ;
        RECT 0.220 5.710 1.010 5.720 ;
        RECT 0.220 5.410 1.040 5.710 ;
        RECT 0.220 5.120 1.070 5.410 ;
        RECT 4.990 5.170 5.310 5.490 ;
        RECT 7.770 5.360 8.090 5.680 ;
        RECT 8.640 5.630 9.030 5.920 ;
        RECT 0.220 4.870 1.040 5.120 ;
        RECT 0.220 1.990 0.860 4.870 ;
        RECT 1.730 4.550 2.050 4.870 ;
        RECT 4.160 4.340 4.480 4.660 ;
        RECT 7.620 4.530 7.940 4.930 ;
        RECT 5.240 4.330 5.450 4.440 ;
        RECT 5.220 4.010 5.480 4.330 ;
        RECT 7.620 4.210 8.090 4.530 ;
        RECT 8.640 4.260 8.980 5.630 ;
        RECT 9.310 4.950 9.580 6.300 ;
        RECT 10.070 6.030 10.390 6.350 ;
        RECT 9.310 4.660 9.690 4.950 ;
        RECT 7.620 4.010 7.940 4.210 ;
        RECT 2.010 3.690 2.240 3.980 ;
        RECT 3.760 3.690 3.990 3.980 ;
        RECT 1.580 2.950 1.900 3.270 ;
        RECT 1.930 2.320 2.140 3.660 ;
        RECT 3.330 2.950 3.650 3.270 ;
        RECT 3.680 2.320 3.890 3.660 ;
        RECT 4.890 3.060 5.210 3.380 ;
        RECT 5.240 2.670 5.450 4.010 ;
        RECT 7.650 4.000 7.940 4.010 ;
        RECT 8.640 3.970 9.030 4.260 ;
        RECT 7.820 3.560 8.140 3.880 ;
        RECT 7.820 3.010 8.140 3.330 ;
        RECT 8.640 2.920 8.980 3.970 ;
        RECT 5.320 2.350 5.550 2.640 ;
        RECT 7.770 2.360 8.090 2.680 ;
        RECT 8.640 2.630 9.030 2.920 ;
        RECT 1.910 2.000 2.170 2.320 ;
        RECT 3.660 2.000 3.920 2.320 ;
        RECT 0.220 1.670 1.170 1.990 ;
        RECT 1.930 1.890 2.140 2.000 ;
        RECT 2.600 1.670 2.920 1.990 ;
        RECT 3.680 1.890 3.890 2.000 ;
        RECT 0.220 0.690 0.860 1.670 ;
        RECT 7.770 1.210 8.090 1.530 ;
        RECT 8.640 1.260 8.980 2.630 ;
        RECT 9.310 2.360 9.580 4.660 ;
        RECT 10.120 3.810 10.440 4.130 ;
        RECT 10.110 3.090 10.430 3.410 ;
        RECT 9.310 2.070 9.690 2.360 ;
        RECT 1.680 0.840 2.000 1.160 ;
        RECT 3.430 0.840 3.750 1.160 ;
        RECT 8.640 0.970 9.030 1.260 ;
        RECT 0.440 0.680 0.860 0.690 ;
        RECT 7.820 0.560 8.140 0.880 ;
        RECT 8.640 0.590 8.980 0.970 ;
        RECT 9.310 0.600 9.580 2.070 ;
        RECT 10.030 0.840 10.350 1.160 ;
        RECT 1.530 0.010 1.850 0.330 ;
        RECT 3.280 0.010 3.600 0.330 ;
      LAYER via ;
        RECT 0.920 5.860 1.180 6.120 ;
        RECT 4.870 6.030 5.130 6.290 ;
        RECT 7.850 6.040 8.110 6.300 ;
        RECT 0.340 4.930 0.930 5.650 ;
        RECT 5.020 5.200 5.280 5.460 ;
        RECT 7.800 5.390 8.060 5.650 ;
        RECT 1.760 4.580 2.020 4.840 ;
        RECT 4.190 4.370 4.450 4.630 ;
        RECT 5.220 4.040 5.480 4.300 ;
        RECT 7.630 4.500 7.890 4.890 ;
        RECT 7.630 4.240 8.060 4.500 ;
        RECT 7.630 4.030 7.890 4.240 ;
        RECT 10.100 6.060 10.360 6.320 ;
        RECT 1.610 2.980 1.870 3.240 ;
        RECT 3.360 2.980 3.620 3.240 ;
        RECT 4.920 3.090 5.180 3.350 ;
        RECT 7.850 3.590 8.110 3.850 ;
        RECT 7.850 3.040 8.110 3.300 ;
        RECT 7.800 2.390 8.060 2.650 ;
        RECT 1.910 2.030 2.170 2.290 ;
        RECT 3.660 2.030 3.920 2.290 ;
        RECT 0.880 1.700 1.140 1.960 ;
        RECT 2.630 1.700 2.890 1.960 ;
        RECT 7.800 1.240 8.060 1.500 ;
        RECT 10.150 3.840 10.410 4.100 ;
        RECT 10.140 3.120 10.400 3.380 ;
        RECT 1.710 0.870 1.970 1.130 ;
        RECT 3.460 0.870 3.720 1.130 ;
        RECT 7.850 0.590 8.110 0.850 ;
        RECT 10.060 0.870 10.320 1.130 ;
        RECT 1.560 0.040 1.820 0.300 ;
        RECT 3.310 0.040 3.570 0.300 ;
      LAYER met2 ;
        RECT 5.000 5.310 5.310 5.500 ;
        RECT 4.960 5.060 5.700 5.310 ;
        RECT 7.330 5.250 7.660 5.460 ;
        RECT 7.770 5.360 8.080 5.690 ;
        RECT 5.450 4.940 5.700 5.060 ;
        RECT 1.730 4.670 2.040 4.880 ;
        RECT 1.730 4.550 4.070 4.670 ;
        RECT 1.880 4.450 4.070 4.550 ;
        RECT 4.160 4.330 4.470 4.660 ;
        RECT 5.480 4.300 5.690 4.380 ;
        RECT 5.190 4.280 5.690 4.300 ;
        RECT 5.140 4.090 5.690 4.280 ;
        RECT 5.140 4.030 5.610 4.090 ;
        RECT 10.120 3.970 10.430 4.140 ;
        RECT 7.950 3.880 10.600 3.970 ;
        RECT 7.820 3.740 10.600 3.880 ;
        RECT 7.820 3.550 8.130 3.740 ;
        RECT 7.820 3.140 8.130 3.340 ;
        RECT 10.110 3.140 10.420 3.420 ;
        RECT 7.690 2.920 10.600 3.140 ;
        RECT 1.830 2.050 2.300 2.300 ;
        RECT 3.580 2.210 4.050 2.300 ;
        RECT 7.330 2.250 7.660 2.460 ;
        RECT 7.770 2.360 8.080 2.690 ;
        RECT 3.580 2.050 5.690 2.210 ;
        RECT 1.880 2.030 2.200 2.050 ;
        RECT 3.630 2.030 5.690 2.050 ;
        RECT 3.920 2.010 5.690 2.030 ;
        RECT 2.350 1.660 2.510 1.840 ;
        RECT 2.600 1.670 2.910 2.000 ;
        RECT 2.330 1.650 2.510 1.660 ;
        RECT 2.110 1.520 2.510 1.650 ;
        RECT 2.110 1.270 2.470 1.520 ;
        RECT 7.330 1.430 7.660 1.640 ;
        RECT 3.630 1.270 5.690 1.410 ;
        RECT 1.650 1.030 2.470 1.270 ;
        RECT 3.400 1.200 5.690 1.270 ;
        RECT 7.770 1.200 8.080 1.530 ;
        RECT 1.650 1.020 2.200 1.030 ;
        RECT 3.400 1.020 3.950 1.200 ;
        RECT 1.690 0.830 2.000 1.020 ;
        RECT 3.440 0.830 3.750 1.020 ;
        RECT 10.030 0.980 10.340 1.170 ;
        RECT 7.680 0.750 10.390 0.980 ;
        RECT 7.820 0.550 8.130 0.750 ;
  END
END sky130_hilas_TA2SignalBiasCell

MACRO sky130_hilas_Tgate4Single01
  CLASS CORE ;
  FOREIGN sky130_hilas_Tgate4Single01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.760 BY 6.410 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPWR
    USE ANALOG ;
    ANTENNADIFFAREA 0.966800 ;
    PORT
      LAYER nwell ;
        RECT 0.120 0.000 2.880 6.410 ;
      LAYER met1 ;
        RECT 0.740 5.490 0.940 6.410 ;
        RECT 0.730 5.200 0.960 5.490 ;
        RECT 0.740 4.410 0.940 5.200 ;
        RECT 0.730 4.120 0.960 4.410 ;
        RECT 0.740 2.290 0.940 4.120 ;
        RECT 0.730 2.000 0.960 2.290 ;
        RECT 0.740 1.210 0.940 2.000 ;
        RECT 0.730 0.920 0.960 1.210 ;
        RECT 0.740 0.000 0.940 0.920 ;
    END
  END VPWR
  PIN INPUT1_2
    USE ANALOG ;
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT 1.640 3.570 1.950 3.690 ;
        RECT 0.870 3.560 1.990 3.570 ;
        RECT 3.210 3.560 3.520 3.690 ;
        RECT 0.000 3.360 3.520 3.560 ;
        RECT 0.870 3.350 1.990 3.360 ;
    END
  END INPUT1_2
  PIN SELECT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT 0.290 4.540 0.610 4.630 ;
        RECT 0.000 4.340 0.610 4.540 ;
    END
  END SELECT2
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 4.250 5.490 4.440 6.410 ;
        RECT 4.230 5.200 4.460 5.490 ;
        RECT 4.250 4.410 4.440 5.200 ;
        RECT 4.230 4.120 4.460 4.410 ;
        RECT 4.250 2.290 4.440 4.120 ;
        RECT 4.230 2.000 4.460 2.290 ;
        RECT 4.250 1.210 4.440 2.000 ;
        RECT 4.230 0.920 4.460 1.210 ;
        RECT 4.250 0.000 4.440 0.920 ;
    END
  END VGND
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.212400 ;
    PORT
      LAYER met2 ;
        RECT 2.560 4.540 2.880 4.560 ;
        RECT 3.570 4.540 3.890 4.570 ;
        RECT 2.510 4.340 4.760 4.540 ;
        RECT 2.560 4.300 2.880 4.340 ;
        RECT 3.570 4.310 3.890 4.340 ;
    END
  END OUTPUT2
  PIN OUTPUT4
    ANTENNADIFFAREA 0.212400 ;
    PORT
      LAYER met2 ;
        RECT 2.560 1.340 2.880 1.360 ;
        RECT 3.570 1.340 3.890 1.370 ;
        RECT 2.510 1.140 4.760 1.340 ;
        RECT 2.560 1.100 2.880 1.140 ;
        RECT 3.570 1.110 3.890 1.140 ;
    END
  END OUTPUT4
  PIN OUTPUT3
    ANTENNADIFFAREA 0.212400 ;
    PORT
      LAYER met2 ;
        RECT 2.560 2.070 2.880 2.110 ;
        RECT 3.570 2.070 3.890 2.100 ;
        RECT 2.510 1.870 4.760 2.070 ;
        RECT 2.560 1.850 2.880 1.870 ;
        RECT 3.570 1.840 3.890 1.870 ;
    END
  END OUTPUT3
  PIN OUTPUT1
    ANTENNADIFFAREA 0.212400 ;
    PORT
      LAYER met2 ;
        RECT 2.560 5.270 2.880 5.310 ;
        RECT 3.570 5.270 3.890 5.300 ;
        RECT 2.510 5.070 4.760 5.270 ;
        RECT 2.560 5.050 2.880 5.070 ;
        RECT 3.570 5.040 3.890 5.070 ;
    END
  END OUTPUT1
  PIN INPUT1_4
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT 1.640 0.370 1.950 0.490 ;
        RECT 0.870 0.360 1.990 0.370 ;
        RECT 3.210 0.360 3.520 0.490 ;
        RECT 0.000 0.160 3.520 0.360 ;
        RECT 0.870 0.150 1.990 0.160 ;
    END
  END INPUT1_4
  PIN SELECT4
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT 0.290 1.340 0.610 1.430 ;
        RECT 0.000 1.140 0.610 1.340 ;
    END
  END SELECT4
  PIN SELECT3
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT 0.000 1.870 0.610 2.070 ;
        RECT 0.290 1.780 0.610 1.870 ;
    END
  END SELECT3
  PIN INPUT1_3
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT 0.870 3.050 1.990 3.060 ;
        RECT 0.000 2.850 3.520 3.050 ;
        RECT 0.870 2.840 1.990 2.850 ;
        RECT 1.640 2.720 1.950 2.840 ;
        RECT 3.210 2.720 3.520 2.850 ;
    END
  END INPUT1_3
  PIN SELECT1
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT 0.000 5.070 0.610 5.270 ;
        RECT 0.290 4.980 0.610 5.070 ;
    END
  END SELECT1
  PIN INPUT1_1
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT 0.870 6.250 1.990 6.260 ;
        RECT 0.000 6.050 3.520 6.250 ;
        RECT 0.870 6.040 1.990 6.050 ;
        RECT 1.640 5.920 1.950 6.040 ;
        RECT 3.210 5.920 3.520 6.050 ;
    END
  END INPUT1_1
  OBS
      LAYER li1 ;
        RECT 1.650 6.190 1.970 6.220 ;
        RECT 3.220 6.190 3.540 6.220 ;
        RECT 0.430 5.850 0.600 6.130 ;
        RECT 1.650 6.000 1.980 6.190 ;
        RECT 2.660 6.050 2.850 6.070 ;
        RECT 1.650 5.960 1.970 6.000 ;
        RECT 0.430 5.810 0.640 5.850 ;
        RECT 0.430 5.790 0.660 5.810 ;
        RECT 1.780 5.800 1.950 5.960 ;
        RECT 2.390 5.880 2.850 6.050 ;
        RECT 3.220 6.000 3.550 6.190 ;
        RECT 3.790 6.050 3.980 6.080 ;
        RECT 3.220 5.960 3.540 6.000 ;
        RECT 2.640 5.870 2.850 5.880 ;
        RECT 2.660 5.840 2.850 5.870 ;
        RECT 3.280 5.800 3.450 5.960 ;
        RECT 3.790 5.880 4.230 6.050 ;
        RECT 3.790 5.850 3.980 5.880 ;
        RECT 0.430 5.770 0.690 5.790 ;
        RECT 0.430 5.720 0.770 5.770 ;
        RECT 0.430 5.660 0.920 5.720 ;
        RECT 0.430 5.630 0.940 5.660 ;
        RECT 0.470 5.600 0.940 5.630 ;
        RECT 0.600 5.550 0.940 5.600 ;
        RECT 0.720 5.540 0.940 5.550 ;
        RECT 0.730 5.510 0.940 5.540 ;
        RECT 0.750 5.430 0.940 5.510 ;
        RECT 2.110 5.430 2.440 5.550 ;
        RECT 4.510 5.460 4.680 6.140 ;
        RECT 0.260 5.380 0.430 5.400 ;
        RECT 0.240 4.950 0.450 5.380 ;
        RECT 0.750 5.260 1.270 5.430 ;
        RECT 0.750 5.230 0.940 5.260 ;
        RECT 1.620 5.250 3.520 5.430 ;
        RECT 4.250 5.420 4.680 5.460 ;
        RECT 3.900 5.260 4.680 5.420 ;
        RECT 3.900 5.250 4.440 5.260 ;
        RECT 4.250 5.230 4.440 5.250 ;
        RECT 0.240 4.230 0.450 4.660 ;
        RECT 0.750 4.350 0.940 4.380 ;
        RECT 4.250 4.360 4.440 4.380 ;
        RECT 0.260 4.210 0.430 4.230 ;
        RECT 0.750 4.180 1.270 4.350 ;
        RECT 1.620 4.180 3.520 4.360 ;
        RECT 3.900 4.350 4.440 4.360 ;
        RECT 3.900 4.190 4.680 4.350 ;
        RECT 0.750 4.100 0.940 4.180 ;
        RECT 0.730 4.070 0.940 4.100 ;
        RECT 0.720 4.060 0.940 4.070 ;
        RECT 2.110 4.060 2.440 4.180 ;
        RECT 4.250 4.150 4.680 4.190 ;
        RECT 0.600 4.010 0.940 4.060 ;
        RECT 0.470 3.980 0.940 4.010 ;
        RECT 0.430 3.950 0.940 3.980 ;
        RECT 0.430 3.890 0.920 3.950 ;
        RECT 0.430 3.840 0.770 3.890 ;
        RECT 0.430 3.820 0.690 3.840 ;
        RECT 0.430 3.800 0.660 3.820 ;
        RECT 0.430 3.760 0.640 3.800 ;
        RECT 0.430 3.480 0.600 3.760 ;
        RECT 1.780 3.650 1.950 3.810 ;
        RECT 2.660 3.740 2.850 3.770 ;
        RECT 2.640 3.730 2.850 3.740 ;
        RECT 1.650 3.610 1.970 3.650 ;
        RECT 1.650 3.420 1.980 3.610 ;
        RECT 2.390 3.560 2.850 3.730 ;
        RECT 3.280 3.650 3.450 3.810 ;
        RECT 3.790 3.730 3.980 3.760 ;
        RECT 2.660 3.540 2.850 3.560 ;
        RECT 3.220 3.610 3.540 3.650 ;
        RECT 3.220 3.420 3.550 3.610 ;
        RECT 3.790 3.560 4.230 3.730 ;
        RECT 3.790 3.530 3.980 3.560 ;
        RECT 4.510 3.470 4.680 4.150 ;
        RECT 1.650 3.390 1.970 3.420 ;
        RECT 3.220 3.390 3.540 3.420 ;
        RECT 1.650 2.990 1.970 3.020 ;
        RECT 3.220 2.990 3.540 3.020 ;
        RECT 0.430 2.650 0.600 2.930 ;
        RECT 1.650 2.800 1.980 2.990 ;
        RECT 2.660 2.850 2.850 2.870 ;
        RECT 1.650 2.760 1.970 2.800 ;
        RECT 0.430 2.610 0.640 2.650 ;
        RECT 0.430 2.590 0.660 2.610 ;
        RECT 1.780 2.600 1.950 2.760 ;
        RECT 2.390 2.680 2.850 2.850 ;
        RECT 3.220 2.800 3.550 2.990 ;
        RECT 3.790 2.850 3.980 2.880 ;
        RECT 3.220 2.760 3.540 2.800 ;
        RECT 2.640 2.670 2.850 2.680 ;
        RECT 2.660 2.640 2.850 2.670 ;
        RECT 3.280 2.600 3.450 2.760 ;
        RECT 3.790 2.680 4.230 2.850 ;
        RECT 3.790 2.650 3.980 2.680 ;
        RECT 0.430 2.570 0.690 2.590 ;
        RECT 0.430 2.520 0.770 2.570 ;
        RECT 0.430 2.460 0.920 2.520 ;
        RECT 0.430 2.430 0.940 2.460 ;
        RECT 0.470 2.400 0.940 2.430 ;
        RECT 0.600 2.350 0.940 2.400 ;
        RECT 0.720 2.340 0.940 2.350 ;
        RECT 0.730 2.310 0.940 2.340 ;
        RECT 0.750 2.230 0.940 2.310 ;
        RECT 2.110 2.230 2.440 2.350 ;
        RECT 4.510 2.260 4.680 2.940 ;
        RECT 0.260 2.180 0.430 2.200 ;
        RECT 0.240 1.750 0.450 2.180 ;
        RECT 0.750 2.060 1.270 2.230 ;
        RECT 0.750 2.030 0.940 2.060 ;
        RECT 1.620 2.050 3.520 2.230 ;
        RECT 4.250 2.220 4.680 2.260 ;
        RECT 3.900 2.060 4.680 2.220 ;
        RECT 3.900 2.050 4.440 2.060 ;
        RECT 4.250 2.030 4.440 2.050 ;
        RECT 0.240 1.030 0.450 1.460 ;
        RECT 0.750 1.150 0.940 1.180 ;
        RECT 4.250 1.160 4.440 1.180 ;
        RECT 0.260 1.010 0.430 1.030 ;
        RECT 0.750 0.980 1.270 1.150 ;
        RECT 1.620 0.980 3.520 1.160 ;
        RECT 3.900 1.150 4.440 1.160 ;
        RECT 3.900 0.990 4.680 1.150 ;
        RECT 0.750 0.900 0.940 0.980 ;
        RECT 0.730 0.870 0.940 0.900 ;
        RECT 0.720 0.860 0.940 0.870 ;
        RECT 2.110 0.860 2.440 0.980 ;
        RECT 4.250 0.950 4.680 0.990 ;
        RECT 0.600 0.810 0.940 0.860 ;
        RECT 0.470 0.780 0.940 0.810 ;
        RECT 0.430 0.750 0.940 0.780 ;
        RECT 0.430 0.690 0.920 0.750 ;
        RECT 0.430 0.640 0.770 0.690 ;
        RECT 0.430 0.620 0.690 0.640 ;
        RECT 0.430 0.600 0.660 0.620 ;
        RECT 0.430 0.560 0.640 0.600 ;
        RECT 0.430 0.280 0.600 0.560 ;
        RECT 1.780 0.450 1.950 0.610 ;
        RECT 2.660 0.540 2.850 0.570 ;
        RECT 2.640 0.530 2.850 0.540 ;
        RECT 1.650 0.410 1.970 0.450 ;
        RECT 1.650 0.220 1.980 0.410 ;
        RECT 2.390 0.360 2.850 0.530 ;
        RECT 3.280 0.450 3.450 0.610 ;
        RECT 3.790 0.530 3.980 0.560 ;
        RECT 2.660 0.340 2.850 0.360 ;
        RECT 3.220 0.410 3.540 0.450 ;
        RECT 3.220 0.220 3.550 0.410 ;
        RECT 3.790 0.360 4.230 0.530 ;
        RECT 3.790 0.330 3.980 0.360 ;
        RECT 4.510 0.270 4.680 0.950 ;
        RECT 1.650 0.190 1.970 0.220 ;
        RECT 3.220 0.190 3.540 0.220 ;
      LAYER mcon ;
        RECT 1.710 6.010 1.880 6.180 ;
        RECT 2.670 5.870 2.840 6.040 ;
        RECT 3.280 6.010 3.450 6.180 ;
        RECT 3.800 5.880 3.970 6.050 ;
        RECT 0.260 5.230 0.430 5.400 ;
        RECT 0.760 5.260 0.930 5.430 ;
        RECT 4.260 5.260 4.430 5.430 ;
        RECT 0.760 4.180 0.930 4.350 ;
        RECT 4.260 4.180 4.430 4.350 ;
        RECT 1.710 3.430 1.880 3.600 ;
        RECT 2.670 3.570 2.840 3.740 ;
        RECT 3.280 3.430 3.450 3.600 ;
        RECT 3.800 3.560 3.970 3.730 ;
        RECT 1.710 2.810 1.880 2.980 ;
        RECT 2.670 2.670 2.840 2.840 ;
        RECT 3.280 2.810 3.450 2.980 ;
        RECT 3.800 2.680 3.970 2.850 ;
        RECT 0.260 2.030 0.430 2.200 ;
        RECT 0.760 2.060 0.930 2.230 ;
        RECT 4.260 2.060 4.430 2.230 ;
        RECT 0.760 0.980 0.930 1.150 ;
        RECT 4.260 0.980 4.430 1.150 ;
        RECT 1.710 0.230 1.880 0.400 ;
        RECT 2.670 0.370 2.840 0.540 ;
        RECT 3.280 0.230 3.450 0.400 ;
        RECT 3.800 0.360 3.970 0.530 ;
      LAYER met1 ;
        RECT 1.640 5.930 1.960 6.250 ;
        RECT 2.640 5.810 2.870 6.100 ;
        RECT 3.210 5.930 3.530 6.250 ;
        RECT 3.770 5.820 4.000 6.110 ;
        RECT 0.230 5.270 0.460 5.460 ;
        RECT 2.660 5.340 2.850 5.810 ;
        RECT 0.230 5.170 0.580 5.270 ;
        RECT 0.240 4.950 0.580 5.170 ;
        RECT 2.590 5.020 2.850 5.340 ;
        RECT 3.770 5.330 3.960 5.820 ;
        RECT 3.590 5.080 3.960 5.330 ;
        RECT 3.590 5.010 3.860 5.080 ;
        RECT 0.240 4.440 0.580 4.660 ;
        RECT 0.230 4.340 0.580 4.440 ;
        RECT 0.230 4.150 0.460 4.340 ;
        RECT 2.590 4.270 2.850 4.590 ;
        RECT 3.590 4.530 3.860 4.600 ;
        RECT 3.590 4.280 3.960 4.530 ;
        RECT 2.660 3.800 2.850 4.270 ;
        RECT 1.640 3.360 1.960 3.680 ;
        RECT 2.640 3.510 2.870 3.800 ;
        RECT 3.770 3.790 3.960 4.280 ;
        RECT 3.210 3.360 3.530 3.680 ;
        RECT 3.770 3.500 4.000 3.790 ;
        RECT 1.640 2.730 1.960 3.050 ;
        RECT 2.640 2.610 2.870 2.900 ;
        RECT 3.210 2.730 3.530 3.050 ;
        RECT 3.770 2.620 4.000 2.910 ;
        RECT 0.230 2.070 0.460 2.260 ;
        RECT 2.660 2.140 2.850 2.610 ;
        RECT 0.230 1.970 0.580 2.070 ;
        RECT 0.240 1.750 0.580 1.970 ;
        RECT 2.590 1.820 2.850 2.140 ;
        RECT 3.770 2.130 3.960 2.620 ;
        RECT 3.590 1.880 3.960 2.130 ;
        RECT 3.590 1.810 3.860 1.880 ;
        RECT 0.240 1.240 0.580 1.460 ;
        RECT 0.230 1.140 0.580 1.240 ;
        RECT 0.230 0.950 0.460 1.140 ;
        RECT 2.590 1.070 2.850 1.390 ;
        RECT 3.590 1.330 3.860 1.400 ;
        RECT 3.590 1.080 3.960 1.330 ;
        RECT 2.660 0.600 2.850 1.070 ;
        RECT 1.640 0.160 1.960 0.480 ;
        RECT 2.640 0.310 2.870 0.600 ;
        RECT 3.770 0.590 3.960 1.080 ;
        RECT 3.210 0.160 3.530 0.480 ;
        RECT 3.770 0.300 4.000 0.590 ;
      LAYER via ;
        RECT 1.670 5.960 1.930 6.220 ;
        RECT 3.240 5.960 3.500 6.220 ;
        RECT 0.320 4.980 0.580 5.240 ;
        RECT 2.590 5.050 2.850 5.310 ;
        RECT 3.600 5.040 3.860 5.300 ;
        RECT 0.320 4.370 0.580 4.630 ;
        RECT 2.590 4.300 2.850 4.560 ;
        RECT 3.600 4.310 3.860 4.570 ;
        RECT 1.670 3.390 1.930 3.650 ;
        RECT 3.240 3.390 3.500 3.650 ;
        RECT 1.670 2.760 1.930 3.020 ;
        RECT 3.240 2.760 3.500 3.020 ;
        RECT 0.320 1.780 0.580 2.040 ;
        RECT 2.590 1.850 2.850 2.110 ;
        RECT 3.600 1.840 3.860 2.100 ;
        RECT 0.320 1.170 0.580 1.430 ;
        RECT 2.590 1.100 2.850 1.360 ;
        RECT 3.600 1.110 3.860 1.370 ;
        RECT 1.670 0.190 1.930 0.450 ;
        RECT 3.240 0.190 3.500 0.450 ;
  END
END sky130_hilas_Tgate4Single01

MACRO sky130_hilas_VinjDecode2to4
  CLASS CORE ;
  FOREIGN sky130_hilas_VinjDecode2to4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.950 BY 6.160 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN OUTPUT00
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 9.570 5.010 9.940 5.090 ;
        RECT 9.570 5.000 10.600 5.010 ;
        RECT 12.480 5.000 12.790 5.160 ;
        RECT 9.570 4.830 12.950 5.000 ;
    END
  END OUTPUT00
  PIN OUTPUT01
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 9.570 3.500 9.940 3.580 ;
        RECT 9.570 3.490 10.600 3.500 ;
        RECT 12.480 3.490 12.790 3.650 ;
        RECT 9.570 3.320 12.950 3.490 ;
    END
  END OUTPUT01
  PIN OUTPUT10
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 9.570 1.990 9.940 2.070 ;
        RECT 9.570 1.980 10.600 1.990 ;
        RECT 12.480 1.980 12.790 2.140 ;
        RECT 9.570 1.810 12.950 1.980 ;
    END
  END OUTPUT10
  PIN OUTPUT11
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 9.570 0.490 9.940 0.570 ;
        RECT 9.570 0.480 10.600 0.490 ;
        RECT 12.480 0.480 12.790 0.640 ;
        RECT 9.570 0.310 12.950 0.480 ;
    END
  END OUTPUT11
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 11.660 0.090 11.930 6.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.180 1.590 3.410 6.120 ;
    END
  END VGND
  PIN VINJ
    ANTENNADIFFAREA 0.914000 ;
    PORT
      LAYER nwell ;
        RECT 6.080 0.000 9.520 6.160 ;
      LAYER met1 ;
        RECT 6.690 5.780 6.910 6.120 ;
        RECT 6.690 5.520 6.920 5.780 ;
        RECT 6.690 5.120 6.910 5.520 ;
        RECT 6.690 4.810 6.940 5.120 ;
        RECT 6.690 4.270 6.910 4.810 ;
        RECT 6.690 4.010 6.920 4.270 ;
        RECT 6.690 3.610 6.910 4.010 ;
        RECT 6.690 3.300 6.940 3.610 ;
        RECT 6.690 2.760 6.910 3.300 ;
        RECT 6.690 2.500 6.920 2.760 ;
        RECT 6.690 2.100 6.910 2.500 ;
        RECT 6.690 1.790 6.940 2.100 ;
        RECT 6.690 1.260 6.910 1.790 ;
        RECT 6.690 1.000 6.920 1.260 ;
        RECT 6.690 0.600 6.910 1.000 ;
        RECT 6.690 0.290 6.940 0.600 ;
        RECT 6.690 0.090 6.910 0.290 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.000 1.500 1.980 6.160 ;
      LAYER met1 ;
        RECT 0.610 5.780 0.830 6.120 ;
        RECT 0.610 5.520 0.840 5.780 ;
        RECT 0.610 5.120 0.830 5.520 ;
        RECT 0.610 4.810 0.860 5.120 ;
        RECT 0.610 4.270 0.830 4.810 ;
        RECT 0.610 4.010 0.840 4.270 ;
        RECT 0.610 3.610 0.830 4.010 ;
        RECT 0.610 3.300 0.860 3.610 ;
        RECT 0.610 2.760 0.830 3.300 ;
        RECT 0.610 2.500 0.840 2.760 ;
        RECT 0.610 2.100 0.830 2.500 ;
        RECT 0.610 1.790 0.860 2.100 ;
        RECT 0.610 1.590 0.830 1.790 ;
    END
  END VINJ
  PIN IN2
    ANTENNAGATEAREA 0.642800 ;
    PORT
      LAYER met2 ;
        RECT 4.560 5.520 4.890 5.580 ;
        RECT 8.710 5.540 9.040 5.620 ;
        RECT 8.440 5.520 9.040 5.540 ;
        RECT 4.560 5.360 9.040 5.520 ;
        RECT 4.560 5.310 4.890 5.360 ;
        RECT 0.000 4.200 4.790 4.220 ;
        RECT 0.000 4.040 4.840 4.200 ;
        RECT 4.570 4.010 4.840 4.040 ;
        RECT 4.570 3.870 4.850 4.010 ;
        RECT 4.620 3.850 4.850 3.870 ;
        RECT 4.540 2.500 4.870 2.560 ;
        RECT 8.710 2.520 9.040 2.600 ;
        RECT 8.440 2.500 9.040 2.520 ;
        RECT 4.540 2.340 9.040 2.500 ;
        RECT 4.540 2.290 4.870 2.340 ;
    END
  END IN2
  PIN IN1
    ANTENNAGATEAREA 0.673600 ;
    PORT
      LAYER met2 ;
        RECT 3.710 5.960 10.110 5.970 ;
        RECT 3.690 5.810 10.110 5.960 ;
        RECT 3.690 5.800 3.960 5.810 ;
        RECT 3.660 5.730 3.960 5.800 ;
        RECT 0.000 5.550 3.960 5.730 ;
        RECT 9.690 5.580 10.110 5.810 ;
        RECT 3.660 5.470 3.930 5.550 ;
        RECT 3.630 4.630 3.960 4.690 ;
        RECT 3.630 4.470 5.270 4.630 ;
        RECT 3.630 4.420 3.960 4.470 ;
        RECT 5.110 4.460 5.270 4.470 ;
        RECT 5.110 4.300 10.110 4.460 ;
        RECT 9.690 4.070 10.110 4.300 ;
    END
  END IN1
  PIN ENABLE
    PORT
      LAYER met2 ;
        RECT 0.000 2.530 3.610 2.710 ;
    END
  END ENABLE
  OBS
      LAYER li1 ;
        RECT 0.620 5.730 0.790 5.870 ;
        RECT 6.700 5.730 6.870 5.870 ;
        RECT 7.430 5.750 7.600 5.830 ;
        RECT 8.240 5.750 8.410 5.830 ;
        RECT 9.780 5.790 9.950 5.910 ;
        RECT 0.620 5.560 0.810 5.730 ;
        RECT 0.620 5.460 0.790 5.560 ;
        RECT 0.190 5.080 0.360 5.180 ;
        RECT 0.170 4.910 0.360 5.080 ;
        RECT 0.190 4.850 0.360 4.910 ;
        RECT 0.610 5.120 0.780 5.180 ;
        RECT 0.610 4.850 0.860 5.120 ;
        RECT 1.350 5.100 1.600 5.180 ;
        RECT 1.350 4.930 2.650 5.100 ;
        RECT 3.210 5.090 3.380 5.720 ;
        RECT 6.700 5.560 6.890 5.730 ;
        RECT 6.700 5.460 6.870 5.560 ;
        RECT 7.430 5.180 7.640 5.750 ;
        RECT 8.200 5.500 8.410 5.750 ;
        RECT 8.800 5.570 8.970 5.670 ;
        RECT 9.740 5.620 9.950 5.790 ;
        RECT 11.670 5.720 11.930 5.790 ;
        RECT 12.470 5.720 12.650 5.850 ;
        RECT 9.780 5.580 9.950 5.620 ;
        RECT 8.200 5.180 8.370 5.500 ;
        RECT 8.770 5.400 8.970 5.570 ;
        RECT 8.800 5.300 8.970 5.400 ;
        RECT 10.340 5.540 11.210 5.710 ;
        RECT 11.670 5.540 12.650 5.720 ;
        RECT 0.620 4.830 0.860 4.850 ;
        RECT 1.430 4.840 1.600 4.930 ;
        RECT 3.130 4.920 3.460 5.090 ;
        RECT 6.270 5.080 6.440 5.180 ;
        RECT 6.250 4.910 6.440 5.080 ;
        RECT 6.270 4.850 6.440 4.910 ;
        RECT 6.690 5.120 6.860 5.180 ;
        RECT 6.690 4.850 6.940 5.120 ;
        RECT 7.430 4.930 7.680 5.180 ;
        RECT 6.700 4.830 6.940 4.850 ;
        RECT 7.510 4.840 7.680 4.930 ;
        RECT 8.160 4.930 8.370 5.180 ;
        RECT 10.340 5.100 10.510 5.540 ;
        RECT 11.670 5.100 11.930 5.540 ;
        RECT 12.470 5.430 12.650 5.540 ;
        RECT 8.880 4.930 10.510 5.100 ;
        RECT 10.960 4.930 11.930 5.100 ;
        RECT 12.380 4.930 12.720 5.100 ;
        RECT 8.160 4.850 8.330 4.930 ;
        RECT 9.650 4.890 9.820 4.930 ;
        RECT 0.620 4.220 0.790 4.360 ;
        RECT 6.700 4.220 6.870 4.360 ;
        RECT 7.430 4.240 7.600 4.320 ;
        RECT 8.240 4.240 8.410 4.320 ;
        RECT 9.780 4.280 9.950 4.400 ;
        RECT 0.620 4.050 0.810 4.220 ;
        RECT 0.620 3.950 0.790 4.050 ;
        RECT 0.190 3.570 0.360 3.670 ;
        RECT 0.170 3.400 0.360 3.570 ;
        RECT 0.190 3.340 0.360 3.400 ;
        RECT 0.610 3.610 0.780 3.670 ;
        RECT 0.610 3.340 0.860 3.610 ;
        RECT 1.350 3.590 1.600 3.670 ;
        RECT 1.350 3.420 2.650 3.590 ;
        RECT 3.210 3.580 3.380 4.210 ;
        RECT 6.700 4.050 6.890 4.220 ;
        RECT 6.700 3.950 6.870 4.050 ;
        RECT 7.430 3.670 7.640 4.240 ;
        RECT 8.200 3.990 8.410 4.240 ;
        RECT 8.800 4.060 8.970 4.160 ;
        RECT 9.740 4.110 9.950 4.280 ;
        RECT 11.670 4.210 11.930 4.280 ;
        RECT 12.470 4.210 12.650 4.340 ;
        RECT 9.780 4.070 9.950 4.110 ;
        RECT 8.200 3.670 8.370 3.990 ;
        RECT 8.770 3.890 8.970 4.060 ;
        RECT 8.800 3.790 8.970 3.890 ;
        RECT 10.340 4.030 11.210 4.200 ;
        RECT 11.670 4.030 12.650 4.210 ;
        RECT 0.620 3.320 0.860 3.340 ;
        RECT 1.430 3.330 1.600 3.420 ;
        RECT 3.130 3.410 3.460 3.580 ;
        RECT 6.270 3.570 6.440 3.670 ;
        RECT 6.250 3.400 6.440 3.570 ;
        RECT 6.270 3.340 6.440 3.400 ;
        RECT 6.690 3.610 6.860 3.670 ;
        RECT 6.690 3.340 6.940 3.610 ;
        RECT 7.430 3.420 7.680 3.670 ;
        RECT 6.700 3.320 6.940 3.340 ;
        RECT 7.510 3.330 7.680 3.420 ;
        RECT 8.160 3.420 8.370 3.670 ;
        RECT 10.340 3.590 10.510 4.030 ;
        RECT 11.670 3.590 11.930 4.030 ;
        RECT 12.470 3.920 12.650 4.030 ;
        RECT 8.880 3.420 10.510 3.590 ;
        RECT 10.960 3.420 11.930 3.590 ;
        RECT 12.380 3.420 12.720 3.590 ;
        RECT 8.160 3.340 8.330 3.420 ;
        RECT 9.650 3.380 9.820 3.420 ;
        RECT 0.620 2.710 0.790 2.850 ;
        RECT 6.700 2.710 6.870 2.850 ;
        RECT 7.430 2.730 7.600 2.810 ;
        RECT 8.240 2.730 8.410 2.810 ;
        RECT 9.780 2.770 9.950 2.890 ;
        RECT 0.620 2.540 0.810 2.710 ;
        RECT 0.620 2.440 0.790 2.540 ;
        RECT 0.190 2.060 0.360 2.160 ;
        RECT 0.170 1.890 0.360 2.060 ;
        RECT 0.190 1.830 0.360 1.890 ;
        RECT 0.610 2.100 0.780 2.160 ;
        RECT 0.610 1.830 0.860 2.100 ;
        RECT 1.350 2.080 1.600 2.160 ;
        RECT 1.350 1.910 2.650 2.080 ;
        RECT 3.210 2.070 3.380 2.700 ;
        RECT 6.700 2.540 6.890 2.710 ;
        RECT 6.700 2.440 6.870 2.540 ;
        RECT 7.430 2.160 7.640 2.730 ;
        RECT 8.200 2.480 8.410 2.730 ;
        RECT 8.800 2.550 8.970 2.650 ;
        RECT 9.740 2.600 9.950 2.770 ;
        RECT 11.670 2.700 11.930 2.770 ;
        RECT 12.470 2.700 12.650 2.830 ;
        RECT 9.780 2.560 9.950 2.600 ;
        RECT 8.200 2.160 8.370 2.480 ;
        RECT 8.770 2.380 8.970 2.550 ;
        RECT 8.800 2.280 8.970 2.380 ;
        RECT 10.340 2.520 11.210 2.690 ;
        RECT 11.670 2.520 12.650 2.700 ;
        RECT 0.620 1.810 0.860 1.830 ;
        RECT 1.430 1.820 1.600 1.910 ;
        RECT 3.130 1.900 3.460 2.070 ;
        RECT 6.270 2.060 6.440 2.160 ;
        RECT 6.250 1.890 6.440 2.060 ;
        RECT 6.270 1.830 6.440 1.890 ;
        RECT 6.690 2.100 6.860 2.160 ;
        RECT 6.690 1.830 6.940 2.100 ;
        RECT 7.430 1.910 7.680 2.160 ;
        RECT 6.700 1.810 6.940 1.830 ;
        RECT 7.510 1.820 7.680 1.910 ;
        RECT 8.160 1.910 8.370 2.160 ;
        RECT 10.340 2.080 10.510 2.520 ;
        RECT 11.670 2.080 11.930 2.520 ;
        RECT 12.470 2.410 12.650 2.520 ;
        RECT 8.880 1.910 10.510 2.080 ;
        RECT 10.960 1.910 11.930 2.080 ;
        RECT 12.380 1.910 12.720 2.080 ;
        RECT 8.160 1.830 8.330 1.910 ;
        RECT 9.650 1.870 9.820 1.910 ;
        RECT 6.700 1.210 6.870 1.350 ;
        RECT 7.430 1.230 7.600 1.310 ;
        RECT 8.240 1.230 8.410 1.310 ;
        RECT 9.780 1.270 9.950 1.390 ;
        RECT 6.700 1.040 6.890 1.210 ;
        RECT 6.700 0.940 6.870 1.040 ;
        RECT 7.430 0.660 7.640 1.230 ;
        RECT 8.200 0.980 8.410 1.230 ;
        RECT 8.800 1.050 8.970 1.150 ;
        RECT 9.740 1.100 9.950 1.270 ;
        RECT 11.670 1.200 11.930 1.270 ;
        RECT 12.470 1.200 12.650 1.330 ;
        RECT 9.780 1.060 9.950 1.100 ;
        RECT 8.200 0.660 8.370 0.980 ;
        RECT 8.770 0.880 8.970 1.050 ;
        RECT 8.800 0.780 8.970 0.880 ;
        RECT 10.340 1.020 11.210 1.190 ;
        RECT 11.670 1.020 12.650 1.200 ;
        RECT 6.270 0.560 6.440 0.660 ;
        RECT 6.250 0.390 6.440 0.560 ;
        RECT 6.270 0.330 6.440 0.390 ;
        RECT 6.690 0.600 6.860 0.660 ;
        RECT 6.690 0.330 6.940 0.600 ;
        RECT 7.430 0.410 7.680 0.660 ;
        RECT 6.700 0.310 6.940 0.330 ;
        RECT 7.510 0.320 7.680 0.410 ;
        RECT 8.160 0.410 8.370 0.660 ;
        RECT 10.340 0.580 10.510 1.020 ;
        RECT 11.670 0.580 11.930 1.020 ;
        RECT 12.470 0.910 12.650 1.020 ;
        RECT 8.880 0.410 10.510 0.580 ;
        RECT 10.960 0.410 11.930 0.580 ;
        RECT 12.380 0.410 12.720 0.580 ;
        RECT 8.160 0.330 8.330 0.410 ;
        RECT 9.650 0.370 9.820 0.410 ;
      LAYER mcon ;
        RECT 0.640 5.560 0.810 5.730 ;
        RECT 6.720 5.560 6.890 5.730 ;
        RECT 3.210 5.200 3.380 5.370 ;
        RECT 0.650 4.880 0.820 5.050 ;
        RECT 1.990 4.930 2.160 5.100 ;
        RECT 6.730 4.880 6.900 5.050 ;
        RECT 11.700 5.220 11.880 5.400 ;
        RECT 0.640 4.050 0.810 4.220 ;
        RECT 6.720 4.050 6.890 4.220 ;
        RECT 3.210 3.690 3.380 3.860 ;
        RECT 0.650 3.370 0.820 3.540 ;
        RECT 1.990 3.420 2.160 3.590 ;
        RECT 6.730 3.370 6.900 3.540 ;
        RECT 11.700 3.710 11.880 3.890 ;
        RECT 0.640 2.540 0.810 2.710 ;
        RECT 6.720 2.540 6.890 2.710 ;
        RECT 3.210 2.180 3.380 2.350 ;
        RECT 0.650 1.860 0.820 2.030 ;
        RECT 1.990 1.910 2.160 2.080 ;
        RECT 6.730 1.860 6.900 2.030 ;
        RECT 11.700 2.200 11.880 2.380 ;
        RECT 6.720 1.040 6.890 1.210 ;
        RECT 6.730 0.360 6.900 0.530 ;
        RECT 11.700 0.700 11.880 0.880 ;
      LAYER met1 ;
        RECT 3.670 5.770 3.940 6.060 ;
        RECT 3.630 5.500 3.960 5.770 ;
        RECT 0.080 4.840 0.390 5.190 ;
        RECT 1.910 4.880 2.230 5.140 ;
        RECT 3.670 4.720 3.940 5.500 ;
        RECT 3.660 4.390 3.940 4.720 ;
        RECT 3.670 4.360 3.940 4.390 ;
        RECT 0.080 3.330 0.390 3.680 ;
        RECT 1.910 3.370 2.230 3.630 ;
        RECT 4.130 3.040 4.400 5.160 ;
        RECT 4.590 4.170 4.860 5.630 ;
        RECT 8.710 5.360 9.040 5.620 ;
        RECT 9.680 5.580 10.110 5.870 ;
        RECT 5.540 5.130 5.830 5.180 ;
        RECT 5.520 4.780 5.830 5.130 ;
        RECT 6.160 4.840 6.470 5.190 ;
        RECT 9.550 4.830 9.940 5.100 ;
        RECT 12.480 4.840 12.790 5.160 ;
        RECT 4.540 3.900 4.870 4.170 ;
        RECT 4.120 2.710 4.400 3.040 ;
        RECT 0.080 1.820 0.390 2.170 ;
        RECT 1.910 1.860 2.230 2.120 ;
        RECT 4.130 1.540 4.400 2.710 ;
        RECT 4.590 2.590 4.860 3.900 ;
        RECT 4.570 2.260 4.860 2.590 ;
        RECT 4.590 2.240 4.860 2.260 ;
        RECT 5.060 3.630 5.330 3.690 ;
        RECT 5.060 3.300 5.340 3.630 ;
        RECT 4.130 1.210 4.430 1.540 ;
        RECT 4.130 1.160 4.400 1.210 ;
        RECT 5.060 1.090 5.330 3.300 ;
        RECT 5.040 0.760 5.330 1.090 ;
        RECT 5.060 0.730 5.330 0.760 ;
        RECT 5.540 2.130 5.830 4.780 ;
        RECT 8.710 3.850 9.040 4.110 ;
        RECT 9.680 4.070 10.110 4.360 ;
        RECT 6.160 3.330 6.470 3.680 ;
        RECT 9.550 3.320 9.940 3.590 ;
        RECT 12.480 3.330 12.790 3.650 ;
        RECT 8.710 2.340 9.040 2.600 ;
        RECT 9.680 2.560 10.110 2.850 ;
        RECT 5.540 1.780 5.840 2.130 ;
        RECT 6.160 1.820 6.470 2.170 ;
        RECT 9.550 1.810 9.940 2.080 ;
        RECT 12.480 1.820 12.790 2.140 ;
        RECT 5.540 0.240 5.830 1.780 ;
        RECT 8.710 0.840 9.040 1.100 ;
        RECT 9.680 1.060 10.110 1.350 ;
        RECT 6.160 0.320 6.470 0.670 ;
        RECT 9.550 0.310 9.940 0.580 ;
        RECT 12.480 0.320 12.790 0.640 ;
      LAYER via ;
        RECT 3.660 5.500 3.930 5.770 ;
        RECT 0.110 4.870 0.370 5.130 ;
        RECT 1.940 4.880 2.200 5.140 ;
        RECT 4.590 5.310 4.860 5.580 ;
        RECT 8.750 5.360 9.010 5.620 ;
        RECT 9.740 5.610 10.000 5.870 ;
        RECT 3.660 4.420 3.930 4.690 ;
        RECT 4.130 4.820 4.400 5.090 ;
        RECT 0.110 3.360 0.370 3.620 ;
        RECT 1.940 3.370 2.200 3.630 ;
        RECT 5.520 4.810 5.810 5.100 ;
        RECT 6.190 4.870 6.450 5.130 ;
        RECT 9.610 4.830 9.870 5.090 ;
        RECT 12.510 4.870 12.770 5.130 ;
        RECT 4.570 3.900 4.840 4.170 ;
        RECT 4.120 2.740 4.390 3.010 ;
        RECT 0.110 1.850 0.370 2.110 ;
        RECT 1.940 1.860 2.200 2.120 ;
        RECT 4.570 2.290 4.840 2.560 ;
        RECT 5.070 3.330 5.340 3.600 ;
        RECT 8.750 3.850 9.010 4.110 ;
        RECT 9.740 4.100 10.000 4.360 ;
        RECT 5.560 3.300 5.820 3.560 ;
        RECT 6.190 3.360 6.450 3.620 ;
        RECT 9.610 3.320 9.870 3.580 ;
        RECT 12.510 3.360 12.770 3.620 ;
        RECT 4.160 1.240 4.430 1.510 ;
        RECT 5.040 0.790 5.310 1.060 ;
        RECT 8.750 2.340 9.010 2.600 ;
        RECT 9.740 2.590 10.000 2.850 ;
        RECT 5.550 1.810 5.840 2.100 ;
        RECT 6.190 1.850 6.450 2.110 ;
        RECT 9.610 1.810 9.870 2.070 ;
        RECT 12.510 1.850 12.770 2.110 ;
        RECT 8.750 0.840 9.010 1.100 ;
        RECT 9.740 1.090 10.000 1.350 ;
        RECT 5.540 0.270 5.830 0.560 ;
        RECT 6.190 0.350 6.450 0.610 ;
        RECT 9.610 0.310 9.870 0.570 ;
        RECT 12.510 0.350 12.770 0.610 ;
      LAYER met2 ;
        RECT 0.080 5.030 0.400 5.130 ;
        RECT 0.070 4.870 0.400 5.030 ;
        RECT 1.910 5.060 2.230 5.140 ;
        RECT 4.100 5.060 4.430 5.090 ;
        RECT 1.910 4.880 4.450 5.060 ;
        RECT 4.100 4.870 4.450 4.880 ;
        RECT 5.490 5.030 5.840 5.100 ;
        RECT 6.160 5.030 6.480 5.130 ;
        RECT 5.490 4.870 6.480 5.030 ;
        RECT 4.100 4.820 4.430 4.870 ;
        RECT 5.490 4.810 5.840 4.870 ;
        RECT 8.710 4.030 9.040 4.110 ;
        RECT 8.440 4.010 9.040 4.030 ;
        RECT 5.120 3.850 9.040 4.010 ;
        RECT 0.080 3.520 0.400 3.620 ;
        RECT 0.070 3.360 0.400 3.520 ;
        RECT 1.910 3.550 2.230 3.630 ;
        RECT 5.120 3.600 5.280 3.850 ;
        RECT 5.040 3.550 5.370 3.600 ;
        RECT 1.910 3.370 5.370 3.550 ;
        RECT 5.040 3.330 5.370 3.370 ;
        RECT 5.530 3.520 5.850 3.560 ;
        RECT 6.160 3.520 6.480 3.620 ;
        RECT 5.530 3.360 6.480 3.520 ;
        RECT 5.530 3.300 5.850 3.360 ;
        RECT 4.090 2.950 4.420 3.010 ;
        RECT 4.090 2.790 10.110 2.950 ;
        RECT 4.090 2.740 4.420 2.790 ;
        RECT 9.690 2.560 10.110 2.790 ;
        RECT 0.080 2.010 0.400 2.110 ;
        RECT 0.070 1.850 0.400 2.010 ;
        RECT 1.910 2.040 2.230 2.120 ;
        RECT 5.520 2.040 5.870 2.100 ;
        RECT 1.910 2.010 6.010 2.040 ;
        RECT 6.160 2.010 6.480 2.110 ;
        RECT 1.910 1.860 6.480 2.010 ;
        RECT 5.520 1.850 6.480 1.860 ;
        RECT 5.520 1.810 5.870 1.850 ;
        RECT 4.130 1.450 4.460 1.510 ;
        RECT 4.130 1.290 10.110 1.450 ;
        RECT 4.130 1.240 4.460 1.290 ;
        RECT 5.010 1.000 5.340 1.060 ;
        RECT 8.710 1.020 9.040 1.100 ;
        RECT 9.690 1.060 10.110 1.290 ;
        RECT 8.440 1.000 9.040 1.020 ;
        RECT 5.010 0.840 9.040 1.000 ;
        RECT 5.010 0.790 5.340 0.840 ;
        RECT 5.510 0.510 5.860 0.560 ;
        RECT 6.160 0.510 6.480 0.610 ;
        RECT 5.510 0.350 6.480 0.510 ;
        RECT 5.510 0.270 5.860 0.350 ;
  END
END sky130_hilas_VinjDecode2to4

MACRO sky130_hilas_TA2Cell_1FG
  CLASS CORE ;
  FOREIGN sky130_hilas_TA2Cell_1FG ;
  ORIGIN 0.000 0.000 ;
  SIZE 34.530 BY 10.100 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 13.570 1.300 14.050 1.310 ;
        RECT 13.570 1.060 14.460 1.300 ;
    END
  END VIN12
  PIN VIN11
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 13.620 4.820 14.460 5.020 ;
    END
  END VIN11
  PIN VIN21
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 28.360 3.390 29.020 3.400 ;
        RECT 28.360 3.160 29.460 3.390 ;
        RECT 28.820 2.960 29.130 3.160 ;
    END
  END VIN21
  PIN VIN22
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 28.780 6.080 29.090 6.240 ;
        RECT 28.350 6.070 29.230 6.080 ;
        RECT 28.280 5.830 29.230 6.070 ;
    END
  END VIN22
  PIN VPWR
    USE ANALOG ;
    ANTENNAGATEAREA 0.408000 ;
    ANTENNADIFFAREA 0.302000 ;
    PORT
      LAYER met2 ;
        RECT 31.750 6.020 32.060 6.250 ;
        RECT 34.000 6.020 34.310 6.270 ;
        RECT 31.620 5.940 34.310 6.020 ;
        RECT 31.620 5.790 34.160 5.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.520 0.050 31.790 0.260 ;
    END
  END VPWR
  PIN VGND
    USE ANALOG ;
    ANTENNAGATEAREA 0.360000 ;
    ANTENNADIFFAREA 1.574400 ;
    PORT
      LAYER nwell ;
        RECT 28.330 6.100 31.640 10.020 ;
        RECT 27.680 6.090 32.810 6.100 ;
        RECT 28.330 5.920 32.810 6.090 ;
        RECT 28.330 3.870 31.640 5.920 ;
      LAYER met2 ;
        RECT 30.250 7.110 30.570 7.370 ;
        RECT 30.290 7.090 31.470 7.110 ;
        RECT 30.290 6.830 31.510 7.090 ;
        RECT 30.290 6.770 31.470 6.830 ;
        RECT 30.250 6.760 31.470 6.770 ;
        RECT 30.250 6.510 30.570 6.760 ;
    END
    PORT
      LAYER met2 ;
        RECT 18.900 0.400 19.220 0.410 ;
        RECT 29.340 0.400 29.670 0.540 ;
        RECT 18.900 0.240 29.670 0.400 ;
        RECT 18.900 0.230 19.590 0.240 ;
        RECT 18.900 0.110 19.220 0.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.190 6.010 13.420 6.090 ;
    END
    PORT
      LAYER met1 ;
        RECT 18.980 6.010 19.210 6.100 ;
    END
  END VGND
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 4.960 5.930 5.280 6.050 ;
        RECT 27.160 5.930 27.480 6.050 ;
        RECT 4.960 5.750 27.480 5.930 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.160 0.050 27.440 0.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.960 6.050 5.240 6.100 ;
        RECT 4.960 5.770 5.280 6.050 ;
      LAYER via ;
        RECT 4.990 5.780 5.250 6.040 ;
    END
  END VINJ
  PIN OUTPUT1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 32.700 3.390 32.810 3.620 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 32.700 2.570 32.810 2.790 ;
    END
  END OUTPUT2
  PIN DRAIN1
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 2.640 5.690 2.950 5.910 ;
        RECT 0.760 5.480 12.290 5.690 ;
        RECT 2.070 5.470 12.290 5.480 ;
        RECT 4.720 5.420 4.790 5.470 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 4.720 0.550 4.800 0.730 ;
    END
  END DRAIN2
  PIN COLSEL2
    PORT
      LAYER met1 ;
        RECT 5.490 6.040 5.680 6.100 ;
    END
  END COLSEL2
  PIN GATE2
    PORT
      LAYER met1 ;
        RECT 11.970 6.010 12.200 6.090 ;
    END
  END GATE2
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT 20.200 6.020 20.430 6.100 ;
    END
  END GATE1
  PIN COLSEL1
    PORT
      LAYER met1 ;
        RECT 26.720 6.020 26.910 6.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 26.720 0.050 26.910 0.100 ;
    END
  END COLSEL1
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 15.480 5.940 16.920 6.100 ;
    END
  END VTUN
  OBS
      LAYER nwell ;
        RECT 0.760 3.870 4.070 10.020 ;
        RECT 5.800 7.580 8.520 9.230 ;
        RECT 5.810 7.540 8.520 7.580 ;
        RECT 5.810 6.210 8.520 6.250 ;
        RECT 5.800 6.100 8.520 6.210 ;
        RECT 4.720 6.090 8.520 6.100 ;
        RECT 4.720 5.420 4.790 5.600 ;
        RECT 5.800 4.560 8.520 6.090 ;
        RECT 11.140 5.320 11.700 7.740 ;
        RECT 20.700 5.320 21.260 7.740 ;
        RECT 23.880 7.580 26.600 9.230 ;
        RECT 23.880 7.540 26.590 7.580 ;
        RECT 23.880 6.210 26.590 6.250 ;
        RECT 23.880 4.560 26.600 6.210 ;
        RECT 29.010 3.160 29.460 3.390 ;
        RECT 27.670 3.030 29.530 3.100 ;
        RECT 4.720 0.550 4.800 0.730 ;
        RECT 31.300 0.000 33.160 1.650 ;
        RECT 33.250 0.500 34.530 6.180 ;
      LAYER li1 ;
        RECT 1.160 9.290 1.360 9.640 ;
        RECT 2.640 9.390 3.170 9.560 ;
        RECT 1.150 9.260 1.360 9.290 ;
        RECT 1.150 8.680 1.370 9.260 ;
        RECT 1.150 8.670 1.360 8.680 ;
        RECT 1.530 8.500 1.720 8.510 ;
        RECT 1.520 8.210 1.720 8.500 ;
        RECT 1.440 7.880 1.730 8.210 ;
        RECT 1.920 7.400 2.090 9.010 ;
        RECT 2.750 8.630 2.920 9.000 ;
        RECT 5.360 8.960 10.420 9.790 ;
        RECT 29.230 9.390 29.760 9.560 ;
        RECT 31.040 9.290 31.240 9.640 ;
        RECT 31.040 9.260 31.250 9.290 ;
        RECT 9.870 8.880 10.350 8.960 ;
        RECT 9.870 8.780 10.200 8.880 ;
        RECT 2.620 8.590 2.940 8.630 ;
        RECT 2.610 8.400 2.940 8.590 ;
        RECT 2.620 8.370 2.940 8.400 ;
        RECT 1.910 7.210 2.090 7.400 ;
        RECT 2.750 7.310 2.920 8.370 ;
        RECT 7.990 8.020 8.220 8.710 ;
        RECT 9.870 8.630 10.020 8.780 ;
        RECT 24.180 8.020 24.410 8.710 ;
        RECT 29.480 8.630 29.650 9.000 ;
        RECT 29.460 8.590 29.780 8.630 ;
        RECT 29.460 8.400 29.790 8.590 ;
        RECT 29.460 8.370 29.780 8.400 ;
        RECT 9.060 7.080 9.250 7.400 ;
        RECT 23.150 7.080 23.340 7.400 ;
        RECT 29.480 7.310 29.650 8.370 ;
        RECT 30.310 7.400 30.480 9.010 ;
        RECT 31.030 8.680 31.250 9.260 ;
        RECT 31.040 8.670 31.250 8.680 ;
        RECT 30.680 8.500 30.870 8.510 ;
        RECT 30.680 8.210 30.880 8.500 ;
        RECT 30.670 7.880 30.960 8.210 ;
        RECT 30.310 7.210 30.490 7.400 ;
        RECT 9.060 6.990 9.340 7.080 ;
        RECT 5.700 6.850 9.340 6.990 ;
        RECT 23.060 6.990 23.340 7.080 ;
        RECT 23.060 6.850 26.700 6.990 ;
        RECT 5.700 6.810 9.250 6.850 ;
        RECT 1.910 6.490 2.090 6.680 ;
        RECT 1.440 5.680 1.730 6.010 ;
        RECT 1.520 5.390 1.720 5.680 ;
        RECT 1.530 5.380 1.720 5.390 ;
        RECT 1.150 5.210 1.360 5.220 ;
        RECT 1.150 4.630 1.370 5.210 ;
        RECT 1.920 4.880 2.090 6.490 ;
        RECT 2.750 5.870 2.920 6.580 ;
        RECT 9.060 6.390 9.250 6.810 ;
        RECT 23.150 6.810 26.700 6.850 ;
        RECT 23.150 6.390 23.340 6.810 ;
        RECT 28.760 6.160 29.080 6.200 ;
        RECT 28.750 6.100 29.080 6.160 ;
        RECT 28.660 5.940 29.080 6.100 ;
        RECT 2.620 5.830 2.940 5.870 ;
        RECT 2.610 5.640 2.940 5.830 ;
        RECT 2.620 5.610 2.940 5.640 ;
        RECT 2.750 4.890 2.920 5.610 ;
        RECT 7.990 5.080 8.220 5.810 ;
        RECT 9.910 5.310 10.230 5.350 ;
        RECT 9.900 5.120 10.230 5.310 ;
        RECT 9.910 5.090 10.230 5.120 ;
        RECT 10.030 4.950 10.050 5.090 ;
        RECT 24.180 5.080 24.410 5.810 ;
        RECT 28.660 5.790 28.900 5.940 ;
        RECT 29.480 5.870 29.650 6.580 ;
        RECT 30.310 6.490 30.490 6.680 ;
        RECT 29.460 5.830 29.780 5.870 ;
        RECT 28.660 5.770 28.830 5.790 ;
        RECT 29.460 5.640 29.790 5.830 ;
        RECT 29.460 5.610 29.780 5.640 ;
        RECT 28.910 5.330 29.230 5.370 ;
        RECT 28.900 5.140 29.230 5.330 ;
        RECT 28.910 5.110 29.230 5.140 ;
        RECT 10.030 4.870 10.380 4.950 ;
        RECT 29.480 4.890 29.650 5.610 ;
        RECT 30.310 4.880 30.480 6.490 ;
        RECT 31.760 6.170 32.080 6.210 ;
        RECT 34.010 6.190 34.330 6.230 ;
        RECT 30.670 5.680 30.960 6.010 ;
        RECT 31.760 5.980 32.090 6.170 ;
        RECT 34.010 6.120 34.340 6.190 ;
        RECT 31.760 5.950 32.080 5.980 ;
        RECT 31.850 5.770 32.050 5.950 ;
        RECT 30.680 5.390 30.880 5.680 ;
        RECT 31.710 5.520 32.030 5.560 ;
        RECT 30.680 5.380 30.870 5.390 ;
        RECT 31.040 5.210 31.250 5.220 ;
        RECT 1.150 4.600 1.360 4.630 ;
        RECT 1.160 4.250 1.360 4.600 ;
        RECT 2.640 4.330 3.170 4.500 ;
        RECT 5.330 4.020 10.380 4.870 ;
        RECT 31.030 4.630 31.250 5.210 ;
        RECT 31.440 5.120 31.610 5.450 ;
        RECT 31.710 5.440 32.040 5.520 ;
        RECT 31.710 5.300 32.050 5.440 ;
        RECT 31.850 5.110 32.050 5.300 ;
        RECT 32.440 5.110 32.990 6.100 ;
        RECT 33.810 5.950 34.440 6.120 ;
        RECT 33.810 5.670 34.170 5.950 ;
        RECT 33.460 5.500 34.170 5.670 ;
        RECT 33.460 4.830 34.160 5.060 ;
        RECT 31.040 4.600 31.250 4.630 ;
        RECT 33.410 4.600 34.160 4.830 ;
        RECT 28.100 4.510 28.420 4.540 ;
        RECT 28.100 4.320 28.430 4.510 ;
        RECT 29.230 4.330 29.760 4.500 ;
        RECT 28.100 4.280 28.420 4.320 ;
        RECT 31.040 4.250 31.240 4.600 ;
        RECT 31.440 4.260 31.610 4.590 ;
        RECT 31.850 4.410 32.050 4.600 ;
        RECT 31.710 4.270 32.050 4.410 ;
        RECT 31.710 4.190 32.040 4.270 ;
        RECT 31.710 4.150 32.030 4.190 ;
        RECT 31.850 3.760 32.050 3.940 ;
        RECT 31.760 3.730 32.080 3.760 ;
        RECT 13.210 2.520 13.410 3.530 ;
        RECT 18.960 2.520 19.250 3.530 ;
        RECT 28.080 2.560 28.260 3.620 ;
        RECT 31.760 3.540 32.090 3.730 ;
        RECT 32.440 3.610 32.990 4.600 ;
        RECT 33.460 4.180 34.160 4.600 ;
        RECT 34.060 3.970 34.380 4.010 ;
        RECT 34.060 3.780 34.390 3.970 ;
        RECT 34.060 3.760 34.380 3.780 ;
        RECT 33.450 3.750 34.380 3.760 ;
        RECT 33.450 3.580 34.150 3.750 ;
        RECT 31.760 3.500 32.080 3.540 ;
        RECT 28.830 3.230 29.150 3.260 ;
        RECT 34.050 3.250 34.370 3.290 ;
        RECT 28.830 3.160 29.160 3.230 ;
        RECT 28.690 3.070 29.160 3.160 ;
        RECT 28.640 3.040 29.160 3.070 ;
        RECT 31.760 3.170 32.080 3.210 ;
        RECT 28.640 3.000 29.150 3.040 ;
        RECT 28.640 2.900 28.860 3.000 ;
        RECT 31.760 2.980 32.090 3.170 ;
        RECT 34.050 3.100 34.380 3.250 ;
        RECT 31.760 2.950 32.080 2.980 ;
        RECT 28.640 2.740 28.810 2.900 ;
        RECT 31.850 2.770 32.050 2.950 ;
        RECT 31.710 2.520 32.030 2.560 ;
        RECT 29.130 2.400 29.210 2.480 ;
        RECT 29.270 2.400 29.460 2.520 ;
        RECT 29.130 2.310 29.460 2.400 ;
        RECT 29.270 2.290 29.460 2.310 ;
        RECT 31.440 2.120 31.610 2.450 ;
        RECT 31.710 2.440 32.040 2.520 ;
        RECT 31.710 2.300 32.050 2.440 ;
        RECT 31.850 2.110 32.050 2.300 ;
        RECT 32.440 2.110 32.990 3.100 ;
        RECT 33.450 3.060 34.380 3.100 ;
        RECT 33.450 3.030 34.370 3.060 ;
        RECT 33.450 2.920 34.150 3.030 ;
        RECT 33.460 2.240 34.160 2.500 ;
        RECT 33.410 2.010 34.160 2.240 ;
        RECT 33.460 1.620 34.160 2.010 ;
        RECT 31.440 1.260 31.610 1.590 ;
        RECT 31.850 1.410 32.050 1.600 ;
        RECT 31.710 1.270 32.050 1.410 ;
        RECT 31.710 1.190 32.040 1.270 ;
        RECT 31.710 1.150 32.030 1.190 ;
        RECT 31.710 0.940 31.890 1.150 ;
        RECT 31.710 0.760 32.050 0.940 ;
        RECT 31.710 0.730 32.080 0.760 ;
        RECT 31.710 0.540 32.090 0.730 ;
        RECT 32.440 0.610 32.990 1.600 ;
        RECT 33.460 1.040 34.170 1.180 ;
        RECT 33.460 1.010 34.290 1.040 ;
        RECT 33.810 1.000 34.290 1.010 ;
        RECT 33.810 0.810 34.300 1.000 ;
        RECT 33.810 0.780 34.290 0.810 ;
        RECT 33.810 0.730 34.170 0.780 ;
        RECT 31.710 0.500 32.080 0.540 ;
        RECT 31.710 0.000 31.890 0.500 ;
        RECT 32.520 0.000 32.690 0.610 ;
        RECT 33.810 0.560 34.440 0.730 ;
      LAYER mcon ;
        RECT 2.990 9.390 3.170 9.560 ;
        RECT 1.180 9.090 1.350 9.260 ;
        RECT 1.530 8.250 1.710 8.440 ;
        RECT 31.050 9.090 31.220 9.260 ;
        RECT 9.970 8.820 10.140 8.990 ;
        RECT 2.710 8.410 2.880 8.580 ;
        RECT 8.020 8.510 8.190 8.680 ;
        RECT 8.020 8.060 8.190 8.230 ;
        RECT 24.210 8.510 24.380 8.680 ;
        RECT 29.520 8.410 29.690 8.580 ;
        RECT 24.210 8.060 24.380 8.230 ;
        RECT 30.690 8.250 30.870 8.440 ;
        RECT 9.160 6.880 9.330 7.050 ;
        RECT 23.070 6.880 23.240 7.050 ;
        RECT 1.530 5.450 1.710 5.640 ;
        RECT 28.850 5.980 29.020 6.150 ;
        RECT 2.710 5.650 2.880 5.820 ;
        RECT 8.020 5.560 8.190 5.730 ;
        RECT 24.210 5.560 24.380 5.730 ;
        RECT 29.520 5.650 29.690 5.820 ;
        RECT 8.020 5.110 8.190 5.280 ;
        RECT 10.000 5.130 10.170 5.300 ;
        RECT 24.210 5.110 24.380 5.280 ;
        RECT 29.000 5.150 29.170 5.320 ;
        RECT 31.820 5.990 31.990 6.160 ;
        RECT 30.690 5.450 30.870 5.640 ;
        RECT 32.760 5.600 32.930 5.770 ;
        RECT 34.070 6.010 34.240 6.180 ;
        RECT 1.180 4.630 1.350 4.800 ;
        RECT 2.990 4.330 3.170 4.500 ;
        RECT 31.770 5.340 31.940 5.510 ;
        RECT 31.050 4.630 31.220 4.800 ;
        RECT 33.420 4.630 33.590 4.800 ;
        RECT 28.160 4.330 28.330 4.500 ;
        RECT 31.770 4.200 31.940 4.370 ;
        RECT 32.760 3.940 32.930 4.110 ;
        RECT 13.220 3.290 13.390 3.460 ;
        RECT 13.230 2.570 13.400 2.740 ;
        RECT 19.010 3.290 19.180 3.460 ;
        RECT 19.010 2.570 19.180 2.740 ;
        RECT 31.820 3.550 31.990 3.720 ;
        RECT 34.120 3.790 34.290 3.960 ;
        RECT 28.890 3.050 29.060 3.220 ;
        RECT 31.820 2.990 31.990 3.160 ;
        RECT 34.110 3.070 34.280 3.240 ;
        RECT 32.760 2.600 32.930 2.770 ;
        RECT 29.280 2.320 29.450 2.490 ;
        RECT 31.770 2.340 31.940 2.510 ;
        RECT 33.420 2.040 33.590 2.210 ;
        RECT 31.770 1.200 31.940 1.370 ;
        RECT 32.760 0.940 32.930 1.110 ;
        RECT 31.820 0.550 31.990 0.720 ;
        RECT 34.030 0.820 34.200 0.990 ;
      LAYER met1 ;
        RECT 1.000 9.320 1.280 9.970 ;
        RECT 1.000 8.720 1.390 9.320 ;
        RECT 1.000 5.170 1.280 8.720 ;
        RECT 1.530 8.510 1.720 9.970 ;
        RECT 2.930 9.150 3.240 9.590 ;
        RECT 8.010 8.760 8.240 9.970 ;
        RECT 9.230 9.000 9.460 9.970 ;
        RECT 1.500 8.480 1.720 8.510 ;
        RECT 1.490 8.210 1.740 8.480 ;
        RECT 2.630 8.340 2.950 8.660 ;
        RECT 1.490 8.200 1.730 8.210 ;
        RECT 1.500 7.960 1.730 8.200 ;
        RECT 7.980 7.970 8.240 8.760 ;
        RECT 9.220 8.750 9.460 9.000 ;
        RECT 9.890 8.750 10.210 9.070 ;
        RECT 1.530 5.930 1.690 7.960 ;
        RECT 1.880 7.400 2.120 7.530 ;
        RECT 1.860 7.080 2.120 7.400 ;
        RECT 1.860 6.480 2.120 6.800 ;
        RECT 1.880 6.360 2.120 6.480 ;
        RECT 1.500 5.690 1.730 5.930 ;
        RECT 1.490 5.680 1.730 5.690 ;
        RECT 1.490 5.410 1.740 5.680 ;
        RECT 2.630 5.580 2.950 5.900 ;
        RECT 8.010 5.820 8.240 7.970 ;
        RECT 9.230 7.110 9.460 8.750 ;
        RECT 9.130 6.820 9.460 7.110 ;
        RECT 1.500 5.380 1.720 5.410 ;
        RECT 1.000 4.570 1.390 5.170 ;
        RECT 1.000 3.920 1.280 4.570 ;
        RECT 1.530 3.920 1.720 5.380 ;
        RECT 7.980 5.030 8.240 5.820 ;
        RECT 2.930 4.300 3.240 4.740 ;
        RECT 8.010 3.920 8.240 5.030 ;
        RECT 9.230 3.920 9.460 6.820 ;
        RECT 9.920 5.060 10.240 5.380 ;
        RECT 11.520 3.930 11.940 9.970 ;
        RECT 20.460 3.920 20.880 9.970 ;
        RECT 22.940 7.110 23.170 9.970 ;
        RECT 24.160 8.760 24.390 9.970 ;
        RECT 29.160 9.150 29.470 9.590 ;
        RECT 24.160 7.970 24.420 8.760 ;
        RECT 29.450 8.340 29.770 8.660 ;
        RECT 30.680 8.510 30.870 9.970 ;
        RECT 31.120 9.320 31.400 9.970 ;
        RECT 31.010 8.720 31.400 9.320 ;
        RECT 30.680 8.480 30.900 8.510 ;
        RECT 30.660 8.210 30.910 8.480 ;
        RECT 30.670 8.200 30.910 8.210 ;
        RECT 22.940 6.820 23.270 7.110 ;
        RECT 22.940 3.920 23.170 6.820 ;
        RECT 24.160 5.820 24.390 7.970 ;
        RECT 30.670 7.960 30.900 8.200 ;
        RECT 30.280 7.400 30.520 7.530 ;
        RECT 30.280 7.080 30.540 7.400 ;
        RECT 30.280 6.480 30.540 6.800 ;
        RECT 30.280 6.360 30.520 6.480 ;
        RECT 27.160 6.050 27.440 6.100 ;
        RECT 24.160 5.030 24.420 5.820 ;
        RECT 27.160 5.750 27.480 6.050 ;
        RECT 28.770 5.910 29.090 6.230 ;
        RECT 30.710 6.100 30.870 7.960 ;
        RECT 31.120 7.120 31.400 8.720 ;
        RECT 31.120 6.800 31.480 7.120 ;
        RECT 31.120 6.100 31.400 6.800 ;
        RECT 31.750 6.100 32.070 6.240 ;
        RECT 30.710 5.960 31.400 6.100 ;
        RECT 30.710 5.930 30.870 5.960 ;
        RECT 29.450 5.580 29.770 5.900 ;
        RECT 30.670 5.690 30.900 5.930 ;
        RECT 30.670 5.680 30.910 5.690 ;
        RECT 30.660 5.410 30.910 5.680 ;
        RECT 28.920 5.080 29.240 5.400 ;
        RECT 30.680 5.380 30.900 5.410 ;
        RECT 24.160 3.920 24.390 5.030 ;
        RECT 28.090 4.250 28.410 4.570 ;
        RECT 29.160 4.300 29.470 4.740 ;
        RECT 29.170 4.240 29.380 4.300 ;
        RECT 29.150 3.920 29.410 4.240 ;
        RECT 30.680 3.920 30.870 5.380 ;
        RECT 31.120 5.170 31.400 5.960 ;
        RECT 31.510 5.950 32.070 6.100 ;
        RECT 31.750 5.920 32.070 5.950 ;
        RECT 32.570 5.830 32.910 6.220 ;
        RECT 31.700 5.270 32.020 5.590 ;
        RECT 32.570 5.540 32.960 5.830 ;
        RECT 31.010 4.570 31.400 5.170 ;
        RECT 31.120 3.920 31.400 4.570 ;
        RECT 31.700 4.120 32.020 4.440 ;
        RECT 32.570 4.170 32.910 5.540 ;
        RECT 33.240 4.860 33.510 6.210 ;
        RECT 34.000 5.940 34.320 6.260 ;
        RECT 33.240 4.570 33.620 4.860 ;
        RECT 13.220 3.280 13.390 3.460 ;
        RECT 19.010 3.280 19.180 3.460 ;
        RECT 13.200 2.690 13.520 2.990 ;
        RECT 28.820 2.970 29.140 3.290 ;
        RECT 13.200 2.580 13.440 2.690 ;
        RECT 18.900 2.620 19.220 2.940 ;
        RECT 13.230 2.570 13.400 2.580 ;
        RECT 13.420 2.520 13.440 2.580 ;
        RECT 19.010 2.570 19.180 2.620 ;
        RECT 29.170 2.580 29.380 3.920 ;
        RECT 32.570 3.880 32.960 4.170 ;
        RECT 31.750 3.470 32.070 3.790 ;
        RECT 31.750 2.920 32.070 3.240 ;
        RECT 32.570 2.830 32.910 3.880 ;
        RECT 29.250 2.260 29.480 2.550 ;
        RECT 31.700 2.270 32.020 2.590 ;
        RECT 32.570 2.540 32.960 2.830 ;
        RECT 31.700 1.120 32.020 1.440 ;
        RECT 32.570 1.170 32.910 2.540 ;
        RECT 33.240 2.270 33.510 4.570 ;
        RECT 34.050 3.720 34.370 4.040 ;
        RECT 34.040 3.000 34.360 3.320 ;
        RECT 33.240 1.980 33.620 2.270 ;
        RECT 32.570 0.880 32.960 1.170 ;
        RECT 18.900 0.110 19.220 0.410 ;
        RECT 29.340 0.250 29.670 0.540 ;
        RECT 31.750 0.470 32.070 0.790 ;
        RECT 32.570 0.500 32.910 0.880 ;
        RECT 33.240 0.510 33.510 1.980 ;
        RECT 33.960 0.750 34.280 1.070 ;
        RECT 29.330 0.220 29.750 0.250 ;
        RECT 30.350 0.240 30.850 0.250 ;
        RECT 30.350 0.220 31.190 0.240 ;
        RECT 29.330 0.110 31.190 0.220 ;
        RECT 29.610 0.080 30.510 0.110 ;
        RECT 30.850 0.050 31.190 0.110 ;
      LAYER via ;
        RECT 2.950 9.180 3.210 9.440 ;
        RECT 2.660 8.370 2.920 8.630 ;
        RECT 9.920 8.780 10.180 9.040 ;
        RECT 1.860 7.110 2.120 7.370 ;
        RECT 1.860 6.510 2.120 6.770 ;
        RECT 2.660 5.610 2.920 5.870 ;
        RECT 2.950 4.450 3.210 4.710 ;
        RECT 9.950 5.090 10.210 5.350 ;
        RECT 29.190 9.180 29.450 9.440 ;
        RECT 29.480 8.370 29.740 8.630 ;
        RECT 30.280 7.110 30.540 7.370 ;
        RECT 30.280 6.510 30.540 6.770 ;
        RECT 27.190 5.770 27.450 6.030 ;
        RECT 28.800 5.940 29.060 6.200 ;
        RECT 31.220 6.830 31.480 7.090 ;
        RECT 29.480 5.610 29.740 5.870 ;
        RECT 28.950 5.110 29.210 5.370 ;
        RECT 28.120 4.280 28.380 4.540 ;
        RECT 29.190 4.450 29.450 4.710 ;
        RECT 29.150 3.950 29.410 4.210 ;
        RECT 31.780 5.950 32.040 6.210 ;
        RECT 31.730 5.300 31.990 5.560 ;
        RECT 31.730 4.150 31.990 4.410 ;
        RECT 34.030 5.970 34.290 6.230 ;
        RECT 28.850 3.000 29.110 3.260 ;
        RECT 13.230 2.710 13.490 2.970 ;
        RECT 18.930 2.650 19.190 2.910 ;
        RECT 31.780 3.500 32.040 3.760 ;
        RECT 31.780 2.950 32.040 3.210 ;
        RECT 31.730 2.300 31.990 2.560 ;
        RECT 31.730 1.150 31.990 1.410 ;
        RECT 34.080 3.750 34.340 4.010 ;
        RECT 34.070 3.030 34.330 3.290 ;
        RECT 18.930 0.130 19.190 0.390 ;
        RECT 29.370 0.260 29.640 0.520 ;
        RECT 31.780 0.500 32.040 0.760 ;
        RECT 33.990 0.780 34.250 1.040 ;
      LAYER met2 ;
        RECT 2.930 9.470 3.240 9.480 ;
        RECT 29.160 9.470 29.470 9.480 ;
        RECT 0.760 9.290 12.290 9.470 ;
        RECT 20.110 9.290 31.640 9.470 ;
        RECT 2.930 9.150 3.240 9.290 ;
        RECT 29.160 9.150 29.470 9.290 ;
        RECT 9.900 8.880 10.210 9.080 ;
        RECT 9.900 8.870 10.500 8.880 ;
        RECT 9.900 8.750 12.290 8.870 ;
        RECT 10.040 8.710 12.290 8.750 ;
        RECT 10.350 8.690 12.290 8.710 ;
        RECT 2.640 8.450 2.950 8.670 ;
        RECT 0.760 8.440 2.950 8.450 ;
        RECT 29.450 8.450 29.760 8.670 ;
        RECT 0.760 8.230 12.290 8.440 ;
        RECT 29.450 8.340 31.640 8.450 ;
        RECT 29.610 8.230 31.640 8.340 ;
        RECT 2.070 8.220 12.290 8.230 ;
        RECT 1.830 7.250 12.290 7.470 ;
        RECT 1.830 7.110 2.150 7.250 ;
        RECT 1.850 6.770 2.110 7.110 ;
        RECT 1.830 6.510 2.150 6.770 ;
        RECT 29.450 5.690 29.760 5.910 ;
        RECT 29.450 5.580 31.640 5.690 ;
        RECT 29.600 5.480 31.640 5.580 ;
        RECT 9.930 5.060 10.240 5.390 ;
        RECT 28.930 5.220 29.240 5.410 ;
        RECT 10.340 4.950 12.290 5.160 ;
        RECT 28.890 4.970 29.610 5.220 ;
        RECT 31.260 5.160 31.590 5.370 ;
        RECT 31.700 5.270 32.010 5.600 ;
        RECT 29.340 4.860 29.610 4.970 ;
        RECT 2.930 4.600 3.240 4.740 ;
        RECT 0.760 4.590 3.240 4.600 ;
        RECT 29.160 4.600 29.470 4.740 ;
        RECT 29.160 4.590 31.640 4.600 ;
        RECT 0.760 4.440 12.290 4.590 ;
        RECT 20.110 4.570 31.640 4.590 ;
        RECT 14.070 4.440 31.640 4.570 ;
        RECT 0.760 4.420 3.240 4.440 ;
        RECT 2.930 4.410 3.240 4.420 ;
        RECT 14.070 4.350 24.210 4.440 ;
        RECT 27.600 4.360 27.950 4.440 ;
        RECT 14.020 3.380 23.030 3.600 ;
        RECT 13.200 2.940 13.520 2.990 ;
        RECT 13.200 2.690 19.220 2.940 ;
        RECT 18.900 2.620 19.220 2.690 ;
        RECT 14.070 1.600 19.730 1.820 ;
        RECT 19.510 1.270 19.730 1.600 ;
        RECT 22.810 1.770 23.030 3.380 ;
        RECT 23.990 3.150 24.210 4.350 ;
        RECT 28.090 4.240 28.400 4.440 ;
        RECT 29.160 4.420 31.640 4.440 ;
        RECT 29.160 4.410 29.470 4.420 ;
        RECT 31.260 4.340 31.590 4.420 ;
        RECT 29.410 4.290 29.610 4.300 ;
        RECT 29.410 4.210 29.630 4.290 ;
        RECT 29.120 4.190 29.630 4.210 ;
        RECT 29.070 3.950 29.630 4.190 ;
        RECT 31.700 4.110 32.010 4.440 ;
        RECT 29.070 3.940 29.540 3.950 ;
        RECT 34.050 3.880 34.360 4.050 ;
        RECT 31.880 3.790 34.530 3.880 ;
        RECT 31.750 3.650 34.530 3.790 ;
        RECT 31.750 3.460 32.060 3.650 ;
        RECT 23.960 3.110 24.210 3.150 ;
        RECT 23.960 2.470 24.220 3.110 ;
        RECT 31.750 3.050 32.060 3.250 ;
        RECT 34.040 3.050 34.350 3.330 ;
        RECT 31.620 2.830 34.530 3.050 ;
        RECT 23.960 2.260 28.090 2.470 ;
        RECT 27.880 2.120 28.090 2.260 ;
        RECT 31.260 2.160 31.590 2.370 ;
        RECT 31.700 2.270 32.010 2.600 ;
        RECT 27.880 1.910 29.900 2.120 ;
        RECT 22.810 1.550 25.660 1.770 ;
        RECT 31.260 1.340 31.590 1.550 ;
        RECT 23.880 1.270 29.900 1.320 ;
        RECT 19.510 1.110 29.900 1.270 ;
        RECT 31.700 1.110 32.010 1.440 ;
        RECT 19.510 1.050 24.270 1.110 ;
        RECT 33.960 0.890 34.270 1.080 ;
        RECT 31.610 0.660 34.320 0.890 ;
        RECT 31.750 0.460 32.060 0.660 ;
  END
END sky130_hilas_TA2Cell_1FG

MACRO sky130_hilas_swc4x1cellOverlap
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x1cellOverlap ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 10.360 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 4.870 6.420 7.590 6.650 ;
        RECT 0.010 2.660 1.740 4.500 ;
        RECT 4.870 3.560 10.080 6.420 ;
        RECT 14.520 4.310 16.250 10.360 ;
        RECT 4.860 0.260 10.080 3.560 ;
        RECT 4.860 0.060 7.580 0.260 ;
      LAYER li1 ;
        RECT 5.270 5.080 7.220 6.250 ;
        RECT 7.620 5.950 7.940 5.960 ;
        RECT 7.620 5.780 8.200 5.950 ;
        RECT 7.620 5.730 7.950 5.780 ;
        RECT 7.620 5.700 7.940 5.730 ;
        RECT 9.480 5.680 9.680 6.030 ;
        RECT 7.620 5.370 7.940 5.410 ;
        RECT 7.620 5.330 7.950 5.370 ;
        RECT 7.620 5.160 8.200 5.330 ;
        RECT 7.620 5.150 7.940 5.160 ;
        RECT 8.750 5.060 8.950 5.660 ;
        RECT 9.480 5.650 9.690 5.680 ;
        RECT 9.470 5.060 9.690 5.650 ;
        RECT 5.270 3.550 7.220 4.720 ;
        RECT 7.620 4.520 7.940 4.530 ;
        RECT 7.620 4.350 8.200 4.520 ;
        RECT 7.620 4.310 7.950 4.350 ;
        RECT 7.620 4.270 7.940 4.310 ;
        RECT 8.750 4.020 8.950 4.620 ;
        RECT 9.470 4.030 9.690 4.620 ;
        RECT 9.480 4.000 9.690 4.030 ;
        RECT 7.620 3.950 7.940 3.980 ;
        RECT 7.620 3.900 7.950 3.950 ;
        RECT 7.620 3.730 8.200 3.900 ;
        RECT 7.620 3.720 7.940 3.730 ;
        RECT 9.480 3.650 9.680 4.000 ;
        RECT 0.430 3.110 0.980 3.540 ;
        RECT 8.870 3.250 9.310 3.420 ;
        RECT 5.260 1.990 7.210 3.160 ;
        RECT 7.620 2.940 7.940 2.950 ;
        RECT 7.620 2.770 8.200 2.940 ;
        RECT 7.620 2.720 7.950 2.770 ;
        RECT 7.620 2.690 7.940 2.720 ;
        RECT 9.480 2.670 9.680 3.020 ;
        RECT 7.620 2.360 7.940 2.400 ;
        RECT 7.620 2.320 7.950 2.360 ;
        RECT 7.620 2.150 8.200 2.320 ;
        RECT 7.620 2.140 7.940 2.150 ;
        RECT 8.750 2.050 8.950 2.650 ;
        RECT 9.480 2.640 9.690 2.670 ;
        RECT 9.470 2.050 9.690 2.640 ;
        RECT 5.260 0.450 7.210 1.620 ;
        RECT 7.620 1.520 7.940 1.530 ;
        RECT 7.620 1.350 8.200 1.520 ;
        RECT 7.620 1.310 7.950 1.350 ;
        RECT 7.620 1.270 7.940 1.310 ;
        RECT 8.750 1.020 8.950 1.620 ;
        RECT 9.470 1.030 9.690 1.620 ;
        RECT 9.480 1.000 9.690 1.030 ;
        RECT 7.620 0.950 7.940 0.980 ;
        RECT 7.620 0.900 7.950 0.950 ;
        RECT 7.620 0.730 8.200 0.900 ;
        RECT 7.620 0.720 7.940 0.730 ;
        RECT 9.480 0.650 9.680 1.000 ;
      LAYER mcon ;
        RECT 5.750 5.910 5.920 6.080 ;
        RECT 5.750 5.570 5.920 5.740 ;
        RECT 7.680 5.740 7.850 5.910 ;
        RECT 8.760 5.450 8.930 5.620 ;
        RECT 5.750 5.230 5.920 5.400 ;
        RECT 7.680 5.190 7.850 5.360 ;
        RECT 9.490 5.480 9.660 5.650 ;
        RECT 5.750 4.380 5.920 4.550 ;
        RECT 7.680 4.320 7.850 4.490 ;
        RECT 5.750 4.040 5.920 4.210 ;
        RECT 8.760 4.060 8.930 4.230 ;
        RECT 9.490 4.030 9.660 4.200 ;
        RECT 5.750 3.700 5.920 3.870 ;
        RECT 7.680 3.770 7.850 3.940 ;
        RECT 0.430 3.190 0.700 3.460 ;
        RECT 9.130 3.250 9.310 3.420 ;
        RECT 5.740 2.820 5.910 2.990 ;
        RECT 7.680 2.730 7.850 2.900 ;
        RECT 5.740 2.480 5.910 2.650 ;
        RECT 8.760 2.440 8.930 2.610 ;
        RECT 5.740 2.140 5.910 2.310 ;
        RECT 7.680 2.180 7.850 2.350 ;
        RECT 9.490 2.470 9.660 2.640 ;
        RECT 5.740 1.280 5.910 1.450 ;
        RECT 7.680 1.320 7.850 1.490 ;
        RECT 5.740 0.940 5.910 1.110 ;
        RECT 8.760 1.060 8.930 1.230 ;
        RECT 9.490 1.030 9.660 1.200 ;
        RECT 5.740 0.600 5.910 0.770 ;
        RECT 7.680 0.770 7.850 0.940 ;
      LAYER met1 ;
        RECT 0.360 0.310 0.760 6.300 ;
        RECT 5.710 5.660 5.970 6.140 ;
        RECT 7.610 5.670 7.930 5.990 ;
        RECT 8.750 5.680 8.910 6.410 ;
        RECT 8.750 5.660 8.950 5.680 ;
        RECT 5.700 5.140 5.970 5.660 ;
        RECT 5.700 4.690 5.960 5.140 ;
        RECT 7.610 5.120 7.930 5.440 ;
        RECT 8.730 5.420 8.960 5.660 ;
        RECT 8.750 5.370 8.960 5.420 ;
        RECT 9.120 5.370 9.310 6.360 ;
        RECT 9.560 5.710 9.720 6.410 ;
        RECT 5.710 4.130 5.970 4.610 ;
        RECT 7.610 4.240 7.930 4.560 ;
        RECT 8.750 4.310 8.910 5.370 ;
        RECT 9.140 5.250 9.310 5.370 ;
        RECT 9.150 4.430 9.310 5.250 ;
        RECT 9.450 5.160 9.720 5.710 ;
        RECT 9.450 5.110 9.730 5.160 ;
        RECT 9.560 5.020 9.730 5.110 ;
        RECT 9.560 4.660 9.720 5.020 ;
        RECT 9.560 4.570 9.730 4.660 ;
        RECT 9.140 4.310 9.310 4.430 ;
        RECT 8.750 4.260 8.960 4.310 ;
        RECT 5.700 3.610 5.970 4.130 ;
        RECT 8.730 4.020 8.960 4.260 ;
        RECT 7.610 3.690 7.930 4.010 ;
        RECT 8.750 4.000 8.950 4.020 ;
        RECT 5.700 3.160 5.960 3.610 ;
        RECT 5.700 2.570 5.960 3.050 ;
        RECT 7.610 2.660 7.930 2.980 ;
        RECT 8.750 2.670 8.910 4.000 ;
        RECT 9.120 3.450 9.310 4.310 ;
        RECT 9.450 4.520 9.730 4.570 ;
        RECT 9.450 3.970 9.720 4.520 ;
        RECT 9.100 3.220 9.340 3.450 ;
        RECT 8.750 2.650 8.950 2.670 ;
        RECT 5.690 2.050 5.960 2.570 ;
        RECT 7.610 2.110 7.930 2.430 ;
        RECT 8.730 2.410 8.960 2.650 ;
        RECT 8.750 2.360 8.960 2.410 ;
        RECT 9.120 2.360 9.310 3.220 ;
        RECT 9.560 2.700 9.720 3.970 ;
        RECT 5.690 1.600 5.950 2.050 ;
        RECT 5.700 1.030 5.960 1.510 ;
        RECT 7.610 1.240 7.930 1.560 ;
        RECT 8.750 1.310 8.910 2.360 ;
        RECT 9.140 2.240 9.310 2.360 ;
        RECT 9.150 1.430 9.310 2.240 ;
        RECT 9.450 2.150 9.720 2.700 ;
        RECT 9.450 2.100 9.730 2.150 ;
        RECT 9.560 2.010 9.730 2.100 ;
        RECT 9.560 1.660 9.720 2.010 ;
        RECT 9.560 1.570 9.730 1.660 ;
        RECT 9.140 1.310 9.310 1.430 ;
        RECT 8.750 1.260 8.960 1.310 ;
        RECT 5.690 0.510 5.960 1.030 ;
        RECT 8.730 1.020 8.960 1.260 ;
        RECT 7.610 0.690 7.930 1.010 ;
        RECT 8.750 1.000 8.950 1.020 ;
        RECT 5.690 0.060 5.950 0.510 ;
        RECT 8.750 0.270 8.910 1.000 ;
        RECT 9.120 0.320 9.310 1.310 ;
        RECT 9.450 1.520 9.730 1.570 ;
        RECT 9.450 0.970 9.720 1.520 ;
        RECT 9.560 0.270 9.720 0.970 ;
      LAYER via ;
        RECT 7.640 5.700 7.900 5.960 ;
        RECT 7.640 5.150 7.900 5.410 ;
        RECT 7.640 4.270 7.900 4.530 ;
        RECT 7.640 3.720 7.900 3.980 ;
        RECT 7.640 2.690 7.900 2.950 ;
        RECT 7.640 2.140 7.900 2.400 ;
        RECT 7.640 1.270 7.900 1.530 ;
        RECT 7.640 0.720 7.900 0.980 ;
      LAYER met2 ;
        RECT 7.610 5.860 7.920 6.000 ;
        RECT 0.000 5.680 10.080 5.860 ;
        RECT 7.610 5.670 7.920 5.680 ;
        RECT 7.610 5.430 7.920 5.450 ;
        RECT 0.000 5.250 10.080 5.430 ;
        RECT 7.610 5.120 7.920 5.250 ;
        RECT 7.610 4.430 7.920 4.560 ;
        RECT 0.000 4.250 10.080 4.430 ;
        RECT 7.610 4.230 7.920 4.250 ;
        RECT 7.610 4.000 7.920 4.010 ;
        RECT 0.000 3.930 7.600 4.000 ;
        RECT 7.610 3.930 10.080 4.000 ;
        RECT 0.000 3.820 10.080 3.930 ;
        RECT 7.610 3.680 7.920 3.820 ;
        RECT 7.610 2.850 7.920 2.990 ;
        RECT 7.610 2.840 10.080 2.850 ;
        RECT 0.020 2.670 10.080 2.840 ;
        RECT 7.610 2.660 7.920 2.670 ;
        RECT 7.610 2.420 7.920 2.440 ;
        RECT 0.020 2.250 10.080 2.420 ;
        RECT 7.520 2.240 10.080 2.250 ;
        RECT 7.610 2.110 7.920 2.240 ;
        RECT 7.610 1.440 7.920 1.560 ;
        RECT 0.020 1.430 7.920 1.440 ;
        RECT 0.020 1.270 10.080 1.430 ;
        RECT 0.800 1.180 2.340 1.270 ;
        RECT 7.520 1.250 10.080 1.270 ;
        RECT 7.610 1.230 7.920 1.250 ;
        RECT 7.610 1.000 7.920 1.010 ;
        RECT 0.020 0.830 10.080 1.000 ;
        RECT 7.610 0.820 10.080 0.830 ;
        RECT 7.610 0.680 7.920 0.820 ;
  END
END sky130_hilas_swc4x1cellOverlap

MACRO sky130_hilas_capacitorSize02
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize02 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.970 BY 5.830 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 7.230 2.620 7.890 3.280 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 0.110 3.200 0.770 3.260 ;
        RECT 1.160 3.200 2.170 3.210 ;
        RECT 0.110 2.700 3.800 3.200 ;
        RECT 0.110 2.690 1.520 2.700 ;
        RECT 0.110 2.600 0.770 2.690 ;
        RECT 3.160 1.580 3.790 2.700 ;
        RECT 3.160 1.570 5.310 1.580 ;
        RECT 1.840 1.270 5.310 1.570 ;
        RECT 1.840 1.100 4.850 1.270 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 0.000 5.280 7.970 5.460 ;
        RECT 0.000 4.850 7.970 5.030 ;
        RECT 0.030 3.850 7.970 4.030 ;
        RECT 0.030 3.420 7.970 3.600 ;
        RECT 0.240 3.080 0.610 3.140 ;
        RECT 0.020 2.800 0.610 3.080 ;
        RECT 0.240 2.740 0.610 2.800 ;
        RECT 7.360 3.100 7.730 3.160 ;
        RECT 7.360 2.820 7.970 3.100 ;
        RECT 7.360 2.760 7.730 2.820 ;
        RECT 0.030 2.270 7.970 2.440 ;
        RECT 0.030 1.850 7.970 2.020 ;
        RECT 0.030 0.870 7.970 1.040 ;
        RECT 0.030 0.430 7.970 0.600 ;
      LAYER via2 ;
        RECT 0.290 2.800 0.570 3.080 ;
        RECT 7.410 2.820 7.690 3.100 ;
      LAYER met3 ;
        RECT 1.460 5.800 3.770 5.830 ;
        RECT 1.460 3.310 5.690 5.800 ;
        RECT 0.020 2.540 0.810 3.290 ;
        RECT 1.460 2.560 7.930 3.310 ;
        RECT 1.460 0.020 5.690 2.560 ;
        RECT 3.740 0.000 5.690 0.020 ;
      LAYER via3 ;
        RECT 0.210 2.690 0.640 3.170 ;
        RECT 7.330 2.710 7.760 3.190 ;
  END
END sky130_hilas_capacitorSize02

MACRO sky130_hilas_TopProtectStructure
  CLASS CORE ;
  FOREIGN sky130_hilas_TopProtectStructure ;
  ORIGIN 0.000 0.000 ;
  SIZE 372.850 BY 389.100 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN IO07
    PORT
      LAYER met1 ;
        RECT 371.600 180.790 372.850 184.680 ;
    END
  END IO07
  PIN IO08
    PORT
      LAYER met1 ;
        RECT 371.600 209.400 372.850 213.290 ;
    END
  END IO08
  PIN IO09
    PORT
      LAYER met1 ;
        RECT 371.580 237.980 372.830 241.870 ;
    END
  END IO09
  PIN IO10
    PORT
      LAYER met1 ;
        RECT 371.600 266.590 372.850 270.480 ;
    END
  END IO10
  PIN IO11
    PORT
      LAYER met1 ;
        RECT 371.590 295.150 372.840 299.040 ;
    END
  END IO11
  PIN IO12
    PORT
      LAYER met1 ;
        RECT 371.590 323.750 372.840 327.640 ;
    END
  END IO12
  PIN IO13
    PORT
      LAYER met1 ;
        RECT 371.600 352.350 372.850 356.240 ;
    END
  END IO13
  PIN IO25
    PORT
      LAYER met1 ;
        RECT 1.250 356.940 2.650 356.950 ;
        RECT 0.000 353.340 2.650 356.940 ;
        RECT 0.000 353.050 4.000 353.340 ;
    END
  END IO25
  PIN IO26
    PORT
      LAYER met1 ;
        RECT 0.010 324.750 2.650 328.360 ;
        RECT 0.010 324.470 4.000 324.750 ;
        RECT 1.250 324.460 4.000 324.470 ;
    END
  END IO26
  PIN IO27
    PORT
      LAYER met1 ;
        RECT 1.250 299.760 2.650 299.770 ;
        RECT 0.000 296.160 2.650 299.760 ;
        RECT 0.000 295.870 4.000 296.160 ;
    END
  END IO27
  PIN IO28
    PORT
      LAYER met1 ;
        RECT 1.260 271.170 2.650 271.180 ;
        RECT 0.020 267.570 2.650 271.170 ;
        RECT 0.020 267.280 4.000 267.570 ;
    END
  END IO28
  PIN IO29
    PORT
      LAYER met1 ;
        RECT 0.010 238.980 2.650 242.590 ;
        RECT 0.010 238.700 4.000 238.980 ;
        RECT 1.250 238.690 4.000 238.700 ;
    END
  END IO29
  PIN IO30
    PORT
      LAYER met1 ;
        RECT 1.250 213.990 2.650 214.000 ;
        RECT 0.000 210.390 2.650 213.990 ;
        RECT 0.000 210.100 4.000 210.390 ;
    END
  END IO30
  PIN IO31
    PORT
      LAYER met1 ;
        RECT 1.250 185.410 2.060 185.420 ;
        RECT 0.010 181.800 2.650 185.410 ;
        RECT 0.010 181.520 4.000 181.800 ;
        RECT 2.060 181.510 4.000 181.520 ;
    END
  END IO31
  PIN IO32
    PORT
      LAYER met1 ;
        RECT 0.040 156.820 2.080 156.830 ;
        RECT 0.040 153.210 2.650 156.820 ;
        RECT 0.040 152.940 4.000 153.210 ;
        RECT 1.270 152.930 4.000 152.940 ;
        RECT 2.060 152.920 4.000 152.930 ;
    END
  END IO32
  PIN IO33
    PORT
      LAYER met1 ;
        RECT 1.260 128.220 2.650 128.230 ;
        RECT 0.020 124.620 2.650 128.220 ;
        RECT 0.020 124.330 4.000 124.620 ;
    END
  END IO33
  PIN IO34
    PORT
      LAYER met1 ;
        RECT 1.260 99.630 2.650 99.640 ;
        RECT 0.010 96.030 2.650 99.630 ;
        RECT 0.010 95.740 4.000 96.030 ;
    END
  END IO34
  PIN IO35
    PORT
      LAYER met1 ;
        RECT 1.260 71.040 2.650 71.050 ;
        RECT 0.010 67.440 2.650 71.040 ;
        RECT 0.010 67.150 4.000 67.440 ;
    END
  END IO35
  PIN IO36
    PORT
      LAYER met1 ;
        RECT 1.270 42.450 2.650 42.460 ;
        RECT 0.020 38.850 2.650 42.450 ;
        RECT 0.020 38.560 4.000 38.850 ;
    END
  END IO36
  PIN IO37
    PORT
      LAYER met1 ;
        RECT 0.020 10.260 2.650 13.870 ;
        RECT 0.020 9.980 4.000 10.260 ;
        RECT 1.250 9.970 4.000 9.980 ;
    END
  END IO37
  PIN VSSA1
    ANTENNADIFFAREA 783.710388 ;
    PORT
      LAYER met2 ;
        RECT 15.930 385.020 101.700 385.780 ;
        RECT 3.420 385.010 101.700 385.020 ;
        RECT 3.290 384.380 101.700 385.010 ;
        RECT 3.290 383.620 16.350 384.380 ;
        RECT 16.400 384.370 17.330 384.380 ;
        RECT 44.990 384.370 45.920 384.380 ;
        RECT 73.580 384.370 74.510 384.380 ;
        RECT 3.290 382.100 5.580 383.620 ;
        RECT 16.650 383.260 16.820 384.370 ;
        RECT 45.240 383.260 45.410 384.370 ;
        RECT 73.830 383.260 74.000 384.370 ;
        RECT 3.740 382.060 5.580 382.100 ;
        RECT 4.180 373.930 5.580 382.060 ;
        RECT 4.150 373.540 5.580 373.930 ;
        RECT 4.150 346.740 5.550 373.540 ;
        RECT 4.150 346.230 5.560 346.740 ;
        RECT 4.150 346.060 6.670 346.230 ;
        RECT 4.150 345.810 5.560 346.060 ;
        RECT 4.150 318.150 5.550 345.810 ;
        RECT 4.150 317.640 5.560 318.150 ;
        RECT 4.150 317.470 6.670 317.640 ;
        RECT 4.150 317.220 5.560 317.470 ;
        RECT 4.150 289.560 5.550 317.220 ;
        RECT 4.150 289.050 5.560 289.560 ;
        RECT 4.150 288.880 6.670 289.050 ;
        RECT 4.150 288.630 5.560 288.880 ;
        RECT 4.150 260.970 5.550 288.630 ;
        RECT 4.150 260.460 5.560 260.970 ;
        RECT 4.150 260.290 6.670 260.460 ;
        RECT 4.150 260.040 5.560 260.290 ;
        RECT 4.150 232.380 5.550 260.040 ;
        RECT 4.150 231.870 5.560 232.380 ;
        RECT 4.150 231.700 6.670 231.870 ;
        RECT 4.150 231.450 5.560 231.700 ;
        RECT 4.150 203.790 5.550 231.450 ;
        RECT 4.150 203.280 5.560 203.790 ;
        RECT 4.150 203.110 6.670 203.280 ;
        RECT 4.150 202.860 5.560 203.110 ;
        RECT 4.150 175.200 5.550 202.860 ;
        RECT 4.150 174.690 5.560 175.200 ;
        RECT 4.150 174.520 6.670 174.690 ;
        RECT 4.150 174.270 5.560 174.520 ;
        RECT 4.150 146.610 5.550 174.270 ;
        RECT 4.150 146.100 5.560 146.610 ;
        RECT 4.150 145.930 6.670 146.100 ;
        RECT 4.150 145.680 5.560 145.930 ;
        RECT 4.150 118.020 5.550 145.680 ;
        RECT 4.150 117.510 5.560 118.020 ;
        RECT 4.150 117.340 6.670 117.510 ;
        RECT 4.150 117.090 5.560 117.340 ;
        RECT 4.150 89.430 5.550 117.090 ;
        RECT 4.150 88.920 5.560 89.430 ;
        RECT 4.150 88.750 6.670 88.920 ;
        RECT 4.150 88.500 5.560 88.750 ;
        RECT 4.150 60.840 5.550 88.500 ;
        RECT 4.150 60.330 5.560 60.840 ;
        RECT 4.150 60.160 6.670 60.330 ;
        RECT 4.150 59.910 5.560 60.160 ;
        RECT 4.150 32.250 5.550 59.910 ;
        RECT 4.150 31.740 5.560 32.250 ;
        RECT 4.150 31.570 6.670 31.740 ;
        RECT 4.150 31.320 5.560 31.570 ;
        RECT 4.150 3.660 5.550 31.320 ;
        RECT 4.150 3.150 5.560 3.660 ;
        RECT 4.150 2.980 6.670 3.150 ;
        RECT 4.150 2.730 5.560 2.980 ;
        RECT 4.150 0.330 5.550 2.730 ;
    END
  END VSSA1
  PIN ANALOG10
    PORT
      LAYER met1 ;
        RECT 23.620 388.670 27.510 389.080 ;
        RECT 23.620 387.910 27.530 388.670 ;
        RECT 23.640 387.870 27.530 387.910 ;
        RECT 23.640 387.280 27.540 387.870 ;
        RECT 23.640 385.930 23.930 387.280 ;
    END
  END ANALOG10
  PIN ANALOG09
    PORT
      LAYER met1 ;
        RECT 52.210 388.670 56.100 389.070 ;
        RECT 52.210 387.900 56.120 388.670 ;
        RECT 52.230 387.870 56.120 387.900 ;
        RECT 52.230 387.280 56.130 387.870 ;
        RECT 52.230 385.930 52.520 387.280 ;
    END
  END ANALOG09
  PIN ANALOG08
    PORT
      LAYER met1 ;
        RECT 80.800 388.670 84.690 389.070 ;
        RECT 80.800 387.900 84.710 388.670 ;
        RECT 80.820 387.870 84.710 387.900 ;
        RECT 80.820 387.280 84.720 387.870 ;
        RECT 80.820 385.930 81.110 387.280 ;
    END
  END ANALOG08
  PIN ANALOG07
    PORT
      LAYER met1 ;
        RECT 122.700 388.690 126.590 389.100 ;
        RECT 122.700 387.930 126.610 388.690 ;
        RECT 122.720 387.890 126.610 387.930 ;
    END
  END ANALOG07
  PIN ANALOG06
    ANTENNAGATEAREA 40.421497 ;
    ANTENNADIFFAREA 920.961548 ;
    PORT
      LAYER nwell ;
        RECT 119.570 373.120 122.310 376.620 ;
        RECT 201.010 370.530 202.740 370.870 ;
        RECT 239.600 370.530 241.330 370.870 ;
        RECT 201.010 368.970 202.760 370.530 ;
        RECT 166.810 367.070 168.580 368.660 ;
        RECT 143.170 359.310 145.200 362.280 ;
        RECT 143.990 359.260 144.530 359.310 ;
        RECT 143.810 358.810 144.530 359.260 ;
        RECT 141.960 358.630 144.530 358.810 ;
        RECT 169.670 354.130 172.170 368.240 ;
        RECT 201.030 367.340 202.760 368.970 ;
        RECT 239.580 368.970 241.330 370.530 ;
        RECT 239.580 367.340 241.310 368.970 ;
        RECT 200.970 364.170 204.280 367.340 ;
        RECT 238.060 364.170 241.370 367.340 ;
        RECT 201.000 363.520 202.750 364.170 ;
        RECT 239.570 363.520 241.320 364.170 ;
        RECT 200.970 361.310 204.280 363.520 ;
        RECT 238.060 361.310 241.370 363.520 ;
        RECT 178.790 361.270 178.820 361.280 ;
        RECT 174.690 360.970 178.820 361.270 ;
        RECT 174.690 360.930 178.790 360.970 ;
        RECT 174.690 354.680 178.800 360.930 ;
        RECT 200.960 360.350 204.280 361.310 ;
        RECT 238.050 360.350 241.370 361.310 ;
        RECT 200.960 358.140 204.270 360.350 ;
        RECT 238.050 358.140 241.360 360.350 ;
        RECT 202.000 357.780 202.560 358.140 ;
        RECT 238.220 357.490 239.500 358.140 ;
        RECT 238.050 354.320 241.360 357.490 ;
        RECT 238.210 351.370 239.490 354.320 ;
        RECT 169.670 344.000 172.170 351.000 ;
        RECT 174.670 344.210 178.090 350.800 ;
        RECT 196.420 346.080 198.980 351.060 ;
        RECT 194.380 346.070 198.980 346.080 ;
        RECT 200.510 346.070 202.740 351.050 ;
        RECT 194.380 344.560 202.740 346.070 ;
        RECT 213.980 344.560 216.540 351.060 ;
        RECT 166.770 334.520 168.540 336.110 ;
        RECT 169.630 334.940 172.130 341.940 ;
        RECT 194.380 341.810 196.940 344.560 ;
        RECT 198.470 341.810 200.700 344.560 ;
        RECT 194.380 341.800 200.700 341.810 ;
        RECT 194.380 341.650 197.030 341.800 ;
        RECT 194.380 341.640 197.210 341.650 ;
        RECT 174.700 341.130 178.120 341.530 ;
        RECT 174.700 335.160 179.850 341.130 ;
        RECT 194.380 339.580 197.030 341.640 ;
        RECT 198.470 339.580 200.700 341.800 ;
        RECT 196.510 339.460 197.030 339.580 ;
        RECT 196.510 339.260 197.020 339.460 ;
        RECT 196.510 338.730 197.030 339.260 ;
        RECT 196.620 335.770 197.030 338.730 ;
        RECT 174.700 335.130 181.120 335.160 ;
        RECT 174.700 334.940 178.120 335.130 ;
        RECT 180.240 334.970 181.120 335.130 ;
        RECT 182.010 333.690 189.850 333.700 ;
        RECT 180.000 333.670 189.850 333.690 ;
        RECT 172.200 328.000 189.850 333.670 ;
        RECT 172.200 327.970 180.040 328.000 ;
        RECT 228.730 325.630 229.580 327.240 ;
        RECT 230.110 326.430 235.160 328.040 ;
        RECT 232.640 325.630 235.160 326.430 ;
        RECT 137.440 318.280 141.360 323.980 ;
        RECT 228.730 321.600 235.160 325.630 ;
        RECT 228.730 321.080 233.990 321.600 ;
        RECT 226.990 320.800 233.990 321.080 ;
        RECT 226.990 319.470 231.680 320.800 ;
        RECT 231.920 319.250 231.990 320.800 ;
        RECT 232.210 320.270 233.990 320.800 ;
        RECT 232.640 320.050 233.990 320.270 ;
        RECT 232.640 319.250 235.160 320.050 ;
        RECT 228.730 318.440 235.160 319.250 ;
        RECT 228.730 318.380 233.990 318.440 ;
        RECT 228.730 317.640 235.160 318.380 ;
        RECT 231.920 317.580 231.990 317.640 ;
        RECT 232.640 317.580 235.160 317.640 ;
        RECT 228.730 312.750 235.160 317.580 ;
        RECT 228.730 311.140 229.580 312.750 ;
        RECT 230.110 311.940 235.160 312.750 ;
        RECT 232.640 311.880 233.990 311.940 ;
        RECT 232.630 311.410 233.990 311.880 ;
      LAYER met3 ;
        RECT 202.010 364.480 202.460 365.230 ;
        RECT 202.010 358.320 202.380 364.480 ;
        RECT 203.050 364.470 203.500 365.220 ;
        RECT 203.130 361.830 203.500 364.470 ;
        RECT 203.130 361.230 203.570 361.830 ;
        RECT 202.010 357.990 202.500 358.320 ;
        RECT 202.060 357.830 202.500 357.990 ;
        RECT 203.130 356.120 203.500 361.230 ;
        RECT 203.120 355.250 203.590 356.120 ;
    END
  END ANALOG06
  PIN ANALOG05
    PORT
      LAYER met1 ;
        RECT 193.410 388.670 197.300 389.080 ;
        RECT 193.410 387.910 197.320 388.670 ;
        RECT 193.430 387.870 197.320 387.910 ;
        RECT 193.430 387.280 197.330 387.870 ;
        RECT 193.430 385.930 193.720 387.280 ;
    END
  END ANALOG05
  PIN ANALOG04
    PORT
      LAYER met1 ;
        RECT 222.010 388.670 225.900 389.080 ;
        RECT 222.010 387.910 225.920 388.670 ;
        RECT 222.030 387.870 225.920 387.910 ;
        RECT 222.020 387.280 225.920 387.870 ;
        RECT 222.020 385.930 222.310 387.280 ;
    END
  END ANALOG04
  PIN ANALOG03
    PORT
      LAYER met1 ;
        RECT 250.600 388.670 254.490 389.080 ;
        RECT 250.600 387.910 254.510 388.670 ;
        RECT 250.620 387.870 254.510 387.910 ;
        RECT 250.610 387.280 254.510 387.870 ;
        RECT 250.610 385.930 250.900 387.280 ;
    END
  END ANALOG03
  PIN ANALOG02
    PORT
      LAYER met1 ;
        RECT 279.190 388.670 283.080 389.080 ;
        RECT 279.190 387.910 283.090 388.670 ;
        RECT 279.200 387.870 283.090 387.910 ;
        RECT 279.200 387.280 283.100 387.870 ;
        RECT 279.200 385.930 279.490 387.280 ;
    END
  END ANALOG02
  PIN ANALOG01
    PORT
      LAYER met1 ;
        RECT 307.780 388.670 311.670 389.070 ;
        RECT 307.780 387.900 311.680 388.670 ;
        RECT 307.790 387.870 311.680 387.900 ;
        RECT 307.790 387.280 311.690 387.870 ;
        RECT 307.790 385.930 308.080 387.280 ;
    END
  END ANALOG01
  PIN ANALOG00
    PORT
      LAYER met1 ;
        RECT 336.370 388.670 340.260 389.070 ;
        RECT 336.370 387.900 340.280 388.670 ;
        RECT 336.390 387.870 340.280 387.900 ;
        RECT 336.380 387.280 340.280 387.870 ;
        RECT 336.380 385.930 336.670 387.280 ;
    END
  END ANALOG00
  PIN VSSA1
    ANTENNAGATEAREA 40.421497 ;
    ANTENNADIFFAREA 909.062256 ;
    PORT
      LAYER met2 ;
        RECT 129.150 385.780 184.620 386.340 ;
        RECT 129.150 385.020 357.260 385.780 ;
        RECT 368.490 385.020 369.680 385.030 ;
        RECT 129.150 384.950 369.680 385.020 ;
        RECT 157.130 384.380 369.680 384.950 ;
        RECT 157.600 384.370 158.530 384.380 ;
        RECT 186.190 384.370 187.120 384.380 ;
        RECT 214.780 384.370 215.710 384.380 ;
        RECT 243.370 384.370 244.300 384.380 ;
        RECT 271.960 384.370 272.890 384.380 ;
        RECT 300.550 384.370 301.480 384.380 ;
        RECT 329.140 384.370 330.070 384.380 ;
        RECT 157.850 383.260 158.020 384.370 ;
        RECT 186.440 383.260 186.610 384.370 ;
        RECT 215.030 383.260 215.200 384.370 ;
        RECT 243.620 383.260 243.790 384.370 ;
        RECT 272.210 383.260 272.380 384.370 ;
        RECT 300.800 383.260 300.970 384.370 ;
        RECT 329.390 383.260 329.560 384.370 ;
        RECT 356.480 383.740 369.680 384.380 ;
        RECT 367.520 382.420 369.680 383.740 ;
        RECT 125.550 380.000 126.230 381.220 ;
        RECT 126.780 380.000 127.230 380.100 ;
        RECT 125.550 379.770 127.230 380.000 ;
        RECT 125.550 378.900 126.230 379.770 ;
        RECT 126.780 379.670 127.230 379.770 ;
        RECT 169.780 377.540 170.230 377.560 ;
        RECT 169.770 377.480 170.250 377.540 ;
        RECT 147.380 377.180 170.250 377.480 ;
        RECT 169.770 377.120 170.250 377.180 ;
        RECT 169.780 377.100 170.230 377.120 ;
        RECT 165.930 376.780 166.380 376.800 ;
        RECT 165.920 376.770 166.400 376.780 ;
        RECT 189.540 376.770 190.960 376.810 ;
        RECT 125.550 375.810 126.230 376.690 ;
        RECT 126.880 376.200 127.310 376.670 ;
        RECT 165.920 376.370 191.010 376.770 ;
        RECT 165.920 376.360 166.400 376.370 ;
        RECT 165.930 376.340 166.380 376.360 ;
        RECT 189.540 376.330 190.960 376.370 ;
        RECT 126.880 376.190 128.820 376.200 ;
        RECT 126.970 375.970 128.820 376.190 ;
        RECT 119.980 375.250 120.300 375.510 ;
        RECT 120.660 375.240 120.970 375.570 ;
        RECT 121.390 375.260 121.710 375.520 ;
        RECT 125.550 375.490 128.910 375.810 ;
        RECT 125.550 375.340 126.230 375.490 ;
        RECT 122.140 375.210 136.790 375.340 ;
        RECT 119.470 375.130 136.790 375.210 ;
        RECT 171.440 375.160 171.940 375.190 ;
        RECT 177.160 375.160 177.660 375.190 ;
        RECT 119.470 374.960 122.280 375.130 ;
        RECT 119.470 374.450 122.140 374.960 ;
        RECT 119.980 374.380 120.300 374.450 ;
        RECT 120.660 374.400 120.970 374.450 ;
        RECT 121.410 374.400 121.730 374.450 ;
        RECT 125.550 374.370 126.230 375.130 ;
        RECT 128.240 375.100 128.820 375.130 ;
        RECT 128.240 375.070 128.560 375.100 ;
        RECT 136.210 374.830 136.450 375.130 ;
        RECT 136.050 374.500 136.450 374.830 ;
        RECT 137.410 374.900 137.720 374.910 ;
        RECT 137.410 374.580 137.830 374.900 ;
        RECT 136.210 374.460 136.450 374.500 ;
        RECT 137.530 374.440 137.830 374.580 ;
        RECT 138.100 374.890 138.410 374.900 ;
        RECT 138.100 374.570 138.560 374.890 ;
        RECT 171.440 374.750 201.600 375.160 ;
        RECT 171.590 374.720 201.600 374.750 ;
        RECT 138.260 374.430 138.560 374.570 ;
        RECT 127.550 374.000 129.080 374.160 ;
        RECT 125.740 373.670 129.080 374.000 ;
        RECT 167.020 374.150 167.520 374.170 ;
        RECT 172.760 374.150 173.200 374.200 ;
        RECT 187.130 374.150 187.630 374.170 ;
        RECT 167.020 373.730 193.530 374.150 ;
        RECT 167.170 373.710 193.530 373.730 ;
        RECT 172.760 373.700 173.200 373.710 ;
        RECT 192.930 373.690 193.430 373.710 ;
        RECT 125.740 373.600 128.010 373.670 ;
        RECT 85.760 373.240 89.850 373.490 ;
        RECT 125.740 373.400 126.140 373.600 ;
        RECT 119.980 373.240 120.300 373.290 ;
        RECT 125.390 373.240 126.140 373.400 ;
        RECT 85.760 371.550 127.730 373.240 ;
        RECT 367.520 373.190 368.800 382.420 ;
        RECT 237.650 372.790 238.420 372.940 ;
        RECT 128.160 372.370 238.420 372.790 ;
        RECT 368.040 372.450 368.800 373.190 ;
        RECT 237.650 372.230 238.420 372.370 ;
        RECT 134.020 371.550 134.490 371.570 ;
        RECT 85.760 370.990 134.490 371.550 ;
        RECT 85.760 370.390 89.850 370.990 ;
        RECT 122.670 370.900 123.110 370.990 ;
        RECT 125.100 370.970 134.490 370.990 ;
        RECT 125.100 370.900 125.820 370.970 ;
        RECT 134.020 370.950 134.490 370.970 ;
        RECT 135.330 370.900 135.640 371.170 ;
        RECT 145.190 370.900 145.500 371.190 ;
        RECT 122.380 370.690 145.610 370.900 ;
        RECT 125.100 369.900 125.780 370.690 ;
        RECT 157.190 370.280 157.500 370.300 ;
        RECT 147.400 370.200 147.720 370.210 ;
        RECT 157.190 370.200 157.510 370.280 ;
        RECT 181.370 370.210 181.690 370.230 ;
        RECT 181.370 370.200 181.700 370.210 ;
        RECT 188.140 370.200 188.460 370.230 ;
        RECT 202.910 370.200 203.230 370.220 ;
        RECT 217.570 370.200 218.130 370.340 ;
        RECT 147.400 369.970 218.130 370.200 ;
        RECT 147.400 369.890 147.720 369.970 ;
        RECT 157.190 369.960 157.500 369.970 ;
        RECT 181.370 369.950 181.700 369.970 ;
        RECT 188.140 369.950 188.460 369.970 ;
        RECT 202.910 369.960 203.230 369.970 ;
        RECT 217.570 369.830 218.130 369.970 ;
        RECT 153.190 369.750 153.560 369.810 ;
        RECT 216.390 369.750 216.930 369.770 ;
        RECT 153.190 369.520 216.930 369.750 ;
        RECT 153.190 369.460 153.560 369.520 ;
        RECT 184.990 369.300 185.270 369.310 ;
        RECT 156.020 369.290 156.330 369.300 ;
        RECT 184.970 369.290 185.290 369.300 ;
        RECT 187.700 369.290 188.020 369.320 ;
        RECT 202.020 369.290 202.340 369.350 ;
        RECT 215.310 369.290 215.850 369.300 ;
        RECT 156.020 369.060 215.850 369.290 ;
        RECT 216.390 369.210 216.930 369.520 ;
        RECT 156.020 369.030 156.350 369.060 ;
        RECT 184.970 369.040 185.290 369.060 ;
        RECT 187.700 369.040 188.020 369.060 ;
        RECT 184.990 369.030 185.270 369.040 ;
        RECT 156.020 369.010 156.330 369.030 ;
        RECT 57.640 368.750 61.020 368.860 ;
        RECT 149.940 368.830 150.260 368.840 ;
        RECT 214.370 368.830 214.900 368.860 ;
        RECT 57.230 368.600 127.730 368.750 ;
        RECT 144.700 368.600 145.100 368.610 ;
        RECT 57.230 368.250 145.100 368.600 ;
        RECT 149.940 368.600 214.900 368.830 ;
        RECT 215.310 368.740 215.850 369.060 ;
        RECT 149.940 368.540 150.260 368.600 ;
        RECT 57.230 366.500 127.730 368.250 ;
        RECT 144.700 368.220 145.100 368.250 ;
        RECT 181.840 368.250 182.160 368.290 ;
        RECT 197.490 368.250 198.770 368.350 ;
        RECT 214.370 368.250 214.900 368.600 ;
        RECT 181.840 368.040 198.770 368.250 ;
        RECT 181.840 368.010 182.160 368.040 ;
        RECT 203.140 366.790 203.450 366.800 ;
        RECT 200.970 366.610 203.450 366.790 ;
        RECT 57.640 366.180 61.020 366.500 ;
        RECT 124.780 366.400 126.050 366.500 ;
        RECT 203.140 366.470 203.450 366.610 ;
        RECT 136.130 366.400 136.430 366.410 ;
        RECT 145.720 366.400 146.010 366.420 ;
        RECT 124.780 366.010 146.040 366.400 ;
        RECT 124.780 365.980 126.050 366.010 ;
        RECT 145.720 365.990 146.010 366.010 ;
        RECT 201.960 364.880 202.540 365.320 ;
        RECT 201.960 364.690 202.600 364.880 ;
        RECT 202.360 364.080 202.600 364.690 ;
        RECT 202.980 364.680 203.560 365.310 ;
        RECT 141.320 363.870 141.640 363.920 ;
        RECT 141.320 363.700 142.060 363.870 ;
        RECT 143.740 363.710 144.050 364.040 ;
        RECT 141.320 363.660 141.640 363.700 ;
        RECT 141.290 362.950 141.610 363.000 ;
        RECT 141.290 362.780 142.060 362.950 ;
        RECT 141.290 362.740 141.610 362.780 ;
        RECT 141.300 362.030 141.620 362.080 ;
        RECT 141.300 361.860 142.060 362.030 ;
        RECT 141.300 361.820 141.620 361.860 ;
        RECT 145.700 361.380 146.020 361.410 ;
        RECT 143.890 361.270 146.120 361.380 ;
        RECT 143.650 361.180 146.120 361.270 ;
        RECT 140.650 361.020 140.970 361.060 ;
        RECT 140.650 360.830 142.080 361.020 ;
        RECT 143.650 360.940 143.960 361.180 ;
        RECT 145.700 361.150 146.020 361.180 ;
        RECT 140.650 360.800 140.970 360.830 ;
        RECT 145.710 360.420 146.030 360.450 ;
        RECT 143.890 360.280 146.120 360.420 ;
        RECT 143.650 360.220 146.120 360.280 ;
        RECT 140.610 360.060 140.930 360.100 ;
        RECT 140.610 359.870 142.080 360.060 ;
        RECT 143.650 359.950 143.960 360.220 ;
        RECT 145.710 360.190 146.030 360.220 ;
        RECT 140.610 359.840 140.930 359.870 ;
        RECT 214.860 359.750 215.170 359.950 ;
        RECT 214.860 359.740 215.460 359.750 ;
        RECT 214.860 359.620 217.250 359.740 ;
        RECT 215.000 359.580 217.250 359.620 ;
        RECT 215.310 359.560 217.250 359.580 ;
        RECT 145.700 359.460 146.020 359.490 ;
        RECT 143.880 359.260 146.120 359.460 ;
        RECT 145.700 359.230 146.020 359.260 ;
        RECT 140.650 359.100 140.970 359.140 ;
        RECT 140.650 358.910 142.080 359.100 ;
        RECT 140.650 358.880 140.970 358.910 ;
        RECT 184.970 358.630 185.280 358.640 ;
        RECT 184.960 358.570 185.290 358.630 ;
        RECT 184.610 358.520 185.290 358.570 ;
        RECT 181.380 358.350 185.290 358.520 ;
        RECT 181.380 358.300 185.280 358.350 ;
        RECT 237.460 353.030 238.240 353.180 ;
        RECT 240.200 353.030 241.100 353.950 ;
        RECT 237.460 352.560 241.100 353.030 ;
        RECT 237.460 352.410 238.240 352.560 ;
        RECT 240.200 351.860 241.100 352.560 ;
        RECT 196.620 350.780 216.360 350.960 ;
        RECT 196.620 350.640 197.040 350.780 ;
        RECT 198.440 350.500 198.750 350.780 ;
        RECT 196.420 350.460 198.750 350.500 ;
        RECT 214.210 350.500 214.520 350.780 ;
        RECT 216.020 350.650 216.360 350.780 ;
        RECT 214.210 350.460 216.540 350.500 ;
        RECT 196.420 350.320 198.600 350.460 ;
        RECT 214.360 350.320 216.540 350.460 ;
        RECT 214.210 350.070 214.520 350.240 ;
        RECT 214.210 349.910 216.540 350.070 ;
        RECT 214.370 349.890 216.540 349.910 ;
        RECT 214.370 348.940 216.540 348.960 ;
        RECT 214.210 348.780 216.540 348.940 ;
        RECT 214.210 348.610 214.520 348.780 ;
        RECT 214.360 348.390 216.540 348.530 ;
        RECT 214.210 348.350 216.540 348.390 ;
        RECT 214.210 348.060 214.520 348.350 ;
        RECT 217.480 348.040 218.080 348.100 ;
        RECT 240.200 348.040 241.100 349.070 ;
        RECT 217.480 347.570 241.100 348.040 ;
        RECT 214.210 347.260 214.520 347.550 ;
        RECT 217.480 347.520 218.080 347.570 ;
        RECT 214.210 347.220 216.540 347.260 ;
        RECT 214.360 347.080 216.540 347.220 ;
        RECT 214.210 346.830 214.520 347.000 ;
        RECT 240.200 346.980 241.100 347.570 ;
        RECT 214.210 346.670 216.540 346.830 ;
        RECT 214.370 346.650 216.540 346.670 ;
        RECT 214.370 345.710 216.540 345.730 ;
        RECT 214.210 345.550 216.540 345.710 ;
        RECT 214.210 345.380 214.520 345.550 ;
        RECT 214.360 345.160 216.540 345.300 ;
        RECT 214.210 345.120 216.540 345.160 ;
        RECT 214.210 344.830 214.520 345.120 ;
        RECT 140.610 344.070 140.920 344.090 ;
        RECT 141.270 344.070 141.580 344.090 ;
        RECT 140.610 343.600 147.930 344.070 ;
        RECT 140.610 343.580 140.920 343.600 ;
        RECT 141.270 343.580 141.580 343.600 ;
        RECT 147.460 342.920 147.930 343.600 ;
        RECT 240.230 342.920 241.130 343.890 ;
        RECT 139.280 342.790 139.540 342.860 ;
        RECT 141.330 342.790 141.650 342.810 ;
        RECT 143.090 342.790 143.420 342.830 ;
        RECT 139.280 342.600 143.420 342.790 ;
        RECT 139.280 342.540 139.540 342.600 ;
        RECT 141.330 342.550 141.650 342.600 ;
        RECT 143.090 342.560 143.420 342.600 ;
        RECT 147.460 342.450 241.130 342.920 ;
        RECT 138.730 342.390 139.050 342.430 ;
        RECT 140.670 342.390 140.990 342.450 ;
        RECT 143.590 342.390 143.910 342.430 ;
        RECT 138.730 342.200 143.910 342.390 ;
        RECT 196.400 342.280 196.710 342.450 ;
        RECT 216.390 342.330 216.960 342.450 ;
        RECT 138.730 342.170 139.050 342.200 ;
        RECT 140.670 342.190 140.990 342.200 ;
        RECT 143.590 342.170 143.910 342.200 ;
        RECT 194.380 342.240 196.710 342.280 ;
        RECT 194.380 342.100 196.560 342.240 ;
        RECT 240.230 341.800 241.130 342.450 ;
        RECT 144.450 340.680 144.740 340.700 ;
        RECT 144.440 340.640 144.760 340.680 ;
        RECT 142.870 340.450 144.760 340.640 ;
        RECT 144.440 340.420 144.760 340.450 ;
        RECT 144.450 340.410 144.740 340.420 ;
        RECT 143.330 340.190 145.320 340.410 ;
        RECT 144.140 339.530 144.450 339.860 ;
        RECT 138.760 338.520 139.050 338.530 ;
        RECT 138.750 338.500 139.070 338.520 ;
        RECT 138.750 338.280 139.750 338.500 ;
        RECT 138.750 338.260 139.070 338.280 ;
        RECT 143.640 338.270 143.960 338.530 ;
        RECT 138.760 338.240 139.050 338.260 ;
        RECT 144.020 338.040 144.340 338.090 ;
        RECT 142.850 338.030 144.340 338.040 ;
        RECT 146.300 338.030 146.620 338.150 ;
        RECT 142.850 337.830 146.620 338.030 ;
        RECT 143.330 337.820 146.310 337.830 ;
        RECT 144.020 337.790 144.340 337.820 ;
        RECT 215.270 337.680 215.820 337.690 ;
        RECT 215.270 337.660 215.830 337.680 ;
        RECT 240.200 337.660 241.100 338.810 ;
        RECT 143.330 337.610 146.310 337.630 ;
        RECT 143.330 337.470 146.630 337.610 ;
        RECT 142.850 337.420 146.630 337.470 ;
        RECT 142.850 337.260 146.020 337.420 ;
        RECT 146.310 337.290 146.630 337.420 ;
        RECT 134.660 336.770 135.070 336.790 ;
        RECT 136.430 336.770 138.420 336.790 ;
        RECT 134.660 336.730 138.420 336.770 ;
        RECT 134.660 336.510 139.750 336.730 ;
        RECT 134.660 336.400 136.810 336.510 ;
        RECT 142.850 336.440 143.060 337.260 ;
        RECT 145.700 337.240 146.020 337.260 ;
        RECT 145.710 337.220 146.000 337.240 ;
        RECT 215.270 337.190 241.100 337.660 ;
        RECT 215.270 337.180 215.830 337.190 ;
        RECT 215.270 337.160 215.820 337.180 ;
        RECT 143.640 336.720 143.960 336.980 ;
        RECT 240.200 336.720 241.100 337.190 ;
        RECT 134.660 336.380 135.070 336.400 ;
        RECT 136.430 336.380 136.800 336.400 ;
        RECT 144.170 335.650 144.480 335.980 ;
        RECT 138.540 335.450 141.250 335.460 ;
        RECT 138.310 335.130 141.250 335.450 ;
        RECT 138.310 334.980 138.930 335.130 ;
        RECT 139.720 334.990 140.030 335.130 ;
        RECT 140.810 334.990 141.120 335.130 ;
        RECT 138.310 333.510 138.660 334.980 ;
        RECT 220.460 334.850 221.020 334.920 ;
        RECT 233.180 334.850 233.860 334.910 ;
        RECT 240.710 334.850 241.370 335.490 ;
        RECT 139.280 334.640 142.440 334.780 ;
        RECT 139.170 334.460 142.440 334.640 ;
        RECT 171.520 334.590 171.850 334.610 ;
        RECT 139.170 334.310 139.480 334.460 ;
        RECT 140.270 334.310 140.580 334.460 ;
        RECT 141.370 334.310 141.680 334.460 ;
        RECT 142.120 333.510 142.440 334.460 ;
        RECT 171.510 334.510 171.860 334.590 ;
        RECT 177.260 334.510 177.580 334.570 ;
        RECT 171.510 334.350 177.580 334.510 ;
        RECT 220.460 334.440 241.370 334.850 ;
        RECT 220.460 334.390 221.020 334.440 ;
        RECT 233.180 334.380 233.860 334.440 ;
        RECT 171.510 334.280 171.860 334.350 ;
        RECT 177.260 334.300 177.580 334.350 ;
        RECT 240.710 334.340 241.370 334.440 ;
        RECT 167.090 333.890 167.420 334.130 ;
        RECT 172.950 334.020 173.250 334.030 ;
        RECT 172.940 333.890 173.260 334.020 ;
        RECT 183.480 333.890 183.760 334.190 ;
        RECT 187.510 333.890 187.810 334.170 ;
        RECT 167.090 333.870 187.810 333.890 ;
        RECT 167.090 333.840 187.800 333.870 ;
        RECT 167.090 333.730 187.740 333.840 ;
        RECT 170.900 333.510 171.340 333.520 ;
        RECT 125.580 333.500 171.340 333.510 ;
        RECT 125.580 333.090 171.360 333.500 ;
        RECT 45.460 332.540 127.730 332.750 ;
        RECT 138.310 332.690 138.660 333.090 ;
        RECT 139.170 332.940 139.480 333.090 ;
        RECT 140.270 332.940 140.580 333.090 ;
        RECT 141.370 332.940 141.680 333.090 ;
        RECT 138.310 332.540 141.260 332.690 ;
        RECT 142.120 332.540 142.440 333.090 ;
        RECT 164.050 333.080 164.530 333.090 ;
        RECT 170.880 333.080 171.360 333.090 ;
        RECT 170.900 333.070 171.340 333.080 ;
        RECT 173.040 332.680 173.350 332.860 ;
        RECT 174.130 332.680 174.440 332.840 ;
        RECT 175.240 332.680 175.550 332.830 ;
        RECT 176.690 332.680 177.000 332.830 ;
        RECT 177.800 332.680 178.110 332.840 ;
        RECT 178.890 332.680 179.200 332.860 ;
        RECT 182.850 332.710 183.160 332.890 ;
        RECT 183.940 332.710 184.250 332.870 ;
        RECT 185.050 332.710 185.360 332.860 ;
        RECT 186.500 332.710 186.810 332.860 ;
        RECT 187.610 332.710 187.920 332.870 ;
        RECT 188.700 332.710 189.010 332.890 ;
        RECT 45.460 332.120 167.540 332.540 ;
        RECT 172.910 332.380 175.850 332.680 ;
        RECT 175.100 332.340 175.850 332.380 ;
        RECT 175.470 332.210 175.850 332.340 ;
        RECT 45.460 330.670 127.730 332.120 ;
        RECT 138.310 331.490 138.660 332.120 ;
        RECT 138.310 331.360 138.690 331.490 ;
        RECT 138.310 331.320 139.060 331.360 ;
        RECT 138.310 331.020 141.250 331.320 ;
        RECT 138.610 330.870 138.920 331.020 ;
        RECT 139.720 330.860 140.030 331.020 ;
        RECT 140.810 330.840 141.120 331.020 ;
        RECT 45.460 190.470 47.540 330.670 ;
        RECT 125.440 330.530 126.710 330.670 ;
        RECT 142.120 330.640 142.440 332.120 ;
        RECT 148.610 331.620 149.440 332.120 ;
        RECT 175.500 331.490 175.850 332.210 ;
        RECT 173.040 331.340 173.350 331.490 ;
        RECT 174.130 331.340 174.440 331.490 ;
        RECT 175.230 331.340 175.850 331.490 ;
        RECT 172.900 331.010 175.850 331.340 ;
        RECT 134.670 330.530 135.080 330.550 ;
        RECT 125.440 330.160 135.080 330.530 ;
        RECT 139.290 330.500 142.440 330.640 ;
        RECT 139.170 330.310 142.440 330.500 ;
        RECT 139.170 330.300 142.350 330.310 ;
        RECT 139.170 330.170 139.480 330.300 ;
        RECT 140.270 330.160 140.580 330.300 ;
        RECT 141.360 330.160 141.670 330.300 ;
        RECT 125.440 329.430 126.710 330.160 ;
        RECT 134.670 330.140 135.080 330.160 ;
        RECT 142.200 330.100 142.490 330.120 ;
        RECT 144.430 330.100 144.740 330.120 ;
        RECT 142.190 329.740 144.740 330.100 ;
        RECT 142.200 329.720 142.490 329.740 ;
        RECT 144.430 329.720 144.740 329.740 ;
        RECT 171.910 328.620 172.220 328.750 ;
        RECT 175.500 328.720 175.850 331.010 ;
        RECT 171.480 328.420 172.220 328.620 ;
        RECT 173.040 328.570 173.350 328.710 ;
        RECT 174.130 328.570 174.440 328.710 ;
        RECT 175.230 328.570 175.850 328.720 ;
        RECT 171.480 328.280 172.080 328.420 ;
        RECT 171.480 327.950 172.230 328.280 ;
        RECT 172.910 328.250 175.850 328.570 ;
        RECT 176.390 332.380 179.330 332.680 ;
        RECT 182.720 332.410 185.660 332.710 ;
        RECT 176.390 332.340 177.140 332.380 ;
        RECT 184.910 332.370 185.660 332.410 ;
        RECT 176.390 332.210 176.770 332.340 ;
        RECT 185.280 332.240 185.660 332.370 ;
        RECT 176.390 331.490 176.740 332.210 ;
        RECT 185.310 331.520 185.660 332.240 ;
        RECT 176.390 331.340 177.010 331.490 ;
        RECT 177.800 331.340 178.110 331.490 ;
        RECT 178.890 331.340 179.200 331.490 ;
        RECT 182.850 331.370 183.160 331.520 ;
        RECT 183.940 331.370 184.250 331.520 ;
        RECT 185.040 331.370 185.660 331.520 ;
        RECT 176.390 331.010 179.340 331.340 ;
        RECT 182.710 331.040 185.660 331.370 ;
        RECT 176.390 328.720 176.740 331.010 ;
        RECT 176.390 328.570 177.010 328.720 ;
        RECT 177.800 328.570 178.110 328.710 ;
        RECT 178.890 328.570 179.200 328.710 ;
        RECT 180.020 328.620 180.330 328.750 ;
        RECT 181.720 328.650 182.030 328.780 ;
        RECT 185.310 328.750 185.660 331.040 ;
        RECT 176.390 328.250 179.330 328.570 ;
        RECT 180.020 328.420 180.760 328.620 ;
        RECT 180.160 328.280 180.760 328.420 ;
        RECT 172.910 328.240 175.620 328.250 ;
        RECT 176.620 328.240 179.330 328.250 ;
        RECT 180.010 327.950 180.760 328.280 ;
        RECT 171.480 327.800 172.080 327.950 ;
        RECT 180.160 327.800 180.760 327.950 ;
        RECT 181.290 328.450 182.030 328.650 ;
        RECT 182.850 328.600 183.160 328.740 ;
        RECT 183.940 328.600 184.250 328.740 ;
        RECT 185.040 328.600 185.660 328.750 ;
        RECT 181.290 328.310 181.890 328.450 ;
        RECT 181.290 327.980 182.040 328.310 ;
        RECT 182.720 328.280 185.660 328.600 ;
        RECT 186.200 332.410 189.140 332.710 ;
        RECT 186.200 332.370 186.950 332.410 ;
        RECT 186.200 332.240 186.580 332.370 ;
        RECT 214.220 332.360 214.820 332.410 ;
        RECT 240.630 332.360 242.730 333.300 ;
        RECT 186.200 331.520 186.550 332.240 ;
        RECT 214.220 331.890 242.730 332.360 ;
        RECT 214.220 331.850 214.820 331.890 ;
        RECT 186.200 331.370 186.820 331.520 ;
        RECT 187.610 331.370 187.920 331.520 ;
        RECT 188.700 331.370 189.010 331.520 ;
        RECT 186.200 331.040 189.150 331.370 ;
        RECT 240.630 331.220 242.730 331.890 ;
        RECT 240.650 331.210 241.420 331.220 ;
        RECT 186.200 328.750 186.550 331.040 ;
        RECT 193.440 329.220 193.750 329.350 ;
        RECT 194.540 329.220 194.850 329.360 ;
        RECT 195.630 329.220 195.940 329.360 ;
        RECT 193.440 329.210 196.620 329.220 ;
        RECT 193.440 329.020 196.710 329.210 ;
        RECT 193.560 328.880 196.710 329.020 ;
        RECT 186.200 328.600 186.820 328.750 ;
        RECT 187.610 328.600 187.920 328.740 ;
        RECT 188.700 328.600 189.010 328.740 ;
        RECT 189.830 328.650 190.140 328.780 ;
        RECT 186.200 328.280 189.140 328.600 ;
        RECT 189.830 328.450 190.570 328.650 ;
        RECT 192.880 328.500 193.190 328.650 ;
        RECT 193.990 328.500 194.300 328.660 ;
        RECT 195.080 328.500 195.390 328.680 ;
        RECT 189.970 328.310 190.570 328.450 ;
        RECT 182.720 328.270 185.430 328.280 ;
        RECT 186.430 328.270 189.140 328.280 ;
        RECT 189.820 327.980 190.570 328.310 ;
        RECT 181.290 327.830 181.890 327.980 ;
        RECT 189.970 327.830 190.570 327.980 ;
        RECT 192.580 328.200 195.520 328.500 ;
        RECT 192.580 328.160 193.330 328.200 ;
        RECT 192.580 328.030 192.960 328.160 ;
        RECT 175.590 327.560 186.490 327.590 ;
        RECT 175.580 327.310 186.490 327.560 ;
        RECT 192.580 327.310 192.930 328.030 ;
        RECT 175.580 327.280 175.920 327.310 ;
        RECT 176.320 327.300 176.660 327.310 ;
        RECT 185.390 327.280 185.730 327.310 ;
        RECT 192.580 327.160 193.200 327.310 ;
        RECT 193.990 327.160 194.300 327.310 ;
        RECT 195.080 327.160 195.390 327.310 ;
        RECT 192.580 326.830 195.530 327.160 ;
        RECT 171.660 326.770 172.160 326.780 ;
        RECT 192.580 326.770 192.930 326.830 ;
        RECT 196.390 326.770 196.710 328.880 ;
        RECT 217.590 326.770 218.150 326.790 ;
        RECT 171.660 326.310 218.150 326.770 ;
        RECT 171.660 326.250 172.180 326.310 ;
        RECT 171.660 326.230 172.160 326.250 ;
        RECT 192.580 325.860 192.930 326.310 ;
        RECT 193.440 326.250 196.710 326.310 ;
        RECT 217.590 326.290 218.150 326.310 ;
        RECT 193.550 326.100 196.710 326.250 ;
        RECT 196.390 325.860 196.710 326.100 ;
        RECT 179.970 325.400 217.050 325.860 ;
        RECT 180.040 325.300 180.560 325.400 ;
        RECT 192.580 324.950 192.930 325.400 ;
        RECT 193.440 325.060 193.750 325.210 ;
        RECT 194.540 325.060 194.850 325.210 ;
        RECT 195.640 325.060 195.950 325.210 ;
        RECT 196.390 325.060 196.710 325.400 ;
        RECT 216.400 325.340 216.960 325.400 ;
        RECT 193.440 324.950 196.710 325.060 ;
        RECT 181.410 324.880 215.960 324.950 ;
        RECT 137.640 324.760 137.990 324.790 ;
        RECT 144.020 324.780 144.350 324.820 ;
        RECT 144.010 324.760 144.360 324.780 ;
        RECT 137.640 324.500 147.670 324.760 ;
        RECT 137.680 324.470 147.670 324.500 ;
        RECT 181.400 324.490 215.960 324.880 ;
        RECT 232.620 324.690 232.950 325.000 ;
        RECT 232.640 324.510 232.930 324.690 ;
        RECT 144.020 324.450 144.350 324.470 ;
        RECT 141.480 324.130 142.080 324.150 ;
        RECT 141.480 324.000 143.820 324.130 ;
        RECT 141.330 323.790 143.820 324.000 ;
        RECT 141.330 323.670 143.860 323.790 ;
        RECT 141.480 323.550 143.860 323.670 ;
        RECT 141.480 323.530 143.820 323.550 ;
        RECT 141.340 323.330 142.080 323.530 ;
        RECT 142.850 323.460 143.510 323.530 ;
        RECT 142.880 323.450 143.480 323.460 ;
        RECT 141.340 323.200 141.650 323.330 ;
        RECT 138.680 322.890 141.840 323.030 ;
        RECT 138.570 322.710 141.840 322.890 ;
        RECT 138.570 322.560 138.880 322.710 ;
        RECT 139.670 322.560 139.980 322.710 ;
        RECT 140.770 322.560 141.080 322.710 ;
        RECT 141.520 321.670 141.840 322.710 ;
        RECT 147.370 322.390 147.660 324.470 ;
        RECT 181.400 324.360 182.050 324.490 ;
        RECT 192.580 324.390 193.200 324.490 ;
        RECT 193.990 324.390 194.300 324.490 ;
        RECT 195.080 324.390 195.390 324.490 ;
        RECT 196.210 324.440 196.520 324.490 ;
        RECT 215.270 324.470 215.830 324.490 ;
        RECT 192.580 324.070 195.520 324.390 ;
        RECT 196.210 324.240 196.950 324.440 ;
        RECT 232.650 324.330 232.930 324.510 ;
        RECT 196.350 324.100 196.950 324.240 ;
        RECT 192.810 324.060 195.520 324.070 ;
        RECT 189.850 324.010 190.370 324.030 ;
        RECT 196.200 324.010 196.950 324.100 ;
        RECT 232.620 324.020 232.950 324.330 ;
        RECT 214.340 324.010 214.900 324.020 ;
        RECT 189.850 323.550 214.990 324.010 ;
        RECT 232.650 323.760 232.930 324.020 ;
        RECT 189.850 323.500 190.380 323.550 ;
        RECT 189.850 323.450 190.370 323.500 ;
        RECT 163.790 322.390 164.110 322.410 ;
        RECT 219.790 322.390 220.950 322.420 ;
        RECT 138.680 321.520 141.840 321.670 ;
        RECT 138.570 321.340 141.840 321.520 ;
        RECT 138.570 321.190 138.880 321.340 ;
        RECT 139.670 321.190 139.980 321.340 ;
        RECT 140.770 321.190 141.080 321.340 ;
        RECT 58.130 317.940 127.730 319.190 ;
        RECT 141.520 318.890 141.840 321.340 ;
        RECT 147.180 321.270 220.950 322.390 ;
        RECT 163.790 321.250 164.110 321.270 ;
        RECT 175.160 321.190 177.080 321.270 ;
        RECT 184.970 321.160 186.900 321.270 ;
        RECT 219.790 321.240 220.950 321.270 ;
        RECT 145.640 318.890 145.950 318.910 ;
        RECT 138.690 318.750 145.950 318.890 ;
        RECT 138.570 318.550 145.950 318.750 ;
        RECT 138.570 318.420 138.880 318.550 ;
        RECT 139.670 318.410 139.980 318.550 ;
        RECT 140.760 318.410 141.070 318.550 ;
        RECT 145.640 318.530 145.950 318.550 ;
        RECT 195.680 317.970 196.070 317.980 ;
        RECT 195.670 317.940 196.070 317.970 ;
        RECT 58.130 317.660 196.070 317.940 ;
        RECT 58.130 317.110 127.730 317.660 ;
        RECT 195.670 317.640 196.070 317.660 ;
        RECT 195.680 317.630 196.070 317.640 ;
        RECT 45.210 186.740 47.810 190.470 ;
        RECT 45.460 186.410 47.540 186.740 ;
        RECT 58.130 104.930 60.210 317.110 ;
        RECT 57.910 100.880 60.700 104.930 ;
        RECT 58.130 100.600 60.210 100.880 ;
      LAYER via2 ;
        RECT 202.080 364.850 202.400 365.170 ;
        RECT 203.110 364.840 203.430 365.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 368.060 173.390 368.800 173.730 ;
        RECT 367.400 172.990 368.810 173.390 ;
        RECT 367.420 172.300 368.800 172.990 ;
        RECT 367.410 171.130 368.810 172.300 ;
    END
  END VSSA1
  PIN VDDA1
    ANTENNADIFFAREA 145.420792 ;
    PORT
      LAYER nwell ;
        RECT 30.800 378.910 42.850 384.850 ;
        RECT 59.390 378.910 71.440 384.850 ;
        RECT 87.980 378.910 100.030 384.850 ;
        RECT 5.080 360.210 11.020 372.260 ;
        RECT 5.080 331.620 11.020 343.670 ;
        RECT 5.080 303.030 11.020 315.080 ;
        RECT 5.080 274.440 11.020 286.490 ;
        RECT 5.080 245.850 11.020 257.900 ;
        RECT 5.080 217.260 11.020 229.310 ;
        RECT 5.080 188.670 11.020 200.720 ;
        RECT 5.080 160.080 11.020 172.130 ;
        RECT 5.080 131.490 11.020 143.540 ;
        RECT 5.080 102.900 11.020 114.950 ;
        RECT 5.080 74.310 11.020 86.360 ;
        RECT 5.080 45.720 11.020 57.770 ;
        RECT 5.080 17.130 11.020 29.180 ;
      LAYER met2 ;
        RECT 42.270 379.480 42.910 382.490 ;
        RECT 70.860 379.480 71.500 382.490 ;
        RECT 99.450 379.480 100.090 382.490 ;
        RECT 15.930 378.650 101.700 379.480 ;
        RECT 10.450 378.080 101.700 378.650 ;
        RECT 10.450 377.250 16.200 378.080 ;
        RECT 41.370 377.950 44.000 378.080 ;
        RECT 69.960 377.950 72.590 378.080 ;
        RECT 98.550 377.950 101.180 378.080 ;
        RECT 41.370 377.440 43.920 377.950 ;
        RECT 69.960 377.440 72.510 377.950 ;
        RECT 98.550 377.440 101.100 377.950 ;
        RECT 41.370 377.370 41.990 377.440 ;
        RECT 69.960 377.370 70.580 377.440 ;
        RECT 98.550 377.370 99.170 377.440 ;
        RECT 10.450 373.410 11.850 377.250 ;
        RECT 10.450 373.330 11.980 373.410 ;
        RECT 10.450 372.320 12.490 373.330 ;
        RECT 7.440 371.680 12.490 372.320 ;
        RECT 10.450 371.400 12.490 371.680 ;
        RECT 10.450 370.780 12.560 371.400 ;
        RECT 10.450 344.820 11.850 370.780 ;
        RECT 10.450 344.740 11.980 344.820 ;
        RECT 10.450 343.730 12.490 344.740 ;
        RECT 7.440 343.090 12.490 343.730 ;
        RECT 10.450 342.810 12.490 343.090 ;
        RECT 10.450 342.190 12.560 342.810 ;
        RECT 10.450 316.230 11.850 342.190 ;
        RECT 10.450 316.150 11.980 316.230 ;
        RECT 10.450 315.140 12.490 316.150 ;
        RECT 7.440 314.500 12.490 315.140 ;
        RECT 10.450 314.220 12.490 314.500 ;
        RECT 10.450 313.600 12.560 314.220 ;
        RECT 10.450 287.640 11.850 313.600 ;
        RECT 10.450 287.560 11.980 287.640 ;
        RECT 10.450 286.550 12.490 287.560 ;
        RECT 7.440 285.910 12.490 286.550 ;
        RECT 10.450 285.630 12.490 285.910 ;
        RECT 10.450 285.010 12.560 285.630 ;
        RECT 10.450 259.050 11.850 285.010 ;
        RECT 10.450 258.970 11.980 259.050 ;
        RECT 10.450 257.960 12.490 258.970 ;
        RECT 7.440 257.320 12.490 257.960 ;
        RECT 10.450 257.040 12.490 257.320 ;
        RECT 10.450 256.420 12.560 257.040 ;
        RECT 10.450 230.460 11.850 256.420 ;
        RECT 10.450 230.380 11.980 230.460 ;
        RECT 10.450 229.370 12.490 230.380 ;
        RECT 7.440 228.730 12.490 229.370 ;
        RECT 10.450 228.450 12.490 228.730 ;
        RECT 10.450 227.830 12.560 228.450 ;
        RECT 10.450 201.870 11.850 227.830 ;
        RECT 10.450 201.790 11.980 201.870 ;
        RECT 10.450 200.780 12.490 201.790 ;
        RECT 7.440 200.140 12.490 200.780 ;
        RECT 10.450 199.860 12.490 200.140 ;
        RECT 10.450 199.240 12.560 199.860 ;
        RECT 10.450 173.280 11.850 199.240 ;
        RECT 10.450 173.200 11.980 173.280 ;
        RECT 10.450 172.190 12.490 173.200 ;
        RECT 7.440 171.550 12.490 172.190 ;
        RECT 10.450 171.270 12.490 171.550 ;
        RECT 10.450 170.650 12.560 171.270 ;
        RECT 10.450 144.690 11.850 170.650 ;
        RECT 10.450 144.610 11.980 144.690 ;
        RECT 10.450 143.600 12.490 144.610 ;
        RECT 7.440 142.960 12.490 143.600 ;
        RECT 10.450 142.680 12.490 142.960 ;
        RECT 10.450 142.060 12.560 142.680 ;
        RECT 10.450 116.100 11.850 142.060 ;
        RECT 10.450 116.020 11.980 116.100 ;
        RECT 10.450 115.010 12.490 116.020 ;
        RECT 7.440 114.370 12.490 115.010 ;
        RECT 10.450 114.090 12.490 114.370 ;
        RECT 10.450 113.470 12.560 114.090 ;
        RECT 10.450 87.510 11.850 113.470 ;
        RECT 10.450 87.430 11.980 87.510 ;
        RECT 10.450 86.420 12.490 87.430 ;
        RECT 7.440 85.780 12.490 86.420 ;
        RECT 10.450 85.500 12.490 85.780 ;
        RECT 10.450 84.880 12.560 85.500 ;
        RECT 10.450 58.920 11.850 84.880 ;
        RECT 10.450 58.840 11.980 58.920 ;
        RECT 10.450 57.830 12.490 58.840 ;
        RECT 7.440 57.190 12.490 57.830 ;
        RECT 10.450 56.910 12.490 57.190 ;
        RECT 10.450 56.290 12.560 56.910 ;
        RECT 10.450 30.330 11.850 56.290 ;
        RECT 10.450 30.250 11.980 30.330 ;
        RECT 10.450 29.240 12.490 30.250 ;
        RECT 7.440 28.600 12.490 29.240 ;
        RECT 10.450 28.320 12.490 28.600 ;
        RECT 10.450 27.700 12.560 28.320 ;
        RECT 10.450 0.000 11.850 27.700 ;
    END
    PORT
      LAYER met2 ;
        RECT 361.080 172.360 362.480 173.140 ;
        RECT 361.070 172.240 362.480 172.360 ;
        RECT 361.060 172.090 362.480 172.240 ;
        RECT 361.060 171.190 362.470 172.090 ;
    END
  END VDDA1
  PIN LADATAOUT01
    PORT
      LAYER met2 ;
        RECT 146.050 6.780 148.070 301.800 ;
        RECT 146.050 5.220 148.080 6.780 ;
        RECT 146.050 5.210 148.070 5.220 ;
    END
  END LADATAOUT01
  PIN LADATAOUT00
    PORT
      LAYER met2 ;
        RECT 141.990 5.210 144.010 301.800 ;
    END
  END LADATAOUT00
  PIN LADATAOUT02
    PORT
      LAYER met2 ;
        RECT 150.020 6.770 152.040 301.800 ;
        RECT 150.010 5.210 152.040 6.770 ;
    END
  END LADATAOUT02
  PIN LADATAOUT03
    PORT
      LAYER met2 ;
        RECT 154.020 6.770 156.040 301.800 ;
        RECT 154.010 5.210 156.040 6.770 ;
    END
  END LADATAOUT03
  PIN LADATAOUT04
    PORT
      LAYER met2 ;
        RECT 158.070 5.210 160.090 301.800 ;
    END
  END LADATAOUT04
  PIN LADATAOUT05
    PORT
      LAYER met2 ;
        RECT 162.080 6.780 164.100 301.800 ;
        RECT 162.070 5.220 164.100 6.780 ;
        RECT 162.080 5.210 164.100 5.220 ;
    END
  END LADATAOUT05
  PIN LADATAOUT06
    PORT
      LAYER met2 ;
        RECT 166.080 5.210 168.100 301.800 ;
    END
  END LADATAOUT06
  PIN LADATAOUT07
    PORT
      LAYER met2 ;
        RECT 170.170 5.210 172.190 301.800 ;
    END
  END LADATAOUT07
  PIN LADATAOUT08
    PORT
      LAYER met2 ;
        RECT 174.300 6.770 176.320 301.800 ;
        RECT 174.290 5.210 176.320 6.770 ;
    END
  END LADATAOUT08
  PIN LADATAOUT09
    PORT
      LAYER met2 ;
        RECT 178.300 6.770 180.320 301.800 ;
        RECT 178.290 5.210 180.320 6.770 ;
    END
  END LADATAOUT09
  PIN LADATAOUT10
    PORT
      LAYER met2 ;
        RECT 182.260 6.770 184.280 301.800 ;
        RECT 182.250 5.210 184.280 6.770 ;
    END
  END LADATAOUT10
  PIN LADATAOUT11
    PORT
      LAYER met2 ;
        RECT 186.310 6.780 188.330 301.800 ;
        RECT 186.310 5.220 188.340 6.780 ;
        RECT 186.310 5.210 188.330 5.220 ;
    END
  END LADATAOUT11
  PIN LADATAOUT12
    PORT
      LAYER met2 ;
        RECT 190.400 5.210 192.420 301.800 ;
    END
  END LADATAOUT12
  PIN LADATAOUT13
    PORT
      LAYER met2 ;
        RECT 194.410 6.760 196.430 301.800 ;
        RECT 194.410 5.210 196.440 6.760 ;
        RECT 194.420 5.200 196.440 5.210 ;
    END
  END LADATAOUT13
  PIN LADATAOUT14
    PORT
      LAYER met2 ;
        RECT 198.450 6.770 200.470 301.800 ;
        RECT 198.450 5.210 200.480 6.770 ;
    END
  END LADATAOUT14
  PIN LADATAOUT15
    PORT
      LAYER met2 ;
        RECT 202.540 6.750 204.560 301.800 ;
        RECT 202.540 5.210 204.570 6.750 ;
        RECT 202.550 5.190 204.570 5.210 ;
    END
  END LADATAOUT15
  PIN LADATA16
    PORT
      LAYER met2 ;
        RECT 206.590 5.210 208.610 301.800 ;
    END
  END LADATA16
  PIN LADATAOUT17
    PORT
      LAYER met2 ;
        RECT 210.560 5.210 212.580 301.800 ;
    END
  END LADATAOUT17
  PIN LADATAOUT18
    PORT
      LAYER met2 ;
        RECT 214.680 5.210 216.700 301.800 ;
    END
  END LADATAOUT18
  PIN LADATAOUT19
    PORT
      LAYER met2 ;
        RECT 218.810 5.200 220.830 301.800 ;
    END
  END LADATAOUT19
  PIN LADATAOUT20
    PORT
      LAYER met2 ;
        RECT 222.820 5.210 224.840 301.800 ;
    END
  END LADATAOUT20
  PIN LADATAOUT21
    PORT
      LAYER met2 ;
        RECT 226.830 6.890 228.850 301.800 ;
        RECT 226.830 5.230 228.870 6.890 ;
    END
  END LADATAOUT21
  PIN LADATAOUT22
    PORT
      LAYER met2 ;
        RECT 230.920 6.870 232.940 301.800 ;
        RECT 230.920 5.210 232.950 6.870 ;
    END
  END LADATAOUT22
  PIN LADATAOUT23
    PORT
      LAYER met2 ;
        RECT 235.090 5.210 237.110 301.800 ;
    END
  END LADATAOUT23
  PIN LADATAOUT24
    PORT
      LAYER met2 ;
        RECT 239.090 6.870 241.110 301.800 ;
        RECT 239.090 5.210 241.120 6.870 ;
    END
  END LADATAOUT24
  PIN LADATAIN00
    PORT
      LAYER met2 ;
        RECT 243.100 6.870 245.120 301.800 ;
        RECT 243.070 5.210 245.120 6.870 ;
    END
  END LADATAIN00
  PIN LADATAIN01
    PORT
      LAYER met2 ;
        RECT 247.060 6.870 249.080 301.800 ;
        RECT 247.050 5.210 249.080 6.870 ;
    END
  END LADATAIN01
  PIN LADATAIN02
    PORT
      LAYER met2 ;
        RECT 251.110 6.870 253.130 301.800 ;
        RECT 251.110 5.210 253.150 6.870 ;
    END
  END LADATAIN02
  PIN LADATAIN03
    PORT
      LAYER met2 ;
        RECT 255.170 6.870 257.190 301.800 ;
        RECT 255.170 5.210 257.210 6.870 ;
    END
  END LADATAIN03
  PIN VCCA
    ANTENNAGATEAREA 1.530100 ;
    ANTENNADIFFAREA 3.709700 ;
    PORT
      LAYER met2 ;
        RECT 243.440 356.810 266.770 357.240 ;
        RECT 199.490 346.340 199.810 346.400 ;
        RECT 203.420 346.340 203.740 346.350 ;
        RECT 209.220 346.340 209.540 346.350 ;
        RECT 213.150 346.340 213.470 346.400 ;
        RECT 199.490 346.160 213.470 346.340 ;
        RECT 199.490 346.110 199.810 346.160 ;
        RECT 203.420 346.090 203.740 346.160 ;
        RECT 209.220 346.090 209.540 346.160 ;
        RECT 213.150 346.110 213.470 346.160 ;
        RECT 199.870 341.500 200.190 341.620 ;
        RECT 199.870 341.360 207.700 341.500 ;
        RECT 197.570 341.280 197.890 341.340 ;
        RECT 200.050 341.310 207.700 341.360 ;
        RECT 200.050 341.290 207.880 341.310 ;
        RECT 201.590 341.280 201.920 341.290 ;
        RECT 197.570 341.110 201.920 341.280 ;
        RECT 197.570 341.060 197.890 341.110 ;
        RECT 201.590 341.050 201.920 341.110 ;
        RECT 207.490 341.100 207.880 341.290 ;
        RECT 196.510 340.750 196.660 340.880 ;
        RECT 194.380 340.730 196.660 340.750 ;
        RECT 194.380 340.570 196.710 340.730 ;
        RECT 196.400 340.460 196.710 340.570 ;
        RECT 196.400 340.400 199.780 340.460 ;
        RECT 196.510 340.370 199.780 340.400 ;
        RECT 199.850 340.370 200.170 340.570 ;
        RECT 196.510 340.320 200.170 340.370 ;
        RECT 194.380 340.310 200.170 340.320 ;
        RECT 194.380 340.180 196.560 340.310 ;
        RECT 199.640 340.210 199.940 340.310 ;
        RECT 194.380 340.140 196.710 340.180 ;
        RECT 196.400 340.070 196.710 340.140 ;
        RECT 196.400 339.990 196.900 340.070 ;
        RECT 198.510 339.990 198.830 340.040 ;
        RECT 193.730 339.830 198.830 339.990 ;
        RECT 196.490 339.810 196.900 339.830 ;
        RECT 196.490 339.710 196.810 339.810 ;
        RECT 198.510 339.780 198.830 339.830 ;
        RECT 199.720 339.230 199.950 339.240 ;
        RECT 199.720 339.200 207.290 339.230 ;
        RECT 197.990 339.060 198.310 339.110 ;
        RECT 193.730 338.930 198.310 339.060 ;
        RECT 199.720 339.030 207.350 339.200 ;
        RECT 199.720 338.930 199.960 339.030 ;
        RECT 193.730 338.900 199.960 338.930 ;
        RECT 196.510 338.750 199.960 338.900 ;
        RECT 207.160 338.830 207.880 339.030 ;
        RECT 207.760 338.820 207.880 338.830 ;
        RECT 196.510 338.730 199.880 338.750 ;
        RECT 199.850 338.550 200.170 338.690 ;
        RECT 199.850 338.530 207.310 338.550 ;
        RECT 207.760 338.530 207.880 338.540 ;
        RECT 199.850 338.430 207.880 338.530 ;
        RECT 199.860 338.330 207.880 338.430 ;
        RECT 199.860 338.320 200.180 338.330 ;
        RECT 196.450 337.370 196.650 337.870 ;
        RECT 199.720 337.370 200.040 337.510 ;
        RECT 196.450 337.250 200.040 337.370 ;
        RECT 196.450 337.220 200.000 337.250 ;
        RECT 193.730 337.170 200.000 337.220 ;
        RECT 193.730 337.060 197.840 337.170 ;
        RECT 196.560 336.930 196.870 337.060 ;
        RECT 197.520 337.010 197.840 337.060 ;
        RECT 196.440 336.780 196.870 336.930 ;
        RECT 196.440 336.660 196.720 336.780 ;
        RECT 197.020 336.320 197.340 336.340 ;
        RECT 196.450 336.290 197.340 336.320 ;
        RECT 193.730 336.130 197.340 336.290 ;
        RECT 207.310 336.270 207.860 336.280 ;
        RECT 196.610 335.990 196.920 336.130 ;
        RECT 197.020 336.080 197.340 336.130 ;
        RECT 199.730 336.260 207.860 336.270 ;
        RECT 196.490 335.860 196.920 335.990 ;
        RECT 199.730 336.050 207.880 336.260 ;
        RECT 199.730 336.040 207.320 336.050 ;
        RECT 199.730 336.030 200.500 336.040 ;
        RECT 199.730 335.860 199.970 336.030 ;
        RECT 196.490 335.780 199.970 335.860 ;
        RECT 196.600 335.620 199.970 335.780 ;
        RECT 243.260 330.870 333.310 330.890 ;
        RECT 198.490 330.370 333.310 330.870 ;
        RECT 243.260 329.970 333.310 330.370 ;
        RECT 197.950 329.470 333.310 329.970 ;
        RECT 243.260 329.070 333.310 329.470 ;
        RECT 197.480 328.800 333.310 329.070 ;
        RECT 197.480 328.570 246.860 328.800 ;
        RECT 197.000 328.160 242.790 328.170 ;
        RECT 197.000 327.670 243.000 328.160 ;
        RECT 240.990 310.370 243.000 327.670 ;
        RECT 244.850 327.580 246.860 328.570 ;
        RECT 248.930 327.580 250.940 328.800 ;
        RECT 253.020 327.580 255.030 328.800 ;
        RECT 264.230 327.580 268.760 327.660 ;
        RECT 243.540 326.430 268.830 327.580 ;
        RECT 244.850 325.380 246.860 326.430 ;
        RECT 248.930 325.380 250.940 326.430 ;
        RECT 253.020 325.380 255.030 326.430 ;
        RECT 264.230 326.410 268.760 326.430 ;
        RECT 243.580 323.290 329.070 325.380 ;
        RECT 240.930 309.850 243.000 310.370 ;
        RECT 244.850 310.370 246.860 323.290 ;
        RECT 240.930 309.720 242.960 309.850 ;
        RECT 244.850 309.720 246.920 310.370 ;
        RECT 248.930 310.350 250.940 323.290 ;
        RECT 253.020 310.370 255.030 323.290 ;
        RECT 244.850 309.680 246.860 309.720 ;
        RECT 248.930 309.700 250.970 310.350 ;
        RECT 252.990 309.790 255.030 310.370 ;
        RECT 252.990 309.720 255.020 309.790 ;
        RECT 248.930 309.620 250.940 309.700 ;
        RECT 326.980 191.860 329.070 323.290 ;
        RECT 331.220 218.330 333.310 328.800 ;
        RECT 331.050 214.620 333.480 218.330 ;
        RECT 326.990 189.960 329.070 191.860 ;
        RECT 326.990 189.840 329.080 189.960 ;
        RECT 326.880 189.780 329.080 189.840 ;
        RECT 326.620 186.100 329.150 189.780 ;
        RECT 326.880 186.080 328.970 186.100 ;
        RECT 263.390 164.230 267.990 165.010 ;
        RECT 263.390 162.550 362.540 164.230 ;
        RECT 263.390 161.260 362.670 162.550 ;
        RECT 263.390 160.440 267.990 161.260 ;
    END
  END VCCA
  OBS
      LAYER nwell ;
        RECT 119.620 380.190 129.310 384.790 ;
        RECT 119.020 378.800 129.310 380.190 ;
        RECT 137.150 378.710 139.370 380.400 ;
        RECT 172.000 378.910 184.050 384.850 ;
        RECT 200.590 378.910 212.640 384.850 ;
        RECT 229.180 378.910 241.230 384.850 ;
        RECT 257.770 378.910 269.820 384.850 ;
        RECT 286.360 378.910 298.410 384.850 ;
        RECT 314.950 378.910 327.000 384.850 ;
        RECT 343.540 378.910 355.590 384.850 ;
        RECT 131.240 375.510 135.240 377.150 ;
        RECT 142.010 376.610 144.720 376.650 ;
        RECT 136.450 375.000 138.060 375.790 ;
        RECT 138.560 375.000 139.070 375.170 ;
        RECT 139.110 375.000 140.260 375.170 ;
        RECT 131.240 371.160 135.240 374.350 ;
        RECT 136.450 373.820 140.450 375.000 ;
        RECT 142.000 374.960 144.720 376.610 ;
        RECT 136.450 373.810 137.240 373.820 ;
        RECT 138.560 373.810 140.450 373.820 ;
        RECT 137.240 373.620 137.510 373.800 ;
        RECT 138.560 373.610 139.070 373.810 ;
        RECT 139.110 373.620 140.260 373.810 ;
        RECT 142.010 373.620 144.720 373.660 ;
        RECT 142.000 370.960 144.720 373.620 ;
        RECT 164.030 368.170 165.800 368.240 ;
        RECT 164.030 366.420 165.800 366.580 ;
        RECT 166.810 365.320 168.580 366.910 ;
        RECT 233.300 366.860 236.610 366.870 ;
        RECT 235.650 366.830 235.840 366.860 ;
        RECT 164.030 364.670 165.800 364.830 ;
        RECT 166.810 363.570 168.580 365.160 ;
        RECT 210.770 364.480 213.490 366.130 ;
        RECT 210.770 364.440 213.480 364.480 ;
        RECT 164.030 362.920 165.800 363.080 ;
        RECT 166.810 361.820 168.580 363.410 ;
        RECT 210.770 363.110 213.480 363.150 ;
        RECT 210.770 363.000 213.490 363.110 ;
        RECT 209.680 362.990 213.490 363.000 ;
        RECT 209.880 362.680 210.200 362.980 ;
        RECT 210.770 361.460 213.490 362.990 ;
        RECT 216.110 362.220 216.670 364.640 ;
        RECT 225.670 362.220 226.230 364.640 ;
        RECT 228.850 364.480 231.570 366.130 ;
        RECT 228.850 364.440 231.560 364.480 ;
        RECT 228.850 363.110 231.560 363.150 ;
        RECT 228.850 361.460 231.570 363.110 ;
        RECT 233.150 363.000 235.910 363.680 ;
        RECT 232.650 362.990 235.910 363.000 ;
        RECT 232.150 362.680 232.470 362.980 ;
        RECT 233.150 362.070 235.910 362.990 ;
        RECT 236.500 362.820 237.780 363.000 ;
        RECT 164.030 361.040 165.800 361.330 ;
        RECT 216.490 360.830 216.910 360.900 ;
        RECT 233.150 360.840 235.910 361.560 ;
        RECT 233.150 360.830 236.600 360.840 ;
        RECT 164.030 359.290 165.800 359.450 ;
        RECT 166.810 358.960 168.580 360.550 ;
        RECT 188.570 358.840 188.580 360.030 ;
        RECT 164.030 357.540 165.800 357.700 ;
        RECT 166.810 357.210 168.580 358.800 ;
        RECT 188.570 358.790 188.620 358.840 ;
        RECT 188.570 358.690 188.630 358.790 ;
        RECT 188.580 357.570 188.630 358.690 ;
        RECT 210.760 358.450 213.480 360.100 ;
        RECT 210.770 358.410 213.480 358.450 ;
        RECT 164.030 355.790 165.800 355.950 ;
        RECT 166.810 355.460 168.580 357.050 ;
        RECT 164.030 354.130 165.800 354.200 ;
        RECT 166.810 353.710 168.580 355.300 ;
        RECT 190.250 353.380 191.980 355.050 ;
        RECT 200.960 354.320 204.270 357.490 ;
        RECT 210.770 357.080 213.480 357.120 ;
        RECT 210.760 356.970 213.480 357.080 ;
        RECT 209.680 356.960 213.480 356.970 ;
        RECT 209.680 356.290 209.750 356.470 ;
        RECT 210.760 355.430 213.480 356.960 ;
        RECT 216.100 356.190 216.660 358.610 ;
        RECT 225.660 356.190 226.220 358.610 ;
        RECT 228.840 358.450 231.560 360.100 ;
        RECT 233.150 358.870 235.910 360.830 ;
        RECT 228.840 358.410 231.550 358.450 ;
        RECT 228.840 357.080 231.550 357.120 ;
        RECT 228.840 355.460 231.560 357.080 ;
        RECT 233.150 356.970 235.910 358.360 ;
        RECT 236.500 356.970 237.780 357.140 ;
        RECT 232.640 356.960 235.910 356.970 ;
        RECT 233.150 356.750 235.910 356.960 ;
        RECT 236.490 356.950 237.780 356.970 ;
        RECT 236.490 356.790 237.770 356.950 ;
        RECT 232.650 355.520 233.100 355.750 ;
        RECT 228.840 355.430 233.170 355.460 ;
        RECT 231.310 355.390 233.170 355.430 ;
        RECT 220.980 353.380 222.710 355.050 ;
        RECT 186.250 351.470 187.980 353.310 ;
        RECT 190.250 351.540 192.010 353.380 ;
        RECT 164.030 350.910 165.800 351.000 ;
        RECT 164.030 349.160 165.800 349.320 ;
        RECT 166.810 348.830 168.580 350.420 ;
        RECT 164.030 347.410 165.800 347.570 ;
        RECT 166.810 347.080 168.580 348.670 ;
        RECT 188.210 348.360 189.940 350.080 ;
        RECT 190.250 348.560 191.980 351.540 ;
        RECT 209.680 351.420 209.760 351.600 ;
        RECT 220.950 351.540 222.710 353.380 ;
        RECT 206.420 349.720 206.540 349.900 ;
        RECT 205.330 349.370 205.920 349.480 ;
        RECT 207.040 349.370 207.630 349.480 ;
        RECT 164.030 345.660 165.800 345.820 ;
        RECT 166.810 345.330 168.580 346.920 ;
        RECT 184.210 346.450 185.940 348.290 ;
        RECT 188.210 346.520 189.970 348.360 ;
        RECT 164.030 344.000 165.800 344.070 ;
        RECT 166.810 343.580 168.580 345.170 ;
        RECT 188.210 343.580 189.940 346.520 ;
        RECT 205.330 346.090 205.920 346.280 ;
        RECT 207.040 346.090 207.630 346.280 ;
        RECT 210.220 344.560 212.450 351.050 ;
        RECT 220.980 348.560 222.710 351.540 ;
        RECT 224.980 351.470 226.710 353.310 ;
        RECT 234.940 351.110 236.800 354.010 ;
        RECT 234.940 351.020 237.770 351.110 ;
        RECT 236.490 350.960 237.770 351.020 ;
        RECT 234.940 350.920 237.770 350.960 ;
        RECT 232.640 349.490 233.090 349.720 ;
        RECT 231.300 349.360 233.160 349.430 ;
        RECT 234.940 347.980 236.800 350.920 ;
        RECT 234.930 347.970 236.800 347.980 ;
        RECT 234.930 344.990 236.790 347.970 ;
        RECT 203.290 344.350 203.880 344.510 ;
        RECT 234.930 341.940 236.790 344.930 ;
        RECT 163.990 341.850 165.760 341.940 ;
        RECT 202.310 341.710 202.690 341.810 ;
        RECT 206.340 341.670 206.740 341.810 ;
        RECT 163.990 340.100 165.760 340.260 ;
        RECT 166.770 339.770 168.540 341.360 ;
        RECT 203.290 341.110 203.880 341.260 ;
        RECT 163.990 338.350 165.760 338.510 ;
        RECT 166.770 338.020 168.540 339.610 ;
        RECT 143.930 337.370 146.300 337.570 ;
        RECT 143.930 335.400 146.860 337.370 ;
        RECT 163.990 336.600 165.760 336.760 ;
        RECT 166.770 336.270 168.540 337.860 ;
        RECT 143.930 334.700 146.300 335.400 ;
        RECT 163.990 334.940 165.760 335.010 ;
      LAYER li1 ;
        RECT 23.660 385.930 23.910 387.390 ;
        RECT 23.700 385.920 23.870 385.930 ;
        RECT 30.340 385.900 30.590 387.380 ;
        RECT 52.250 385.930 52.500 387.390 ;
        RECT 52.290 385.920 52.460 385.930 ;
        RECT 58.930 385.900 59.180 387.380 ;
        RECT 80.840 385.930 81.090 387.390 ;
        RECT 80.880 385.920 81.050 385.930 ;
        RECT 87.520 385.900 87.770 387.380 ;
        RECT 150.290 386.690 150.510 387.810 ;
        RECT 150.240 386.500 150.570 386.690 ;
        RECT 157.030 386.500 157.270 387.850 ;
        RECT 164.860 386.300 165.110 387.390 ;
        RECT 171.540 386.300 171.790 387.380 ;
        RECT 129.530 386.030 184.270 386.300 ;
        RECT 129.530 385.900 153.870 386.030 ;
        RECT 162.560 385.900 184.270 386.030 ;
        RECT 193.450 385.930 193.700 387.390 ;
        RECT 193.490 385.920 193.660 385.930 ;
        RECT 200.130 385.900 200.380 387.380 ;
        RECT 222.040 385.930 222.290 387.390 ;
        RECT 222.080 385.920 222.250 385.930 ;
        RECT 228.720 385.900 228.970 387.380 ;
        RECT 250.630 385.930 250.880 387.390 ;
        RECT 250.670 385.920 250.840 385.930 ;
        RECT 257.310 385.900 257.560 387.380 ;
        RECT 279.220 385.930 279.470 387.390 ;
        RECT 279.260 385.920 279.430 385.930 ;
        RECT 285.900 385.900 286.150 387.380 ;
        RECT 307.810 385.930 308.060 387.390 ;
        RECT 307.850 385.920 308.020 385.930 ;
        RECT 314.490 385.900 314.740 387.380 ;
        RECT 336.400 385.930 336.650 387.390 ;
        RECT 336.440 385.920 336.610 385.930 ;
        RECT 343.080 385.900 343.330 387.380 ;
        RECT 16.480 385.180 43.860 385.690 ;
        RECT 16.480 383.250 17.280 385.180 ;
        RECT 17.860 384.730 18.030 384.810 ;
        RECT 29.100 384.730 29.330 384.820 ;
        RECT 17.860 384.720 29.330 384.730 ;
        RECT 16.480 378.670 16.990 383.250 ;
        RECT 17.850 379.250 29.330 384.720 ;
        RECT 17.780 379.080 29.330 379.250 ;
        RECT 17.850 379.020 18.040 379.080 ;
        RECT 29.100 378.840 29.330 379.080 ;
        RECT 17.730 378.670 19.530 378.680 ;
        RECT 29.890 378.670 30.400 385.180 ;
        RECT 31.160 384.290 42.410 384.460 ;
        RECT 31.160 379.420 31.330 384.290 ;
        RECT 31.720 383.960 41.830 383.980 ;
        RECT 31.720 383.920 41.850 383.960 ;
        RECT 31.670 383.750 41.850 383.920 ;
        RECT 31.720 379.730 41.850 383.750 ;
        RECT 42.240 382.530 42.410 384.290 ;
        RECT 31.720 379.650 41.830 379.730 ;
        RECT 31.150 379.350 31.330 379.420 ;
        RECT 42.240 379.350 42.850 382.530 ;
        RECT 31.150 379.180 42.850 379.350 ;
        RECT 42.310 379.070 42.850 379.180 ;
        RECT 43.310 378.830 43.860 385.180 ;
        RECT 43.300 378.670 43.860 378.830 ;
        RECT 16.480 378.330 43.860 378.670 ;
        RECT 45.070 385.180 72.450 385.690 ;
        RECT 45.070 383.250 45.870 385.180 ;
        RECT 46.450 384.730 46.620 384.810 ;
        RECT 57.690 384.730 57.920 384.820 ;
        RECT 46.450 384.720 57.920 384.730 ;
        RECT 45.070 378.670 45.580 383.250 ;
        RECT 46.440 379.250 57.920 384.720 ;
        RECT 46.370 379.080 57.920 379.250 ;
        RECT 46.440 379.020 46.630 379.080 ;
        RECT 57.690 378.840 57.920 379.080 ;
        RECT 46.320 378.670 48.120 378.680 ;
        RECT 58.480 378.670 58.990 385.180 ;
        RECT 59.750 384.290 71.000 384.460 ;
        RECT 59.750 379.420 59.920 384.290 ;
        RECT 60.310 383.960 70.420 383.980 ;
        RECT 60.310 383.920 70.440 383.960 ;
        RECT 60.260 383.750 70.440 383.920 ;
        RECT 60.310 379.730 70.440 383.750 ;
        RECT 70.830 382.530 71.000 384.290 ;
        RECT 60.310 379.650 70.420 379.730 ;
        RECT 59.740 379.350 59.920 379.420 ;
        RECT 70.830 379.350 71.440 382.530 ;
        RECT 59.740 379.180 71.440 379.350 ;
        RECT 70.900 379.070 71.440 379.180 ;
        RECT 71.900 378.830 72.450 385.180 ;
        RECT 71.890 378.670 72.450 378.830 ;
        RECT 45.070 378.330 72.450 378.670 ;
        RECT 73.660 385.180 101.040 385.690 ;
        RECT 73.660 383.250 74.460 385.180 ;
        RECT 75.040 384.730 75.210 384.810 ;
        RECT 86.280 384.730 86.510 384.820 ;
        RECT 75.040 384.720 86.510 384.730 ;
        RECT 73.660 378.670 74.170 383.250 ;
        RECT 75.030 379.250 86.510 384.720 ;
        RECT 74.960 379.080 86.510 379.250 ;
        RECT 75.030 379.020 75.220 379.080 ;
        RECT 86.280 378.840 86.510 379.080 ;
        RECT 74.910 378.670 76.710 378.680 ;
        RECT 87.070 378.670 87.580 385.180 ;
        RECT 88.340 384.290 99.590 384.460 ;
        RECT 88.340 379.420 88.510 384.290 ;
        RECT 88.900 383.960 99.010 383.980 ;
        RECT 88.900 383.920 99.030 383.960 ;
        RECT 88.850 383.750 99.030 383.920 ;
        RECT 88.900 379.730 99.030 383.750 ;
        RECT 99.420 382.530 99.590 384.290 ;
        RECT 88.900 379.650 99.010 379.730 ;
        RECT 88.330 379.350 88.510 379.420 ;
        RECT 99.420 379.350 100.030 382.530 ;
        RECT 88.330 379.180 100.030 379.350 ;
        RECT 99.490 379.070 100.030 379.180 ;
        RECT 100.490 378.830 101.040 385.180 ;
        RECT 119.480 379.100 119.650 379.770 ;
        RECT 100.480 378.670 101.040 378.830 ;
        RECT 73.660 378.330 101.040 378.670 ;
        RECT 16.510 378.160 43.860 378.330 ;
        RECT 45.100 378.160 72.450 378.330 ;
        RECT 73.690 378.160 101.040 378.330 ;
        RECT 129.530 378.300 129.700 385.900 ;
        RECT 184.100 385.690 184.270 385.900 ;
        RECT 157.680 385.180 185.060 385.690 ;
        RECT 157.680 383.250 158.480 385.180 ;
        RECT 159.060 384.730 159.230 384.810 ;
        RECT 170.300 384.730 170.530 384.820 ;
        RECT 159.060 384.720 170.530 384.730 ;
        RECT 138.840 379.230 139.070 379.920 ;
        RECT 157.680 378.670 158.190 383.250 ;
        RECT 159.050 379.250 170.530 384.720 ;
        RECT 158.980 379.080 170.530 379.250 ;
        RECT 159.050 379.020 159.240 379.080 ;
        RECT 170.300 378.840 170.530 379.080 ;
        RECT 158.930 378.670 160.730 378.680 ;
        RECT 171.090 378.670 171.600 385.180 ;
        RECT 172.360 384.290 183.610 384.460 ;
        RECT 172.360 379.420 172.530 384.290 ;
        RECT 172.920 383.960 183.030 383.980 ;
        RECT 172.920 383.920 183.050 383.960 ;
        RECT 172.870 383.750 183.050 383.920 ;
        RECT 172.920 379.730 183.050 383.750 ;
        RECT 183.440 382.530 183.610 384.290 ;
        RECT 172.920 379.650 183.030 379.730 ;
        RECT 172.350 379.350 172.530 379.420 ;
        RECT 183.440 379.350 184.050 382.530 ;
        RECT 172.350 379.180 184.050 379.350 ;
        RECT 183.510 379.070 184.050 379.180 ;
        RECT 184.100 378.820 184.270 385.180 ;
        RECT 184.510 378.830 185.060 385.180 ;
        RECT 184.500 378.670 185.060 378.830 ;
        RECT 157.680 378.330 185.060 378.670 ;
        RECT 186.270 385.180 213.650 385.690 ;
        RECT 186.270 383.250 187.070 385.180 ;
        RECT 187.650 384.730 187.820 384.810 ;
        RECT 198.890 384.730 199.120 384.820 ;
        RECT 187.650 384.720 199.120 384.730 ;
        RECT 186.270 378.670 186.780 383.250 ;
        RECT 187.640 379.250 199.120 384.720 ;
        RECT 187.570 379.080 199.120 379.250 ;
        RECT 187.640 379.020 187.830 379.080 ;
        RECT 198.890 378.840 199.120 379.080 ;
        RECT 187.520 378.670 189.320 378.680 ;
        RECT 199.680 378.670 200.190 385.180 ;
        RECT 200.950 384.290 212.200 384.460 ;
        RECT 200.950 379.420 201.120 384.290 ;
        RECT 201.510 383.960 211.620 383.980 ;
        RECT 201.510 383.920 211.640 383.960 ;
        RECT 201.460 383.750 211.640 383.920 ;
        RECT 201.510 379.730 211.640 383.750 ;
        RECT 212.030 382.530 212.200 384.290 ;
        RECT 201.510 379.650 211.620 379.730 ;
        RECT 200.940 379.350 201.120 379.420 ;
        RECT 212.030 379.350 212.640 382.530 ;
        RECT 200.940 379.180 212.640 379.350 ;
        RECT 212.100 379.070 212.640 379.180 ;
        RECT 213.100 378.830 213.650 385.180 ;
        RECT 213.090 378.670 213.650 378.830 ;
        RECT 186.270 378.330 213.650 378.670 ;
        RECT 214.860 385.180 242.240 385.690 ;
        RECT 214.860 383.250 215.660 385.180 ;
        RECT 216.240 384.730 216.410 384.810 ;
        RECT 227.480 384.730 227.710 384.820 ;
        RECT 216.240 384.720 227.710 384.730 ;
        RECT 214.860 378.670 215.370 383.250 ;
        RECT 216.230 379.250 227.710 384.720 ;
        RECT 216.160 379.080 227.710 379.250 ;
        RECT 216.230 379.020 216.420 379.080 ;
        RECT 227.480 378.840 227.710 379.080 ;
        RECT 216.110 378.670 217.910 378.680 ;
        RECT 228.270 378.670 228.780 385.180 ;
        RECT 229.540 384.290 240.790 384.460 ;
        RECT 229.540 379.420 229.710 384.290 ;
        RECT 230.100 383.960 240.210 383.980 ;
        RECT 230.100 383.920 240.230 383.960 ;
        RECT 230.050 383.750 240.230 383.920 ;
        RECT 230.100 379.730 240.230 383.750 ;
        RECT 240.620 382.530 240.790 384.290 ;
        RECT 230.100 379.650 240.210 379.730 ;
        RECT 229.530 379.350 229.710 379.420 ;
        RECT 240.620 379.350 241.230 382.530 ;
        RECT 229.530 379.180 241.230 379.350 ;
        RECT 240.690 379.070 241.230 379.180 ;
        RECT 241.690 378.830 242.240 385.180 ;
        RECT 241.680 378.670 242.240 378.830 ;
        RECT 214.860 378.330 242.240 378.670 ;
        RECT 243.450 385.180 270.830 385.690 ;
        RECT 243.450 383.250 244.250 385.180 ;
        RECT 244.830 384.730 245.000 384.810 ;
        RECT 256.070 384.730 256.300 384.820 ;
        RECT 244.830 384.720 256.300 384.730 ;
        RECT 243.450 378.670 243.960 383.250 ;
        RECT 244.820 379.250 256.300 384.720 ;
        RECT 244.750 379.080 256.300 379.250 ;
        RECT 244.820 379.020 245.010 379.080 ;
        RECT 256.070 378.840 256.300 379.080 ;
        RECT 244.700 378.670 246.500 378.680 ;
        RECT 256.860 378.670 257.370 385.180 ;
        RECT 258.130 384.290 269.380 384.460 ;
        RECT 258.130 379.420 258.300 384.290 ;
        RECT 258.690 383.960 268.800 383.980 ;
        RECT 258.690 383.920 268.820 383.960 ;
        RECT 258.640 383.750 268.820 383.920 ;
        RECT 258.690 379.730 268.820 383.750 ;
        RECT 269.210 382.530 269.380 384.290 ;
        RECT 258.690 379.650 268.800 379.730 ;
        RECT 258.120 379.350 258.300 379.420 ;
        RECT 269.210 379.350 269.820 382.530 ;
        RECT 258.120 379.180 269.820 379.350 ;
        RECT 269.280 379.070 269.820 379.180 ;
        RECT 270.280 378.830 270.830 385.180 ;
        RECT 270.270 378.670 270.830 378.830 ;
        RECT 243.450 378.330 270.830 378.670 ;
        RECT 272.040 385.180 299.420 385.690 ;
        RECT 272.040 383.250 272.840 385.180 ;
        RECT 273.420 384.730 273.590 384.810 ;
        RECT 284.660 384.730 284.890 384.820 ;
        RECT 273.420 384.720 284.890 384.730 ;
        RECT 272.040 378.670 272.550 383.250 ;
        RECT 273.410 379.250 284.890 384.720 ;
        RECT 273.340 379.080 284.890 379.250 ;
        RECT 273.410 379.020 273.600 379.080 ;
        RECT 284.660 378.840 284.890 379.080 ;
        RECT 273.290 378.670 275.090 378.680 ;
        RECT 285.450 378.670 285.960 385.180 ;
        RECT 286.720 384.290 297.970 384.460 ;
        RECT 286.720 379.420 286.890 384.290 ;
        RECT 287.280 383.960 297.390 383.980 ;
        RECT 287.280 383.920 297.410 383.960 ;
        RECT 287.230 383.750 297.410 383.920 ;
        RECT 287.280 379.730 297.410 383.750 ;
        RECT 297.800 382.530 297.970 384.290 ;
        RECT 287.280 379.650 297.390 379.730 ;
        RECT 286.710 379.350 286.890 379.420 ;
        RECT 297.800 379.350 298.410 382.530 ;
        RECT 286.710 379.180 298.410 379.350 ;
        RECT 297.870 379.070 298.410 379.180 ;
        RECT 298.870 378.830 299.420 385.180 ;
        RECT 298.860 378.670 299.420 378.830 ;
        RECT 272.040 378.330 299.420 378.670 ;
        RECT 300.630 385.180 328.010 385.690 ;
        RECT 300.630 383.250 301.430 385.180 ;
        RECT 302.010 384.730 302.180 384.810 ;
        RECT 313.250 384.730 313.480 384.820 ;
        RECT 302.010 384.720 313.480 384.730 ;
        RECT 300.630 378.670 301.140 383.250 ;
        RECT 302.000 379.250 313.480 384.720 ;
        RECT 301.930 379.080 313.480 379.250 ;
        RECT 302.000 379.020 302.190 379.080 ;
        RECT 313.250 378.840 313.480 379.080 ;
        RECT 301.880 378.670 303.680 378.680 ;
        RECT 314.040 378.670 314.550 385.180 ;
        RECT 315.310 384.290 326.560 384.460 ;
        RECT 315.310 379.420 315.480 384.290 ;
        RECT 315.870 383.960 325.980 383.980 ;
        RECT 315.870 383.920 326.000 383.960 ;
        RECT 315.820 383.750 326.000 383.920 ;
        RECT 315.870 379.730 326.000 383.750 ;
        RECT 326.390 382.530 326.560 384.290 ;
        RECT 315.870 379.650 325.980 379.730 ;
        RECT 315.300 379.350 315.480 379.420 ;
        RECT 326.390 379.350 327.000 382.530 ;
        RECT 315.300 379.180 327.000 379.350 ;
        RECT 326.460 379.070 327.000 379.180 ;
        RECT 327.460 378.830 328.010 385.180 ;
        RECT 327.450 378.670 328.010 378.830 ;
        RECT 300.630 378.330 328.010 378.670 ;
        RECT 329.220 385.180 356.600 385.690 ;
        RECT 329.220 383.250 330.020 385.180 ;
        RECT 330.600 384.730 330.770 384.810 ;
        RECT 341.840 384.730 342.070 384.820 ;
        RECT 330.600 384.720 342.070 384.730 ;
        RECT 329.220 378.670 329.730 383.250 ;
        RECT 330.590 379.250 342.070 384.720 ;
        RECT 330.520 379.080 342.070 379.250 ;
        RECT 330.590 379.020 330.780 379.080 ;
        RECT 341.840 378.840 342.070 379.080 ;
        RECT 330.470 378.670 332.270 378.680 ;
        RECT 342.630 378.670 343.140 385.180 ;
        RECT 343.900 384.290 355.150 384.460 ;
        RECT 343.900 379.420 344.070 384.290 ;
        RECT 344.460 383.960 354.570 383.980 ;
        RECT 344.460 383.920 354.590 383.960 ;
        RECT 344.410 383.750 354.590 383.920 ;
        RECT 344.460 379.730 354.590 383.750 ;
        RECT 354.980 382.530 355.150 384.290 ;
        RECT 344.460 379.650 354.570 379.730 ;
        RECT 343.890 379.350 344.070 379.420 ;
        RECT 354.980 379.350 355.590 382.530 ;
        RECT 343.890 379.180 355.590 379.350 ;
        RECT 355.050 379.070 355.590 379.180 ;
        RECT 356.050 378.830 356.600 385.180 ;
        RECT 356.040 378.670 356.600 378.830 ;
        RECT 329.220 378.330 356.600 378.670 ;
        RECT 157.710 378.160 185.060 378.330 ;
        RECT 186.300 378.160 213.650 378.330 ;
        RECT 214.890 378.160 242.240 378.330 ;
        RECT 243.480 378.160 270.830 378.330 ;
        RECT 272.070 378.160 299.420 378.330 ;
        RECT 300.660 378.160 328.010 378.330 ;
        RECT 329.250 378.160 356.600 378.330 ;
        RECT 16.510 378.140 17.200 378.160 ;
        RECT 17.710 378.150 19.510 378.160 ;
        RECT 45.100 378.140 45.790 378.160 ;
        RECT 46.300 378.150 48.100 378.160 ;
        RECT 73.690 378.140 74.380 378.160 ;
        RECT 74.890 378.150 76.690 378.160 ;
        RECT 157.710 378.140 158.400 378.160 ;
        RECT 158.910 378.150 160.710 378.160 ;
        RECT 186.300 378.140 186.990 378.160 ;
        RECT 187.500 378.150 189.300 378.160 ;
        RECT 214.890 378.140 215.580 378.160 ;
        RECT 216.090 378.150 217.890 378.160 ;
        RECT 243.480 378.140 244.170 378.160 ;
        RECT 244.680 378.150 246.480 378.160 ;
        RECT 272.070 378.140 272.760 378.160 ;
        RECT 273.270 378.150 275.070 378.160 ;
        RECT 300.660 378.140 301.350 378.160 ;
        RECT 301.860 378.150 303.660 378.160 ;
        RECT 329.250 378.140 329.940 378.160 ;
        RECT 330.450 378.150 332.250 378.160 ;
        RECT 155.970 377.960 158.330 378.130 ;
        RECT 119.440 376.310 119.610 376.640 ;
        RECT 119.680 376.200 119.770 376.340 ;
        RECT 120.840 376.310 121.010 376.640 ;
        RECT 119.570 376.020 120.570 376.200 ;
        RECT 121.060 376.190 121.140 376.340 ;
        RECT 122.770 376.230 123.440 376.400 ;
        RECT 120.970 376.020 121.980 376.190 ;
        RECT 131.580 375.840 134.890 376.820 ;
        RECT 120.640 375.490 120.960 375.530 ;
        RECT 120.630 375.340 120.960 375.490 ;
        RECT 119.900 375.170 121.980 375.340 ;
        RECT 122.510 375.310 123.180 375.480 ;
        RECT 136.830 375.200 137.000 375.530 ;
        RECT 137.510 375.200 137.680 375.530 ;
        RECT 144.190 375.480 144.420 376.170 ;
        RECT 120.080 374.760 121.900 374.930 ;
        RECT 120.640 374.650 120.960 374.690 ;
        RECT 120.630 374.520 120.960 374.650 ;
        RECT 119.900 374.350 121.980 374.520 ;
        RECT 122.690 374.510 122.900 374.940 ;
        RECT 136.030 374.750 136.350 374.790 ;
        RECT 136.020 374.560 136.350 374.750 ;
        RECT 136.900 374.640 137.070 374.990 ;
        RECT 137.390 374.830 137.710 374.870 ;
        RECT 137.380 374.640 137.710 374.830 ;
        RECT 138.080 374.820 138.400 374.860 ;
        RECT 136.030 374.530 136.350 374.560 ;
        RECT 122.710 374.490 122.880 374.510 ;
        RECT 136.470 374.380 137.070 374.640 ;
        RECT 137.390 374.610 137.710 374.640 ;
        RECT 138.070 374.630 138.400 374.820 ;
        RECT 138.080 374.600 138.400 374.630 ;
        RECT 145.400 374.400 145.570 374.420 ;
        RECT 122.510 373.880 123.180 374.050 ;
        RECT 119.900 373.510 120.570 373.680 ;
        RECT 121.300 373.510 121.980 373.680 ;
        RECT 122.180 373.390 122.370 373.530 ;
        RECT 122.180 373.300 123.450 373.390 ;
        RECT 4.240 372.720 11.770 373.270 ;
        RECT 122.310 373.220 123.450 373.300 ;
        RECT 131.580 373.040 134.890 374.020 ;
        RECT 122.300 372.790 122.470 372.830 ;
        RECT 122.300 372.760 122.680 372.790 ;
        RECT 2.550 359.750 4.030 360.000 ;
        RECT 4.240 359.810 4.750 372.720 ;
        RECT 11.100 372.710 11.770 372.720 ;
        RECT 7.400 371.820 10.860 372.260 ;
        RECT 5.470 371.720 10.860 371.820 ;
        RECT 5.470 371.650 10.750 371.720 ;
        RECT 5.470 360.740 5.640 371.650 ;
        RECT 5.970 371.240 10.200 371.260 ;
        RECT 5.950 361.130 10.280 371.240 ;
        RECT 6.010 361.080 6.180 361.130 ;
        RECT 10.580 360.740 10.750 371.650 ;
        RECT 5.470 360.570 10.750 360.740 ;
        RECT 10.510 360.560 10.750 360.570 ;
        RECT 11.260 359.810 11.770 372.710 ;
        RECT 119.900 372.390 120.570 372.560 ;
        RECT 120.870 372.430 121.040 372.760 ;
        RECT 122.300 372.570 122.690 372.760 ;
        RECT 122.780 372.610 123.450 372.780 ;
        RECT 121.100 372.390 121.980 372.560 ;
        RECT 122.300 372.530 122.680 372.570 ;
        RECT 122.300 372.500 122.470 372.530 ;
        RECT 120.620 371.850 120.940 371.890 ;
        RECT 122.050 371.870 122.370 371.910 ;
        RECT 120.610 371.720 120.940 371.850 ;
        RECT 122.040 371.720 122.370 371.870 ;
        RECT 119.890 371.550 123.470 371.720 ;
        RECT 131.580 371.490 134.890 372.470 ;
        RECT 135.530 371.520 135.700 374.170 ;
        RECT 136.900 373.980 137.070 374.380 ;
        RECT 142.510 374.230 145.570 374.400 ;
        RECT 145.400 373.580 145.570 374.230 ;
        RECT 145.400 373.410 146.670 373.580 ;
        RECT 144.190 372.490 144.420 373.180 ;
        RECT 119.830 371.270 120.150 371.310 ;
        RECT 120.760 371.270 121.080 371.310 ;
        RECT 121.460 371.270 121.780 371.310 ;
        RECT 122.200 371.270 122.520 371.310 ;
        RECT 119.820 371.080 120.150 371.270 ;
        RECT 120.750 371.080 121.080 371.270 ;
        RECT 121.450 371.080 121.780 371.270 ;
        RECT 122.190 371.100 122.520 371.270 ;
        RECT 122.910 371.260 123.230 371.300 ;
        RECT 122.900 371.100 123.230 371.260 ;
        RECT 135.530 371.130 135.710 371.520 ;
        RECT 144.190 371.480 144.420 372.170 ;
        RECT 145.400 371.150 145.570 373.410 ;
        RECT 147.520 372.190 147.690 373.080 ;
        RECT 122.190 371.080 123.230 371.100 ;
        RECT 135.310 371.090 135.710 371.130 ;
        RECT 145.170 371.110 145.570 371.150 ;
        RECT 119.830 371.050 120.150 371.080 ;
        RECT 120.760 371.050 121.080 371.080 ;
        RECT 121.460 371.050 121.780 371.080 ;
        RECT 122.200 371.050 123.230 371.080 ;
        RECT 119.940 371.040 123.230 371.050 ;
        RECT 119.940 370.880 123.370 371.040 ;
        RECT 135.300 370.900 135.710 371.090 ;
        RECT 145.160 371.000 145.570 371.110 ;
        RECT 145.160 370.920 145.490 371.000 ;
        RECT 122.520 370.870 123.370 370.880 ;
        RECT 135.310 370.870 135.710 370.900 ;
        RECT 145.170 370.890 145.490 370.920 ;
        RECT 135.530 370.790 135.710 370.870 ;
        RECT 144.600 369.750 146.120 369.760 ;
        RECT 144.600 368.960 146.150 369.750 ;
        RECT 201.790 369.140 202.340 369.570 ;
        RECT 240.000 369.140 240.550 369.570 ;
        RECT 168.470 368.190 168.820 368.290 ;
        RECT 172.060 368.240 172.230 368.280 ;
        RECT 171.080 368.220 172.230 368.240 ;
        RECT 170.130 368.190 170.590 368.220 ;
        RECT 167.060 368.020 167.820 368.190 ;
        RECT 168.070 368.020 169.240 368.190 ;
        RECT 169.480 368.050 170.590 368.190 ;
        RECT 171.040 368.050 172.230 368.220 ;
        RECT 169.480 368.020 170.300 368.050 ;
        RECT 167.060 368.010 167.290 368.020 ;
        RECT 167.020 367.570 167.290 368.010 ;
        RECT 170.040 367.880 170.300 368.020 ;
        RECT 168.500 367.570 168.830 367.830 ;
        RECT 169.450 367.780 169.740 367.810 ;
        RECT 169.410 367.610 169.740 367.780 ;
        RECT 169.450 367.570 169.740 367.610 ;
        RECT 170.040 367.710 171.220 367.880 ;
        RECT 170.040 367.570 170.300 367.710 ;
        RECT 166.470 367.430 166.640 367.490 ;
        RECT 166.440 367.210 166.660 367.430 ;
        RECT 166.990 367.390 167.320 367.570 ;
        RECT 167.570 367.400 169.730 367.570 ;
        RECT 169.970 367.400 170.300 367.570 ;
        RECT 170.440 367.560 171.220 367.710 ;
        RECT 170.070 367.350 170.300 367.400 ;
        RECT 166.470 367.160 166.640 367.210 ;
        RECT 170.070 367.120 170.240 367.350 ;
        RECT 170.590 367.210 170.800 367.540 ;
        RECT 171.040 367.270 171.220 367.560 ;
        RECT 171.500 367.550 171.830 367.720 ;
        RECT 169.860 367.110 170.240 367.120 ;
        RECT 169.860 367.050 170.330 367.110 ;
        RECT 171.580 367.090 171.760 367.550 ;
        RECT 171.770 367.370 172.390 367.540 ;
        RECT 201.790 367.410 202.340 367.840 ;
        RECT 240.000 367.410 240.550 367.840 ;
        RECT 169.520 367.000 170.330 367.050 ;
        RECT 169.510 366.940 170.330 367.000 ;
        RECT 169.510 366.880 170.250 366.940 ;
        RECT 170.800 366.920 171.760 367.090 ;
        RECT 169.860 366.830 170.250 366.880 ;
        RECT 168.470 366.440 168.820 366.540 ;
        RECT 172.060 366.490 172.230 366.530 ;
        RECT 171.080 366.470 172.230 366.490 ;
        RECT 170.130 366.440 170.590 366.470 ;
        RECT 167.060 366.270 167.820 366.440 ;
        RECT 168.070 366.270 169.240 366.440 ;
        RECT 169.480 366.300 170.590 366.440 ;
        RECT 171.040 366.300 172.230 366.470 ;
        RECT 169.480 366.270 170.300 366.300 ;
        RECT 167.060 366.260 167.290 366.270 ;
        RECT 167.020 365.820 167.290 366.260 ;
        RECT 170.040 366.130 170.300 366.270 ;
        RECT 168.500 365.820 168.830 366.080 ;
        RECT 169.450 366.030 169.740 366.060 ;
        RECT 169.410 365.860 169.740 366.030 ;
        RECT 169.450 365.820 169.740 365.860 ;
        RECT 170.040 365.960 171.220 366.130 ;
        RECT 170.040 365.820 170.300 365.960 ;
        RECT 166.470 365.680 166.640 365.740 ;
        RECT 166.440 365.460 166.660 365.680 ;
        RECT 166.990 365.640 167.320 365.820 ;
        RECT 167.570 365.650 169.730 365.820 ;
        RECT 169.970 365.650 170.300 365.820 ;
        RECT 170.440 365.810 171.220 365.960 ;
        RECT 170.070 365.600 170.300 365.650 ;
        RECT 166.470 365.410 166.640 365.460 ;
        RECT 170.070 365.370 170.240 365.600 ;
        RECT 170.590 365.460 170.800 365.790 ;
        RECT 171.040 365.520 171.220 365.810 ;
        RECT 171.500 365.800 171.830 365.970 ;
        RECT 192.570 365.800 193.240 366.670 ;
        RECT 201.370 366.610 201.570 366.960 ;
        RECT 202.850 366.710 203.380 366.880 ;
        RECT 238.960 366.710 239.490 366.880 ;
        RECT 201.360 366.580 201.570 366.610 ;
        RECT 201.360 366.000 201.580 366.580 ;
        RECT 201.360 365.990 201.570 366.000 ;
        RECT 201.740 365.820 201.930 365.830 ;
        RECT 169.860 365.360 170.240 365.370 ;
        RECT 169.860 365.300 170.330 365.360 ;
        RECT 171.580 365.340 171.760 365.800 ;
        RECT 171.770 365.620 172.390 365.790 ;
        RECT 201.730 365.530 201.930 365.820 ;
        RECT 169.520 365.250 170.330 365.300 ;
        RECT 169.510 365.190 170.330 365.250 ;
        RECT 169.510 365.130 170.250 365.190 ;
        RECT 170.800 365.170 171.760 365.340 ;
        RECT 201.670 365.200 201.940 365.530 ;
        RECT 169.860 365.080 170.250 365.130 ;
        RECT 143.740 364.950 144.060 364.990 ;
        RECT 144.830 364.960 145.150 365.000 ;
        RECT 143.740 364.880 144.070 364.950 ;
        RECT 143.740 364.730 144.110 364.880 ;
        RECT 143.910 364.550 144.110 364.730 ;
        RECT 144.500 364.550 144.700 364.880 ;
        RECT 144.830 364.770 145.160 364.960 ;
        RECT 144.830 364.740 145.150 364.770 ;
        RECT 168.470 364.690 168.820 364.790 ;
        RECT 172.060 364.740 172.230 364.780 ;
        RECT 171.080 364.720 172.230 364.740 ;
        RECT 202.130 364.720 202.300 366.330 ;
        RECT 170.130 364.690 170.590 364.720 ;
        RECT 167.060 364.520 167.820 364.690 ;
        RECT 168.070 364.520 169.240 364.690 ;
        RECT 169.480 364.550 170.590 364.690 ;
        RECT 171.040 364.550 172.230 364.720 ;
        RECT 169.480 364.520 170.300 364.550 ;
        RECT 202.120 364.530 202.300 364.720 ;
        RECT 202.960 364.630 203.130 366.320 ;
        RECT 203.550 366.130 203.880 366.300 ;
        RECT 204.850 365.820 206.950 366.670 ;
        RECT 240.770 366.610 240.970 366.960 ;
        RECT 240.770 366.580 240.980 366.610 ;
        RECT 208.280 366.320 208.470 366.550 ;
        RECT 208.560 366.270 209.440 366.440 ;
        RECT 208.750 365.880 208.940 365.990 ;
        RECT 208.640 365.760 208.940 365.880 ;
        RECT 209.270 365.880 209.440 366.270 ;
        RECT 208.640 365.710 208.860 365.760 ;
        RECT 209.270 365.710 209.660 365.880 ;
        RECT 203.550 365.340 203.880 365.510 ;
        RECT 204.900 365.340 205.250 365.510 ;
        RECT 211.070 365.090 211.300 365.610 ;
        RECT 207.350 364.920 207.670 364.960 ;
        RECT 208.600 364.920 209.680 365.090 ;
        RECT 210.010 364.920 211.300 365.090 ;
        RECT 229.150 364.920 229.380 365.610 ;
        RECT 234.430 365.490 234.750 365.530 ;
        RECT 234.430 365.300 234.760 365.490 ;
        RECT 234.430 365.270 234.750 365.300 ;
        RECT 207.340 364.730 207.670 364.920 ;
        RECT 233.340 364.860 233.980 365.040 ;
        RECT 234.360 364.870 234.710 365.040 ;
        RECT 234.810 365.030 235.000 365.140 ;
        RECT 234.810 364.910 235.140 365.030 ;
        RECT 234.890 364.830 235.140 364.910 ;
        RECT 203.550 364.550 203.880 364.720 ;
        RECT 204.900 364.550 205.240 364.720 ;
        RECT 207.350 364.700 207.670 364.730 ;
        RECT 167.060 364.510 167.290 364.520 ;
        RECT 143.360 364.240 143.690 364.410 ;
        RECT 142.200 364.040 142.520 364.080 ;
        RECT 167.020 364.070 167.290 364.510 ;
        RECT 170.040 364.380 170.300 364.520 ;
        RECT 168.500 364.070 168.830 364.330 ;
        RECT 169.450 364.280 169.740 364.310 ;
        RECT 169.410 364.110 169.740 364.280 ;
        RECT 169.450 364.070 169.740 364.110 ;
        RECT 170.040 364.210 171.220 364.380 ;
        RECT 208.280 364.330 208.470 364.560 ;
        RECT 233.740 364.480 233.910 364.490 ;
        RECT 233.740 364.440 234.140 364.480 ;
        RECT 170.040 364.070 170.300 364.210 ;
        RECT 142.200 363.850 142.530 364.040 ;
        RECT 143.750 363.960 144.070 364.000 ;
        RECT 144.840 363.970 145.160 364.010 ;
        RECT 143.750 363.890 144.080 363.960 ;
        RECT 144.090 363.890 144.260 363.940 ;
        RECT 144.580 363.890 144.770 363.930 ;
        RECT 143.750 363.860 144.260 363.890 ;
        RECT 144.510 363.860 144.770 363.890 ;
        RECT 142.200 363.820 142.520 363.850 ;
        RECT 142.220 363.750 142.430 363.820 ;
        RECT 143.750 363.740 144.770 363.860 ;
        RECT 144.840 363.780 145.170 363.970 ;
        RECT 166.470 363.930 166.640 363.990 ;
        RECT 144.840 363.750 145.160 363.780 ;
        RECT 143.920 363.700 144.770 363.740 ;
        RECT 166.440 363.710 166.660 363.930 ;
        RECT 166.990 363.890 167.320 364.070 ;
        RECT 167.570 363.900 169.730 364.070 ;
        RECT 169.970 363.900 170.300 364.070 ;
        RECT 170.440 364.060 171.220 364.210 ;
        RECT 170.070 363.850 170.300 363.900 ;
        RECT 143.920 363.610 144.710 363.700 ;
        RECT 166.470 363.660 166.640 363.710 ;
        RECT 170.070 363.620 170.240 363.850 ;
        RECT 170.590 363.710 170.800 364.040 ;
        RECT 171.040 363.770 171.220 364.060 ;
        RECT 171.500 364.050 171.830 364.220 ;
        RECT 208.580 364.130 208.660 364.300 ;
        RECT 143.920 363.560 144.270 363.610 ;
        RECT 144.510 363.560 144.710 363.610 ;
        RECT 169.860 363.610 170.240 363.620 ;
        RECT 144.090 363.550 144.270 363.560 ;
        RECT 169.860 363.550 170.330 363.610 ;
        RECT 171.580 363.590 171.760 364.050 ;
        RECT 171.770 363.870 172.390 364.040 ;
        RECT 209.140 363.980 209.350 364.410 ;
        RECT 209.160 363.960 209.330 363.980 ;
        RECT 169.520 363.500 170.330 363.550 ;
        RECT 169.510 363.440 170.330 363.500 ;
        RECT 143.370 363.250 143.700 363.420 ;
        RECT 169.510 363.380 170.250 363.440 ;
        RECT 170.800 363.420 171.760 363.590 ;
        RECT 169.860 363.330 170.250 363.380 ;
        RECT 142.180 363.120 142.500 363.160 ;
        RECT 142.180 362.930 142.510 363.120 ;
        RECT 201.780 363.110 202.330 363.540 ;
        RECT 207.340 363.230 207.660 363.270 ;
        RECT 208.290 363.260 208.480 363.490 ;
        RECT 208.610 363.390 208.660 363.560 ;
        RECT 208.750 363.440 208.940 363.670 ;
        RECT 209.750 363.560 209.920 364.130 ;
        RECT 214.030 363.980 214.220 364.300 ;
        RECT 228.120 363.980 228.310 364.300 ;
        RECT 233.740 364.250 234.150 364.440 ;
        RECT 234.350 364.410 234.540 364.520 ;
        RECT 234.350 364.290 234.690 364.410 ;
        RECT 233.740 364.220 234.140 364.250 ;
        RECT 234.400 364.240 234.690 364.290 ;
        RECT 233.740 364.190 233.910 364.220 ;
        RECT 234.970 364.150 235.140 364.830 ;
        RECT 239.210 364.630 239.380 366.320 ;
        RECT 240.040 364.720 240.210 366.330 ;
        RECT 240.760 366.000 240.980 366.580 ;
        RECT 240.770 365.990 240.980 366.000 ;
        RECT 240.410 365.820 240.600 365.830 ;
        RECT 240.410 365.530 240.610 365.820 ;
        RECT 240.400 365.200 240.690 365.530 ;
        RECT 240.040 364.530 240.220 364.720 ;
        RECT 214.030 363.890 214.310 363.980 ;
        RECT 210.670 363.750 214.310 363.890 ;
        RECT 228.030 363.890 228.310 363.980 ;
        RECT 228.030 363.750 231.670 363.890 ;
        RECT 210.670 363.710 214.220 363.750 ;
        RECT 209.030 363.530 209.080 363.540 ;
        RECT 209.660 363.530 209.740 363.540 ;
        RECT 209.030 363.490 209.740 363.530 ;
        RECT 209.030 363.450 209.760 363.490 ;
        RECT 208.990 363.330 209.830 363.450 ;
        RECT 214.030 363.290 214.220 363.710 ;
        RECT 228.120 363.710 231.670 363.750 ;
        RECT 228.120 363.290 228.310 363.710 ;
        RECT 233.360 363.360 233.570 363.790 ;
        RECT 233.380 363.340 233.550 363.360 ;
        RECT 143.750 362.970 144.070 363.010 ;
        RECT 144.840 362.980 145.160 363.020 ;
        RECT 142.180 362.900 142.500 362.930 ;
        RECT 143.750 362.900 144.080 362.970 ;
        RECT 143.750 362.750 144.120 362.900 ;
        RECT 143.920 362.570 144.120 362.750 ;
        RECT 144.510 362.570 144.710 362.900 ;
        RECT 144.840 362.790 145.170 362.980 ;
        RECT 168.470 362.940 168.820 363.040 ;
        RECT 172.060 362.990 172.230 363.030 ;
        RECT 171.080 362.970 172.230 362.990 ;
        RECT 202.120 362.970 202.300 363.110 ;
        RECT 170.130 362.940 170.590 362.970 ;
        RECT 144.840 362.760 145.160 362.790 ;
        RECT 167.060 362.770 167.820 362.940 ;
        RECT 168.070 362.770 169.240 362.940 ;
        RECT 169.480 362.800 170.590 362.940 ;
        RECT 171.040 362.800 172.230 362.970 ;
        RECT 169.480 362.770 170.300 362.800 ;
        RECT 167.060 362.760 167.290 362.770 ;
        RECT 143.370 362.260 143.700 362.430 ;
        RECT 167.020 362.320 167.290 362.760 ;
        RECT 170.040 362.630 170.300 362.770 ;
        RECT 168.500 362.320 168.830 362.580 ;
        RECT 169.450 362.530 169.740 362.560 ;
        RECT 169.410 362.360 169.740 362.530 ;
        RECT 169.450 362.320 169.740 362.360 ;
        RECT 170.040 362.460 171.220 362.630 ;
        RECT 170.040 362.320 170.300 362.460 ;
        RECT 143.660 362.180 143.980 362.220 ;
        RECT 166.470 362.180 166.640 362.240 ;
        RECT 142.160 362.130 142.480 362.170 ;
        RECT 142.160 361.940 142.490 362.130 ;
        RECT 143.660 362.010 143.990 362.180 ;
        RECT 144.960 362.080 145.280 362.120 ;
        RECT 143.660 361.960 144.140 362.010 ;
        RECT 142.160 361.910 142.480 361.940 ;
        RECT 143.830 361.830 144.140 361.960 ;
        RECT 143.810 361.810 144.140 361.830 ;
        RECT 143.970 361.680 144.140 361.810 ;
        RECT 144.650 361.680 144.820 362.010 ;
        RECT 144.960 361.890 145.290 362.080 ;
        RECT 166.440 361.960 166.660 362.180 ;
        RECT 166.990 362.140 167.320 362.320 ;
        RECT 167.570 362.150 169.730 362.320 ;
        RECT 169.970 362.150 170.300 362.320 ;
        RECT 170.440 362.310 171.220 362.460 ;
        RECT 170.070 362.100 170.300 362.150 ;
        RECT 166.470 361.910 166.640 361.960 ;
        RECT 144.960 361.860 145.280 361.890 ;
        RECT 170.070 361.870 170.240 362.100 ;
        RECT 170.590 361.960 170.800 362.290 ;
        RECT 171.040 362.020 171.220 362.310 ;
        RECT 171.500 362.300 171.830 362.470 ;
        RECT 169.860 361.860 170.240 361.870 ;
        RECT 169.860 361.800 170.330 361.860 ;
        RECT 171.580 361.840 171.760 362.300 ;
        RECT 171.770 362.120 172.390 362.290 ;
        RECT 201.670 362.160 201.940 362.490 ;
        RECT 201.730 361.870 201.930 362.160 ;
        RECT 201.740 361.860 201.930 361.870 ;
        RECT 169.520 361.750 170.330 361.800 ;
        RECT 169.510 361.690 170.330 361.750 ;
        RECT 169.510 361.630 170.250 361.690 ;
        RECT 170.800 361.670 171.760 361.840 ;
        RECT 202.130 361.810 202.300 362.970 ;
        RECT 201.360 361.690 201.570 361.700 ;
        RECT 143.330 361.570 143.760 361.590 ;
        RECT 169.860 361.580 170.250 361.630 ;
        RECT 143.310 361.400 143.760 361.570 ;
        RECT 143.330 361.380 143.760 361.400 ;
        RECT 143.660 361.190 143.980 361.230 ;
        RECT 143.660 361.020 143.990 361.190 ;
        RECT 144.960 361.090 145.280 361.130 ;
        RECT 201.360 361.110 201.580 361.690 ;
        RECT 201.780 361.380 202.330 361.810 ;
        RECT 202.130 361.360 202.300 361.380 ;
        RECT 202.960 361.370 203.130 363.060 ;
        RECT 203.550 362.970 203.880 363.140 ;
        RECT 204.900 362.970 205.240 363.140 ;
        RECT 207.330 363.040 207.660 363.230 ;
        RECT 233.880 363.220 234.070 363.330 ;
        RECT 233.880 363.100 234.300 363.220 ;
        RECT 207.340 363.010 207.660 363.040 ;
        RECT 233.780 363.050 234.300 363.100 ;
        RECT 234.650 363.050 235.910 363.230 ;
        RECT 238.980 363.110 239.300 363.130 ;
        RECT 239.990 363.110 240.540 363.540 ;
        RECT 236.730 363.070 237.050 363.110 ;
        RECT 233.780 362.970 233.970 363.050 ;
        RECT 233.760 362.940 233.970 362.970 ;
        RECT 233.750 362.930 233.970 362.940 ;
        RECT 235.140 362.930 235.470 363.050 ;
        RECT 233.630 362.880 233.970 362.930 ;
        RECT 233.500 362.850 233.970 362.880 ;
        RECT 236.730 362.880 237.060 363.070 ;
        RECT 238.980 363.020 239.550 363.110 ;
        RECT 236.730 362.850 237.050 362.880 ;
        RECT 233.460 362.820 233.970 362.850 ;
        RECT 208.600 362.600 209.680 362.770 ;
        RECT 210.000 362.670 211.240 362.770 ;
        RECT 233.460 362.760 233.950 362.820 ;
        RECT 233.460 362.710 233.800 362.760 ;
        RECT 234.430 362.730 234.750 362.770 ;
        RECT 210.000 362.600 211.300 362.670 ;
        RECT 203.550 362.180 203.880 362.350 ;
        RECT 204.900 362.180 205.250 362.350 ;
        RECT 210.330 362.280 210.500 362.340 ;
        RECT 208.740 361.980 208.930 362.090 ;
        RECT 210.310 362.070 210.520 362.280 ;
        RECT 210.330 362.000 210.500 362.070 ;
        RECT 211.070 361.980 211.300 362.600 ;
        RECT 229.150 361.980 229.380 362.710 ;
        RECT 233.460 362.690 233.720 362.710 ;
        RECT 233.460 362.670 233.690 362.690 ;
        RECT 233.460 362.630 233.670 362.670 ;
        RECT 233.460 362.350 233.630 362.630 ;
        RECT 234.430 362.540 234.760 362.730 ;
        RECT 234.810 362.670 234.980 362.680 ;
        RECT 234.810 362.630 235.140 362.670 ;
        RECT 234.430 362.510 234.750 362.540 ;
        RECT 234.810 362.440 235.150 362.630 ;
        RECT 235.790 362.610 235.980 362.720 ;
        RECT 236.820 362.670 237.020 362.850 ;
        RECT 235.670 362.600 235.980 362.610 ;
        RECT 235.420 362.490 235.980 362.600 ;
        RECT 234.810 362.410 235.140 362.440 ;
        RECT 235.420 362.430 235.800 362.490 ;
        RECT 234.810 362.380 234.980 362.410 ;
        RECT 236.500 362.160 236.670 362.490 ;
        RECT 236.680 362.420 237.000 362.460 ;
        RECT 236.680 362.340 237.010 362.420 ;
        RECT 236.680 362.200 237.020 362.340 ;
        RECT 236.820 362.010 237.020 362.200 ;
        RECT 237.410 362.010 237.960 363.000 ;
        RECT 238.780 362.940 239.550 363.020 ;
        RECT 240.040 362.970 240.220 363.110 ;
        RECT 238.780 362.870 239.380 362.940 ;
        RECT 238.780 362.850 239.110 362.870 ;
        RECT 238.780 362.570 239.140 362.850 ;
        RECT 238.430 362.400 239.140 362.570 ;
        RECT 208.640 361.860 208.930 361.980 ;
        RECT 209.200 361.970 209.660 361.980 ;
        RECT 208.640 361.810 208.850 361.860 ;
        RECT 209.200 361.820 209.670 361.970 ;
        RECT 209.200 361.810 209.660 361.820 ;
        RECT 203.550 361.390 203.880 361.560 ;
        RECT 204.900 361.390 205.250 361.560 ;
        RECT 208.310 361.470 208.500 361.580 ;
        RECT 209.200 361.470 209.390 361.810 ;
        RECT 233.340 361.660 233.980 361.840 ;
        RECT 234.360 361.670 234.710 361.840 ;
        RECT 234.810 361.830 235.000 361.940 ;
        RECT 234.810 361.710 235.140 361.830 ;
        RECT 238.430 361.730 239.130 361.960 ;
        RECT 234.890 361.630 235.140 361.710 ;
        RECT 208.310 361.350 209.390 361.470 ;
        RECT 208.430 361.290 209.390 361.350 ;
        RECT 233.740 361.280 233.910 361.290 ;
        RECT 143.660 360.970 144.140 361.020 ;
        RECT 143.830 360.840 144.140 360.970 ;
        RECT 143.810 360.820 144.140 360.840 ;
        RECT 143.970 360.690 144.140 360.820 ;
        RECT 144.650 360.690 144.820 361.020 ;
        RECT 144.960 360.900 145.290 361.090 ;
        RECT 201.360 361.080 201.570 361.110 ;
        RECT 144.960 360.870 145.280 360.900 ;
        RECT 169.860 360.740 170.250 360.790 ;
        RECT 169.510 360.680 170.250 360.740 ;
        RECT 169.510 360.620 170.330 360.680 ;
        RECT 143.330 360.580 143.760 360.600 ;
        RECT 143.310 360.410 143.760 360.580 ;
        RECT 169.520 360.570 170.330 360.620 ;
        RECT 169.860 360.510 170.330 360.570 ;
        RECT 170.800 360.530 171.760 360.700 ;
        RECT 169.860 360.500 170.240 360.510 ;
        RECT 166.470 360.410 166.640 360.460 ;
        RECT 143.330 360.390 143.760 360.410 ;
        RECT 143.660 360.200 143.980 360.240 ;
        RECT 143.660 360.030 143.990 360.200 ;
        RECT 166.440 360.190 166.660 360.410 ;
        RECT 170.070 360.270 170.240 360.500 ;
        RECT 144.960 360.100 145.280 360.140 ;
        RECT 166.470 360.130 166.640 360.190 ;
        RECT 143.660 359.980 144.140 360.030 ;
        RECT 143.830 359.900 144.140 359.980 ;
        RECT 143.830 359.850 144.300 359.900 ;
        RECT 143.810 359.830 144.300 359.850 ;
        RECT 4.240 359.300 11.770 359.810 ;
        RECT 143.970 359.810 144.300 359.830 ;
        RECT 143.970 359.700 144.360 359.810 ;
        RECT 144.650 359.700 144.820 360.030 ;
        RECT 144.960 359.910 145.290 360.100 ;
        RECT 166.990 360.050 167.320 360.230 ;
        RECT 170.070 360.220 170.300 360.270 ;
        RECT 167.570 360.050 169.730 360.220 ;
        RECT 169.970 360.050 170.300 360.220 ;
        RECT 170.590 360.080 170.800 360.410 ;
        RECT 171.040 360.060 171.220 360.350 ;
        RECT 171.580 360.070 171.760 360.530 ;
        RECT 172.750 360.520 172.920 360.940 ;
        RECT 173.560 360.820 173.800 360.850 ;
        RECT 173.230 360.650 173.800 360.820 ;
        RECT 174.040 360.650 175.380 360.820 ;
        RECT 175.830 360.650 176.790 360.820 ;
        RECT 173.560 360.610 173.800 360.650 ;
        RECT 176.340 360.640 176.510 360.650 ;
        RECT 172.680 360.300 172.850 360.340 ;
        RECT 171.770 360.080 172.390 360.250 ;
        RECT 172.620 360.130 172.850 360.300 ;
        RECT 175.970 360.200 176.310 360.380 ;
        RECT 144.960 359.880 145.280 359.910 ;
        RECT 144.130 359.620 144.360 359.700 ;
        RECT 167.020 359.610 167.290 360.050 ;
        RECT 168.500 359.790 168.830 360.050 ;
        RECT 169.450 360.010 169.740 360.050 ;
        RECT 169.410 359.840 169.740 360.010 ;
        RECT 169.450 359.810 169.740 359.840 ;
        RECT 170.040 359.910 170.300 360.050 ;
        RECT 170.440 359.910 171.220 360.060 ;
        RECT 143.330 359.590 143.760 359.610 ;
        RECT 143.310 359.420 143.760 359.590 ;
        RECT 167.060 359.600 167.290 359.610 ;
        RECT 170.040 359.740 171.220 359.910 ;
        RECT 171.500 359.900 171.830 360.070 ;
        RECT 172.680 359.780 172.850 360.130 ;
        RECT 172.920 359.910 173.110 360.140 ;
        RECT 173.210 360.030 173.580 360.200 ;
        RECT 174.040 360.030 176.790 360.200 ;
        RECT 177.320 359.960 177.490 360.890 ;
        RECT 177.720 360.050 177.890 360.940 ;
        RECT 201.370 360.930 201.570 361.080 ;
        RECT 233.460 361.000 233.630 361.280 ;
        RECT 233.740 361.240 234.140 361.280 ;
        RECT 233.740 361.050 234.150 361.240 ;
        RECT 234.350 361.210 234.540 361.320 ;
        RECT 234.970 361.250 235.140 361.630 ;
        RECT 238.380 361.500 239.130 361.730 ;
        RECT 234.350 361.090 234.690 361.210 ;
        RECT 233.740 361.020 234.140 361.050 ;
        RECT 234.400 361.040 234.690 361.090 ;
        RECT 234.810 361.190 235.140 361.250 ;
        RECT 201.360 360.730 201.570 360.930 ;
        RECT 202.850 360.850 203.380 360.980 ;
        RECT 202.840 360.810 203.380 360.850 ;
        RECT 233.460 360.960 233.670 361.000 ;
        RECT 233.740 360.990 233.910 361.020 ;
        RECT 234.810 361.000 235.150 361.190 ;
        RECT 235.420 361.140 235.800 361.200 ;
        RECT 235.420 361.030 235.980 361.140 ;
        RECT 235.670 361.020 235.980 361.030 ;
        RECT 236.500 361.020 236.670 361.350 ;
        RECT 236.820 361.310 237.020 361.500 ;
        RECT 236.680 361.170 237.020 361.310 ;
        RECT 236.680 361.090 237.010 361.170 ;
        RECT 236.680 361.050 237.000 361.090 ;
        RECT 233.460 360.940 233.690 360.960 ;
        RECT 234.810 360.950 235.140 361.000 ;
        RECT 233.460 360.920 233.720 360.940 ;
        RECT 233.460 360.870 233.800 360.920 ;
        RECT 235.790 360.910 235.980 361.020 ;
        RECT 233.460 360.810 233.950 360.870 ;
        RECT 201.360 360.580 201.560 360.730 ;
        RECT 202.840 360.680 203.370 360.810 ;
        RECT 233.460 360.780 233.970 360.810 ;
        RECT 233.500 360.750 233.970 360.780 ;
        RECT 233.630 360.700 233.970 360.750 ;
        RECT 233.750 360.690 233.970 360.700 ;
        RECT 233.760 360.660 233.970 360.690 ;
        RECT 201.350 360.550 201.560 360.580 ;
        RECT 201.350 359.970 201.570 360.550 ;
        RECT 201.350 359.960 201.560 359.970 ;
        RECT 201.730 359.790 201.920 359.800 ;
        RECT 170.040 359.600 170.300 359.740 ;
        RECT 167.060 359.430 167.820 359.600 ;
        RECT 168.070 359.430 169.240 359.600 ;
        RECT 169.480 359.570 170.300 359.600 ;
        RECT 169.480 359.430 170.590 359.570 ;
        RECT 143.330 359.400 143.760 359.420 ;
        RECT 168.470 359.330 168.820 359.430 ;
        RECT 170.130 359.400 170.590 359.430 ;
        RECT 171.040 359.400 172.230 359.570 ;
        RECT 201.720 359.500 201.920 359.790 ;
        RECT 171.080 359.380 172.230 359.400 ;
        RECT 172.060 359.340 172.230 359.380 ;
        RECT 2.540 353.280 4.000 353.320 ;
        RECT 2.540 353.110 4.010 353.280 ;
        RECT 2.540 353.070 4.000 353.110 ;
        RECT 4.240 346.690 4.750 359.300 ;
        RECT 5.110 358.510 11.090 358.740 ;
        RECT 5.200 347.450 10.850 358.510 ;
        RECT 11.260 348.940 11.770 359.300 ;
        RECT 169.860 358.990 170.250 359.040 ;
        RECT 172.680 359.020 172.850 359.370 ;
        RECT 169.510 358.930 170.250 358.990 ;
        RECT 169.510 358.870 170.330 358.930 ;
        RECT 169.520 358.820 170.330 358.870 ;
        RECT 169.860 358.760 170.330 358.820 ;
        RECT 170.800 358.780 171.760 358.950 ;
        RECT 172.620 358.850 172.850 359.020 ;
        RECT 172.920 359.010 173.110 359.240 ;
        RECT 173.210 358.950 173.580 359.120 ;
        RECT 174.040 358.950 176.790 359.120 ;
        RECT 172.680 358.810 172.850 358.850 ;
        RECT 169.860 358.750 170.240 358.760 ;
        RECT 166.470 358.660 166.640 358.710 ;
        RECT 166.440 358.440 166.660 358.660 ;
        RECT 170.070 358.520 170.240 358.750 ;
        RECT 166.470 358.380 166.640 358.440 ;
        RECT 166.990 358.300 167.320 358.480 ;
        RECT 170.070 358.470 170.300 358.520 ;
        RECT 167.570 358.300 169.730 358.470 ;
        RECT 169.970 358.300 170.300 358.470 ;
        RECT 170.590 358.330 170.800 358.660 ;
        RECT 171.040 358.310 171.220 358.600 ;
        RECT 171.580 358.320 171.760 358.780 ;
        RECT 175.970 358.770 176.310 358.950 ;
        RECT 171.770 358.330 172.390 358.500 ;
        RECT 167.020 357.860 167.290 358.300 ;
        RECT 168.500 358.040 168.830 358.300 ;
        RECT 169.450 358.260 169.740 358.300 ;
        RECT 169.410 358.090 169.740 358.260 ;
        RECT 169.450 358.060 169.740 358.090 ;
        RECT 170.040 358.160 170.300 358.300 ;
        RECT 170.440 358.160 171.220 358.310 ;
        RECT 167.060 357.850 167.290 357.860 ;
        RECT 170.040 357.990 171.220 358.160 ;
        RECT 171.500 358.150 171.830 358.320 ;
        RECT 172.750 358.210 172.920 358.630 ;
        RECT 173.560 358.500 173.800 358.540 ;
        RECT 176.340 358.500 176.510 358.510 ;
        RECT 173.230 358.330 173.800 358.500 ;
        RECT 174.040 358.330 175.380 358.500 ;
        RECT 175.830 358.330 176.790 358.500 ;
        RECT 173.560 358.300 173.800 358.330 ;
        RECT 177.320 358.260 177.490 359.190 ;
        RECT 201.640 359.170 201.930 359.500 ;
        RECT 177.720 358.210 177.890 359.100 ;
        RECT 202.120 358.690 202.290 360.300 ;
        RECT 202.110 358.500 202.290 358.690 ;
        RECT 202.950 358.600 203.120 360.290 ;
        RECT 210.320 359.830 215.380 360.660 ;
        RECT 233.360 359.840 233.570 360.590 ;
        RECT 233.780 360.580 233.970 360.660 ;
        RECT 235.140 360.580 235.470 360.700 ;
        RECT 236.820 360.660 237.020 360.840 ;
        RECT 236.730 360.630 237.050 360.660 ;
        RECT 233.780 360.530 234.300 360.580 ;
        RECT 233.880 360.410 234.300 360.530 ;
        RECT 233.880 360.300 234.070 360.410 ;
        RECT 234.650 360.400 235.910 360.580 ;
        RECT 236.730 360.440 237.060 360.630 ;
        RECT 237.410 360.510 237.960 361.500 ;
        RECT 238.430 361.080 239.130 361.500 ;
        RECT 239.210 361.370 239.380 362.870 ;
        RECT 240.040 361.810 240.210 362.970 ;
        RECT 240.400 362.160 240.690 362.490 ;
        RECT 240.410 361.870 240.610 362.160 ;
        RECT 240.410 361.860 240.600 361.870 ;
        RECT 239.990 361.380 240.540 361.810 ;
        RECT 240.770 361.690 240.980 361.700 ;
        RECT 240.040 361.360 240.210 361.380 ;
        RECT 240.760 361.110 240.980 361.690 ;
        RECT 240.770 361.080 240.980 361.110 ;
        RECT 238.960 360.850 239.490 360.980 ;
        RECT 240.770 360.930 240.970 361.080 ;
        RECT 238.950 360.810 239.490 360.850 ;
        RECT 238.950 360.680 239.480 360.810 ;
        RECT 240.760 360.730 240.970 360.930 ;
        RECT 239.030 360.660 239.350 360.680 ;
        RECT 238.420 360.650 239.350 360.660 ;
        RECT 238.420 360.480 239.120 360.650 ;
        RECT 240.760 360.580 240.960 360.730 ;
        RECT 240.760 360.550 240.970 360.580 ;
        RECT 236.730 360.400 237.050 360.440 ;
        RECT 239.200 360.190 239.370 360.290 ;
        RECT 233.880 360.020 234.070 360.130 ;
        RECT 236.730 360.070 237.050 360.110 ;
        RECT 233.880 359.900 234.300 360.020 ;
        RECT 233.780 359.850 234.300 359.900 ;
        RECT 234.650 359.850 235.910 360.030 ;
        RECT 236.730 359.880 237.060 360.070 ;
        RECT 239.020 360.000 239.370 360.190 ;
        RECT 236.730 359.850 237.050 359.880 ;
        RECT 214.830 359.750 215.310 359.830 ;
        RECT 233.780 359.770 233.970 359.850 ;
        RECT 214.830 359.650 215.160 359.750 ;
        RECT 233.760 359.740 233.970 359.770 ;
        RECT 233.750 359.730 233.970 359.740 ;
        RECT 235.140 359.730 235.470 359.850 ;
        RECT 233.630 359.680 233.970 359.730 ;
        RECT 233.500 359.650 233.970 359.680 ;
        RECT 236.820 359.670 237.020 359.850 ;
        RECT 207.580 359.460 207.900 359.500 ;
        RECT 207.570 359.270 207.900 359.460 ;
        RECT 207.580 359.240 207.900 359.270 ;
        RECT 212.950 358.890 213.180 359.580 ;
        RECT 214.830 359.500 214.980 359.650 ;
        RECT 233.460 359.620 233.970 359.650 ;
        RECT 229.140 358.890 229.370 359.580 ;
        RECT 233.460 359.560 233.950 359.620 ;
        RECT 233.460 359.510 233.800 359.560 ;
        RECT 233.460 359.490 233.720 359.510 ;
        RECT 233.460 359.470 233.690 359.490 ;
        RECT 233.460 359.430 233.670 359.470 ;
        RECT 234.420 359.460 234.740 359.500 ;
        RECT 233.460 359.150 233.630 359.430 ;
        RECT 233.740 359.410 233.910 359.440 ;
        RECT 233.740 359.380 234.140 359.410 ;
        RECT 234.420 359.390 234.750 359.460 ;
        RECT 233.740 359.190 234.150 359.380 ;
        RECT 234.400 359.340 234.750 359.390 ;
        RECT 234.350 359.270 234.750 359.340 ;
        RECT 234.810 359.430 235.140 359.480 ;
        RECT 234.350 359.240 234.740 359.270 ;
        RECT 234.810 359.240 235.150 359.430 ;
        RECT 235.790 359.410 235.980 359.520 ;
        RECT 235.670 359.400 235.980 359.410 ;
        RECT 235.420 359.290 235.980 359.400 ;
        RECT 234.350 359.220 234.690 359.240 ;
        RECT 233.740 359.150 234.140 359.190 ;
        RECT 233.740 359.140 233.910 359.150 ;
        RECT 234.350 359.110 234.540 359.220 ;
        RECT 234.810 359.180 235.140 359.240 ;
        RECT 235.420 359.230 235.800 359.290 ;
        RECT 234.970 358.800 235.140 359.180 ;
        RECT 236.500 359.160 236.670 359.490 ;
        RECT 236.680 359.420 237.000 359.460 ;
        RECT 236.680 359.340 237.010 359.420 ;
        RECT 236.680 359.200 237.020 359.340 ;
        RECT 236.820 359.010 237.020 359.200 ;
        RECT 237.410 359.010 237.960 360.000 ;
        RECT 238.420 359.930 239.370 360.000 ;
        RECT 238.420 359.820 239.120 359.930 ;
        RECT 238.430 359.140 239.130 359.400 ;
        RECT 238.380 358.910 239.130 359.140 ;
        RECT 233.340 358.590 233.980 358.770 ;
        RECT 234.360 358.590 234.710 358.760 ;
        RECT 234.890 358.720 235.140 358.800 ;
        RECT 234.810 358.600 235.140 358.720 ;
        RECT 232.400 358.520 232.720 358.560 ;
        RECT 232.390 358.330 232.720 358.520 ;
        RECT 234.810 358.490 235.000 358.600 ;
        RECT 238.430 358.520 239.130 358.910 ;
        RECT 239.200 358.600 239.370 359.930 ;
        RECT 240.030 358.690 240.200 360.300 ;
        RECT 240.750 359.970 240.970 360.550 ;
        RECT 240.760 359.960 240.970 359.970 ;
        RECT 240.400 359.790 240.590 359.800 ;
        RECT 240.400 359.500 240.600 359.790 ;
        RECT 240.390 359.170 240.680 359.500 ;
        RECT 240.030 358.500 240.210 358.690 ;
        RECT 232.400 358.320 232.720 358.330 ;
        RECT 232.390 358.300 232.720 358.320 ;
        RECT 170.040 357.850 170.300 357.990 ;
        RECT 214.020 357.950 214.210 358.270 ;
        RECT 228.110 357.950 228.300 358.270 ;
        RECT 232.390 357.990 232.560 358.300 ;
        RECT 214.020 357.860 214.300 357.950 ;
        RECT 167.060 357.680 167.820 357.850 ;
        RECT 168.070 357.680 169.240 357.850 ;
        RECT 169.480 357.820 170.300 357.850 ;
        RECT 169.480 357.680 170.590 357.820 ;
        RECT 168.470 357.580 168.820 357.680 ;
        RECT 170.130 357.650 170.590 357.680 ;
        RECT 171.040 357.650 172.230 357.820 ;
        RECT 171.080 357.630 172.230 357.650 ;
        RECT 172.060 357.590 172.230 357.630 ;
        RECT 172.750 357.320 172.920 357.740 ;
        RECT 173.560 357.620 173.800 357.650 ;
        RECT 173.230 357.450 173.800 357.620 ;
        RECT 174.040 357.450 175.380 357.620 ;
        RECT 175.830 357.450 176.790 357.620 ;
        RECT 173.560 357.410 173.800 357.450 ;
        RECT 176.340 357.440 176.510 357.450 ;
        RECT 169.860 357.240 170.250 357.290 ;
        RECT 169.510 357.180 170.250 357.240 ;
        RECT 169.510 357.120 170.330 357.180 ;
        RECT 169.520 357.070 170.330 357.120 ;
        RECT 169.860 357.010 170.330 357.070 ;
        RECT 170.800 357.030 171.760 357.200 ;
        RECT 172.680 357.100 172.850 357.140 ;
        RECT 169.860 357.000 170.240 357.010 ;
        RECT 166.470 356.910 166.640 356.960 ;
        RECT 166.440 356.690 166.660 356.910 ;
        RECT 170.070 356.770 170.240 357.000 ;
        RECT 166.470 356.630 166.640 356.690 ;
        RECT 166.990 356.550 167.320 356.730 ;
        RECT 170.070 356.720 170.300 356.770 ;
        RECT 167.570 356.550 169.730 356.720 ;
        RECT 169.970 356.550 170.300 356.720 ;
        RECT 170.590 356.580 170.800 356.910 ;
        RECT 171.040 356.560 171.220 356.850 ;
        RECT 171.580 356.570 171.760 357.030 ;
        RECT 172.620 356.930 172.850 357.100 ;
        RECT 175.970 357.000 176.310 357.180 ;
        RECT 171.770 356.580 172.390 356.750 ;
        RECT 172.680 356.580 172.850 356.930 ;
        RECT 172.920 356.710 173.110 356.940 ;
        RECT 173.210 356.830 173.580 357.000 ;
        RECT 174.040 356.830 176.790 357.000 ;
        RECT 177.320 356.760 177.490 357.690 ;
        RECT 177.720 356.850 177.890 357.740 ;
        RECT 210.660 357.720 214.300 357.860 ;
        RECT 228.020 357.860 228.300 357.950 ;
        RECT 228.020 357.720 231.660 357.860 ;
        RECT 233.460 357.800 233.630 358.080 ;
        RECT 234.810 358.020 234.980 358.050 ;
        RECT 236.500 358.020 236.670 358.350 ;
        RECT 236.820 358.310 237.020 358.500 ;
        RECT 236.680 358.170 237.020 358.310 ;
        RECT 236.680 358.090 237.010 358.170 ;
        RECT 236.680 358.050 237.000 358.090 ;
        RECT 234.810 357.990 235.140 358.020 ;
        RECT 234.810 357.800 235.150 357.990 ;
        RECT 235.420 357.940 235.800 358.000 ;
        RECT 235.420 357.830 235.980 357.940 ;
        RECT 235.670 357.820 235.980 357.830 ;
        RECT 233.460 357.760 233.670 357.800 ;
        RECT 234.810 357.760 235.140 357.800 ;
        RECT 233.460 357.740 233.690 357.760 ;
        RECT 234.810 357.750 234.980 357.760 ;
        RECT 210.660 357.680 214.210 357.720 ;
        RECT 214.020 357.260 214.210 357.680 ;
        RECT 228.110 357.680 231.660 357.720 ;
        RECT 232.550 357.690 232.870 357.730 ;
        RECT 228.110 357.260 228.300 357.680 ;
        RECT 232.540 357.500 232.870 357.690 ;
        RECT 233.460 357.720 233.720 357.740 ;
        RECT 233.460 357.670 233.800 357.720 ;
        RECT 235.790 357.710 235.980 357.820 ;
        RECT 233.460 357.610 233.950 357.670 ;
        RECT 236.820 357.660 237.020 357.840 ;
        RECT 236.730 357.630 237.050 357.660 ;
        RECT 233.460 357.580 233.970 357.610 ;
        RECT 233.500 357.550 233.970 357.580 ;
        RECT 233.630 357.500 233.970 357.550 ;
        RECT 232.550 357.470 232.870 357.500 ;
        RECT 233.750 357.490 233.970 357.500 ;
        RECT 233.760 357.460 233.970 357.490 ;
        RECT 233.780 357.380 233.970 357.460 ;
        RECT 235.140 357.380 235.470 357.500 ;
        RECT 236.730 357.440 237.060 357.630 ;
        RECT 237.410 357.510 237.960 358.500 ;
        RECT 238.430 357.940 239.140 358.080 ;
        RECT 238.430 357.910 239.260 357.940 ;
        RECT 238.780 357.900 239.260 357.910 ;
        RECT 238.780 357.710 239.270 357.900 ;
        RECT 238.780 357.680 239.260 357.710 ;
        RECT 238.780 357.630 239.140 357.680 ;
        RECT 238.780 357.460 239.110 357.630 ;
        RECT 236.730 357.400 237.050 357.440 ;
        RECT 233.780 357.330 234.300 357.380 ;
        RECT 233.880 357.210 234.300 357.330 ;
        RECT 202.110 356.940 202.290 357.130 ;
        RECT 233.880 357.100 234.070 357.210 ;
        RECT 234.650 357.200 235.910 357.380 ;
        RECT 239.220 357.370 239.550 357.540 ;
        RECT 233.380 357.070 233.550 357.090 ;
        RECT 238.970 357.080 239.290 357.100 ;
        RECT 167.020 356.110 167.290 356.550 ;
        RECT 168.500 356.290 168.830 356.550 ;
        RECT 169.450 356.510 169.740 356.550 ;
        RECT 169.410 356.340 169.740 356.510 ;
        RECT 169.450 356.310 169.740 356.340 ;
        RECT 170.040 356.410 170.300 356.550 ;
        RECT 170.440 356.410 171.220 356.560 ;
        RECT 167.060 356.100 167.290 356.110 ;
        RECT 170.040 356.240 171.220 356.410 ;
        RECT 171.500 356.400 171.830 356.570 ;
        RECT 170.040 356.100 170.300 356.240 ;
        RECT 167.060 355.930 167.820 356.100 ;
        RECT 168.070 355.930 169.240 356.100 ;
        RECT 169.480 356.070 170.300 356.100 ;
        RECT 169.480 355.930 170.590 356.070 ;
        RECT 168.470 355.830 168.820 355.930 ;
        RECT 170.130 355.900 170.590 355.930 ;
        RECT 171.040 355.900 172.230 356.070 ;
        RECT 171.080 355.880 172.230 355.900 ;
        RECT 172.060 355.840 172.230 355.880 ;
        RECT 172.680 355.820 172.850 356.170 ;
        RECT 201.640 356.130 201.930 356.460 ;
        RECT 172.620 355.650 172.850 355.820 ;
        RECT 172.920 355.810 173.110 356.040 ;
        RECT 173.210 355.750 173.580 355.920 ;
        RECT 174.040 355.750 176.790 355.920 ;
        RECT 172.680 355.610 172.850 355.650 ;
        RECT 175.970 355.570 176.310 355.750 ;
        RECT 169.860 355.490 170.250 355.540 ;
        RECT 169.510 355.430 170.250 355.490 ;
        RECT 169.510 355.370 170.330 355.430 ;
        RECT 169.520 355.320 170.330 355.370 ;
        RECT 169.860 355.260 170.330 355.320 ;
        RECT 170.800 355.280 171.760 355.450 ;
        RECT 169.860 355.250 170.240 355.260 ;
        RECT 166.470 355.160 166.640 355.210 ;
        RECT 166.440 354.940 166.660 355.160 ;
        RECT 170.070 355.020 170.240 355.250 ;
        RECT 166.470 354.880 166.640 354.940 ;
        RECT 166.990 354.800 167.320 354.980 ;
        RECT 170.070 354.970 170.300 355.020 ;
        RECT 167.570 354.800 169.730 354.970 ;
        RECT 169.970 354.800 170.300 354.970 ;
        RECT 170.590 354.830 170.800 355.160 ;
        RECT 171.040 354.810 171.220 355.100 ;
        RECT 171.580 354.820 171.760 355.280 ;
        RECT 172.750 355.010 172.920 355.430 ;
        RECT 173.560 355.300 173.800 355.340 ;
        RECT 176.340 355.300 176.510 355.310 ;
        RECT 173.230 355.130 173.800 355.300 ;
        RECT 174.040 355.130 175.380 355.300 ;
        RECT 175.830 355.130 176.790 355.300 ;
        RECT 173.560 355.100 173.800 355.130 ;
        RECT 177.320 355.060 177.490 355.990 ;
        RECT 177.720 355.010 177.890 355.900 ;
        RECT 201.720 355.840 201.920 356.130 ;
        RECT 201.730 355.830 201.920 355.840 ;
        RECT 201.350 355.660 201.560 355.670 ;
        RECT 201.350 355.080 201.570 355.660 ;
        RECT 202.120 355.330 202.290 356.940 ;
        RECT 202.950 355.340 203.120 357.030 ;
        RECT 231.740 356.870 232.060 356.900 ;
        RECT 207.580 356.700 207.900 356.740 ;
        RECT 207.570 356.510 207.900 356.700 ;
        RECT 231.740 356.680 232.070 356.870 ;
        RECT 207.580 356.480 207.900 356.510 ;
        RECT 212.950 355.950 213.180 356.680 ;
        RECT 214.870 356.180 215.190 356.220 ;
        RECT 214.860 355.990 215.190 356.180 ;
        RECT 214.870 355.960 215.190 355.990 ;
        RECT 214.990 355.820 215.010 355.960 ;
        RECT 229.140 355.950 229.370 356.680 ;
        RECT 231.740 356.640 232.060 356.680 ;
        RECT 233.360 356.640 233.570 357.070 ;
        RECT 236.720 357.040 237.040 357.080 ;
        RECT 236.720 356.850 237.050 357.040 ;
        RECT 238.970 356.990 239.540 357.080 ;
        RECT 236.720 356.820 237.040 356.850 ;
        RECT 234.420 356.700 234.740 356.740 ;
        RECT 234.420 356.510 234.750 356.700 ;
        RECT 236.810 356.640 237.010 356.820 ;
        RECT 234.420 356.480 234.740 356.510 ;
        RECT 233.740 356.210 233.910 356.240 ;
        RECT 233.740 356.180 234.140 356.210 ;
        RECT 233.740 355.990 234.150 356.180 ;
        RECT 234.400 356.140 234.690 356.190 ;
        RECT 234.350 356.020 234.690 356.140 ;
        RECT 214.990 355.740 215.340 355.820 ;
        RECT 201.350 355.050 201.560 355.080 ;
        RECT 171.770 354.830 172.390 355.000 ;
        RECT 167.020 354.360 167.290 354.800 ;
        RECT 168.500 354.540 168.830 354.800 ;
        RECT 169.450 354.760 169.740 354.800 ;
        RECT 169.410 354.590 169.740 354.760 ;
        RECT 169.450 354.560 169.740 354.590 ;
        RECT 170.040 354.660 170.300 354.800 ;
        RECT 170.440 354.660 171.220 354.810 ;
        RECT 167.060 354.350 167.290 354.360 ;
        RECT 170.040 354.490 171.220 354.660 ;
        RECT 171.500 354.650 171.830 354.820 ;
        RECT 201.360 354.700 201.560 355.050 ;
        RECT 202.840 354.780 203.370 354.950 ;
        RECT 210.290 354.890 215.340 355.740 ;
        RECT 231.720 354.920 231.900 355.980 ;
        RECT 233.740 355.950 234.140 355.990 ;
        RECT 233.740 355.940 233.910 355.950 ;
        RECT 234.350 355.910 234.540 356.020 ;
        RECT 232.470 355.590 232.790 355.620 ;
        RECT 234.970 355.600 235.140 356.280 ;
        RECT 236.490 356.130 236.660 356.460 ;
        RECT 236.670 356.390 236.990 356.430 ;
        RECT 236.670 356.310 237.000 356.390 ;
        RECT 236.670 356.170 237.010 356.310 ;
        RECT 236.810 355.980 237.010 356.170 ;
        RECT 237.400 355.980 237.950 356.970 ;
        RECT 238.770 356.910 239.540 356.990 ;
        RECT 240.030 356.940 240.210 357.130 ;
        RECT 238.770 356.840 239.370 356.910 ;
        RECT 238.770 356.820 239.100 356.840 ;
        RECT 238.770 356.540 239.130 356.820 ;
        RECT 238.420 356.370 239.130 356.540 ;
        RECT 238.420 355.700 239.120 355.930 ;
        RECT 232.470 355.520 232.800 355.590 ;
        RECT 232.330 355.400 232.800 355.520 ;
        RECT 232.330 355.390 232.790 355.400 ;
        RECT 233.340 355.390 233.980 355.570 ;
        RECT 234.360 355.390 234.710 355.560 ;
        RECT 234.890 355.520 235.140 355.600 ;
        RECT 234.810 355.400 235.140 355.520 ;
        RECT 238.370 355.470 239.120 355.700 ;
        RECT 232.450 355.360 232.790 355.390 ;
        RECT 232.450 355.290 232.500 355.360 ;
        RECT 234.810 355.290 235.000 355.400 ;
        RECT 232.370 354.960 232.540 355.290 ;
        RECT 236.490 354.990 236.660 355.320 ;
        RECT 236.810 355.280 237.010 355.470 ;
        RECT 236.670 355.140 237.010 355.280 ;
        RECT 236.670 355.060 237.000 355.140 ;
        RECT 236.670 355.020 236.990 355.060 ;
        RECT 232.770 354.760 232.850 354.840 ;
        RECT 232.910 354.760 233.100 354.880 ;
        RECT 232.770 354.670 233.100 354.760 ;
        RECT 232.910 354.650 233.100 354.670 ;
        RECT 236.810 354.630 237.010 354.810 ;
        RECT 236.720 354.600 237.040 354.630 ;
        RECT 170.040 354.350 170.300 354.490 ;
        RECT 236.720 354.410 237.050 354.600 ;
        RECT 237.400 354.480 237.950 355.470 ;
        RECT 238.420 355.050 239.120 355.470 ;
        RECT 239.200 355.340 239.370 356.840 ;
        RECT 240.030 355.330 240.200 356.940 ;
        RECT 240.390 356.130 240.680 356.460 ;
        RECT 240.400 355.840 240.600 356.130 ;
        RECT 240.400 355.830 240.590 355.840 ;
        RECT 240.760 355.660 240.970 355.670 ;
        RECT 240.750 355.080 240.970 355.660 ;
        RECT 240.760 355.050 240.970 355.080 ;
        RECT 238.950 354.780 239.480 354.950 ;
        RECT 239.020 354.650 239.350 354.780 ;
        RECT 240.760 354.700 240.960 355.050 ;
        RECT 239.020 354.630 239.340 354.650 ;
        RECT 238.410 354.620 239.340 354.630 ;
        RECT 238.410 354.450 239.110 354.620 ;
        RECT 167.060 354.180 167.820 354.350 ;
        RECT 168.070 354.180 169.240 354.350 ;
        RECT 169.480 354.320 170.300 354.350 ;
        RECT 169.480 354.180 170.590 354.320 ;
        RECT 168.470 354.080 168.820 354.180 ;
        RECT 170.130 354.150 170.590 354.180 ;
        RECT 171.040 354.150 172.230 354.320 ;
        RECT 171.080 354.130 172.230 354.150 ;
        RECT 172.060 354.090 172.230 354.130 ;
        RECT 218.170 353.390 218.370 354.400 ;
        RECT 223.920 353.390 224.210 354.400 ;
        RECT 236.720 354.370 237.040 354.410 ;
        RECT 239.010 354.120 239.330 354.160 ;
        RECT 236.720 354.040 237.040 354.080 ;
        RECT 236.720 353.850 237.050 354.040 ;
        RECT 239.010 353.970 239.340 354.120 ;
        RECT 236.720 353.820 237.040 353.850 ;
        RECT 236.810 353.640 237.010 353.820 ;
        RECT 232.390 352.490 232.710 352.530 ;
        RECT 187.010 351.920 187.560 352.350 ;
        RECT 191.040 351.990 191.590 352.420 ;
        RECT 221.370 351.990 221.920 352.420 ;
        RECT 225.400 351.920 225.950 352.350 ;
        RECT 232.380 352.300 232.710 352.490 ;
        RECT 232.390 352.290 232.710 352.300 ;
        RECT 232.380 352.270 232.710 352.290 ;
        RECT 232.380 351.960 232.550 352.270 ;
        RECT 232.540 351.660 232.860 351.700 ;
        RECT 232.530 351.470 232.860 351.660 ;
        RECT 235.350 351.490 235.530 353.540 ;
        RECT 236.080 353.280 236.410 353.450 ;
        RECT 236.160 351.500 236.330 353.280 ;
        RECT 236.490 353.130 236.660 353.460 ;
        RECT 236.670 353.390 236.990 353.430 ;
        RECT 236.670 353.310 237.000 353.390 ;
        RECT 236.670 353.170 237.010 353.310 ;
        RECT 236.810 352.980 237.010 353.170 ;
        RECT 237.400 352.980 237.950 353.970 ;
        RECT 238.410 353.930 239.340 353.970 ;
        RECT 238.410 353.900 239.330 353.930 ;
        RECT 238.410 353.790 239.110 353.900 ;
        RECT 238.420 353.110 239.120 353.370 ;
        RECT 238.370 352.880 239.120 353.110 ;
        RECT 238.420 352.490 239.120 352.880 ;
        RECT 236.490 351.990 236.660 352.320 ;
        RECT 236.810 352.280 237.010 352.470 ;
        RECT 236.670 352.140 237.010 352.280 ;
        RECT 236.670 352.060 237.000 352.140 ;
        RECT 236.670 352.020 236.990 352.060 ;
        RECT 236.810 351.630 237.010 351.810 ;
        RECT 236.720 351.600 237.040 351.630 ;
        RECT 232.540 351.440 232.860 351.470 ;
        RECT 236.720 351.410 237.050 351.600 ;
        RECT 237.400 351.480 237.950 352.470 ;
        RECT 238.420 351.910 239.130 352.050 ;
        RECT 238.420 351.880 239.250 351.910 ;
        RECT 238.770 351.870 239.250 351.880 ;
        RECT 238.770 351.680 239.260 351.870 ;
        RECT 238.770 351.650 239.250 351.680 ;
        RECT 238.770 351.600 239.130 351.650 ;
        RECT 238.770 351.430 239.100 351.600 ;
        RECT 236.720 351.370 237.040 351.410 ;
        RECT 239.210 351.340 239.540 351.510 ;
        RECT 231.730 350.840 232.050 350.870 ;
        RECT 198.420 350.710 198.740 350.750 ;
        RECT 169.860 350.610 170.250 350.660 ;
        RECT 169.510 350.550 170.250 350.610 ;
        RECT 169.510 350.490 170.330 350.550 ;
        RECT 169.520 350.440 170.330 350.490 ;
        RECT 169.860 350.380 170.330 350.440 ;
        RECT 170.800 350.400 171.760 350.570 ;
        RECT 169.860 350.370 170.240 350.380 ;
        RECT 166.470 350.280 166.640 350.330 ;
        RECT 166.440 350.060 166.660 350.280 ;
        RECT 170.070 350.140 170.240 350.370 ;
        RECT 166.470 350.000 166.640 350.060 ;
        RECT 166.990 349.920 167.320 350.100 ;
        RECT 170.070 350.090 170.300 350.140 ;
        RECT 167.570 349.920 169.730 350.090 ;
        RECT 169.970 349.920 170.300 350.090 ;
        RECT 170.590 349.950 170.800 350.280 ;
        RECT 171.040 349.930 171.220 350.220 ;
        RECT 171.580 349.940 171.760 350.400 ;
        RECT 171.770 349.950 172.390 350.120 ;
        RECT 172.730 350.050 172.900 350.470 ;
        RECT 173.540 350.350 173.780 350.380 ;
        RECT 173.210 350.180 173.780 350.350 ;
        RECT 174.020 350.180 175.360 350.350 ;
        RECT 175.810 350.180 176.770 350.350 ;
        RECT 173.540 350.140 173.780 350.180 ;
        RECT 176.320 350.170 176.490 350.180 ;
        RECT 167.020 349.480 167.290 349.920 ;
        RECT 168.500 349.660 168.830 349.920 ;
        RECT 169.450 349.880 169.740 349.920 ;
        RECT 169.410 349.710 169.740 349.880 ;
        RECT 169.450 349.680 169.740 349.710 ;
        RECT 170.040 349.780 170.300 349.920 ;
        RECT 170.440 349.780 171.220 349.930 ;
        RECT 167.060 349.470 167.290 349.480 ;
        RECT 170.040 349.610 171.220 349.780 ;
        RECT 171.500 349.770 171.830 349.940 ;
        RECT 172.660 349.830 172.830 349.870 ;
        RECT 172.600 349.660 172.830 349.830 ;
        RECT 175.950 349.730 176.290 349.910 ;
        RECT 170.040 349.470 170.300 349.610 ;
        RECT 167.060 349.300 167.820 349.470 ;
        RECT 168.070 349.300 169.240 349.470 ;
        RECT 169.480 349.440 170.300 349.470 ;
        RECT 169.480 349.300 170.590 349.440 ;
        RECT 168.470 349.200 168.820 349.300 ;
        RECT 170.130 349.270 170.590 349.300 ;
        RECT 171.040 349.270 172.230 349.440 ;
        RECT 172.660 349.310 172.830 349.660 ;
        RECT 172.900 349.440 173.090 349.670 ;
        RECT 173.190 349.560 173.560 349.730 ;
        RECT 174.020 349.560 176.770 349.730 ;
        RECT 177.300 349.490 177.470 350.420 ;
        RECT 177.700 349.580 177.870 350.470 ;
        RECT 196.820 350.320 197.020 350.670 ;
        RECT 198.410 350.590 198.740 350.710 ;
        RECT 198.300 350.490 198.740 350.590 ;
        RECT 214.220 350.710 214.540 350.750 ;
        RECT 214.220 350.590 214.550 350.710 ;
        RECT 214.220 350.490 214.660 350.590 ;
        RECT 198.300 350.420 198.640 350.490 ;
        RECT 214.320 350.420 214.660 350.490 ;
        RECT 196.810 350.290 197.020 350.320 ;
        RECT 215.940 350.320 216.140 350.670 ;
        RECT 231.730 350.650 232.060 350.840 ;
        RECT 231.730 350.610 232.050 350.650 ;
        RECT 196.810 349.700 197.030 350.290 ;
        RECT 197.550 349.700 197.750 350.300 ;
        RECT 198.420 350.160 198.740 350.200 ;
        RECT 198.410 349.970 198.740 350.160 ;
        RECT 198.300 349.940 198.740 349.970 ;
        RECT 214.220 350.160 214.540 350.200 ;
        RECT 214.220 349.970 214.550 350.160 ;
        RECT 214.220 349.940 214.660 349.970 ;
        RECT 198.300 349.800 198.640 349.940 ;
        RECT 214.320 349.800 214.660 349.940 ;
        RECT 215.210 349.700 215.410 350.300 ;
        RECT 215.940 350.290 216.150 350.320 ;
        RECT 215.930 349.700 216.150 350.290 ;
        RECT 171.080 349.250 172.230 349.270 ;
        RECT 172.060 349.210 172.230 349.250 ;
        RECT 11.250 348.920 11.770 348.940 ;
        RECT 5.200 347.440 10.910 347.450 ;
        RECT 5.120 347.270 10.910 347.440 ;
        RECT 5.210 347.260 10.910 347.270 ;
        RECT 10.680 347.190 10.850 347.260 ;
        RECT 11.250 347.140 11.780 348.920 ;
        RECT 169.860 348.860 170.250 348.910 ;
        RECT 169.510 348.800 170.250 348.860 ;
        RECT 169.510 348.740 170.330 348.800 ;
        RECT 169.520 348.690 170.330 348.740 ;
        RECT 169.860 348.630 170.330 348.690 ;
        RECT 170.800 348.650 171.760 348.820 ;
        RECT 169.860 348.620 170.240 348.630 ;
        RECT 166.470 348.530 166.640 348.580 ;
        RECT 166.440 348.310 166.660 348.530 ;
        RECT 170.070 348.390 170.240 348.620 ;
        RECT 166.470 348.250 166.640 348.310 ;
        RECT 166.990 348.170 167.320 348.350 ;
        RECT 170.070 348.340 170.300 348.390 ;
        RECT 167.570 348.170 169.730 348.340 ;
        RECT 169.970 348.170 170.300 348.340 ;
        RECT 170.590 348.200 170.800 348.530 ;
        RECT 171.040 348.180 171.220 348.470 ;
        RECT 171.580 348.190 171.760 348.650 ;
        RECT 172.660 348.550 172.830 348.900 ;
        RECT 172.600 348.380 172.830 348.550 ;
        RECT 172.900 348.540 173.090 348.770 ;
        RECT 173.190 348.480 173.560 348.650 ;
        RECT 174.020 348.480 176.770 348.650 ;
        RECT 171.770 348.200 172.390 348.370 ;
        RECT 172.660 348.340 172.830 348.380 ;
        RECT 175.950 348.300 176.290 348.480 ;
        RECT 167.020 347.730 167.290 348.170 ;
        RECT 168.500 347.910 168.830 348.170 ;
        RECT 169.450 348.130 169.740 348.170 ;
        RECT 169.410 347.960 169.740 348.130 ;
        RECT 169.450 347.930 169.740 347.960 ;
        RECT 170.040 348.030 170.300 348.170 ;
        RECT 170.440 348.030 171.220 348.180 ;
        RECT 167.060 347.720 167.290 347.730 ;
        RECT 170.040 347.860 171.220 348.030 ;
        RECT 171.500 348.020 171.830 348.190 ;
        RECT 170.040 347.720 170.300 347.860 ;
        RECT 172.730 347.740 172.900 348.160 ;
        RECT 173.540 348.030 173.780 348.070 ;
        RECT 176.320 348.030 176.490 348.040 ;
        RECT 173.210 347.860 173.780 348.030 ;
        RECT 174.020 347.860 175.360 348.030 ;
        RECT 175.810 347.860 176.770 348.030 ;
        RECT 173.540 347.830 173.780 347.860 ;
        RECT 177.300 347.790 177.470 348.720 ;
        RECT 177.700 347.740 177.870 348.630 ;
        RECT 196.810 348.560 197.030 349.150 ;
        RECT 196.810 348.530 197.020 348.560 ;
        RECT 197.550 348.550 197.750 349.150 ;
        RECT 199.560 349.070 199.730 349.600 ;
        RECT 203.500 349.080 203.670 349.610 ;
        RECT 209.290 349.080 209.460 349.610 ;
        RECT 213.230 349.070 213.400 349.600 ;
        RECT 198.300 348.910 198.640 349.050 ;
        RECT 214.320 348.910 214.660 349.050 ;
        RECT 198.300 348.880 198.740 348.910 ;
        RECT 198.410 348.690 198.740 348.880 ;
        RECT 198.420 348.650 198.740 348.690 ;
        RECT 214.220 348.880 214.660 348.910 ;
        RECT 214.220 348.690 214.550 348.880 ;
        RECT 214.220 348.650 214.540 348.690 ;
        RECT 215.210 348.550 215.410 349.150 ;
        RECT 215.930 348.560 216.150 349.150 ;
        RECT 231.710 348.890 231.890 349.950 ;
        RECT 232.460 349.560 232.780 349.590 ;
        RECT 232.460 349.490 232.790 349.560 ;
        RECT 232.320 349.370 232.790 349.490 ;
        RECT 232.320 349.360 232.780 349.370 ;
        RECT 232.440 349.330 232.780 349.360 ;
        RECT 232.440 349.260 232.490 349.330 ;
        RECT 232.360 348.930 232.530 349.260 ;
        RECT 232.760 348.730 232.840 348.810 ;
        RECT 232.900 348.730 233.090 348.850 ;
        RECT 232.760 348.640 233.090 348.730 ;
        RECT 232.900 348.620 233.090 348.640 ;
        RECT 196.820 348.180 197.020 348.530 ;
        RECT 215.940 348.530 216.150 348.560 ;
        RECT 198.300 348.360 198.640 348.430 ;
        RECT 198.300 348.260 198.740 348.360 ;
        RECT 198.410 348.140 198.740 348.260 ;
        RECT 198.420 348.100 198.740 348.140 ;
        RECT 197.190 347.720 197.630 347.890 ;
        RECT 167.060 347.550 167.820 347.720 ;
        RECT 168.070 347.550 169.240 347.720 ;
        RECT 169.480 347.690 170.300 347.720 ;
        RECT 169.480 347.550 170.590 347.690 ;
        RECT 168.470 347.450 168.820 347.550 ;
        RECT 170.130 347.520 170.590 347.550 ;
        RECT 171.040 347.520 172.230 347.690 ;
        RECT 171.080 347.500 172.230 347.520 ;
        RECT 172.060 347.460 172.230 347.500 ;
        RECT 198.420 347.470 198.740 347.510 ;
        RECT 11.260 347.120 11.780 347.140 ;
        RECT 4.240 346.400 6.680 346.690 ;
        RECT 11.260 346.610 11.770 347.120 ;
        RECT 169.860 347.110 170.250 347.160 ;
        RECT 169.510 347.050 170.250 347.110 ;
        RECT 169.510 346.990 170.330 347.050 ;
        RECT 169.520 346.940 170.330 346.990 ;
        RECT 169.860 346.880 170.330 346.940 ;
        RECT 170.800 346.900 171.760 347.070 ;
        RECT 169.860 346.870 170.240 346.880 ;
        RECT 166.470 346.780 166.640 346.830 ;
        RECT 11.260 346.400 11.790 346.610 ;
        RECT 166.440 346.560 166.660 346.780 ;
        RECT 170.070 346.640 170.240 346.870 ;
        RECT 166.470 346.500 166.640 346.560 ;
        RECT 166.990 346.420 167.320 346.600 ;
        RECT 170.070 346.590 170.300 346.640 ;
        RECT 167.570 346.420 169.730 346.590 ;
        RECT 169.970 346.420 170.300 346.590 ;
        RECT 170.590 346.450 170.800 346.780 ;
        RECT 171.040 346.430 171.220 346.720 ;
        RECT 171.580 346.440 171.760 346.900 ;
        RECT 172.730 346.850 172.900 347.270 ;
        RECT 173.540 347.150 173.780 347.180 ;
        RECT 173.210 346.980 173.780 347.150 ;
        RECT 174.020 346.980 175.360 347.150 ;
        RECT 175.810 346.980 176.770 347.150 ;
        RECT 173.540 346.940 173.780 346.980 ;
        RECT 176.320 346.970 176.490 346.980 ;
        RECT 172.660 346.630 172.830 346.670 ;
        RECT 171.770 346.450 172.390 346.620 ;
        RECT 172.600 346.460 172.830 346.630 ;
        RECT 175.950 346.530 176.290 346.710 ;
        RECT 4.240 345.920 11.790 346.400 ;
        RECT 167.020 345.980 167.290 346.420 ;
        RECT 168.500 346.160 168.830 346.420 ;
        RECT 169.450 346.380 169.740 346.420 ;
        RECT 169.410 346.210 169.740 346.380 ;
        RECT 169.450 346.180 169.740 346.210 ;
        RECT 170.040 346.280 170.300 346.420 ;
        RECT 170.440 346.280 171.220 346.430 ;
        RECT 167.060 345.970 167.290 345.980 ;
        RECT 170.040 346.110 171.220 346.280 ;
        RECT 171.500 346.270 171.830 346.440 ;
        RECT 172.660 346.110 172.830 346.460 ;
        RECT 172.900 346.240 173.090 346.470 ;
        RECT 173.190 346.360 173.560 346.530 ;
        RECT 174.020 346.360 176.770 346.530 ;
        RECT 177.300 346.290 177.470 347.220 ;
        RECT 177.700 346.380 177.870 347.270 ;
        RECT 184.970 346.900 185.520 347.330 ;
        RECT 189.000 346.970 189.550 347.400 ;
        RECT 196.820 347.080 197.020 347.430 ;
        RECT 198.410 347.350 198.740 347.470 ;
        RECT 198.300 347.250 198.740 347.350 ;
        RECT 198.300 347.180 198.640 347.250 ;
        RECT 199.560 347.230 199.730 348.240 ;
        RECT 203.490 347.370 203.660 348.380 ;
        RECT 209.300 347.370 209.470 348.380 ;
        RECT 214.320 348.360 214.660 348.430 ;
        RECT 214.220 348.260 214.660 348.360 ;
        RECT 213.230 347.230 213.400 348.240 ;
        RECT 214.220 348.140 214.550 348.260 ;
        RECT 215.940 348.180 216.140 348.530 ;
        RECT 235.350 348.440 235.530 350.490 ;
        RECT 236.080 350.230 236.410 350.400 ;
        RECT 236.160 348.450 236.330 350.230 ;
        RECT 214.220 348.100 214.540 348.140 ;
        RECT 215.330 347.720 215.770 347.890 ;
        RECT 214.220 347.470 214.540 347.510 ;
        RECT 214.220 347.350 214.550 347.470 ;
        RECT 214.220 347.250 214.660 347.350 ;
        RECT 214.320 347.180 214.660 347.250 ;
        RECT 196.810 347.050 197.020 347.080 ;
        RECT 215.940 347.080 216.140 347.430 ;
        RECT 196.810 346.460 197.030 347.050 ;
        RECT 197.550 346.460 197.750 347.060 ;
        RECT 198.420 346.920 198.740 346.960 ;
        RECT 198.410 346.730 198.740 346.920 ;
        RECT 198.300 346.700 198.740 346.730 ;
        RECT 214.220 346.920 214.540 346.960 ;
        RECT 214.220 346.730 214.550 346.920 ;
        RECT 214.220 346.700 214.660 346.730 ;
        RECT 198.300 346.560 198.640 346.700 ;
        RECT 214.320 346.560 214.660 346.700 ;
        RECT 215.210 346.460 215.410 347.060 ;
        RECT 215.940 347.050 216.150 347.080 ;
        RECT 215.930 346.460 216.150 347.050 ;
        RECT 170.040 345.970 170.300 346.110 ;
        RECT 4.240 345.890 11.600 345.920 ;
        RECT 167.060 345.800 167.820 345.970 ;
        RECT 168.070 345.800 169.240 345.970 ;
        RECT 169.480 345.940 170.300 345.970 ;
        RECT 169.480 345.800 170.590 345.940 ;
        RECT 168.470 345.700 168.820 345.800 ;
        RECT 170.130 345.770 170.590 345.800 ;
        RECT 171.040 345.770 172.230 345.940 ;
        RECT 171.080 345.750 172.230 345.770 ;
        RECT 172.060 345.710 172.230 345.750 ;
        RECT 196.380 345.730 196.700 345.770 ;
        RECT 169.860 345.360 170.250 345.410 ;
        RECT 169.510 345.300 170.250 345.360 ;
        RECT 172.660 345.350 172.830 345.700 ;
        RECT 169.510 345.240 170.330 345.300 ;
        RECT 169.520 345.190 170.330 345.240 ;
        RECT 169.860 345.130 170.330 345.190 ;
        RECT 170.800 345.150 171.760 345.320 ;
        RECT 172.600 345.180 172.830 345.350 ;
        RECT 172.900 345.340 173.090 345.570 ;
        RECT 173.190 345.280 173.560 345.450 ;
        RECT 174.020 345.280 176.770 345.450 ;
        RECT 169.860 345.120 170.240 345.130 ;
        RECT 166.470 345.030 166.640 345.080 ;
        RECT 166.440 344.810 166.660 345.030 ;
        RECT 170.070 344.890 170.240 345.120 ;
        RECT 166.470 344.750 166.640 344.810 ;
        RECT 4.240 344.130 11.770 344.680 ;
        RECT 166.990 344.670 167.320 344.850 ;
        RECT 170.070 344.840 170.300 344.890 ;
        RECT 167.570 344.670 169.730 344.840 ;
        RECT 169.970 344.670 170.300 344.840 ;
        RECT 170.590 344.700 170.800 345.030 ;
        RECT 171.040 344.680 171.220 344.970 ;
        RECT 171.580 344.690 171.760 345.150 ;
        RECT 172.660 345.140 172.830 345.180 ;
        RECT 175.950 345.100 176.290 345.280 ;
        RECT 171.770 344.700 172.390 344.870 ;
        RECT 167.020 344.230 167.290 344.670 ;
        RECT 168.500 344.410 168.830 344.670 ;
        RECT 169.450 344.630 169.740 344.670 ;
        RECT 169.410 344.460 169.740 344.630 ;
        RECT 169.450 344.430 169.740 344.460 ;
        RECT 170.040 344.530 170.300 344.670 ;
        RECT 170.440 344.530 171.220 344.680 ;
        RECT 2.550 331.160 4.030 331.410 ;
        RECT 4.240 331.220 4.750 344.130 ;
        RECT 11.100 344.120 11.770 344.130 ;
        RECT 7.400 343.230 10.860 343.670 ;
        RECT 5.470 343.130 10.860 343.230 ;
        RECT 5.470 343.060 10.750 343.130 ;
        RECT 5.470 332.150 5.640 343.060 ;
        RECT 5.970 342.650 10.200 342.670 ;
        RECT 5.950 332.540 10.280 342.650 ;
        RECT 6.010 332.490 6.180 332.540 ;
        RECT 10.580 332.150 10.750 343.060 ;
        RECT 5.470 331.980 10.750 332.150 ;
        RECT 10.510 331.970 10.750 331.980 ;
        RECT 11.260 331.220 11.770 344.120 ;
        RECT 167.060 344.220 167.290 344.230 ;
        RECT 170.040 344.360 171.220 344.530 ;
        RECT 171.500 344.520 171.830 344.690 ;
        RECT 172.730 344.540 172.900 344.960 ;
        RECT 173.540 344.830 173.780 344.870 ;
        RECT 176.320 344.830 176.490 344.840 ;
        RECT 173.210 344.660 173.780 344.830 ;
        RECT 174.020 344.660 175.360 344.830 ;
        RECT 175.810 344.660 176.770 344.830 ;
        RECT 173.540 344.630 173.780 344.660 ;
        RECT 177.300 344.590 177.470 345.520 ;
        RECT 177.700 344.540 177.870 345.430 ;
        RECT 194.780 345.340 194.980 345.690 ;
        RECT 196.370 345.610 196.700 345.730 ;
        RECT 196.260 345.510 196.700 345.610 ;
        RECT 196.260 345.440 196.600 345.510 ;
        RECT 194.770 345.310 194.980 345.340 ;
        RECT 196.810 345.330 197.030 345.920 ;
        RECT 194.770 344.720 194.990 345.310 ;
        RECT 195.510 344.720 195.710 345.320 ;
        RECT 196.810 345.300 197.020 345.330 ;
        RECT 197.550 345.320 197.750 345.920 ;
        RECT 198.300 345.680 198.640 345.820 ;
        RECT 214.320 345.680 214.660 345.820 ;
        RECT 198.300 345.650 198.740 345.680 ;
        RECT 198.410 345.460 198.740 345.650 ;
        RECT 198.420 345.420 198.740 345.460 ;
        RECT 214.220 345.650 214.660 345.680 ;
        RECT 214.220 345.460 214.550 345.650 ;
        RECT 214.220 345.420 214.540 345.460 ;
        RECT 215.210 345.320 215.410 345.920 ;
        RECT 215.930 345.330 216.150 345.920 ;
        RECT 235.340 345.460 235.520 347.510 ;
        RECT 236.070 347.250 236.400 347.420 ;
        RECT 236.150 345.470 236.320 347.250 ;
        RECT 196.380 345.180 196.700 345.220 ;
        RECT 196.370 344.990 196.700 345.180 ;
        RECT 196.260 344.960 196.700 344.990 ;
        RECT 196.260 344.820 196.600 344.960 ;
        RECT 196.820 344.950 197.020 345.300 ;
        RECT 215.940 345.300 216.150 345.330 ;
        RECT 198.300 345.130 198.640 345.200 ;
        RECT 214.320 345.130 214.660 345.200 ;
        RECT 198.300 345.030 198.740 345.130 ;
        RECT 198.410 344.910 198.740 345.030 ;
        RECT 198.420 344.870 198.740 344.910 ;
        RECT 214.220 345.030 214.660 345.130 ;
        RECT 214.220 344.910 214.550 345.030 ;
        RECT 215.940 344.950 216.140 345.300 ;
        RECT 214.220 344.870 214.540 344.910 ;
        RECT 170.040 344.220 170.300 344.360 ;
        RECT 167.060 344.050 167.820 344.220 ;
        RECT 168.070 344.050 169.240 344.220 ;
        RECT 169.480 344.190 170.300 344.220 ;
        RECT 169.480 344.050 170.590 344.190 ;
        RECT 168.470 343.950 168.820 344.050 ;
        RECT 170.130 344.020 170.590 344.050 ;
        RECT 171.040 344.020 172.230 344.190 ;
        RECT 171.080 344.000 172.230 344.020 ;
        RECT 172.060 343.960 172.230 344.000 ;
        RECT 194.770 343.600 194.990 344.190 ;
        RECT 194.770 343.570 194.980 343.600 ;
        RECT 195.510 343.590 195.710 344.190 ;
        RECT 196.260 343.950 196.600 344.090 ;
        RECT 197.650 344.030 197.820 344.560 ;
        RECT 201.670 344.060 201.840 344.590 ;
        RECT 196.260 343.920 196.700 343.950 ;
        RECT 196.370 343.730 196.700 343.920 ;
        RECT 196.380 343.690 196.700 343.730 ;
        RECT 194.780 343.220 194.980 343.570 ;
        RECT 196.260 343.400 196.600 343.470 ;
        RECT 196.260 343.300 196.700 343.400 ;
        RECT 196.370 343.180 196.700 343.300 ;
        RECT 196.380 343.140 196.700 343.180 ;
        RECT 195.150 342.760 195.590 342.930 ;
        RECT 196.380 342.490 196.700 342.530 ;
        RECT 194.780 342.100 194.980 342.450 ;
        RECT 196.370 342.370 196.700 342.490 ;
        RECT 196.260 342.270 196.700 342.370 ;
        RECT 196.260 342.200 196.600 342.270 ;
        RECT 197.640 342.170 197.810 343.360 ;
        RECT 201.660 342.130 201.830 343.300 ;
        RECT 235.340 342.410 235.520 344.460 ;
        RECT 236.070 344.200 236.400 344.370 ;
        RECT 236.150 342.420 236.320 344.200 ;
        RECT 194.770 342.070 194.980 342.100 ;
        RECT 169.820 341.550 170.210 341.600 ;
        RECT 169.470 341.490 170.210 341.550 ;
        RECT 169.470 341.430 170.290 341.490 ;
        RECT 169.480 341.380 170.290 341.430 ;
        RECT 169.820 341.320 170.290 341.380 ;
        RECT 170.760 341.340 171.720 341.510 ;
        RECT 194.770 341.480 194.990 342.070 ;
        RECT 195.510 341.480 195.710 342.080 ;
        RECT 196.380 341.940 196.700 341.980 ;
        RECT 196.370 341.750 196.700 341.940 ;
        RECT 196.260 341.720 196.700 341.750 ;
        RECT 196.260 341.580 196.600 341.720 ;
        RECT 169.820 341.310 170.200 341.320 ;
        RECT 166.430 341.220 166.600 341.270 ;
        RECT 166.400 341.000 166.620 341.220 ;
        RECT 170.030 341.080 170.200 341.310 ;
        RECT 166.430 340.940 166.600 341.000 ;
        RECT 166.950 340.860 167.280 341.040 ;
        RECT 170.030 341.030 170.260 341.080 ;
        RECT 167.530 340.860 169.690 341.030 ;
        RECT 169.930 340.860 170.260 341.030 ;
        RECT 170.550 340.890 170.760 341.220 ;
        RECT 171.000 340.870 171.180 341.160 ;
        RECT 171.540 340.880 171.720 341.340 ;
        RECT 171.730 340.890 172.350 341.060 ;
        RECT 144.160 339.830 144.330 340.470 ;
        RECT 144.710 339.830 144.880 340.470 ;
        RECT 145.350 340.270 145.520 340.470 ;
        RECT 145.900 340.270 146.070 340.470 ;
        RECT 166.980 340.420 167.250 340.860 ;
        RECT 168.460 340.600 168.790 340.860 ;
        RECT 169.410 340.820 169.700 340.860 ;
        RECT 169.370 340.650 169.700 340.820 ;
        RECT 169.410 340.620 169.700 340.650 ;
        RECT 170.000 340.720 170.260 340.860 ;
        RECT 170.400 340.720 171.180 340.870 ;
        RECT 167.020 340.410 167.250 340.420 ;
        RECT 170.000 340.550 171.180 340.720 ;
        RECT 171.460 340.710 171.790 340.880 ;
        RECT 172.760 340.780 172.930 341.200 ;
        RECT 173.570 341.080 173.810 341.110 ;
        RECT 173.240 340.910 173.810 341.080 ;
        RECT 174.050 340.910 175.390 341.080 ;
        RECT 175.840 340.910 176.800 341.080 ;
        RECT 173.570 340.870 173.810 340.910 ;
        RECT 176.350 340.900 176.520 340.910 ;
        RECT 172.690 340.560 172.860 340.600 ;
        RECT 170.000 340.410 170.260 340.550 ;
        RECT 145.350 340.240 145.690 340.270 ;
        RECT 145.900 340.240 146.340 340.270 ;
        RECT 167.020 340.240 167.780 340.410 ;
        RECT 168.030 340.240 169.200 340.410 ;
        RECT 169.440 340.380 170.260 340.410 ;
        RECT 172.630 340.390 172.860 340.560 ;
        RECT 175.980 340.460 176.320 340.640 ;
        RECT 169.440 340.240 170.550 340.380 ;
        RECT 145.350 340.050 145.700 340.240 ;
        RECT 145.900 340.050 146.350 340.240 ;
        RECT 168.430 340.140 168.780 340.240 ;
        RECT 170.090 340.210 170.550 340.240 ;
        RECT 171.000 340.210 172.190 340.380 ;
        RECT 171.040 340.190 172.190 340.210 ;
        RECT 172.020 340.150 172.190 340.190 ;
        RECT 145.350 340.010 145.690 340.050 ;
        RECT 145.900 340.010 146.340 340.050 ;
        RECT 172.690 340.040 172.860 340.390 ;
        RECT 172.930 340.170 173.120 340.400 ;
        RECT 173.220 340.290 173.590 340.460 ;
        RECT 174.050 340.290 176.800 340.460 ;
        RECT 177.330 340.220 177.500 341.150 ;
        RECT 177.730 340.310 177.900 341.200 ;
        RECT 208.200 341.170 209.660 341.290 ;
        RECT 208.010 341.120 209.660 341.170 ;
        RECT 208.010 340.950 208.340 341.120 ;
        RECT 194.770 340.350 194.990 340.940 ;
        RECT 194.770 340.320 194.980 340.350 ;
        RECT 195.510 340.340 195.710 340.940 ;
        RECT 208.010 340.910 208.330 340.950 ;
        RECT 209.490 340.890 209.660 341.120 ;
        RECT 196.260 340.700 196.600 340.840 ;
        RECT 196.260 340.670 196.700 340.700 ;
        RECT 196.370 340.480 196.700 340.670 ;
        RECT 208.340 340.490 208.680 340.890 ;
        RECT 208.850 340.720 209.180 340.890 ;
        RECT 209.400 340.720 209.740 340.890 ;
        RECT 208.930 340.550 209.100 340.720 ;
        RECT 209.490 340.550 209.660 340.720 ;
        RECT 196.380 340.440 196.700 340.480 ;
        RECT 208.160 340.380 208.680 340.490 ;
        RECT 208.850 340.380 209.180 340.550 ;
        RECT 209.400 340.380 209.740 340.550 ;
        RECT 144.150 339.800 144.470 339.830 ;
        RECT 144.710 339.800 145.170 339.830 ;
        RECT 144.150 339.610 144.480 339.800 ;
        RECT 144.710 339.610 145.180 339.800 ;
        RECT 144.150 339.570 144.470 339.610 ;
        RECT 144.710 339.570 145.170 339.610 ;
        RECT 144.160 338.070 144.330 339.570 ;
        RECT 144.710 338.070 144.880 339.570 ;
        RECT 145.350 338.070 145.520 340.010 ;
        RECT 145.900 338.070 146.070 340.010 ;
        RECT 194.780 339.970 194.980 340.320 ;
        RECT 208.160 340.270 208.490 340.380 ;
        RECT 208.160 340.230 208.480 340.270 ;
        RECT 196.260 340.150 196.600 340.220 ;
        RECT 208.930 340.150 209.180 340.380 ;
        RECT 210.060 340.300 210.570 340.970 ;
        RECT 196.260 340.050 196.700 340.150 ;
        RECT 196.370 339.930 196.700 340.050 ;
        RECT 196.380 339.890 196.700 339.930 ;
        RECT 208.930 339.980 209.600 340.150 ;
        RECT 208.160 339.860 208.480 339.900 ;
        RECT 169.820 339.800 170.210 339.850 ;
        RECT 169.470 339.740 170.210 339.800 ;
        RECT 169.470 339.680 170.290 339.740 ;
        RECT 169.480 339.630 170.290 339.680 ;
        RECT 169.820 339.570 170.290 339.630 ;
        RECT 170.760 339.590 171.720 339.760 ;
        RECT 208.160 339.750 208.490 339.860 ;
        RECT 208.930 339.750 209.180 339.980 ;
        RECT 208.160 339.640 208.680 339.750 ;
        RECT 169.820 339.560 170.200 339.570 ;
        RECT 146.450 338.710 146.620 339.560 ;
        RECT 166.430 339.470 166.600 339.520 ;
        RECT 166.400 339.250 166.620 339.470 ;
        RECT 170.030 339.330 170.200 339.560 ;
        RECT 166.430 339.190 166.600 339.250 ;
        RECT 166.950 339.110 167.280 339.290 ;
        RECT 170.030 339.280 170.260 339.330 ;
        RECT 167.530 339.110 169.690 339.280 ;
        RECT 169.930 339.110 170.260 339.280 ;
        RECT 170.550 339.140 170.760 339.470 ;
        RECT 171.000 339.120 171.180 339.410 ;
        RECT 171.540 339.130 171.720 339.590 ;
        RECT 171.730 339.140 172.350 339.310 ;
        RECT 172.690 339.280 172.860 339.630 ;
        RECT 166.980 338.670 167.250 339.110 ;
        RECT 168.460 338.850 168.790 339.110 ;
        RECT 169.410 339.070 169.700 339.110 ;
        RECT 169.370 338.900 169.700 339.070 ;
        RECT 169.410 338.870 169.700 338.900 ;
        RECT 170.000 338.970 170.260 339.110 ;
        RECT 170.400 338.970 171.180 339.120 ;
        RECT 167.020 338.660 167.250 338.670 ;
        RECT 170.000 338.800 171.180 338.970 ;
        RECT 171.460 338.960 171.790 339.130 ;
        RECT 172.630 339.110 172.860 339.280 ;
        RECT 172.930 339.270 173.120 339.500 ;
        RECT 173.220 339.210 173.590 339.380 ;
        RECT 174.050 339.210 176.800 339.380 ;
        RECT 172.690 339.070 172.860 339.110 ;
        RECT 175.980 339.030 176.320 339.210 ;
        RECT 170.000 338.660 170.260 338.800 ;
        RECT 167.020 338.490 167.780 338.660 ;
        RECT 168.030 338.490 169.200 338.660 ;
        RECT 169.440 338.630 170.260 338.660 ;
        RECT 169.440 338.490 170.550 338.630 ;
        RECT 168.430 338.390 168.780 338.490 ;
        RECT 170.090 338.460 170.550 338.490 ;
        RECT 171.000 338.460 172.190 338.630 ;
        RECT 172.760 338.470 172.930 338.890 ;
        RECT 173.570 338.760 173.810 338.800 ;
        RECT 176.350 338.760 176.520 338.770 ;
        RECT 173.240 338.590 173.810 338.760 ;
        RECT 174.050 338.590 175.390 338.760 ;
        RECT 175.840 338.590 176.800 338.760 ;
        RECT 173.570 338.560 173.810 338.590 ;
        RECT 177.330 338.520 177.500 339.450 ;
        RECT 177.730 338.470 177.900 339.360 ;
        RECT 208.340 339.240 208.680 339.640 ;
        RECT 208.850 339.580 209.180 339.750 ;
        RECT 209.400 339.580 209.740 339.750 ;
        RECT 208.930 339.410 209.100 339.580 ;
        RECT 209.490 339.410 209.660 339.580 ;
        RECT 208.850 339.240 209.180 339.410 ;
        RECT 209.400 339.240 209.740 339.410 ;
        RECT 208.010 339.180 208.330 339.220 ;
        RECT 208.010 339.010 208.340 339.180 ;
        RECT 209.490 339.010 209.660 339.240 ;
        RECT 210.060 339.160 210.570 339.830 ;
        RECT 208.010 338.960 209.660 339.010 ;
        RECT 208.200 338.840 209.660 338.960 ;
        RECT 171.040 338.440 172.190 338.460 ;
        RECT 172.020 338.400 172.190 338.440 ;
        RECT 208.200 338.400 209.660 338.520 ;
        RECT 208.010 338.350 209.660 338.400 ;
        RECT 208.010 338.180 208.340 338.350 ;
        RECT 208.010 338.140 208.330 338.180 ;
        RECT 209.490 338.120 209.660 338.350 ;
        RECT 146.340 338.080 146.770 338.100 ;
        RECT 143.530 338.000 143.700 338.020 ;
        RECT 143.510 337.880 143.720 338.000 ;
        RECT 146.340 337.910 146.790 338.080 ;
        RECT 169.820 338.050 170.210 338.100 ;
        RECT 169.470 337.990 170.210 338.050 ;
        RECT 169.470 337.930 170.290 337.990 ;
        RECT 146.340 337.890 146.770 337.910 ;
        RECT 169.480 337.880 170.290 337.930 ;
        RECT 143.510 337.570 143.910 337.880 ;
        RECT 169.820 337.820 170.290 337.880 ;
        RECT 170.760 337.840 171.720 338.010 ;
        RECT 169.820 337.810 170.200 337.820 ;
        RECT 166.430 337.720 166.600 337.770 ;
        RECT 143.700 337.450 143.910 337.570 ;
        RECT 146.350 337.540 146.780 337.560 ;
        RECT 143.720 337.430 143.890 337.450 ;
        RECT 144.170 335.950 144.340 337.420 ;
        RECT 144.170 335.920 144.500 335.950 ;
        RECT 144.720 335.940 144.890 337.430 ;
        RECT 141.970 335.720 142.480 335.900 ;
        RECT 141.910 335.690 142.480 335.720 ;
        RECT 141.900 335.500 142.480 335.690 ;
        RECT 141.910 335.460 142.480 335.500 ;
        RECT 138.600 335.250 138.920 335.280 ;
        RECT 139.700 335.260 140.020 335.290 ;
        RECT 140.790 335.260 141.110 335.290 ;
        RECT 138.590 335.190 138.920 335.250 ;
        RECT 139.690 335.190 140.020 335.260 ;
        RECT 137.160 332.790 137.330 335.190 ;
        RECT 137.710 332.790 137.880 335.190 ;
        RECT 138.260 332.790 138.430 335.190 ;
        RECT 138.590 335.060 138.980 335.190 ;
        RECT 138.600 335.020 138.980 335.060 ;
        RECT 138.810 332.720 138.980 335.020 ;
        RECT 139.360 334.610 139.530 335.190 ;
        RECT 139.690 335.070 140.080 335.190 ;
        RECT 140.780 335.070 141.110 335.260 ;
        RECT 141.970 335.250 142.480 335.460 ;
        RECT 141.920 335.220 142.480 335.250 ;
        RECT 144.170 335.730 144.510 335.920 ;
        RECT 144.720 335.910 145.190 335.940 ;
        RECT 144.170 335.690 144.500 335.730 ;
        RECT 144.720 335.720 145.200 335.910 ;
        RECT 139.700 335.030 140.080 335.070 ;
        RECT 140.790 335.030 141.110 335.070 ;
        RECT 141.910 335.030 142.490 335.220 ;
        RECT 139.150 334.580 139.530 334.610 ;
        RECT 139.140 334.390 139.530 334.580 ;
        RECT 139.150 334.350 139.530 334.390 ;
        RECT 139.360 333.240 139.530 334.350 ;
        RECT 139.150 333.210 139.530 333.240 ;
        RECT 139.140 333.020 139.530 333.210 ;
        RECT 139.150 332.980 139.530 333.020 ;
        RECT 139.360 332.720 139.530 332.980 ;
        RECT 139.910 332.720 140.080 335.030 ;
        RECT 141.920 334.990 142.490 335.030 ;
        RECT 141.980 334.890 142.490 334.990 ;
        RECT 144.170 334.930 144.340 335.690 ;
        RECT 144.720 335.680 145.190 335.720 ;
        RECT 144.720 334.930 144.890 335.680 ;
        RECT 145.350 335.170 145.520 337.420 ;
        RECT 145.350 335.140 145.670 335.170 ;
        RECT 145.350 334.950 145.680 335.140 ;
        RECT 145.900 335.110 146.070 337.430 ;
        RECT 146.350 337.370 146.800 337.540 ;
        RECT 166.400 337.500 166.620 337.720 ;
        RECT 170.030 337.580 170.200 337.810 ;
        RECT 166.430 337.440 166.600 337.500 ;
        RECT 146.350 337.350 146.780 337.370 ;
        RECT 166.950 337.360 167.280 337.540 ;
        RECT 170.030 337.530 170.260 337.580 ;
        RECT 167.530 337.360 169.690 337.530 ;
        RECT 169.930 337.360 170.260 337.530 ;
        RECT 170.550 337.390 170.760 337.720 ;
        RECT 171.000 337.370 171.180 337.660 ;
        RECT 171.540 337.380 171.720 337.840 ;
        RECT 172.760 337.580 172.930 338.000 ;
        RECT 173.570 337.880 173.810 337.910 ;
        RECT 173.240 337.710 173.810 337.880 ;
        RECT 174.050 337.710 175.390 337.880 ;
        RECT 175.840 337.710 176.800 337.880 ;
        RECT 173.570 337.670 173.810 337.710 ;
        RECT 176.350 337.700 176.520 337.710 ;
        RECT 171.730 337.390 172.350 337.560 ;
        RECT 166.980 336.920 167.250 337.360 ;
        RECT 168.460 337.100 168.790 337.360 ;
        RECT 169.410 337.320 169.700 337.360 ;
        RECT 169.370 337.150 169.700 337.320 ;
        RECT 169.410 337.120 169.700 337.150 ;
        RECT 170.000 337.220 170.260 337.360 ;
        RECT 170.400 337.220 171.180 337.370 ;
        RECT 167.020 336.910 167.250 336.920 ;
        RECT 170.000 337.050 171.180 337.220 ;
        RECT 171.460 337.210 171.790 337.380 ;
        RECT 172.690 337.360 172.860 337.400 ;
        RECT 172.630 337.190 172.860 337.360 ;
        RECT 175.980 337.260 176.320 337.440 ;
        RECT 170.000 336.910 170.260 337.050 ;
        RECT 146.440 336.160 146.610 336.830 ;
        RECT 167.020 336.740 167.780 336.910 ;
        RECT 168.030 336.740 169.200 336.910 ;
        RECT 169.440 336.880 170.260 336.910 ;
        RECT 169.440 336.740 170.550 336.880 ;
        RECT 168.430 336.640 168.780 336.740 ;
        RECT 170.090 336.710 170.550 336.740 ;
        RECT 171.000 336.710 172.190 336.880 ;
        RECT 172.690 336.840 172.860 337.190 ;
        RECT 172.930 336.970 173.120 337.200 ;
        RECT 173.220 337.090 173.590 337.260 ;
        RECT 174.050 337.090 176.800 337.260 ;
        RECT 177.330 337.020 177.500 337.950 ;
        RECT 177.730 337.110 177.900 338.000 ;
        RECT 208.340 337.720 208.680 338.120 ;
        RECT 208.850 337.950 209.180 338.120 ;
        RECT 209.400 337.950 209.740 338.120 ;
        RECT 208.930 337.780 209.100 337.950 ;
        RECT 209.490 337.780 209.660 337.950 ;
        RECT 208.160 337.610 208.680 337.720 ;
        RECT 208.850 337.610 209.180 337.780 ;
        RECT 209.400 337.610 209.740 337.780 ;
        RECT 208.160 337.500 208.490 337.610 ;
        RECT 208.160 337.460 208.480 337.500 ;
        RECT 208.930 337.380 209.180 337.610 ;
        RECT 210.060 337.530 210.570 338.200 ;
        RECT 208.930 337.210 209.600 337.380 ;
        RECT 208.160 337.090 208.480 337.130 ;
        RECT 196.570 337.030 196.890 337.070 ;
        RECT 196.570 336.860 196.900 337.030 ;
        RECT 208.160 336.980 208.490 337.090 ;
        RECT 208.930 336.980 209.180 337.210 ;
        RECT 208.160 336.870 208.680 336.980 ;
        RECT 196.480 336.840 196.900 336.860 ;
        RECT 171.040 336.690 172.190 336.710 ;
        RECT 172.020 336.650 172.190 336.690 ;
        RECT 196.480 336.810 196.890 336.840 ;
        RECT 169.820 336.300 170.210 336.350 ;
        RECT 169.470 336.240 170.210 336.300 ;
        RECT 169.470 336.180 170.290 336.240 ;
        RECT 169.480 336.130 170.290 336.180 ;
        RECT 169.820 336.070 170.290 336.130 ;
        RECT 170.760 336.090 171.720 336.260 ;
        RECT 169.820 336.060 170.200 336.070 ;
        RECT 166.430 335.970 166.600 336.020 ;
        RECT 166.400 335.750 166.620 335.970 ;
        RECT 170.030 335.830 170.200 336.060 ;
        RECT 166.430 335.690 166.600 335.750 ;
        RECT 166.950 335.610 167.280 335.790 ;
        RECT 170.030 335.780 170.260 335.830 ;
        RECT 167.530 335.610 169.690 335.780 ;
        RECT 169.930 335.610 170.260 335.780 ;
        RECT 170.550 335.640 170.760 335.970 ;
        RECT 171.000 335.620 171.180 335.910 ;
        RECT 171.540 335.630 171.720 336.090 ;
        RECT 172.690 336.080 172.860 336.430 ;
        RECT 172.630 335.910 172.860 336.080 ;
        RECT 172.930 336.070 173.120 336.300 ;
        RECT 173.220 336.010 173.590 336.180 ;
        RECT 174.050 336.010 176.800 336.180 ;
        RECT 172.690 335.870 172.860 335.910 ;
        RECT 175.980 335.830 176.320 336.010 ;
        RECT 171.730 335.640 172.350 335.810 ;
        RECT 166.980 335.170 167.250 335.610 ;
        RECT 168.460 335.350 168.790 335.610 ;
        RECT 169.410 335.570 169.700 335.610 ;
        RECT 169.370 335.400 169.700 335.570 ;
        RECT 169.410 335.370 169.700 335.400 ;
        RECT 170.000 335.470 170.260 335.610 ;
        RECT 170.400 335.470 171.180 335.620 ;
        RECT 167.020 335.160 167.250 335.170 ;
        RECT 170.000 335.300 171.180 335.470 ;
        RECT 171.460 335.460 171.790 335.630 ;
        RECT 170.000 335.160 170.260 335.300 ;
        RECT 172.760 335.270 172.930 335.690 ;
        RECT 173.570 335.560 173.810 335.600 ;
        RECT 176.350 335.560 176.520 335.570 ;
        RECT 173.240 335.390 173.810 335.560 ;
        RECT 174.050 335.390 175.390 335.560 ;
        RECT 175.840 335.390 176.800 335.560 ;
        RECT 173.570 335.360 173.810 335.390 ;
        RECT 177.330 335.320 177.500 336.250 ;
        RECT 177.730 335.270 177.900 336.160 ;
        RECT 196.480 336.110 196.660 336.810 ;
        RECT 208.340 336.470 208.680 336.870 ;
        RECT 208.850 336.810 209.180 336.980 ;
        RECT 209.400 336.810 209.740 336.980 ;
        RECT 208.930 336.640 209.100 336.810 ;
        RECT 209.490 336.640 209.660 336.810 ;
        RECT 208.850 336.470 209.180 336.640 ;
        RECT 209.400 336.470 209.740 336.640 ;
        RECT 208.010 336.410 208.330 336.450 ;
        RECT 208.010 336.240 208.340 336.410 ;
        RECT 209.490 336.240 209.660 336.470 ;
        RECT 210.060 336.390 210.570 337.060 ;
        RECT 208.010 336.190 209.660 336.240 ;
        RECT 196.480 336.070 196.940 336.110 ;
        RECT 208.200 336.070 209.660 336.190 ;
        RECT 196.480 335.940 196.950 336.070 ;
        RECT 196.620 335.880 196.950 335.940 ;
        RECT 196.620 335.850 196.940 335.880 ;
        RECT 145.900 335.080 146.380 335.110 ;
        RECT 145.350 334.910 145.670 334.950 ;
        RECT 145.900 334.930 146.390 335.080 ;
        RECT 167.020 334.990 167.780 335.160 ;
        RECT 168.030 334.990 169.200 335.160 ;
        RECT 169.440 335.130 170.260 335.160 ;
        RECT 169.440 334.990 170.550 335.130 ;
        RECT 146.060 334.890 146.390 334.930 ;
        RECT 168.430 334.890 168.780 334.990 ;
        RECT 170.090 334.960 170.550 334.990 ;
        RECT 171.000 334.960 172.190 335.130 ;
        RECT 171.040 334.940 172.190 334.960 ;
        RECT 172.020 334.900 172.190 334.940 ;
        RECT 146.060 334.850 146.380 334.890 ;
        RECT 140.250 334.580 140.570 334.610 ;
        RECT 141.350 334.580 141.670 334.610 ;
        RECT 140.240 334.390 140.570 334.580 ;
        RECT 141.340 334.390 141.670 334.580 ;
        RECT 140.250 334.350 140.570 334.390 ;
        RECT 141.350 334.350 141.670 334.390 ;
        RECT 142.270 333.480 142.440 334.700 ;
        RECT 172.500 333.460 172.820 333.500 ;
        RECT 173.590 333.460 173.910 333.500 ;
        RECT 172.500 333.440 172.830 333.460 ;
        RECT 173.590 333.440 173.920 333.460 ;
        RECT 174.690 333.450 175.010 333.490 ;
        RECT 174.690 333.440 175.020 333.450 ;
        RECT 172.440 333.270 172.830 333.440 ;
        RECT 172.440 333.240 172.820 333.270 ;
        RECT 140.250 333.210 140.570 333.240 ;
        RECT 141.350 333.210 141.670 333.240 ;
        RECT 140.240 333.100 140.570 333.210 ;
        RECT 141.340 333.100 141.670 333.210 ;
        RECT 140.240 333.020 140.630 333.100 ;
        RECT 140.250 332.980 140.630 333.020 ;
        RECT 140.460 332.720 140.630 332.980 ;
        RECT 141.010 332.720 141.180 333.100 ;
        RECT 141.340 333.020 141.730 333.100 ;
        RECT 141.350 332.980 141.730 333.020 ;
        RECT 141.560 332.720 141.730 332.980 ;
        RECT 138.600 332.480 138.920 332.510 ;
        RECT 139.700 332.480 140.020 332.510 ;
        RECT 140.790 332.480 141.110 332.510 ;
        RECT 138.590 332.410 138.920 332.480 ;
        RECT 139.690 332.410 140.020 332.480 ;
        RECT 4.240 330.710 11.770 331.220 ;
        RECT 2.540 324.690 4.000 324.730 ;
        RECT 2.540 324.520 4.010 324.690 ;
        RECT 2.540 324.480 4.000 324.520 ;
        RECT 4.240 318.100 4.750 330.710 ;
        RECT 5.110 329.920 11.090 330.150 ;
        RECT 5.200 318.860 10.850 329.920 ;
        RECT 11.260 320.350 11.770 330.710 ;
        RECT 137.160 330.010 137.330 332.410 ;
        RECT 137.710 330.010 137.880 332.410 ;
        RECT 138.260 330.010 138.430 332.410 ;
        RECT 138.590 332.290 138.980 332.410 ;
        RECT 138.600 332.250 138.980 332.290 ;
        RECT 138.810 331.170 138.980 332.250 ;
        RECT 138.590 331.140 138.980 331.170 ;
        RECT 138.580 330.950 138.980 331.140 ;
        RECT 138.590 330.910 138.980 330.950 ;
        RECT 138.810 330.010 138.980 330.910 ;
        RECT 139.360 330.470 139.530 332.410 ;
        RECT 139.690 332.290 140.080 332.410 ;
        RECT 140.780 332.290 141.110 332.480 ;
        RECT 139.700 332.250 140.080 332.290 ;
        RECT 140.790 332.250 141.110 332.290 ;
        RECT 139.910 331.160 140.080 332.250 ;
        RECT 148.600 331.200 149.360 331.620 ;
        RECT 139.700 331.130 140.080 331.160 ;
        RECT 139.690 330.940 140.080 331.130 ;
        RECT 140.790 331.110 141.110 331.140 ;
        RECT 139.700 330.900 140.080 330.940 ;
        RECT 140.780 330.920 141.110 331.110 ;
        RECT 139.150 330.440 139.530 330.470 ;
        RECT 139.140 330.250 139.530 330.440 ;
        RECT 139.150 330.210 139.530 330.250 ;
        RECT 139.360 330.010 139.530 330.210 ;
        RECT 139.910 330.010 140.080 330.900 ;
        RECT 140.790 330.880 141.110 330.920 ;
        RECT 140.250 330.430 140.570 330.460 ;
        RECT 141.340 330.430 141.660 330.460 ;
        RECT 140.240 330.240 140.570 330.430 ;
        RECT 141.330 330.240 141.660 330.430 ;
        RECT 148.620 330.410 149.360 331.200 ;
        RECT 172.440 330.720 172.610 333.240 ;
        RECT 172.990 332.820 173.160 333.440 ;
        RECT 173.540 333.270 173.920 333.440 ;
        RECT 173.540 333.240 173.910 333.270 ;
        RECT 172.990 332.780 173.370 332.820 ;
        RECT 172.990 332.590 173.380 332.780 ;
        RECT 172.990 332.560 173.370 332.590 ;
        RECT 172.990 331.450 173.160 332.560 ;
        RECT 172.990 331.410 173.370 331.450 ;
        RECT 172.990 331.220 173.380 331.410 ;
        RECT 172.990 331.190 173.370 331.220 ;
        RECT 172.440 330.680 172.810 330.720 ;
        RECT 172.440 330.490 172.820 330.680 ;
        RECT 172.440 330.460 172.810 330.490 ;
        RECT 140.250 330.200 140.570 330.240 ;
        RECT 141.340 330.200 141.660 330.240 ;
        RECT 172.440 329.350 172.610 330.460 ;
        RECT 172.440 329.310 172.810 329.350 ;
        RECT 172.440 329.120 172.820 329.310 ;
        RECT 172.440 329.090 172.810 329.120 ;
        RECT 171.670 328.730 172.180 328.810 ;
        RECT 171.670 328.710 172.190 328.730 ;
        RECT 171.670 328.670 172.240 328.710 ;
        RECT 171.670 328.480 172.250 328.670 ;
        RECT 171.680 328.450 172.240 328.480 ;
        RECT 171.680 328.240 172.190 328.450 ;
        RECT 171.680 328.200 172.250 328.240 ;
        RECT 171.680 328.010 172.260 328.200 ;
        RECT 172.440 328.120 172.610 329.090 ;
        RECT 172.990 328.670 173.160 331.190 ;
        RECT 173.540 330.720 173.710 333.240 ;
        RECT 174.090 332.800 174.260 333.440 ;
        RECT 174.640 333.260 175.020 333.440 ;
        RECT 174.640 333.230 175.010 333.260 ;
        RECT 174.090 332.760 174.460 332.800 ;
        RECT 174.090 332.570 174.470 332.760 ;
        RECT 174.090 332.540 174.460 332.570 ;
        RECT 174.090 331.450 174.260 332.540 ;
        RECT 174.090 331.410 174.460 331.450 ;
        RECT 174.090 331.220 174.470 331.410 ;
        RECT 174.090 331.190 174.460 331.220 ;
        RECT 173.540 330.680 173.910 330.720 ;
        RECT 173.540 330.490 173.920 330.680 ;
        RECT 173.540 330.460 173.910 330.490 ;
        RECT 173.540 329.350 173.710 330.460 ;
        RECT 173.540 329.310 173.910 329.350 ;
        RECT 173.540 329.120 173.920 329.310 ;
        RECT 173.540 329.090 173.910 329.120 ;
        RECT 172.990 328.630 173.370 328.670 ;
        RECT 172.990 328.440 173.380 328.630 ;
        RECT 172.990 328.410 173.370 328.440 ;
        RECT 172.990 328.110 173.160 328.410 ;
        RECT 173.540 328.110 173.710 329.090 ;
        RECT 174.090 328.670 174.260 331.190 ;
        RECT 174.640 330.720 174.810 333.230 ;
        RECT 175.190 332.790 175.360 333.440 ;
        RECT 175.190 332.750 175.570 332.790 ;
        RECT 175.190 332.560 175.580 332.750 ;
        RECT 175.730 332.710 175.900 333.470 ;
        RECT 176.340 332.710 176.510 333.470 ;
        RECT 177.230 333.450 177.550 333.490 ;
        RECT 178.330 333.460 178.650 333.500 ;
        RECT 179.420 333.460 179.740 333.500 ;
        RECT 182.310 333.490 182.630 333.530 ;
        RECT 183.400 333.490 183.720 333.530 ;
        RECT 182.310 333.470 182.640 333.490 ;
        RECT 183.400 333.470 183.730 333.490 ;
        RECT 184.500 333.480 184.820 333.520 ;
        RECT 184.500 333.470 184.830 333.480 ;
        RECT 177.220 333.440 177.550 333.450 ;
        RECT 178.320 333.440 178.650 333.460 ;
        RECT 179.410 333.440 179.740 333.460 ;
        RECT 176.880 332.790 177.050 333.440 ;
        RECT 177.220 333.260 177.600 333.440 ;
        RECT 177.230 333.230 177.600 333.260 ;
        RECT 176.670 332.750 177.050 332.790 ;
        RECT 176.660 332.560 177.050 332.750 ;
        RECT 175.190 332.530 175.570 332.560 ;
        RECT 176.670 332.530 177.050 332.560 ;
        RECT 175.190 331.450 175.360 332.530 ;
        RECT 176.880 331.450 177.050 332.530 ;
        RECT 175.190 331.410 175.560 331.450 ;
        RECT 176.680 331.410 177.050 331.450 ;
        RECT 175.190 331.220 175.570 331.410 ;
        RECT 176.670 331.220 177.050 331.410 ;
        RECT 175.190 331.190 175.560 331.220 ;
        RECT 176.680 331.190 177.050 331.220 ;
        RECT 174.640 330.680 175.010 330.720 ;
        RECT 174.640 330.490 175.020 330.680 ;
        RECT 174.640 330.460 175.010 330.490 ;
        RECT 174.640 329.350 174.810 330.460 ;
        RECT 174.640 329.310 175.010 329.350 ;
        RECT 174.640 329.120 175.020 329.310 ;
        RECT 174.640 329.090 175.010 329.120 ;
        RECT 174.090 328.630 174.460 328.670 ;
        RECT 174.090 328.440 174.470 328.630 ;
        RECT 174.090 328.410 174.460 328.440 ;
        RECT 174.090 328.110 174.260 328.410 ;
        RECT 174.640 328.110 174.810 329.090 ;
        RECT 175.190 328.680 175.360 331.190 ;
        RECT 176.880 328.680 177.050 331.190 ;
        RECT 177.430 330.720 177.600 333.230 ;
        RECT 177.980 332.800 178.150 333.440 ;
        RECT 178.320 333.270 178.700 333.440 ;
        RECT 178.330 333.240 178.700 333.270 ;
        RECT 177.780 332.760 178.150 332.800 ;
        RECT 177.770 332.570 178.150 332.760 ;
        RECT 177.780 332.540 178.150 332.570 ;
        RECT 177.980 331.450 178.150 332.540 ;
        RECT 177.780 331.410 178.150 331.450 ;
        RECT 177.770 331.220 178.150 331.410 ;
        RECT 177.780 331.190 178.150 331.220 ;
        RECT 177.230 330.680 177.600 330.720 ;
        RECT 177.220 330.490 177.600 330.680 ;
        RECT 177.230 330.460 177.600 330.490 ;
        RECT 177.430 329.350 177.600 330.460 ;
        RECT 177.230 329.310 177.600 329.350 ;
        RECT 177.220 329.120 177.600 329.310 ;
        RECT 177.230 329.090 177.600 329.120 ;
        RECT 175.190 328.640 175.560 328.680 ;
        RECT 176.680 328.640 177.050 328.680 ;
        RECT 175.190 328.450 175.570 328.640 ;
        RECT 176.670 328.450 177.050 328.640 ;
        RECT 175.190 328.420 175.560 328.450 ;
        RECT 176.680 328.420 177.050 328.450 ;
        RECT 175.190 328.110 175.360 328.420 ;
        RECT 176.880 328.110 177.050 328.420 ;
        RECT 177.430 328.110 177.600 329.090 ;
        RECT 177.980 328.670 178.150 331.190 ;
        RECT 178.530 330.720 178.700 333.240 ;
        RECT 179.080 332.820 179.250 333.440 ;
        RECT 179.410 333.270 179.800 333.440 ;
        RECT 179.420 333.240 179.800 333.270 ;
        RECT 178.870 332.780 179.250 332.820 ;
        RECT 178.860 332.590 179.250 332.780 ;
        RECT 178.870 332.560 179.250 332.590 ;
        RECT 179.080 331.450 179.250 332.560 ;
        RECT 178.870 331.410 179.250 331.450 ;
        RECT 178.860 331.220 179.250 331.410 ;
        RECT 178.870 331.190 179.250 331.220 ;
        RECT 178.330 330.680 178.700 330.720 ;
        RECT 178.320 330.490 178.700 330.680 ;
        RECT 178.330 330.460 178.700 330.490 ;
        RECT 178.530 329.350 178.700 330.460 ;
        RECT 178.330 329.310 178.700 329.350 ;
        RECT 178.320 329.120 178.700 329.310 ;
        RECT 178.330 329.090 178.700 329.120 ;
        RECT 177.780 328.630 178.150 328.670 ;
        RECT 177.770 328.440 178.150 328.630 ;
        RECT 177.780 328.410 178.150 328.440 ;
        RECT 177.980 328.110 178.150 328.410 ;
        RECT 178.530 328.110 178.700 329.090 ;
        RECT 179.080 328.670 179.250 331.190 ;
        RECT 179.630 330.720 179.800 333.240 ;
        RECT 179.430 330.680 179.800 330.720 ;
        RECT 179.420 330.490 179.800 330.680 ;
        RECT 179.430 330.460 179.800 330.490 ;
        RECT 179.630 329.350 179.800 330.460 ;
        RECT 179.430 329.310 179.800 329.350 ;
        RECT 179.420 329.120 179.800 329.310 ;
        RECT 179.430 329.090 179.800 329.120 ;
        RECT 178.870 328.630 179.250 328.670 ;
        RECT 178.860 328.440 179.250 328.630 ;
        RECT 178.870 328.410 179.250 328.440 ;
        RECT 179.080 328.110 179.250 328.410 ;
        RECT 179.630 328.120 179.800 329.090 ;
        RECT 182.250 333.300 182.640 333.470 ;
        RECT 182.250 333.270 182.630 333.300 ;
        RECT 182.250 330.750 182.420 333.270 ;
        RECT 182.800 332.850 182.970 333.470 ;
        RECT 183.350 333.300 183.730 333.470 ;
        RECT 183.350 333.270 183.720 333.300 ;
        RECT 182.800 332.810 183.180 332.850 ;
        RECT 182.800 332.620 183.190 332.810 ;
        RECT 182.800 332.590 183.180 332.620 ;
        RECT 182.800 331.480 182.970 332.590 ;
        RECT 182.800 331.440 183.180 331.480 ;
        RECT 182.800 331.250 183.190 331.440 ;
        RECT 182.800 331.220 183.180 331.250 ;
        RECT 182.250 330.710 182.620 330.750 ;
        RECT 182.250 330.520 182.630 330.710 ;
        RECT 182.250 330.490 182.620 330.520 ;
        RECT 182.250 329.380 182.420 330.490 ;
        RECT 182.250 329.340 182.620 329.380 ;
        RECT 182.250 329.150 182.630 329.340 ;
        RECT 182.250 329.120 182.620 329.150 ;
        RECT 180.060 328.730 180.570 328.810 ;
        RECT 180.050 328.710 180.570 328.730 ;
        RECT 180.000 328.670 180.570 328.710 ;
        RECT 179.990 328.480 180.570 328.670 ;
        RECT 181.480 328.760 181.990 328.840 ;
        RECT 181.480 328.740 182.000 328.760 ;
        RECT 181.480 328.700 182.050 328.740 ;
        RECT 181.480 328.510 182.060 328.700 ;
        RECT 181.490 328.480 182.050 328.510 ;
        RECT 180.000 328.450 180.560 328.480 ;
        RECT 180.050 328.240 180.560 328.450 ;
        RECT 179.990 328.200 180.560 328.240 ;
        RECT 179.980 328.010 180.560 328.200 ;
        RECT 171.680 327.980 172.250 328.010 ;
        RECT 179.990 327.980 180.560 328.010 ;
        RECT 171.680 327.800 172.190 327.980 ;
        RECT 180.050 327.800 180.560 327.980 ;
        RECT 181.490 328.270 182.000 328.480 ;
        RECT 181.490 328.230 182.060 328.270 ;
        RECT 181.490 328.040 182.070 328.230 ;
        RECT 182.250 328.150 182.420 329.120 ;
        RECT 182.800 328.700 182.970 331.220 ;
        RECT 183.350 330.750 183.520 333.270 ;
        RECT 183.900 332.830 184.070 333.470 ;
        RECT 184.450 333.290 184.830 333.470 ;
        RECT 184.450 333.260 184.820 333.290 ;
        RECT 183.900 332.790 184.270 332.830 ;
        RECT 183.900 332.600 184.280 332.790 ;
        RECT 183.900 332.570 184.270 332.600 ;
        RECT 183.900 331.480 184.070 332.570 ;
        RECT 183.900 331.440 184.270 331.480 ;
        RECT 183.900 331.250 184.280 331.440 ;
        RECT 183.900 331.220 184.270 331.250 ;
        RECT 183.350 330.710 183.720 330.750 ;
        RECT 183.350 330.520 183.730 330.710 ;
        RECT 183.350 330.490 183.720 330.520 ;
        RECT 183.350 329.380 183.520 330.490 ;
        RECT 183.350 329.340 183.720 329.380 ;
        RECT 183.350 329.150 183.730 329.340 ;
        RECT 183.350 329.120 183.720 329.150 ;
        RECT 182.800 328.660 183.180 328.700 ;
        RECT 182.800 328.470 183.190 328.660 ;
        RECT 182.800 328.440 183.180 328.470 ;
        RECT 182.800 328.140 182.970 328.440 ;
        RECT 183.350 328.140 183.520 329.120 ;
        RECT 183.900 328.700 184.070 331.220 ;
        RECT 184.450 330.750 184.620 333.260 ;
        RECT 185.000 332.820 185.170 333.470 ;
        RECT 185.000 332.780 185.380 332.820 ;
        RECT 185.000 332.590 185.390 332.780 ;
        RECT 185.540 332.740 185.710 333.500 ;
        RECT 186.150 332.740 186.320 333.500 ;
        RECT 187.040 333.480 187.360 333.520 ;
        RECT 188.140 333.490 188.460 333.530 ;
        RECT 189.230 333.490 189.550 333.530 ;
        RECT 187.030 333.470 187.360 333.480 ;
        RECT 188.130 333.470 188.460 333.490 ;
        RECT 189.220 333.470 189.550 333.490 ;
        RECT 186.690 332.820 186.860 333.470 ;
        RECT 187.030 333.290 187.410 333.470 ;
        RECT 187.040 333.260 187.410 333.290 ;
        RECT 186.480 332.780 186.860 332.820 ;
        RECT 186.470 332.590 186.860 332.780 ;
        RECT 185.000 332.560 185.380 332.590 ;
        RECT 186.480 332.560 186.860 332.590 ;
        RECT 185.000 331.480 185.170 332.560 ;
        RECT 186.690 331.480 186.860 332.560 ;
        RECT 185.000 331.440 185.370 331.480 ;
        RECT 186.490 331.440 186.860 331.480 ;
        RECT 185.000 331.250 185.380 331.440 ;
        RECT 186.480 331.250 186.860 331.440 ;
        RECT 185.000 331.220 185.370 331.250 ;
        RECT 186.490 331.220 186.860 331.250 ;
        RECT 184.450 330.710 184.820 330.750 ;
        RECT 184.450 330.520 184.830 330.710 ;
        RECT 184.450 330.490 184.820 330.520 ;
        RECT 184.450 329.380 184.620 330.490 ;
        RECT 184.450 329.340 184.820 329.380 ;
        RECT 184.450 329.150 184.830 329.340 ;
        RECT 184.450 329.120 184.820 329.150 ;
        RECT 183.900 328.660 184.270 328.700 ;
        RECT 183.900 328.470 184.280 328.660 ;
        RECT 183.900 328.440 184.270 328.470 ;
        RECT 183.900 328.140 184.070 328.440 ;
        RECT 184.450 328.140 184.620 329.120 ;
        RECT 185.000 328.710 185.170 331.220 ;
        RECT 186.690 328.710 186.860 331.220 ;
        RECT 187.240 330.750 187.410 333.260 ;
        RECT 187.790 332.830 187.960 333.470 ;
        RECT 188.130 333.300 188.510 333.470 ;
        RECT 188.140 333.270 188.510 333.300 ;
        RECT 187.590 332.790 187.960 332.830 ;
        RECT 187.580 332.600 187.960 332.790 ;
        RECT 187.590 332.570 187.960 332.600 ;
        RECT 187.790 331.480 187.960 332.570 ;
        RECT 187.590 331.440 187.960 331.480 ;
        RECT 187.580 331.250 187.960 331.440 ;
        RECT 187.590 331.220 187.960 331.250 ;
        RECT 187.040 330.710 187.410 330.750 ;
        RECT 187.030 330.520 187.410 330.710 ;
        RECT 187.040 330.490 187.410 330.520 ;
        RECT 187.240 329.380 187.410 330.490 ;
        RECT 187.040 329.340 187.410 329.380 ;
        RECT 187.030 329.150 187.410 329.340 ;
        RECT 187.040 329.120 187.410 329.150 ;
        RECT 185.000 328.670 185.370 328.710 ;
        RECT 186.490 328.670 186.860 328.710 ;
        RECT 185.000 328.480 185.380 328.670 ;
        RECT 186.480 328.480 186.860 328.670 ;
        RECT 185.000 328.450 185.370 328.480 ;
        RECT 186.490 328.450 186.860 328.480 ;
        RECT 185.000 328.140 185.170 328.450 ;
        RECT 186.690 328.140 186.860 328.450 ;
        RECT 187.240 328.140 187.410 329.120 ;
        RECT 187.790 328.700 187.960 331.220 ;
        RECT 188.340 330.750 188.510 333.270 ;
        RECT 188.890 332.850 189.060 333.470 ;
        RECT 189.220 333.300 189.610 333.470 ;
        RECT 189.230 333.270 189.610 333.300 ;
        RECT 188.680 332.810 189.060 332.850 ;
        RECT 188.670 332.620 189.060 332.810 ;
        RECT 188.680 332.590 189.060 332.620 ;
        RECT 188.890 331.480 189.060 332.590 ;
        RECT 188.680 331.440 189.060 331.480 ;
        RECT 188.670 331.250 189.060 331.440 ;
        RECT 188.680 331.220 189.060 331.250 ;
        RECT 188.140 330.710 188.510 330.750 ;
        RECT 188.130 330.520 188.510 330.710 ;
        RECT 188.140 330.490 188.510 330.520 ;
        RECT 188.340 329.380 188.510 330.490 ;
        RECT 188.140 329.340 188.510 329.380 ;
        RECT 188.130 329.150 188.510 329.340 ;
        RECT 188.140 329.120 188.510 329.150 ;
        RECT 187.590 328.660 187.960 328.700 ;
        RECT 187.580 328.470 187.960 328.660 ;
        RECT 187.590 328.440 187.960 328.470 ;
        RECT 187.790 328.140 187.960 328.440 ;
        RECT 188.340 328.140 188.510 329.120 ;
        RECT 188.890 328.700 189.060 331.220 ;
        RECT 189.440 330.750 189.610 333.270 ;
        RECT 189.240 330.710 189.610 330.750 ;
        RECT 189.230 330.520 189.610 330.710 ;
        RECT 189.240 330.490 189.610 330.520 ;
        RECT 189.440 329.380 189.610 330.490 ;
        RECT 189.240 329.340 189.610 329.380 ;
        RECT 189.230 329.150 189.610 329.340 ;
        RECT 189.240 329.120 189.610 329.150 ;
        RECT 188.680 328.660 189.060 328.700 ;
        RECT 188.670 328.470 189.060 328.660 ;
        RECT 188.680 328.440 189.060 328.470 ;
        RECT 188.890 328.140 189.060 328.440 ;
        RECT 189.440 328.150 189.610 329.120 ;
        RECT 189.870 328.760 190.380 328.840 ;
        RECT 189.860 328.740 190.380 328.760 ;
        RECT 189.810 328.700 190.380 328.740 ;
        RECT 189.800 328.510 190.380 328.700 ;
        RECT 189.810 328.480 190.370 328.510 ;
        RECT 189.860 328.270 190.370 328.480 ;
        RECT 189.800 328.230 190.370 328.270 ;
        RECT 189.790 328.040 190.370 328.230 ;
        RECT 181.490 328.010 182.060 328.040 ;
        RECT 189.800 328.010 190.370 328.040 ;
        RECT 181.490 327.830 182.000 328.010 ;
        RECT 189.860 327.830 190.370 328.010 ;
        RECT 191.430 327.110 191.600 329.510 ;
        RECT 191.980 327.110 192.150 329.510 ;
        RECT 192.530 327.110 192.700 329.510 ;
        RECT 193.080 328.610 193.250 329.510 ;
        RECT 193.630 329.310 193.800 329.510 ;
        RECT 193.420 329.270 193.800 329.310 ;
        RECT 193.410 329.080 193.800 329.270 ;
        RECT 193.420 329.050 193.800 329.080 ;
        RECT 192.860 328.570 193.250 328.610 ;
        RECT 192.850 328.380 193.250 328.570 ;
        RECT 192.860 328.350 193.250 328.380 ;
        RECT 193.080 327.270 193.250 328.350 ;
        RECT 192.870 327.230 193.250 327.270 ;
        RECT 192.860 327.110 193.250 327.230 ;
        RECT 193.630 327.110 193.800 329.050 ;
        RECT 194.180 328.620 194.350 329.510 ;
        RECT 194.520 329.280 194.840 329.320 ;
        RECT 195.610 329.280 195.930 329.320 ;
        RECT 194.510 329.090 194.840 329.280 ;
        RECT 195.600 329.090 195.930 329.280 ;
        RECT 194.520 329.060 194.840 329.090 ;
        RECT 195.610 329.060 195.930 329.090 ;
        RECT 193.970 328.580 194.350 328.620 ;
        RECT 195.060 328.600 195.380 328.640 ;
        RECT 193.960 328.390 194.350 328.580 ;
        RECT 195.050 328.410 195.380 328.600 ;
        RECT 193.970 328.360 194.350 328.390 ;
        RECT 195.060 328.380 195.380 328.410 ;
        RECT 194.180 327.270 194.350 328.360 ;
        RECT 193.970 327.230 194.350 327.270 ;
        RECT 195.060 327.230 195.380 327.270 ;
        RECT 193.960 327.110 194.350 327.230 ;
        RECT 192.860 327.040 193.190 327.110 ;
        RECT 193.960 327.040 194.290 327.110 ;
        RECT 195.050 327.040 195.380 327.230 ;
        RECT 192.870 327.010 193.190 327.040 ;
        RECT 193.970 327.010 194.290 327.040 ;
        RECT 195.060 327.010 195.380 327.040 ;
        RECT 191.430 324.330 191.600 326.730 ;
        RECT 191.980 324.330 192.150 326.730 ;
        RECT 192.530 324.330 192.700 326.730 ;
        RECT 193.080 324.500 193.250 326.800 ;
        RECT 193.630 326.540 193.800 326.800 ;
        RECT 193.420 326.500 193.800 326.540 ;
        RECT 193.410 326.310 193.800 326.500 ;
        RECT 193.420 326.280 193.800 326.310 ;
        RECT 193.630 325.170 193.800 326.280 ;
        RECT 193.420 325.130 193.800 325.170 ;
        RECT 193.410 324.940 193.800 325.130 ;
        RECT 193.420 324.910 193.800 324.940 ;
        RECT 192.870 324.460 193.250 324.500 ;
        RECT 192.860 324.330 193.250 324.460 ;
        RECT 193.630 324.330 193.800 324.910 ;
        RECT 194.180 324.490 194.350 326.800 ;
        RECT 194.730 326.540 194.900 326.800 ;
        RECT 194.520 326.500 194.900 326.540 ;
        RECT 194.510 326.420 194.900 326.500 ;
        RECT 195.280 326.420 195.450 326.800 ;
        RECT 195.830 326.540 196.000 326.800 ;
        RECT 195.620 326.500 196.000 326.540 ;
        RECT 195.610 326.420 196.000 326.500 ;
        RECT 194.510 326.310 194.840 326.420 ;
        RECT 195.610 326.310 195.940 326.420 ;
        RECT 194.520 326.280 194.840 326.310 ;
        RECT 195.620 326.280 195.940 326.310 ;
        RECT 194.520 325.130 194.840 325.170 ;
        RECT 195.620 325.130 195.940 325.170 ;
        RECT 194.510 324.940 194.840 325.130 ;
        RECT 195.610 324.940 195.940 325.130 ;
        RECT 194.520 324.910 194.840 324.940 ;
        RECT 195.620 324.910 195.940 324.940 ;
        RECT 196.540 324.820 196.710 326.040 ;
        RECT 227.070 325.530 227.300 325.640 ;
        RECT 226.970 325.360 231.630 325.530 ;
        RECT 229.950 325.080 230.280 325.250 ;
        RECT 230.910 325.080 231.240 325.250 ;
        RECT 231.870 325.080 232.200 325.250 ;
        RECT 232.830 325.080 233.160 325.250 ;
        RECT 232.680 325.020 232.870 325.030 ;
        RECT 228.190 324.840 231.990 324.850 ;
        RECT 232.650 324.840 232.910 325.020 ;
        RECT 228.190 324.700 232.910 324.840 ;
        RECT 228.190 324.680 232.670 324.700 ;
        RECT 231.760 324.670 232.670 324.680 ;
        RECT 196.250 324.530 196.760 324.630 ;
        RECT 231.760 324.570 231.990 324.670 ;
        RECT 196.190 324.490 196.760 324.530 ;
        RECT 193.970 324.450 194.350 324.490 ;
        RECT 195.060 324.450 195.380 324.490 ;
        RECT 193.960 324.330 194.350 324.450 ;
        RECT 192.860 324.270 193.190 324.330 ;
        RECT 192.870 324.240 193.190 324.270 ;
        RECT 193.960 324.260 194.290 324.330 ;
        RECT 195.050 324.260 195.380 324.450 ;
        RECT 196.180 324.300 196.760 324.490 ;
        RECT 229.950 324.400 230.280 324.570 ;
        RECT 230.910 324.400 231.240 324.570 ;
        RECT 231.760 324.400 232.200 324.570 ;
        RECT 232.830 324.400 233.160 324.570 ;
        RECT 196.190 324.270 196.750 324.300 ;
        RECT 193.970 324.230 194.290 324.260 ;
        RECT 195.060 324.230 195.380 324.260 ;
        RECT 141.370 323.970 141.880 324.150 ;
        RECT 196.240 324.060 196.750 324.270 ;
        RECT 196.180 324.020 196.750 324.060 ;
        RECT 231.760 324.210 231.990 324.400 ;
        RECT 232.680 324.350 232.870 324.360 ;
        RECT 232.650 324.210 232.910 324.350 ;
        RECT 231.760 324.030 232.910 324.210 ;
        RECT 141.310 323.940 141.880 323.970 ;
        RECT 138.200 323.530 138.370 323.840 ;
        RECT 138.000 323.500 138.370 323.530 ;
        RECT 137.990 323.310 138.370 323.500 ;
        RECT 138.000 323.270 138.370 323.310 ;
        RECT 138.200 320.760 138.370 323.270 ;
        RECT 138.750 322.860 138.920 323.840 ;
        RECT 139.300 323.540 139.470 323.840 ;
        RECT 139.100 323.510 139.470 323.540 ;
        RECT 139.090 323.320 139.470 323.510 ;
        RECT 139.100 323.280 139.470 323.320 ;
        RECT 138.550 322.830 138.920 322.860 ;
        RECT 138.540 322.640 138.920 322.830 ;
        RECT 138.550 322.600 138.920 322.640 ;
        RECT 138.750 321.490 138.920 322.600 ;
        RECT 138.550 321.460 138.920 321.490 ;
        RECT 138.540 321.270 138.920 321.460 ;
        RECT 138.550 321.230 138.920 321.270 ;
        RECT 138.000 320.730 138.370 320.760 ;
        RECT 137.990 320.540 138.370 320.730 ;
        RECT 138.000 320.500 138.370 320.540 ;
        RECT 11.250 320.330 11.770 320.350 ;
        RECT 5.200 318.850 10.910 318.860 ;
        RECT 5.120 318.680 10.910 318.850 ;
        RECT 5.210 318.670 10.910 318.680 ;
        RECT 10.680 318.600 10.850 318.670 ;
        RECT 11.250 318.550 11.780 320.330 ;
        RECT 138.200 319.420 138.370 320.500 ;
        RECT 137.990 319.390 138.370 319.420 ;
        RECT 11.260 318.530 11.780 318.550 ;
        RECT 4.240 317.810 6.680 318.100 ;
        RECT 11.260 318.020 11.770 318.530 ;
        RECT 137.660 318.480 137.830 319.240 ;
        RECT 137.980 319.200 138.370 319.390 ;
        RECT 137.990 319.160 138.370 319.200 ;
        RECT 138.200 318.510 138.370 319.160 ;
        RECT 138.750 318.720 138.920 321.230 ;
        RECT 139.300 320.760 139.470 323.280 ;
        RECT 139.850 322.860 140.020 323.840 ;
        RECT 140.400 323.540 140.570 323.840 ;
        RECT 140.190 323.510 140.570 323.540 ;
        RECT 140.180 323.320 140.570 323.510 ;
        RECT 140.190 323.280 140.570 323.320 ;
        RECT 139.650 322.830 140.020 322.860 ;
        RECT 139.640 322.640 140.020 322.830 ;
        RECT 139.650 322.600 140.020 322.640 ;
        RECT 139.850 321.490 140.020 322.600 ;
        RECT 139.650 321.460 140.020 321.490 ;
        RECT 139.640 321.270 140.020 321.460 ;
        RECT 139.650 321.230 140.020 321.270 ;
        RECT 139.100 320.730 139.470 320.760 ;
        RECT 139.090 320.540 139.470 320.730 ;
        RECT 139.100 320.500 139.470 320.540 ;
        RECT 139.300 319.410 139.470 320.500 ;
        RECT 139.100 319.380 139.470 319.410 ;
        RECT 139.090 319.190 139.470 319.380 ;
        RECT 139.100 319.150 139.470 319.190 ;
        RECT 138.550 318.690 138.920 318.720 ;
        RECT 138.540 318.510 138.920 318.690 ;
        RECT 139.300 318.510 139.470 319.150 ;
        RECT 139.850 318.710 140.020 321.230 ;
        RECT 140.400 320.760 140.570 323.280 ;
        RECT 140.950 322.860 141.120 323.830 ;
        RECT 141.300 323.750 141.880 323.940 ;
        RECT 196.170 323.830 196.750 324.020 ;
        RECT 227.070 323.920 227.300 324.030 ;
        RECT 231.760 324.000 232.770 324.030 ;
        RECT 196.180 323.800 196.750 323.830 ;
        RECT 141.310 323.710 141.880 323.750 ;
        RECT 141.370 323.500 141.880 323.710 ;
        RECT 196.240 323.620 196.750 323.800 ;
        RECT 226.970 323.750 231.450 323.920 ;
        RECT 231.760 323.640 231.990 324.000 ;
        RECT 141.320 323.470 141.880 323.500 ;
        RECT 229.950 323.470 230.280 323.640 ;
        RECT 230.910 323.470 231.240 323.640 ;
        RECT 231.760 323.470 232.200 323.640 ;
        RECT 232.830 323.470 233.160 323.640 ;
        RECT 141.310 323.280 141.890 323.470 ;
        RECT 141.320 323.240 141.890 323.280 ;
        RECT 231.760 323.240 231.990 323.470 ;
        RECT 141.370 323.220 141.890 323.240 ;
        RECT 141.380 323.140 141.890 323.220 ;
        RECT 228.220 323.070 231.990 323.240 ;
        RECT 231.760 322.960 231.990 323.070 ;
        RECT 140.750 322.830 141.120 322.860 ;
        RECT 140.740 322.640 141.120 322.830 ;
        RECT 140.750 322.600 141.120 322.640 ;
        RECT 140.950 321.490 141.120 322.600 ;
        RECT 142.950 322.510 145.340 322.880 ;
        RECT 229.950 322.790 230.280 322.960 ;
        RECT 230.910 322.790 231.240 322.960 ;
        RECT 231.760 322.790 232.200 322.960 ;
        RECT 232.830 322.900 233.160 322.960 ;
        RECT 232.480 322.880 233.160 322.900 ;
        RECT 232.460 322.790 233.160 322.880 ;
        RECT 140.750 321.460 141.120 321.490 ;
        RECT 140.740 321.270 141.120 321.460 ;
        RECT 140.750 321.230 141.120 321.270 ;
        RECT 140.190 320.730 140.570 320.760 ;
        RECT 140.180 320.540 140.570 320.730 ;
        RECT 140.190 320.500 140.570 320.540 ;
        RECT 140.400 319.390 140.570 320.500 ;
        RECT 140.190 319.360 140.570 319.390 ;
        RECT 140.180 319.170 140.570 319.360 ;
        RECT 140.190 319.130 140.570 319.170 ;
        RECT 139.650 318.680 140.020 318.710 ;
        RECT 139.640 318.510 140.020 318.680 ;
        RECT 140.400 318.510 140.570 319.130 ;
        RECT 140.950 318.710 141.120 321.230 ;
        RECT 143.000 319.250 145.340 322.510 ;
        RECT 227.070 322.320 227.300 322.430 ;
        RECT 226.970 322.150 231.470 322.320 ;
        RECT 231.760 322.030 231.990 322.790 ;
        RECT 232.460 322.710 232.910 322.790 ;
        RECT 232.480 322.690 232.910 322.710 ;
        RECT 229.950 321.860 230.280 322.030 ;
        RECT 230.910 321.860 231.240 322.030 ;
        RECT 231.760 321.860 232.200 322.030 ;
        RECT 232.830 321.860 233.160 322.030 ;
        RECT 231.760 321.630 231.990 321.860 ;
        RECT 228.230 321.460 231.990 321.630 ;
        RECT 231.760 321.350 231.990 321.460 ;
        RECT 228.530 321.270 228.960 321.290 ;
        RECT 228.510 321.100 228.960 321.270 ;
        RECT 229.950 321.180 230.280 321.350 ;
        RECT 230.910 321.180 231.240 321.350 ;
        RECT 231.760 321.180 232.200 321.350 ;
        RECT 232.830 321.290 233.160 321.350 ;
        RECT 232.480 321.270 233.160 321.290 ;
        RECT 232.460 321.180 233.160 321.270 ;
        RECT 228.530 321.080 228.960 321.100 ;
        RECT 227.070 320.700 227.300 320.810 ;
        RECT 226.970 320.530 231.470 320.700 ;
        RECT 231.760 320.030 231.990 321.180 ;
        RECT 232.460 321.100 232.910 321.180 ;
        RECT 232.480 321.080 232.910 321.100 ;
        RECT 228.220 320.020 231.990 320.030 ;
        RECT 228.210 319.860 231.990 320.020 ;
        RECT 228.210 319.850 228.540 319.860 ;
        RECT 230.130 319.850 230.460 319.860 ;
        RECT 231.090 319.850 231.420 319.860 ;
        RECT 230.750 319.410 231.180 319.430 ;
        RECT 143.000 319.240 145.330 319.250 ;
        RECT 230.750 319.240 231.200 319.410 ;
        RECT 230.750 319.220 231.180 319.240 ;
        RECT 227.070 319.100 227.300 319.210 ;
        RECT 226.970 318.930 231.420 319.100 ;
        RECT 231.760 318.870 231.990 319.860 ;
        RECT 232.470 319.660 232.900 319.680 ;
        RECT 232.450 319.490 232.900 319.660 ;
        RECT 232.470 319.470 232.900 319.490 ;
        RECT 140.740 318.680 141.120 318.710 ;
        RECT 229.950 318.700 230.280 318.870 ;
        RECT 230.910 318.700 231.240 318.870 ;
        RECT 231.760 318.700 232.200 318.870 ;
        RECT 232.830 318.700 233.160 318.870 ;
        RECT 140.730 318.510 141.120 318.680 ;
        RECT 138.540 318.500 138.870 318.510 ;
        RECT 138.550 318.460 138.870 318.500 ;
        RECT 139.640 318.490 139.970 318.510 ;
        RECT 140.730 318.490 141.060 318.510 ;
        RECT 139.650 318.450 139.970 318.490 ;
        RECT 140.740 318.450 141.060 318.490 ;
        RECT 231.760 318.410 231.990 318.700 ;
        RECT 228.200 318.240 231.990 318.410 ;
        RECT 231.760 318.190 231.990 318.240 ;
        RECT 229.950 318.020 230.280 318.190 ;
        RECT 230.910 318.020 231.240 318.190 ;
        RECT 231.760 318.020 232.200 318.190 ;
        RECT 232.830 318.060 233.160 318.190 ;
        RECT 232.480 318.040 233.160 318.060 ;
        RECT 232.460 318.020 233.160 318.040 ;
        RECT 11.260 317.810 11.790 318.020 ;
        RECT 4.240 317.330 11.790 317.810 ;
        RECT 227.070 317.480 227.300 317.590 ;
        RECT 4.240 317.300 11.600 317.330 ;
        RECT 226.970 317.310 231.470 317.480 ;
        RECT 231.760 317.200 231.990 318.020 ;
        RECT 232.460 317.870 232.910 318.020 ;
        RECT 232.480 317.850 232.910 317.870 ;
        RECT 232.180 317.830 232.610 317.850 ;
        RECT 232.160 317.660 232.610 317.830 ;
        RECT 232.180 317.640 232.610 317.660 ;
        RECT 229.950 317.030 230.280 317.200 ;
        RECT 230.910 317.030 231.240 317.200 ;
        RECT 231.760 317.030 232.200 317.200 ;
        RECT 232.830 317.030 233.160 317.200 ;
        RECT 231.760 316.790 231.990 317.030 ;
        RECT 228.200 316.620 231.990 316.790 ;
        RECT 231.760 316.520 231.990 316.620 ;
        RECT 229.950 316.350 230.280 316.520 ;
        RECT 230.910 316.350 231.240 316.520 ;
        RECT 231.760 316.350 232.200 316.520 ;
        RECT 232.830 316.450 233.160 316.520 ;
        RECT 232.470 316.430 233.160 316.450 ;
        RECT 232.450 316.350 233.160 316.430 ;
        RECT 4.240 315.540 11.770 316.090 ;
        RECT 227.070 315.880 227.300 315.990 ;
        RECT 226.970 315.710 231.390 315.880 ;
        RECT 231.760 315.590 231.990 316.350 ;
        RECT 232.450 316.260 232.900 316.350 ;
        RECT 232.470 316.240 232.900 316.260 ;
        RECT 2.550 302.570 4.030 302.820 ;
        RECT 4.240 302.630 4.750 315.540 ;
        RECT 11.100 315.530 11.770 315.540 ;
        RECT 7.400 314.640 10.860 315.080 ;
        RECT 5.470 314.540 10.860 314.640 ;
        RECT 5.470 314.470 10.750 314.540 ;
        RECT 5.470 303.560 5.640 314.470 ;
        RECT 5.970 314.060 10.200 314.080 ;
        RECT 5.950 303.950 10.280 314.060 ;
        RECT 6.010 303.900 6.180 303.950 ;
        RECT 10.580 303.560 10.750 314.470 ;
        RECT 5.470 303.390 10.750 303.560 ;
        RECT 10.510 303.380 10.750 303.390 ;
        RECT 11.260 302.630 11.770 315.530 ;
        RECT 229.950 315.420 230.280 315.590 ;
        RECT 230.910 315.420 231.240 315.590 ;
        RECT 231.760 315.420 232.200 315.590 ;
        RECT 232.830 315.420 233.160 315.590 ;
        RECT 231.760 315.200 231.990 315.420 ;
        RECT 228.200 315.030 232.000 315.200 ;
        RECT 231.760 314.910 231.990 315.030 ;
        RECT 229.950 314.740 230.280 314.910 ;
        RECT 230.910 314.740 231.240 314.910 ;
        RECT 231.760 314.740 232.200 314.910 ;
        RECT 227.070 314.250 227.300 314.370 ;
        RECT 226.970 314.080 231.430 314.250 ;
        RECT 231.760 313.980 231.990 314.740 ;
        RECT 232.270 314.390 232.480 314.820 ;
        RECT 232.830 314.740 233.160 314.910 ;
        RECT 232.290 314.370 232.460 314.390 ;
        RECT 229.950 313.810 230.280 313.980 ;
        RECT 230.910 313.810 231.240 313.980 ;
        RECT 231.760 313.810 232.200 313.980 ;
        RECT 232.830 313.810 233.160 313.980 ;
        RECT 231.760 313.590 231.990 313.810 ;
        RECT 228.200 313.420 231.990 313.590 ;
        RECT 229.950 313.130 230.280 313.300 ;
        RECT 230.910 313.130 231.240 313.300 ;
        RECT 231.870 313.130 232.200 313.300 ;
        RECT 232.830 313.250 233.160 313.300 ;
        RECT 232.470 313.230 233.160 313.250 ;
        RECT 232.450 313.130 233.160 313.230 ;
        RECT 232.450 313.060 232.900 313.130 ;
        RECT 232.470 313.040 232.900 313.060 ;
        RECT 233.180 312.250 233.550 327.120 ;
        RECT 233.180 312.000 233.560 312.250 ;
        RECT 229.230 311.520 229.660 311.540 ;
        RECT 230.170 311.520 230.600 311.540 ;
        RECT 232.430 311.520 232.860 311.540 ;
        RECT 229.210 311.350 229.660 311.520 ;
        RECT 230.150 311.350 230.600 311.520 ;
        RECT 231.120 311.500 231.550 311.520 ;
        RECT 229.230 311.330 229.660 311.350 ;
        RECT 230.170 311.330 230.600 311.350 ;
        RECT 231.100 311.330 231.550 311.500 ;
        RECT 232.410 311.350 232.860 311.520 ;
        RECT 232.430 311.330 232.860 311.350 ;
        RECT 231.120 311.310 231.550 311.330 ;
        RECT 4.240 302.120 11.770 302.630 ;
        RECT 2.540 296.100 4.000 296.140 ;
        RECT 2.540 295.930 4.010 296.100 ;
        RECT 2.540 295.890 4.000 295.930 ;
        RECT 4.240 289.510 4.750 302.120 ;
        RECT 5.110 301.330 11.090 301.560 ;
        RECT 5.200 290.270 10.850 301.330 ;
        RECT 11.260 291.760 11.770 302.120 ;
        RECT 11.250 291.740 11.770 291.760 ;
        RECT 5.200 290.260 10.910 290.270 ;
        RECT 5.120 290.090 10.910 290.260 ;
        RECT 5.210 290.080 10.910 290.090 ;
        RECT 10.680 290.010 10.850 290.080 ;
        RECT 11.250 289.960 11.780 291.740 ;
        RECT 11.260 289.940 11.780 289.960 ;
        RECT 4.240 289.220 6.680 289.510 ;
        RECT 11.260 289.430 11.770 289.940 ;
        RECT 11.260 289.220 11.790 289.430 ;
        RECT 4.240 288.740 11.790 289.220 ;
        RECT 4.240 288.710 11.600 288.740 ;
        RECT 4.240 286.950 11.770 287.500 ;
        RECT 2.550 273.980 4.030 274.230 ;
        RECT 4.240 274.040 4.750 286.950 ;
        RECT 11.100 286.940 11.770 286.950 ;
        RECT 7.400 286.050 10.860 286.490 ;
        RECT 5.470 285.950 10.860 286.050 ;
        RECT 5.470 285.880 10.750 285.950 ;
        RECT 5.470 274.970 5.640 285.880 ;
        RECT 5.970 285.470 10.200 285.490 ;
        RECT 5.950 275.360 10.280 285.470 ;
        RECT 6.010 275.310 6.180 275.360 ;
        RECT 10.580 274.970 10.750 285.880 ;
        RECT 5.470 274.800 10.750 274.970 ;
        RECT 10.510 274.790 10.750 274.800 ;
        RECT 11.260 274.040 11.770 286.940 ;
        RECT 4.240 273.530 11.770 274.040 ;
        RECT 2.540 267.510 4.000 267.550 ;
        RECT 2.540 267.340 4.010 267.510 ;
        RECT 2.540 267.300 4.000 267.340 ;
        RECT 4.240 260.920 4.750 273.530 ;
        RECT 5.110 272.740 11.090 272.970 ;
        RECT 5.200 261.680 10.850 272.740 ;
        RECT 11.260 263.170 11.770 273.530 ;
        RECT 11.250 263.150 11.770 263.170 ;
        RECT 5.200 261.670 10.910 261.680 ;
        RECT 5.120 261.500 10.910 261.670 ;
        RECT 5.210 261.490 10.910 261.500 ;
        RECT 10.680 261.420 10.850 261.490 ;
        RECT 11.250 261.370 11.780 263.150 ;
        RECT 11.260 261.350 11.780 261.370 ;
        RECT 4.240 260.630 6.680 260.920 ;
        RECT 11.260 260.840 11.770 261.350 ;
        RECT 11.260 260.630 11.790 260.840 ;
        RECT 4.240 260.150 11.790 260.630 ;
        RECT 4.240 260.120 11.600 260.150 ;
        RECT 4.240 258.360 11.770 258.910 ;
        RECT 2.550 245.390 4.030 245.640 ;
        RECT 4.240 245.450 4.750 258.360 ;
        RECT 11.100 258.350 11.770 258.360 ;
        RECT 7.400 257.460 10.860 257.900 ;
        RECT 5.470 257.360 10.860 257.460 ;
        RECT 5.470 257.290 10.750 257.360 ;
        RECT 5.470 246.380 5.640 257.290 ;
        RECT 5.970 256.880 10.200 256.900 ;
        RECT 5.950 246.770 10.280 256.880 ;
        RECT 6.010 246.720 6.180 246.770 ;
        RECT 10.580 246.380 10.750 257.290 ;
        RECT 5.470 246.210 10.750 246.380 ;
        RECT 10.510 246.200 10.750 246.210 ;
        RECT 11.260 245.450 11.770 258.350 ;
        RECT 4.240 244.940 11.770 245.450 ;
        RECT 2.540 238.920 4.000 238.960 ;
        RECT 2.540 238.750 4.010 238.920 ;
        RECT 2.540 238.710 4.000 238.750 ;
        RECT 4.240 232.330 4.750 244.940 ;
        RECT 5.110 244.150 11.090 244.380 ;
        RECT 5.200 233.090 10.850 244.150 ;
        RECT 11.260 234.580 11.770 244.940 ;
        RECT 11.250 234.560 11.770 234.580 ;
        RECT 5.200 233.080 10.910 233.090 ;
        RECT 5.120 232.910 10.910 233.080 ;
        RECT 5.210 232.900 10.910 232.910 ;
        RECT 10.680 232.830 10.850 232.900 ;
        RECT 11.250 232.780 11.780 234.560 ;
        RECT 11.260 232.760 11.780 232.780 ;
        RECT 4.240 232.040 6.680 232.330 ;
        RECT 11.260 232.250 11.770 232.760 ;
        RECT 11.260 232.040 11.790 232.250 ;
        RECT 4.240 231.560 11.790 232.040 ;
        RECT 4.240 231.530 11.600 231.560 ;
        RECT 4.240 229.770 11.770 230.320 ;
        RECT 2.550 216.800 4.030 217.050 ;
        RECT 4.240 216.860 4.750 229.770 ;
        RECT 11.100 229.760 11.770 229.770 ;
        RECT 7.400 228.870 10.860 229.310 ;
        RECT 5.470 228.770 10.860 228.870 ;
        RECT 5.470 228.700 10.750 228.770 ;
        RECT 5.470 217.790 5.640 228.700 ;
        RECT 5.970 228.290 10.200 228.310 ;
        RECT 5.950 218.180 10.280 228.290 ;
        RECT 6.010 218.130 6.180 218.180 ;
        RECT 10.580 217.790 10.750 228.700 ;
        RECT 5.470 217.620 10.750 217.790 ;
        RECT 10.510 217.610 10.750 217.620 ;
        RECT 11.260 216.860 11.770 229.760 ;
        RECT 4.240 216.350 11.770 216.860 ;
        RECT 2.540 210.330 4.000 210.370 ;
        RECT 2.540 210.160 4.010 210.330 ;
        RECT 2.540 210.120 4.000 210.160 ;
        RECT 4.240 203.740 4.750 216.350 ;
        RECT 5.110 215.560 11.090 215.790 ;
        RECT 5.200 204.500 10.850 215.560 ;
        RECT 11.260 205.990 11.770 216.350 ;
        RECT 11.250 205.970 11.770 205.990 ;
        RECT 5.200 204.490 10.910 204.500 ;
        RECT 5.120 204.320 10.910 204.490 ;
        RECT 5.210 204.310 10.910 204.320 ;
        RECT 10.680 204.240 10.850 204.310 ;
        RECT 11.250 204.190 11.780 205.970 ;
        RECT 11.260 204.170 11.780 204.190 ;
        RECT 4.240 203.450 6.680 203.740 ;
        RECT 11.260 203.660 11.770 204.170 ;
        RECT 11.260 203.450 11.790 203.660 ;
        RECT 4.240 202.970 11.790 203.450 ;
        RECT 4.240 202.940 11.600 202.970 ;
        RECT 4.240 201.180 11.770 201.730 ;
        RECT 2.550 188.210 4.030 188.460 ;
        RECT 4.240 188.270 4.750 201.180 ;
        RECT 11.100 201.170 11.770 201.180 ;
        RECT 7.400 200.280 10.860 200.720 ;
        RECT 5.470 200.180 10.860 200.280 ;
        RECT 5.470 200.110 10.750 200.180 ;
        RECT 5.470 189.200 5.640 200.110 ;
        RECT 5.970 199.700 10.200 199.720 ;
        RECT 5.950 189.590 10.280 199.700 ;
        RECT 6.010 189.540 6.180 189.590 ;
        RECT 10.580 189.200 10.750 200.110 ;
        RECT 5.470 189.030 10.750 189.200 ;
        RECT 10.510 189.020 10.750 189.030 ;
        RECT 11.260 188.270 11.770 201.170 ;
        RECT 4.240 187.760 11.770 188.270 ;
        RECT 2.540 181.740 4.000 181.780 ;
        RECT 2.540 181.570 4.010 181.740 ;
        RECT 2.540 181.530 4.000 181.570 ;
        RECT 4.240 175.150 4.750 187.760 ;
        RECT 5.110 186.970 11.090 187.200 ;
        RECT 5.200 175.910 10.850 186.970 ;
        RECT 11.260 177.400 11.770 187.760 ;
        RECT 11.250 177.380 11.770 177.400 ;
        RECT 5.200 175.900 10.910 175.910 ;
        RECT 5.120 175.730 10.910 175.900 ;
        RECT 5.210 175.720 10.910 175.730 ;
        RECT 10.680 175.650 10.850 175.720 ;
        RECT 11.250 175.600 11.780 177.380 ;
        RECT 11.260 175.580 11.780 175.600 ;
        RECT 4.240 174.860 6.680 175.150 ;
        RECT 11.260 175.070 11.770 175.580 ;
        RECT 11.260 174.860 11.790 175.070 ;
        RECT 4.240 174.380 11.790 174.860 ;
        RECT 4.240 174.350 11.600 174.380 ;
        RECT 4.240 172.590 11.770 173.140 ;
        RECT 2.550 159.620 4.030 159.870 ;
        RECT 4.240 159.680 4.750 172.590 ;
        RECT 11.100 172.580 11.770 172.590 ;
        RECT 7.400 171.690 10.860 172.130 ;
        RECT 5.470 171.590 10.860 171.690 ;
        RECT 5.470 171.520 10.750 171.590 ;
        RECT 5.470 160.610 5.640 171.520 ;
        RECT 5.970 171.110 10.200 171.130 ;
        RECT 5.950 161.000 10.280 171.110 ;
        RECT 6.010 160.950 6.180 161.000 ;
        RECT 10.580 160.610 10.750 171.520 ;
        RECT 5.470 160.440 10.750 160.610 ;
        RECT 10.510 160.430 10.750 160.440 ;
        RECT 11.260 159.680 11.770 172.580 ;
        RECT 4.240 159.170 11.770 159.680 ;
        RECT 2.540 153.150 4.000 153.190 ;
        RECT 2.540 152.980 4.010 153.150 ;
        RECT 2.540 152.940 4.000 152.980 ;
        RECT 4.240 146.560 4.750 159.170 ;
        RECT 5.110 158.380 11.090 158.610 ;
        RECT 5.200 147.320 10.850 158.380 ;
        RECT 11.260 148.810 11.770 159.170 ;
        RECT 11.250 148.790 11.770 148.810 ;
        RECT 5.200 147.310 10.910 147.320 ;
        RECT 5.120 147.140 10.910 147.310 ;
        RECT 5.210 147.130 10.910 147.140 ;
        RECT 10.680 147.060 10.850 147.130 ;
        RECT 11.250 147.010 11.780 148.790 ;
        RECT 11.260 146.990 11.780 147.010 ;
        RECT 4.240 146.270 6.680 146.560 ;
        RECT 11.260 146.480 11.770 146.990 ;
        RECT 11.260 146.270 11.790 146.480 ;
        RECT 4.240 145.790 11.790 146.270 ;
        RECT 4.240 145.760 11.600 145.790 ;
        RECT 4.240 144.000 11.770 144.550 ;
        RECT 2.550 131.030 4.030 131.280 ;
        RECT 4.240 131.090 4.750 144.000 ;
        RECT 11.100 143.990 11.770 144.000 ;
        RECT 7.400 143.100 10.860 143.540 ;
        RECT 5.470 143.000 10.860 143.100 ;
        RECT 5.470 142.930 10.750 143.000 ;
        RECT 5.470 132.020 5.640 142.930 ;
        RECT 5.970 142.520 10.200 142.540 ;
        RECT 5.950 132.410 10.280 142.520 ;
        RECT 6.010 132.360 6.180 132.410 ;
        RECT 10.580 132.020 10.750 142.930 ;
        RECT 5.470 131.850 10.750 132.020 ;
        RECT 10.510 131.840 10.750 131.850 ;
        RECT 11.260 131.090 11.770 143.990 ;
        RECT 4.240 130.580 11.770 131.090 ;
        RECT 2.540 124.560 4.000 124.600 ;
        RECT 2.540 124.390 4.010 124.560 ;
        RECT 2.540 124.350 4.000 124.390 ;
        RECT 4.240 117.970 4.750 130.580 ;
        RECT 5.110 129.790 11.090 130.020 ;
        RECT 5.200 118.730 10.850 129.790 ;
        RECT 11.260 120.220 11.770 130.580 ;
        RECT 11.250 120.200 11.770 120.220 ;
        RECT 5.200 118.720 10.910 118.730 ;
        RECT 5.120 118.550 10.910 118.720 ;
        RECT 5.210 118.540 10.910 118.550 ;
        RECT 10.680 118.470 10.850 118.540 ;
        RECT 11.250 118.420 11.780 120.200 ;
        RECT 11.260 118.400 11.780 118.420 ;
        RECT 4.240 117.680 6.680 117.970 ;
        RECT 11.260 117.890 11.770 118.400 ;
        RECT 11.260 117.680 11.790 117.890 ;
        RECT 4.240 117.200 11.790 117.680 ;
        RECT 4.240 117.170 11.600 117.200 ;
        RECT 4.240 115.410 11.770 115.960 ;
        RECT 2.550 102.440 4.030 102.690 ;
        RECT 4.240 102.500 4.750 115.410 ;
        RECT 11.100 115.400 11.770 115.410 ;
        RECT 7.400 114.510 10.860 114.950 ;
        RECT 5.470 114.410 10.860 114.510 ;
        RECT 5.470 114.340 10.750 114.410 ;
        RECT 5.470 103.430 5.640 114.340 ;
        RECT 5.970 113.930 10.200 113.950 ;
        RECT 5.950 103.820 10.280 113.930 ;
        RECT 6.010 103.770 6.180 103.820 ;
        RECT 10.580 103.430 10.750 114.340 ;
        RECT 5.470 103.260 10.750 103.430 ;
        RECT 10.510 103.250 10.750 103.260 ;
        RECT 11.260 102.500 11.770 115.400 ;
        RECT 4.240 101.990 11.770 102.500 ;
        RECT 2.540 95.970 4.000 96.010 ;
        RECT 2.540 95.800 4.010 95.970 ;
        RECT 2.540 95.760 4.000 95.800 ;
        RECT 4.240 89.380 4.750 101.990 ;
        RECT 5.110 101.200 11.090 101.430 ;
        RECT 5.200 90.140 10.850 101.200 ;
        RECT 11.260 91.630 11.770 101.990 ;
        RECT 11.250 91.610 11.770 91.630 ;
        RECT 5.200 90.130 10.910 90.140 ;
        RECT 5.120 89.960 10.910 90.130 ;
        RECT 5.210 89.950 10.910 89.960 ;
        RECT 10.680 89.880 10.850 89.950 ;
        RECT 11.250 89.830 11.780 91.610 ;
        RECT 11.260 89.810 11.780 89.830 ;
        RECT 4.240 89.090 6.680 89.380 ;
        RECT 11.260 89.300 11.770 89.810 ;
        RECT 11.260 89.090 11.790 89.300 ;
        RECT 4.240 88.610 11.790 89.090 ;
        RECT 4.240 88.580 11.600 88.610 ;
        RECT 4.240 86.820 11.770 87.370 ;
        RECT 2.550 73.850 4.030 74.100 ;
        RECT 4.240 73.910 4.750 86.820 ;
        RECT 11.100 86.810 11.770 86.820 ;
        RECT 7.400 85.920 10.860 86.360 ;
        RECT 5.470 85.820 10.860 85.920 ;
        RECT 5.470 85.750 10.750 85.820 ;
        RECT 5.470 74.840 5.640 85.750 ;
        RECT 5.970 85.340 10.200 85.360 ;
        RECT 5.950 75.230 10.280 85.340 ;
        RECT 6.010 75.180 6.180 75.230 ;
        RECT 10.580 74.840 10.750 85.750 ;
        RECT 5.470 74.670 10.750 74.840 ;
        RECT 10.510 74.660 10.750 74.670 ;
        RECT 11.260 73.910 11.770 86.810 ;
        RECT 4.240 73.400 11.770 73.910 ;
        RECT 2.540 67.380 4.000 67.420 ;
        RECT 2.540 67.210 4.010 67.380 ;
        RECT 2.540 67.170 4.000 67.210 ;
        RECT 4.240 60.790 4.750 73.400 ;
        RECT 5.110 72.610 11.090 72.840 ;
        RECT 5.200 61.550 10.850 72.610 ;
        RECT 11.260 63.040 11.770 73.400 ;
        RECT 11.250 63.020 11.770 63.040 ;
        RECT 5.200 61.540 10.910 61.550 ;
        RECT 5.120 61.370 10.910 61.540 ;
        RECT 5.210 61.360 10.910 61.370 ;
        RECT 10.680 61.290 10.850 61.360 ;
        RECT 11.250 61.240 11.780 63.020 ;
        RECT 11.260 61.220 11.780 61.240 ;
        RECT 4.240 60.500 6.680 60.790 ;
        RECT 11.260 60.710 11.770 61.220 ;
        RECT 11.260 60.500 11.790 60.710 ;
        RECT 4.240 60.020 11.790 60.500 ;
        RECT 4.240 59.990 11.600 60.020 ;
        RECT 4.240 58.230 11.770 58.780 ;
        RECT 2.550 45.260 4.030 45.510 ;
        RECT 4.240 45.320 4.750 58.230 ;
        RECT 11.100 58.220 11.770 58.230 ;
        RECT 7.400 57.330 10.860 57.770 ;
        RECT 5.470 57.230 10.860 57.330 ;
        RECT 5.470 57.160 10.750 57.230 ;
        RECT 5.470 46.250 5.640 57.160 ;
        RECT 5.970 56.750 10.200 56.770 ;
        RECT 5.950 46.640 10.280 56.750 ;
        RECT 6.010 46.590 6.180 46.640 ;
        RECT 10.580 46.250 10.750 57.160 ;
        RECT 5.470 46.080 10.750 46.250 ;
        RECT 10.510 46.070 10.750 46.080 ;
        RECT 11.260 45.320 11.770 58.220 ;
        RECT 4.240 44.810 11.770 45.320 ;
        RECT 2.540 38.790 4.000 38.830 ;
        RECT 2.540 38.620 4.010 38.790 ;
        RECT 2.540 38.580 4.000 38.620 ;
        RECT 4.240 32.200 4.750 44.810 ;
        RECT 5.110 44.020 11.090 44.250 ;
        RECT 5.200 32.960 10.850 44.020 ;
        RECT 11.260 34.450 11.770 44.810 ;
        RECT 11.250 34.430 11.770 34.450 ;
        RECT 5.200 32.950 10.910 32.960 ;
        RECT 5.120 32.780 10.910 32.950 ;
        RECT 5.210 32.770 10.910 32.780 ;
        RECT 10.680 32.700 10.850 32.770 ;
        RECT 11.250 32.650 11.780 34.430 ;
        RECT 11.260 32.630 11.780 32.650 ;
        RECT 4.240 31.910 6.680 32.200 ;
        RECT 11.260 32.120 11.770 32.630 ;
        RECT 11.260 31.910 11.790 32.120 ;
        RECT 4.240 31.430 11.790 31.910 ;
        RECT 4.240 31.400 11.600 31.430 ;
        RECT 4.240 29.640 11.770 30.190 ;
        RECT 2.550 16.670 4.030 16.920 ;
        RECT 4.240 16.730 4.750 29.640 ;
        RECT 11.100 29.630 11.770 29.640 ;
        RECT 7.400 28.740 10.860 29.180 ;
        RECT 5.470 28.640 10.860 28.740 ;
        RECT 5.470 28.570 10.750 28.640 ;
        RECT 5.470 17.660 5.640 28.570 ;
        RECT 5.970 28.160 10.200 28.180 ;
        RECT 5.950 18.050 10.280 28.160 ;
        RECT 6.010 18.000 6.180 18.050 ;
        RECT 10.580 17.660 10.750 28.570 ;
        RECT 5.470 17.490 10.750 17.660 ;
        RECT 10.510 17.480 10.750 17.490 ;
        RECT 11.260 16.730 11.770 29.630 ;
        RECT 4.240 16.220 11.770 16.730 ;
        RECT 2.540 10.200 4.000 10.240 ;
        RECT 2.540 10.030 4.010 10.200 ;
        RECT 2.540 9.990 4.000 10.030 ;
        RECT 4.240 3.610 4.750 16.220 ;
        RECT 5.110 15.430 11.090 15.660 ;
        RECT 5.200 4.370 10.850 15.430 ;
        RECT 11.260 5.860 11.770 16.220 ;
        RECT 11.250 5.840 11.770 5.860 ;
        RECT 5.200 4.360 10.910 4.370 ;
        RECT 5.120 4.190 10.910 4.360 ;
        RECT 5.210 4.180 10.910 4.190 ;
        RECT 10.680 4.110 10.850 4.180 ;
        RECT 11.250 4.060 11.780 5.840 ;
        RECT 11.260 4.040 11.780 4.060 ;
        RECT 4.240 3.320 6.680 3.610 ;
        RECT 11.260 3.530 11.770 4.040 ;
        RECT 11.260 3.320 11.790 3.530 ;
        RECT 4.240 2.840 11.790 3.320 ;
        RECT 4.240 2.810 11.600 2.840 ;
      LAYER mcon ;
        RECT 150.320 387.610 150.490 387.780 ;
        RECT 23.700 386.870 23.870 387.040 ;
        RECT 23.700 386.510 23.870 386.680 ;
        RECT 23.700 386.140 23.870 386.310 ;
        RECT 30.380 387.190 30.550 387.360 ;
        RECT 30.380 386.830 30.550 387.000 ;
        RECT 30.380 386.470 30.550 386.640 ;
        RECT 30.380 386.110 30.550 386.280 ;
        RECT 52.290 386.870 52.460 387.040 ;
        RECT 52.290 386.510 52.460 386.680 ;
        RECT 52.290 386.140 52.460 386.310 ;
        RECT 58.970 387.190 59.140 387.360 ;
        RECT 58.970 386.830 59.140 387.000 ;
        RECT 58.970 386.470 59.140 386.640 ;
        RECT 58.970 386.110 59.140 386.280 ;
        RECT 80.880 386.870 81.050 387.040 ;
        RECT 80.880 386.510 81.050 386.680 ;
        RECT 80.880 386.140 81.050 386.310 ;
        RECT 87.560 387.190 87.730 387.360 ;
        RECT 87.560 386.830 87.730 387.000 ;
        RECT 150.320 387.250 150.490 387.420 ;
        RECT 150.320 386.890 150.490 387.060 ;
        RECT 87.560 386.470 87.730 386.640 ;
        RECT 150.320 386.530 150.490 386.700 ;
        RECT 157.070 387.440 157.240 387.610 ;
        RECT 157.070 387.080 157.240 387.250 ;
        RECT 157.070 386.720 157.240 386.890 ;
        RECT 164.900 386.870 165.070 387.040 ;
        RECT 164.900 386.510 165.070 386.680 ;
        RECT 87.560 386.110 87.730 386.280 ;
        RECT 164.900 386.140 165.070 386.310 ;
        RECT 171.580 387.190 171.750 387.360 ;
        RECT 171.580 386.830 171.750 387.000 ;
        RECT 171.580 386.470 171.750 386.640 ;
        RECT 193.490 386.870 193.660 387.040 ;
        RECT 193.490 386.510 193.660 386.680 ;
        RECT 171.580 386.110 171.750 386.280 ;
        RECT 129.870 385.920 153.770 386.090 ;
        RECT 162.650 385.920 183.820 386.090 ;
        RECT 193.490 386.140 193.660 386.310 ;
        RECT 200.170 387.190 200.340 387.360 ;
        RECT 200.170 386.830 200.340 387.000 ;
        RECT 200.170 386.470 200.340 386.640 ;
        RECT 200.170 386.110 200.340 386.280 ;
        RECT 222.080 386.870 222.250 387.040 ;
        RECT 222.080 386.510 222.250 386.680 ;
        RECT 222.080 386.140 222.250 386.310 ;
        RECT 228.760 387.190 228.930 387.360 ;
        RECT 228.760 386.830 228.930 387.000 ;
        RECT 228.760 386.470 228.930 386.640 ;
        RECT 228.760 386.110 228.930 386.280 ;
        RECT 250.670 386.870 250.840 387.040 ;
        RECT 250.670 386.510 250.840 386.680 ;
        RECT 250.670 386.140 250.840 386.310 ;
        RECT 257.350 387.190 257.520 387.360 ;
        RECT 257.350 386.830 257.520 387.000 ;
        RECT 257.350 386.470 257.520 386.640 ;
        RECT 257.350 386.110 257.520 386.280 ;
        RECT 279.260 386.870 279.430 387.040 ;
        RECT 279.260 386.510 279.430 386.680 ;
        RECT 279.260 386.140 279.430 386.310 ;
        RECT 285.940 387.190 286.110 387.360 ;
        RECT 285.940 386.830 286.110 387.000 ;
        RECT 285.940 386.470 286.110 386.640 ;
        RECT 285.940 386.110 286.110 386.280 ;
        RECT 307.850 386.870 308.020 387.040 ;
        RECT 307.850 386.510 308.020 386.680 ;
        RECT 307.850 386.140 308.020 386.310 ;
        RECT 314.530 387.190 314.700 387.360 ;
        RECT 314.530 386.830 314.700 387.000 ;
        RECT 314.530 386.470 314.700 386.640 ;
        RECT 314.530 386.110 314.700 386.280 ;
        RECT 336.440 386.870 336.610 387.040 ;
        RECT 336.440 386.510 336.610 386.680 ;
        RECT 336.440 386.140 336.610 386.310 ;
        RECT 343.120 387.190 343.290 387.360 ;
        RECT 343.120 386.830 343.290 387.000 ;
        RECT 343.120 386.470 343.290 386.640 ;
        RECT 343.120 386.110 343.290 386.280 ;
        RECT 16.560 385.520 18.420 385.530 ;
        RECT 16.560 385.350 18.430 385.520 ;
        RECT 39.920 385.340 43.080 385.520 ;
        RECT 16.600 383.260 16.780 385.160 ;
        RECT 17.000 383.250 17.180 385.160 ;
        RECT 18.190 384.220 29.170 384.390 ;
        RECT 18.190 383.600 29.170 383.770 ;
        RECT 18.200 382.980 29.180 383.150 ;
        RECT 18.220 382.400 29.200 382.570 ;
        RECT 18.230 381.810 29.210 381.980 ;
        RECT 18.230 381.210 29.210 381.380 ;
        RECT 18.180 380.610 29.160 380.780 ;
        RECT 18.190 380.000 29.170 380.170 ;
        RECT 18.180 379.400 29.160 379.570 ;
        RECT 31.920 383.460 41.370 383.630 ;
        RECT 31.910 382.710 41.300 382.880 ;
        RECT 31.940 381.990 41.340 382.160 ;
        RECT 31.950 381.330 41.320 381.500 ;
        RECT 31.940 380.680 41.390 380.850 ;
        RECT 31.950 380.040 41.340 380.210 ;
        RECT 43.490 384.360 43.690 385.290 ;
        RECT 42.420 379.120 42.770 382.420 ;
        RECT 45.150 385.520 47.010 385.530 ;
        RECT 45.150 385.350 47.020 385.520 ;
        RECT 68.510 385.340 71.670 385.520 ;
        RECT 45.190 383.260 45.370 385.160 ;
        RECT 45.590 383.250 45.770 385.160 ;
        RECT 46.780 384.220 57.760 384.390 ;
        RECT 46.780 383.600 57.760 383.770 ;
        RECT 46.790 382.980 57.770 383.150 ;
        RECT 46.810 382.400 57.790 382.570 ;
        RECT 46.820 381.810 57.800 381.980 ;
        RECT 46.820 381.210 57.800 381.380 ;
        RECT 46.770 380.610 57.750 380.780 ;
        RECT 46.780 380.000 57.760 380.170 ;
        RECT 46.770 379.400 57.750 379.570 ;
        RECT 60.510 383.460 69.960 383.630 ;
        RECT 60.500 382.710 69.890 382.880 ;
        RECT 60.530 381.990 69.930 382.160 ;
        RECT 60.540 381.330 69.910 381.500 ;
        RECT 60.530 380.680 69.980 380.850 ;
        RECT 60.540 380.040 69.930 380.210 ;
        RECT 72.080 384.360 72.280 385.290 ;
        RECT 71.010 379.120 71.360 382.420 ;
        RECT 73.740 385.520 75.600 385.530 ;
        RECT 73.740 385.350 75.610 385.520 ;
        RECT 97.100 385.340 100.260 385.520 ;
        RECT 73.780 383.260 73.960 385.160 ;
        RECT 74.180 383.250 74.360 385.160 ;
        RECT 75.370 384.220 86.350 384.390 ;
        RECT 75.370 383.600 86.350 383.770 ;
        RECT 75.380 382.980 86.360 383.150 ;
        RECT 75.400 382.400 86.380 382.570 ;
        RECT 75.410 381.810 86.390 381.980 ;
        RECT 75.410 381.210 86.390 381.380 ;
        RECT 75.360 380.610 86.340 380.780 ;
        RECT 75.370 380.000 86.350 380.170 ;
        RECT 75.360 379.400 86.340 379.570 ;
        RECT 89.100 383.460 98.550 383.630 ;
        RECT 89.090 382.710 98.480 382.880 ;
        RECT 89.120 381.990 98.520 382.160 ;
        RECT 89.130 381.330 98.500 381.500 ;
        RECT 89.120 380.680 98.570 380.850 ;
        RECT 89.130 380.040 98.520 380.210 ;
        RECT 100.670 384.360 100.870 385.290 ;
        RECT 99.600 379.120 99.950 382.420 ;
        RECT 119.480 379.350 119.650 379.520 ;
        RECT 157.760 385.520 159.620 385.530 ;
        RECT 157.760 385.350 159.630 385.520 ;
        RECT 181.120 385.340 184.280 385.520 ;
        RECT 157.800 383.260 157.980 385.160 ;
        RECT 158.200 383.250 158.380 385.160 ;
        RECT 159.390 384.220 170.370 384.390 ;
        RECT 159.390 383.600 170.370 383.770 ;
        RECT 138.870 379.710 139.040 379.880 ;
        RECT 138.870 379.260 139.040 379.430 ;
        RECT 159.400 382.980 170.380 383.150 ;
        RECT 159.420 382.400 170.400 382.570 ;
        RECT 159.430 381.810 170.410 381.980 ;
        RECT 159.430 381.210 170.410 381.380 ;
        RECT 159.380 380.610 170.360 380.780 ;
        RECT 159.390 380.000 170.370 380.170 ;
        RECT 159.380 379.400 170.360 379.570 ;
        RECT 173.120 383.460 182.570 383.630 ;
        RECT 173.110 382.710 182.500 382.880 ;
        RECT 173.140 381.990 182.540 382.160 ;
        RECT 173.150 381.330 182.520 381.500 ;
        RECT 173.140 380.680 182.590 380.850 ;
        RECT 173.150 380.040 182.540 380.210 ;
        RECT 183.620 379.120 183.970 382.420 ;
        RECT 184.690 384.360 184.890 385.290 ;
        RECT 186.350 385.520 188.210 385.530 ;
        RECT 186.350 385.350 188.220 385.520 ;
        RECT 209.710 385.340 212.870 385.520 ;
        RECT 186.390 383.260 186.570 385.160 ;
        RECT 186.790 383.250 186.970 385.160 ;
        RECT 187.980 384.220 198.960 384.390 ;
        RECT 187.980 383.600 198.960 383.770 ;
        RECT 187.990 382.980 198.970 383.150 ;
        RECT 188.010 382.400 198.990 382.570 ;
        RECT 188.020 381.810 199.000 381.980 ;
        RECT 188.020 381.210 199.000 381.380 ;
        RECT 187.970 380.610 198.950 380.780 ;
        RECT 187.980 380.000 198.960 380.170 ;
        RECT 187.970 379.400 198.950 379.570 ;
        RECT 201.710 383.460 211.160 383.630 ;
        RECT 201.700 382.710 211.090 382.880 ;
        RECT 201.730 381.990 211.130 382.160 ;
        RECT 201.740 381.330 211.110 381.500 ;
        RECT 201.730 380.680 211.180 380.850 ;
        RECT 201.740 380.040 211.130 380.210 ;
        RECT 213.280 384.360 213.480 385.290 ;
        RECT 212.210 379.120 212.560 382.420 ;
        RECT 214.940 385.520 216.800 385.530 ;
        RECT 214.940 385.350 216.810 385.520 ;
        RECT 238.300 385.340 241.460 385.520 ;
        RECT 214.980 383.260 215.160 385.160 ;
        RECT 215.380 383.250 215.560 385.160 ;
        RECT 216.570 384.220 227.550 384.390 ;
        RECT 216.570 383.600 227.550 383.770 ;
        RECT 216.580 382.980 227.560 383.150 ;
        RECT 216.600 382.400 227.580 382.570 ;
        RECT 216.610 381.810 227.590 381.980 ;
        RECT 216.610 381.210 227.590 381.380 ;
        RECT 216.560 380.610 227.540 380.780 ;
        RECT 216.570 380.000 227.550 380.170 ;
        RECT 216.560 379.400 227.540 379.570 ;
        RECT 230.300 383.460 239.750 383.630 ;
        RECT 230.290 382.710 239.680 382.880 ;
        RECT 230.320 381.990 239.720 382.160 ;
        RECT 230.330 381.330 239.700 381.500 ;
        RECT 230.320 380.680 239.770 380.850 ;
        RECT 230.330 380.040 239.720 380.210 ;
        RECT 241.870 384.360 242.070 385.290 ;
        RECT 240.800 379.120 241.150 382.420 ;
        RECT 243.530 385.520 245.390 385.530 ;
        RECT 243.530 385.350 245.400 385.520 ;
        RECT 266.890 385.340 270.050 385.520 ;
        RECT 243.570 383.260 243.750 385.160 ;
        RECT 243.970 383.250 244.150 385.160 ;
        RECT 245.160 384.220 256.140 384.390 ;
        RECT 245.160 383.600 256.140 383.770 ;
        RECT 245.170 382.980 256.150 383.150 ;
        RECT 245.190 382.400 256.170 382.570 ;
        RECT 245.200 381.810 256.180 381.980 ;
        RECT 245.200 381.210 256.180 381.380 ;
        RECT 245.150 380.610 256.130 380.780 ;
        RECT 245.160 380.000 256.140 380.170 ;
        RECT 245.150 379.400 256.130 379.570 ;
        RECT 258.890 383.460 268.340 383.630 ;
        RECT 258.880 382.710 268.270 382.880 ;
        RECT 258.910 381.990 268.310 382.160 ;
        RECT 258.920 381.330 268.290 381.500 ;
        RECT 258.910 380.680 268.360 380.850 ;
        RECT 258.920 380.040 268.310 380.210 ;
        RECT 270.460 384.360 270.660 385.290 ;
        RECT 269.390 379.120 269.740 382.420 ;
        RECT 272.120 385.520 273.980 385.530 ;
        RECT 272.120 385.350 273.990 385.520 ;
        RECT 295.480 385.340 298.640 385.520 ;
        RECT 272.160 383.260 272.340 385.160 ;
        RECT 272.560 383.250 272.740 385.160 ;
        RECT 273.750 384.220 284.730 384.390 ;
        RECT 273.750 383.600 284.730 383.770 ;
        RECT 273.760 382.980 284.740 383.150 ;
        RECT 273.780 382.400 284.760 382.570 ;
        RECT 273.790 381.810 284.770 381.980 ;
        RECT 273.790 381.210 284.770 381.380 ;
        RECT 273.740 380.610 284.720 380.780 ;
        RECT 273.750 380.000 284.730 380.170 ;
        RECT 273.740 379.400 284.720 379.570 ;
        RECT 287.480 383.460 296.930 383.630 ;
        RECT 287.470 382.710 296.860 382.880 ;
        RECT 287.500 381.990 296.900 382.160 ;
        RECT 287.510 381.330 296.880 381.500 ;
        RECT 287.500 380.680 296.950 380.850 ;
        RECT 287.510 380.040 296.900 380.210 ;
        RECT 299.050 384.360 299.250 385.290 ;
        RECT 297.980 379.120 298.330 382.420 ;
        RECT 300.710 385.520 302.570 385.530 ;
        RECT 300.710 385.350 302.580 385.520 ;
        RECT 324.070 385.340 327.230 385.520 ;
        RECT 300.750 383.260 300.930 385.160 ;
        RECT 301.150 383.250 301.330 385.160 ;
        RECT 302.340 384.220 313.320 384.390 ;
        RECT 302.340 383.600 313.320 383.770 ;
        RECT 302.350 382.980 313.330 383.150 ;
        RECT 302.370 382.400 313.350 382.570 ;
        RECT 302.380 381.810 313.360 381.980 ;
        RECT 302.380 381.210 313.360 381.380 ;
        RECT 302.330 380.610 313.310 380.780 ;
        RECT 302.340 380.000 313.320 380.170 ;
        RECT 302.330 379.400 313.310 379.570 ;
        RECT 316.070 383.460 325.520 383.630 ;
        RECT 316.060 382.710 325.450 382.880 ;
        RECT 316.090 381.990 325.490 382.160 ;
        RECT 316.100 381.330 325.470 381.500 ;
        RECT 316.090 380.680 325.540 380.850 ;
        RECT 316.100 380.040 325.490 380.210 ;
        RECT 327.640 384.360 327.840 385.290 ;
        RECT 326.570 379.120 326.920 382.420 ;
        RECT 329.300 385.520 331.160 385.530 ;
        RECT 329.300 385.350 331.170 385.520 ;
        RECT 352.660 385.340 355.820 385.520 ;
        RECT 329.340 383.260 329.520 385.160 ;
        RECT 329.740 383.250 329.920 385.160 ;
        RECT 330.930 384.220 341.910 384.390 ;
        RECT 330.930 383.600 341.910 383.770 ;
        RECT 330.940 382.980 341.920 383.150 ;
        RECT 330.960 382.400 341.940 382.570 ;
        RECT 330.970 381.810 341.950 381.980 ;
        RECT 330.970 381.210 341.950 381.380 ;
        RECT 330.920 380.610 341.900 380.780 ;
        RECT 330.930 380.000 341.910 380.170 ;
        RECT 330.920 379.400 341.900 379.570 ;
        RECT 344.660 383.460 354.110 383.630 ;
        RECT 344.650 382.710 354.040 382.880 ;
        RECT 344.680 381.990 354.080 382.160 ;
        RECT 344.690 381.330 354.060 381.500 ;
        RECT 344.680 380.680 354.130 380.850 ;
        RECT 344.690 380.040 354.080 380.210 ;
        RECT 356.230 384.360 356.430 385.290 ;
        RECT 355.160 379.120 355.510 382.420 ;
        RECT 156.340 377.960 156.510 378.130 ;
        RECT 156.710 377.960 156.880 378.130 ;
        RECT 157.070 377.960 157.240 378.130 ;
        RECT 157.430 377.960 157.600 378.130 ;
        RECT 157.790 377.960 157.970 378.130 ;
        RECT 158.160 377.960 158.330 378.130 ;
        RECT 133.150 376.590 133.320 376.760 ;
        RECT 123.020 376.230 123.190 376.400 ;
        RECT 120.150 376.020 120.320 376.190 ;
        RECT 121.560 376.020 121.730 376.190 ;
        RECT 133.150 375.900 133.320 376.070 ;
        RECT 144.220 375.960 144.390 376.130 ;
        RECT 120.150 375.170 120.320 375.340 ;
        RECT 120.730 375.310 120.900 375.480 ;
        RECT 121.560 375.170 121.730 375.340 ;
        RECT 122.760 375.310 122.930 375.480 ;
        RECT 144.220 375.510 144.390 375.680 ;
        RECT 120.330 374.760 120.500 374.930 ;
        RECT 121.390 374.760 121.560 374.930 ;
        RECT 120.150 374.350 120.320 374.520 ;
        RECT 120.730 374.470 120.900 374.640 ;
        RECT 121.560 374.350 121.730 374.520 ;
        RECT 136.120 374.570 136.290 374.740 ;
        RECT 137.480 374.650 137.650 374.820 ;
        RECT 138.170 374.640 138.340 374.810 ;
        RECT 122.760 373.880 122.930 374.050 ;
        RECT 133.150 373.790 133.320 373.960 ;
        RECT 120.150 373.510 120.320 373.680 ;
        RECT 121.560 373.510 121.730 373.680 ;
        RECT 122.190 373.330 122.360 373.500 ;
        RECT 4.640 372.900 5.570 373.100 ;
        RECT 133.150 373.100 133.320 373.270 ;
        RECT 4.410 369.330 4.590 372.490 ;
        RECT 7.510 371.830 10.810 372.180 ;
        RECT 2.570 359.790 2.740 359.960 ;
        RECT 2.930 359.790 3.100 359.960 ;
        RECT 3.290 359.790 3.460 359.960 ;
        RECT 3.650 359.790 3.820 359.960 ;
        RECT 6.300 361.330 6.470 370.780 ;
        RECT 7.050 361.320 7.220 370.710 ;
        RECT 7.770 361.350 7.940 370.750 ;
        RECT 8.430 361.360 8.600 370.730 ;
        RECT 9.080 361.350 9.250 370.800 ;
        RECT 9.720 361.360 9.890 370.750 ;
        RECT 120.150 372.390 120.320 372.560 ;
        RECT 122.420 372.580 122.590 372.750 ;
        RECT 123.030 372.610 123.200 372.780 ;
        RECT 121.560 372.390 121.730 372.560 ;
        RECT 133.150 372.240 133.320 372.410 ;
        RECT 120.710 371.670 120.880 371.840 ;
        RECT 122.140 371.690 122.310 371.860 ;
        RECT 133.150 371.550 133.320 371.720 ;
        RECT 144.220 372.970 144.390 373.140 ;
        RECT 144.220 372.520 144.390 372.690 ;
        RECT 144.220 371.960 144.390 372.130 ;
        RECT 119.920 371.090 120.090 371.260 ;
        RECT 120.850 371.090 121.020 371.260 ;
        RECT 121.550 371.090 121.720 371.260 ;
        RECT 122.290 371.090 122.460 371.260 ;
        RECT 123.000 371.080 123.170 371.250 ;
        RECT 144.220 371.510 144.390 371.680 ;
        RECT 147.520 372.880 147.690 373.050 ;
        RECT 135.400 370.910 135.570 371.080 ;
        RECT 145.260 370.930 145.430 371.100 ;
        RECT 144.670 368.990 145.100 369.730 ;
        RECT 202.070 369.220 202.340 369.490 ;
        RECT 240.000 369.220 240.270 369.490 ;
        RECT 168.550 368.060 168.760 368.270 ;
        RECT 167.080 367.690 167.250 367.860 ;
        RECT 169.510 367.590 169.680 367.760 ;
        RECT 170.550 367.630 170.720 367.800 ;
        RECT 171.590 367.290 171.760 367.460 ;
        RECT 202.070 367.490 202.340 367.760 ;
        RECT 240.000 367.490 240.270 367.760 ;
        RECT 171.590 366.930 171.760 367.100 ;
        RECT 168.550 366.310 168.760 366.520 ;
        RECT 167.080 365.940 167.250 366.110 ;
        RECT 169.510 365.840 169.680 366.010 ;
        RECT 170.550 365.880 170.720 366.050 ;
        RECT 192.960 365.830 193.220 366.650 ;
        RECT 203.200 366.710 203.380 366.880 ;
        RECT 201.390 366.410 201.560 366.580 ;
        RECT 171.590 365.540 171.760 365.710 ;
        RECT 201.740 365.570 201.920 365.760 ;
        RECT 171.590 365.180 171.760 365.350 ;
        RECT 143.800 364.770 143.970 364.940 ;
        RECT 144.890 364.780 145.060 364.950 ;
        RECT 168.550 364.560 168.760 364.770 ;
        RECT 204.910 365.860 205.230 366.650 ;
        RECT 208.290 366.350 208.460 366.520 ;
        RECT 240.780 366.410 240.950 366.580 ;
        RECT 208.760 365.790 208.930 365.960 ;
        RECT 211.100 365.410 211.270 365.580 ;
        RECT 211.100 364.960 211.270 365.130 ;
        RECT 229.180 365.410 229.350 365.580 ;
        RECT 234.490 365.310 234.660 365.480 ;
        RECT 229.180 364.960 229.350 365.130 ;
        RECT 207.440 364.740 207.610 364.910 ;
        RECT 234.820 364.940 234.990 365.110 ;
        RECT 167.080 364.190 167.250 364.360 ;
        RECT 169.510 364.090 169.680 364.260 ;
        RECT 208.290 364.360 208.460 364.530 ;
        RECT 142.260 363.860 142.430 364.030 ;
        RECT 143.810 363.780 143.980 363.950 ;
        RECT 144.590 363.730 144.760 363.900 ;
        RECT 144.900 363.790 145.070 363.960 ;
        RECT 170.550 364.130 170.720 364.300 ;
        RECT 171.590 363.790 171.760 363.960 ;
        RECT 171.590 363.430 171.760 363.600 ;
        RECT 202.060 363.190 202.330 363.460 ;
        RECT 208.300 363.290 208.470 363.460 ;
        RECT 208.760 363.470 208.930 363.640 ;
        RECT 233.880 364.260 234.050 364.430 ;
        RECT 234.360 364.320 234.530 364.490 ;
        RECT 240.420 365.570 240.600 365.760 ;
        RECT 214.130 363.780 214.300 363.950 ;
        RECT 228.040 363.780 228.210 363.950 ;
        RECT 142.240 362.940 142.410 363.110 ;
        RECT 143.810 362.790 143.980 362.960 ;
        RECT 144.900 362.800 145.070 362.970 ;
        RECT 168.550 362.810 168.760 363.020 ;
        RECT 167.080 362.440 167.250 362.610 ;
        RECT 169.510 362.340 169.680 362.510 ;
        RECT 142.220 361.950 142.390 362.120 ;
        RECT 143.720 362.000 143.890 362.170 ;
        RECT 145.020 361.900 145.190 362.070 ;
        RECT 170.550 362.380 170.720 362.550 ;
        RECT 171.590 362.040 171.760 362.210 ;
        RECT 201.740 361.930 201.920 362.120 ;
        RECT 171.590 361.680 171.760 361.850 ;
        RECT 202.060 361.460 202.330 361.730 ;
        RECT 207.430 363.050 207.600 363.220 ;
        RECT 233.890 363.130 234.060 363.300 ;
        RECT 239.990 363.190 240.260 363.460 ;
        RECT 236.790 362.890 236.960 363.060 ;
        RECT 211.100 362.460 211.270 362.630 ;
        RECT 208.750 361.890 208.920 362.060 ;
        RECT 211.100 362.010 211.270 362.180 ;
        RECT 229.180 362.460 229.350 362.630 ;
        RECT 234.490 362.550 234.660 362.720 ;
        RECT 234.880 362.450 235.050 362.620 ;
        RECT 235.800 362.520 235.970 362.690 ;
        RECT 237.730 362.500 237.900 362.670 ;
        RECT 239.040 362.910 239.210 363.080 ;
        RECT 229.180 362.010 229.350 362.180 ;
        RECT 236.740 362.240 236.910 362.410 ;
        RECT 208.320 361.380 208.490 361.550 ;
        RECT 234.820 361.740 234.990 361.910 ;
        RECT 143.720 361.010 143.890 361.180 ;
        RECT 201.390 361.110 201.560 361.280 ;
        RECT 145.020 360.910 145.190 361.080 ;
        RECT 172.750 360.770 172.920 360.940 ;
        RECT 171.590 360.520 171.760 360.690 ;
        RECT 173.590 360.650 173.760 360.820 ;
        RECT 174.340 360.650 174.510 360.820 ;
        RECT 143.720 360.020 143.890 360.190 ;
        RECT 144.160 359.630 144.330 359.800 ;
        RECT 145.020 359.920 145.190 360.090 ;
        RECT 171.590 360.160 171.760 360.330 ;
        RECT 177.320 360.320 177.490 360.490 ;
        RECT 167.080 359.760 167.250 359.930 ;
        RECT 169.510 359.860 169.680 360.030 ;
        RECT 170.550 359.820 170.720 359.990 ;
        RECT 172.930 359.940 173.100 360.110 ;
        RECT 177.720 360.770 177.890 360.940 ;
        RECT 233.880 361.060 234.050 361.230 ;
        RECT 234.360 361.120 234.530 361.290 ;
        RECT 238.390 361.530 238.560 361.700 ;
        RECT 203.200 360.850 203.380 360.980 ;
        RECT 203.190 360.810 203.380 360.850 ;
        RECT 234.880 361.010 235.050 361.180 ;
        RECT 235.800 360.940 235.970 361.110 ;
        RECT 236.740 361.100 236.910 361.270 ;
        RECT 240.420 361.930 240.600 362.120 ;
        RECT 239.990 361.460 240.260 361.730 ;
        RECT 240.780 361.110 240.950 361.280 ;
        RECT 237.730 360.840 237.900 361.010 ;
        RECT 238.960 360.860 239.140 360.980 ;
        RECT 238.960 360.850 239.260 360.860 ;
        RECT 203.190 360.680 203.370 360.810 ;
        RECT 177.720 360.410 177.890 360.580 ;
        RECT 201.380 360.380 201.550 360.550 ;
        RECT 168.550 359.350 168.760 359.560 ;
        RECT 201.730 359.540 201.910 359.730 ;
        RECT 2.890 353.110 3.060 353.280 ;
        RECT 3.250 353.110 3.420 353.280 ;
        RECT 3.620 353.110 3.790 353.280 ;
        RECT 4.410 347.830 4.580 347.840 ;
        RECT 4.400 345.970 4.580 347.830 ;
        RECT 5.540 347.600 5.710 358.580 ;
        RECT 6.160 347.600 6.330 358.580 ;
        RECT 6.780 347.610 6.950 358.590 ;
        RECT 7.360 347.630 7.530 358.610 ;
        RECT 7.950 347.640 8.120 358.620 ;
        RECT 8.550 347.640 8.720 358.620 ;
        RECT 9.150 347.590 9.320 358.570 ;
        RECT 9.760 347.600 9.930 358.580 ;
        RECT 10.360 347.590 10.530 358.570 ;
        RECT 171.590 358.770 171.760 358.940 ;
        RECT 172.930 359.040 173.100 359.210 ;
        RECT 177.320 358.660 177.490 358.830 ;
        RECT 171.590 358.410 171.760 358.580 ;
        RECT 167.080 358.010 167.250 358.180 ;
        RECT 169.510 358.110 169.680 358.280 ;
        RECT 170.550 358.070 170.720 358.240 ;
        RECT 173.590 358.330 173.760 358.500 ;
        RECT 174.340 358.330 174.510 358.500 ;
        RECT 176.340 358.340 176.510 358.510 ;
        RECT 177.720 358.930 177.890 359.100 ;
        RECT 177.720 358.570 177.890 358.740 ;
        RECT 214.930 359.690 215.100 359.860 ;
        RECT 233.380 360.120 233.550 360.310 ;
        RECT 233.890 360.330 234.060 360.500 ;
        RECT 236.790 360.450 236.960 360.620 ;
        RECT 238.950 360.690 239.260 360.850 ;
        RECT 240.770 360.380 240.940 360.550 ;
        RECT 233.890 359.930 234.060 360.100 ;
        RECT 236.790 359.890 236.960 360.060 ;
        RECT 239.080 359.970 239.250 360.140 ;
        RECT 207.670 359.280 207.840 359.450 ;
        RECT 212.980 359.380 213.150 359.550 ;
        RECT 212.980 358.930 213.150 359.100 ;
        RECT 229.170 359.380 229.340 359.550 ;
        RECT 237.730 359.500 237.900 359.670 ;
        RECT 233.880 359.200 234.050 359.370 ;
        RECT 234.480 359.310 234.650 359.450 ;
        RECT 234.360 359.280 234.650 359.310 ;
        RECT 234.360 359.140 234.530 359.280 ;
        RECT 234.880 359.250 235.050 359.420 ;
        RECT 235.800 359.320 235.970 359.490 ;
        RECT 229.170 358.930 229.340 359.100 ;
        RECT 236.740 359.240 236.910 359.410 ;
        RECT 238.390 358.940 238.560 359.110 ;
        RECT 232.490 358.340 232.660 358.510 ;
        RECT 234.820 358.520 234.990 358.690 ;
        RECT 240.410 359.540 240.590 359.730 ;
        RECT 168.550 357.600 168.760 357.810 ;
        RECT 214.120 357.750 214.290 357.920 ;
        RECT 172.750 357.570 172.920 357.740 ;
        RECT 173.590 357.450 173.760 357.620 ;
        RECT 174.340 357.450 174.510 357.620 ;
        RECT 171.590 357.020 171.760 357.190 ;
        RECT 177.320 357.120 177.490 357.290 ;
        RECT 171.590 356.660 171.760 356.830 ;
        RECT 172.930 356.740 173.100 356.910 ;
        RECT 177.720 357.570 177.890 357.740 ;
        RECT 228.030 357.750 228.200 357.920 ;
        RECT 236.740 358.100 236.910 358.270 ;
        RECT 234.880 357.810 235.050 357.980 ;
        RECT 235.800 357.740 235.970 357.910 ;
        RECT 237.730 357.840 237.900 358.010 ;
        RECT 177.720 357.210 177.890 357.380 ;
        RECT 232.640 357.510 232.810 357.680 ;
        RECT 236.790 357.450 236.960 357.620 ;
        RECT 239.000 357.720 239.170 357.890 ;
        RECT 233.890 357.130 234.060 357.300 ;
        RECT 167.080 356.260 167.250 356.430 ;
        RECT 169.510 356.360 169.680 356.530 ;
        RECT 170.550 356.320 170.720 356.490 ;
        RECT 168.550 355.850 168.760 356.060 ;
        RECT 172.930 355.840 173.100 356.010 ;
        RECT 201.730 355.900 201.910 356.090 ;
        RECT 177.320 355.460 177.490 355.630 ;
        RECT 171.590 355.270 171.760 355.440 ;
        RECT 171.590 354.910 171.760 355.080 ;
        RECT 173.590 355.130 173.760 355.300 ;
        RECT 174.340 355.130 174.510 355.300 ;
        RECT 176.340 355.140 176.510 355.310 ;
        RECT 177.720 355.730 177.890 355.900 ;
        RECT 177.720 355.370 177.890 355.540 ;
        RECT 233.380 356.920 233.550 357.090 ;
        RECT 207.670 356.520 207.840 356.690 ;
        RECT 231.800 356.690 231.970 356.860 ;
        RECT 212.980 356.430 213.150 356.600 ;
        RECT 236.780 356.860 236.950 357.030 ;
        RECT 229.170 356.430 229.340 356.600 ;
        RECT 234.480 356.520 234.650 356.690 ;
        RECT 237.720 356.470 237.890 356.640 ;
        RECT 239.030 356.880 239.200 357.050 ;
        RECT 212.980 355.980 213.150 356.150 ;
        RECT 214.960 356.000 215.130 356.170 ;
        RECT 229.170 355.980 229.340 356.150 ;
        RECT 233.880 356.000 234.050 356.170 ;
        RECT 201.380 355.080 201.550 355.250 ;
        RECT 167.080 354.510 167.250 354.680 ;
        RECT 169.510 354.610 169.680 354.780 ;
        RECT 170.550 354.570 170.720 354.740 ;
        RECT 203.190 354.780 203.370 354.950 ;
        RECT 234.360 355.940 234.530 356.110 ;
        RECT 236.730 356.210 236.900 356.380 ;
        RECT 232.530 355.410 232.700 355.580 ;
        RECT 234.820 355.320 234.990 355.490 ;
        RECT 238.380 355.500 238.550 355.670 ;
        RECT 236.730 355.070 236.900 355.240 ;
        RECT 240.410 355.900 240.590 356.090 ;
        RECT 240.770 355.080 240.940 355.250 ;
        RECT 232.920 354.680 233.090 354.850 ;
        RECT 237.720 354.810 237.890 354.980 ;
        RECT 236.780 354.420 236.950 354.590 ;
        RECT 238.950 354.830 239.130 354.950 ;
        RECT 238.950 354.780 239.250 354.830 ;
        RECT 239.080 354.660 239.250 354.780 ;
        RECT 168.550 354.100 168.760 354.310 ;
        RECT 218.180 354.160 218.350 354.330 ;
        RECT 218.190 353.440 218.360 353.610 ;
        RECT 223.970 354.160 224.140 354.330 ;
        RECT 236.780 353.860 236.950 354.030 ;
        RECT 239.070 353.940 239.240 354.110 ;
        RECT 223.970 353.440 224.140 353.610 ;
        RECT 187.290 352.000 187.560 352.270 ;
        RECT 191.320 352.070 191.590 352.340 ;
        RECT 221.370 352.070 221.640 352.340 ;
        RECT 232.480 352.310 232.650 352.480 ;
        RECT 225.400 352.000 225.670 352.270 ;
        RECT 232.630 351.480 232.800 351.650 ;
        RECT 237.720 353.470 237.890 353.640 ;
        RECT 236.730 353.210 236.900 353.380 ;
        RECT 238.380 352.910 238.550 353.080 ;
        RECT 236.730 352.070 236.900 352.240 ;
        RECT 237.720 351.810 237.890 351.980 ;
        RECT 236.780 351.420 236.950 351.590 ;
        RECT 238.990 351.690 239.160 351.860 ;
        RECT 171.590 350.390 171.760 350.560 ;
        RECT 171.590 350.030 171.760 350.200 ;
        RECT 172.730 350.300 172.900 350.470 ;
        RECT 173.570 350.180 173.740 350.350 ;
        RECT 174.320 350.180 174.490 350.350 ;
        RECT 167.080 349.630 167.250 349.800 ;
        RECT 169.510 349.730 169.680 349.900 ;
        RECT 170.550 349.690 170.720 349.860 ;
        RECT 177.300 349.850 177.470 350.020 ;
        RECT 168.550 349.220 168.760 349.430 ;
        RECT 172.910 349.470 173.080 349.640 ;
        RECT 177.700 350.300 177.870 350.470 ;
        RECT 198.510 350.530 198.680 350.700 ;
        RECT 214.280 350.530 214.450 350.700 ;
        RECT 177.700 349.940 177.870 350.110 ;
        RECT 231.790 350.660 231.960 350.830 ;
        RECT 196.840 350.120 197.010 350.290 ;
        RECT 197.570 350.090 197.740 350.260 ;
        RECT 198.510 349.980 198.680 350.150 ;
        RECT 214.280 349.980 214.450 350.150 ;
        RECT 215.220 350.090 215.390 350.260 ;
        RECT 215.950 350.120 216.120 350.290 ;
        RECT 199.560 349.430 199.730 349.600 ;
        RECT 171.590 348.640 171.760 348.810 ;
        RECT 171.590 348.280 171.760 348.450 ;
        RECT 172.910 348.570 173.080 348.740 ;
        RECT 177.300 348.190 177.470 348.360 ;
        RECT 167.080 347.880 167.250 348.050 ;
        RECT 169.510 347.980 169.680 348.150 ;
        RECT 170.550 347.940 170.720 348.110 ;
        RECT 173.570 347.860 173.740 348.030 ;
        RECT 174.320 347.860 174.490 348.030 ;
        RECT 176.320 347.870 176.490 348.040 ;
        RECT 177.700 348.460 177.870 348.630 ;
        RECT 196.840 348.560 197.010 348.730 ;
        RECT 203.500 349.440 203.670 349.610 ;
        RECT 209.290 349.440 209.460 349.610 ;
        RECT 213.230 349.430 213.400 349.600 ;
        RECT 197.570 348.590 197.740 348.760 ;
        RECT 198.510 348.700 198.680 348.870 ;
        RECT 214.280 348.700 214.450 348.870 ;
        RECT 215.220 348.590 215.390 348.760 ;
        RECT 232.520 349.380 232.690 349.550 ;
        RECT 215.950 348.560 216.120 348.730 ;
        RECT 232.910 348.650 233.080 348.820 ;
        RECT 177.700 348.100 177.870 348.270 ;
        RECT 198.510 348.150 198.680 348.320 ;
        RECT 199.560 347.840 199.730 348.010 ;
        RECT 168.550 347.470 168.760 347.680 ;
        RECT 4.770 346.410 6.680 346.590 ;
        RECT 172.730 347.100 172.900 347.270 ;
        RECT 171.590 346.890 171.760 347.060 ;
        RECT 173.570 346.980 173.740 347.150 ;
        RECT 174.320 346.980 174.490 347.150 ;
        RECT 171.590 346.530 171.760 346.700 ;
        RECT 177.300 346.650 177.470 346.820 ;
        RECT 4.770 346.010 6.670 346.190 ;
        RECT 167.080 346.130 167.250 346.300 ;
        RECT 169.510 346.230 169.680 346.400 ;
        RECT 170.550 346.190 170.720 346.360 ;
        RECT 172.910 346.270 173.080 346.440 ;
        RECT 177.700 347.100 177.870 347.270 ;
        RECT 177.700 346.740 177.870 346.910 ;
        RECT 185.250 346.980 185.520 347.250 ;
        RECT 189.280 347.050 189.550 347.320 ;
        RECT 198.510 347.290 198.680 347.460 ;
        RECT 199.560 347.480 199.730 347.650 ;
        RECT 203.490 347.980 203.660 348.150 ;
        RECT 203.490 347.620 203.660 347.790 ;
        RECT 209.300 347.980 209.470 348.150 ;
        RECT 209.300 347.620 209.470 347.790 ;
        RECT 214.280 348.150 214.450 348.320 ;
        RECT 213.230 347.840 213.400 348.010 ;
        RECT 215.590 347.720 215.770 347.890 ;
        RECT 213.230 347.480 213.400 347.650 ;
        RECT 214.280 347.290 214.450 347.460 ;
        RECT 196.840 346.880 197.010 347.050 ;
        RECT 197.570 346.850 197.740 347.020 ;
        RECT 198.510 346.740 198.680 346.910 ;
        RECT 214.280 346.740 214.450 346.910 ;
        RECT 215.220 346.850 215.390 347.020 ;
        RECT 215.950 346.880 216.120 347.050 ;
        RECT 168.550 345.720 168.760 345.930 ;
        RECT 171.590 345.140 171.760 345.310 ;
        RECT 172.910 345.370 173.080 345.540 ;
        RECT 177.300 344.990 177.470 345.160 ;
        RECT 171.590 344.780 171.760 344.950 ;
        RECT 4.640 344.310 5.570 344.510 ;
        RECT 167.080 344.380 167.250 344.550 ;
        RECT 169.510 344.480 169.680 344.650 ;
        RECT 170.550 344.440 170.720 344.610 ;
        RECT 173.570 344.660 173.740 344.830 ;
        RECT 174.320 344.660 174.490 344.830 ;
        RECT 176.320 344.670 176.490 344.840 ;
        RECT 177.700 345.260 177.870 345.430 ;
        RECT 196.470 345.550 196.640 345.720 ;
        RECT 177.700 344.900 177.870 345.070 ;
        RECT 196.840 345.330 197.010 345.500 ;
        RECT 197.570 345.360 197.740 345.530 ;
        RECT 198.510 345.470 198.680 345.640 ;
        RECT 214.280 345.470 214.450 345.640 ;
        RECT 194.800 345.140 194.970 345.310 ;
        RECT 215.220 345.360 215.390 345.530 ;
        RECT 215.950 345.330 216.120 345.500 ;
        RECT 195.530 345.110 195.700 345.280 ;
        RECT 196.470 345.000 196.640 345.170 ;
        RECT 198.510 344.920 198.680 345.090 ;
        RECT 214.280 344.920 214.450 345.090 ;
        RECT 4.410 340.740 4.590 343.900 ;
        RECT 7.510 343.240 10.810 343.590 ;
        RECT 2.570 331.200 2.740 331.370 ;
        RECT 2.930 331.200 3.100 331.370 ;
        RECT 3.290 331.200 3.460 331.370 ;
        RECT 3.650 331.200 3.820 331.370 ;
        RECT 6.300 332.740 6.470 342.190 ;
        RECT 7.050 332.730 7.220 342.120 ;
        RECT 7.770 332.760 7.940 342.160 ;
        RECT 8.430 332.770 8.600 342.140 ;
        RECT 9.080 332.760 9.250 342.210 ;
        RECT 9.720 332.770 9.890 342.160 ;
        RECT 197.650 344.390 197.820 344.560 ;
        RECT 168.550 343.970 168.760 344.180 ;
        RECT 194.800 343.600 194.970 343.770 ;
        RECT 201.670 344.420 201.840 344.590 ;
        RECT 195.530 343.630 195.700 343.800 ;
        RECT 196.470 343.740 196.640 343.910 ;
        RECT 196.470 343.190 196.640 343.360 ;
        RECT 197.640 343.190 197.810 343.360 ;
        RECT 197.640 342.530 197.810 342.700 ;
        RECT 196.470 342.310 196.640 342.480 ;
        RECT 201.660 343.130 201.830 343.300 ;
        RECT 201.660 342.490 201.830 342.660 ;
        RECT 194.800 341.900 194.970 342.070 ;
        RECT 171.550 341.330 171.720 341.500 ;
        RECT 195.530 341.870 195.700 342.040 ;
        RECT 196.470 341.760 196.640 341.930 ;
        RECT 171.550 340.970 171.720 341.140 ;
        RECT 172.760 341.030 172.930 341.200 ;
        RECT 167.040 340.570 167.210 340.740 ;
        RECT 169.470 340.670 169.640 340.840 ;
        RECT 170.510 340.630 170.680 340.800 ;
        RECT 173.600 340.910 173.770 341.080 ;
        RECT 174.350 340.910 174.520 341.080 ;
        RECT 145.430 340.060 145.600 340.230 ;
        RECT 146.080 340.060 146.250 340.230 ;
        RECT 168.510 340.160 168.720 340.370 ;
        RECT 177.330 340.580 177.500 340.750 ;
        RECT 172.940 340.200 173.110 340.370 ;
        RECT 177.730 341.030 177.900 341.200 ;
        RECT 208.070 340.960 208.240 341.130 ;
        RECT 177.730 340.670 177.900 340.840 ;
        RECT 194.800 340.350 194.970 340.520 ;
        RECT 195.530 340.380 195.700 340.550 ;
        RECT 196.470 340.490 196.640 340.660 ;
        RECT 210.230 340.550 210.400 340.720 ;
        RECT 144.210 339.620 144.380 339.790 ;
        RECT 144.910 339.620 145.080 339.790 ;
        RECT 208.220 340.280 208.390 340.450 ;
        RECT 196.470 339.940 196.640 340.110 ;
        RECT 208.970 339.980 209.140 340.150 ;
        RECT 171.550 339.580 171.720 339.750 ;
        RECT 208.220 339.680 208.390 339.850 ;
        RECT 146.450 339.390 146.620 339.560 ;
        RECT 171.550 339.220 171.720 339.390 ;
        RECT 167.040 338.820 167.210 338.990 ;
        RECT 169.470 338.920 169.640 339.090 ;
        RECT 170.510 338.880 170.680 339.050 ;
        RECT 172.940 339.300 173.110 339.470 ;
        RECT 177.330 338.920 177.500 339.090 ;
        RECT 168.510 338.410 168.720 338.620 ;
        RECT 173.600 338.590 173.770 338.760 ;
        RECT 174.350 338.590 174.520 338.760 ;
        RECT 176.350 338.600 176.520 338.770 ;
        RECT 177.730 339.190 177.900 339.360 ;
        RECT 210.230 339.410 210.400 339.580 ;
        RECT 177.730 338.830 177.900 339.000 ;
        RECT 208.070 339.000 208.240 339.170 ;
        RECT 208.070 338.190 208.240 338.360 ;
        RECT 143.530 337.850 143.700 338.020 ;
        RECT 146.620 337.910 146.790 338.080 ;
        RECT 171.550 337.830 171.720 338.000 ;
        RECT 142.000 335.510 142.170 335.680 ;
        RECT 138.690 335.070 138.860 335.240 ;
        RECT 139.790 335.080 139.960 335.250 ;
        RECT 140.880 335.080 141.050 335.250 ;
        RECT 144.240 335.740 144.410 335.910 ;
        RECT 144.930 335.730 145.100 335.900 ;
        RECT 142.010 335.040 142.180 335.210 ;
        RECT 139.240 334.400 139.410 334.570 ;
        RECT 139.240 333.030 139.410 333.200 ;
        RECT 145.410 334.960 145.580 335.130 ;
        RECT 146.630 337.370 146.800 337.540 ;
        RECT 171.550 337.470 171.720 337.640 ;
        RECT 172.760 337.830 172.930 338.000 ;
        RECT 173.600 337.710 173.770 337.880 ;
        RECT 174.350 337.710 174.520 337.880 ;
        RECT 167.040 337.070 167.210 337.240 ;
        RECT 169.470 337.170 169.640 337.340 ;
        RECT 170.510 337.130 170.680 337.300 ;
        RECT 177.330 337.380 177.500 337.550 ;
        RECT 168.510 336.660 168.720 336.870 ;
        RECT 172.940 337.000 173.110 337.170 ;
        RECT 177.730 337.830 177.900 338.000 ;
        RECT 210.230 337.780 210.400 337.950 ;
        RECT 177.730 337.470 177.900 337.640 ;
        RECT 208.220 337.510 208.390 337.680 ;
        RECT 208.970 337.210 209.140 337.380 ;
        RECT 196.630 336.850 196.800 337.020 ;
        RECT 208.220 336.910 208.390 337.080 ;
        RECT 146.440 336.410 146.610 336.580 ;
        RECT 171.550 336.080 171.720 336.250 ;
        RECT 172.940 336.100 173.110 336.270 ;
        RECT 171.550 335.720 171.720 335.890 ;
        RECT 177.330 335.720 177.500 335.890 ;
        RECT 167.040 335.320 167.210 335.490 ;
        RECT 169.470 335.420 169.640 335.590 ;
        RECT 170.510 335.380 170.680 335.550 ;
        RECT 173.600 335.390 173.770 335.560 ;
        RECT 174.350 335.390 174.520 335.560 ;
        RECT 176.350 335.400 176.520 335.570 ;
        RECT 177.730 335.990 177.900 336.160 ;
        RECT 210.230 336.640 210.400 336.810 ;
        RECT 208.070 336.230 208.240 336.400 ;
        RECT 196.680 335.890 196.850 336.060 ;
        RECT 177.730 335.630 177.900 335.800 ;
        RECT 146.120 334.900 146.290 335.070 ;
        RECT 168.510 334.910 168.720 335.120 ;
        RECT 140.340 334.400 140.510 334.570 ;
        RECT 141.440 334.400 141.610 334.570 ;
        RECT 142.270 334.530 142.440 334.700 ;
        RECT 142.270 333.840 142.440 334.010 ;
        RECT 172.560 333.280 172.730 333.450 ;
        RECT 140.340 333.030 140.510 333.200 ;
        RECT 141.440 333.030 141.610 333.200 ;
        RECT 2.890 324.520 3.060 324.690 ;
        RECT 3.250 324.520 3.420 324.690 ;
        RECT 3.620 324.520 3.790 324.690 ;
        RECT 4.410 319.240 4.580 319.250 ;
        RECT 4.400 317.380 4.580 319.240 ;
        RECT 5.540 319.010 5.710 329.990 ;
        RECT 6.160 319.010 6.330 329.990 ;
        RECT 6.780 319.020 6.950 330.000 ;
        RECT 7.360 319.040 7.530 330.020 ;
        RECT 7.950 319.050 8.120 330.030 ;
        RECT 8.550 319.050 8.720 330.030 ;
        RECT 9.150 319.000 9.320 329.980 ;
        RECT 9.760 319.010 9.930 329.990 ;
        RECT 10.360 319.000 10.530 329.980 ;
        RECT 138.690 332.300 138.860 332.470 ;
        RECT 138.680 330.960 138.850 331.130 ;
        RECT 139.790 332.300 139.960 332.470 ;
        RECT 140.880 332.300 141.050 332.470 ;
        RECT 148.820 331.280 148.990 331.620 ;
        RECT 149.190 331.280 149.360 331.620 ;
        RECT 139.790 330.950 139.960 331.120 ;
        RECT 140.880 330.930 141.050 331.100 ;
        RECT 139.240 330.260 139.410 330.430 ;
        RECT 140.340 330.250 140.510 330.420 ;
        RECT 141.430 330.250 141.600 330.420 ;
        RECT 173.650 333.280 173.820 333.450 ;
        RECT 173.110 332.600 173.280 332.770 ;
        RECT 173.110 331.230 173.280 331.400 ;
        RECT 172.550 330.500 172.720 330.670 ;
        RECT 172.550 329.130 172.720 329.300 ;
        RECT 171.980 328.490 172.150 328.660 ;
        RECT 171.990 328.020 172.160 328.190 ;
        RECT 174.750 333.270 174.920 333.440 ;
        RECT 174.200 332.580 174.370 332.750 ;
        RECT 174.200 331.230 174.370 331.400 ;
        RECT 173.650 330.500 173.820 330.670 ;
        RECT 173.650 329.130 173.820 329.300 ;
        RECT 173.110 328.450 173.280 328.620 ;
        RECT 175.730 333.300 175.900 333.470 ;
        RECT 175.730 332.940 175.900 333.110 ;
        RECT 175.310 332.570 175.480 332.740 ;
        RECT 176.340 333.300 176.510 333.470 ;
        RECT 176.340 332.940 176.510 333.110 ;
        RECT 177.320 333.270 177.490 333.440 ;
        RECT 176.760 332.570 176.930 332.740 ;
        RECT 175.300 331.230 175.470 331.400 ;
        RECT 176.770 331.230 176.940 331.400 ;
        RECT 174.750 330.500 174.920 330.670 ;
        RECT 174.750 329.130 174.920 329.300 ;
        RECT 174.200 328.450 174.370 328.620 ;
        RECT 178.420 333.280 178.590 333.450 ;
        RECT 177.870 332.580 178.040 332.750 ;
        RECT 177.870 331.230 178.040 331.400 ;
        RECT 177.320 330.500 177.490 330.670 ;
        RECT 177.320 329.130 177.490 329.300 ;
        RECT 175.300 328.460 175.470 328.630 ;
        RECT 176.770 328.460 176.940 328.630 ;
        RECT 179.510 333.280 179.680 333.450 ;
        RECT 178.960 332.600 179.130 332.770 ;
        RECT 178.960 331.230 179.130 331.400 ;
        RECT 178.420 330.500 178.590 330.670 ;
        RECT 178.420 329.130 178.590 329.300 ;
        RECT 177.870 328.450 178.040 328.620 ;
        RECT 179.520 330.500 179.690 330.670 ;
        RECT 179.520 329.130 179.690 329.300 ;
        RECT 178.960 328.450 179.130 328.620 ;
        RECT 182.370 333.310 182.540 333.480 ;
        RECT 183.460 333.310 183.630 333.480 ;
        RECT 182.920 332.630 183.090 332.800 ;
        RECT 182.920 331.260 183.090 331.430 ;
        RECT 182.360 330.530 182.530 330.700 ;
        RECT 182.360 329.160 182.530 329.330 ;
        RECT 180.090 328.490 180.260 328.660 ;
        RECT 181.790 328.520 181.960 328.690 ;
        RECT 180.080 328.020 180.250 328.190 ;
        RECT 181.800 328.050 181.970 328.220 ;
        RECT 184.560 333.300 184.730 333.470 ;
        RECT 184.010 332.610 184.180 332.780 ;
        RECT 184.010 331.260 184.180 331.430 ;
        RECT 183.460 330.530 183.630 330.700 ;
        RECT 183.460 329.160 183.630 329.330 ;
        RECT 182.920 328.480 183.090 328.650 ;
        RECT 185.540 333.330 185.710 333.500 ;
        RECT 185.540 332.970 185.710 333.140 ;
        RECT 185.120 332.600 185.290 332.770 ;
        RECT 186.150 333.330 186.320 333.500 ;
        RECT 186.150 332.970 186.320 333.140 ;
        RECT 187.130 333.300 187.300 333.470 ;
        RECT 186.570 332.600 186.740 332.770 ;
        RECT 185.110 331.260 185.280 331.430 ;
        RECT 186.580 331.260 186.750 331.430 ;
        RECT 184.560 330.530 184.730 330.700 ;
        RECT 184.560 329.160 184.730 329.330 ;
        RECT 184.010 328.480 184.180 328.650 ;
        RECT 188.230 333.310 188.400 333.480 ;
        RECT 187.680 332.610 187.850 332.780 ;
        RECT 187.680 331.260 187.850 331.430 ;
        RECT 187.130 330.530 187.300 330.700 ;
        RECT 187.130 329.160 187.300 329.330 ;
        RECT 185.110 328.490 185.280 328.660 ;
        RECT 186.580 328.490 186.750 328.660 ;
        RECT 189.320 333.310 189.490 333.480 ;
        RECT 188.770 332.630 188.940 332.800 ;
        RECT 188.770 331.260 188.940 331.430 ;
        RECT 188.230 330.530 188.400 330.700 ;
        RECT 188.230 329.160 188.400 329.330 ;
        RECT 187.680 328.480 187.850 328.650 ;
        RECT 189.330 330.530 189.500 330.700 ;
        RECT 189.330 329.160 189.500 329.330 ;
        RECT 188.770 328.480 188.940 328.650 ;
        RECT 189.900 328.520 190.070 328.690 ;
        RECT 189.890 328.050 190.060 328.220 ;
        RECT 193.510 329.090 193.680 329.260 ;
        RECT 192.950 328.390 193.120 328.560 ;
        RECT 192.960 327.050 193.130 327.220 ;
        RECT 194.610 329.100 194.780 329.270 ;
        RECT 195.700 329.100 195.870 329.270 ;
        RECT 194.060 328.400 194.230 328.570 ;
        RECT 195.150 328.420 195.320 328.590 ;
        RECT 194.060 327.050 194.230 327.220 ;
        RECT 195.150 327.050 195.320 327.220 ;
        RECT 193.510 326.320 193.680 326.490 ;
        RECT 193.510 324.950 193.680 325.120 ;
        RECT 192.960 324.280 193.130 324.450 ;
        RECT 194.610 326.320 194.780 326.490 ;
        RECT 195.710 326.320 195.880 326.490 ;
        RECT 196.540 325.870 196.710 326.040 ;
        RECT 196.540 325.510 196.710 325.680 ;
        RECT 194.610 324.950 194.780 325.120 ;
        RECT 195.710 324.950 195.880 325.120 ;
        RECT 227.100 325.460 227.270 325.630 ;
        RECT 232.690 324.760 232.860 324.930 ;
        RECT 194.060 324.270 194.230 324.440 ;
        RECT 195.150 324.270 195.320 324.440 ;
        RECT 196.280 324.310 196.450 324.480 ;
        RECT 232.690 324.090 232.860 324.260 ;
        RECT 138.090 323.320 138.260 323.490 ;
        RECT 139.190 323.330 139.360 323.500 ;
        RECT 138.640 322.650 138.810 322.820 ;
        RECT 138.640 321.280 138.810 321.450 ;
        RECT 138.090 320.550 138.260 320.720 ;
        RECT 138.080 319.210 138.250 319.380 ;
        RECT 137.660 318.840 137.830 319.010 ;
        RECT 4.770 317.820 6.680 318.000 ;
        RECT 140.280 323.330 140.450 323.500 ;
        RECT 139.740 322.650 139.910 322.820 ;
        RECT 139.740 321.280 139.910 321.450 ;
        RECT 139.190 320.550 139.360 320.720 ;
        RECT 139.190 319.200 139.360 319.370 ;
        RECT 138.640 318.510 138.810 318.680 ;
        RECT 141.400 323.760 141.570 323.930 ;
        RECT 196.270 323.840 196.440 324.010 ;
        RECT 227.100 323.850 227.270 324.020 ;
        RECT 141.410 323.290 141.580 323.460 ;
        RECT 140.840 322.650 141.010 322.820 ;
        RECT 140.840 321.280 141.010 321.450 ;
        RECT 140.280 320.550 140.450 320.720 ;
        RECT 140.280 319.180 140.450 319.350 ;
        RECT 139.740 318.500 139.910 318.670 ;
        RECT 143.010 319.310 143.180 322.830 ;
        RECT 143.370 319.310 143.540 322.830 ;
        RECT 143.730 319.310 143.900 322.830 ;
        RECT 144.420 319.310 144.590 322.830 ;
        RECT 144.780 319.310 144.950 322.830 ;
        RECT 145.140 319.310 145.310 322.830 ;
        RECT 227.100 322.250 227.270 322.420 ;
        RECT 227.100 320.630 227.270 320.800 ;
        RECT 231.030 319.240 231.200 319.410 ;
        RECT 227.100 319.030 227.270 319.200 ;
        RECT 140.830 318.500 141.000 318.670 ;
        RECT 4.770 317.420 6.670 317.600 ;
        RECT 227.100 317.410 227.270 317.580 ;
        RECT 4.640 315.720 5.570 315.920 ;
        RECT 227.100 315.810 227.270 315.980 ;
        RECT 4.410 312.150 4.590 315.310 ;
        RECT 7.510 314.650 10.810 315.000 ;
        RECT 2.570 302.610 2.740 302.780 ;
        RECT 2.930 302.610 3.100 302.780 ;
        RECT 3.290 302.610 3.460 302.780 ;
        RECT 3.650 302.610 3.820 302.780 ;
        RECT 6.300 304.150 6.470 313.600 ;
        RECT 7.050 304.140 7.220 313.530 ;
        RECT 7.770 304.170 7.940 313.570 ;
        RECT 8.430 304.180 8.600 313.550 ;
        RECT 9.080 304.170 9.250 313.620 ;
        RECT 9.720 304.180 9.890 313.570 ;
        RECT 227.100 314.190 227.270 314.360 ;
        RECT 233.380 312.100 233.550 327.050 ;
        RECT 2.890 295.930 3.060 296.100 ;
        RECT 3.250 295.930 3.420 296.100 ;
        RECT 3.620 295.930 3.790 296.100 ;
        RECT 4.410 290.650 4.580 290.660 ;
        RECT 4.400 288.790 4.580 290.650 ;
        RECT 5.540 290.420 5.710 301.400 ;
        RECT 6.160 290.420 6.330 301.400 ;
        RECT 6.780 290.430 6.950 301.410 ;
        RECT 7.360 290.450 7.530 301.430 ;
        RECT 7.950 290.460 8.120 301.440 ;
        RECT 8.550 290.460 8.720 301.440 ;
        RECT 9.150 290.410 9.320 301.390 ;
        RECT 9.760 290.420 9.930 301.400 ;
        RECT 10.360 290.410 10.530 301.390 ;
        RECT 4.770 289.230 6.680 289.410 ;
        RECT 4.770 288.830 6.670 289.010 ;
        RECT 4.640 287.130 5.570 287.330 ;
        RECT 4.410 283.560 4.590 286.720 ;
        RECT 7.510 286.060 10.810 286.410 ;
        RECT 2.570 274.020 2.740 274.190 ;
        RECT 2.930 274.020 3.100 274.190 ;
        RECT 3.290 274.020 3.460 274.190 ;
        RECT 3.650 274.020 3.820 274.190 ;
        RECT 6.300 275.560 6.470 285.010 ;
        RECT 7.050 275.550 7.220 284.940 ;
        RECT 7.770 275.580 7.940 284.980 ;
        RECT 8.430 275.590 8.600 284.960 ;
        RECT 9.080 275.580 9.250 285.030 ;
        RECT 9.720 275.590 9.890 284.980 ;
        RECT 2.890 267.340 3.060 267.510 ;
        RECT 3.250 267.340 3.420 267.510 ;
        RECT 3.620 267.340 3.790 267.510 ;
        RECT 4.410 262.060 4.580 262.070 ;
        RECT 4.400 260.200 4.580 262.060 ;
        RECT 5.540 261.830 5.710 272.810 ;
        RECT 6.160 261.830 6.330 272.810 ;
        RECT 6.780 261.840 6.950 272.820 ;
        RECT 7.360 261.860 7.530 272.840 ;
        RECT 7.950 261.870 8.120 272.850 ;
        RECT 8.550 261.870 8.720 272.850 ;
        RECT 9.150 261.820 9.320 272.800 ;
        RECT 9.760 261.830 9.930 272.810 ;
        RECT 10.360 261.820 10.530 272.800 ;
        RECT 4.770 260.640 6.680 260.820 ;
        RECT 4.770 260.240 6.670 260.420 ;
        RECT 4.640 258.540 5.570 258.740 ;
        RECT 4.410 254.970 4.590 258.130 ;
        RECT 7.510 257.470 10.810 257.820 ;
        RECT 2.570 245.430 2.740 245.600 ;
        RECT 2.930 245.430 3.100 245.600 ;
        RECT 3.290 245.430 3.460 245.600 ;
        RECT 3.650 245.430 3.820 245.600 ;
        RECT 6.300 246.970 6.470 256.420 ;
        RECT 7.050 246.960 7.220 256.350 ;
        RECT 7.770 246.990 7.940 256.390 ;
        RECT 8.430 247.000 8.600 256.370 ;
        RECT 9.080 246.990 9.250 256.440 ;
        RECT 9.720 247.000 9.890 256.390 ;
        RECT 2.890 238.750 3.060 238.920 ;
        RECT 3.250 238.750 3.420 238.920 ;
        RECT 3.620 238.750 3.790 238.920 ;
        RECT 4.410 233.470 4.580 233.480 ;
        RECT 4.400 231.610 4.580 233.470 ;
        RECT 5.540 233.240 5.710 244.220 ;
        RECT 6.160 233.240 6.330 244.220 ;
        RECT 6.780 233.250 6.950 244.230 ;
        RECT 7.360 233.270 7.530 244.250 ;
        RECT 7.950 233.280 8.120 244.260 ;
        RECT 8.550 233.280 8.720 244.260 ;
        RECT 9.150 233.230 9.320 244.210 ;
        RECT 9.760 233.240 9.930 244.220 ;
        RECT 10.360 233.230 10.530 244.210 ;
        RECT 4.770 232.050 6.680 232.230 ;
        RECT 4.770 231.650 6.670 231.830 ;
        RECT 4.640 229.950 5.570 230.150 ;
        RECT 4.410 226.380 4.590 229.540 ;
        RECT 7.510 228.880 10.810 229.230 ;
        RECT 2.570 216.840 2.740 217.010 ;
        RECT 2.930 216.840 3.100 217.010 ;
        RECT 3.290 216.840 3.460 217.010 ;
        RECT 3.650 216.840 3.820 217.010 ;
        RECT 6.300 218.380 6.470 227.830 ;
        RECT 7.050 218.370 7.220 227.760 ;
        RECT 7.770 218.400 7.940 227.800 ;
        RECT 8.430 218.410 8.600 227.780 ;
        RECT 9.080 218.400 9.250 227.850 ;
        RECT 9.720 218.410 9.890 227.800 ;
        RECT 2.890 210.160 3.060 210.330 ;
        RECT 3.250 210.160 3.420 210.330 ;
        RECT 3.620 210.160 3.790 210.330 ;
        RECT 4.410 204.880 4.580 204.890 ;
        RECT 4.400 203.020 4.580 204.880 ;
        RECT 5.540 204.650 5.710 215.630 ;
        RECT 6.160 204.650 6.330 215.630 ;
        RECT 6.780 204.660 6.950 215.640 ;
        RECT 7.360 204.680 7.530 215.660 ;
        RECT 7.950 204.690 8.120 215.670 ;
        RECT 8.550 204.690 8.720 215.670 ;
        RECT 9.150 204.640 9.320 215.620 ;
        RECT 9.760 204.650 9.930 215.630 ;
        RECT 10.360 204.640 10.530 215.620 ;
        RECT 4.770 203.460 6.680 203.640 ;
        RECT 4.770 203.060 6.670 203.240 ;
        RECT 4.640 201.360 5.570 201.560 ;
        RECT 4.410 197.790 4.590 200.950 ;
        RECT 7.510 200.290 10.810 200.640 ;
        RECT 2.570 188.250 2.740 188.420 ;
        RECT 2.930 188.250 3.100 188.420 ;
        RECT 3.290 188.250 3.460 188.420 ;
        RECT 3.650 188.250 3.820 188.420 ;
        RECT 6.300 189.790 6.470 199.240 ;
        RECT 7.050 189.780 7.220 199.170 ;
        RECT 7.770 189.810 7.940 199.210 ;
        RECT 8.430 189.820 8.600 199.190 ;
        RECT 9.080 189.810 9.250 199.260 ;
        RECT 9.720 189.820 9.890 199.210 ;
        RECT 2.890 181.570 3.060 181.740 ;
        RECT 3.250 181.570 3.420 181.740 ;
        RECT 3.620 181.570 3.790 181.740 ;
        RECT 4.410 176.290 4.580 176.300 ;
        RECT 4.400 174.430 4.580 176.290 ;
        RECT 5.540 176.060 5.710 187.040 ;
        RECT 6.160 176.060 6.330 187.040 ;
        RECT 6.780 176.070 6.950 187.050 ;
        RECT 7.360 176.090 7.530 187.070 ;
        RECT 7.950 176.100 8.120 187.080 ;
        RECT 8.550 176.100 8.720 187.080 ;
        RECT 9.150 176.050 9.320 187.030 ;
        RECT 9.760 176.060 9.930 187.040 ;
        RECT 10.360 176.050 10.530 187.030 ;
        RECT 4.770 174.870 6.680 175.050 ;
        RECT 4.770 174.470 6.670 174.650 ;
        RECT 4.640 172.770 5.570 172.970 ;
        RECT 4.410 169.200 4.590 172.360 ;
        RECT 7.510 171.700 10.810 172.050 ;
        RECT 2.570 159.660 2.740 159.830 ;
        RECT 2.930 159.660 3.100 159.830 ;
        RECT 3.290 159.660 3.460 159.830 ;
        RECT 3.650 159.660 3.820 159.830 ;
        RECT 6.300 161.200 6.470 170.650 ;
        RECT 7.050 161.190 7.220 170.580 ;
        RECT 7.770 161.220 7.940 170.620 ;
        RECT 8.430 161.230 8.600 170.600 ;
        RECT 9.080 161.220 9.250 170.670 ;
        RECT 9.720 161.230 9.890 170.620 ;
        RECT 2.890 152.980 3.060 153.150 ;
        RECT 3.250 152.980 3.420 153.150 ;
        RECT 3.620 152.980 3.790 153.150 ;
        RECT 4.410 147.700 4.580 147.710 ;
        RECT 4.400 145.840 4.580 147.700 ;
        RECT 5.540 147.470 5.710 158.450 ;
        RECT 6.160 147.470 6.330 158.450 ;
        RECT 6.780 147.480 6.950 158.460 ;
        RECT 7.360 147.500 7.530 158.480 ;
        RECT 7.950 147.510 8.120 158.490 ;
        RECT 8.550 147.510 8.720 158.490 ;
        RECT 9.150 147.460 9.320 158.440 ;
        RECT 9.760 147.470 9.930 158.450 ;
        RECT 10.360 147.460 10.530 158.440 ;
        RECT 4.770 146.280 6.680 146.460 ;
        RECT 4.770 145.880 6.670 146.060 ;
        RECT 4.640 144.180 5.570 144.380 ;
        RECT 4.410 140.610 4.590 143.770 ;
        RECT 7.510 143.110 10.810 143.460 ;
        RECT 2.570 131.070 2.740 131.240 ;
        RECT 2.930 131.070 3.100 131.240 ;
        RECT 3.290 131.070 3.460 131.240 ;
        RECT 3.650 131.070 3.820 131.240 ;
        RECT 6.300 132.610 6.470 142.060 ;
        RECT 7.050 132.600 7.220 141.990 ;
        RECT 7.770 132.630 7.940 142.030 ;
        RECT 8.430 132.640 8.600 142.010 ;
        RECT 9.080 132.630 9.250 142.080 ;
        RECT 9.720 132.640 9.890 142.030 ;
        RECT 2.890 124.390 3.060 124.560 ;
        RECT 3.250 124.390 3.420 124.560 ;
        RECT 3.620 124.390 3.790 124.560 ;
        RECT 4.410 119.110 4.580 119.120 ;
        RECT 4.400 117.250 4.580 119.110 ;
        RECT 5.540 118.880 5.710 129.860 ;
        RECT 6.160 118.880 6.330 129.860 ;
        RECT 6.780 118.890 6.950 129.870 ;
        RECT 7.360 118.910 7.530 129.890 ;
        RECT 7.950 118.920 8.120 129.900 ;
        RECT 8.550 118.920 8.720 129.900 ;
        RECT 9.150 118.870 9.320 129.850 ;
        RECT 9.760 118.880 9.930 129.860 ;
        RECT 10.360 118.870 10.530 129.850 ;
        RECT 4.770 117.690 6.680 117.870 ;
        RECT 4.770 117.290 6.670 117.470 ;
        RECT 4.640 115.590 5.570 115.790 ;
        RECT 4.410 112.020 4.590 115.180 ;
        RECT 7.510 114.520 10.810 114.870 ;
        RECT 2.570 102.480 2.740 102.650 ;
        RECT 2.930 102.480 3.100 102.650 ;
        RECT 3.290 102.480 3.460 102.650 ;
        RECT 3.650 102.480 3.820 102.650 ;
        RECT 6.300 104.020 6.470 113.470 ;
        RECT 7.050 104.010 7.220 113.400 ;
        RECT 7.770 104.040 7.940 113.440 ;
        RECT 8.430 104.050 8.600 113.420 ;
        RECT 9.080 104.040 9.250 113.490 ;
        RECT 9.720 104.050 9.890 113.440 ;
        RECT 2.890 95.800 3.060 95.970 ;
        RECT 3.250 95.800 3.420 95.970 ;
        RECT 3.620 95.800 3.790 95.970 ;
        RECT 4.410 90.520 4.580 90.530 ;
        RECT 4.400 88.660 4.580 90.520 ;
        RECT 5.540 90.290 5.710 101.270 ;
        RECT 6.160 90.290 6.330 101.270 ;
        RECT 6.780 90.300 6.950 101.280 ;
        RECT 7.360 90.320 7.530 101.300 ;
        RECT 7.950 90.330 8.120 101.310 ;
        RECT 8.550 90.330 8.720 101.310 ;
        RECT 9.150 90.280 9.320 101.260 ;
        RECT 9.760 90.290 9.930 101.270 ;
        RECT 10.360 90.280 10.530 101.260 ;
        RECT 4.770 89.100 6.680 89.280 ;
        RECT 4.770 88.700 6.670 88.880 ;
        RECT 4.640 87.000 5.570 87.200 ;
        RECT 4.410 83.430 4.590 86.590 ;
        RECT 7.510 85.930 10.810 86.280 ;
        RECT 2.570 73.890 2.740 74.060 ;
        RECT 2.930 73.890 3.100 74.060 ;
        RECT 3.290 73.890 3.460 74.060 ;
        RECT 3.650 73.890 3.820 74.060 ;
        RECT 6.300 75.430 6.470 84.880 ;
        RECT 7.050 75.420 7.220 84.810 ;
        RECT 7.770 75.450 7.940 84.850 ;
        RECT 8.430 75.460 8.600 84.830 ;
        RECT 9.080 75.450 9.250 84.900 ;
        RECT 9.720 75.460 9.890 84.850 ;
        RECT 2.890 67.210 3.060 67.380 ;
        RECT 3.250 67.210 3.420 67.380 ;
        RECT 3.620 67.210 3.790 67.380 ;
        RECT 4.410 61.930 4.580 61.940 ;
        RECT 4.400 60.070 4.580 61.930 ;
        RECT 5.540 61.700 5.710 72.680 ;
        RECT 6.160 61.700 6.330 72.680 ;
        RECT 6.780 61.710 6.950 72.690 ;
        RECT 7.360 61.730 7.530 72.710 ;
        RECT 7.950 61.740 8.120 72.720 ;
        RECT 8.550 61.740 8.720 72.720 ;
        RECT 9.150 61.690 9.320 72.670 ;
        RECT 9.760 61.700 9.930 72.680 ;
        RECT 10.360 61.690 10.530 72.670 ;
        RECT 4.770 60.510 6.680 60.690 ;
        RECT 4.770 60.110 6.670 60.290 ;
        RECT 4.640 58.410 5.570 58.610 ;
        RECT 4.410 54.840 4.590 58.000 ;
        RECT 7.510 57.340 10.810 57.690 ;
        RECT 2.570 45.300 2.740 45.470 ;
        RECT 2.930 45.300 3.100 45.470 ;
        RECT 3.290 45.300 3.460 45.470 ;
        RECT 3.650 45.300 3.820 45.470 ;
        RECT 6.300 46.840 6.470 56.290 ;
        RECT 7.050 46.830 7.220 56.220 ;
        RECT 7.770 46.860 7.940 56.260 ;
        RECT 8.430 46.870 8.600 56.240 ;
        RECT 9.080 46.860 9.250 56.310 ;
        RECT 9.720 46.870 9.890 56.260 ;
        RECT 2.890 38.620 3.060 38.790 ;
        RECT 3.250 38.620 3.420 38.790 ;
        RECT 3.620 38.620 3.790 38.790 ;
        RECT 4.410 33.340 4.580 33.350 ;
        RECT 4.400 31.480 4.580 33.340 ;
        RECT 5.540 33.110 5.710 44.090 ;
        RECT 6.160 33.110 6.330 44.090 ;
        RECT 6.780 33.120 6.950 44.100 ;
        RECT 7.360 33.140 7.530 44.120 ;
        RECT 7.950 33.150 8.120 44.130 ;
        RECT 8.550 33.150 8.720 44.130 ;
        RECT 9.150 33.100 9.320 44.080 ;
        RECT 9.760 33.110 9.930 44.090 ;
        RECT 10.360 33.100 10.530 44.080 ;
        RECT 4.770 31.920 6.680 32.100 ;
        RECT 4.770 31.520 6.670 31.700 ;
        RECT 4.640 29.820 5.570 30.020 ;
        RECT 4.410 26.250 4.590 29.410 ;
        RECT 7.510 28.750 10.810 29.100 ;
        RECT 2.570 16.710 2.740 16.880 ;
        RECT 2.930 16.710 3.100 16.880 ;
        RECT 3.290 16.710 3.460 16.880 ;
        RECT 3.650 16.710 3.820 16.880 ;
        RECT 6.300 18.250 6.470 27.700 ;
        RECT 7.050 18.240 7.220 27.630 ;
        RECT 7.770 18.270 7.940 27.670 ;
        RECT 8.430 18.280 8.600 27.650 ;
        RECT 9.080 18.270 9.250 27.720 ;
        RECT 9.720 18.280 9.890 27.670 ;
        RECT 2.890 10.030 3.060 10.200 ;
        RECT 3.250 10.030 3.420 10.200 ;
        RECT 3.620 10.030 3.790 10.200 ;
        RECT 4.410 4.750 4.580 4.760 ;
        RECT 4.400 2.890 4.580 4.750 ;
        RECT 5.540 4.520 5.710 15.500 ;
        RECT 6.160 4.520 6.330 15.500 ;
        RECT 6.780 4.530 6.950 15.510 ;
        RECT 7.360 4.550 7.530 15.530 ;
        RECT 7.950 4.560 8.120 15.540 ;
        RECT 8.550 4.560 8.720 15.540 ;
        RECT 9.150 4.510 9.320 15.490 ;
        RECT 9.760 4.520 9.930 15.500 ;
        RECT 10.360 4.510 10.530 15.490 ;
        RECT 4.770 3.330 6.680 3.510 ;
        RECT 4.770 2.930 6.670 3.110 ;
      LAYER met1 ;
        RECT 164.820 388.670 168.710 389.080 ;
        RECT 150.210 387.820 152.620 388.460 ;
        RECT 30.280 387.250 30.630 387.410 ;
        RECT 58.870 387.250 59.220 387.410 ;
        RECT 87.460 387.250 87.810 387.410 ;
        RECT 30.270 386.300 30.640 387.250 ;
        RECT 58.860 386.300 59.230 387.250 ;
        RECT 87.450 386.300 87.820 387.250 ;
        RECT 150.230 386.470 150.640 387.820 ;
        RECT 156.960 387.160 157.370 387.930 ;
        RECT 164.820 387.910 168.730 388.670 ;
        RECT 156.690 386.890 157.370 387.160 ;
        RECT 164.840 387.870 168.730 387.910 ;
        RECT 164.840 387.280 168.740 387.870 ;
        RECT 156.690 386.460 158.380 386.890 ;
        RECT 29.920 385.930 32.390 386.300 ;
        RECT 58.510 385.930 60.980 386.300 ;
        RECT 87.100 385.930 89.570 386.300 ;
        RECT 129.480 386.280 153.850 386.300 ;
        RECT 16.370 385.130 18.740 385.760 ;
        RECT 16.400 383.170 17.350 385.130 ;
        RECT 18.100 385.110 18.680 385.130 ;
        RECT 28.480 384.470 32.390 385.930 ;
        RECT 39.710 385.280 43.840 385.680 ;
        RECT 39.710 385.190 43.850 385.280 ;
        RECT 18.770 384.460 32.390 384.470 ;
        RECT 16.630 377.500 17.350 383.170 ;
        RECT 18.100 383.900 32.390 384.460 ;
        RECT 43.320 384.290 43.850 385.190 ;
        RECT 44.960 385.130 47.330 385.760 ;
        RECT 18.100 379.600 41.450 383.900 ;
        RECT 44.990 383.170 45.940 385.130 ;
        RECT 46.690 385.110 47.270 385.130 ;
        RECT 57.070 384.470 60.980 385.930 ;
        RECT 68.300 385.280 72.430 385.680 ;
        RECT 68.300 385.190 72.440 385.280 ;
        RECT 47.360 384.460 60.980 384.470 ;
        RECT 42.220 382.480 42.790 382.490 ;
        RECT 18.100 379.320 32.390 379.600 ;
        RECT 28.480 377.770 32.390 379.320 ;
        RECT 42.220 379.060 42.840 382.480 ;
        RECT 42.220 379.050 42.790 379.060 ;
        RECT 28.460 376.230 32.410 377.770 ;
        RECT 41.390 377.420 41.950 377.920 ;
        RECT 45.220 377.500 45.940 383.170 ;
        RECT 46.690 383.900 60.980 384.460 ;
        RECT 71.910 384.290 72.440 385.190 ;
        RECT 73.550 385.130 75.920 385.760 ;
        RECT 46.690 379.600 70.040 383.900 ;
        RECT 73.580 383.170 74.530 385.130 ;
        RECT 75.280 385.110 75.860 385.130 ;
        RECT 85.660 384.470 89.570 385.930 ;
        RECT 129.420 385.890 153.850 386.280 ;
        RECT 96.890 385.280 101.020 385.680 ;
        RECT 96.890 385.190 101.030 385.280 ;
        RECT 75.950 384.460 89.570 384.470 ;
        RECT 70.810 382.480 71.380 382.490 ;
        RECT 46.690 379.320 60.980 379.600 ;
        RECT 57.070 377.770 60.980 379.320 ;
        RECT 70.810 379.060 71.430 382.480 ;
        RECT 70.810 379.050 71.380 379.060 ;
        RECT 41.400 377.200 41.950 377.420 ;
        RECT 57.050 377.000 61.000 377.770 ;
        RECT 69.980 377.420 70.540 377.920 ;
        RECT 73.810 377.500 74.530 383.170 ;
        RECT 75.280 383.900 89.570 384.460 ;
        RECT 100.500 384.290 101.030 385.190 ;
        RECT 75.280 379.600 98.630 383.900 ;
        RECT 99.400 382.480 99.970 382.490 ;
        RECT 75.280 379.320 89.570 379.600 ;
        RECT 85.660 377.770 89.570 379.320 ;
        RECT 99.400 379.060 100.020 382.480 ;
        RECT 126.760 379.640 127.260 380.120 ;
        RECT 119.440 379.260 119.680 379.620 ;
        RECT 99.400 379.050 99.970 379.060 ;
        RECT 69.990 377.200 70.540 377.420 ;
        RECT 57.060 376.230 61.010 377.000 ;
        RECT 85.640 376.230 89.590 377.770 ;
        RECT 98.570 377.420 99.130 377.920 ;
        RECT 98.580 377.200 99.130 377.420 ;
        RECT 98.860 376.490 99.030 376.610 ;
        RECT 4.650 373.250 5.640 373.260 ;
        RECT 4.250 372.730 5.640 373.250 ;
        RECT 4.250 369.120 4.740 372.730 ;
        RECT 7.450 372.200 10.870 372.250 ;
        RECT 7.440 371.630 10.880 372.200 ;
        RECT 6.030 361.800 10.330 370.860 ;
        RECT 12.010 370.810 12.730 371.360 ;
        RECT 12.010 370.800 12.510 370.810 ;
        RECT 29.140 365.590 32.370 376.230 ;
        RECT 57.730 369.000 60.960 376.230 ;
        RECT 86.320 373.290 89.550 376.230 ;
        RECT 85.890 370.550 89.720 373.290 ;
        RECT 98.510 369.930 99.030 376.490 ;
        RECT 98.450 369.420 99.100 369.930 ;
        RECT 57.570 366.110 61.070 369.000 ;
        RECT 26.970 361.970 32.370 365.590 ;
        RECT 14.530 361.890 17.920 361.960 ;
        RECT 12.160 361.810 12.930 361.820 ;
        RECT 13.560 361.810 17.920 361.890 ;
        RECT 12.160 361.800 17.920 361.810 ;
        RECT 3.630 360.050 17.920 361.800 ;
        RECT 26.970 361.790 29.910 361.970 ;
        RECT 98.510 361.740 99.030 369.420 ;
        RECT 101.910 365.510 102.320 376.720 ;
        RECT 126.860 376.680 127.250 379.640 ;
        RECT 129.420 377.640 129.830 385.890 ;
        RECT 156.020 385.760 158.380 386.460 ;
        RECT 164.840 386.300 165.130 387.280 ;
        RECT 171.480 387.250 171.830 387.410 ;
        RECT 200.070 387.250 200.420 387.410 ;
        RECT 228.660 387.250 229.010 387.410 ;
        RECT 257.250 387.250 257.600 387.410 ;
        RECT 285.840 387.250 286.190 387.410 ;
        RECT 314.430 387.250 314.780 387.410 ;
        RECT 343.020 387.250 343.370 387.410 ;
        RECT 171.470 386.300 171.840 387.250 ;
        RECT 200.060 386.300 200.430 387.250 ;
        RECT 228.650 386.300 229.020 387.250 ;
        RECT 257.240 386.300 257.610 387.250 ;
        RECT 285.830 386.300 286.200 387.250 ;
        RECT 314.420 386.300 314.790 387.250 ;
        RECT 343.010 386.300 343.380 387.250 ;
        RECT 162.650 386.290 184.010 386.300 ;
        RECT 162.590 385.900 184.010 386.290 ;
        RECT 199.710 385.930 202.180 386.300 ;
        RECT 228.300 385.930 230.770 386.300 ;
        RECT 256.890 385.930 259.360 386.300 ;
        RECT 285.480 385.930 287.950 386.300 ;
        RECT 314.070 385.930 316.540 386.300 ;
        RECT 342.660 385.930 345.130 386.300 ;
        RECT 162.590 385.890 183.850 385.900 ;
        RECT 156.020 385.130 159.940 385.760 ;
        RECT 152.860 380.480 154.200 380.930 ;
        RECT 156.020 380.480 158.550 385.130 ;
        RECT 159.300 385.110 159.880 385.130 ;
        RECT 169.680 384.470 173.590 385.890 ;
        RECT 180.910 385.280 185.040 385.680 ;
        RECT 180.910 385.190 185.050 385.280 ;
        RECT 159.970 384.460 173.590 384.470 ;
        RECT 159.300 383.900 173.590 384.460 ;
        RECT 184.520 384.290 185.050 385.190 ;
        RECT 186.160 385.130 188.530 385.760 ;
        RECT 159.300 380.480 182.650 383.900 ;
        RECT 186.190 383.170 187.140 385.130 ;
        RECT 187.890 385.110 188.470 385.130 ;
        RECT 198.270 384.470 202.180 385.930 ;
        RECT 209.500 385.280 213.630 385.680 ;
        RECT 209.500 385.190 213.640 385.280 ;
        RECT 188.560 384.460 202.180 384.470 ;
        RECT 152.860 380.060 182.650 380.480 ;
        RECT 138.830 379.180 139.090 379.970 ;
        RECT 152.860 379.920 154.200 380.060 ;
        RECT 147.450 379.320 150.220 379.560 ;
        RECT 147.450 378.910 147.690 379.320 ;
        RECT 120.020 376.270 120.280 376.570 ;
        RECT 122.880 376.430 123.140 376.620 ;
        RECT 122.880 376.300 123.250 376.430 ;
        RECT 120.020 376.250 120.430 376.270 ;
        RECT 120.050 375.960 120.430 376.250 ;
        RECT 121.460 375.960 122.490 376.270 ;
        RECT 122.960 376.200 123.250 376.300 ;
        RECT 120.010 375.400 120.270 375.540 ;
        RECT 120.010 375.220 120.360 375.400 ;
        RECT 120.650 375.240 120.970 375.560 ;
        RECT 121.420 375.400 121.680 375.550 ;
        RECT 121.420 375.230 121.760 375.400 ;
        RECT 120.120 375.170 120.360 375.220 ;
        RECT 121.530 375.170 121.760 375.230 ;
        RECT 120.060 375.090 121.810 375.170 ;
        RECT 120.010 374.770 121.810 375.090 ;
        RECT 120.060 374.670 121.810 374.770 ;
        RECT 120.010 374.510 121.810 374.670 ;
        RECT 120.010 374.350 120.360 374.510 ;
        RECT 120.650 374.400 120.970 374.510 ;
        RECT 121.440 374.370 121.760 374.510 ;
        RECT 120.120 374.290 120.360 374.350 ;
        RECT 121.530 374.290 121.760 374.370 ;
        RECT 120.120 373.320 120.350 373.740 ;
        RECT 120.010 373.000 120.350 373.320 ;
        RECT 120.120 372.330 120.350 373.000 ;
        RECT 121.530 372.330 121.760 373.740 ;
        RECT 122.250 373.560 122.490 375.960 ;
        RECT 126.860 376.190 127.330 376.680 ;
        RECT 128.410 376.230 130.890 377.000 ;
        RECT 126.860 376.180 127.310 376.190 ;
        RECT 122.970 375.510 123.240 375.640 ;
        RECT 122.650 375.280 123.330 375.510 ;
        RECT 122.910 375.220 123.330 375.280 ;
        RECT 122.630 374.660 122.950 374.980 ;
        RECT 122.680 374.430 122.910 374.660 ;
        RECT 123.100 374.280 123.330 375.220 ;
        RECT 122.970 374.100 123.330 374.280 ;
        RECT 122.970 374.080 123.240 374.100 ;
        RECT 122.650 373.850 123.240 374.080 ;
        RECT 122.160 373.270 122.490 373.560 ;
        RECT 122.250 373.190 122.490 373.270 ;
        RECT 122.350 372.500 122.670 372.820 ;
        RECT 122.970 372.810 123.240 373.850 ;
        RECT 122.970 372.580 123.300 372.810 ;
        RECT 120.630 371.600 120.950 371.920 ;
        RECT 122.060 371.620 122.380 371.940 ;
        RECT 119.840 371.020 120.160 371.340 ;
        RECT 120.770 371.020 121.090 371.340 ;
        RECT 121.470 371.020 121.790 371.340 ;
        RECT 122.210 371.020 122.530 371.340 ;
        RECT 122.920 371.010 123.240 371.330 ;
        RECT 124.960 370.620 125.250 371.680 ;
        RECT 101.790 365.040 102.320 365.510 ;
        RECT 98.310 361.010 99.030 361.740 ;
        RECT 2.680 360.040 17.920 360.050 ;
        RECT 2.520 359.690 17.920 360.040 ;
        RECT 2.680 359.680 17.920 359.690 ;
        RECT 3.630 359.330 17.920 359.680 ;
        RECT 4.000 357.890 17.920 359.330 ;
        RECT 5.460 348.180 10.610 357.890 ;
        RECT 12.160 357.870 13.560 357.890 ;
        RECT 4.170 348.090 4.800 348.150 ;
        RECT 4.170 347.510 4.820 348.090 ;
        RECT 5.470 347.510 10.610 348.180 ;
        RECT 4.170 346.760 4.800 347.510 ;
        RECT 4.170 346.040 12.430 346.760 ;
        RECT 4.170 345.810 6.760 346.040 ;
        RECT 4.170 345.780 4.800 345.810 ;
        RECT 4.650 344.660 5.640 344.670 ;
        RECT 4.250 344.140 5.640 344.660 ;
        RECT 4.250 340.530 4.740 344.140 ;
        RECT 7.450 343.610 10.870 343.660 ;
        RECT 7.440 343.040 10.880 343.610 ;
        RECT 6.030 333.210 10.330 342.270 ;
        RECT 12.010 342.220 12.730 342.770 ;
        RECT 12.010 342.210 12.510 342.220 ;
        RECT 12.160 333.210 13.560 333.230 ;
        RECT 23.700 333.210 25.960 333.250 ;
        RECT 3.630 331.460 25.960 333.210 ;
        RECT 2.680 331.450 25.960 331.460 ;
        RECT 2.520 331.100 25.960 331.450 ;
        RECT 2.680 331.090 25.960 331.100 ;
        RECT 3.630 330.740 25.960 331.090 ;
        RECT 4.000 329.980 25.960 330.740 ;
        RECT 4.000 329.300 13.560 329.980 ;
        RECT 23.700 329.940 25.960 329.980 ;
        RECT 5.460 319.590 10.610 329.300 ;
        RECT 12.160 329.290 13.560 329.300 ;
        RECT 12.160 329.280 12.930 329.290 ;
        RECT 98.510 325.660 99.030 361.010 ;
        RECT 101.910 360.790 102.320 365.040 ;
        RECT 101.770 360.200 102.390 360.790 ;
        RECT 98.430 325.060 99.060 325.660 ;
        RECT 101.910 324.640 102.320 360.200 ;
        RECT 101.860 324.140 102.340 324.640 ;
        RECT 4.170 319.500 4.800 319.560 ;
        RECT 4.170 318.920 4.820 319.500 ;
        RECT 5.470 318.920 10.610 319.590 ;
        RECT 4.170 318.170 4.800 318.920 ;
        RECT 4.170 317.450 12.430 318.170 ;
        RECT 126.860 318.070 127.250 376.180 ;
        RECT 128.270 375.040 128.530 375.360 ;
        RECT 128.280 372.820 128.520 375.040 ;
        RECT 129.020 374.720 130.180 376.230 ;
        RECT 133.120 376.180 133.360 376.820 ;
        RECT 138.330 376.260 138.570 376.670 ;
        RECT 133.120 375.920 133.350 376.180 ;
        RECT 133.110 375.700 133.350 375.920 ;
        RECT 144.170 375.420 144.440 376.670 ;
        RECT 148.880 375.780 149.140 376.670 ;
        RECT 136.040 374.720 136.360 374.820 ;
        RECT 137.400 374.720 137.720 374.900 ;
        RECT 138.090 374.720 138.410 374.890 ;
        RECT 149.980 374.720 150.220 379.320 ;
        RECT 156.020 379.260 158.550 380.060 ;
        RECT 159.300 379.600 182.650 380.060 ;
        RECT 183.420 382.480 183.990 382.490 ;
        RECT 159.300 379.320 173.590 379.600 ;
        RECT 153.290 378.990 158.550 379.260 ;
        RECT 156.020 378.390 158.550 378.990 ;
        RECT 155.900 377.570 158.550 378.390 ;
        RECT 156.050 374.720 156.320 377.570 ;
        RECT 157.830 377.500 158.550 377.570 ;
        RECT 165.960 376.810 166.380 379.320 ;
        RECT 169.680 377.770 173.590 379.320 ;
        RECT 165.920 376.330 166.400 376.810 ;
        RECT 169.660 376.240 173.610 377.770 ;
        RECT 129.020 373.590 156.380 374.720 ;
        RECT 167.050 373.700 167.490 374.200 ;
        RECT 129.020 373.390 156.570 373.590 ;
        RECT 133.120 373.380 133.360 373.390 ;
        RECT 133.120 373.120 133.350 373.380 ;
        RECT 133.110 372.900 133.350 373.120 ;
        RECT 128.190 372.340 128.610 372.820 ;
        RECT 133.120 371.830 133.360 372.470 ;
        RECT 133.120 371.570 133.350 371.830 ;
        RECT 134.080 371.580 134.370 373.390 ;
        RECT 147.440 373.270 147.680 373.390 ;
        RECT 144.180 373.210 144.440 373.230 ;
        RECT 133.110 371.350 133.350 371.570 ;
        RECT 134.060 370.910 134.470 371.580 ;
        RECT 135.320 370.840 135.640 371.160 ;
        RECT 138.320 370.620 138.560 372.500 ;
        RECT 144.140 370.620 144.450 373.210 ;
        RECT 147.440 371.980 147.720 373.270 ;
        RECT 145.180 370.860 145.500 371.180 ;
        RECT 147.440 370.220 147.680 371.980 ;
        RECT 148.100 370.800 148.350 372.670 ;
        RECT 148.100 370.620 148.360 370.800 ;
        RECT 147.390 369.880 147.730 370.220 ;
        RECT 144.640 369.780 145.130 369.790 ;
        RECT 143.730 364.700 144.050 365.020 ;
        RECT 140.710 361.090 140.940 364.570 ;
        RECT 141.380 363.950 141.600 364.570 ;
        RECT 141.350 363.630 141.610 363.950 ;
        RECT 142.190 363.790 142.510 364.110 ;
        RECT 143.740 363.710 144.060 364.030 ;
        RECT 141.380 363.030 141.600 363.630 ;
        RECT 141.320 362.710 141.600 363.030 ;
        RECT 142.170 362.870 142.490 363.190 ;
        RECT 143.740 362.720 144.060 363.040 ;
        RECT 141.380 362.110 141.600 362.710 ;
        RECT 141.330 361.790 141.600 362.110 ;
        RECT 142.150 361.880 142.470 362.200 ;
        RECT 143.650 361.930 143.970 362.250 ;
        RECT 140.680 360.770 140.940 361.090 ;
        RECT 140.710 360.130 140.940 360.770 ;
        RECT 140.640 359.810 140.940 360.130 ;
        RECT 140.710 359.170 140.940 359.810 ;
        RECT 140.680 358.850 140.940 359.170 ;
        RECT 140.710 344.100 140.940 358.850 ;
        RECT 141.380 344.100 141.600 361.790 ;
        RECT 143.480 361.600 143.800 361.640 ;
        RECT 143.250 361.370 143.800 361.600 ;
        RECT 143.480 361.320 143.800 361.370 ;
        RECT 143.650 360.940 143.970 361.260 ;
        RECT 143.480 360.610 143.800 360.650 ;
        RECT 143.250 360.380 143.800 360.610 ;
        RECT 143.480 360.330 143.800 360.380 ;
        RECT 143.650 359.950 143.970 360.270 ;
        RECT 144.070 359.900 144.290 368.840 ;
        RECT 144.630 368.630 145.140 369.780 ;
        RECT 149.980 368.850 150.220 373.390 ;
        RECT 153.260 369.820 153.570 373.390 ;
        RECT 155.050 371.990 156.380 373.390 ;
        RECT 153.180 369.450 153.570 369.820 ;
        RECT 156.050 369.310 156.320 371.990 ;
        RECT 157.220 370.310 157.470 373.460 ;
        RECT 164.260 370.960 164.580 371.010 ;
        RECT 164.170 370.670 164.580 370.960 ;
        RECT 157.180 369.950 157.510 370.310 ;
        RECT 156.010 369.000 156.350 369.310 ;
        RECT 144.580 368.530 145.140 368.630 ;
        RECT 149.930 368.530 150.270 368.850 ;
        RECT 144.050 359.830 144.290 359.900 ;
        RECT 144.470 368.130 145.140 368.530 ;
        RECT 164.170 368.240 164.410 370.670 ;
        RECT 167.110 368.660 167.420 373.700 ;
        RECT 170.340 372.480 173.570 376.240 ;
        RECT 177.190 374.720 177.630 375.220 ;
        RECT 167.050 368.240 167.420 368.660 ;
        RECT 164.170 368.170 164.510 368.240 ;
        RECT 167.050 368.180 167.520 368.240 ;
        RECT 144.470 368.100 145.130 368.130 ;
        RECT 144.470 363.960 144.690 368.100 ;
        RECT 164.170 367.170 164.410 368.170 ;
        RECT 166.310 367.160 166.720 367.490 ;
        RECT 167.050 367.100 167.420 368.180 ;
        RECT 168.470 368.020 168.820 368.310 ;
        RECT 168.470 368.000 168.670 368.020 ;
        RECT 169.430 367.810 169.740 367.820 ;
        RECT 169.430 367.540 169.750 367.810 ;
        RECT 169.450 367.530 169.740 367.540 ;
        RECT 167.050 366.980 167.290 367.100 ;
        RECT 169.990 366.980 170.300 368.670 ;
        RECT 170.470 367.600 170.790 367.880 ;
        RECT 170.470 367.580 170.830 367.600 ;
        RECT 170.550 367.270 170.830 367.580 ;
        RECT 167.050 366.490 167.290 366.910 ;
        RECT 145.690 365.980 146.040 366.440 ;
        RECT 164.270 366.420 164.510 366.490 ;
        RECT 167.050 366.430 167.520 366.490 ;
        RECT 162.120 366.000 162.490 366.310 ;
        RECT 145.090 365.620 145.340 365.740 ;
        RECT 145.060 365.160 145.380 365.620 ;
        RECT 145.090 365.030 145.340 365.160 ;
        RECT 144.820 364.710 145.340 365.030 ;
        RECT 145.090 364.370 145.340 364.710 ;
        RECT 145.090 364.050 145.380 364.370 ;
        RECT 145.090 364.040 145.340 364.050 ;
        RECT 144.470 363.670 144.790 363.960 ;
        RECT 144.830 363.720 145.340 364.040 ;
        RECT 144.050 359.730 144.390 359.830 ;
        RECT 143.480 359.620 143.800 359.660 ;
        RECT 143.250 359.390 143.800 359.620 ;
        RECT 143.480 359.340 143.800 359.390 ;
        RECT 144.070 359.600 144.390 359.730 ;
        RECT 140.600 343.570 140.940 344.100 ;
        RECT 141.260 343.570 141.600 344.100 ;
        RECT 139.290 342.830 139.520 342.900 ;
        RECT 139.250 342.570 139.570 342.830 ;
        RECT 138.800 342.460 139.030 342.500 ;
        RECT 138.760 342.140 139.030 342.460 ;
        RECT 129.450 340.900 130.170 341.600 ;
        RECT 129.460 335.750 130.120 340.900 ;
        RECT 138.800 338.620 139.030 342.140 ;
        RECT 139.290 340.100 139.520 342.570 ;
        RECT 140.710 342.480 140.940 343.570 ;
        RECT 141.380 342.840 141.600 343.570 ;
        RECT 143.140 342.860 143.410 342.900 ;
        RECT 141.360 342.520 141.620 342.840 ;
        RECT 143.120 342.530 143.410 342.860 ;
        RECT 140.700 342.160 140.960 342.480 ;
        RECT 142.590 340.990 142.880 341.020 ;
        RECT 139.290 339.730 140.020 340.100 ;
        RECT 138.800 338.550 139.060 338.620 ;
        RECT 138.780 338.540 139.060 338.550 ;
        RECT 138.750 338.230 139.070 338.540 ;
        RECT 134.650 336.370 135.080 336.800 ;
        RECT 129.460 335.030 130.200 335.750 ;
        RECT 134.700 330.560 135.070 336.370 ;
        RECT 138.610 334.990 138.930 335.310 ;
        RECT 139.290 334.640 139.520 339.730 ;
        RECT 143.140 339.560 143.410 342.530 ;
        RECT 143.020 339.310 143.410 339.560 ;
        RECT 143.620 342.460 143.860 342.500 ;
        RECT 143.620 342.140 143.880 342.460 ;
        RECT 143.620 339.000 143.860 342.140 ;
        RECT 143.020 338.770 143.860 339.000 ;
        RECT 143.620 338.560 143.860 338.770 ;
        RECT 144.070 339.860 144.290 359.600 ;
        RECT 144.470 340.710 144.690 363.670 ;
        RECT 145.090 363.450 145.340 363.720 ;
        RECT 145.090 363.130 145.380 363.450 ;
        RECT 145.090 363.050 145.340 363.130 ;
        RECT 144.830 362.730 145.340 363.050 ;
        RECT 145.090 362.530 145.340 362.730 ;
        RECT 145.090 362.210 145.350 362.530 ;
        RECT 145.090 362.150 145.340 362.210 ;
        RECT 144.950 361.830 145.340 362.150 ;
        RECT 145.090 361.160 145.340 361.830 ;
        RECT 144.950 360.840 145.340 361.160 ;
        RECT 145.090 360.170 145.340 360.840 ;
        RECT 144.950 359.850 145.340 360.170 ;
        RECT 145.090 341.860 145.340 359.850 ;
        RECT 145.710 361.440 145.970 365.980 ;
        RECT 161.480 364.280 161.870 364.650 ;
        RECT 160.900 362.790 161.290 363.180 ;
        RECT 145.710 361.120 145.990 361.440 ;
        RECT 160.260 361.200 160.650 361.580 ;
        RECT 160.290 361.190 160.630 361.200 ;
        RECT 145.710 360.480 145.970 361.120 ;
        RECT 159.650 361.000 159.990 361.010 ;
        RECT 159.640 360.610 160.000 361.000 ;
        RECT 145.710 360.160 146.000 360.480 ;
        RECT 145.710 359.520 145.970 360.160 ;
        RECT 145.710 359.200 145.990 359.520 ;
        RECT 145.090 341.840 145.350 341.860 ;
        RECT 145.080 341.560 145.360 341.840 ;
        RECT 145.090 341.540 145.350 341.560 ;
        RECT 144.430 340.390 144.750 340.710 ;
        RECT 144.070 339.540 144.460 339.860 ;
        RECT 143.620 338.240 143.930 338.560 ;
        RECT 143.620 338.080 143.860 338.240 ;
        RECT 144.070 338.100 144.290 339.540 ;
        RECT 143.500 337.880 143.860 338.080 ;
        RECT 143.500 337.570 143.920 337.880 ;
        RECT 144.030 337.780 144.310 338.100 ;
        RECT 143.620 337.370 143.920 337.570 ;
        RECT 143.620 337.010 143.860 337.370 ;
        RECT 143.620 336.690 143.930 337.010 ;
        RECT 141.920 335.430 142.240 335.750 ;
        RECT 139.710 335.000 140.030 335.320 ;
        RECT 140.800 335.000 141.120 335.320 ;
        RECT 141.930 334.960 142.250 335.280 ;
        RECT 139.160 334.320 139.520 334.640 ;
        RECT 140.260 334.320 140.580 334.640 ;
        RECT 141.360 334.320 141.680 334.640 ;
        RECT 139.290 333.270 139.520 334.320 ;
        RECT 142.210 334.300 142.500 334.730 ;
        RECT 142.210 334.280 142.680 334.300 ;
        RECT 142.220 333.980 142.680 334.280 ;
        RECT 142.220 333.450 142.500 333.980 ;
        RECT 142.230 333.420 142.500 333.450 ;
        RECT 139.160 332.950 139.520 333.270 ;
        RECT 140.260 332.950 140.580 333.270 ;
        RECT 141.360 332.950 141.680 333.270 ;
        RECT 138.610 332.220 138.930 332.540 ;
        RECT 139.290 332.230 139.520 332.950 ;
        RECT 139.710 332.230 140.030 332.540 ;
        RECT 140.800 332.230 141.120 332.540 ;
        RECT 139.290 332.000 141.740 332.230 ;
        RECT 141.420 331.670 141.740 332.000 ;
        RECT 138.600 330.880 138.920 331.200 ;
        RECT 139.710 330.870 140.030 331.190 ;
        RECT 140.800 330.850 141.120 331.170 ;
        RECT 134.660 330.130 135.090 330.560 ;
        RECT 139.160 330.180 139.480 330.500 ;
        RECT 140.260 330.170 140.580 330.490 ;
        RECT 141.350 330.170 141.670 330.490 ;
        RECT 142.180 330.100 142.510 330.130 ;
        RECT 142.040 330.020 142.510 330.100 ;
        RECT 141.800 329.780 142.510 330.020 ;
        RECT 142.180 329.710 142.510 329.780 ;
        RECT 137.670 324.470 137.960 324.820 ;
        RECT 137.680 319.180 137.940 324.470 ;
        RECT 143.620 324.110 143.860 336.690 ;
        RECT 144.070 335.980 144.290 337.780 ;
        RECT 144.470 335.980 144.690 340.390 ;
        RECT 145.090 339.860 145.340 341.540 ;
        RECT 145.360 339.980 145.680 340.300 ;
        RECT 144.840 339.540 145.340 339.860 ;
        RECT 144.070 335.660 144.690 335.980 ;
        RECT 145.090 335.970 145.340 339.540 ;
        RECT 145.710 337.530 145.970 359.200 ;
        RECT 159.030 359.050 159.390 359.440 ;
        RECT 158.380 357.510 158.790 357.910 ;
        RECT 157.850 355.950 158.210 356.340 ;
        RECT 157.270 350.890 157.600 350.910 ;
        RECT 157.210 350.470 157.600 350.890 ;
        RECT 156.640 349.280 156.970 349.300 ;
        RECT 156.590 348.890 156.980 349.280 ;
        RECT 156.020 347.730 156.350 347.740 ;
        RECT 155.990 347.340 156.350 347.730 ;
        RECT 155.370 345.860 155.760 346.260 ;
        RECT 154.700 340.690 155.130 341.090 ;
        RECT 146.010 339.980 146.330 340.300 ;
        RECT 146.390 338.680 146.680 339.590 ;
        RECT 154.040 339.120 154.450 339.520 ;
        RECT 146.300 338.110 146.620 338.150 ;
        RECT 146.300 337.880 146.860 338.110 ;
        RECT 146.300 337.830 146.620 337.880 ;
        RECT 146.310 337.570 146.630 337.610 ;
        RECT 145.700 337.210 146.010 337.530 ;
        RECT 146.310 337.340 146.860 337.570 ;
        RECT 153.430 337.480 153.820 337.880 ;
        RECT 146.310 337.290 146.630 337.340 ;
        RECT 144.070 324.810 144.290 335.660 ;
        RECT 144.470 332.570 144.690 335.660 ;
        RECT 144.860 335.650 145.340 335.970 ;
        RECT 145.090 335.200 145.340 335.650 ;
        RECT 145.090 334.880 145.660 335.200 ;
        RECT 144.470 332.090 144.760 332.570 ;
        RECT 144.470 330.130 144.690 332.090 ;
        RECT 144.450 329.710 144.710 330.130 ;
        RECT 144.470 325.090 144.690 329.710 ;
        RECT 145.090 326.470 145.340 334.880 ;
        RECT 145.050 326.070 145.350 326.470 ;
        RECT 144.470 324.950 144.710 325.090 ;
        RECT 144.030 324.460 144.340 324.810 ;
        RECT 144.480 324.320 144.710 324.950 ;
        RECT 141.320 323.680 141.640 324.000 ;
        RECT 138.010 323.240 138.330 323.560 ;
        RECT 139.110 323.250 139.430 323.570 ;
        RECT 140.200 323.250 140.520 323.570 ;
        RECT 142.830 323.550 143.860 324.110 ;
        RECT 144.470 324.290 144.710 324.320 ;
        RECT 141.330 323.210 141.650 323.530 ;
        RECT 142.830 323.440 143.620 323.550 ;
        RECT 144.470 322.900 144.690 324.290 ;
        RECT 138.560 322.570 138.880 322.890 ;
        RECT 139.660 322.570 139.980 322.890 ;
        RECT 140.760 322.570 141.080 322.890 ;
        RECT 138.560 321.200 138.880 321.520 ;
        RECT 139.660 321.200 139.980 321.520 ;
        RECT 140.760 321.200 141.080 321.520 ;
        RECT 138.010 320.470 138.330 320.790 ;
        RECT 139.110 320.470 139.430 320.790 ;
        RECT 140.200 320.470 140.520 320.790 ;
        RECT 137.630 318.370 137.940 319.180 ;
        RECT 138.000 319.130 138.320 319.450 ;
        RECT 139.110 319.120 139.430 319.440 ;
        RECT 140.200 319.100 140.520 319.420 ;
        RECT 142.940 319.220 145.360 322.900 ;
        RECT 145.710 318.930 145.970 337.210 ;
        RECT 146.380 336.660 146.650 336.840 ;
        RECT 146.360 336.340 146.680 336.660 ;
        RECT 146.380 336.170 146.650 336.340 ;
        RECT 152.740 336.040 153.150 336.430 ;
        RECT 146.050 334.820 146.370 335.140 ;
        RECT 148.530 330.890 149.460 332.540 ;
        RECT 148.620 330.410 149.360 330.890 ;
        RECT 138.560 318.430 138.880 318.750 ;
        RECT 139.660 318.420 139.980 318.740 ;
        RECT 140.750 318.420 141.070 318.740 ;
        RECT 145.620 318.520 145.970 318.930 ;
        RECT 137.680 318.170 137.940 318.370 ;
        RECT 126.690 317.550 127.250 318.070 ;
        RECT 4.170 317.220 6.760 317.450 ;
        RECT 4.170 317.190 4.800 317.220 ;
        RECT 4.650 316.070 5.640 316.080 ;
        RECT 4.250 315.550 5.640 316.070 ;
        RECT 4.250 311.940 4.740 315.550 ;
        RECT 7.450 315.020 10.870 315.070 ;
        RECT 7.440 314.450 10.880 315.020 ;
        RECT 6.030 304.620 10.330 313.680 ;
        RECT 12.010 313.630 12.730 314.180 ;
        RECT 12.010 313.620 12.510 313.630 ;
        RECT 152.800 312.700 153.130 336.040 ;
        RECT 152.750 312.690 153.180 312.700 ;
        RECT 152.720 312.230 153.210 312.690 ;
        RECT 152.750 312.210 153.180 312.230 ;
        RECT 153.450 311.910 153.780 337.480 ;
        RECT 153.360 311.420 153.850 311.910 ;
        RECT 154.100 311.200 154.430 339.120 ;
        RECT 154.070 310.740 154.470 311.200 ;
        RECT 153.860 310.250 154.440 310.360 ;
        RECT 154.770 310.250 155.100 340.690 ;
        RECT 155.410 314.830 155.740 345.860 ;
        RECT 155.410 310.370 155.730 314.830 ;
        RECT 156.020 310.980 156.350 347.340 ;
        RECT 156.640 311.230 156.970 348.890 ;
        RECT 157.270 312.260 157.600 350.470 ;
        RECT 157.870 312.560 158.200 355.950 ;
        RECT 158.450 313.130 158.780 357.510 ;
        RECT 159.060 314.160 159.390 359.050 ;
        RECT 159.650 314.770 159.980 360.610 ;
        RECT 160.290 315.440 160.620 361.190 ;
        RECT 160.910 316.090 161.240 362.790 ;
        RECT 161.510 316.720 161.840 364.280 ;
        RECT 162.140 317.330 162.470 366.000 ;
        RECT 166.310 365.410 166.720 365.740 ;
        RECT 167.050 365.230 167.290 366.430 ;
        RECT 168.470 366.270 168.820 366.560 ;
        RECT 168.470 366.250 168.670 366.270 ;
        RECT 169.430 366.060 169.740 366.070 ;
        RECT 169.430 365.790 169.750 366.060 ;
        RECT 169.450 365.780 169.740 365.790 ;
        RECT 169.990 365.230 170.300 366.920 ;
        RECT 170.470 365.850 170.790 366.130 ;
        RECT 170.470 365.830 170.830 365.850 ;
        RECT 170.550 365.520 170.830 365.830 ;
        RECT 167.050 364.740 167.290 365.160 ;
        RECT 164.270 364.670 164.510 364.740 ;
        RECT 167.050 364.680 167.520 364.740 ;
        RECT 166.310 363.660 166.720 363.990 ;
        RECT 167.050 363.480 167.290 364.680 ;
        RECT 168.470 364.520 168.820 364.810 ;
        RECT 168.470 364.500 168.670 364.520 ;
        RECT 169.430 364.310 169.740 364.320 ;
        RECT 169.430 364.040 169.750 364.310 ;
        RECT 169.450 364.030 169.740 364.040 ;
        RECT 169.990 363.480 170.300 365.170 ;
        RECT 170.470 364.100 170.790 364.380 ;
        RECT 170.470 364.080 170.830 364.100 ;
        RECT 170.550 363.770 170.830 364.080 ;
        RECT 167.050 362.990 167.290 363.410 ;
        RECT 164.270 362.920 164.510 362.990 ;
        RECT 167.050 362.930 167.520 362.990 ;
        RECT 166.310 361.910 166.720 362.240 ;
        RECT 167.050 361.730 167.290 362.930 ;
        RECT 168.470 362.770 168.820 363.060 ;
        RECT 168.470 362.750 168.670 362.770 ;
        RECT 169.430 362.560 169.740 362.570 ;
        RECT 169.430 362.290 169.750 362.560 ;
        RECT 169.450 362.280 169.740 362.290 ;
        RECT 169.990 361.730 170.300 363.420 ;
        RECT 170.470 362.350 170.790 362.630 ;
        RECT 170.470 362.330 170.830 362.350 ;
        RECT 170.550 362.020 170.830 362.330 ;
        RECT 164.270 361.080 164.510 361.290 ;
        RECT 167.210 361.070 167.520 361.300 ;
        RECT 166.310 360.130 166.720 360.460 ;
        RECT 164.270 359.380 164.510 359.450 ;
        RECT 167.050 359.440 167.290 360.640 ;
        RECT 169.450 360.080 169.740 360.090 ;
        RECT 169.430 359.810 169.750 360.080 ;
        RECT 169.430 359.800 169.740 359.810 ;
        RECT 168.470 359.600 168.670 359.620 ;
        RECT 167.050 359.380 167.520 359.440 ;
        RECT 167.050 358.960 167.290 359.380 ;
        RECT 168.470 359.310 168.820 359.600 ;
        RECT 169.990 358.950 170.300 360.640 ;
        RECT 170.550 360.040 170.830 360.350 ;
        RECT 170.470 360.020 170.830 360.040 ;
        RECT 170.470 359.740 170.790 360.020 ;
        RECT 166.310 358.380 166.720 358.710 ;
        RECT 164.270 357.630 164.510 357.700 ;
        RECT 167.050 357.690 167.290 358.890 ;
        RECT 169.450 358.330 169.740 358.340 ;
        RECT 169.430 358.060 169.750 358.330 ;
        RECT 169.430 358.050 169.740 358.060 ;
        RECT 168.470 357.850 168.670 357.870 ;
        RECT 167.050 357.630 167.520 357.690 ;
        RECT 167.050 357.210 167.290 357.630 ;
        RECT 168.470 357.560 168.820 357.850 ;
        RECT 169.990 357.200 170.300 358.890 ;
        RECT 170.550 358.290 170.830 358.600 ;
        RECT 170.470 358.270 170.830 358.290 ;
        RECT 170.470 357.990 170.790 358.270 ;
        RECT 166.310 356.630 166.720 356.960 ;
        RECT 164.270 355.880 164.510 355.950 ;
        RECT 167.050 355.940 167.290 357.140 ;
        RECT 169.450 356.580 169.740 356.590 ;
        RECT 169.430 356.310 169.750 356.580 ;
        RECT 169.430 356.300 169.740 356.310 ;
        RECT 168.470 356.100 168.670 356.120 ;
        RECT 167.050 355.880 167.520 355.940 ;
        RECT 167.050 355.460 167.290 355.880 ;
        RECT 168.470 355.810 168.820 356.100 ;
        RECT 169.990 355.450 170.300 357.140 ;
        RECT 170.550 356.540 170.830 356.850 ;
        RECT 170.470 356.520 170.830 356.540 ;
        RECT 170.470 356.240 170.790 356.520 ;
        RECT 164.170 354.200 164.410 355.090 ;
        RECT 166.310 354.880 166.720 355.210 ;
        RECT 167.050 355.160 167.290 355.390 ;
        RECT 164.170 354.130 164.510 354.200 ;
        RECT 167.050 354.190 167.420 355.160 ;
        RECT 169.450 354.830 169.740 354.840 ;
        RECT 169.430 354.560 169.750 354.830 ;
        RECT 169.430 354.550 169.740 354.560 ;
        RECT 168.470 354.350 168.670 354.370 ;
        RECT 167.050 354.130 167.520 354.190 ;
        RECT 164.170 351.000 164.410 354.130 ;
        RECT 167.050 353.710 167.420 354.130 ;
        RECT 168.470 354.060 168.820 354.350 ;
        RECT 167.110 351.000 167.420 353.710 ;
        RECT 169.990 353.700 170.300 355.390 ;
        RECT 170.550 354.790 170.830 355.100 ;
        RECT 170.470 354.770 170.830 354.790 ;
        RECT 170.470 354.490 170.790 354.770 ;
        RECT 164.170 350.950 164.510 351.000 ;
        RECT 164.170 350.720 164.410 350.950 ;
        RECT 167.110 350.940 167.520 351.000 ;
        RECT 167.110 350.650 167.420 350.940 ;
        RECT 166.310 350.000 166.720 350.330 ;
        RECT 164.270 349.250 164.510 349.320 ;
        RECT 167.050 349.310 167.290 350.510 ;
        RECT 169.450 349.950 169.740 349.960 ;
        RECT 169.430 349.680 169.750 349.950 ;
        RECT 169.430 349.670 169.740 349.680 ;
        RECT 168.470 349.470 168.670 349.490 ;
        RECT 167.050 349.250 167.520 349.310 ;
        RECT 167.050 348.830 167.290 349.250 ;
        RECT 168.470 349.180 168.820 349.470 ;
        RECT 169.990 348.820 170.300 350.510 ;
        RECT 170.550 349.910 170.830 350.220 ;
        RECT 170.470 349.890 170.830 349.910 ;
        RECT 170.470 349.610 170.790 349.890 ;
        RECT 166.310 348.250 166.720 348.580 ;
        RECT 164.270 347.500 164.510 347.570 ;
        RECT 167.050 347.560 167.290 348.760 ;
        RECT 169.450 348.200 169.740 348.210 ;
        RECT 169.430 347.930 169.750 348.200 ;
        RECT 169.430 347.920 169.740 347.930 ;
        RECT 168.470 347.720 168.670 347.740 ;
        RECT 167.050 347.500 167.520 347.560 ;
        RECT 167.050 347.080 167.290 347.500 ;
        RECT 168.470 347.430 168.820 347.720 ;
        RECT 169.990 347.070 170.300 348.760 ;
        RECT 170.550 348.160 170.830 348.470 ;
        RECT 170.470 348.140 170.830 348.160 ;
        RECT 170.470 347.860 170.790 348.140 ;
        RECT 166.310 346.500 166.720 346.830 ;
        RECT 164.270 345.750 164.510 345.820 ;
        RECT 167.050 345.810 167.290 347.010 ;
        RECT 169.450 346.450 169.740 346.460 ;
        RECT 169.430 346.180 169.750 346.450 ;
        RECT 169.430 346.170 169.740 346.180 ;
        RECT 168.470 345.970 168.670 345.990 ;
        RECT 167.050 345.750 167.520 345.810 ;
        RECT 167.050 345.330 167.290 345.750 ;
        RECT 168.470 345.680 168.820 345.970 ;
        RECT 169.990 345.320 170.300 347.010 ;
        RECT 170.550 346.410 170.830 346.720 ;
        RECT 170.470 346.390 170.830 346.410 ;
        RECT 170.470 346.110 170.790 346.390 ;
        RECT 164.170 344.100 164.410 344.960 ;
        RECT 166.310 344.750 166.720 345.080 ;
        RECT 167.050 345.030 167.290 345.260 ;
        RECT 167.050 344.100 167.420 345.030 ;
        RECT 169.450 344.700 169.740 344.710 ;
        RECT 169.430 344.430 169.750 344.700 ;
        RECT 169.430 344.420 169.740 344.430 ;
        RECT 168.470 344.220 168.670 344.240 ;
        RECT 164.170 341.190 164.510 344.100 ;
        RECT 167.050 343.580 167.520 344.100 ;
        RECT 168.470 343.930 168.820 344.220 ;
        RECT 167.110 341.450 167.520 343.580 ;
        RECT 169.990 343.570 170.300 345.260 ;
        RECT 170.550 344.660 170.830 344.970 ;
        RECT 170.470 344.640 170.830 344.660 ;
        RECT 170.470 344.360 170.790 344.640 ;
        RECT 171.540 341.940 171.830 372.480 ;
        RECT 173.000 361.000 173.190 372.480 ;
        RECT 172.720 360.510 173.190 361.000 ;
        RECT 173.580 360.860 173.950 360.880 ;
        RECT 173.530 360.600 173.950 360.860 ;
        RECT 173.580 360.590 173.950 360.600 ;
        RECT 172.540 360.070 172.860 360.350 ;
        RECT 173.000 360.170 173.190 360.510 ;
        RECT 172.900 359.880 173.190 360.170 ;
        RECT 173.000 359.270 173.190 359.880 ;
        RECT 172.540 358.800 172.860 359.080 ;
        RECT 172.900 358.980 173.190 359.270 ;
        RECT 173.000 358.640 173.190 358.980 ;
        RECT 172.720 358.150 173.190 358.640 ;
        RECT 173.580 358.550 173.950 358.560 ;
        RECT 173.530 358.290 173.950 358.550 ;
        RECT 173.580 358.270 173.950 358.290 ;
        RECT 173.000 357.800 173.190 358.150 ;
        RECT 172.720 357.310 173.190 357.800 ;
        RECT 173.580 357.660 173.950 357.680 ;
        RECT 173.530 357.400 173.950 357.660 ;
        RECT 173.580 357.390 173.950 357.400 ;
        RECT 172.540 356.870 172.860 357.150 ;
        RECT 173.000 356.970 173.190 357.310 ;
        RECT 172.900 356.680 173.190 356.970 ;
        RECT 173.000 356.070 173.190 356.680 ;
        RECT 172.540 355.600 172.860 355.880 ;
        RECT 172.900 355.780 173.190 356.070 ;
        RECT 173.000 355.440 173.190 355.780 ;
        RECT 172.720 354.950 173.190 355.440 ;
        RECT 173.580 355.350 173.950 355.360 ;
        RECT 173.530 355.090 173.950 355.350 ;
        RECT 173.580 355.070 173.950 355.090 ;
        RECT 173.000 351.180 173.190 354.950 ;
        RECT 174.310 351.280 174.540 361.220 ;
        RECT 177.280 361.000 177.530 374.720 ;
        RECT 178.980 374.680 179.710 379.600 ;
        RECT 183.420 379.060 184.040 382.480 ;
        RECT 184.130 381.400 185.110 381.550 ;
        RECT 183.420 379.050 183.990 379.060 ;
        RECT 182.590 377.420 183.150 377.920 ;
        RECT 182.600 377.200 183.150 377.420 ;
        RECT 181.980 376.630 182.590 376.770 ;
        RECT 179.140 364.290 179.310 374.680 ;
        RECT 181.960 374.670 183.140 376.630 ;
        RECT 181.160 373.760 183.140 374.670 ;
        RECT 184.140 374.150 185.110 381.400 ;
        RECT 186.420 377.500 187.140 383.170 ;
        RECT 187.890 383.900 202.180 384.460 ;
        RECT 212.810 384.290 213.640 385.190 ;
        RECT 214.750 385.130 217.120 385.760 ;
        RECT 187.890 383.650 211.240 383.900 ;
        RECT 212.810 383.650 213.530 384.290 ;
        RECT 187.890 382.930 213.530 383.650 ;
        RECT 214.780 383.170 215.730 385.130 ;
        RECT 216.480 385.110 217.060 385.130 ;
        RECT 226.860 384.470 230.770 385.930 ;
        RECT 238.090 385.280 242.220 385.680 ;
        RECT 238.090 385.190 242.230 385.280 ;
        RECT 217.150 384.460 230.770 384.470 ;
        RECT 187.890 379.600 211.240 382.930 ;
        RECT 212.010 382.480 212.580 382.490 ;
        RECT 187.890 379.320 202.180 379.600 ;
        RECT 197.480 377.770 202.180 379.320 ;
        RECT 181.160 373.580 182.970 373.760 ;
        RECT 184.120 373.680 185.130 374.150 ;
        RECT 186.400 373.600 187.120 377.460 ;
        RECT 189.530 376.310 191.000 376.840 ;
        RECT 187.160 373.700 187.600 374.200 ;
        RECT 181.160 372.890 181.890 373.580 ;
        RECT 181.360 369.950 181.700 370.240 ;
        RECT 181.410 369.920 181.670 369.950 ;
        RECT 179.530 366.390 179.790 366.710 ;
        RECT 179.560 364.160 179.750 366.390 ;
        RECT 181.430 364.140 181.640 369.920 ;
        RECT 185.000 369.320 185.260 369.330 ;
        RECT 184.980 369.020 185.280 369.320 ;
        RECT 185.000 369.010 185.260 369.020 ;
        RECT 181.830 367.990 182.170 368.310 ;
        RECT 181.900 364.160 182.090 367.990 ;
        RECT 182.270 365.900 182.560 366.220 ;
        RECT 182.310 364.140 182.520 365.900 ;
        RECT 183.310 365.420 183.650 365.740 ;
        RECT 183.390 364.170 183.570 365.420 ;
        RECT 176.040 360.840 176.380 360.890 ;
        RECT 176.040 360.820 176.600 360.840 ;
        RECT 175.920 360.650 176.600 360.820 ;
        RECT 176.040 360.610 176.600 360.650 ;
        RECT 176.040 360.570 176.380 360.610 ;
        RECT 177.280 359.930 177.920 361.000 ;
        RECT 177.280 359.220 177.530 359.930 ;
        RECT 176.040 358.540 176.380 358.580 ;
        RECT 176.040 358.500 176.600 358.540 ;
        RECT 175.920 358.330 176.600 358.500 ;
        RECT 176.040 358.310 176.600 358.330 ;
        RECT 176.040 358.260 176.380 358.310 ;
        RECT 177.280 358.150 177.920 359.220 ;
        RECT 185.030 358.780 185.230 369.010 ;
        RECT 187.260 364.120 187.490 373.700 ;
        RECT 188.160 369.930 188.440 370.250 ;
        RECT 187.720 369.020 188.000 369.340 ;
        RECT 185.010 358.650 185.230 358.780 ;
        RECT 184.960 358.320 185.290 358.650 ;
        RECT 187.490 358.210 187.500 358.370 ;
        RECT 177.280 357.800 177.530 358.150 ;
        RECT 176.040 357.640 176.380 357.690 ;
        RECT 176.040 357.620 176.600 357.640 ;
        RECT 175.920 357.450 176.600 357.620 ;
        RECT 176.040 357.410 176.600 357.450 ;
        RECT 176.040 357.370 176.380 357.410 ;
        RECT 177.280 356.730 177.920 357.800 ;
        RECT 187.750 357.480 187.970 369.020 ;
        RECT 187.740 357.410 187.970 357.480 ;
        RECT 187.730 356.810 187.930 357.410 ;
        RECT 188.180 356.960 188.410 369.930 ;
        RECT 189.550 363.930 189.970 376.310 ;
        RECT 190.580 363.930 191.000 376.310 ;
        RECT 197.480 376.230 202.200 377.770 ;
        RECT 192.960 373.660 193.400 374.160 ;
        RECT 193.060 366.680 193.290 373.660 ;
        RECT 197.480 368.410 198.760 376.230 ;
        RECT 198.930 372.480 202.160 376.230 ;
        RECT 197.480 368.330 198.780 368.410 ;
        RECT 197.470 368.030 198.780 368.330 ;
        RECT 194.250 367.380 194.550 367.700 ;
        RECT 192.930 366.670 193.290 366.680 ;
        RECT 192.900 365.780 193.290 366.670 ;
        RECT 193.060 364.120 193.290 365.780 ;
        RECT 194.280 364.120 194.510 367.380 ;
        RECT 200.560 366.830 200.990 367.170 ;
        RECT 200.800 364.160 200.990 366.830 ;
        RECT 201.240 366.640 201.520 372.480 ;
        RECT 201.240 366.040 201.600 366.640 ;
        RECT 201.240 364.070 201.520 366.040 ;
        RECT 201.740 365.830 201.930 367.280 ;
        RECT 202.010 366.950 202.400 370.540 ;
        RECT 202.940 369.930 203.200 370.250 ;
        RECT 201.710 365.800 201.930 365.830 ;
        RECT 201.700 365.530 201.950 365.800 ;
        RECT 201.700 365.520 201.940 365.530 ;
        RECT 201.710 365.340 201.940 365.520 ;
        RECT 202.080 365.340 202.270 366.950 ;
        RECT 202.960 366.910 203.180 369.930 ;
        RECT 202.960 366.470 203.450 366.910 ;
        RECT 204.930 366.710 205.270 379.600 ;
        RECT 209.430 379.470 209.800 379.480 ;
        RECT 209.380 379.020 209.880 379.470 ;
        RECT 212.010 379.060 212.630 382.480 ;
        RECT 212.010 379.050 212.580 379.060 ;
        RECT 205.580 370.610 205.900 370.980 ;
        RECT 204.880 366.630 205.270 366.710 ;
        RECT 202.960 365.340 203.180 366.470 ;
        RECT 204.870 365.860 205.270 366.630 ;
        RECT 204.880 365.790 205.270 365.860 ;
        RECT 201.710 365.280 202.590 365.340 ;
        RECT 201.740 364.260 201.900 365.280 ;
        RECT 201.910 364.650 202.590 365.280 ;
        RECT 202.950 364.650 203.630 365.340 ;
        RECT 202.090 364.510 202.330 364.650 ;
        RECT 201.330 361.740 201.490 363.430 ;
        RECT 201.740 362.410 201.900 363.430 ;
        RECT 201.710 362.170 201.940 362.410 ;
        RECT 201.700 362.160 201.940 362.170 ;
        RECT 201.700 361.890 201.950 362.160 ;
        RECT 201.710 361.860 201.930 361.890 ;
        RECT 201.320 361.650 201.490 361.740 ;
        RECT 201.320 361.600 201.600 361.650 ;
        RECT 201.330 361.250 201.600 361.600 ;
        RECT 201.740 361.250 201.930 361.860 ;
        RECT 201.320 361.050 201.600 361.250 ;
        RECT 201.320 360.610 201.490 361.050 ;
        RECT 201.320 360.060 201.590 360.610 ;
        RECT 201.310 360.010 201.590 360.060 ;
        RECT 201.730 360.410 201.930 361.250 ;
        RECT 202.000 360.920 202.390 364.510 ;
        RECT 204.930 364.010 205.270 365.790 ;
        RECT 205.600 365.230 205.870 370.610 ;
        RECT 209.430 366.870 209.800 379.020 ;
        RECT 211.180 377.420 211.740 377.920 ;
        RECT 215.010 377.500 215.730 383.170 ;
        RECT 216.480 383.900 230.770 384.460 ;
        RECT 241.700 384.290 242.230 385.190 ;
        RECT 243.340 385.130 245.710 385.760 ;
        RECT 216.480 379.600 239.830 383.900 ;
        RECT 243.370 383.170 244.320 385.130 ;
        RECT 245.070 385.110 245.650 385.130 ;
        RECT 255.450 384.470 259.360 385.930 ;
        RECT 266.680 385.280 270.810 385.680 ;
        RECT 266.680 385.190 270.820 385.280 ;
        RECT 245.740 384.460 259.360 384.470 ;
        RECT 240.600 382.480 241.170 382.490 ;
        RECT 216.480 379.320 230.770 379.600 ;
        RECT 226.420 377.770 230.770 379.320 ;
        RECT 211.190 377.200 211.740 377.420 ;
        RECT 226.420 376.230 230.790 377.770 ;
        RECT 210.220 375.570 210.680 376.000 ;
        RECT 206.090 366.820 206.250 366.870 ;
        RECT 206.500 366.810 206.690 366.870 ;
        RECT 208.370 366.580 208.580 366.870 ;
        RECT 208.260 366.290 208.580 366.580 ;
        RECT 205.600 364.730 206.280 365.230 ;
        RECT 205.600 364.080 205.870 364.730 ;
        RECT 207.360 364.670 207.680 364.990 ;
        RECT 208.370 364.590 208.580 366.290 ;
        RECT 208.840 366.020 209.030 366.870 ;
        RECT 208.730 365.730 209.030 366.020 ;
        RECT 208.260 364.300 208.580 364.590 ;
        RECT 206.730 364.050 206.990 364.110 ;
        RECT 208.370 364.080 208.580 364.300 ;
        RECT 206.730 363.790 207.090 364.050 ;
        RECT 206.850 363.630 207.090 363.790 ;
        RECT 208.840 363.700 209.030 365.730 ;
        RECT 209.250 364.410 209.800 366.870 ;
        RECT 209.130 363.900 209.800 364.410 ;
        RECT 208.390 363.520 208.580 363.570 ;
        RECT 207.350 362.980 207.670 363.300 ;
        RECT 208.270 363.230 208.580 363.520 ;
        RECT 208.730 363.410 209.030 363.700 ;
        RECT 208.390 361.610 208.580 363.230 ;
        RECT 208.840 362.120 209.030 363.410 ;
        RECT 208.720 361.830 209.030 362.120 ;
        RECT 208.070 361.320 208.080 361.330 ;
        RECT 208.290 361.320 208.580 361.610 ;
        RECT 203.140 360.880 203.450 361.220 ;
        RECT 203.130 360.780 203.450 360.880 ;
        RECT 206.090 360.840 206.250 360.870 ;
        RECT 206.500 360.840 206.690 360.870 ;
        RECT 205.960 360.820 206.250 360.840 ;
        RECT 206.490 360.820 206.690 360.840 ;
        RECT 208.380 360.820 208.610 361.320 ;
        RECT 208.840 360.820 209.030 361.830 ;
        RECT 209.250 360.820 209.800 363.900 ;
        RECT 210.240 363.000 210.610 375.570 ;
        RECT 226.420 372.480 230.750 376.230 ;
        RECT 210.990 370.860 211.440 371.290 ;
        RECT 210.040 362.980 210.200 363.000 ;
        RECT 209.880 362.680 210.200 362.980 ;
        RECT 210.240 362.940 210.640 363.000 ;
        RECT 203.130 360.440 203.440 360.780 ;
        RECT 201.310 359.920 201.480 360.010 ;
        RECT 201.320 358.230 201.480 359.920 ;
        RECT 201.730 359.800 201.920 360.410 ;
        RECT 201.700 359.770 201.920 359.800 ;
        RECT 201.690 359.500 201.940 359.770 ;
        RECT 201.690 359.490 201.930 359.500 ;
        RECT 201.700 359.250 201.930 359.490 ;
        RECT 201.730 358.230 201.890 359.250 ;
        RECT 202.080 358.440 202.320 358.820 ;
        RECT 187.740 356.780 187.970 356.810 ;
        RECT 177.280 356.020 177.530 356.730 ;
        RECT 176.040 355.340 176.380 355.380 ;
        RECT 176.040 355.300 176.600 355.340 ;
        RECT 175.920 355.130 176.600 355.300 ;
        RECT 176.040 355.110 176.600 355.130 ;
        RECT 176.040 355.060 176.380 355.110 ;
        RECT 177.280 354.950 177.920 356.020 ;
        RECT 177.280 351.290 177.530 354.950 ;
        RECT 187.750 353.580 187.970 356.780 ;
        RECT 201.320 355.710 201.480 357.400 ;
        RECT 201.730 356.380 201.890 357.400 ;
        RECT 202.080 356.810 202.320 357.190 ;
        RECT 201.700 356.140 201.930 356.380 ;
        RECT 201.690 356.130 201.930 356.140 ;
        RECT 201.690 355.860 201.940 356.130 ;
        RECT 201.700 355.830 201.920 355.860 ;
        RECT 201.310 355.620 201.480 355.710 ;
        RECT 201.310 355.570 201.590 355.620 ;
        RECT 201.320 355.020 201.590 355.570 ;
        RECT 201.320 354.380 201.480 355.020 ;
        RECT 201.730 354.380 201.920 355.830 ;
        RECT 203.130 354.750 203.440 355.190 ;
        RECT 205.960 354.790 206.240 360.820 ;
        RECT 206.490 360.780 206.680 360.820 ;
        RECT 207.590 359.210 207.910 359.530 ;
        RECT 206.730 358.050 206.990 358.370 ;
        RECT 206.730 357.450 206.990 357.770 ;
        RECT 207.590 356.450 207.910 356.770 ;
        RECT 206.490 354.790 206.680 354.850 ;
        RECT 187.750 353.490 188.100 353.580 ;
        RECT 172.980 350.680 173.190 351.180 ;
        RECT 174.290 350.870 174.540 351.280 ;
        RECT 177.260 350.870 177.530 351.290 ;
        RECT 179.040 351.440 179.320 352.550 ;
        RECT 179.570 351.860 179.760 352.460 ;
        RECT 181.570 352.020 181.960 352.040 ;
        RECT 181.560 351.930 181.960 352.020 ;
        RECT 181.410 351.920 181.960 351.930 ;
        RECT 179.570 351.670 181.170 351.860 ;
        RECT 179.040 351.160 180.760 351.440 ;
        RECT 180.560 350.930 180.760 351.160 ;
        RECT 172.980 350.530 173.170 350.680 ;
        RECT 172.700 350.040 173.170 350.530 ;
        RECT 173.560 350.390 173.930 350.410 ;
        RECT 173.510 350.130 173.930 350.390 ;
        RECT 173.560 350.120 173.930 350.130 ;
        RECT 172.520 349.600 172.840 349.880 ;
        RECT 172.980 349.700 173.170 350.040 ;
        RECT 172.880 349.410 173.170 349.700 ;
        RECT 172.980 348.800 173.170 349.410 ;
        RECT 172.520 348.330 172.840 348.610 ;
        RECT 172.880 348.510 173.170 348.800 ;
        RECT 172.980 348.170 173.170 348.510 ;
        RECT 172.700 347.680 173.170 348.170 ;
        RECT 173.560 348.080 173.930 348.090 ;
        RECT 173.510 347.820 173.930 348.080 ;
        RECT 173.560 347.800 173.930 347.820 ;
        RECT 172.980 347.330 173.170 347.680 ;
        RECT 172.700 346.840 173.170 347.330 ;
        RECT 173.560 347.190 173.930 347.210 ;
        RECT 173.510 346.930 173.930 347.190 ;
        RECT 173.560 346.920 173.930 346.930 ;
        RECT 172.520 346.400 172.840 346.680 ;
        RECT 172.980 346.500 173.170 346.840 ;
        RECT 172.880 346.210 173.170 346.500 ;
        RECT 172.980 345.600 173.170 346.210 ;
        RECT 172.520 345.130 172.840 345.410 ;
        RECT 172.880 345.310 173.170 345.600 ;
        RECT 172.980 345.010 173.170 345.310 ;
        RECT 174.290 345.050 174.520 350.870 ;
        RECT 177.260 350.530 177.510 350.870 ;
        RECT 180.570 350.630 180.730 350.930 ;
        RECT 180.980 350.550 181.170 351.670 ;
        RECT 181.380 351.680 181.960 351.920 ;
        RECT 181.380 351.660 181.950 351.680 ;
        RECT 181.380 351.650 181.570 351.660 ;
        RECT 181.380 350.810 181.550 351.650 ;
        RECT 186.050 351.590 186.280 352.500 ;
        RECT 185.530 351.520 186.280 351.590 ;
        RECT 185.500 351.360 186.280 351.520 ;
        RECT 187.230 351.460 187.620 353.320 ;
        RECT 187.750 353.270 188.260 353.490 ;
        RECT 190.580 351.690 191.000 352.690 ;
        RECT 190.580 351.510 191.010 351.690 ;
        RECT 191.260 351.530 191.650 353.390 ;
        RECT 185.500 350.910 185.910 351.360 ;
        RECT 181.380 350.540 181.540 350.810 ;
        RECT 176.020 350.370 176.360 350.420 ;
        RECT 176.020 350.350 176.580 350.370 ;
        RECT 175.900 350.180 176.580 350.350 ;
        RECT 176.020 350.140 176.580 350.180 ;
        RECT 176.020 350.100 176.360 350.140 ;
        RECT 177.260 349.460 177.900 350.530 ;
        RECT 185.500 350.420 185.880 350.910 ;
        RECT 187.250 350.560 187.490 351.460 ;
        RECT 190.580 351.120 191.020 351.510 ;
        RECT 193.060 351.300 193.290 352.500 ;
        RECT 190.610 350.910 191.020 351.120 ;
        RECT 190.610 350.400 191.010 350.910 ;
        RECT 193.050 350.560 193.290 351.300 ;
        RECT 194.280 351.610 194.510 352.500 ;
        RECT 194.280 351.230 195.040 351.610 ;
        RECT 200.800 351.480 200.990 352.460 ;
        RECT 194.660 350.770 195.040 351.230 ;
        RECT 198.970 351.110 199.250 351.430 ;
        RECT 199.400 351.290 200.990 351.480 ;
        RECT 196.780 350.930 196.940 351.050 ;
        RECT 196.630 350.790 196.940 350.930 ;
        RECT 196.620 350.640 196.940 350.790 ;
        RECT 196.780 350.350 196.940 350.640 ;
        RECT 196.780 349.800 197.050 350.350 ;
        RECT 196.770 349.750 197.050 349.800 ;
        RECT 197.190 350.010 197.380 351.000 ;
        RECT 197.590 350.320 197.750 351.050 ;
        RECT 198.430 350.460 198.750 350.780 ;
        RECT 199.000 350.630 199.160 351.110 ;
        RECT 199.400 351.060 199.590 351.290 ;
        RECT 201.240 351.100 201.520 352.550 ;
        RECT 209.430 352.110 209.800 360.820 ;
        RECT 210.240 356.970 210.610 362.940 ;
        RECT 209.920 356.920 210.200 356.970 ;
        RECT 210.240 356.920 210.640 356.970 ;
        RECT 209.920 356.910 210.640 356.920 ;
        RECT 209.920 356.640 210.610 356.910 ;
        RECT 209.400 351.650 209.850 352.110 ;
        RECT 209.430 351.610 209.800 351.650 ;
        RECT 210.240 351.520 210.610 356.640 ;
        RECT 199.850 351.090 201.520 351.100 ;
        RECT 199.400 350.960 199.770 351.060 ;
        RECT 199.370 350.550 199.770 350.960 ;
        RECT 199.810 350.820 201.520 351.090 ;
        RECT 210.210 351.060 210.650 351.520 ;
        RECT 211.010 351.060 211.380 370.860 ;
        RECT 217.560 369.810 218.140 370.370 ;
        RECT 214.350 368.240 214.910 368.890 ;
        RECT 215.300 368.730 215.860 369.310 ;
        RECT 216.380 369.190 216.940 369.780 ;
        RECT 214.370 366.870 214.870 368.240 ;
        RECT 211.880 365.780 212.310 366.220 ;
        RECT 199.810 350.630 199.970 350.820 ;
        RECT 197.550 350.300 197.750 350.320 ;
        RECT 197.540 350.060 197.770 350.300 ;
        RECT 197.540 350.010 197.750 350.060 ;
        RECT 197.190 349.890 197.360 350.010 ;
        RECT 196.770 349.660 196.940 349.750 ;
        RECT 177.260 348.750 177.510 349.460 ;
        RECT 196.780 349.190 196.940 349.660 ;
        RECT 196.770 349.100 196.940 349.190 ;
        RECT 196.770 349.050 197.050 349.100 ;
        RECT 176.020 348.070 176.360 348.110 ;
        RECT 176.020 348.030 176.580 348.070 ;
        RECT 175.900 347.860 176.580 348.030 ;
        RECT 176.020 347.840 176.580 347.860 ;
        RECT 176.020 347.790 176.360 347.840 ;
        RECT 177.260 347.680 177.900 348.750 ;
        RECT 196.780 348.500 197.050 349.050 ;
        RECT 197.190 348.960 197.350 349.890 ;
        RECT 197.190 348.840 197.360 348.960 ;
        RECT 197.590 348.840 197.750 350.010 ;
        RECT 198.430 349.910 198.750 350.230 ;
        RECT 199.530 349.670 199.770 350.550 ;
        RECT 199.520 349.010 199.790 349.670 ;
        RECT 177.260 347.330 177.510 347.680 ;
        RECT 176.020 347.170 176.360 347.220 ;
        RECT 176.020 347.150 176.580 347.170 ;
        RECT 175.900 346.980 176.580 347.150 ;
        RECT 176.020 346.940 176.580 346.980 ;
        RECT 176.020 346.900 176.360 346.940 ;
        RECT 177.260 346.260 177.900 347.330 ;
        RECT 185.190 346.440 185.580 348.300 ;
        RECT 189.220 346.510 189.610 348.370 ;
        RECT 196.780 347.110 196.940 348.500 ;
        RECT 197.190 347.920 197.380 348.840 ;
        RECT 197.540 348.790 197.750 348.840 ;
        RECT 197.540 348.550 197.770 348.790 ;
        RECT 198.430 348.620 198.750 348.940 ;
        RECT 197.550 348.530 197.750 348.550 ;
        RECT 197.160 347.900 197.400 347.920 ;
        RECT 197.590 347.900 197.750 348.530 ;
        RECT 198.430 348.070 198.750 348.390 ;
        RECT 197.160 347.710 197.750 347.900 ;
        RECT 197.160 347.690 197.400 347.710 ;
        RECT 196.780 346.560 197.050 347.110 ;
        RECT 196.770 346.510 197.050 346.560 ;
        RECT 197.190 346.770 197.380 347.690 ;
        RECT 197.590 347.080 197.750 347.710 ;
        RECT 198.430 347.220 198.750 347.540 ;
        RECT 197.550 347.060 197.750 347.080 ;
        RECT 197.540 346.820 197.770 347.060 ;
        RECT 197.540 346.770 197.750 346.820 ;
        RECT 197.190 346.650 197.360 346.770 ;
        RECT 196.770 346.420 196.940 346.510 ;
        RECT 177.260 345.550 177.510 346.260 ;
        RECT 172.980 344.970 173.190 345.010 ;
        RECT 172.700 344.480 173.190 344.970 ;
        RECT 173.560 344.880 173.930 344.890 ;
        RECT 173.510 344.620 173.930 344.880 ;
        RECT 173.560 344.600 173.930 344.620 ;
        RECT 172.980 344.260 173.190 344.480 ;
        RECT 174.290 344.260 174.540 345.050 ;
        RECT 176.020 344.870 176.360 344.910 ;
        RECT 176.020 344.830 176.580 344.870 ;
        RECT 175.900 344.660 176.580 344.830 ;
        RECT 176.020 344.640 176.580 344.660 ;
        RECT 176.020 344.590 176.360 344.640 ;
        RECT 177.260 344.480 177.900 345.550 ;
        RECT 194.740 345.370 194.900 346.070 ;
        RECT 177.260 344.260 177.530 344.480 ;
        RECT 164.270 340.950 164.510 341.190 ;
        RECT 166.270 340.940 166.680 341.270 ;
        RECT 167.010 340.920 167.520 341.450 ;
        RECT 164.230 340.190 164.470 340.260 ;
        RECT 167.010 340.250 167.250 340.920 ;
        RECT 169.410 340.890 169.700 340.900 ;
        RECT 169.390 340.620 169.710 340.890 ;
        RECT 169.390 340.610 169.700 340.620 ;
        RECT 168.430 340.410 168.630 340.430 ;
        RECT 167.010 340.190 167.480 340.250 ;
        RECT 167.010 339.770 167.250 340.190 ;
        RECT 168.430 340.120 168.780 340.410 ;
        RECT 169.950 339.760 170.260 341.450 ;
        RECT 171.500 341.190 171.830 341.940 ;
        RECT 173.000 341.480 173.190 344.260 ;
        RECT 174.310 343.970 174.540 344.260 ;
        RECT 174.220 343.490 174.550 343.970 ;
        RECT 174.310 341.480 174.540 343.490 ;
        RECT 177.280 341.480 177.530 344.260 ;
        RECT 173.000 341.260 173.200 341.480 ;
        RECT 170.510 340.850 170.790 341.160 ;
        RECT 170.430 340.830 170.790 340.850 ;
        RECT 170.430 340.550 170.750 340.830 ;
        RECT 166.270 339.190 166.680 339.520 ;
        RECT 164.230 338.440 164.470 338.510 ;
        RECT 167.010 338.500 167.250 339.700 ;
        RECT 169.410 339.140 169.700 339.150 ;
        RECT 169.390 338.870 169.710 339.140 ;
        RECT 169.390 338.860 169.700 338.870 ;
        RECT 168.430 338.660 168.630 338.680 ;
        RECT 167.010 338.440 167.480 338.500 ;
        RECT 167.010 338.020 167.250 338.440 ;
        RECT 168.430 338.370 168.780 338.660 ;
        RECT 169.950 338.010 170.260 339.700 ;
        RECT 170.510 339.100 170.790 339.410 ;
        RECT 170.430 339.080 170.790 339.100 ;
        RECT 170.430 338.800 170.750 339.080 ;
        RECT 166.270 337.440 166.680 337.770 ;
        RECT 164.230 336.690 164.470 336.760 ;
        RECT 167.010 336.750 167.250 337.950 ;
        RECT 169.410 337.390 169.700 337.400 ;
        RECT 169.390 337.120 169.710 337.390 ;
        RECT 169.390 337.110 169.700 337.120 ;
        RECT 168.430 336.910 168.630 336.930 ;
        RECT 167.010 336.690 167.480 336.750 ;
        RECT 167.010 336.270 167.250 336.690 ;
        RECT 168.430 336.620 168.780 336.910 ;
        RECT 169.950 336.260 170.260 337.950 ;
        RECT 170.510 337.350 170.790 337.660 ;
        RECT 170.430 337.330 170.790 337.350 ;
        RECT 170.430 337.050 170.750 337.330 ;
        RECT 166.270 335.690 166.680 336.020 ;
        RECT 167.010 335.260 167.250 336.200 ;
        RECT 169.410 335.640 169.700 335.650 ;
        RECT 169.390 335.370 169.710 335.640 ;
        RECT 169.390 335.360 169.700 335.370 ;
        RECT 164.170 335.010 164.410 335.190 ;
        RECT 164.170 334.940 164.470 335.010 ;
        RECT 167.010 335.000 167.420 335.260 ;
        RECT 168.430 335.160 168.630 335.180 ;
        RECT 167.010 334.940 167.480 335.000 ;
        RECT 164.170 322.560 164.410 334.940 ;
        RECT 167.010 334.520 167.420 334.940 ;
        RECT 168.430 334.870 168.780 335.160 ;
        RECT 167.110 334.110 167.420 334.520 ;
        RECT 169.950 334.510 170.260 336.200 ;
        RECT 170.510 335.600 170.790 335.910 ;
        RECT 170.430 335.580 170.790 335.600 ;
        RECT 170.430 335.300 170.750 335.580 ;
        RECT 171.500 335.240 171.790 341.190 ;
        RECT 172.730 340.770 173.200 341.260 ;
        RECT 173.590 341.120 173.960 341.140 ;
        RECT 173.540 340.860 173.960 341.120 ;
        RECT 174.310 340.880 174.550 341.480 ;
        RECT 177.280 341.260 177.540 341.480 ;
        RECT 176.050 341.100 176.390 341.150 ;
        RECT 176.050 341.080 176.610 341.100 ;
        RECT 177.280 341.090 177.930 341.260 ;
        RECT 175.930 340.910 176.610 341.080 ;
        RECT 173.590 340.850 173.960 340.860 ;
        RECT 172.550 340.330 172.870 340.610 ;
        RECT 173.010 340.430 173.200 340.770 ;
        RECT 172.910 340.140 173.200 340.430 ;
        RECT 173.010 339.530 173.200 340.140 ;
        RECT 172.550 339.060 172.870 339.340 ;
        RECT 172.910 339.240 173.200 339.530 ;
        RECT 173.010 338.900 173.200 339.240 ;
        RECT 172.730 338.410 173.200 338.900 ;
        RECT 173.590 338.810 173.960 338.820 ;
        RECT 173.540 338.550 173.960 338.810 ;
        RECT 173.590 338.530 173.960 338.550 ;
        RECT 173.010 338.060 173.200 338.410 ;
        RECT 172.730 337.570 173.200 338.060 ;
        RECT 173.590 337.920 173.960 337.940 ;
        RECT 173.540 337.660 173.960 337.920 ;
        RECT 173.590 337.650 173.960 337.660 ;
        RECT 172.550 337.130 172.870 337.410 ;
        RECT 173.010 337.230 173.200 337.570 ;
        RECT 172.910 336.940 173.200 337.230 ;
        RECT 173.010 336.330 173.200 336.940 ;
        RECT 172.550 335.860 172.870 336.140 ;
        RECT 172.910 336.040 173.200 336.330 ;
        RECT 173.010 335.700 173.200 336.040 ;
        RECT 171.500 334.940 171.830 335.240 ;
        RECT 172.730 335.210 173.200 335.700 ;
        RECT 173.590 335.610 173.960 335.620 ;
        RECT 173.540 335.350 173.960 335.610 ;
        RECT 173.590 335.330 173.960 335.350 ;
        RECT 173.000 334.990 173.200 335.210 ;
        RECT 174.320 334.990 174.550 340.880 ;
        RECT 176.050 340.870 176.610 340.910 ;
        RECT 176.050 340.830 176.390 340.870 ;
        RECT 177.290 340.190 177.930 341.090 ;
        RECT 180.600 341.030 180.760 345.080 ;
        RECT 183.350 341.440 183.590 345.160 ;
        RECT 183.330 341.190 183.720 341.440 ;
        RECT 183.470 340.940 183.720 341.190 ;
        RECT 185.530 340.810 185.910 345.300 ;
        RECT 187.280 341.420 187.520 345.160 ;
        RECT 187.280 341.150 187.750 341.420 ;
        RECT 187.480 340.920 187.750 341.150 ;
        RECT 189.560 340.790 189.960 345.320 ;
        RECT 193.080 342.650 193.320 345.160 ;
        RECT 194.740 344.820 195.010 345.370 ;
        RECT 194.730 344.770 195.010 344.820 ;
        RECT 195.150 345.030 195.340 346.020 ;
        RECT 195.550 345.340 195.710 346.070 ;
        RECT 196.780 345.960 196.940 346.420 ;
        RECT 196.770 345.870 196.940 345.960 ;
        RECT 196.770 345.820 197.050 345.870 ;
        RECT 196.390 345.480 196.710 345.800 ;
        RECT 195.510 345.320 195.710 345.340 ;
        RECT 195.500 345.080 195.730 345.320 ;
        RECT 196.780 345.270 197.050 345.820 ;
        RECT 197.190 345.730 197.350 346.650 ;
        RECT 197.590 346.080 197.750 346.770 ;
        RECT 198.430 346.670 198.750 346.990 ;
        RECT 199.530 346.420 199.770 349.010 ;
        RECT 199.520 346.100 199.780 346.420 ;
        RECT 199.530 346.080 199.770 346.100 ;
        RECT 201.710 346.080 202.090 351.060 ;
        RECT 203.460 349.650 203.700 351.060 ;
        RECT 205.740 350.690 206.140 351.060 ;
        RECT 206.820 350.690 207.220 351.060 ;
        RECT 205.740 350.470 207.220 350.690 ;
        RECT 203.450 348.990 203.710 349.650 ;
        RECT 203.460 346.380 203.700 348.990 ;
        RECT 197.190 345.610 197.360 345.730 ;
        RECT 197.590 345.610 197.860 346.080 ;
        RECT 195.500 345.030 195.710 345.080 ;
        RECT 195.150 344.910 195.320 345.030 ;
        RECT 194.730 344.680 194.900 344.770 ;
        RECT 194.740 344.230 194.900 344.680 ;
        RECT 194.730 344.140 194.900 344.230 ;
        RECT 194.730 344.090 195.010 344.140 ;
        RECT 194.740 343.540 195.010 344.090 ;
        RECT 195.150 344.000 195.310 344.910 ;
        RECT 195.150 343.880 195.320 344.000 ;
        RECT 195.550 343.880 195.710 345.030 ;
        RECT 196.390 344.930 196.710 345.250 ;
        RECT 196.780 344.570 196.940 345.270 ;
        RECT 197.190 344.620 197.380 345.610 ;
        RECT 197.540 345.320 197.860 345.610 ;
        RECT 198.430 345.390 198.750 345.710 ;
        RECT 197.550 345.300 197.860 345.320 ;
        RECT 197.590 344.570 197.860 345.300 ;
        RECT 198.430 344.840 198.750 345.160 ;
        RECT 193.080 342.410 193.660 342.650 ;
        RECT 193.420 341.070 193.660 342.410 ;
        RECT 194.740 342.130 194.900 343.540 ;
        RECT 195.150 342.960 195.340 343.880 ;
        RECT 195.500 343.830 195.710 343.880 ;
        RECT 195.500 343.590 195.730 343.830 ;
        RECT 196.390 343.660 196.710 343.980 ;
        RECT 195.510 343.570 195.710 343.590 ;
        RECT 195.120 342.930 195.360 342.960 ;
        RECT 195.550 342.930 195.710 343.570 ;
        RECT 196.390 343.110 196.710 343.430 ;
        RECT 195.120 342.760 195.710 342.930 ;
        RECT 195.120 342.730 195.360 342.760 ;
        RECT 194.740 341.580 195.010 342.130 ;
        RECT 194.730 341.530 195.010 341.580 ;
        RECT 195.150 341.790 195.340 342.730 ;
        RECT 195.550 342.100 195.710 342.760 ;
        RECT 196.390 342.240 196.710 342.560 ;
        RECT 195.510 342.080 195.710 342.100 ;
        RECT 195.500 341.840 195.730 342.080 ;
        RECT 195.500 341.790 195.710 341.840 ;
        RECT 195.150 341.670 195.320 341.790 ;
        RECT 194.730 341.440 194.900 341.530 ;
        RECT 194.740 340.980 194.900 341.440 ;
        RECT 194.730 340.890 194.900 340.980 ;
        RECT 194.730 340.840 195.010 340.890 ;
        RECT 194.740 340.290 195.010 340.840 ;
        RECT 195.150 340.750 195.310 341.670 ;
        RECT 195.150 340.630 195.320 340.750 ;
        RECT 195.550 340.630 195.710 341.790 ;
        RECT 196.390 341.690 196.710 342.010 ;
        RECT 197.610 341.810 197.860 344.570 ;
        RECT 199.530 344.560 200.050 346.080 ;
        RECT 197.380 341.740 197.540 341.810 ;
        RECT 197.610 341.740 197.980 341.810 ;
        RECT 198.190 341.740 198.350 341.810 ;
        RECT 197.610 341.370 197.860 341.740 ;
        RECT 199.670 341.650 200.050 344.560 ;
        RECT 201.620 344.560 202.090 346.080 ;
        RECT 203.450 346.080 203.710 346.380 ;
        RECT 203.450 346.060 204.100 346.080 ;
        RECT 203.460 344.560 204.100 346.060 ;
        RECT 205.740 344.560 206.140 350.470 ;
        RECT 206.820 344.560 207.220 350.470 ;
        RECT 209.260 349.650 209.500 351.060 ;
        RECT 210.240 351.010 210.610 351.060 ;
        RECT 209.250 348.990 209.510 349.650 ;
        RECT 210.870 349.160 211.380 351.060 ;
        RECT 209.260 346.380 209.500 348.990 ;
        RECT 210.870 348.740 211.390 349.160 ;
        RECT 210.870 348.730 211.380 348.740 ;
        RECT 209.250 346.060 209.510 346.380 ;
        RECT 209.260 344.560 209.500 346.060 ;
        RECT 210.870 344.560 211.250 348.730 ;
        RECT 197.590 341.340 197.870 341.370 ;
        RECT 197.580 341.060 197.880 341.340 ;
        RECT 199.670 341.330 200.160 341.650 ;
        RECT 201.620 341.340 201.890 344.560 ;
        RECT 202.310 341.710 202.690 341.810 ;
        RECT 197.590 341.040 197.870 341.060 ;
        RECT 177.290 339.480 177.540 340.190 ;
        RECT 178.630 339.760 178.950 340.100 ;
        RECT 176.050 338.800 176.390 338.840 ;
        RECT 176.050 338.760 176.610 338.800 ;
        RECT 175.930 338.590 176.610 338.760 ;
        RECT 176.050 338.570 176.610 338.590 ;
        RECT 176.050 338.520 176.390 338.570 ;
        RECT 177.290 338.410 177.930 339.480 ;
        RECT 177.290 338.060 177.540 338.410 ;
        RECT 176.050 337.900 176.390 337.950 ;
        RECT 176.050 337.880 176.610 337.900 ;
        RECT 175.930 337.710 176.610 337.880 ;
        RECT 176.050 337.670 176.610 337.710 ;
        RECT 176.050 337.630 176.390 337.670 ;
        RECT 177.290 336.990 177.930 338.060 ;
        RECT 177.290 336.280 177.540 336.990 ;
        RECT 176.050 335.600 176.390 335.640 ;
        RECT 176.050 335.560 176.610 335.600 ;
        RECT 175.930 335.390 176.610 335.560 ;
        RECT 176.050 335.370 176.610 335.390 ;
        RECT 176.050 335.320 176.390 335.370 ;
        RECT 177.290 335.310 177.930 336.280 ;
        RECT 177.280 335.210 177.930 335.310 ;
        RECT 177.280 334.990 177.540 335.210 ;
        RECT 178.710 335.000 178.920 339.760 ;
        RECT 194.740 339.590 194.900 340.290 ;
        RECT 195.150 339.640 195.340 340.630 ;
        RECT 195.500 340.580 195.710 340.630 ;
        RECT 195.500 340.340 195.730 340.580 ;
        RECT 196.390 340.410 196.710 340.730 ;
        RECT 195.510 340.320 195.710 340.340 ;
        RECT 195.550 339.590 195.710 340.320 ;
        RECT 196.390 340.100 196.710 340.180 ;
        RECT 196.390 339.860 196.870 340.100 ;
        RECT 196.510 339.780 196.870 339.860 ;
        RECT 196.510 339.090 196.720 339.780 ;
        RECT 197.610 339.580 197.860 341.040 ;
        RECT 199.670 340.600 200.050 341.330 ;
        RECT 201.600 341.030 201.910 341.340 ;
        RECT 199.670 340.280 200.140 340.600 ;
        RECT 198.540 340.010 198.800 340.070 ;
        RECT 198.530 339.750 198.800 340.010 ;
        RECT 196.510 338.770 196.850 339.090 ;
        RECT 198.020 338.820 198.280 339.140 ;
        RECT 196.510 338.730 196.720 338.770 ;
        RECT 179.970 338.070 180.360 338.320 ;
        RECT 179.250 336.970 179.590 337.310 ;
        RECT 179.290 336.950 179.510 336.970 ;
        RECT 171.540 334.620 171.830 334.940 ;
        RECT 172.040 334.640 172.380 334.960 ;
        RECT 171.510 334.270 171.860 334.620 ;
        RECT 167.070 333.780 167.440 334.110 ;
        RECT 171.540 333.810 171.830 334.270 ;
        RECT 172.040 334.030 172.290 334.640 ;
        RECT 173.000 334.050 173.190 334.990 ;
        RECT 177.280 334.580 177.530 334.990 ;
        RECT 178.680 334.680 178.960 335.000 ;
        RECT 179.290 334.670 179.490 336.950 ;
        RECT 179.750 335.130 179.940 335.490 ;
        RECT 177.250 334.290 177.590 334.580 ;
        RECT 179.250 334.350 179.530 334.670 ;
        RECT 179.710 334.660 179.990 335.130 ;
        RECT 167.110 332.570 167.420 333.780 ;
        RECT 170.970 333.530 171.830 333.810 ;
        RECT 170.890 333.520 171.830 333.530 ;
        RECT 171.990 333.920 172.290 334.030 ;
        RECT 170.890 333.050 171.350 333.520 ;
        RECT 167.060 332.090 167.480 332.570 ;
        RECT 171.990 332.410 172.180 333.920 ;
        RECT 172.940 333.730 173.260 334.050 ;
        RECT 175.620 333.710 175.880 333.780 ;
        RECT 176.360 333.710 176.620 333.780 ;
        RECT 172.490 333.210 172.810 333.530 ;
        RECT 173.580 333.210 173.900 333.530 ;
        RECT 174.680 333.200 175.000 333.520 ;
        RECT 173.040 332.530 173.360 332.850 ;
        RECT 174.130 332.510 174.450 332.830 ;
        RECT 175.240 332.680 175.560 332.820 ;
        RECT 175.620 332.680 176.620 333.710 ;
        RECT 177.240 333.200 177.560 333.520 ;
        RECT 178.340 333.210 178.660 333.530 ;
        RECT 179.430 333.210 179.750 333.530 ;
        RECT 180.180 333.440 180.360 338.070 ;
        RECT 196.560 336.780 196.880 337.100 ;
        RECT 197.550 336.980 197.810 337.300 ;
        RECT 196.610 335.820 196.930 336.140 ;
        RECT 197.050 336.050 197.310 336.370 ;
        RECT 181.500 334.600 181.760 334.630 ;
        RECT 181.480 334.300 181.780 334.600 ;
        RECT 181.500 334.290 181.760 334.300 ;
        RECT 180.180 333.140 180.660 333.440 ;
        RECT 181.510 333.370 181.730 334.290 ;
        RECT 183.470 334.160 183.720 335.390 ;
        RECT 187.480 334.180 187.750 335.410 ;
        RECT 190.300 334.610 190.730 335.010 ;
        RECT 183.460 333.900 183.780 334.160 ;
        RECT 187.480 333.870 187.830 334.180 ;
        RECT 185.430 333.630 185.690 333.810 ;
        RECT 186.170 333.630 186.430 333.810 ;
        RECT 180.260 333.030 180.660 333.140 ;
        RECT 181.450 332.970 181.790 333.370 ;
        RECT 182.300 333.240 182.620 333.560 ;
        RECT 183.390 333.240 183.710 333.560 ;
        RECT 184.490 333.230 184.810 333.550 ;
        RECT 181.510 332.890 181.730 332.970 ;
        RECT 176.680 332.680 177.000 332.820 ;
        RECT 175.240 332.500 175.880 332.680 ;
        RECT 171.550 332.090 172.180 332.410 ;
        RECT 175.380 332.360 175.880 332.500 ;
        RECT 171.550 331.990 171.990 332.090 ;
        RECT 173.040 331.160 173.360 331.480 ;
        RECT 174.130 331.160 174.450 331.480 ;
        RECT 175.230 331.340 175.550 331.480 ;
        RECT 175.620 331.340 175.880 332.360 ;
        RECT 175.230 331.160 175.880 331.340 ;
        RECT 175.380 331.020 175.880 331.160 ;
        RECT 172.480 330.430 172.800 330.750 ;
        RECT 173.580 330.430 173.900 330.750 ;
        RECT 174.680 330.430 175.000 330.750 ;
        RECT 172.480 329.060 172.800 329.380 ;
        RECT 173.580 329.060 173.900 329.380 ;
        RECT 174.680 329.060 175.000 329.380 ;
        RECT 171.910 328.560 172.230 328.740 ;
        RECT 171.760 328.420 172.230 328.560 ;
        RECT 171.760 328.270 172.080 328.420 ;
        RECT 173.040 328.380 173.360 328.700 ;
        RECT 174.130 328.380 174.450 328.700 ;
        RECT 175.230 328.570 175.550 328.710 ;
        RECT 175.620 328.570 175.880 331.020 ;
        RECT 175.230 328.390 175.880 328.570 ;
        RECT 171.760 327.950 172.240 328.270 ;
        RECT 175.380 328.250 175.880 328.390 ;
        RECT 171.760 326.810 172.080 327.950 ;
        RECT 175.620 327.590 175.880 328.250 ;
        RECT 176.360 332.500 177.000 332.680 ;
        RECT 177.790 332.510 178.110 332.830 ;
        RECT 178.880 332.530 179.200 332.850 ;
        RECT 182.850 332.560 183.170 332.880 ;
        RECT 183.940 332.540 184.260 332.860 ;
        RECT 185.050 332.700 185.370 332.850 ;
        RECT 185.430 332.700 186.430 333.630 ;
        RECT 187.050 333.230 187.370 333.550 ;
        RECT 188.150 333.240 188.470 333.560 ;
        RECT 189.240 333.240 189.560 333.560 ;
        RECT 186.490 332.700 186.810 332.850 ;
        RECT 185.050 332.530 185.690 332.700 ;
        RECT 176.360 332.360 176.860 332.500 ;
        RECT 185.190 332.380 185.690 332.530 ;
        RECT 176.360 331.330 176.620 332.360 ;
        RECT 176.690 331.330 177.010 331.480 ;
        RECT 176.360 331.160 177.010 331.330 ;
        RECT 177.790 331.160 178.110 331.480 ;
        RECT 178.880 331.160 179.200 331.480 ;
        RECT 182.850 331.190 183.170 331.510 ;
        RECT 183.940 331.190 184.260 331.510 ;
        RECT 185.040 331.360 185.360 331.510 ;
        RECT 185.430 331.360 185.690 332.380 ;
        RECT 185.040 331.190 185.690 331.360 ;
        RECT 176.360 331.010 176.860 331.160 ;
        RECT 185.190 331.040 185.690 331.190 ;
        RECT 176.360 328.560 176.620 331.010 ;
        RECT 177.240 330.430 177.560 330.750 ;
        RECT 178.340 330.430 178.660 330.750 ;
        RECT 179.440 330.430 179.760 330.750 ;
        RECT 182.290 330.460 182.610 330.780 ;
        RECT 183.390 330.460 183.710 330.780 ;
        RECT 184.490 330.460 184.810 330.780 ;
        RECT 177.240 329.060 177.560 329.380 ;
        RECT 178.340 329.060 178.660 329.380 ;
        RECT 179.440 329.060 179.760 329.380 ;
        RECT 182.290 329.090 182.610 329.410 ;
        RECT 183.390 329.090 183.710 329.410 ;
        RECT 184.490 329.090 184.810 329.410 ;
        RECT 176.690 328.560 177.010 328.710 ;
        RECT 176.360 328.390 177.010 328.560 ;
        RECT 176.360 328.240 176.860 328.390 ;
        RECT 177.790 328.380 178.110 328.700 ;
        RECT 178.880 328.380 179.200 328.700 ;
        RECT 180.010 328.580 180.330 328.740 ;
        RECT 180.010 328.420 180.470 328.580 ;
        RECT 181.720 328.570 182.040 328.770 ;
        RECT 180.130 328.270 180.470 328.420 ;
        RECT 176.360 327.610 176.620 328.240 ;
        RECT 180.000 327.950 180.470 328.270 ;
        RECT 175.610 327.250 175.890 327.590 ;
        RECT 176.350 327.270 176.630 327.610 ;
        RECT 171.640 326.210 172.180 326.810 ;
        RECT 175.620 325.840 175.880 327.250 ;
        RECT 176.360 325.840 176.620 327.270 ;
        RECT 163.770 321.240 164.420 322.560 ;
        RECT 175.620 322.410 176.620 325.840 ;
        RECT 180.130 325.790 180.470 327.950 ;
        RECT 181.560 328.450 182.040 328.570 ;
        RECT 181.560 328.300 181.900 328.450 ;
        RECT 182.850 328.410 183.170 328.730 ;
        RECT 183.940 328.410 184.260 328.730 ;
        RECT 185.040 328.590 185.360 328.740 ;
        RECT 185.430 328.590 185.690 331.040 ;
        RECT 185.040 328.420 185.690 328.590 ;
        RECT 181.560 327.980 182.050 328.300 ;
        RECT 185.190 328.270 185.690 328.420 ;
        RECT 180.070 325.270 180.530 325.790 ;
        RECT 181.560 324.900 181.900 327.980 ;
        RECT 185.430 327.590 185.690 328.270 ;
        RECT 186.170 332.530 186.810 332.700 ;
        RECT 187.600 332.540 187.920 332.860 ;
        RECT 188.690 332.560 189.010 332.880 ;
        RECT 190.340 332.820 190.690 334.610 ;
        RECT 192.160 334.050 192.380 335.370 ;
        RECT 193.420 334.650 193.650 335.370 ;
        RECT 193.420 334.420 196.630 334.650 ;
        RECT 193.420 334.410 193.650 334.420 ;
        RECT 191.870 333.810 192.380 334.050 ;
        RECT 191.870 332.560 192.100 333.810 ;
        RECT 196.400 333.450 196.630 334.420 ;
        RECT 196.350 333.050 196.660 333.450 ;
        RECT 186.170 332.380 186.670 332.530 ;
        RECT 186.170 331.350 186.430 332.380 ;
        RECT 191.760 332.120 192.220 332.560 ;
        RECT 186.500 331.350 186.820 331.510 ;
        RECT 186.170 331.190 186.820 331.350 ;
        RECT 187.600 331.190 187.920 331.510 ;
        RECT 188.690 331.190 189.010 331.510 ;
        RECT 186.170 331.030 186.670 331.190 ;
        RECT 186.170 328.590 186.430 331.030 ;
        RECT 187.050 330.460 187.370 330.780 ;
        RECT 188.150 330.460 188.470 330.780 ;
        RECT 189.250 330.460 189.570 330.780 ;
        RECT 196.400 329.880 196.630 333.050 ;
        RECT 196.270 329.660 196.630 329.880 ;
        RECT 196.070 329.430 196.630 329.660 ;
        RECT 196.070 329.420 196.610 329.430 ;
        RECT 187.050 329.090 187.370 329.410 ;
        RECT 188.150 329.090 188.470 329.410 ;
        RECT 189.250 329.090 189.570 329.410 ;
        RECT 193.430 329.020 193.750 329.340 ;
        RECT 194.530 329.030 194.850 329.350 ;
        RECT 195.620 329.030 195.940 329.350 ;
        RECT 186.500 328.590 186.820 328.740 ;
        RECT 186.170 328.420 186.820 328.590 ;
        RECT 186.170 328.270 186.670 328.420 ;
        RECT 187.600 328.410 187.920 328.730 ;
        RECT 188.690 328.410 189.010 328.730 ;
        RECT 189.820 328.610 190.140 328.770 ;
        RECT 189.820 328.450 190.250 328.610 ;
        RECT 189.980 328.300 190.250 328.450 ;
        RECT 192.870 328.320 193.190 328.640 ;
        RECT 193.980 328.330 194.300 328.650 ;
        RECT 195.070 328.350 195.390 328.670 ;
        RECT 185.420 327.250 185.700 327.590 ;
        RECT 185.430 326.070 185.690 327.250 ;
        RECT 186.170 326.070 186.430 328.270 ;
        RECT 189.810 327.980 190.250 328.300 ;
        RECT 197.050 328.210 197.300 336.050 ;
        RECT 197.550 329.110 197.800 336.980 ;
        RECT 198.030 330.020 198.280 338.820 ;
        RECT 198.530 330.910 198.780 339.750 ;
        RECT 199.670 339.580 200.050 340.280 ;
        RECT 201.620 339.580 201.890 341.030 ;
        RECT 203.700 339.580 204.100 344.560 ;
        RECT 211.890 343.990 212.260 365.780 ;
        RECT 214.200 364.010 214.870 366.870 ;
        RECT 214.100 363.720 214.870 364.010 ;
        RECT 212.320 362.890 212.530 363.000 ;
        RECT 212.790 362.920 212.980 363.000 ;
        RECT 213.200 362.940 213.410 363.000 ;
        RECT 214.200 360.840 214.870 363.720 ;
        RECT 212.970 359.630 213.200 360.840 ;
        RECT 214.190 359.940 214.870 360.840 ;
        RECT 214.190 359.870 215.170 359.940 ;
        RECT 212.940 358.840 213.200 359.630 ;
        RECT 214.180 359.620 215.170 359.870 ;
        RECT 212.330 356.960 212.560 357.080 ;
        RECT 212.970 356.690 213.200 358.840 ;
        RECT 214.190 357.980 214.870 359.620 ;
        RECT 214.090 357.690 214.870 357.980 ;
        RECT 212.940 355.900 213.200 356.690 ;
        RECT 212.970 354.790 213.200 355.900 ;
        RECT 214.190 354.790 214.870 357.690 ;
        RECT 214.880 355.930 215.200 356.250 ;
        RECT 213.190 349.670 213.430 351.060 ;
        RECT 214.370 350.780 214.870 354.790 ;
        RECT 215.300 351.050 215.800 368.730 ;
        RECT 216.430 356.960 216.930 369.190 ;
        RECT 216.430 356.880 217.160 356.960 ;
        RECT 214.210 350.460 214.870 350.780 ;
        RECT 214.370 350.230 214.870 350.460 ;
        RECT 215.210 350.300 215.800 351.050 ;
        RECT 216.020 350.940 216.180 351.050 ;
        RECT 216.020 350.660 216.350 350.940 ;
        RECT 216.020 350.350 216.180 350.660 ;
        RECT 214.210 349.910 214.870 350.230 ;
        RECT 215.190 350.060 215.800 350.300 ;
        RECT 213.170 349.010 213.440 349.670 ;
        RECT 213.190 346.420 213.430 349.010 ;
        RECT 214.370 348.940 214.870 349.910 ;
        RECT 214.210 348.620 214.870 348.940 ;
        RECT 215.210 348.790 215.800 350.060 ;
        RECT 215.910 349.800 216.180 350.350 ;
        RECT 215.910 349.750 216.190 349.800 ;
        RECT 216.020 349.660 216.190 349.750 ;
        RECT 216.020 349.190 216.180 349.660 ;
        RECT 216.020 349.100 216.190 349.190 ;
        RECT 214.370 348.390 214.870 348.620 ;
        RECT 215.190 348.550 215.800 348.790 ;
        RECT 214.210 348.070 214.870 348.390 ;
        RECT 214.370 347.540 214.870 348.070 ;
        RECT 214.210 347.220 214.870 347.540 ;
        RECT 214.370 346.990 214.870 347.220 ;
        RECT 215.210 347.060 215.800 348.550 ;
        RECT 215.910 349.050 216.190 349.100 ;
        RECT 215.910 348.500 216.180 349.050 ;
        RECT 216.020 347.110 216.180 348.500 ;
        RECT 214.210 346.670 214.870 346.990 ;
        RECT 215.190 346.820 215.800 347.060 ;
        RECT 213.180 346.100 213.440 346.420 ;
        RECT 213.190 344.560 213.430 346.100 ;
        RECT 214.370 345.710 214.870 346.670 ;
        RECT 214.210 345.390 214.870 345.710 ;
        RECT 215.210 345.560 215.800 346.820 ;
        RECT 215.910 346.560 216.180 347.110 ;
        RECT 215.910 346.510 216.190 346.560 ;
        RECT 216.020 346.420 216.190 346.510 ;
        RECT 216.020 345.960 216.180 346.420 ;
        RECT 216.020 345.870 216.190 345.960 ;
        RECT 214.370 345.160 214.870 345.390 ;
        RECT 215.190 345.320 215.800 345.560 ;
        RECT 214.210 344.840 214.870 345.160 ;
        RECT 211.850 343.480 212.340 343.990 ;
        RECT 211.890 343.450 212.260 343.480 ;
        RECT 206.340 341.530 206.740 341.810 ;
        RECT 208.000 340.880 208.320 341.200 ;
        RECT 208.150 340.200 208.470 340.520 ;
        RECT 208.150 339.610 208.470 339.930 ;
        RECT 208.000 338.930 208.320 339.250 ;
        RECT 199.880 338.620 200.140 338.720 ;
        RECT 199.790 338.400 200.140 338.620 ;
        RECT 199.790 337.540 199.950 338.400 ;
        RECT 208.000 338.110 208.320 338.430 ;
        RECT 199.750 337.220 200.010 337.540 ;
        RECT 208.150 337.430 208.470 337.750 ;
        RECT 199.790 337.120 199.950 337.220 ;
        RECT 208.150 336.840 208.470 337.160 ;
        RECT 208.000 336.160 208.320 336.480 ;
        RECT 202.310 335.760 202.690 335.860 ;
        RECT 208.940 335.760 209.170 341.810 ;
        RECT 210.200 337.460 210.430 341.810 ;
        RECT 210.160 337.450 210.440 337.460 ;
        RECT 210.160 337.130 210.460 337.450 ;
        RECT 210.200 335.760 210.430 337.130 ;
        RECT 214.370 332.410 214.870 344.840 ;
        RECT 215.210 344.570 215.800 345.320 ;
        RECT 215.910 345.820 216.190 345.870 ;
        RECT 215.910 345.270 216.180 345.820 ;
        RECT 216.020 344.570 216.180 345.270 ;
        RECT 215.300 337.690 215.800 344.570 ;
        RECT 216.430 342.920 216.930 356.880 ;
        RECT 217.560 348.090 218.060 369.810 ;
        RECT 226.420 368.210 227.700 372.480 ;
        RECT 226.410 366.870 227.700 368.210 ;
        RECT 220.440 362.850 220.860 363.000 ;
        RECT 221.470 362.850 221.890 363.000 ;
        RECT 225.170 362.920 225.400 363.000 ;
        RECT 220.440 362.710 221.890 362.850 ;
        RECT 225.430 360.840 225.850 366.870 ;
        RECT 226.420 366.380 227.700 366.870 ;
        RECT 227.910 364.010 228.140 366.870 ;
        RECT 229.130 365.660 229.360 366.870 ;
        RECT 229.130 364.870 229.390 365.660 ;
        RECT 234.290 365.560 234.480 379.600 ;
        RECT 240.600 379.060 241.220 382.480 ;
        RECT 240.600 379.050 241.170 379.060 ;
        RECT 239.770 377.420 240.330 377.920 ;
        RECT 243.600 377.500 244.320 383.170 ;
        RECT 245.070 383.900 259.360 384.460 ;
        RECT 270.290 384.290 270.820 385.190 ;
        RECT 271.930 385.130 274.300 385.760 ;
        RECT 245.070 379.600 268.420 383.900 ;
        RECT 271.960 383.170 272.910 385.130 ;
        RECT 273.660 385.110 274.240 385.130 ;
        RECT 284.040 384.470 287.950 385.930 ;
        RECT 295.270 385.280 299.400 385.680 ;
        RECT 295.270 385.190 299.410 385.280 ;
        RECT 274.330 384.460 287.950 384.470 ;
        RECT 269.190 382.480 269.760 382.490 ;
        RECT 245.070 379.320 259.360 379.600 ;
        RECT 255.450 377.770 259.360 379.320 ;
        RECT 269.190 379.060 269.810 382.480 ;
        RECT 269.190 379.050 269.760 379.060 ;
        RECT 239.780 377.200 240.330 377.420 ;
        RECT 236.450 376.090 236.640 376.100 ;
        RECT 243.580 376.090 244.300 377.460 ;
        RECT 255.430 376.230 259.380 377.770 ;
        RECT 268.360 377.420 268.920 377.920 ;
        RECT 272.190 377.500 272.910 383.170 ;
        RECT 273.660 383.900 287.950 384.460 ;
        RECT 298.880 384.290 299.410 385.190 ;
        RECT 300.520 385.130 302.890 385.760 ;
        RECT 273.660 379.600 297.010 383.900 ;
        RECT 300.550 383.170 301.500 385.130 ;
        RECT 302.250 385.110 302.830 385.130 ;
        RECT 312.630 384.470 316.540 385.930 ;
        RECT 323.860 385.280 327.990 385.680 ;
        RECT 323.860 385.190 328.000 385.280 ;
        RECT 302.920 384.460 316.540 384.470 ;
        RECT 297.780 382.480 298.350 382.490 ;
        RECT 273.660 379.320 287.950 379.600 ;
        RECT 284.040 377.770 287.950 379.320 ;
        RECT 297.780 379.060 298.400 382.480 ;
        RECT 297.780 379.050 298.350 379.060 ;
        RECT 268.370 377.200 268.920 377.420 ;
        RECT 284.020 377.000 287.970 377.770 ;
        RECT 296.950 377.420 297.510 377.920 ;
        RECT 300.780 377.500 301.500 383.170 ;
        RECT 302.250 383.900 316.540 384.460 ;
        RECT 327.470 384.290 328.000 385.190 ;
        RECT 329.110 385.130 331.480 385.760 ;
        RECT 302.250 379.600 325.600 383.900 ;
        RECT 329.140 383.170 330.090 385.130 ;
        RECT 330.840 385.110 331.420 385.130 ;
        RECT 341.220 384.470 345.130 385.930 ;
        RECT 352.450 385.280 356.580 385.680 ;
        RECT 352.450 385.190 356.590 385.280 ;
        RECT 331.510 384.460 345.130 384.470 ;
        RECT 326.370 382.480 326.940 382.490 ;
        RECT 302.250 379.320 316.540 379.600 ;
        RECT 312.630 377.770 316.540 379.320 ;
        RECT 326.370 379.060 326.990 382.480 ;
        RECT 326.370 379.050 326.940 379.060 ;
        RECT 296.960 377.200 297.510 377.420 ;
        RECT 284.030 376.230 287.980 377.000 ;
        RECT 312.610 376.230 316.560 377.770 ;
        RECT 325.540 377.420 326.100 377.920 ;
        RECT 329.370 377.500 330.090 383.170 ;
        RECT 330.840 383.900 345.130 384.460 ;
        RECT 356.060 384.290 356.590 385.190 ;
        RECT 330.840 379.600 354.190 383.900 ;
        RECT 354.960 382.480 355.530 382.490 ;
        RECT 330.840 379.320 345.130 379.600 ;
        RECT 341.220 377.770 345.130 379.320 ;
        RECT 354.960 379.060 355.580 382.480 ;
        RECT 354.960 379.050 355.530 379.060 ;
        RECT 325.550 377.200 326.100 377.420 ;
        RECT 341.200 376.230 345.150 377.770 ;
        RECT 354.130 377.420 354.690 377.920 ;
        RECT 354.140 377.200 354.690 377.420 ;
        RECT 236.450 375.740 244.300 376.090 ;
        RECT 236.450 373.610 236.640 375.740 ;
        RECT 256.110 375.550 259.340 376.230 ;
        RECT 255.350 375.270 259.340 375.550 ;
        RECT 255.330 375.070 259.340 375.270 ;
        RECT 237.630 372.880 238.450 372.970 ;
        RECT 237.570 372.190 238.450 372.880 ;
        RECT 235.650 366.830 235.840 366.870 ;
        RECT 234.290 365.450 234.740 365.560 ;
        RECT 234.290 365.380 234.900 365.450 ;
        RECT 234.150 365.280 234.900 365.380 ;
        RECT 234.050 365.240 234.900 365.280 ;
        RECT 230.780 365.200 230.980 365.230 ;
        RECT 226.870 363.430 227.220 363.910 ;
        RECT 227.910 363.720 228.240 364.010 ;
        RECT 225.420 360.820 225.850 360.840 ;
        RECT 222.880 360.230 223.350 360.720 ;
        RECT 218.100 357.000 218.420 357.300 ;
        RECT 218.150 356.880 218.380 356.960 ;
        RECT 220.440 356.810 221.880 356.970 ;
        RECT 218.180 354.150 218.350 354.330 ;
        RECT 218.160 353.560 218.480 353.860 ;
        RECT 218.160 353.450 218.400 353.560 ;
        RECT 218.190 353.440 218.360 353.450 ;
        RECT 218.380 353.390 218.400 353.450 ;
        RECT 221.310 351.530 221.700 353.390 ;
        RECT 217.510 347.530 218.060 348.090 ;
        RECT 216.420 342.360 216.940 342.920 ;
        RECT 215.290 337.170 215.810 337.690 ;
        RECT 214.210 331.840 214.870 332.410 ;
        RECT 198.480 330.330 198.850 330.910 ;
        RECT 197.950 329.440 198.320 330.020 ;
        RECT 197.460 328.530 197.830 329.110 ;
        RECT 181.470 324.380 181.990 324.900 ;
        RECT 185.430 322.470 186.430 326.070 ;
        RECT 189.980 324.020 190.250 327.980 ;
        RECT 192.880 326.980 193.200 327.300 ;
        RECT 193.980 326.980 194.300 327.300 ;
        RECT 195.070 326.980 195.390 327.300 ;
        RECT 195.720 326.570 196.050 327.990 ;
        RECT 196.990 327.640 197.340 328.210 ;
        RECT 193.430 326.250 193.750 326.570 ;
        RECT 194.530 326.250 194.850 326.570 ;
        RECT 195.630 326.250 196.050 326.570 ;
        RECT 195.720 325.200 196.050 326.250 ;
        RECT 196.500 326.070 196.770 326.100 ;
        RECT 196.490 325.540 196.770 326.070 ;
        RECT 196.490 325.240 196.950 325.540 ;
        RECT 193.430 324.880 193.750 325.200 ;
        RECT 194.530 324.880 194.850 325.200 ;
        RECT 195.630 324.880 196.050 325.200 ;
        RECT 192.880 324.210 193.200 324.530 ;
        RECT 193.980 324.200 194.300 324.520 ;
        RECT 195.070 324.200 195.390 324.520 ;
        RECT 189.870 323.460 190.360 324.020 ;
        RECT 185.430 322.430 187.450 322.470 ;
        RECT 175.140 322.370 177.070 322.410 ;
        RECT 174.600 321.180 177.070 322.370 ;
        RECT 162.120 316.950 162.490 317.330 ;
        RECT 161.470 316.330 161.860 316.720 ;
        RECT 160.870 315.700 161.250 316.090 ;
        RECT 160.280 315.070 160.630 315.440 ;
        RECT 159.640 314.390 160.000 314.770 ;
        RECT 159.050 314.150 159.390 314.160 ;
        RECT 159.030 313.780 159.410 314.150 ;
        RECT 159.050 313.770 159.380 313.780 ;
        RECT 157.270 311.930 157.620 312.260 ;
        RECT 157.290 311.870 157.620 311.930 ;
        RECT 156.000 310.650 156.350 310.980 ;
        RECT 156.000 310.580 156.330 310.650 ;
        RECT 153.860 309.920 155.100 310.250 ;
        RECT 155.390 309.950 155.830 310.370 ;
        RECT 153.860 309.810 154.440 309.920 ;
        RECT 174.600 309.690 175.540 321.180 ;
        RECT 184.950 321.150 187.450 322.430 ;
        RECT 186.560 311.150 187.450 321.150 ;
        RECT 195.720 318.000 196.050 324.880 ;
        RECT 196.480 325.220 196.950 325.240 ;
        RECT 196.480 324.790 196.770 325.220 ;
        RECT 196.200 324.240 196.520 324.560 ;
        RECT 196.190 323.770 196.510 324.090 ;
        RECT 214.370 323.530 214.870 331.840 ;
        RECT 215.300 324.440 215.800 337.170 ;
        RECT 216.430 325.310 216.930 342.360 ;
        RECT 217.560 326.820 218.060 347.530 ;
        RECT 220.450 334.380 221.030 334.940 ;
        RECT 220.480 334.370 220.990 334.380 ;
        RECT 217.560 326.260 218.120 326.820 ;
        RECT 217.560 326.130 218.060 326.260 ;
        RECT 220.480 322.500 220.980 334.370 ;
        RECT 219.850 321.220 220.980 322.500 ;
        RECT 195.660 317.610 196.090 318.000 ;
        RECT 222.930 316.880 223.330 360.230 ;
        RECT 223.850 359.620 224.270 359.980 ;
        RECT 222.920 316.420 223.390 316.880 ;
        RECT 223.860 316.080 224.250 359.620 ;
        RECT 224.770 357.230 225.220 357.660 ;
        RECT 224.790 356.970 225.180 357.230 ;
        RECT 225.420 356.980 225.840 360.820 ;
        RECT 225.420 356.970 226.010 356.980 ;
        RECT 224.790 356.890 225.390 356.970 ;
        RECT 223.830 315.610 224.290 316.080 ;
        RECT 224.790 315.260 225.180 356.890 ;
        RECT 225.420 356.670 226.030 356.970 ;
        RECT 225.420 354.790 226.010 356.670 ;
        RECT 225.630 353.320 226.010 354.790 ;
        RECT 225.340 351.460 226.010 353.320 ;
        RECT 224.770 314.800 225.240 315.260 ;
        RECT 225.630 314.460 226.010 351.460 ;
        RECT 226.970 333.440 227.200 363.430 ;
        RECT 227.910 360.840 228.140 363.720 ;
        RECT 229.130 362.720 229.360 364.870 ;
        RECT 230.690 364.700 231.000 365.200 ;
        RECT 234.050 364.960 234.480 365.240 ;
        RECT 229.130 361.930 229.390 362.720 ;
        RECT 229.130 360.840 229.360 361.930 ;
        RECT 230.780 361.450 230.980 364.700 ;
        RECT 234.230 364.550 234.480 364.960 ;
        RECT 234.710 365.170 234.900 365.240 ;
        RECT 234.710 364.880 235.020 365.170 ;
        RECT 233.810 364.190 234.130 364.510 ;
        RECT 234.230 364.460 234.560 364.550 ;
        RECT 234.290 364.260 234.560 364.460 ;
        RECT 233.360 363.630 233.580 363.790 ;
        RECT 233.360 363.570 233.700 363.630 ;
        RECT 233.350 363.310 233.700 363.570 ;
        RECT 233.770 363.360 233.970 363.680 ;
        RECT 231.140 363.250 231.340 363.290 ;
        RECT 233.350 363.280 233.580 363.310 ;
        RECT 233.770 363.070 234.090 363.360 ;
        RECT 231.690 362.920 231.880 363.000 ;
        RECT 232.130 362.980 232.410 363.000 ;
        RECT 232.130 362.920 232.470 362.980 ;
        RECT 232.150 362.680 232.470 362.920 ;
        RECT 233.770 362.070 233.970 363.070 ;
        RECT 234.290 362.800 234.480 364.260 ;
        RECT 234.710 363.930 234.900 364.880 ;
        RECT 235.340 364.080 235.600 364.400 ;
        RECT 236.090 364.120 236.370 366.870 ;
        RECT 236.090 363.800 236.540 364.120 ;
        RECT 235.340 363.480 235.600 363.800 ;
        RECT 234.650 363.230 234.840 363.290 ;
        RECT 235.710 363.260 235.970 363.560 ;
        RECT 235.690 363.240 235.970 363.260 ;
        RECT 235.690 363.000 235.880 363.240 ;
        RECT 236.090 363.000 236.370 363.800 ;
        RECT 237.280 363.640 237.470 363.680 ;
        RECT 236.720 363.000 237.040 363.140 ;
        RECT 237.570 363.120 238.280 372.190 ;
        RECT 255.150 371.370 259.500 375.070 ;
        RECT 284.700 370.890 287.930 376.230 ;
        RECT 239.940 366.950 240.330 370.540 ;
        RECT 238.890 366.470 239.200 366.910 ;
        RECT 240.410 365.830 240.600 367.280 ;
        RECT 240.850 366.640 241.010 367.280 ;
        RECT 284.400 366.840 287.950 370.890 ;
        RECT 240.740 366.090 241.010 366.640 ;
        RECT 240.740 366.040 241.020 366.090 ;
        RECT 240.850 365.950 241.020 366.040 ;
        RECT 240.410 365.800 240.630 365.830 ;
        RECT 240.390 365.530 240.640 365.800 ;
        RECT 240.400 365.520 240.640 365.530 ;
        RECT 240.400 365.280 240.630 365.520 ;
        RECT 240.010 364.510 240.250 364.850 ;
        RECT 235.690 362.860 236.370 363.000 ;
        RECT 234.290 362.480 234.740 362.800 ;
        RECT 235.690 362.750 235.880 362.860 ;
        RECT 234.290 362.180 234.480 362.480 ;
        RECT 234.810 362.380 235.130 362.700 ;
        RECT 235.690 362.670 236.000 362.750 ;
        RECT 235.670 362.460 236.000 362.670 ;
        RECT 235.670 362.380 235.900 362.460 ;
        RECT 234.150 362.080 234.480 362.180 ;
        RECT 234.050 361.760 234.480 362.080 ;
        RECT 227.900 360.820 228.140 360.840 ;
        RECT 229.120 360.820 229.360 360.840 ;
        RECT 233.770 361.310 233.970 361.560 ;
        RECT 234.230 361.460 234.480 361.760 ;
        RECT 234.710 361.970 234.900 362.250 ;
        RECT 234.710 361.680 235.020 361.970 ;
        RECT 234.230 361.350 234.420 361.460 ;
        RECT 233.770 360.990 234.130 361.310 ;
        RECT 234.230 361.260 234.560 361.350 ;
        RECT 234.330 361.060 234.560 361.260 ;
        RECT 234.710 361.250 234.900 361.680 ;
        RECT 227.900 357.980 228.130 360.820 ;
        RECT 229.120 359.630 229.350 360.820 ;
        RECT 233.360 360.430 233.580 360.590 ;
        RECT 233.770 360.560 233.970 360.990 ;
        RECT 234.710 360.930 235.130 361.250 ;
        RECT 235.670 361.170 235.900 361.250 ;
        RECT 235.670 360.960 236.000 361.170 ;
        RECT 234.710 360.730 234.900 360.930 ;
        RECT 235.690 360.880 236.000 360.960 ;
        RECT 235.690 360.870 235.880 360.880 ;
        RECT 235.650 360.840 235.880 360.870 ;
        RECT 236.090 360.840 236.370 362.860 ;
        RECT 236.480 362.850 237.040 363.000 ;
        RECT 236.720 362.820 237.040 362.850 ;
        RECT 237.540 363.110 238.280 363.120 ;
        RECT 236.670 362.170 236.990 362.490 ;
        RECT 237.280 362.070 237.470 362.120 ;
        RECT 237.540 361.760 238.480 363.110 ;
        RECT 238.970 362.840 239.290 363.160 ;
        RECT 237.280 361.510 237.470 361.560 ;
        RECT 237.540 361.470 238.590 361.760 ;
        RECT 236.670 361.020 236.990 361.340 ;
        RECT 235.640 360.800 235.880 360.840 ;
        RECT 233.360 360.370 233.700 360.430 ;
        RECT 233.350 360.060 233.700 360.370 ;
        RECT 233.360 360.000 233.700 360.060 ;
        RECT 233.770 360.270 234.090 360.560 ;
        RECT 235.690 360.390 235.880 360.800 ;
        RECT 236.080 360.820 236.370 360.840 ;
        RECT 235.690 360.370 235.970 360.390 ;
        RECT 233.770 360.160 233.970 360.270 ;
        RECT 233.360 359.840 233.580 360.000 ;
        RECT 233.770 359.870 234.090 360.160 ;
        RECT 235.710 360.060 235.970 360.370 ;
        RECT 235.690 360.040 235.970 360.060 ;
        RECT 229.120 358.840 229.380 359.630 ;
        RECT 233.770 359.440 233.970 359.870 ;
        RECT 234.710 359.530 234.900 359.700 ;
        RECT 234.410 359.500 234.900 359.530 ;
        RECT 235.690 359.550 235.880 360.040 ;
        RECT 233.770 359.120 234.130 359.440 ;
        RECT 234.410 359.370 235.130 359.500 ;
        RECT 235.690 359.470 236.000 359.550 ;
        RECT 234.330 359.210 235.130 359.370 ;
        RECT 234.330 359.170 234.560 359.210 ;
        RECT 233.770 358.870 233.970 359.120 ;
        RECT 234.230 359.080 234.560 359.170 ;
        RECT 234.710 359.180 235.130 359.210 ;
        RECT 235.670 359.260 236.000 359.470 ;
        RECT 235.670 359.180 235.900 359.260 ;
        RECT 227.900 357.690 228.230 357.980 ;
        RECT 227.900 354.790 228.130 357.690 ;
        RECT 229.120 356.690 229.350 358.840 ;
        RECT 234.230 358.670 234.420 359.080 ;
        RECT 232.410 358.270 232.730 358.590 ;
        RECT 234.050 358.420 234.420 358.670 ;
        RECT 234.710 358.750 234.900 359.180 ;
        RECT 234.710 358.460 235.020 358.750 ;
        RECT 232.560 357.440 232.880 357.760 ;
        RECT 233.770 357.360 233.970 358.360 ;
        RECT 234.050 358.350 234.410 358.420 ;
        RECT 234.150 358.250 234.410 358.350 ;
        RECT 234.710 358.180 234.900 358.460 ;
        RECT 235.330 358.050 235.590 358.370 ;
        RECT 236.080 358.090 236.360 360.820 ;
        RECT 236.720 360.370 237.040 360.690 ;
        RECT 237.280 360.440 237.470 360.480 ;
        RECT 236.720 359.820 237.040 360.140 ;
        RECT 237.280 359.950 237.470 359.990 ;
        RECT 236.670 359.170 236.990 359.490 ;
        RECT 237.540 359.170 238.480 361.470 ;
        RECT 238.890 360.940 239.200 361.220 ;
        RECT 238.890 360.880 239.340 360.940 ;
        RECT 239.930 360.920 240.320 364.510 ;
        RECT 240.440 364.260 240.600 365.280 ;
        RECT 240.850 364.260 241.010 365.950 ;
        RECT 313.290 365.260 316.520 376.230 ;
        RECT 240.440 362.410 240.600 363.430 ;
        RECT 240.400 362.170 240.630 362.410 ;
        RECT 240.400 362.160 240.640 362.170 ;
        RECT 240.390 361.890 240.640 362.160 ;
        RECT 240.410 361.860 240.630 361.890 ;
        RECT 240.410 361.250 240.600 361.860 ;
        RECT 240.850 361.740 241.010 363.430 ;
        RECT 313.090 362.730 316.680 365.260 ;
        RECT 341.880 361.770 345.110 376.230 ;
        RECT 240.850 361.650 241.020 361.740 ;
        RECT 238.880 360.620 239.340 360.880 ;
        RECT 238.880 360.440 239.190 360.620 ;
        RECT 240.400 360.410 240.600 361.250 ;
        RECT 240.740 361.600 241.020 361.650 ;
        RECT 240.740 361.050 241.010 361.600 ;
        RECT 240.840 360.610 241.010 361.050 ;
        RECT 240.730 360.410 241.010 360.610 ;
        RECT 239.010 359.900 239.330 360.220 ;
        RECT 240.400 359.800 240.590 360.410 ;
        RECT 240.730 360.060 241.000 360.410 ;
        RECT 240.730 360.010 241.010 360.060 ;
        RECT 240.840 359.920 241.010 360.010 ;
        RECT 240.400 359.770 240.620 359.800 ;
        RECT 240.380 359.500 240.630 359.770 ;
        RECT 240.390 359.490 240.630 359.500 ;
        RECT 240.390 359.250 240.620 359.490 ;
        RECT 237.280 358.870 237.470 358.920 ;
        RECT 237.540 358.880 238.590 359.170 ;
        RECT 234.810 357.730 235.130 358.050 ;
        RECT 235.670 357.970 235.900 358.050 ;
        RECT 235.330 357.450 235.590 357.770 ;
        RECT 235.670 357.760 236.000 357.970 ;
        RECT 235.690 357.680 236.000 357.760 ;
        RECT 236.080 357.770 236.530 358.090 ;
        RECT 236.670 358.020 236.990 358.340 ;
        RECT 237.280 358.310 237.470 358.360 ;
        RECT 231.140 357.240 231.340 357.280 ;
        RECT 233.350 357.120 233.580 357.150 ;
        RECT 231.690 356.970 231.880 357.000 ;
        RECT 232.130 356.970 232.410 357.000 ;
        RECT 231.680 356.950 231.880 356.970 ;
        RECT 232.120 356.950 232.410 356.970 ;
        RECT 231.680 356.930 231.870 356.950 ;
        RECT 231.680 356.890 232.050 356.930 ;
        RECT 229.120 355.900 229.380 356.690 ;
        RECT 231.730 356.610 232.050 356.890 ;
        RECT 232.120 356.920 232.400 356.950 ;
        RECT 232.120 356.620 232.440 356.920 ;
        RECT 233.350 356.860 233.700 357.120 ;
        RECT 233.360 356.800 233.700 356.860 ;
        RECT 233.770 357.070 234.090 357.360 ;
        RECT 234.290 357.150 234.610 357.450 ;
        RECT 234.650 357.240 234.840 357.300 ;
        RECT 235.690 357.190 235.880 357.680 ;
        RECT 235.690 357.170 235.970 357.190 ;
        RECT 235.710 357.150 235.970 357.170 ;
        RECT 234.290 357.120 234.720 357.150 ;
        RECT 235.320 357.140 235.970 357.150 ;
        RECT 236.080 357.140 236.360 357.770 ;
        RECT 236.720 357.370 237.040 357.690 ;
        RECT 237.540 357.410 238.480 358.880 ;
        RECT 240.000 358.440 240.240 358.820 ;
        RECT 240.430 358.230 240.590 359.250 ;
        RECT 240.840 358.230 241.000 359.920 ;
        RECT 341.570 358.150 345.330 361.770 ;
        RECT 355.920 361.080 359.330 361.400 ;
        RECT 238.930 357.650 239.250 357.970 ;
        RECT 355.920 357.850 362.560 361.080 ;
        RECT 237.540 357.400 238.280 357.410 ;
        RECT 235.320 357.120 236.360 357.140 ;
        RECT 234.290 357.090 236.360 357.120 ;
        RECT 232.810 356.500 233.020 356.710 ;
        RECT 233.360 356.640 233.580 356.800 ;
        RECT 233.770 356.750 233.970 357.070 ;
        RECT 234.440 357.040 236.360 357.090 ;
        RECT 234.470 357.010 236.360 357.040 ;
        RECT 234.500 356.990 236.360 357.010 ;
        RECT 234.570 356.980 235.530 356.990 ;
        RECT 235.710 356.870 236.360 356.990 ;
        RECT 236.490 357.110 236.760 357.160 ;
        RECT 236.490 356.970 237.030 357.110 ;
        RECT 237.570 357.090 238.280 357.400 ;
        RECT 235.810 356.830 236.360 356.870 ;
        RECT 234.410 356.500 234.730 356.770 ;
        RECT 232.810 356.180 233.140 356.500 ;
        RECT 234.410 356.450 234.900 356.500 ;
        RECT 229.120 354.790 229.350 355.900 ;
        RECT 232.460 355.330 232.780 355.650 ;
        RECT 232.810 354.940 233.020 356.180 ;
        RECT 233.810 355.920 234.130 356.240 ;
        RECT 234.330 355.970 234.560 356.170 ;
        RECT 234.230 355.880 234.560 355.970 ;
        RECT 234.230 355.470 234.420 355.880 ;
        RECT 234.050 355.220 234.420 355.470 ;
        RECT 234.710 355.550 234.900 356.450 ;
        RECT 234.710 355.260 235.020 355.550 ;
        RECT 234.050 355.150 234.410 355.220 ;
        RECT 234.150 355.050 234.410 355.150 ;
        RECT 234.710 354.980 234.900 355.260 ;
        RECT 232.890 354.620 233.120 354.910 ;
        RECT 235.640 354.790 235.830 354.840 ;
        RECT 236.080 354.790 236.360 356.830 ;
        RECT 236.470 356.820 237.030 356.970 ;
        RECT 236.710 356.790 237.030 356.820 ;
        RECT 237.530 357.080 238.280 357.090 ;
        RECT 237.280 356.750 237.470 356.790 ;
        RECT 236.660 356.140 236.980 356.460 ;
        RECT 237.530 355.730 238.470 357.080 ;
        RECT 238.960 356.810 239.280 357.130 ;
        RECT 240.000 356.810 240.240 357.190 ;
        RECT 240.430 356.380 240.590 357.400 ;
        RECT 240.390 356.140 240.620 356.380 ;
        RECT 240.390 356.130 240.630 356.140 ;
        RECT 240.380 355.860 240.630 356.130 ;
        RECT 240.400 355.830 240.620 355.860 ;
        RECT 237.530 355.440 238.580 355.730 ;
        RECT 236.660 354.990 236.980 355.310 ;
        RECT 236.710 354.340 237.030 354.660 ;
        RECT 236.710 353.790 237.030 354.110 ;
        RECT 236.660 353.140 236.980 353.460 ;
        RECT 237.530 353.190 238.470 355.440 ;
        RECT 238.880 354.910 239.190 355.190 ;
        RECT 238.880 354.750 239.330 354.910 ;
        RECT 239.010 354.590 239.330 354.750 ;
        RECT 240.400 354.380 240.590 355.830 ;
        RECT 240.840 355.710 241.000 357.400 ;
        RECT 240.840 355.620 241.010 355.710 ;
        RECT 240.730 355.570 241.010 355.620 ;
        RECT 240.730 355.020 241.000 355.570 ;
        RECT 240.840 354.380 241.000 355.020 ;
        RECT 239.000 353.870 239.320 354.190 ;
        RECT 237.440 353.140 238.470 353.190 ;
        RECT 237.440 352.850 238.580 353.140 ;
        RECT 232.400 352.240 232.720 352.560 ;
        RECT 237.440 352.400 238.470 352.850 ;
        RECT 236.660 351.990 236.980 352.310 ;
        RECT 237.530 352.040 237.870 352.400 ;
        RECT 237.530 351.750 237.920 352.040 ;
        RECT 232.550 351.410 232.870 351.730 ;
        RECT 234.300 351.120 234.630 351.410 ;
        RECT 236.710 351.340 237.030 351.660 ;
        RECT 237.530 351.370 237.870 351.750 ;
        RECT 238.200 351.380 238.470 352.400 ;
        RECT 238.920 351.620 239.240 351.940 ;
        RECT 234.290 351.090 234.710 351.120 ;
        RECT 235.310 351.110 235.810 351.120 ;
        RECT 235.310 351.090 236.150 351.110 ;
        RECT 234.290 350.980 236.150 351.090 ;
        RECT 231.680 350.920 231.870 350.970 ;
        RECT 232.120 350.920 232.400 350.970 ;
        RECT 234.570 350.950 235.470 350.980 ;
        RECT 235.810 350.920 236.150 350.980 ;
        RECT 236.480 350.920 236.750 351.130 ;
        RECT 231.720 350.580 232.040 350.900 ;
        RECT 232.800 350.470 233.010 350.680 ;
        RECT 232.800 350.150 233.130 350.470 ;
        RECT 232.450 349.300 232.770 349.620 ;
        RECT 232.800 348.910 233.010 350.150 ;
        RECT 232.880 348.590 233.110 348.880 ;
        RECT 233.160 334.360 233.880 334.930 ;
        RECT 226.970 333.210 227.210 333.440 ;
        RECT 226.970 325.660 227.200 333.210 ;
        RECT 233.220 327.350 233.730 334.360 ;
        RECT 264.240 327.690 268.660 357.800 ;
        RECT 355.920 357.360 359.330 357.850 ;
        RECT 347.510 332.490 349.830 332.570 ;
        RECT 347.510 329.260 362.550 332.490 ;
        RECT 347.510 329.200 349.830 329.260 ;
        RECT 233.080 327.300 233.730 327.350 ;
        RECT 233.070 327.120 233.730 327.300 ;
        RECT 233.040 327.110 233.730 327.120 ;
        RECT 233.040 326.740 233.640 327.110 ;
        RECT 226.970 325.430 227.330 325.660 ;
        RECT 226.970 324.050 227.200 325.430 ;
        RECT 232.620 324.870 232.940 325.010 ;
        RECT 233.040 324.870 233.620 326.740 ;
        RECT 264.210 326.370 268.680 327.690 ;
        RECT 232.620 324.690 233.620 324.870 ;
        RECT 232.690 324.340 233.620 324.690 ;
        RECT 226.970 323.820 227.330 324.050 ;
        RECT 232.620 324.020 233.620 324.340 ;
        RECT 232.690 323.880 233.620 324.020 ;
        RECT 226.970 322.450 227.200 323.820 ;
        RECT 233.040 323.100 233.620 323.880 ;
        RECT 232.630 322.910 232.950 322.960 ;
        RECT 232.400 322.680 232.950 322.910 ;
        RECT 232.630 322.640 232.950 322.680 ;
        RECT 233.090 322.500 233.620 323.100 ;
        RECT 233.050 322.490 233.620 322.500 ;
        RECT 226.970 322.220 227.330 322.450 ;
        RECT 226.970 320.830 227.200 322.220 ;
        RECT 233.040 321.490 233.620 322.490 ;
        RECT 232.630 321.300 232.950 321.350 ;
        RECT 228.450 321.240 228.960 321.300 ;
        RECT 228.450 321.070 230.690 321.240 ;
        RECT 232.400 321.070 232.950 321.300 ;
        RECT 228.680 321.040 230.690 321.070 ;
        RECT 226.970 320.600 227.330 320.830 ;
        RECT 226.970 319.230 227.200 320.600 ;
        RECT 227.790 319.520 228.110 319.690 ;
        RECT 227.790 319.430 229.530 319.520 ;
        RECT 227.990 319.340 229.530 319.430 ;
        RECT 226.970 319.000 227.330 319.230 ;
        RECT 226.970 317.610 227.200 319.000 ;
        RECT 230.520 317.790 230.690 321.040 ;
        RECT 232.630 321.030 232.950 321.070 ;
        RECT 233.090 320.890 233.620 321.490 ;
        RECT 233.040 319.880 233.620 320.890 ;
        RECT 232.620 319.690 232.940 319.740 ;
        RECT 232.390 319.460 232.940 319.690 ;
        RECT 230.750 319.220 231.260 319.440 ;
        RECT 232.620 319.420 232.940 319.460 ;
        RECT 233.080 319.280 233.620 319.880 ;
        RECT 230.970 319.210 231.260 319.220 ;
        RECT 233.040 318.260 233.620 319.280 ;
        RECT 232.630 318.070 232.950 318.120 ;
        RECT 232.400 317.860 232.950 318.070 ;
        RECT 232.100 317.840 232.950 317.860 ;
        RECT 232.100 317.640 232.610 317.840 ;
        RECT 232.630 317.800 232.950 317.840 ;
        RECT 233.090 317.660 233.620 318.260 ;
        RECT 232.100 317.630 232.390 317.640 ;
        RECT 226.970 317.380 227.330 317.610 ;
        RECT 226.970 316.010 227.200 317.380 ;
        RECT 233.040 316.650 233.620 317.660 ;
        RECT 232.620 316.460 232.940 316.510 ;
        RECT 232.390 316.230 232.940 316.460 ;
        RECT 232.620 316.190 232.940 316.230 ;
        RECT 233.080 316.050 233.620 316.650 ;
        RECT 226.970 315.780 227.330 316.010 ;
        RECT 225.600 314.000 226.040 314.460 ;
        RECT 226.970 314.390 227.200 315.780 ;
        RECT 232.210 314.540 232.530 314.860 ;
        RECT 226.970 314.160 227.330 314.390 ;
        RECT 232.260 314.310 232.490 314.540 ;
        RECT 233.040 314.180 233.620 316.050 ;
        RECT 226.970 314.090 227.200 314.160 ;
        RECT 232.620 313.260 232.940 313.310 ;
        RECT 232.390 313.030 232.940 313.260 ;
        RECT 232.620 312.990 232.940 313.030 ;
        RECT 233.080 311.970 233.620 314.180 ;
        RECT 229.380 311.550 229.700 311.600 ;
        RECT 230.320 311.550 230.640 311.600 ;
        RECT 229.150 311.320 229.700 311.550 ;
        RECT 230.090 311.320 230.640 311.550 ;
        RECT 231.270 311.530 231.590 311.580 ;
        RECT 232.580 311.550 232.900 311.600 ;
        RECT 229.380 311.280 229.700 311.320 ;
        RECT 230.320 311.280 230.640 311.320 ;
        RECT 231.040 311.300 231.590 311.530 ;
        RECT 232.350 311.320 232.900 311.550 ;
        RECT 231.270 311.260 231.590 311.300 ;
        RECT 232.580 311.280 232.900 311.320 ;
        RECT 186.560 310.420 187.480 311.150 ;
        RECT 186.530 309.690 187.450 310.420 ;
        RECT 12.160 304.620 12.930 304.640 ;
        RECT 27.610 304.620 29.840 304.700 ;
        RECT 3.630 302.870 29.840 304.620 ;
        RECT 2.680 302.860 29.840 302.870 ;
        RECT 2.520 302.510 29.840 302.860 ;
        RECT 2.680 302.500 29.840 302.510 ;
        RECT 3.630 302.150 29.840 302.500 ;
        RECT 4.000 301.390 29.840 302.150 ;
        RECT 4.000 300.710 13.570 301.390 ;
        RECT 27.610 301.240 29.840 301.390 ;
        RECT 5.460 291.000 10.610 300.710 ;
        RECT 12.160 300.690 13.570 300.710 ;
        RECT 12.930 300.680 13.570 300.690 ;
        RECT 4.170 290.910 4.800 290.970 ;
        RECT 4.170 290.330 4.820 290.910 ;
        RECT 5.470 290.330 10.610 291.000 ;
        RECT 4.170 289.580 4.800 290.330 ;
        RECT 4.170 288.860 12.430 289.580 ;
        RECT 4.170 288.630 6.760 288.860 ;
        RECT 4.170 288.600 4.800 288.630 ;
        RECT 4.650 287.480 5.640 287.490 ;
        RECT 4.250 286.960 5.640 287.480 ;
        RECT 4.250 283.350 4.740 286.960 ;
        RECT 7.450 286.430 10.870 286.480 ;
        RECT 7.440 285.860 10.880 286.430 ;
        RECT 6.030 276.030 10.330 285.090 ;
        RECT 12.010 285.040 12.730 285.590 ;
        RECT 12.010 285.030 12.510 285.040 ;
        RECT 12.160 276.040 12.930 276.050 ;
        RECT 12.160 276.030 13.560 276.040 ;
        RECT 32.120 276.030 34.530 276.130 ;
        RECT 3.630 274.280 34.530 276.030 ;
        RECT 2.680 274.270 34.530 274.280 ;
        RECT 2.520 273.920 34.530 274.270 ;
        RECT 2.680 273.910 34.530 273.920 ;
        RECT 3.630 273.560 34.530 273.910 ;
        RECT 4.000 272.800 34.530 273.560 ;
        RECT 4.000 272.120 13.560 272.800 ;
        RECT 32.120 272.700 34.530 272.800 ;
        RECT 5.460 262.410 10.610 272.120 ;
        RECT 12.160 272.100 13.560 272.120 ;
        RECT 4.170 262.320 4.800 262.380 ;
        RECT 4.170 261.740 4.820 262.320 ;
        RECT 5.470 261.740 10.610 262.410 ;
        RECT 4.170 260.990 4.800 261.740 ;
        RECT 4.170 260.270 12.430 260.990 ;
        RECT 4.170 260.040 6.760 260.270 ;
        RECT 4.170 260.010 4.800 260.040 ;
        RECT 4.650 258.890 5.640 258.900 ;
        RECT 4.250 258.370 5.640 258.890 ;
        RECT 4.250 254.760 4.740 258.370 ;
        RECT 7.450 257.840 10.870 257.890 ;
        RECT 7.440 257.270 10.880 257.840 ;
        RECT 6.030 247.440 10.330 256.500 ;
        RECT 12.010 256.450 12.730 257.000 ;
        RECT 12.010 256.440 12.510 256.450 ;
        RECT 12.160 247.440 13.570 247.460 ;
        RECT 36.680 247.440 38.950 247.510 ;
        RECT 3.630 245.690 38.950 247.440 ;
        RECT 2.680 245.680 38.950 245.690 ;
        RECT 2.520 245.330 38.950 245.680 ;
        RECT 2.680 245.320 38.950 245.330 ;
        RECT 3.630 244.970 38.950 245.320 ;
        RECT 4.000 244.210 38.950 244.970 ;
        RECT 4.000 243.530 13.570 244.210 ;
        RECT 36.680 244.110 38.950 244.210 ;
        RECT 5.460 233.820 10.610 243.530 ;
        RECT 12.160 243.520 13.570 243.530 ;
        RECT 12.160 243.510 12.930 243.520 ;
        RECT 4.170 233.730 4.800 233.790 ;
        RECT 4.170 233.150 4.820 233.730 ;
        RECT 5.470 233.150 10.610 233.820 ;
        RECT 4.170 232.400 4.800 233.150 ;
        RECT 4.170 231.680 12.430 232.400 ;
        RECT 4.170 231.450 6.760 231.680 ;
        RECT 4.170 231.420 4.800 231.450 ;
        RECT 4.650 230.300 5.640 230.310 ;
        RECT 4.250 229.780 5.640 230.300 ;
        RECT 4.250 226.170 4.740 229.780 ;
        RECT 7.450 229.250 10.870 229.300 ;
        RECT 7.440 228.680 10.880 229.250 ;
        RECT 6.030 218.850 10.330 227.910 ;
        RECT 12.010 227.860 12.730 228.410 ;
        RECT 12.010 227.850 12.510 227.860 ;
        RECT 12.160 218.850 13.560 218.870 ;
        RECT 41.040 218.850 43.290 218.910 ;
        RECT 3.630 217.100 43.290 218.850 ;
        RECT 2.680 217.090 43.290 217.100 ;
        RECT 2.520 216.740 43.290 217.090 ;
        RECT 2.680 216.730 43.290 216.740 ;
        RECT 3.630 216.380 43.290 216.730 ;
        RECT 4.000 215.620 43.290 216.380 ;
        RECT 4.000 214.940 13.560 215.620 ;
        RECT 41.040 215.540 43.290 215.620 ;
        RECT 5.460 205.230 10.610 214.940 ;
        RECT 12.160 214.930 13.560 214.940 ;
        RECT 12.160 214.920 12.930 214.930 ;
        RECT 4.170 205.140 4.800 205.200 ;
        RECT 4.170 204.560 4.820 205.140 ;
        RECT 5.470 204.560 10.610 205.230 ;
        RECT 4.170 203.810 4.800 204.560 ;
        RECT 4.170 203.090 12.430 203.810 ;
        RECT 4.170 202.860 6.760 203.090 ;
        RECT 4.170 202.830 4.800 202.860 ;
        RECT 4.650 201.710 5.640 201.720 ;
        RECT 4.250 201.190 5.640 201.710 ;
        RECT 4.250 197.580 4.740 201.190 ;
        RECT 7.450 200.660 10.870 200.710 ;
        RECT 7.440 200.090 10.880 200.660 ;
        RECT 6.030 190.260 10.330 199.320 ;
        RECT 12.010 199.270 12.730 199.820 ;
        RECT 12.010 199.260 12.510 199.270 ;
        RECT 12.160 190.260 13.560 190.280 ;
        RECT 45.360 190.260 47.610 190.370 ;
        RECT 3.630 188.510 47.760 190.260 ;
        RECT 2.680 188.500 47.760 188.510 ;
        RECT 2.520 188.150 47.760 188.500 ;
        RECT 2.680 188.140 47.760 188.150 ;
        RECT 3.630 187.790 47.760 188.140 ;
        RECT 4.000 187.030 47.760 187.790 ;
        RECT 4.000 186.350 13.560 187.030 ;
        RECT 45.360 186.920 47.610 187.030 ;
        RECT 5.460 176.640 10.610 186.350 ;
        RECT 12.160 186.340 13.560 186.350 ;
        RECT 12.160 186.330 12.930 186.340 ;
        RECT 4.170 176.550 4.800 176.610 ;
        RECT 4.170 175.970 4.820 176.550 ;
        RECT 5.470 175.970 10.610 176.640 ;
        RECT 4.170 175.220 4.800 175.970 ;
        RECT 4.170 174.500 12.430 175.220 ;
        RECT 4.170 174.270 6.760 174.500 ;
        RECT 4.170 174.240 4.800 174.270 ;
        RECT 4.650 173.120 5.640 173.130 ;
        RECT 4.250 172.600 5.640 173.120 ;
        RECT 4.250 168.990 4.740 172.600 ;
        RECT 7.450 172.070 10.870 172.120 ;
        RECT 7.440 171.500 10.880 172.070 ;
        RECT 6.030 161.670 10.330 170.730 ;
        RECT 12.010 170.680 12.730 171.230 ;
        RECT 12.010 170.670 12.510 170.680 ;
        RECT 264.240 165.070 268.660 326.370 ;
        RECT 343.340 303.900 345.700 304.030 ;
        RECT 343.340 300.670 362.570 303.900 ;
        RECT 343.340 300.570 345.700 300.670 ;
        RECT 339.330 275.310 341.610 275.470 ;
        RECT 339.330 272.080 362.550 275.310 ;
        RECT 339.330 271.970 341.610 272.080 ;
        RECT 335.030 246.720 337.450 246.840 ;
        RECT 335.030 243.490 362.550 246.720 ;
        RECT 335.030 243.330 337.450 243.490 ;
        RECT 331.140 218.130 333.410 218.240 ;
        RECT 331.140 214.900 362.560 218.130 ;
        RECT 331.140 214.770 333.410 214.900 ;
        RECT 326.740 189.540 329.040 189.620 ;
        RECT 326.740 186.310 362.560 189.540 ;
        RECT 326.740 186.210 329.040 186.310 ;
        RECT 12.160 161.680 12.930 161.690 ;
        RECT 12.160 161.670 13.560 161.680 ;
        RECT 49.420 161.670 51.830 161.770 ;
        RECT 3.630 159.920 51.830 161.670 ;
        RECT 263.320 161.330 268.660 165.070 ;
        RECT 263.320 160.370 268.080 161.330 ;
        RECT 2.680 159.910 51.830 159.920 ;
        RECT 2.520 159.560 51.830 159.910 ;
        RECT 2.680 159.550 51.830 159.560 ;
        RECT 3.630 159.200 51.830 159.550 ;
        RECT 4.000 158.440 51.830 159.200 ;
        RECT 4.000 157.760 13.560 158.440 ;
        RECT 49.420 158.260 51.830 158.440 ;
        RECT 5.460 148.050 10.610 157.760 ;
        RECT 12.160 157.740 13.560 157.760 ;
        RECT 4.170 147.960 4.800 148.020 ;
        RECT 4.170 147.380 4.820 147.960 ;
        RECT 5.470 147.380 10.610 148.050 ;
        RECT 4.170 146.630 4.800 147.380 ;
        RECT 4.170 145.910 12.430 146.630 ;
        RECT 4.170 145.680 6.760 145.910 ;
        RECT 4.170 145.650 4.800 145.680 ;
        RECT 4.650 144.530 5.640 144.540 ;
        RECT 4.250 144.010 5.640 144.530 ;
        RECT 4.250 140.400 4.740 144.010 ;
        RECT 7.450 143.480 10.870 143.530 ;
        RECT 7.440 142.910 10.880 143.480 ;
        RECT 6.030 133.080 10.330 142.140 ;
        RECT 12.010 142.090 12.730 142.640 ;
        RECT 12.010 142.080 12.510 142.090 ;
        RECT 12.160 133.090 12.930 133.100 ;
        RECT 12.160 133.080 13.560 133.090 ;
        RECT 53.700 133.080 56.160 133.150 ;
        RECT 3.630 131.330 56.160 133.080 ;
        RECT 2.680 131.320 56.160 131.330 ;
        RECT 2.520 130.970 56.160 131.320 ;
        RECT 2.680 130.960 56.160 130.970 ;
        RECT 3.630 130.610 56.160 130.960 ;
        RECT 4.000 129.850 56.160 130.610 ;
        RECT 4.000 129.170 13.560 129.850 ;
        RECT 53.700 129.800 56.160 129.850 ;
        RECT 5.460 119.460 10.610 129.170 ;
        RECT 12.160 129.150 13.560 129.170 ;
        RECT 4.170 119.370 4.800 119.430 ;
        RECT 4.170 118.790 4.820 119.370 ;
        RECT 5.470 118.790 10.610 119.460 ;
        RECT 4.170 118.040 4.800 118.790 ;
        RECT 4.170 117.320 12.430 118.040 ;
        RECT 4.170 117.090 6.760 117.320 ;
        RECT 4.170 117.060 4.800 117.090 ;
        RECT 4.650 115.940 5.640 115.950 ;
        RECT 4.250 115.420 5.640 115.940 ;
        RECT 4.250 111.810 4.740 115.420 ;
        RECT 7.450 114.890 10.870 114.940 ;
        RECT 7.440 114.320 10.880 114.890 ;
        RECT 6.030 104.490 10.330 113.550 ;
        RECT 12.010 113.500 12.730 114.050 ;
        RECT 12.010 113.490 12.510 113.500 ;
        RECT 12.910 104.510 13.550 104.520 ;
        RECT 12.160 104.490 13.550 104.510 ;
        RECT 58.070 104.490 60.470 104.630 ;
        RECT 3.630 102.740 60.470 104.490 ;
        RECT 2.680 102.730 60.470 102.740 ;
        RECT 2.520 102.380 60.470 102.730 ;
        RECT 2.680 102.370 60.470 102.380 ;
        RECT 3.630 102.020 60.470 102.370 ;
        RECT 4.000 101.260 60.470 102.020 ;
        RECT 4.000 100.580 13.550 101.260 ;
        RECT 58.070 101.160 60.470 101.260 ;
        RECT 5.460 90.870 10.610 100.580 ;
        RECT 12.160 100.560 12.930 100.580 ;
        RECT 4.170 90.780 4.800 90.840 ;
        RECT 4.170 90.200 4.820 90.780 ;
        RECT 5.470 90.200 10.610 90.870 ;
        RECT 4.170 89.450 4.800 90.200 ;
        RECT 4.170 88.730 12.430 89.450 ;
        RECT 4.170 88.500 6.760 88.730 ;
        RECT 4.170 88.470 4.800 88.500 ;
        RECT 4.650 87.350 5.640 87.360 ;
        RECT 4.250 86.830 5.640 87.350 ;
        RECT 4.250 83.220 4.740 86.830 ;
        RECT 7.450 86.300 10.870 86.350 ;
        RECT 7.440 85.730 10.880 86.300 ;
        RECT 6.030 75.900 10.330 84.960 ;
        RECT 12.010 84.910 12.730 85.460 ;
        RECT 12.010 84.900 12.510 84.910 ;
        RECT 12.160 75.900 13.550 75.920 ;
        RECT 62.010 75.900 64.500 75.980 ;
        RECT 3.630 74.150 64.500 75.900 ;
        RECT 2.680 74.140 64.500 74.150 ;
        RECT 2.520 73.790 64.500 74.140 ;
        RECT 2.680 73.780 64.500 73.790 ;
        RECT 3.630 73.430 64.500 73.780 ;
        RECT 4.000 72.670 64.500 73.430 ;
        RECT 4.000 71.990 13.550 72.670 ;
        RECT 62.010 72.480 64.500 72.670 ;
        RECT 5.460 62.280 10.610 71.990 ;
        RECT 12.160 71.980 13.550 71.990 ;
        RECT 12.160 71.970 12.930 71.980 ;
        RECT 4.170 62.190 4.800 62.250 ;
        RECT 4.170 61.610 4.820 62.190 ;
        RECT 5.470 61.610 10.610 62.280 ;
        RECT 4.170 60.860 4.800 61.610 ;
        RECT 4.170 60.140 12.430 60.860 ;
        RECT 4.170 59.910 6.760 60.140 ;
        RECT 4.170 59.880 4.800 59.910 ;
        RECT 4.650 58.760 5.640 58.770 ;
        RECT 4.250 58.240 5.640 58.760 ;
        RECT 4.250 54.630 4.740 58.240 ;
        RECT 7.450 57.710 10.870 57.760 ;
        RECT 7.440 57.140 10.880 57.710 ;
        RECT 6.030 47.310 10.330 56.370 ;
        RECT 12.010 56.320 12.730 56.870 ;
        RECT 12.010 56.310 12.510 56.320 ;
        RECT 12.160 47.320 12.930 47.330 ;
        RECT 12.160 47.310 13.570 47.320 ;
        RECT 66.480 47.310 68.830 47.410 ;
        RECT 3.630 45.560 68.830 47.310 ;
        RECT 2.680 45.550 68.830 45.560 ;
        RECT 2.520 45.200 68.830 45.550 ;
        RECT 2.680 45.190 68.830 45.200 ;
        RECT 3.630 44.840 68.830 45.190 ;
        RECT 4.000 44.080 68.830 44.840 ;
        RECT 4.000 43.400 13.570 44.080 ;
        RECT 66.480 43.950 68.830 44.080 ;
        RECT 5.460 33.690 10.610 43.400 ;
        RECT 12.160 43.380 13.570 43.400 ;
        RECT 4.170 33.600 4.800 33.660 ;
        RECT 4.170 33.020 4.820 33.600 ;
        RECT 5.470 33.020 10.610 33.690 ;
        RECT 4.170 32.270 4.800 33.020 ;
        RECT 4.170 31.550 12.430 32.270 ;
        RECT 4.170 31.320 6.760 31.550 ;
        RECT 4.170 31.290 4.800 31.320 ;
        RECT 4.650 30.170 5.640 30.180 ;
        RECT 4.250 29.650 5.640 30.170 ;
        RECT 4.250 26.040 4.740 29.650 ;
        RECT 7.450 29.120 10.870 29.170 ;
        RECT 7.440 28.550 10.880 29.120 ;
        RECT 6.030 18.720 10.330 27.780 ;
        RECT 12.010 27.730 12.730 28.280 ;
        RECT 12.010 27.720 12.510 27.730 ;
        RECT 12.930 18.740 13.570 18.750 ;
        RECT 12.160 18.720 13.570 18.740 ;
        RECT 70.480 18.720 73.190 18.780 ;
        RECT 3.630 16.970 73.190 18.720 ;
        RECT 2.680 16.960 73.190 16.970 ;
        RECT 2.520 16.610 73.190 16.960 ;
        RECT 2.680 16.600 73.190 16.610 ;
        RECT 3.630 16.250 73.190 16.600 ;
        RECT 4.000 15.490 73.190 16.250 ;
        RECT 4.000 14.810 13.570 15.490 ;
        RECT 70.480 15.370 73.190 15.490 ;
        RECT 5.460 5.100 10.610 14.810 ;
        RECT 12.160 14.790 12.930 14.810 ;
        RECT 4.170 5.010 4.800 5.070 ;
        RECT 4.170 4.430 4.820 5.010 ;
        RECT 5.470 4.430 10.610 5.100 ;
        RECT 4.170 3.680 4.800 4.430 ;
        RECT 4.170 2.960 12.430 3.680 ;
        RECT 4.170 2.730 6.760 2.960 ;
        RECT 4.170 2.700 4.800 2.730 ;
      LAYER via ;
        RECT 16.590 385.280 18.620 385.610 ;
        RECT 16.530 384.420 17.230 385.040 ;
        RECT 39.980 385.280 42.970 385.630 ;
        RECT 45.180 385.280 47.210 385.610 ;
        RECT 43.410 384.480 43.760 385.240 ;
        RECT 45.120 384.420 45.820 385.040 ;
        RECT 68.570 385.280 71.560 385.630 ;
        RECT 73.770 385.280 75.800 385.610 ;
        RECT 42.380 379.190 42.800 382.360 ;
        RECT 41.410 377.370 41.930 377.890 ;
        RECT 72.000 384.480 72.350 385.240 ;
        RECT 73.710 384.420 74.410 385.040 ;
        RECT 129.970 385.980 153.770 386.240 ;
        RECT 97.160 385.280 100.150 385.630 ;
        RECT 70.970 379.190 71.390 382.360 ;
        RECT 70.000 377.370 70.520 377.890 ;
        RECT 100.590 384.480 100.940 385.240 ;
        RECT 99.560 379.190 99.980 382.360 ;
        RECT 126.810 379.690 127.200 380.080 ;
        RECT 98.590 377.370 99.110 377.890 ;
        RECT 4.690 372.820 5.450 373.170 ;
        RECT 4.300 369.390 4.650 372.380 ;
        RECT 7.570 371.790 10.740 372.210 ;
        RECT 12.040 370.820 12.560 371.340 ;
        RECT 86.320 370.730 89.550 372.980 ;
        RECT 98.510 369.450 99.030 369.820 ;
        RECT 57.730 366.240 60.960 368.490 ;
        RECT 27.310 361.970 29.560 365.200 ;
        RECT 15.780 358.570 17.640 361.800 ;
        RECT 162.650 385.980 183.510 386.240 ;
        RECT 157.790 385.280 159.820 385.610 ;
        RECT 157.730 384.420 158.430 385.040 ;
        RECT 181.180 385.280 184.170 385.630 ;
        RECT 186.380 385.280 188.410 385.610 ;
        RECT 184.610 384.480 184.960 385.240 ;
        RECT 186.320 384.420 187.020 385.040 ;
        RECT 209.770 385.280 212.760 385.630 ;
        RECT 214.970 385.280 217.000 385.610 ;
        RECT 120.020 376.280 120.280 376.540 ;
        RECT 122.880 376.330 123.140 376.590 ;
        RECT 126.890 376.240 127.280 376.630 ;
        RECT 120.010 375.250 120.270 375.510 ;
        RECT 120.680 375.270 120.940 375.530 ;
        RECT 121.420 375.260 121.680 375.520 ;
        RECT 120.010 374.800 120.270 375.060 ;
        RECT 121.420 374.820 121.680 375.080 ;
        RECT 120.010 374.380 120.270 374.640 ;
        RECT 120.680 374.430 120.940 374.690 ;
        RECT 121.440 374.400 121.700 374.660 ;
        RECT 120.010 373.030 120.270 373.290 ;
        RECT 122.660 374.690 122.920 374.950 ;
        RECT 122.380 372.530 122.640 372.790 ;
        RECT 120.660 371.630 120.920 371.890 ;
        RECT 122.090 371.650 122.350 371.910 ;
        RECT 119.870 371.050 120.130 371.310 ;
        RECT 120.800 371.050 121.060 371.310 ;
        RECT 121.500 371.050 121.760 371.310 ;
        RECT 122.240 371.050 122.500 371.310 ;
        RECT 122.950 371.040 123.210 371.300 ;
        RECT 101.850 365.070 102.260 365.480 ;
        RECT 98.370 361.130 98.890 361.650 ;
        RECT 4.320 346.000 4.650 348.030 ;
        RECT 4.890 345.940 5.510 346.640 ;
        RECT 4.690 344.230 5.450 344.580 ;
        RECT 4.300 340.800 4.650 343.790 ;
        RECT 7.570 343.200 10.740 343.620 ;
        RECT 12.040 342.230 12.560 342.750 ;
        RECT 23.830 329.980 25.910 333.210 ;
        RECT 101.900 360.280 102.310 360.690 ;
        RECT 98.470 325.110 98.990 325.630 ;
        RECT 101.900 324.170 102.310 324.610 ;
        RECT 4.320 317.410 4.650 319.440 ;
        RECT 128.270 375.070 128.530 375.330 ;
        RECT 136.070 374.530 136.330 374.790 ;
        RECT 137.430 374.610 137.690 374.870 ;
        RECT 138.120 374.600 138.380 374.860 ;
        RECT 169.800 377.120 170.220 377.540 ;
        RECT 165.950 376.360 166.370 376.780 ;
        RECT 171.470 374.750 171.910 375.190 ;
        RECT 167.050 373.730 167.490 374.170 ;
        RECT 177.190 374.750 177.630 375.190 ;
        RECT 183.580 379.190 184.000 382.360 ;
        RECT 182.610 377.370 183.130 377.890 ;
        RECT 179.010 374.720 179.450 375.160 ;
        RECT 172.760 373.730 173.200 374.170 ;
        RECT 128.190 372.370 128.610 372.790 ;
        RECT 134.140 370.970 134.430 371.550 ;
        RECT 135.350 370.870 135.610 371.130 ;
        RECT 145.210 370.890 145.470 371.150 ;
        RECT 147.430 369.910 147.690 370.170 ;
        RECT 143.760 364.730 144.020 364.990 ;
        RECT 141.350 363.660 141.610 363.920 ;
        RECT 142.220 363.820 142.480 364.080 ;
        RECT 143.770 363.740 144.030 364.000 ;
        RECT 141.320 362.740 141.580 363.000 ;
        RECT 142.200 362.900 142.460 363.160 ;
        RECT 143.770 362.750 144.030 363.010 ;
        RECT 141.330 361.820 141.590 362.080 ;
        RECT 142.180 361.910 142.440 362.170 ;
        RECT 143.680 361.960 143.940 362.220 ;
        RECT 140.680 360.800 140.940 361.060 ;
        RECT 140.640 359.840 140.900 360.100 ;
        RECT 140.680 358.880 140.940 359.140 ;
        RECT 143.510 361.350 143.770 361.610 ;
        RECT 143.680 360.970 143.940 361.230 ;
        RECT 143.510 360.360 143.770 360.620 ;
        RECT 143.680 359.980 143.940 360.240 ;
        RECT 153.220 369.480 153.530 369.790 ;
        RECT 164.290 370.710 164.550 370.970 ;
        RECT 157.220 370.020 157.480 370.280 ;
        RECT 156.050 369.030 156.320 369.290 ;
        RECT 144.720 368.250 145.070 368.600 ;
        RECT 149.970 368.560 150.230 368.820 ;
        RECT 166.420 367.190 166.680 367.450 ;
        RECT 168.520 368.030 168.780 368.290 ;
        RECT 169.460 367.550 169.720 367.810 ;
        RECT 170.500 367.590 170.760 367.850 ;
        RECT 170.560 367.310 170.820 367.570 ;
        RECT 145.740 366.010 146.000 366.400 ;
        RECT 162.140 366.020 162.470 366.280 ;
        RECT 145.100 365.190 145.360 365.590 ;
        RECT 144.850 364.740 145.110 365.000 ;
        RECT 145.120 364.080 145.380 364.340 ;
        RECT 144.860 363.750 145.120 364.010 ;
        RECT 143.510 359.370 143.770 359.630 ;
        RECT 140.640 343.600 140.900 344.070 ;
        RECT 141.280 343.600 141.540 344.070 ;
        RECT 139.280 342.570 139.540 342.830 ;
        RECT 138.760 342.170 139.020 342.430 ;
        RECT 129.480 340.920 130.140 341.580 ;
        RECT 141.360 342.550 141.620 342.810 ;
        RECT 143.120 342.560 143.390 342.830 ;
        RECT 140.700 342.190 140.960 342.450 ;
        RECT 138.780 338.260 139.040 338.520 ;
        RECT 134.690 336.400 135.060 336.770 ;
        RECT 129.520 335.060 130.180 335.720 ;
        RECT 138.640 335.020 138.900 335.280 ;
        RECT 143.620 342.170 143.880 342.430 ;
        RECT 145.120 363.160 145.380 363.420 ;
        RECT 144.860 362.760 145.120 363.020 ;
        RECT 145.090 362.240 145.350 362.500 ;
        RECT 144.980 361.860 145.240 362.120 ;
        RECT 144.980 360.870 145.240 361.130 ;
        RECT 144.980 359.880 145.240 360.140 ;
        RECT 161.510 364.300 161.840 364.630 ;
        RECT 160.940 362.820 161.270 363.150 ;
        RECT 145.730 361.150 145.990 361.410 ;
        RECT 160.300 361.220 160.630 361.550 ;
        RECT 159.660 360.650 159.990 360.980 ;
        RECT 145.740 360.190 146.000 360.450 ;
        RECT 145.730 359.230 145.990 359.490 ;
        RECT 145.090 341.570 145.350 341.830 ;
        RECT 144.470 340.420 144.730 340.680 ;
        RECT 144.170 339.570 144.430 339.830 ;
        RECT 143.670 338.270 143.930 338.530 ;
        RECT 144.050 337.810 144.310 338.070 ;
        RECT 143.670 336.720 143.930 336.980 ;
        RECT 141.950 335.460 142.210 335.720 ;
        RECT 139.740 335.030 140.000 335.290 ;
        RECT 140.830 335.030 141.090 335.290 ;
        RECT 141.960 334.990 142.220 335.250 ;
        RECT 139.190 334.350 139.450 334.610 ;
        RECT 140.290 334.350 140.550 334.610 ;
        RECT 141.390 334.350 141.650 334.610 ;
        RECT 139.190 332.980 139.450 333.240 ;
        RECT 140.290 332.980 140.550 333.240 ;
        RECT 141.390 332.980 141.650 333.240 ;
        RECT 138.640 332.250 138.900 332.510 ;
        RECT 139.740 332.250 140.000 332.510 ;
        RECT 140.830 332.250 141.090 332.510 ;
        RECT 138.630 330.910 138.890 331.170 ;
        RECT 139.740 330.900 140.000 331.160 ;
        RECT 140.830 330.880 141.090 331.140 ;
        RECT 134.680 330.160 135.050 330.530 ;
        RECT 139.190 330.210 139.450 330.470 ;
        RECT 140.290 330.200 140.550 330.460 ;
        RECT 141.380 330.200 141.640 330.460 ;
        RECT 142.220 329.740 142.480 330.100 ;
        RECT 137.670 324.500 137.960 324.790 ;
        RECT 145.390 340.010 145.650 340.270 ;
        RECT 144.870 339.570 145.130 339.830 ;
        RECT 159.050 359.080 159.380 359.410 ;
        RECT 158.420 357.550 158.750 357.880 ;
        RECT 157.860 355.980 158.190 356.310 ;
        RECT 157.240 350.510 157.570 350.840 ;
        RECT 156.610 348.920 156.940 349.250 ;
        RECT 155.990 347.370 156.320 347.700 ;
        RECT 155.390 345.890 155.720 346.220 ;
        RECT 154.750 340.720 155.080 341.050 ;
        RECT 146.040 340.010 146.300 340.270 ;
        RECT 146.410 338.990 146.670 339.250 ;
        RECT 154.080 339.150 154.410 339.480 ;
        RECT 146.330 337.860 146.590 338.120 ;
        RECT 145.730 337.240 145.990 337.500 ;
        RECT 146.340 337.320 146.600 337.580 ;
        RECT 153.460 337.510 153.790 337.840 ;
        RECT 144.200 335.690 144.460 335.950 ;
        RECT 144.890 335.680 145.150 335.940 ;
        RECT 145.370 334.910 145.630 335.170 ;
        RECT 144.490 332.120 144.750 332.540 ;
        RECT 144.450 329.740 144.710 330.100 ;
        RECT 145.070 326.110 145.330 326.440 ;
        RECT 144.040 324.490 144.330 324.780 ;
        RECT 141.350 323.710 141.610 323.970 ;
        RECT 138.040 323.270 138.300 323.530 ;
        RECT 139.140 323.280 139.400 323.540 ;
        RECT 140.230 323.280 140.490 323.540 ;
        RECT 141.360 323.240 141.620 323.500 ;
        RECT 142.880 323.480 143.480 324.080 ;
        RECT 138.590 322.600 138.850 322.860 ;
        RECT 139.690 322.600 139.950 322.860 ;
        RECT 140.790 322.600 141.050 322.860 ;
        RECT 138.590 321.230 138.850 321.490 ;
        RECT 139.690 321.230 139.950 321.490 ;
        RECT 140.790 321.230 141.050 321.490 ;
        RECT 138.040 320.500 138.300 320.760 ;
        RECT 139.140 320.500 139.400 320.760 ;
        RECT 140.230 320.500 140.490 320.760 ;
        RECT 138.030 319.160 138.290 319.420 ;
        RECT 139.140 319.150 139.400 319.410 ;
        RECT 140.230 319.130 140.490 319.390 ;
        RECT 146.390 336.370 146.650 336.630 ;
        RECT 152.780 336.070 153.110 336.400 ;
        RECT 146.080 334.850 146.340 335.110 ;
        RECT 148.740 331.710 149.320 332.420 ;
        RECT 138.590 318.460 138.850 318.720 ;
        RECT 139.690 318.450 139.950 318.710 ;
        RECT 140.780 318.450 141.040 318.710 ;
        RECT 145.660 318.550 145.920 318.890 ;
        RECT 4.890 317.350 5.510 318.050 ;
        RECT 126.750 317.610 127.140 318.000 ;
        RECT 4.690 315.640 5.450 315.990 ;
        RECT 4.300 312.210 4.650 315.200 ;
        RECT 7.570 314.610 10.740 315.030 ;
        RECT 12.040 313.640 12.560 314.160 ;
        RECT 152.750 312.240 153.180 312.670 ;
        RECT 153.400 311.450 153.830 311.880 ;
        RECT 154.070 310.770 154.470 311.170 ;
        RECT 153.900 309.830 154.410 310.340 ;
        RECT 166.420 365.440 166.680 365.700 ;
        RECT 168.520 366.280 168.780 366.540 ;
        RECT 169.460 365.800 169.720 366.060 ;
        RECT 170.500 365.840 170.760 366.100 ;
        RECT 170.560 365.560 170.820 365.820 ;
        RECT 166.420 363.690 166.680 363.950 ;
        RECT 168.520 364.530 168.780 364.790 ;
        RECT 169.460 364.050 169.720 364.310 ;
        RECT 170.500 364.090 170.760 364.350 ;
        RECT 170.560 363.810 170.820 364.070 ;
        RECT 166.420 361.940 166.680 362.200 ;
        RECT 168.520 362.780 168.780 363.040 ;
        RECT 169.460 362.300 169.720 362.560 ;
        RECT 170.500 362.340 170.760 362.600 ;
        RECT 170.560 362.060 170.820 362.320 ;
        RECT 166.420 360.170 166.680 360.430 ;
        RECT 169.460 359.810 169.720 360.070 ;
        RECT 168.520 359.330 168.780 359.590 ;
        RECT 170.560 360.050 170.820 360.310 ;
        RECT 170.500 359.770 170.760 360.030 ;
        RECT 166.420 358.420 166.680 358.680 ;
        RECT 169.460 358.060 169.720 358.320 ;
        RECT 168.520 357.580 168.780 357.840 ;
        RECT 170.560 358.300 170.820 358.560 ;
        RECT 170.500 358.020 170.760 358.280 ;
        RECT 166.420 356.670 166.680 356.930 ;
        RECT 169.460 356.310 169.720 356.570 ;
        RECT 168.520 355.830 168.780 356.090 ;
        RECT 170.560 356.550 170.820 356.810 ;
        RECT 170.500 356.270 170.760 356.530 ;
        RECT 166.420 354.920 166.680 355.180 ;
        RECT 169.460 354.560 169.720 354.820 ;
        RECT 168.520 354.080 168.780 354.340 ;
        RECT 170.560 354.800 170.820 355.060 ;
        RECT 170.500 354.520 170.760 354.780 ;
        RECT 166.420 350.040 166.680 350.300 ;
        RECT 169.460 349.680 169.720 349.940 ;
        RECT 168.520 349.200 168.780 349.460 ;
        RECT 170.560 349.920 170.820 350.180 ;
        RECT 170.500 349.640 170.760 349.900 ;
        RECT 166.420 348.290 166.680 348.550 ;
        RECT 169.460 347.930 169.720 348.190 ;
        RECT 168.520 347.450 168.780 347.710 ;
        RECT 170.560 348.170 170.820 348.430 ;
        RECT 170.500 347.890 170.760 348.150 ;
        RECT 166.420 346.540 166.680 346.800 ;
        RECT 169.460 346.180 169.720 346.440 ;
        RECT 168.520 345.700 168.780 345.960 ;
        RECT 170.560 346.420 170.820 346.680 ;
        RECT 170.500 346.140 170.760 346.400 ;
        RECT 166.420 344.790 166.680 345.050 ;
        RECT 169.460 344.430 169.720 344.690 ;
        RECT 168.520 343.950 168.780 344.210 ;
        RECT 170.560 344.670 170.820 344.930 ;
        RECT 170.500 344.390 170.760 344.650 ;
        RECT 173.660 360.600 173.920 360.860 ;
        RECT 172.570 360.080 172.830 360.340 ;
        RECT 172.570 358.810 172.830 359.070 ;
        RECT 173.660 358.290 173.920 358.550 ;
        RECT 173.660 357.400 173.920 357.660 ;
        RECT 172.570 356.880 172.830 357.140 ;
        RECT 172.570 355.610 172.830 355.870 ;
        RECT 173.660 355.090 173.920 355.350 ;
        RECT 213.200 384.480 213.550 385.240 ;
        RECT 214.910 384.420 215.610 385.040 ;
        RECT 238.360 385.280 241.350 385.630 ;
        RECT 243.560 385.280 245.590 385.610 ;
        RECT 184.150 373.720 185.100 374.130 ;
        RECT 189.570 376.360 190.920 376.780 ;
        RECT 187.160 373.730 187.600 374.170 ;
        RECT 181.410 369.950 181.670 370.210 ;
        RECT 179.530 366.420 179.790 366.680 ;
        RECT 185.000 369.040 185.260 369.300 ;
        RECT 181.870 368.020 182.130 368.280 ;
        RECT 182.290 365.930 182.550 366.190 ;
        RECT 183.350 365.450 183.610 365.710 ;
        RECT 176.070 360.600 176.330 360.860 ;
        RECT 176.070 358.290 176.330 358.550 ;
        RECT 188.170 369.960 188.430 370.220 ;
        RECT 187.730 369.050 187.990 369.310 ;
        RECT 184.990 358.350 185.260 358.620 ;
        RECT 176.070 357.400 176.330 357.660 ;
        RECT 192.960 373.690 193.400 374.130 ;
        RECT 201.290 374.720 201.570 375.160 ;
        RECT 197.510 368.060 198.730 368.320 ;
        RECT 194.270 367.410 194.530 367.670 ;
        RECT 200.600 366.870 200.860 367.130 ;
        RECT 202.940 369.960 203.200 370.220 ;
        RECT 202.050 369.090 202.310 369.350 ;
        RECT 203.160 366.500 203.420 366.760 ;
        RECT 209.460 379.060 209.830 379.430 ;
        RECT 212.170 379.190 212.590 382.360 ;
        RECT 205.610 370.670 205.870 370.940 ;
        RECT 202.050 364.880 202.310 365.140 ;
        RECT 203.070 364.890 203.330 365.150 ;
        RECT 211.200 377.370 211.720 377.890 ;
        RECT 241.790 384.480 242.140 385.240 ;
        RECT 243.500 384.420 244.200 385.040 ;
        RECT 266.950 385.280 269.940 385.630 ;
        RECT 272.150 385.280 274.180 385.610 ;
        RECT 210.280 375.600 210.650 375.970 ;
        RECT 205.820 364.770 206.250 365.200 ;
        RECT 207.390 364.700 207.650 364.960 ;
        RECT 206.730 363.820 206.990 364.080 ;
        RECT 207.380 363.010 207.640 363.270 ;
        RECT 203.160 360.930 203.420 361.190 ;
        RECT 211.050 370.890 211.420 371.260 ;
        RECT 209.910 362.700 210.170 362.960 ;
        RECT 203.150 360.470 203.410 360.730 ;
        RECT 176.070 355.090 176.330 355.350 ;
        RECT 203.150 354.900 203.410 355.160 ;
        RECT 207.620 359.240 207.880 359.500 ;
        RECT 206.730 358.080 206.990 358.340 ;
        RECT 206.730 357.480 206.990 357.740 ;
        RECT 207.620 356.480 207.880 356.740 ;
        RECT 173.640 350.130 173.900 350.390 ;
        RECT 172.550 349.610 172.810 349.870 ;
        RECT 172.550 348.340 172.810 348.600 ;
        RECT 173.640 347.820 173.900 348.080 ;
        RECT 173.640 346.930 173.900 347.190 ;
        RECT 172.550 346.410 172.810 346.670 ;
        RECT 172.550 345.140 172.810 345.400 ;
        RECT 181.630 351.710 181.910 351.990 ;
        RECT 176.050 350.130 176.310 350.390 ;
        RECT 198.980 351.140 199.240 351.400 ;
        RECT 196.660 350.660 196.920 350.920 ;
        RECT 198.460 350.490 198.720 350.750 ;
        RECT 209.950 356.650 210.210 356.910 ;
        RECT 209.470 351.690 209.840 352.060 ;
        RECT 210.240 351.100 210.610 351.470 ;
        RECT 217.600 369.840 218.100 370.340 ;
        RECT 214.380 368.280 214.880 368.780 ;
        RECT 215.330 368.770 215.830 369.270 ;
        RECT 216.410 369.240 216.910 369.740 ;
        RECT 211.930 365.820 212.300 366.190 ;
        RECT 176.050 347.820 176.310 348.080 ;
        RECT 198.460 349.940 198.720 350.200 ;
        RECT 176.050 346.930 176.310 347.190 ;
        RECT 198.460 348.650 198.720 348.910 ;
        RECT 198.460 348.100 198.720 348.360 ;
        RECT 198.460 347.250 198.720 347.510 ;
        RECT 173.640 344.620 173.900 344.880 ;
        RECT 176.050 344.620 176.310 344.880 ;
        RECT 166.380 340.980 166.640 341.240 ;
        RECT 169.420 340.620 169.680 340.880 ;
        RECT 168.480 340.140 168.740 340.400 ;
        RECT 174.260 343.520 174.520 343.930 ;
        RECT 170.520 340.860 170.780 341.120 ;
        RECT 170.460 340.580 170.720 340.840 ;
        RECT 166.380 339.230 166.640 339.490 ;
        RECT 169.420 338.870 169.680 339.130 ;
        RECT 168.480 338.390 168.740 338.650 ;
        RECT 170.520 339.110 170.780 339.370 ;
        RECT 170.460 338.830 170.720 339.090 ;
        RECT 166.380 337.480 166.640 337.740 ;
        RECT 169.420 337.120 169.680 337.380 ;
        RECT 168.480 336.640 168.740 336.900 ;
        RECT 170.520 337.360 170.780 337.620 ;
        RECT 170.460 337.080 170.720 337.340 ;
        RECT 166.380 335.730 166.640 335.990 ;
        RECT 169.420 335.370 169.680 335.630 ;
        RECT 168.480 334.890 168.740 335.150 ;
        RECT 170.520 335.610 170.780 335.870 ;
        RECT 170.460 335.330 170.720 335.590 ;
        RECT 173.670 340.860 173.930 341.120 ;
        RECT 172.580 340.340 172.840 340.600 ;
        RECT 172.580 339.070 172.840 339.330 ;
        RECT 173.670 338.550 173.930 338.810 ;
        RECT 173.670 337.660 173.930 337.920 ;
        RECT 172.580 337.140 172.840 337.400 ;
        RECT 172.580 335.870 172.840 336.130 ;
        RECT 173.670 335.350 173.930 335.610 ;
        RECT 176.080 340.860 176.340 341.120 ;
        RECT 196.420 345.510 196.680 345.770 ;
        RECT 198.460 346.700 198.720 346.960 ;
        RECT 199.520 346.130 199.780 346.390 ;
        RECT 196.420 344.960 196.680 345.220 ;
        RECT 198.460 345.420 198.720 345.680 ;
        RECT 198.460 344.870 198.720 345.130 ;
        RECT 196.420 343.690 196.680 343.950 ;
        RECT 196.420 343.140 196.680 343.400 ;
        RECT 196.420 342.270 196.680 342.530 ;
        RECT 196.420 341.720 196.680 341.980 ;
        RECT 203.450 346.090 203.710 346.350 ;
        RECT 210.980 348.770 211.350 349.140 ;
        RECT 209.250 346.090 209.510 346.350 ;
        RECT 199.900 341.360 200.160 341.620 ;
        RECT 197.600 341.070 197.860 341.330 ;
        RECT 178.660 339.800 178.920 340.060 ;
        RECT 176.080 338.550 176.340 338.810 ;
        RECT 176.080 337.660 176.340 337.920 ;
        RECT 176.080 335.350 176.340 335.610 ;
        RECT 196.420 340.440 196.680 340.700 ;
        RECT 196.420 340.070 196.680 340.150 ;
        RECT 196.420 339.890 196.870 340.070 ;
        RECT 196.610 339.810 196.870 339.890 ;
        RECT 201.620 341.050 201.890 341.310 ;
        RECT 199.880 340.310 200.140 340.570 ;
        RECT 198.540 339.780 198.800 340.040 ;
        RECT 196.590 338.800 196.850 339.060 ;
        RECT 198.020 338.850 198.280 339.110 ;
        RECT 179.290 337.020 179.550 337.280 ;
        RECT 172.080 334.670 172.340 334.930 ;
        RECT 171.540 334.300 171.830 334.590 ;
        RECT 167.100 333.790 167.410 334.100 ;
        RECT 178.690 334.710 178.950 334.970 ;
        RECT 179.720 334.700 179.980 334.960 ;
        RECT 177.290 334.300 177.550 334.560 ;
        RECT 179.260 334.380 179.520 334.640 ;
        RECT 170.910 333.080 171.330 333.500 ;
        RECT 167.060 332.120 167.480 332.540 ;
        RECT 172.970 333.760 173.230 334.020 ;
        RECT 172.520 333.240 172.780 333.500 ;
        RECT 173.610 333.240 173.870 333.500 ;
        RECT 174.710 333.230 174.970 333.490 ;
        RECT 173.070 332.560 173.330 332.820 ;
        RECT 174.160 332.540 174.420 332.800 ;
        RECT 175.270 332.530 175.530 332.790 ;
        RECT 177.270 333.230 177.530 333.490 ;
        RECT 178.370 333.240 178.630 333.500 ;
        RECT 179.460 333.240 179.720 333.500 ;
        RECT 196.590 336.810 196.850 337.070 ;
        RECT 197.550 337.010 197.810 337.270 ;
        RECT 196.640 335.850 196.900 336.110 ;
        RECT 197.050 336.080 197.310 336.340 ;
        RECT 181.500 334.320 181.760 334.580 ;
        RECT 180.300 333.070 180.630 333.400 ;
        RECT 190.340 334.630 190.690 334.980 ;
        RECT 183.490 333.900 183.750 334.160 ;
        RECT 187.530 333.870 187.800 334.140 ;
        RECT 181.450 333.000 181.790 333.340 ;
        RECT 182.330 333.270 182.590 333.530 ;
        RECT 183.420 333.270 183.680 333.530 ;
        RECT 184.520 333.260 184.780 333.520 ;
        RECT 171.590 332.030 171.910 332.350 ;
        RECT 173.070 331.190 173.330 331.450 ;
        RECT 174.160 331.190 174.420 331.450 ;
        RECT 175.260 331.190 175.520 331.450 ;
        RECT 172.510 330.460 172.770 330.720 ;
        RECT 173.610 330.460 173.870 330.720 ;
        RECT 174.710 330.460 174.970 330.720 ;
        RECT 172.510 329.090 172.770 329.350 ;
        RECT 173.610 329.090 173.870 329.350 ;
        RECT 174.710 329.090 174.970 329.350 ;
        RECT 171.940 328.450 172.200 328.710 ;
        RECT 173.070 328.410 173.330 328.670 ;
        RECT 174.160 328.410 174.420 328.670 ;
        RECT 175.260 328.420 175.520 328.680 ;
        RECT 171.950 327.980 172.210 328.240 ;
        RECT 176.710 332.530 176.970 332.790 ;
        RECT 177.820 332.540 178.080 332.800 ;
        RECT 178.910 332.560 179.170 332.820 ;
        RECT 182.880 332.590 183.140 332.850 ;
        RECT 183.970 332.570 184.230 332.830 ;
        RECT 185.080 332.560 185.340 332.820 ;
        RECT 187.080 333.260 187.340 333.520 ;
        RECT 188.180 333.270 188.440 333.530 ;
        RECT 189.270 333.270 189.530 333.530 ;
        RECT 176.720 331.190 176.980 331.450 ;
        RECT 177.820 331.190 178.080 331.450 ;
        RECT 178.910 331.190 179.170 331.450 ;
        RECT 182.880 331.220 183.140 331.480 ;
        RECT 183.970 331.220 184.230 331.480 ;
        RECT 185.070 331.220 185.330 331.480 ;
        RECT 177.270 330.460 177.530 330.720 ;
        RECT 178.370 330.460 178.630 330.720 ;
        RECT 179.470 330.460 179.730 330.720 ;
        RECT 182.320 330.490 182.580 330.750 ;
        RECT 183.420 330.490 183.680 330.750 ;
        RECT 184.520 330.490 184.780 330.750 ;
        RECT 177.270 329.090 177.530 329.350 ;
        RECT 178.370 329.090 178.630 329.350 ;
        RECT 179.470 329.090 179.730 329.350 ;
        RECT 182.320 329.120 182.580 329.380 ;
        RECT 183.420 329.120 183.680 329.380 ;
        RECT 184.520 329.120 184.780 329.380 ;
        RECT 176.720 328.420 176.980 328.680 ;
        RECT 177.820 328.410 178.080 328.670 ;
        RECT 178.910 328.410 179.170 328.670 ;
        RECT 180.040 328.450 180.300 328.710 ;
        RECT 180.030 327.980 180.290 328.240 ;
        RECT 175.610 327.280 175.890 327.560 ;
        RECT 176.350 327.300 176.630 327.580 ;
        RECT 171.690 326.250 172.150 326.710 ;
        RECT 181.750 328.480 182.010 328.740 ;
        RECT 182.880 328.440 183.140 328.700 ;
        RECT 183.970 328.440 184.230 328.700 ;
        RECT 185.070 328.450 185.330 328.710 ;
        RECT 181.760 328.010 182.020 328.270 ;
        RECT 180.070 325.300 180.530 325.760 ;
        RECT 186.520 332.560 186.780 332.820 ;
        RECT 187.630 332.570 187.890 332.830 ;
        RECT 188.720 332.590 188.980 332.850 ;
        RECT 190.380 332.860 190.640 333.180 ;
        RECT 196.370 333.080 196.630 333.420 ;
        RECT 191.800 332.150 192.180 332.530 ;
        RECT 186.530 331.220 186.790 331.480 ;
        RECT 187.630 331.220 187.890 331.480 ;
        RECT 188.720 331.220 188.980 331.480 ;
        RECT 187.080 330.490 187.340 330.750 ;
        RECT 188.180 330.490 188.440 330.750 ;
        RECT 189.280 330.490 189.540 330.750 ;
        RECT 187.080 329.120 187.340 329.380 ;
        RECT 188.180 329.120 188.440 329.380 ;
        RECT 189.280 329.120 189.540 329.380 ;
        RECT 193.460 329.050 193.720 329.310 ;
        RECT 194.560 329.060 194.820 329.320 ;
        RECT 195.650 329.060 195.910 329.320 ;
        RECT 186.530 328.450 186.790 328.710 ;
        RECT 187.630 328.440 187.890 328.700 ;
        RECT 188.720 328.440 188.980 328.700 ;
        RECT 189.850 328.480 190.110 328.740 ;
        RECT 192.900 328.350 193.160 328.610 ;
        RECT 194.010 328.360 194.270 328.620 ;
        RECT 195.100 328.380 195.360 328.640 ;
        RECT 185.420 327.280 185.700 327.560 ;
        RECT 189.840 328.010 190.100 328.270 ;
        RECT 214.880 359.650 215.140 359.910 ;
        RECT 214.910 355.960 215.170 356.220 ;
        RECT 214.240 350.490 214.500 350.750 ;
        RECT 216.060 350.670 216.320 350.930 ;
        RECT 214.240 349.940 214.500 350.200 ;
        RECT 214.240 348.650 214.500 348.910 ;
        RECT 214.240 348.100 214.500 348.360 ;
        RECT 214.240 347.250 214.500 347.510 ;
        RECT 214.240 346.700 214.500 346.960 ;
        RECT 213.180 346.130 213.440 346.390 ;
        RECT 214.240 345.420 214.500 345.680 ;
        RECT 214.240 344.870 214.500 345.130 ;
        RECT 211.910 343.520 212.280 343.930 ;
        RECT 208.030 340.910 208.290 341.170 ;
        RECT 208.180 340.230 208.440 340.490 ;
        RECT 208.180 339.640 208.440 339.900 ;
        RECT 208.030 338.960 208.290 339.220 ;
        RECT 199.880 338.430 200.140 338.690 ;
        RECT 208.030 338.140 208.290 338.400 ;
        RECT 199.750 337.250 200.010 337.510 ;
        RECT 208.180 337.460 208.440 337.720 ;
        RECT 208.180 336.870 208.440 337.130 ;
        RECT 208.030 336.190 208.290 336.450 ;
        RECT 210.170 337.160 210.440 337.430 ;
        RECT 226.410 366.900 227.690 368.180 ;
        RECT 240.760 379.190 241.180 382.360 ;
        RECT 239.790 377.370 240.310 377.890 ;
        RECT 270.380 384.480 270.730 385.240 ;
        RECT 272.090 384.420 272.790 385.040 ;
        RECT 295.540 385.280 298.530 385.630 ;
        RECT 300.740 385.280 302.770 385.610 ;
        RECT 269.350 379.190 269.770 382.360 ;
        RECT 268.380 377.370 268.900 377.890 ;
        RECT 298.970 384.480 299.320 385.240 ;
        RECT 300.680 384.420 301.380 385.040 ;
        RECT 324.130 385.280 327.120 385.630 ;
        RECT 329.330 385.280 331.360 385.610 ;
        RECT 297.940 379.190 298.360 382.360 ;
        RECT 296.970 377.370 297.490 377.890 ;
        RECT 327.560 384.480 327.910 385.240 ;
        RECT 329.270 384.420 329.970 385.040 ;
        RECT 352.720 385.280 355.710 385.630 ;
        RECT 326.530 379.190 326.950 382.360 ;
        RECT 325.560 377.370 326.080 377.890 ;
        RECT 356.150 384.480 356.500 385.240 ;
        RECT 355.120 379.190 355.540 382.360 ;
        RECT 354.150 377.370 354.670 377.890 ;
        RECT 237.680 372.230 238.390 372.940 ;
        RECT 226.900 363.460 227.160 363.880 ;
        RECT 222.900 360.260 223.300 360.660 ;
        RECT 218.130 357.020 218.390 357.280 ;
        RECT 218.190 353.580 218.450 353.840 ;
        RECT 217.510 347.560 218.010 348.060 ;
        RECT 216.430 342.370 216.930 342.840 ;
        RECT 215.300 337.180 215.800 337.680 ;
        RECT 214.250 331.880 214.750 332.380 ;
        RECT 198.520 330.370 198.780 330.870 ;
        RECT 197.980 329.470 198.240 329.970 ;
        RECT 197.510 328.570 197.770 329.070 ;
        RECT 181.500 324.410 181.960 324.870 ;
        RECT 192.910 327.010 193.170 327.270 ;
        RECT 194.010 327.010 194.270 327.270 ;
        RECT 195.100 327.010 195.360 327.270 ;
        RECT 197.030 327.670 197.290 328.170 ;
        RECT 193.460 326.280 193.720 326.540 ;
        RECT 194.560 326.280 194.820 326.540 ;
        RECT 195.660 326.280 195.920 326.540 ;
        RECT 193.460 324.910 193.720 325.170 ;
        RECT 194.560 324.910 194.820 325.170 ;
        RECT 195.660 324.910 195.920 325.170 ;
        RECT 192.910 324.240 193.170 324.500 ;
        RECT 194.010 324.230 194.270 324.490 ;
        RECT 195.100 324.230 195.360 324.490 ;
        RECT 189.890 323.500 190.350 323.960 ;
        RECT 163.820 321.270 164.080 322.390 ;
        RECT 175.930 322.330 177.050 322.350 ;
        RECT 175.190 321.230 177.050 322.330 ;
        RECT 175.190 321.210 176.310 321.230 ;
        RECT 185.000 321.180 186.860 322.370 ;
        RECT 162.140 316.980 162.470 317.310 ;
        RECT 161.520 316.360 161.850 316.690 ;
        RECT 160.890 315.730 161.220 316.060 ;
        RECT 160.290 315.100 160.620 315.430 ;
        RECT 159.650 314.420 159.980 314.750 ;
        RECT 159.050 313.800 159.380 314.130 ;
        RECT 158.450 313.160 158.780 313.490 ;
        RECT 157.870 312.590 158.200 312.920 ;
        RECT 157.290 311.900 157.620 312.230 ;
        RECT 156.640 311.260 156.970 311.590 ;
        RECT 156.000 310.610 156.330 310.950 ;
        RECT 155.420 309.970 155.790 310.340 ;
        RECT 196.230 324.270 196.490 324.530 ;
        RECT 196.220 323.800 196.480 324.060 ;
        RECT 220.490 334.400 220.990 334.900 ;
        RECT 217.620 326.290 218.120 326.790 ;
        RECT 216.430 325.340 216.930 325.800 ;
        RECT 215.300 324.470 215.800 324.930 ;
        RECT 214.370 323.560 214.870 324.020 ;
        RECT 219.910 321.270 220.850 322.390 ;
        RECT 195.700 317.640 196.030 317.970 ;
        RECT 223.880 359.620 224.240 359.980 ;
        RECT 223.930 357.020 224.190 357.280 ;
        RECT 224.800 357.250 225.190 357.640 ;
        RECT 223.890 353.520 224.150 353.780 ;
        RECT 223.890 351.000 224.150 351.260 ;
        RECT 222.960 316.450 223.360 316.850 ;
        RECT 223.870 315.650 224.260 316.040 ;
        RECT 225.630 356.690 226.010 356.950 ;
        RECT 224.800 314.830 225.190 315.220 ;
        RECT 230.730 364.740 230.990 365.170 ;
        RECT 234.150 365.090 234.410 365.350 ;
        RECT 234.450 365.270 234.710 365.530 ;
        RECT 233.840 364.220 234.100 364.480 ;
        RECT 233.440 363.340 233.700 363.600 ;
        RECT 232.180 362.700 232.440 362.960 ;
        RECT 235.340 364.110 235.600 364.370 ;
        RECT 236.280 363.830 236.540 364.090 ;
        RECT 235.340 363.510 235.600 363.770 ;
        RECT 235.710 363.270 235.970 363.530 ;
        RECT 256.110 372.040 259.340 374.100 ;
        RECT 238.920 366.500 239.180 366.760 ;
        RECT 284.700 367.150 286.760 370.450 ;
        RECT 234.450 362.510 234.710 362.770 ;
        RECT 234.840 362.410 235.100 362.670 ;
        RECT 234.150 361.890 234.410 362.150 ;
        RECT 233.840 361.020 234.100 361.280 ;
        RECT 234.840 360.960 235.100 361.220 ;
        RECT 236.750 362.850 237.010 363.110 ;
        RECT 236.700 362.200 236.960 362.460 ;
        RECT 239.000 362.870 239.260 363.130 ;
        RECT 236.700 361.050 236.960 361.310 ;
        RECT 233.440 360.030 233.700 360.400 ;
        RECT 235.710 360.070 235.970 360.360 ;
        RECT 233.840 359.150 234.100 359.410 ;
        RECT 234.440 359.240 234.700 359.500 ;
        RECT 234.840 359.210 235.100 359.470 ;
        RECT 232.440 358.300 232.700 358.560 ;
        RECT 232.590 357.470 232.850 357.730 ;
        RECT 234.150 358.280 234.410 358.540 ;
        RECT 235.330 358.080 235.590 358.340 ;
        RECT 236.750 360.400 237.010 360.660 ;
        RECT 236.750 359.850 237.010 360.110 ;
        RECT 236.700 359.200 236.960 359.460 ;
        RECT 238.920 360.930 239.180 361.190 ;
        RECT 313.290 362.900 316.520 364.960 ;
        RECT 239.050 360.730 239.310 360.910 ;
        RECT 238.910 360.650 239.310 360.730 ;
        RECT 238.910 360.470 239.170 360.650 ;
        RECT 239.040 359.930 239.300 360.190 ;
        RECT 234.840 357.760 235.100 358.020 ;
        RECT 235.330 357.480 235.590 357.740 ;
        RECT 236.270 357.800 236.530 358.060 ;
        RECT 236.700 358.050 236.960 358.310 ;
        RECT 231.760 356.640 232.020 356.900 ;
        RECT 232.150 356.640 232.410 356.900 ;
        RECT 233.440 356.830 233.700 357.090 ;
        RECT 234.320 357.170 234.580 357.430 ;
        RECT 235.710 356.900 235.970 357.160 ;
        RECT 236.750 357.400 237.010 357.660 ;
        RECT 341.880 358.490 345.110 360.540 ;
        RECT 238.960 357.680 239.220 357.940 ;
        RECT 356.220 357.850 358.210 361.080 ;
        RECT 232.880 356.210 233.140 356.470 ;
        RECT 234.440 356.480 234.700 356.740 ;
        RECT 232.490 355.360 232.750 355.620 ;
        RECT 233.840 355.950 234.100 356.210 ;
        RECT 234.150 355.080 234.410 355.340 ;
        RECT 236.740 356.820 237.000 357.080 ;
        RECT 236.690 356.170 236.950 356.430 ;
        RECT 238.990 356.840 239.250 357.100 ;
        RECT 236.690 355.020 236.950 355.280 ;
        RECT 236.740 354.370 237.000 354.630 ;
        RECT 236.740 353.820 237.000 354.080 ;
        RECT 236.690 353.170 236.950 353.430 ;
        RECT 238.910 354.900 239.170 355.160 ;
        RECT 239.040 354.620 239.300 354.880 ;
        RECT 264.480 356.870 266.700 357.190 ;
        RECT 239.030 353.900 239.290 354.160 ;
        RECT 232.430 352.270 232.690 352.530 ;
        RECT 237.490 352.440 238.200 353.150 ;
        RECT 236.690 352.020 236.950 352.280 ;
        RECT 232.580 351.440 232.840 351.700 ;
        RECT 234.330 351.130 234.600 351.390 ;
        RECT 236.740 351.370 237.000 351.630 ;
        RECT 238.950 351.650 239.210 351.910 ;
        RECT 231.750 350.610 232.010 350.870 ;
        RECT 232.870 350.180 233.130 350.440 ;
        RECT 232.480 349.330 232.740 349.590 ;
        RECT 233.290 334.390 233.800 334.900 ;
        RECT 347.670 329.260 349.760 332.490 ;
        RECT 232.650 324.720 232.910 324.980 ;
        RECT 264.320 326.480 268.600 327.570 ;
        RECT 232.650 324.050 232.910 324.310 ;
        RECT 232.660 322.670 232.920 322.930 ;
        RECT 227.820 319.430 228.080 319.690 ;
        RECT 232.660 321.060 232.920 321.320 ;
        RECT 232.650 319.450 232.910 319.710 ;
        RECT 232.660 317.830 232.920 318.090 ;
        RECT 232.650 316.220 232.910 316.480 ;
        RECT 225.620 314.040 226.000 314.420 ;
        RECT 232.240 314.570 232.500 314.830 ;
        RECT 232.650 313.020 232.910 313.280 ;
        RECT 229.410 311.310 229.670 311.570 ;
        RECT 230.350 311.310 230.610 311.570 ;
        RECT 231.300 311.290 231.560 311.550 ;
        RECT 232.610 311.310 232.870 311.570 ;
        RECT 27.730 301.390 29.810 304.620 ;
        RECT 4.320 288.820 4.650 290.850 ;
        RECT 4.890 288.760 5.510 289.460 ;
        RECT 4.690 287.050 5.450 287.400 ;
        RECT 4.300 283.620 4.650 286.610 ;
        RECT 7.570 286.020 10.740 286.440 ;
        RECT 12.040 285.050 12.560 285.570 ;
        RECT 32.360 272.800 34.440 276.030 ;
        RECT 4.320 260.230 4.650 262.260 ;
        RECT 4.890 260.170 5.510 260.870 ;
        RECT 4.690 258.460 5.450 258.810 ;
        RECT 4.300 255.030 4.650 258.020 ;
        RECT 7.570 257.430 10.740 257.850 ;
        RECT 12.040 256.460 12.560 256.980 ;
        RECT 36.770 244.210 38.850 247.440 ;
        RECT 4.320 231.640 4.650 233.670 ;
        RECT 4.890 231.580 5.510 232.280 ;
        RECT 4.690 229.870 5.450 230.220 ;
        RECT 4.300 226.440 4.650 229.430 ;
        RECT 7.570 228.840 10.740 229.260 ;
        RECT 12.040 227.870 12.560 228.390 ;
        RECT 41.110 215.620 43.190 218.850 ;
        RECT 4.320 203.050 4.650 205.080 ;
        RECT 4.890 202.990 5.510 203.690 ;
        RECT 4.690 201.280 5.450 201.630 ;
        RECT 4.300 197.850 4.650 200.840 ;
        RECT 7.570 200.250 10.740 200.670 ;
        RECT 12.040 199.280 12.560 199.800 ;
        RECT 4.320 174.460 4.650 176.490 ;
        RECT 4.890 174.400 5.510 175.100 ;
        RECT 4.690 172.690 5.450 173.040 ;
        RECT 4.300 169.260 4.650 172.250 ;
        RECT 7.570 171.660 10.740 172.080 ;
        RECT 12.040 170.690 12.560 171.210 ;
        RECT 343.420 300.670 345.510 303.900 ;
        RECT 339.440 272.080 341.530 275.310 ;
        RECT 335.190 243.490 337.280 246.720 ;
        RECT 331.250 214.900 333.340 218.130 ;
        RECT 49.650 158.440 51.730 161.670 ;
        RECT 263.500 160.540 267.920 164.960 ;
        RECT 4.320 145.870 4.650 147.900 ;
        RECT 4.890 145.810 5.510 146.510 ;
        RECT 4.690 144.100 5.450 144.450 ;
        RECT 4.300 140.670 4.650 143.660 ;
        RECT 7.570 143.070 10.740 143.490 ;
        RECT 12.040 142.100 12.560 142.620 ;
        RECT 4.320 117.280 4.650 119.310 ;
        RECT 4.890 117.220 5.510 117.920 ;
        RECT 4.690 115.510 5.450 115.860 ;
        RECT 4.300 112.080 4.650 115.070 ;
        RECT 7.570 114.480 10.740 114.900 ;
        RECT 12.040 113.510 12.560 114.030 ;
        RECT 58.270 101.260 60.350 104.490 ;
        RECT 4.320 88.690 4.650 90.720 ;
        RECT 4.890 88.630 5.510 89.330 ;
        RECT 4.690 86.920 5.450 87.270 ;
        RECT 4.300 83.490 4.650 86.480 ;
        RECT 7.570 85.890 10.740 86.310 ;
        RECT 12.040 84.920 12.560 85.440 ;
        RECT 62.240 72.670 64.320 75.900 ;
        RECT 4.320 60.100 4.650 62.130 ;
        RECT 4.890 60.040 5.510 60.740 ;
        RECT 4.690 58.330 5.450 58.680 ;
        RECT 4.300 54.900 4.650 57.890 ;
        RECT 7.570 57.300 10.740 57.720 ;
        RECT 12.040 56.330 12.560 56.850 ;
        RECT 66.680 44.080 68.760 47.310 ;
        RECT 4.320 31.510 4.650 33.540 ;
        RECT 4.890 31.450 5.510 32.150 ;
        RECT 4.690 29.740 5.450 30.090 ;
        RECT 4.300 26.310 4.650 29.300 ;
        RECT 7.570 28.710 10.740 29.130 ;
        RECT 12.040 27.740 12.560 28.260 ;
        RECT 70.980 15.490 73.060 18.720 ;
        RECT 4.320 2.920 4.650 4.950 ;
        RECT 4.890 2.860 5.510 3.560 ;
      LAYER met2 ;
        RECT 183.470 380.050 184.110 382.490 ;
        RECT 129.150 379.480 184.620 380.050 ;
        RECT 212.060 379.480 212.700 382.490 ;
        RECT 240.650 380.780 241.290 382.490 ;
        RECT 240.270 379.480 241.290 380.780 ;
        RECT 269.240 379.480 269.880 382.490 ;
        RECT 297.830 379.480 298.470 382.490 ;
        RECT 326.420 379.480 327.060 382.490 ;
        RECT 355.010 379.480 355.650 382.490 ;
        RECT 129.150 378.720 357.260 379.480 ;
        RECT 129.150 378.650 362.510 378.720 ;
        RECT 157.130 378.080 362.510 378.650 ;
        RECT 182.570 377.950 185.200 378.080 ;
        RECT 211.160 377.950 213.790 378.080 ;
        RECT 239.750 377.950 242.380 378.080 ;
        RECT 268.340 377.950 270.970 378.080 ;
        RECT 296.930 377.950 299.560 378.080 ;
        RECT 325.520 377.950 328.150 378.080 ;
        RECT 125.400 377.800 127.880 377.810 ;
        RECT 125.400 377.410 129.350 377.800 ;
        RECT 127.670 377.040 129.350 377.410 ;
        RECT 145.330 377.710 146.080 377.720 ;
        RECT 145.330 377.410 146.950 377.710 ;
        RECT 145.330 377.240 145.570 377.410 ;
        RECT 146.650 377.190 146.950 377.410 ;
        RECT 182.570 377.440 185.120 377.950 ;
        RECT 211.160 377.440 213.710 377.950 ;
        RECT 239.750 377.440 242.300 377.950 ;
        RECT 268.340 377.440 270.890 377.950 ;
        RECT 296.930 377.440 299.480 377.950 ;
        RECT 325.520 377.440 328.070 377.950 ;
        RECT 354.110 377.440 362.510 378.080 ;
        RECT 182.570 377.370 183.190 377.440 ;
        RECT 211.160 377.370 211.780 377.440 ;
        RECT 239.750 377.370 240.370 377.440 ;
        RECT 268.340 377.370 268.960 377.440 ;
        RECT 296.930 377.370 297.550 377.440 ;
        RECT 325.520 377.370 326.140 377.440 ;
        RECT 354.110 377.370 354.730 377.440 ;
        RECT 355.840 377.320 362.510 377.440 ;
        RECT 119.990 376.280 120.310 376.540 ;
        RECT 122.850 376.440 123.170 376.590 ;
        RECT 120.370 376.200 123.260 376.440 ;
        RECT 210.230 375.970 210.670 375.990 ;
        RECT 240.270 375.970 241.130 376.650 ;
        RECT 210.230 375.600 241.130 375.970 ;
        RECT 210.230 375.580 210.670 375.600 ;
        RECT 122.630 374.660 122.950 374.980 ;
        RECT 122.650 373.620 122.920 374.660 ;
        RECT 240.270 374.550 241.130 375.600 ;
        RECT 120.130 373.610 122.920 373.620 ;
        RECT 119.470 373.390 122.920 373.610 ;
        RECT 119.470 373.380 122.400 373.390 ;
        RECT 254.960 372.810 259.760 374.900 ;
        RECT 211.010 371.260 211.430 371.280 ;
        RECT 240.240 371.260 241.100 372.560 ;
        RECT 164.270 370.940 164.570 371.000 ;
        RECT 205.590 370.940 205.890 370.970 ;
        RECT 164.270 370.710 205.960 370.940 ;
        RECT 211.010 370.890 241.100 371.260 ;
        RECT 211.010 370.870 211.430 370.890 ;
        RECT 164.270 370.680 164.570 370.710 ;
        RECT 205.590 370.630 205.890 370.710 ;
        RECT 240.240 370.460 241.100 370.890 ;
        RECT 243.260 370.750 259.810 372.810 ;
        RECT 361.100 371.810 362.500 377.320 ;
        RECT 98.460 369.880 99.080 369.900 ;
        RECT 98.460 369.510 127.610 369.880 ;
        RECT 98.460 369.440 99.080 369.510 ;
        RECT 125.100 369.400 125.610 369.510 ;
        RECT 125.100 369.110 128.200 369.400 ;
        RECT 125.610 369.100 128.200 369.110 ;
        RECT 284.550 368.680 287.860 370.740 ;
        RECT 168.520 367.520 168.780 368.320 ;
        RECT 169.440 367.810 169.760 367.820 ;
        RECT 169.430 367.800 169.760 367.810 ;
        RECT 170.470 367.800 170.790 367.850 ;
        RECT 169.430 367.600 174.750 367.800 ;
        RECT 194.260 367.670 194.540 367.690 ;
        RECT 169.430 367.550 169.760 367.600 ;
        RECT 170.470 367.590 170.790 367.600 ;
        RECT 169.440 367.530 169.760 367.550 ;
        RECT 170.520 367.520 170.860 367.580 ;
        RECT 166.250 367.160 166.710 367.480 ;
        RECT 168.420 367.300 170.860 367.520 ;
        RECT 174.550 367.100 174.750 367.600 ;
        RECT 194.240 367.640 194.560 367.670 ;
        RECT 226.380 367.640 227.720 368.180 ;
        RECT 194.240 367.430 227.720 367.640 ;
        RECT 194.240 367.410 194.560 367.430 ;
        RECT 194.260 367.390 194.540 367.410 ;
        RECT 200.570 367.100 200.880 367.160 ;
        RECT 163.470 366.920 163.570 366.990 ;
        RECT 163.080 366.750 163.640 366.920 ;
        RECT 174.550 366.900 200.880 367.100 ;
        RECT 226.380 366.900 227.720 367.430 ;
        RECT 200.570 366.840 200.880 366.900 ;
        RECT 238.890 366.790 239.200 366.800 ;
        RECT 240.240 366.790 241.100 368.170 ;
        RECT 162.110 366.190 162.500 366.280 ;
        RECT 163.080 366.190 163.250 366.750 ;
        RECT 163.470 366.670 163.570 366.750 ;
        RECT 179.500 366.630 179.820 366.680 ;
        RECT 162.110 366.020 163.260 366.190 ;
        RECT 168.520 365.770 168.780 366.570 ;
        RECT 174.500 366.430 179.870 366.630 ;
        RECT 238.890 366.610 241.370 366.790 ;
        RECT 243.260 366.620 288.180 368.680 ;
        RECT 238.890 366.470 239.200 366.610 ;
        RECT 169.440 366.060 169.760 366.070 ;
        RECT 169.430 366.050 169.760 366.060 ;
        RECT 170.470 366.050 170.790 366.100 ;
        RECT 174.500 366.050 174.700 366.430 ;
        RECT 179.500 366.420 179.820 366.430 ;
        RECT 208.140 366.370 208.460 366.390 ;
        RECT 182.260 366.190 182.570 366.200 ;
        RECT 205.730 366.190 205.810 366.370 ;
        RECT 208.140 366.190 217.250 366.370 ;
        RECT 225.080 366.190 234.200 366.370 ;
        RECT 240.240 366.190 241.100 366.610 ;
        RECT 182.260 366.160 182.580 366.190 ;
        RECT 169.430 365.850 174.700 366.050 ;
        RECT 175.010 365.960 182.580 366.160 ;
        RECT 169.430 365.800 169.760 365.850 ;
        RECT 170.470 365.840 170.790 365.850 ;
        RECT 169.440 365.780 169.760 365.800 ;
        RECT 170.520 365.770 170.860 365.830 ;
        RECT 145.080 365.590 145.370 365.610 ;
        RECT 101.810 365.460 102.290 365.490 ;
        RECT 27.100 364.260 29.740 365.440 ;
        RECT 101.810 365.080 127.600 365.460 ;
        RECT 132.630 365.190 145.390 365.590 ;
        RECT 166.250 365.410 166.710 365.730 ;
        RECT 168.420 365.550 170.860 365.770 ;
        RECT 101.810 365.060 102.290 365.080 ;
        RECT 27.020 362.500 127.330 364.260 ;
        RECT 132.630 362.500 133.030 365.190 ;
        RECT 145.080 365.180 145.370 365.190 ;
        RECT 163.470 365.090 163.570 365.240 ;
        RECT 143.060 364.620 143.660 364.790 ;
        RECT 143.730 364.700 144.040 365.030 ;
        RECT 144.820 364.800 145.130 365.040 ;
        RECT 163.080 364.920 163.640 365.090 ;
        RECT 144.820 364.710 145.140 364.800 ;
        RECT 144.920 364.630 145.140 364.710 ;
        RECT 161.510 364.650 161.840 364.660 ;
        RECT 161.490 364.550 161.860 364.650 ;
        RECT 163.080 364.550 163.250 364.920 ;
        RECT 136.430 364.510 136.800 364.520 ;
        RECT 134.640 364.280 136.800 364.510 ;
        RECT 161.490 364.380 163.250 364.550 ;
        RECT 141.890 364.340 141.960 364.380 ;
        RECT 141.890 364.280 142.030 364.340 ;
        RECT 145.090 364.290 145.410 364.340 ;
        RECT 134.640 364.150 142.060 364.280 ;
        RECT 134.640 363.450 135.260 364.150 ;
        RECT 136.430 364.110 142.060 364.150 ;
        RECT 143.870 364.120 145.470 364.290 ;
        RECT 161.490 364.270 161.860 364.380 ;
        RECT 163.080 364.370 163.250 364.380 ;
        RECT 142.190 363.790 142.500 364.120 ;
        RECT 145.090 364.080 145.410 364.120 ;
        RECT 144.830 363.810 145.140 364.050 ;
        RECT 168.520 364.020 168.780 364.820 ;
        RECT 169.440 364.310 169.760 364.320 ;
        RECT 169.430 364.300 169.760 364.310 ;
        RECT 170.470 364.300 170.790 364.350 ;
        RECT 175.010 364.300 175.210 365.960 ;
        RECT 182.260 365.930 182.580 365.960 ;
        RECT 211.890 366.070 241.100 366.190 ;
        RECT 182.260 365.920 182.570 365.930 ;
        RECT 211.890 365.820 240.990 366.070 ;
        RECT 211.890 365.790 212.300 365.820 ;
        RECT 183.320 365.680 183.640 365.720 ;
        RECT 169.430 364.100 175.210 364.300 ;
        RECT 175.560 365.480 183.720 365.680 ;
        RECT 169.430 364.050 169.760 364.100 ;
        RECT 170.470 364.090 170.790 364.100 ;
        RECT 169.440 364.030 169.760 364.050 ;
        RECT 170.520 364.020 170.860 364.080 ;
        RECT 143.070 363.630 143.670 363.800 ;
        RECT 144.830 363.720 145.150 363.810 ;
        RECT 144.930 363.640 145.150 363.720 ;
        RECT 166.250 363.660 166.710 363.980 ;
        RECT 168.420 363.800 170.860 364.020 ;
        RECT 136.430 363.450 136.800 363.490 ;
        RECT 27.020 362.100 133.030 362.500 ;
        RECT 134.110 363.360 136.800 363.450 ;
        RECT 145.090 363.370 145.410 363.420 ;
        RECT 134.110 363.190 142.060 363.360 ;
        RECT 143.870 363.200 145.470 363.370 ;
        RECT 163.470 363.360 163.570 363.490 ;
        RECT 134.110 363.080 136.800 363.190 ;
        RECT 134.110 362.970 135.260 363.080 ;
        RECT 134.110 362.520 135.220 362.970 ;
        RECT 142.170 362.870 142.480 363.200 ;
        RECT 145.090 363.160 145.410 363.200 ;
        RECT 163.040 363.190 163.640 363.360 ;
        RECT 160.910 363.070 161.300 363.170 ;
        RECT 163.040 363.070 163.210 363.190 ;
        RECT 163.470 363.170 163.570 363.190 ;
        RECT 143.070 362.640 143.670 362.810 ;
        RECT 143.740 362.720 144.050 363.050 ;
        RECT 144.830 362.820 145.140 363.060 ;
        RECT 160.910 362.900 163.210 363.070 ;
        RECT 144.830 362.730 145.150 362.820 ;
        RECT 160.910 362.800 161.300 362.900 ;
        RECT 144.930 362.650 145.150 362.730 ;
        RECT 136.430 362.520 136.800 362.560 ;
        RECT 134.110 362.440 136.800 362.520 ;
        RECT 145.060 362.450 145.380 362.500 ;
        RECT 134.110 362.410 142.060 362.440 ;
        RECT 134.110 362.270 142.100 362.410 ;
        RECT 143.870 362.280 145.470 362.450 ;
        RECT 134.110 362.150 136.800 362.270 ;
        RECT 134.110 362.110 135.010 362.150 ;
        RECT 27.020 362.010 127.330 362.100 ;
        RECT 14.870 359.920 17.760 361.880 ;
        RECT 27.100 361.840 29.740 362.010 ;
        RECT 98.340 361.590 98.960 361.680 ;
        RECT 125.070 361.590 126.340 362.010 ;
        RECT 98.340 361.180 127.280 361.590 ;
        RECT 98.340 361.090 98.960 361.180 ;
        RECT 101.810 360.690 102.350 360.720 ;
        RECT 101.810 360.280 127.240 360.690 ;
        RECT 101.810 360.240 102.350 360.280 ;
        RECT 14.840 358.060 126.960 359.920 ;
        RECT 125.500 357.560 126.770 358.060 ;
        RECT 134.110 357.560 134.480 362.110 ;
        RECT 142.150 361.880 142.460 362.210 ;
        RECT 143.170 361.810 143.540 362.000 ;
        RECT 143.650 361.930 143.960 362.260 ;
        RECT 145.060 362.240 145.380 362.280 ;
        RECT 168.520 362.270 168.780 363.070 ;
        RECT 169.440 362.560 169.760 362.570 ;
        RECT 169.430 362.550 169.760 362.560 ;
        RECT 170.470 362.550 170.790 362.600 ;
        RECT 175.560 362.550 175.760 365.480 ;
        RECT 183.320 365.440 183.640 365.480 ;
        RECT 234.420 365.350 234.730 365.570 ;
        RECT 234.120 365.240 236.610 365.350 ;
        RECT 205.800 365.170 206.270 365.230 ;
        RECT 234.120 365.220 234.440 365.240 ;
        RECT 234.580 365.220 236.610 365.240 ;
        RECT 230.700 365.180 230.990 365.190 ;
        RECT 230.700 365.170 231.000 365.180 ;
        RECT 233.340 365.170 236.610 365.220 ;
        RECT 241.230 365.170 241.680 365.190 ;
        RECT 205.800 364.740 241.690 365.170 ;
        RECT 207.370 364.670 217.250 364.740 ;
        RECT 230.700 364.730 231.000 364.740 ;
        RECT 230.700 364.710 230.990 364.730 ;
        RECT 207.540 364.640 217.250 364.670 ;
        RECT 312.940 364.600 316.870 365.050 ;
        RECT 233.810 364.240 234.120 364.520 ;
        RECT 233.340 364.190 234.120 364.240 ;
        RECT 169.430 362.350 175.760 362.550 ;
        RECT 178.710 363.680 179.000 363.860 ;
        RECT 206.700 363.820 207.020 364.080 ;
        RECT 233.340 364.040 233.910 364.190 ;
        RECT 235.310 364.110 235.630 364.370 ;
        RECT 236.250 364.010 236.570 364.090 ;
        RECT 240.730 364.060 241.090 364.070 ;
        RECT 207.090 363.910 217.250 363.950 ;
        RECT 207.080 363.720 217.250 363.910 ;
        RECT 226.880 363.880 227.180 363.900 ;
        RECT 235.260 363.880 236.570 364.010 ;
        RECT 240.170 363.880 241.090 364.060 ;
        RECT 226.870 363.780 241.090 363.880 ;
        RECT 169.430 362.300 169.760 362.350 ;
        RECT 170.470 362.340 170.790 362.350 ;
        RECT 169.440 362.280 169.760 362.300 ;
        RECT 170.520 362.270 170.860 362.330 ;
        RECT 144.950 361.830 145.260 362.160 ;
        RECT 166.250 361.910 166.710 362.230 ;
        RECT 168.420 362.050 170.860 362.270 ;
        RECT 163.470 361.640 163.570 361.740 ;
        RECT 143.480 361.580 143.800 361.640 ;
        RECT 135.590 361.420 142.080 361.440 ;
        RECT 125.500 357.190 134.480 357.560 ;
        RECT 135.300 361.250 142.080 361.420 ;
        RECT 143.170 361.390 143.800 361.580 ;
        RECT 143.480 361.320 143.800 361.390 ;
        RECT 160.270 361.470 160.660 361.560 ;
        RECT 163.210 361.470 163.640 361.640 ;
        RECT 160.270 361.300 163.840 361.470 ;
        RECT 135.300 361.070 136.800 361.250 ;
        RECT 160.270 361.210 160.660 361.300 ;
        RECT 163.210 361.280 163.380 361.300 ;
        RECT 135.300 360.480 135.960 361.070 ;
        RECT 136.430 361.030 136.800 361.070 ;
        RECT 143.170 360.820 143.540 361.010 ;
        RECT 144.950 360.840 145.260 361.170 ;
        RECT 159.630 360.900 160.020 361.010 ;
        RECT 163.470 360.900 163.570 360.950 ;
        RECT 159.630 360.730 163.840 360.900 ;
        RECT 173.630 360.840 173.950 360.890 ;
        RECT 176.040 360.840 176.360 360.860 ;
        RECT 178.710 360.840 178.890 363.680 ;
        RECT 226.870 363.460 241.130 363.780 ;
        RECT 226.880 363.440 227.180 363.460 ;
        RECT 233.410 363.410 233.730 363.460 ;
        RECT 235.680 363.410 236.000 363.460 ;
        RECT 233.030 363.340 233.730 363.410 ;
        RECT 207.360 362.980 207.670 363.310 ;
        RECT 230.400 363.060 230.450 363.260 ;
        RECT 233.030 363.210 233.640 363.340 ;
        RECT 235.540 363.270 236.000 363.410 ;
        RECT 235.540 363.210 235.910 363.270 ;
        RECT 237.720 363.210 237.790 363.410 ;
        RECT 209.880 362.970 210.200 362.980 ;
        RECT 207.530 362.860 217.250 362.970 ;
        RECT 232.150 362.860 232.470 362.980 ;
        RECT 207.530 362.780 232.470 362.860 ;
        RECT 209.880 362.680 232.470 362.780 ;
        RECT 233.250 362.730 233.560 362.970 ;
        RECT 236.720 362.920 237.030 363.150 ;
        RECT 238.970 362.920 239.280 363.170 ;
        RECT 240.170 363.120 241.130 363.460 ;
        RECT 236.590 362.840 239.280 362.920 ;
        RECT 234.420 362.590 234.730 362.810 ;
        RECT 234.810 362.590 235.120 362.710 ;
        RECT 236.590 362.690 239.130 362.840 ;
        RECT 209.680 362.320 209.760 362.500 ;
        RECT 234.420 362.480 236.610 362.590 ;
        RECT 234.570 362.440 236.610 362.480 ;
        RECT 233.900 362.430 236.610 362.440 ;
        RECT 233.030 362.380 236.610 362.430 ;
        RECT 230.400 362.080 230.460 362.280 ;
        RECT 233.030 362.230 235.910 362.380 ;
        RECT 233.900 362.220 235.020 362.230 ;
        RECT 234.120 362.120 234.440 362.150 ;
        RECT 234.120 362.020 234.580 362.120 ;
        RECT 235.090 362.080 235.160 362.230 ;
        RECT 236.230 362.060 236.560 362.270 ;
        RECT 236.670 362.170 236.980 362.500 ;
        RECT 203.060 361.250 203.660 361.810 ;
        RECT 206.660 361.640 211.890 361.870 ;
        RECT 212.260 361.640 221.410 361.870 ;
        RECT 233.340 361.820 235.220 362.020 ;
        RECT 234.310 361.760 234.580 361.820 ;
        RECT 240.230 361.690 241.130 363.120 ;
        RECT 243.260 362.540 316.870 364.600 ;
        RECT 312.940 362.530 316.870 362.540 ;
        RECT 221.120 361.540 221.410 361.640 ;
        RECT 229.100 361.540 230.240 361.620 ;
        RECT 205.730 361.320 205.810 361.500 ;
        RECT 208.040 361.490 208.200 361.510 ;
        RECT 221.120 361.490 230.240 361.540 ;
        RECT 230.400 361.490 230.460 361.550 ;
        RECT 234.140 361.490 234.300 361.510 ;
        RECT 208.040 361.440 217.250 361.490 ;
        RECT 208.160 361.340 217.250 361.440 ;
        RECT 221.120 361.440 234.300 361.490 ;
        RECT 221.120 361.410 234.180 361.440 ;
        RECT 221.120 361.400 235.020 361.410 ;
        RECT 235.090 361.400 235.160 361.550 ;
        RECT 221.120 361.340 235.910 361.400 ;
        RECT 221.120 361.330 221.410 361.340 ;
        RECT 232.570 361.260 232.920 361.340 ;
        RECT 203.140 361.080 203.450 361.220 ;
        RECT 233.030 361.200 235.910 361.340 ;
        RECT 236.230 361.240 236.560 361.450 ;
        RECT 200.970 360.900 203.450 361.080 ;
        RECT 233.810 361.190 235.120 361.200 ;
        RECT 233.810 361.040 234.120 361.190 ;
        RECT 203.140 360.890 203.450 360.900 ;
        RECT 143.480 360.590 143.800 360.650 ;
        RECT 159.630 360.630 160.020 360.730 ;
        RECT 163.470 360.630 163.570 360.730 ;
        RECT 173.630 360.670 178.890 360.840 ;
        RECT 206.670 360.820 211.890 361.040 ;
        RECT 212.260 360.820 220.470 361.040 ;
        RECT 233.340 360.990 234.120 361.040 ;
        RECT 203.130 360.760 203.440 360.770 ;
        RECT 173.630 360.650 176.360 360.670 ;
        RECT 135.300 360.290 142.080 360.480 ;
        RECT 143.170 360.400 143.800 360.590 ;
        RECT 173.630 360.570 173.950 360.650 ;
        RECT 176.040 360.600 176.360 360.650 ;
        RECT 200.960 360.580 203.440 360.760 ;
        RECT 143.480 360.330 143.800 360.400 ;
        RECT 135.300 360.110 136.800 360.290 ;
        RECT 135.300 360.100 135.970 360.110 ;
        RECT 135.300 360.060 135.960 360.100 ;
        RECT 136.430 360.070 136.800 360.110 ;
        RECT 125.500 356.560 126.770 357.190 ;
        RECT 23.730 353.400 127.250 355.480 ;
        RECT 23.730 333.290 25.810 353.400 ;
        RECT 125.440 352.800 126.710 353.400 ;
        RECT 135.300 352.800 135.670 360.060 ;
        RECT 143.170 359.830 143.540 360.020 ;
        RECT 144.950 359.850 145.260 360.180 ;
        RECT 166.250 360.140 166.710 360.460 ;
        RECT 203.130 360.440 203.440 360.580 ;
        RECT 168.420 360.100 170.860 360.320 ;
        RECT 143.480 359.600 143.800 359.660 ;
        RECT 125.440 352.430 135.670 352.800 ;
        RECT 136.430 359.330 142.080 359.520 ;
        RECT 143.170 359.410 143.800 359.600 ;
        RECT 143.480 359.340 143.800 359.410 ;
        RECT 159.020 359.330 159.410 359.430 ;
        RECT 125.440 351.810 126.710 352.430 ;
        RECT 27.890 348.520 127.730 350.600 ;
        RECT 23.660 329.920 26.000 333.290 ;
        RECT 23.730 329.050 25.810 329.920 ;
        RECT 27.890 304.690 29.970 348.520 ;
        RECT 125.500 347.960 126.770 348.520 ;
        RECT 136.430 347.960 136.800 359.330 ;
        RECT 159.020 359.160 163.840 359.330 ;
        RECT 168.520 359.300 168.780 360.100 ;
        RECT 169.440 360.070 169.760 360.090 ;
        RECT 169.430 360.020 169.760 360.070 ;
        RECT 170.520 360.040 170.860 360.100 ;
        RECT 172.280 360.060 172.870 360.360 ;
        RECT 208.130 360.160 217.250 360.340 ;
        RECT 172.280 360.040 172.630 360.060 ;
        RECT 170.470 360.020 170.790 360.030 ;
        RECT 172.280 360.020 172.480 360.040 ;
        RECT 169.430 359.820 172.480 360.020 ;
        RECT 169.430 359.810 169.760 359.820 ;
        RECT 169.440 359.800 169.760 359.810 ;
        RECT 170.470 359.770 170.790 359.820 ;
        RECT 207.600 359.320 207.910 359.540 ;
        RECT 205.720 359.310 207.910 359.320 ;
        RECT 159.020 359.060 159.410 359.160 ;
        RECT 163.290 359.000 163.640 359.160 ;
        RECT 205.720 359.100 217.250 359.310 ;
        RECT 207.030 359.090 217.250 359.100 ;
        RECT 172.530 359.020 172.870 359.090 ;
        RECT 163.470 358.880 163.570 359.000 ;
        RECT 172.230 358.790 172.870 359.020 ;
        RECT 178.270 358.790 179.000 358.970 ;
        RECT 220.250 358.940 220.470 360.820 ;
        RECT 221.190 360.770 229.180 360.970 ;
        RECT 233.340 360.840 233.910 360.990 ;
        RECT 234.380 360.860 234.600 361.190 ;
        RECT 234.810 360.920 235.120 361.190 ;
        RECT 236.670 361.010 236.980 361.340 ;
        RECT 238.890 361.080 239.200 361.220 ;
        RECT 238.890 360.900 241.370 361.080 ;
        RECT 238.890 360.890 239.330 360.900 ;
        RECT 234.400 360.850 234.600 360.860 ;
        RECT 239.020 360.780 239.330 360.890 ;
        RECT 222.870 360.560 223.330 360.690 ;
        RECT 228.960 360.640 229.180 360.770 ;
        RECT 236.850 360.760 239.500 360.780 ;
        RECT 236.850 360.690 241.360 360.760 ;
        RECT 228.960 360.560 230.240 360.640 ;
        RECT 222.870 360.440 230.240 360.560 ;
        RECT 222.870 360.360 229.450 360.440 ;
        RECT 230.400 360.370 230.450 360.570 ;
        RECT 234.600 360.440 236.320 360.640 ;
        RECT 236.720 360.580 241.360 360.690 ;
        RECT 236.720 360.550 239.500 360.580 ;
        RECT 233.030 360.400 233.640 360.420 ;
        RECT 222.870 360.240 223.330 360.360 ;
        RECT 228.960 360.340 229.180 360.360 ;
        RECT 233.030 360.340 233.730 360.400 ;
        RECT 234.600 360.360 236.310 360.440 ;
        RECT 236.720 360.360 237.030 360.550 ;
        RECT 237.670 360.420 237.780 360.520 ;
        RECT 238.880 360.440 239.190 360.550 ;
        RECT 225.070 360.160 234.190 360.340 ;
        RECT 235.540 360.220 236.000 360.360 ;
        RECT 235.680 360.210 236.000 360.220 ;
        RECT 227.780 360.090 228.000 360.100 ;
        RECT 221.200 359.910 228.030 360.090 ;
        RECT 228.960 360.050 229.180 360.160 ;
        RECT 228.930 360.010 229.180 360.050 ;
        RECT 228.930 359.910 229.190 360.010 ;
        RECT 221.200 359.840 230.240 359.910 ;
        RECT 230.400 359.860 230.450 360.060 ;
        RECT 233.030 360.030 233.730 360.160 ;
        RECT 235.540 360.070 236.000 360.210 ;
        RECT 233.030 360.010 233.640 360.030 ;
        RECT 235.540 360.010 235.910 360.070 ;
        RECT 236.110 359.910 236.310 360.360 ;
        RECT 237.670 360.290 237.790 360.420 ;
        RECT 237.720 360.220 237.790 360.290 ;
        RECT 341.740 360.260 345.240 360.800 ;
        RECT 236.720 359.950 237.030 360.150 ;
        RECT 237.720 360.010 237.790 360.210 ;
        RECT 239.010 359.950 239.320 360.230 ;
        RECT 223.880 359.710 230.240 359.840 ;
        RECT 234.600 359.710 236.310 359.910 ;
        RECT 236.590 359.730 239.500 359.950 ;
        RECT 223.880 359.590 224.240 359.710 ;
        RECT 221.200 358.940 224.710 359.110 ;
        RECT 220.250 358.930 224.710 358.940 ;
        RECT 227.740 358.930 228.030 359.710 ;
        RECT 228.930 359.370 229.190 359.710 ;
        RECT 233.340 359.440 233.910 359.590 ;
        RECT 233.340 359.390 234.120 359.440 ;
        RECT 228.930 359.230 233.060 359.370 ;
        RECT 233.810 359.240 234.120 359.390 ;
        RECT 234.410 359.320 234.720 359.540 ;
        RECT 234.810 359.320 235.120 359.510 ;
        RECT 236.110 359.320 236.310 359.710 ;
        RECT 234.410 359.240 236.600 359.320 ;
        RECT 233.810 359.230 236.600 359.240 ;
        RECT 228.930 359.160 236.600 359.230 ;
        RECT 236.670 359.170 236.980 359.500 ;
        RECT 237.670 359.470 237.780 359.690 ;
        RECT 232.850 359.100 236.600 359.160 ;
        RECT 166.250 358.390 166.710 358.710 ;
        RECT 168.420 358.350 170.860 358.570 ;
        RECT 158.390 357.800 158.810 357.890 ;
        RECT 158.390 357.630 163.290 357.800 ;
        RECT 158.390 357.540 158.810 357.630 ;
        RECT 163.120 357.450 163.290 357.630 ;
        RECT 168.520 357.550 168.780 358.350 ;
        RECT 169.440 358.320 169.760 358.340 ;
        RECT 169.430 358.270 169.760 358.320 ;
        RECT 170.520 358.290 170.860 358.350 ;
        RECT 170.470 358.270 170.790 358.280 ;
        RECT 172.230 358.270 172.430 358.790 ;
        RECT 178.270 358.580 178.450 358.790 ;
        RECT 220.250 358.730 230.240 358.930 ;
        RECT 230.400 358.880 230.460 359.080 ;
        RECT 232.850 359.030 235.910 359.100 ;
        RECT 236.110 359.060 236.560 359.100 ;
        RECT 232.850 359.020 233.060 359.030 ;
        RECT 233.900 359.020 235.020 359.030 ;
        RECT 232.850 358.810 234.860 359.020 ;
        RECT 235.090 358.880 235.160 359.030 ;
        RECT 220.250 358.720 221.850 358.730 ;
        RECT 169.430 358.070 172.430 358.270 ;
        RECT 173.630 358.500 173.950 358.580 ;
        RECT 176.110 358.550 178.450 358.580 ;
        RECT 176.040 358.500 178.450 358.550 ;
        RECT 224.480 358.520 224.710 358.730 ;
        RECT 227.740 358.670 228.030 358.730 ;
        RECT 227.740 358.520 230.630 358.670 ;
        RECT 236.110 358.660 236.310 359.060 ;
        RECT 240.200 358.660 241.100 359.330 ;
        RECT 173.630 358.420 178.450 358.500 ;
        RECT 173.630 358.310 176.360 358.420 ;
        RECT 176.840 358.410 178.450 358.420 ;
        RECT 177.540 358.400 178.450 358.410 ;
        RECT 207.440 358.360 211.890 358.520 ;
        RECT 207.410 358.340 211.890 358.360 ;
        RECT 212.260 358.450 230.630 358.520 ;
        RECT 212.260 358.420 229.450 358.450 ;
        RECT 232.420 358.440 232.730 358.600 ;
        RECT 212.260 358.340 230.240 358.420 ;
        RECT 206.700 358.320 230.240 358.340 ;
        RECT 173.630 358.260 173.950 358.310 ;
        RECT 176.040 358.290 176.360 358.310 ;
        RECT 169.430 358.060 169.760 358.070 ;
        RECT 169.440 358.050 169.760 358.060 ;
        RECT 170.470 358.020 170.790 358.070 ;
        RECT 173.630 357.640 173.950 357.690 ;
        RECT 176.040 357.640 176.360 357.660 ;
        RECT 173.630 357.620 176.360 357.640 ;
        RECT 178.370 357.640 178.920 357.820 ;
        RECT 202.000 357.780 202.560 358.320 ;
        RECT 206.700 358.120 217.250 358.320 ;
        RECT 224.480 358.170 224.700 358.320 ;
        RECT 229.150 358.220 230.240 358.320 ;
        RECT 230.400 358.220 230.460 358.350 ;
        RECT 231.990 358.220 232.870 358.440 ;
        RECT 233.340 358.410 235.220 358.610 ;
        RECT 234.120 358.280 234.440 358.410 ;
        RECT 228.850 358.210 234.850 358.220 ;
        RECT 228.850 358.200 235.020 358.210 ;
        RECT 235.090 358.200 235.160 358.350 ;
        RECT 235.300 358.200 235.620 358.340 ;
        RECT 236.110 358.230 241.100 358.660 ;
        RECT 228.850 358.170 235.910 358.200 ;
        RECT 206.700 358.080 207.020 358.120 ;
        RECT 206.810 357.740 207.070 357.980 ;
        RECT 178.370 357.620 178.550 357.640 ;
        RECT 173.630 357.460 178.550 357.620 ;
        RECT 206.700 357.630 207.070 357.740 ;
        RECT 206.700 357.480 207.020 357.630 ;
        RECT 173.630 357.450 176.360 357.460 ;
        RECT 163.120 357.280 163.640 357.450 ;
        RECT 173.630 357.370 173.950 357.450 ;
        RECT 176.040 357.400 176.360 357.450 ;
        RECT 163.470 357.130 163.570 357.280 ;
        RECT 172.390 357.150 172.870 357.160 ;
        RECT 166.250 356.640 166.710 356.960 ;
        RECT 172.260 356.860 172.870 357.150 ;
        RECT 168.420 356.600 170.860 356.820 ;
        RECT 157.830 356.230 158.220 356.320 ;
        RECT 157.830 356.060 163.200 356.230 ;
        RECT 157.830 355.970 158.220 356.060 ;
        RECT 163.040 355.950 163.200 356.060 ;
        RECT 163.040 355.650 163.210 355.950 ;
        RECT 168.520 355.800 168.780 356.600 ;
        RECT 169.440 356.570 169.760 356.590 ;
        RECT 169.430 356.520 169.760 356.570 ;
        RECT 170.520 356.540 170.860 356.600 ;
        RECT 172.260 356.710 172.580 356.860 ;
        RECT 207.410 356.780 207.640 358.120 ;
        RECT 224.480 358.010 235.910 358.170 ;
        RECT 224.480 357.950 229.240 358.010 ;
        RECT 233.030 358.000 235.910 358.010 ;
        RECT 236.110 358.060 236.310 358.230 ;
        RECT 233.900 357.990 235.120 358.000 ;
        RECT 224.800 357.650 225.190 357.670 ;
        RECT 209.680 357.450 209.760 357.630 ;
        RECT 224.790 357.540 225.200 357.650 ;
        RECT 232.570 357.580 232.880 357.770 ;
        RECT 234.810 357.720 235.120 357.990 ;
        RECT 236.110 357.980 236.560 358.060 ;
        RECT 236.670 358.010 236.980 358.230 ;
        RECT 235.250 357.800 236.560 357.980 ;
        RECT 235.250 357.630 236.430 357.800 ;
        RECT 238.930 357.790 239.240 357.980 ;
        RECT 224.790 357.440 229.450 357.540 ;
        RECT 224.790 357.340 230.240 357.440 ;
        RECT 224.790 357.300 225.200 357.340 ;
        RECT 229.220 357.300 230.240 357.340 ;
        RECT 230.400 357.300 230.450 357.370 ;
        RECT 232.530 357.330 233.080 357.580 ;
        RECT 235.300 357.540 235.620 357.630 ;
        RECT 236.110 357.540 236.310 357.630 ;
        RECT 236.580 357.560 239.290 357.790 ;
        RECT 234.600 357.450 236.310 357.540 ;
        RECT 234.290 357.300 236.310 357.450 ;
        RECT 236.720 357.360 237.030 357.560 ;
        RECT 218.100 357.240 236.310 357.300 ;
        RECT 240.200 357.240 241.100 358.230 ;
        RECT 243.260 358.210 345.330 360.260 ;
        RECT 218.100 357.150 234.610 357.240 ;
        RECT 235.540 357.160 235.910 357.220 ;
        RECT 218.100 357.000 218.420 357.150 ;
        RECT 223.900 357.000 224.220 357.150 ;
        RECT 233.030 357.090 233.640 357.150 ;
        RECT 233.030 357.020 233.730 357.090 ;
        RECT 235.540 357.020 236.000 357.160 ;
        RECT 225.620 356.950 226.020 356.960 ;
        RECT 209.920 356.800 210.240 356.920 ;
        RECT 225.600 356.890 226.040 356.950 ;
        RECT 233.410 356.940 233.730 357.020 ;
        RECT 225.600 356.800 229.450 356.890 ;
        RECT 231.730 356.800 232.040 356.930 ;
        RECT 232.120 356.800 232.440 356.920 ;
        RECT 170.470 356.520 170.790 356.530 ;
        RECT 172.260 356.520 172.460 356.710 ;
        RECT 207.410 356.560 207.910 356.780 ;
        RECT 209.920 356.620 232.440 356.800 ;
        RECT 233.240 356.830 233.730 356.940 ;
        RECT 235.680 356.900 236.000 357.020 ;
        RECT 236.110 356.890 236.310 357.240 ;
        RECT 236.710 356.890 237.020 357.120 ;
        RECT 237.720 357.020 237.790 357.220 ;
        RECT 238.960 356.890 239.270 357.140 ;
        RECT 233.240 356.700 233.550 356.830 ;
        RECT 234.600 356.780 236.310 356.890 ;
        RECT 169.430 356.320 172.460 356.520 ;
        RECT 205.720 356.350 217.250 356.560 ;
        RECT 229.100 356.510 230.240 356.620 ;
        RECT 231.730 356.600 232.040 356.620 ;
        RECT 234.410 356.570 236.310 356.780 ;
        RECT 236.580 356.810 239.270 356.890 ;
        RECT 236.580 356.660 239.120 356.810 ;
        RECT 234.410 356.560 236.300 356.570 ;
        RECT 207.030 356.340 217.250 356.350 ;
        RECT 169.430 356.310 169.760 356.320 ;
        RECT 169.440 356.300 169.760 356.310 ;
        RECT 170.470 356.270 170.790 356.320 ;
        RECT 172.530 355.820 172.870 355.890 ;
        RECT 207.410 355.840 207.640 356.340 ;
        RECT 209.680 356.290 209.750 356.340 ;
        RECT 232.710 356.300 233.180 356.550 ;
        RECT 234.410 356.450 236.600 356.560 ;
        RECT 214.890 355.930 215.200 356.260 ;
        RECT 232.850 356.210 233.170 356.300 ;
        RECT 233.340 356.240 233.910 356.390 ;
        RECT 234.560 356.350 236.600 356.450 ;
        RECT 233.340 356.190 234.120 356.240 ;
        RECT 215.300 355.910 217.250 356.030 ;
        RECT 233.810 355.910 234.120 356.190 ;
        RECT 234.350 356.070 234.570 356.090 ;
        RECT 172.390 355.770 172.870 355.820 ;
        RECT 163.470 355.650 163.570 355.700 ;
        RECT 163.040 355.480 163.640 355.650 ;
        RECT 172.190 355.590 172.870 355.770 ;
        RECT 163.470 355.380 163.570 355.480 ;
        RECT 166.250 354.890 166.710 355.210 ;
        RECT 168.420 354.850 170.860 355.070 ;
        RECT 168.520 354.050 168.780 354.850 ;
        RECT 169.440 354.820 169.760 354.840 ;
        RECT 169.430 354.770 169.760 354.820 ;
        RECT 170.520 354.790 170.860 354.850 ;
        RECT 170.470 354.770 170.790 354.780 ;
        RECT 172.190 354.770 172.370 355.590 ;
        RECT 173.630 355.300 173.950 355.380 ;
        RECT 176.040 355.320 176.360 355.350 ;
        RECT 176.040 355.300 178.650 355.320 ;
        RECT 173.630 355.140 178.650 355.300 ;
        RECT 203.040 355.230 203.660 355.760 ;
        RECT 206.660 355.610 207.640 355.840 ;
        RECT 208.250 355.710 211.890 355.910 ;
        RECT 212.260 355.730 229.450 355.910 ;
        RECT 232.230 355.750 232.660 355.760 ;
        RECT 212.260 355.710 230.240 355.730 ;
        RECT 208.030 355.460 208.190 355.480 ;
        RECT 208.250 355.460 208.450 355.710 ;
        RECT 218.580 355.690 219.420 355.710 ;
        RECT 229.190 355.530 230.240 355.710 ;
        RECT 232.230 355.520 233.100 355.750 ;
        RECT 234.300 355.730 234.570 356.070 ;
        RECT 236.220 356.030 236.550 356.240 ;
        RECT 236.660 356.140 236.970 356.470 ;
        RECT 353.440 356.190 359.150 361.830 ;
        RECT 353.000 356.150 359.150 356.190 ;
        RECT 243.260 355.690 359.150 356.150 ;
        RECT 232.460 355.460 232.770 355.520 ;
        RECT 234.130 355.460 234.290 355.480 ;
        RECT 208.030 355.410 217.250 355.460 ;
        RECT 225.070 355.440 234.290 355.460 ;
        RECT 208.150 355.310 217.250 355.410 ;
        RECT 219.030 355.410 234.290 355.440 ;
        RECT 219.030 355.310 235.220 355.410 ;
        RECT 173.630 355.110 176.360 355.140 ;
        RECT 173.630 355.060 173.950 355.110 ;
        RECT 176.040 355.090 176.360 355.110 ;
        RECT 169.430 354.570 172.380 354.770 ;
        RECT 169.430 354.560 169.760 354.570 ;
        RECT 169.440 354.550 169.760 354.560 ;
        RECT 170.470 354.520 170.790 354.570 ;
        RECT 178.470 352.950 178.650 355.140 ;
        RECT 203.130 355.050 203.440 355.190 ;
        RECT 200.960 354.870 203.440 355.050 ;
        RECT 208.250 355.010 208.450 355.310 ;
        RECT 219.030 355.220 229.170 355.310 ;
        RECT 232.560 355.230 232.910 355.310 ;
        RECT 203.130 354.860 203.440 354.870 ;
        RECT 206.670 354.860 208.450 355.010 ;
        RECT 206.670 354.790 208.420 354.860 ;
        RECT 218.980 354.250 227.990 354.470 ;
        RECT 218.160 353.810 218.480 353.860 ;
        RECT 218.160 353.560 224.180 353.810 ;
        RECT 223.860 353.490 224.180 353.560 ;
        RECT 178.470 352.770 179.010 352.950 ;
        RECT 219.030 352.470 224.690 352.690 ;
        RECT 218.530 352.170 219.010 352.180 ;
        RECT 181.610 352.010 181.930 352.020 ;
        RECT 209.420 352.010 209.880 352.080 ;
        RECT 181.610 351.730 209.880 352.010 ;
        RECT 218.530 351.930 219.420 352.170 ;
        RECT 224.470 352.140 224.690 352.470 ;
        RECT 227.770 352.640 227.990 354.250 ;
        RECT 228.950 354.020 229.170 355.220 ;
        RECT 233.340 355.210 235.220 355.310 ;
        RECT 236.220 355.210 236.550 355.420 ;
        RECT 234.120 355.170 234.440 355.210 ;
        RECT 234.120 355.160 234.570 355.170 ;
        RECT 234.120 355.080 234.590 355.160 ;
        RECT 234.370 354.830 234.590 355.080 ;
        RECT 236.660 354.980 236.970 355.310 ;
        RECT 238.880 355.050 239.190 355.190 ;
        RECT 238.880 354.870 241.360 355.050 ;
        RECT 238.880 354.860 239.320 354.870 ;
        RECT 234.390 354.820 234.590 354.830 ;
        RECT 239.010 354.750 239.320 354.860 ;
        RECT 236.840 354.660 239.490 354.750 ;
        RECT 236.710 354.520 239.490 354.660 ;
        RECT 236.710 354.330 237.020 354.520 ;
        RECT 233.320 354.030 233.640 354.270 ;
        RECT 237.660 354.260 237.770 354.490 ;
        RECT 228.920 353.980 229.170 354.020 ;
        RECT 228.920 353.340 229.180 353.980 ;
        RECT 236.710 353.920 237.020 354.120 ;
        RECT 239.000 353.920 239.310 354.200 ;
        RECT 236.580 353.700 239.490 353.920 ;
        RECT 243.260 353.790 358.990 355.690 ;
        RECT 228.920 353.130 233.050 353.340 ;
        RECT 232.840 352.990 233.050 353.130 ;
        RECT 236.220 353.030 236.550 353.240 ;
        RECT 236.660 353.140 236.970 353.470 ;
        RECT 237.660 353.440 237.770 353.660 ;
        RECT 232.840 352.780 234.860 352.990 ;
        RECT 227.770 352.420 230.620 352.640 ;
        RECT 232.410 352.410 232.720 352.570 ;
        RECT 231.980 352.190 232.860 352.410 ;
        RECT 236.220 352.210 236.550 352.420 ;
        RECT 228.840 352.140 234.860 352.190 ;
        RECT 224.470 351.980 234.860 352.140 ;
        RECT 236.660 351.980 236.970 352.310 ;
        RECT 224.470 351.920 229.230 351.980 ;
        RECT 238.920 351.760 239.230 351.950 ;
        RECT 181.610 351.680 181.930 351.730 ;
        RECT 209.420 351.670 209.880 351.730 ;
        RECT 209.680 351.420 209.760 351.600 ;
        RECT 232.560 351.550 232.870 351.740 ;
        RECT 210.210 351.410 210.640 351.490 ;
        RECT 198.950 351.150 210.640 351.410 ;
        RECT 232.520 351.300 233.070 351.550 ;
        RECT 236.570 351.530 239.280 351.760 ;
        RECT 198.950 351.140 199.270 351.150 ;
        RECT 210.210 351.080 210.640 351.150 ;
        RECT 223.860 351.270 224.180 351.280 ;
        RECT 234.300 351.270 234.630 351.410 ;
        RECT 236.710 351.330 237.020 351.530 ;
        RECT 347.660 351.410 349.750 351.590 ;
        RECT 223.860 351.110 234.630 351.270 ;
        RECT 223.860 351.100 224.550 351.110 ;
        RECT 223.860 350.980 224.180 351.100 ;
        RECT 157.220 350.760 157.590 350.880 ;
        RECT 163.470 350.760 163.570 350.820 ;
        RECT 157.220 350.590 163.570 350.760 ;
        RECT 157.220 350.480 157.590 350.590 ;
        RECT 163.470 350.500 163.570 350.590 ;
        RECT 231.720 350.570 232.030 350.900 ;
        RECT 173.610 350.370 173.930 350.420 ;
        RECT 176.020 350.370 176.340 350.390 ;
        RECT 173.610 350.350 178.090 350.370 ;
        RECT 178.390 350.350 178.570 350.360 ;
        RECT 166.250 350.010 166.710 350.330 ;
        RECT 173.610 350.240 178.570 350.350 ;
        RECT 198.860 350.320 214.100 350.500 ;
        RECT 232.700 350.270 233.170 350.520 ;
        RECT 173.610 350.200 180.400 350.240 ;
        RECT 168.420 349.970 170.860 350.190 ;
        RECT 173.610 350.180 176.340 350.200 ;
        RECT 173.610 350.100 173.930 350.180 ;
        RECT 176.020 350.130 176.340 350.180 ;
        RECT 178.050 350.170 180.400 350.200 ;
        RECT 178.390 350.060 180.400 350.170 ;
        RECT 198.440 350.070 198.750 350.240 ;
        RECT 232.840 350.180 233.160 350.270 ;
        RECT 156.580 349.170 156.970 349.260 ;
        RECT 168.520 349.170 168.780 349.970 ;
        RECT 169.440 349.940 169.760 349.960 ;
        RECT 169.430 349.890 169.760 349.940 ;
        RECT 170.520 349.910 170.860 349.970 ;
        RECT 196.420 349.910 198.750 350.070 ;
        RECT 198.890 350.060 198.980 350.070 ;
        RECT 213.980 350.060 214.070 350.070 ;
        RECT 170.470 349.890 170.790 349.900 ;
        RECT 196.420 349.890 198.590 349.910 ;
        RECT 169.430 349.690 172.850 349.890 ;
        RECT 198.860 349.880 214.100 350.060 ;
        RECT 169.430 349.680 169.760 349.690 ;
        RECT 169.440 349.670 169.760 349.680 ;
        RECT 170.470 349.640 170.790 349.690 ;
        RECT 172.370 349.660 172.850 349.690 ;
        RECT 172.510 349.590 172.850 349.660 ;
        RECT 232.220 349.720 232.650 349.730 ;
        RECT 232.220 349.490 233.090 349.720 ;
        RECT 232.450 349.290 232.760 349.490 ;
        RECT 243.260 349.320 349.750 351.410 ;
        RECT 156.580 349.070 163.540 349.170 ;
        RECT 156.580 349.050 163.570 349.070 ;
        RECT 156.580 349.000 163.640 349.050 ;
        RECT 210.950 349.040 211.390 349.160 ;
        RECT 156.580 348.910 156.970 349.000 ;
        RECT 163.250 348.880 163.640 349.000 ;
        RECT 210.820 348.960 211.390 349.040 ;
        RECT 196.420 348.940 198.590 348.960 ;
        RECT 163.470 348.750 163.570 348.880 ;
        RECT 196.420 348.780 198.750 348.940 ;
        RECT 198.860 348.780 214.100 348.960 ;
        RECT 166.250 348.260 166.710 348.580 ;
        RECT 172.510 348.550 172.850 348.620 ;
        RECT 198.440 348.610 198.750 348.780 ;
        RECT 210.940 348.760 211.390 348.780 ;
        RECT 210.940 348.700 211.340 348.760 ;
        RECT 172.370 348.500 172.850 348.550 ;
        RECT 200.110 348.530 211.340 348.700 ;
        RECT 172.170 348.490 172.850 348.500 ;
        RECT 168.420 348.220 170.860 348.440 ;
        RECT 125.500 347.590 136.800 347.960 ;
        RECT 155.960 347.620 156.350 347.700 ;
        RECT 125.500 346.990 126.770 347.590 ;
        RECT 155.960 347.450 163.140 347.620 ;
        RECT 155.960 347.370 156.350 347.450 ;
        RECT 162.990 347.380 163.140 347.450 ;
        RECT 168.520 347.420 168.780 348.220 ;
        RECT 169.440 348.190 169.760 348.210 ;
        RECT 169.430 348.140 169.760 348.190 ;
        RECT 170.520 348.160 170.860 348.220 ;
        RECT 172.150 348.320 172.850 348.490 ;
        RECT 196.420 348.390 198.600 348.530 ;
        RECT 196.420 348.350 198.750 348.390 ;
        RECT 198.860 348.350 214.100 348.530 ;
        RECT 170.470 348.140 170.790 348.150 ;
        RECT 172.150 348.140 172.350 348.320 ;
        RECT 169.430 347.940 172.350 348.140 ;
        RECT 178.130 348.110 180.460 348.270 ;
        RECT 173.610 348.030 173.930 348.110 ;
        RECT 176.090 348.090 180.460 348.110 ;
        RECT 176.090 348.080 178.310 348.090 ;
        RECT 176.020 348.030 178.310 348.080 ;
        RECT 198.440 348.060 198.750 348.350 ;
        RECT 173.610 347.950 178.310 348.030 ;
        RECT 169.430 347.930 169.760 347.940 ;
        RECT 169.440 347.920 169.760 347.930 ;
        RECT 170.470 347.890 170.790 347.940 ;
        RECT 173.610 347.840 176.340 347.950 ;
        RECT 176.820 347.940 178.310 347.950 ;
        RECT 177.520 347.930 178.310 347.940 ;
        RECT 173.610 347.790 173.930 347.840 ;
        RECT 176.020 347.820 176.340 347.840 ;
        RECT 162.990 347.270 163.160 347.380 ;
        RECT 163.470 347.270 163.570 347.320 ;
        RECT 162.990 347.100 163.640 347.270 ;
        RECT 198.440 347.260 198.750 347.550 ;
        RECT 196.420 347.220 198.750 347.260 ;
        RECT 173.610 347.170 173.930 347.220 ;
        RECT 176.020 347.170 176.340 347.190 ;
        RECT 173.610 347.150 176.340 347.170 ;
        RECT 173.610 347.140 178.330 347.150 ;
        RECT 163.470 347.000 163.570 347.100 ;
        RECT 173.610 347.000 178.340 347.140 ;
        RECT 196.420 347.080 198.600 347.220 ;
        RECT 198.870 347.080 214.090 347.260 ;
        RECT 173.610 346.990 180.440 347.000 ;
        RECT 173.610 346.980 176.340 346.990 ;
        RECT 173.610 346.900 173.930 346.980 ;
        RECT 176.020 346.930 176.340 346.980 ;
        RECT 166.250 346.510 166.710 346.830 ;
        RECT 178.160 346.820 180.440 346.990 ;
        RECT 198.440 346.830 198.750 347.000 ;
        RECT 168.420 346.470 170.860 346.690 ;
        RECT 172.370 346.670 172.850 346.690 ;
        RECT 155.350 346.140 155.770 346.230 ;
        RECT 155.350 345.970 163.160 346.140 ;
        RECT 155.350 345.870 155.770 345.970 ;
        RECT 27.670 301.280 29.970 304.690 ;
        RECT 27.890 300.950 29.970 301.280 ;
        RECT 32.230 343.810 127.730 345.780 ;
        RECT 162.990 345.480 163.160 345.970 ;
        RECT 168.520 345.670 168.780 346.470 ;
        RECT 169.440 346.440 169.760 346.460 ;
        RECT 169.430 346.390 169.760 346.440 ;
        RECT 170.520 346.410 170.860 346.470 ;
        RECT 170.470 346.390 170.790 346.400 ;
        RECT 172.100 346.390 172.850 346.670 ;
        RECT 196.420 346.670 198.750 346.830 ;
        RECT 196.420 346.650 198.590 346.670 ;
        RECT 198.860 346.650 214.100 346.830 ;
        RECT 169.430 346.340 172.590 346.390 ;
        RECT 169.430 346.190 172.450 346.340 ;
        RECT 169.430 346.180 169.760 346.190 ;
        RECT 169.440 346.170 169.760 346.180 ;
        RECT 170.470 346.140 170.790 346.190 ;
        RECT 196.400 345.730 196.710 345.810 ;
        RECT 196.400 345.710 198.590 345.730 ;
        RECT 163.470 345.480 163.570 345.570 ;
        RECT 196.400 345.550 198.750 345.710 ;
        RECT 198.870 345.550 214.090 345.730 ;
        RECT 196.400 345.520 196.710 345.550 ;
        RECT 194.380 345.480 196.710 345.520 ;
        RECT 162.990 345.310 163.640 345.480 ;
        RECT 172.510 345.350 172.850 345.420 ;
        RECT 163.470 345.250 163.570 345.310 ;
        RECT 172.140 345.120 172.850 345.350 ;
        RECT 194.380 345.340 196.560 345.480 ;
        RECT 198.440 345.380 198.750 345.550 ;
        RECT 196.420 345.260 198.600 345.300 ;
        RECT 196.400 345.160 198.600 345.260 ;
        RECT 196.400 345.120 198.750 345.160 ;
        RECT 198.890 345.130 214.070 345.300 ;
        RECT 166.250 344.760 166.710 345.080 ;
        RECT 168.420 344.720 170.860 344.940 ;
        RECT 168.520 343.920 168.780 344.720 ;
        RECT 169.440 344.690 169.760 344.710 ;
        RECT 169.430 344.640 169.760 344.690 ;
        RECT 170.520 344.660 170.860 344.720 ;
        RECT 170.470 344.640 170.790 344.650 ;
        RECT 172.140 344.640 172.340 345.120 ;
        RECT 196.400 345.090 196.710 345.120 ;
        RECT 198.440 345.090 198.750 345.120 ;
        RECT 169.430 344.440 172.340 344.640 ;
        RECT 173.610 344.830 173.930 344.910 ;
        RECT 176.020 344.850 176.340 344.880 ;
        RECT 178.120 344.860 180.420 345.040 ;
        RECT 194.380 344.930 196.710 345.090 ;
        RECT 194.380 344.910 196.550 344.930 ;
        RECT 196.840 344.900 204.450 345.090 ;
        RECT 178.120 344.850 178.320 344.860 ;
        RECT 176.020 344.830 178.320 344.850 ;
        RECT 198.440 344.830 198.750 344.900 ;
        RECT 173.610 344.670 178.320 344.830 ;
        RECT 173.610 344.640 176.340 344.670 ;
        RECT 173.610 344.590 173.930 344.640 ;
        RECT 176.020 344.620 176.340 344.640 ;
        RECT 169.430 344.430 169.760 344.440 ;
        RECT 169.440 344.420 169.760 344.430 ;
        RECT 170.470 344.390 170.790 344.440 ;
        RECT 194.380 343.980 196.550 344.000 ;
        RECT 174.230 343.930 174.540 343.950 ;
        RECT 194.380 343.930 196.710 343.980 ;
        RECT 196.820 343.930 204.450 344.000 ;
        RECT 211.870 343.930 212.320 343.960 ;
        RECT 32.230 343.700 135.140 343.810 ;
        RECT 32.230 276.210 34.310 343.700 ;
        RECT 125.440 343.440 135.140 343.700 ;
        RECT 174.230 343.520 212.320 343.930 ;
        RECT 243.260 343.920 345.610 346.010 ;
        RECT 174.230 343.500 174.540 343.520 ;
        RECT 125.440 342.770 126.710 343.440 ;
        RECT 134.770 342.090 135.140 343.440 ;
        RECT 194.380 343.430 196.560 343.520 ;
        RECT 211.870 343.500 212.320 343.520 ;
        RECT 194.380 343.390 196.710 343.430 ;
        RECT 196.400 343.100 196.710 343.390 ;
        RECT 196.850 343.380 196.940 343.410 ;
        RECT 196.820 343.270 196.940 343.380 ;
        RECT 196.820 342.120 196.970 342.290 ;
        RECT 134.770 342.080 136.800 342.090 ;
        RECT 134.770 341.900 137.020 342.080 ;
        RECT 134.770 341.840 138.420 341.900 ;
        RECT 196.400 341.850 196.710 342.020 ;
        RECT 134.770 341.720 139.750 341.840 ;
        RECT 145.070 341.830 145.370 341.850 ;
        RECT 145.060 341.810 145.380 341.830 ;
        RECT 136.430 341.680 139.750 341.720 ;
        RECT 136.800 341.620 139.750 341.680 ;
        RECT 129.430 341.430 130.200 341.620 ;
        RECT 142.840 341.590 145.380 341.810 ;
        RECT 163.430 341.680 163.530 341.760 ;
        RECT 194.380 341.690 196.710 341.850 ;
        RECT 136.430 341.430 136.820 341.450 ;
        RECT 129.430 341.390 136.820 341.430 ;
        RECT 129.430 341.180 139.740 341.390 ;
        RECT 36.770 339.780 127.730 341.080 ;
        RECT 129.430 341.060 136.810 341.180 ;
        RECT 142.840 341.150 143.060 341.590 ;
        RECT 145.060 341.570 145.380 341.590 ;
        RECT 145.070 341.550 145.370 341.570 ;
        RECT 163.180 341.510 163.600 341.680 ;
        RECT 194.380 341.670 196.550 341.690 ;
        RECT 196.820 341.680 203.680 341.850 ;
        RECT 203.980 341.710 204.450 341.870 ;
        RECT 203.980 341.700 204.440 341.710 ;
        RECT 196.850 341.670 196.940 341.680 ;
        RECT 163.180 341.410 163.560 341.510 ;
        RECT 163.180 341.190 163.460 341.410 ;
        RECT 196.470 341.340 197.200 341.520 ;
        RECT 129.430 340.880 130.200 341.060 ;
        RECT 136.430 341.040 136.800 341.060 ;
        RECT 154.710 340.970 155.120 341.070 ;
        RECT 163.180 340.970 163.450 341.190 ;
        RECT 154.710 340.800 163.450 340.970 ;
        RECT 166.210 340.950 166.670 341.270 ;
        RECT 168.380 340.910 170.820 341.130 ;
        RECT 154.710 340.710 155.120 340.800 ;
        RECT 163.180 340.790 163.350 340.800 ;
        RECT 146.170 340.300 146.860 340.380 ;
        RECT 145.360 339.970 145.670 340.300 ;
        RECT 146.010 340.170 146.860 340.300 ;
        RECT 146.010 339.970 146.320 340.170 ;
        RECT 168.480 340.110 168.740 340.910 ;
        RECT 169.400 340.880 169.720 340.900 ;
        RECT 169.390 340.830 169.720 340.880 ;
        RECT 170.480 340.850 170.820 340.910 ;
        RECT 173.640 341.100 173.960 341.150 ;
        RECT 176.050 341.100 176.370 341.120 ;
        RECT 173.640 341.090 178.120 341.100 ;
        RECT 206.980 341.090 207.120 341.100 ;
        RECT 173.640 340.930 178.250 341.090 ;
        RECT 173.640 340.910 176.370 340.930 ;
        RECT 177.940 340.910 178.250 340.930 ;
        RECT 170.430 340.830 170.750 340.840 ;
        RECT 173.640 340.830 173.960 340.910 ;
        RECT 176.050 340.860 176.370 340.910 ;
        RECT 169.390 340.630 172.470 340.830 ;
        RECT 178.070 340.730 180.420 340.910 ;
        RECT 196.820 340.720 204.450 340.890 ;
        RECT 206.980 340.760 207.130 341.090 ;
        RECT 208.000 340.870 208.310 341.200 ;
        RECT 169.390 340.620 169.720 340.630 ;
        RECT 169.400 340.610 169.720 340.620 ;
        RECT 170.430 340.580 170.750 340.630 ;
        RECT 172.270 340.620 172.470 340.630 ;
        RECT 172.270 340.390 172.880 340.620 ;
        RECT 196.850 340.570 196.940 340.720 ;
        RECT 206.980 340.560 208.190 340.760 ;
        RECT 208.300 340.520 210.590 340.610 ;
        RECT 172.540 340.320 172.880 340.390 ;
        RECT 208.150 340.450 210.590 340.520 ;
        RECT 178.710 340.100 179.880 340.250 ;
        RECT 208.150 340.190 208.460 340.450 ;
        RECT 36.770 339.410 131.490 339.780 ;
        RECT 143.330 339.750 144.040 339.960 ;
        RECT 144.990 339.860 146.860 339.940 ;
        RECT 163.430 339.920 163.530 340.010 ;
        RECT 144.840 339.720 146.860 339.860 ;
        RECT 163.120 339.750 163.600 339.920 ;
        RECT 178.650 339.770 178.930 340.100 ;
        RECT 207.090 339.940 208.290 340.000 ;
        RECT 207.090 339.900 208.460 339.940 ;
        RECT 207.080 339.820 208.460 339.900 ;
        RECT 144.840 339.530 145.150 339.720 ;
        RECT 36.770 339.000 127.730 339.410 ;
        RECT 32.020 272.610 34.590 276.210 ;
        RECT 32.230 272.570 34.310 272.610 ;
        RECT 36.770 247.590 38.850 339.000 ;
        RECT 125.500 338.670 126.770 339.000 ;
        RECT 131.120 337.750 131.490 339.410 ;
        RECT 154.050 339.400 154.440 339.510 ;
        RECT 163.120 339.460 163.290 339.750 ;
        RECT 163.430 339.690 163.530 339.750 ;
        RECT 208.010 339.700 208.460 339.820 ;
        RECT 208.010 339.680 208.040 339.700 ;
        RECT 208.150 339.680 208.460 339.700 ;
        RECT 208.150 339.610 210.590 339.680 ;
        RECT 163.120 339.400 163.280 339.460 ;
        RECT 146.380 339.220 146.700 339.280 ;
        RECT 154.050 339.240 163.280 339.400 ;
        RECT 154.050 339.230 162.930 339.240 ;
        RECT 146.380 339.010 146.860 339.220 ;
        RECT 154.050 339.130 154.440 339.230 ;
        RECT 166.210 339.200 166.670 339.520 ;
        RECT 196.440 339.390 197.020 339.570 ;
        RECT 208.300 339.520 210.590 339.610 ;
        RECT 168.380 339.160 170.820 339.380 ;
        RECT 172.540 339.280 172.880 339.350 ;
        RECT 172.400 339.240 172.880 339.280 ;
        RECT 146.380 338.960 146.700 339.010 ;
        RECT 143.330 338.390 143.580 338.610 ;
        RECT 168.480 338.360 168.740 339.160 ;
        RECT 169.400 339.130 169.720 339.150 ;
        RECT 169.390 339.080 169.720 339.130 ;
        RECT 170.480 339.100 170.820 339.160 ;
        RECT 170.430 339.080 170.750 339.090 ;
        RECT 172.260 339.080 172.880 339.240 ;
        RECT 169.390 339.050 172.880 339.080 ;
        RECT 169.390 338.880 172.580 339.050 ;
        RECT 169.390 338.870 169.720 338.880 ;
        RECT 169.400 338.860 169.720 338.870 ;
        RECT 170.430 338.830 170.750 338.880 ;
        RECT 178.050 338.840 179.840 338.960 ;
        RECT 208.000 338.930 208.310 339.260 ;
        RECT 243.260 339.040 341.530 341.130 ;
        RECT 173.640 338.760 173.960 338.840 ;
        RECT 176.120 338.810 179.840 338.840 ;
        RECT 176.050 338.780 179.840 338.810 ;
        RECT 176.050 338.760 178.230 338.780 ;
        RECT 173.640 338.680 178.230 338.760 ;
        RECT 173.640 338.570 176.370 338.680 ;
        RECT 176.850 338.670 178.230 338.680 ;
        RECT 177.550 338.660 178.230 338.670 ;
        RECT 173.640 338.520 173.960 338.570 ;
        RECT 176.050 338.550 176.370 338.570 ;
        RECT 177.910 338.630 178.230 338.660 ;
        RECT 177.910 338.550 178.090 338.630 ;
        RECT 163.430 338.110 163.530 338.260 ;
        RECT 163.040 337.940 163.600 338.110 ;
        RECT 196.470 338.100 197.020 338.280 ;
        RECT 208.000 338.100 208.310 338.430 ;
        RECT 163.040 337.900 163.210 337.940 ;
        RECT 173.640 337.900 173.960 337.950 ;
        RECT 176.050 337.900 176.370 337.920 ;
        RECT 153.440 337.860 153.810 337.870 ;
        RECT 163.040 337.860 163.200 337.900 ;
        RECT 131.120 337.570 137.070 337.750 ;
        RECT 153.440 337.690 163.200 337.860 ;
        RECT 173.640 337.880 176.370 337.900 ;
        RECT 131.120 337.500 137.140 337.570 ;
        RECT 138.530 337.500 139.750 337.510 ;
        RECT 131.120 337.380 139.750 337.500 ;
        RECT 153.440 337.480 153.810 337.690 ;
        RECT 166.210 337.450 166.670 337.770 ;
        RECT 173.640 337.720 178.160 337.880 ;
        RECT 173.640 337.710 176.370 337.720 ;
        RECT 173.640 337.630 173.960 337.710 ;
        RECT 176.050 337.660 176.370 337.710 ;
        RECT 177.980 337.670 178.160 337.720 ;
        RECT 207.070 337.710 208.070 337.870 ;
        RECT 208.300 337.750 210.590 337.840 ;
        RECT 208.150 337.680 210.590 337.750 ;
        RECT 168.380 337.410 170.820 337.630 ;
        RECT 177.980 337.490 179.870 337.670 ;
        RECT 208.150 337.420 208.460 337.680 ;
        RECT 136.430 337.340 139.750 337.380 ;
        RECT 136.790 337.290 139.750 337.340 ;
        RECT 143.330 336.850 143.580 337.070 ;
        RECT 41.120 335.640 127.730 336.820 ;
        RECT 146.360 336.610 146.680 336.660 ;
        RECT 168.480 336.610 168.740 337.410 ;
        RECT 169.400 337.380 169.720 337.400 ;
        RECT 169.390 337.330 169.720 337.380 ;
        RECT 170.480 337.350 170.820 337.410 ;
        RECT 170.430 337.330 170.750 337.340 ;
        RECT 172.400 337.330 172.880 337.420 ;
        RECT 210.140 337.350 210.470 337.440 ;
        RECT 169.390 337.130 172.880 337.330 ;
        RECT 169.390 337.120 169.720 337.130 ;
        RECT 169.400 337.110 169.720 337.120 ;
        RECT 170.430 337.080 170.750 337.130 ;
        RECT 172.340 337.120 172.880 337.130 ;
        RECT 179.260 337.260 179.580 337.300 ;
        RECT 172.340 337.040 172.630 337.120 ;
        RECT 179.260 337.050 179.870 337.260 ;
        RECT 203.790 337.180 210.470 337.350 ;
        RECT 179.260 336.980 179.720 337.050 ;
        RECT 208.150 336.910 208.460 337.170 ;
        RECT 210.140 337.150 210.470 337.180 ;
        RECT 207.080 336.730 208.080 336.900 ;
        RECT 208.150 336.840 210.590 336.910 ;
        RECT 208.300 336.750 210.590 336.840 ;
        RECT 207.080 336.720 208.020 336.730 ;
        RECT 146.360 336.400 146.860 336.610 ;
        RECT 146.360 336.340 146.680 336.400 ;
        RECT 152.750 336.320 153.140 336.420 ;
        RECT 163.430 336.390 163.530 336.510 ;
        RECT 162.950 336.320 163.600 336.390 ;
        RECT 152.750 336.220 163.600 336.320 ;
        RECT 152.750 336.150 163.240 336.220 ;
        RECT 163.430 336.190 163.530 336.220 ;
        RECT 172.320 336.160 172.620 336.200 ;
        RECT 208.000 336.160 208.310 336.490 ;
        RECT 143.330 336.070 143.600 336.080 ;
        RECT 129.430 335.640 130.230 335.780 ;
        RECT 142.080 335.750 142.680 335.900 ;
        RECT 143.330 335.860 144.080 336.070 ;
        RECT 152.750 336.050 153.140 336.150 ;
        RECT 163.070 336.130 163.240 336.150 ;
        RECT 172.310 336.150 172.620 336.160 ;
        RECT 145.030 335.970 146.860 336.050 ;
        RECT 41.120 335.140 130.230 335.640 ;
        RECT 141.930 335.420 142.680 335.750 ;
        RECT 144.860 335.840 146.860 335.970 ;
        RECT 144.860 335.640 145.170 335.840 ;
        RECT 166.210 335.700 166.670 336.020 ;
        RECT 168.380 335.660 170.820 335.880 ;
        RECT 142.080 335.280 142.680 335.420 ;
        RECT 41.120 334.740 127.730 335.140 ;
        RECT 129.430 335.010 130.230 335.140 ;
        RECT 141.940 335.080 142.680 335.280 ;
        RECT 143.330 335.080 145.290 335.300 ;
        RECT 141.940 334.950 142.250 335.080 ;
        RECT 145.340 334.870 145.650 335.200 ;
        RECT 146.180 335.140 146.860 335.220 ;
        RECT 146.050 335.010 146.860 335.140 ;
        RECT 146.050 334.810 146.360 335.010 ;
        RECT 168.480 334.860 168.740 335.660 ;
        RECT 169.400 335.630 169.720 335.650 ;
        RECT 169.390 335.580 169.720 335.630 ;
        RECT 170.480 335.600 170.820 335.660 ;
        RECT 172.310 335.850 172.880 336.150 ;
        RECT 170.430 335.580 170.750 335.590 ;
        RECT 172.310 335.580 172.510 335.850 ;
        RECT 169.390 335.380 172.510 335.580 ;
        RECT 173.640 335.560 173.960 335.640 ;
        RECT 176.050 335.580 176.370 335.610 ;
        RECT 178.220 335.580 179.850 335.710 ;
        RECT 176.050 335.560 179.850 335.580 ;
        RECT 173.640 335.530 179.850 335.560 ;
        RECT 173.640 335.400 178.400 335.530 ;
        RECT 169.390 335.370 169.720 335.380 ;
        RECT 169.400 335.360 169.720 335.370 ;
        RECT 170.430 335.330 170.750 335.380 ;
        RECT 173.640 335.370 176.370 335.400 ;
        RECT 173.640 335.320 173.960 335.370 ;
        RECT 176.050 335.350 176.370 335.370 ;
        RECT 172.050 334.880 172.370 334.930 ;
        RECT 178.660 334.880 178.980 334.980 ;
        RECT 36.610 244.020 39.000 247.590 ;
        RECT 36.770 243.490 38.850 244.020 ;
        RECT 41.120 218.980 43.200 334.740 ;
        RECT 125.500 334.580 126.770 334.740 ;
        RECT 172.050 334.720 178.980 334.880 ;
        RECT 172.050 334.670 172.370 334.720 ;
        RECT 178.660 334.700 178.980 334.720 ;
        RECT 179.690 334.860 180.010 335.170 ;
        RECT 190.310 334.880 190.720 334.990 ;
        RECT 183.340 334.860 190.720 334.880 ;
        RECT 179.690 334.720 190.720 334.860 ;
        RECT 179.690 334.690 180.010 334.720 ;
        RECT 183.260 334.650 190.720 334.720 ;
        RECT 179.250 334.640 179.530 334.650 ;
        RECT 179.230 334.550 179.550 334.640 ;
        RECT 190.310 334.620 190.720 334.650 ;
        RECT 181.470 334.550 181.790 334.580 ;
        RECT 179.200 334.390 181.790 334.550 ;
        RECT 179.230 334.380 179.550 334.390 ;
        RECT 179.250 334.370 179.530 334.380 ;
        RECT 181.470 334.320 181.790 334.390 ;
        RECT 181.490 334.310 181.770 334.320 ;
        RECT 243.260 333.840 337.440 335.930 ;
        RECT 172.490 333.400 172.800 333.540 ;
        RECT 173.580 333.400 173.890 333.540 ;
        RECT 174.680 333.400 174.990 333.530 ;
        RECT 171.810 333.390 174.990 333.400 ;
        RECT 171.720 333.200 174.990 333.390 ;
        RECT 177.250 333.400 177.560 333.530 ;
        RECT 178.350 333.400 178.660 333.540 ;
        RECT 179.440 333.400 179.750 333.540 ;
        RECT 182.300 333.430 182.610 333.570 ;
        RECT 183.390 333.430 183.700 333.570 ;
        RECT 184.490 333.430 184.800 333.560 ;
        RECT 180.270 333.400 180.650 333.430 ;
        RECT 181.620 333.420 184.800 333.430 ;
        RECT 177.250 333.200 180.650 333.400 ;
        RECT 181.530 333.340 184.800 333.420 ;
        RECT 171.720 333.060 174.870 333.200 ;
        RECT 177.370 333.060 180.650 333.200 ;
        RECT 171.720 332.380 172.040 333.060 ;
        RECT 171.570 332.000 172.040 332.380 ;
        RECT 171.720 330.610 172.040 332.000 ;
        RECT 180.200 333.040 180.650 333.060 ;
        RECT 181.420 333.230 184.800 333.340 ;
        RECT 187.060 333.430 187.370 333.560 ;
        RECT 188.160 333.430 188.470 333.570 ;
        RECT 189.250 333.430 189.560 333.570 ;
        RECT 187.060 333.420 190.240 333.430 ;
        RECT 196.350 333.420 196.650 333.440 ;
        RECT 187.060 333.230 190.330 333.420 ;
        RECT 181.420 333.090 184.680 333.230 ;
        RECT 187.180 333.200 190.330 333.230 ;
        RECT 187.180 333.090 190.670 333.200 ;
        RECT 172.480 330.610 172.790 330.760 ;
        RECT 173.580 330.610 173.890 330.760 ;
        RECT 174.680 330.610 174.990 330.760 ;
        RECT 171.720 330.430 174.990 330.610 ;
        RECT 177.250 330.610 177.560 330.760 ;
        RECT 178.350 330.610 178.660 330.760 ;
        RECT 179.450 330.610 179.760 330.760 ;
        RECT 180.200 330.610 180.520 333.040 ;
        RECT 181.420 333.000 181.850 333.090 ;
        RECT 177.250 330.430 180.520 330.610 ;
        RECT 171.720 330.280 174.880 330.430 ;
        RECT 177.360 330.280 180.520 330.430 ;
        RECT 171.720 329.240 172.040 330.280 ;
        RECT 172.480 329.240 172.790 329.390 ;
        RECT 173.580 329.240 173.890 329.390 ;
        RECT 174.680 329.240 174.990 329.390 ;
        RECT 171.720 329.060 174.990 329.240 ;
        RECT 177.250 329.240 177.560 329.390 ;
        RECT 178.350 329.240 178.660 329.390 ;
        RECT 179.450 329.240 179.760 329.390 ;
        RECT 180.200 329.240 180.520 330.280 ;
        RECT 177.250 329.060 180.520 329.240 ;
        RECT 171.720 328.920 174.880 329.060 ;
        RECT 177.360 328.920 180.520 329.060 ;
        RECT 181.530 330.640 181.850 333.000 ;
        RECT 190.010 332.840 190.670 333.090 ;
        RECT 195.640 333.080 196.660 333.420 ;
        RECT 196.350 333.060 196.660 333.080 ;
        RECT 182.290 330.640 182.600 330.790 ;
        RECT 183.390 330.640 183.700 330.790 ;
        RECT 184.490 330.640 184.800 330.790 ;
        RECT 181.530 330.460 184.800 330.640 ;
        RECT 187.060 330.640 187.370 330.790 ;
        RECT 188.160 330.640 188.470 330.790 ;
        RECT 189.260 330.640 189.570 330.790 ;
        RECT 190.010 330.640 190.330 332.840 ;
        RECT 191.760 332.120 192.210 332.550 ;
        RECT 187.060 330.460 190.330 330.640 ;
        RECT 181.530 330.310 184.690 330.460 ;
        RECT 187.170 330.310 190.330 330.460 ;
        RECT 181.530 329.270 181.850 330.310 ;
        RECT 182.290 329.270 182.600 329.420 ;
        RECT 183.390 329.270 183.700 329.420 ;
        RECT 184.490 329.270 184.800 329.420 ;
        RECT 181.530 329.090 184.800 329.270 ;
        RECT 187.060 329.270 187.370 329.420 ;
        RECT 188.160 329.270 188.470 329.420 ;
        RECT 189.260 329.270 189.570 329.420 ;
        RECT 190.010 329.270 190.330 330.310 ;
        RECT 187.060 329.090 190.330 329.270 ;
        RECT 181.530 328.950 184.690 329.090 ;
        RECT 187.170 328.950 190.330 329.090 ;
        RECT 49.620 326.520 127.730 328.600 ;
        RECT 136.390 327.140 136.760 327.150 ;
        RECT 135.070 326.760 137.680 327.140 ;
        RECT 40.940 215.460 43.390 218.980 ;
        RECT 41.120 215.340 43.200 215.460 ;
        RECT 49.620 161.840 51.700 326.520 ;
        RECT 125.500 326.320 126.770 326.520 ;
        RECT 135.070 326.320 135.450 326.760 ;
        RECT 136.390 326.740 136.760 326.760 ;
        RECT 145.060 326.440 145.340 326.450 ;
        RECT 125.500 325.940 135.450 326.320 ;
        RECT 141.470 326.110 145.360 326.440 ;
        RECT 145.060 326.090 145.340 326.110 ;
        RECT 98.440 325.590 99.040 325.640 ;
        RECT 125.500 325.590 126.770 325.940 ;
        RECT 98.440 325.150 127.780 325.590 ;
        RECT 98.440 325.080 99.040 325.150 ;
        RECT 125.500 325.140 126.770 325.150 ;
        RECT 101.870 324.610 102.330 324.620 ;
        RECT 101.870 324.170 127.740 324.610 ;
        RECT 101.870 324.150 102.330 324.170 ;
        RECT 137.940 323.700 140.650 323.710 ;
        RECT 53.870 321.370 127.730 323.450 ;
        RECT 137.710 323.380 140.650 323.700 ;
        RECT 137.710 323.230 138.330 323.380 ;
        RECT 139.120 323.240 139.430 323.380 ;
        RECT 140.210 323.240 140.520 323.380 ;
        RECT 49.200 158.170 51.910 161.840 ;
        RECT 49.620 157.450 51.700 158.170 ;
        RECT 53.870 133.220 55.950 321.370 ;
        RECT 125.500 321.090 126.770 321.370 ;
        RECT 125.500 320.710 135.470 321.090 ;
        RECT 125.500 320.120 126.770 320.710 ;
        RECT 135.090 319.860 135.470 320.710 ;
        RECT 137.710 320.940 138.060 323.230 ;
        RECT 228.870 322.910 229.070 322.920 ;
        RECT 232.630 322.910 232.950 322.960 ;
        RECT 228.870 322.760 232.950 322.910 ;
        RECT 137.710 320.610 140.660 320.940 ;
        RECT 137.710 320.460 138.330 320.610 ;
        RECT 139.120 320.460 139.430 320.610 ;
        RECT 140.210 320.460 140.520 320.610 ;
        RECT 136.390 319.860 136.760 319.870 ;
        RECT 137.710 319.860 138.060 320.460 ;
        RECT 135.090 319.740 138.060 319.860 ;
        RECT 135.090 319.610 138.090 319.740 ;
        RECT 135.090 319.570 138.460 319.610 ;
        RECT 227.820 319.590 228.080 319.720 ;
        RECT 135.090 319.480 140.650 319.570 ;
        RECT 136.390 319.460 136.760 319.480 ;
        RECT 137.710 319.270 140.650 319.480 ;
        RECT 227.750 319.400 228.080 319.590 ;
        RECT 138.010 319.120 138.320 319.270 ;
        RECT 139.120 319.110 139.430 319.270 ;
        RECT 140.210 319.090 140.520 319.270 ;
        RECT 162.090 317.310 162.510 317.320 ;
        RECT 162.090 317.060 202.360 317.310 ;
        RECT 162.090 316.980 202.370 317.060 ;
        RECT 162.090 316.970 162.510 316.980 ;
        RECT 196.330 316.960 202.370 316.980 ;
        RECT 161.490 316.690 161.870 316.700 ;
        RECT 125.370 314.580 126.640 316.460 ;
        RECT 161.490 316.360 198.290 316.690 ;
        RECT 161.490 316.350 161.870 316.360 ;
        RECT 192.220 316.350 198.290 316.360 ;
        RECT 160.850 316.060 161.270 316.070 ;
        RECT 160.850 315.730 194.210 316.060 ;
        RECT 160.850 315.720 161.270 315.730 ;
        RECT 160.260 315.420 160.660 315.440 ;
        RECT 160.260 315.090 190.200 315.420 ;
        RECT 160.260 315.080 160.660 315.090 ;
        RECT 159.600 314.750 160.010 314.760 ;
        RECT 159.590 314.420 186.110 314.750 ;
        RECT 159.600 314.400 160.010 314.420 ;
        RECT 62.280 312.070 127.730 314.150 ;
        RECT 159.020 314.130 159.430 314.140 ;
        RECT 159.020 314.110 182.090 314.130 ;
        RECT 159.020 313.800 182.100 314.110 ;
        RECT 159.020 313.790 159.430 313.800 ;
        RECT 158.420 313.480 158.810 313.490 ;
        RECT 158.420 313.160 178.110 313.480 ;
        RECT 158.520 313.150 178.110 313.160 ;
        RECT 157.840 312.870 158.230 312.920 ;
        RECT 152.700 312.660 153.240 312.700 ;
        RECT 139.870 312.620 153.240 312.660 ;
        RECT 139.820 312.230 153.240 312.620 ;
        RECT 157.840 312.590 174.200 312.870 ;
        RECT 158.100 312.540 174.200 312.590 ;
        RECT 53.540 129.740 56.280 133.220 ;
        RECT 53.870 128.930 55.950 129.740 ;
        RECT 62.280 76.150 64.360 312.070 ;
        RECT 125.440 309.830 126.710 311.710 ;
        RECT 139.820 310.350 141.830 312.230 ;
        RECT 152.700 312.200 153.240 312.230 ;
        RECT 157.260 311.900 170.000 312.230 ;
        RECT 153.350 311.820 153.890 311.890 ;
        RECT 143.920 311.390 153.890 311.820 ;
        RECT 163.870 311.600 165.890 311.620 ;
        RECT 156.710 311.590 165.920 311.600 ;
        RECT 143.920 310.380 145.900 311.390 ;
        RECT 156.610 311.270 165.920 311.590 ;
        RECT 156.610 311.260 157.000 311.270 ;
        RECT 154.030 311.010 154.520 311.210 ;
        RECT 148.420 310.990 154.520 311.010 ;
        RECT 147.850 310.710 154.520 310.990 ;
        RECT 147.850 310.610 154.430 310.710 ;
        RECT 155.970 310.610 161.950 310.950 ;
        RECT 147.850 310.380 149.830 310.610 ;
        RECT 153.860 310.380 154.510 310.390 ;
        RECT 139.800 309.690 141.830 310.350 ;
        RECT 143.870 309.720 145.900 310.380 ;
        RECT 147.830 309.720 149.860 310.380 ;
        RECT 151.830 309.750 154.510 310.380 ;
        RECT 155.360 310.360 155.910 310.380 ;
        RECT 155.360 309.930 157.910 310.360 ;
        RECT 159.920 310.350 161.960 310.610 ;
        RECT 151.830 309.720 153.860 309.750 ;
        RECT 155.880 309.700 157.910 309.930 ;
        RECT 159.910 309.690 161.960 310.350 ;
        RECT 163.840 309.720 165.920 311.270 ;
        RECT 167.950 310.600 169.980 311.900 ;
        RECT 167.950 310.310 169.990 310.600 ;
        RECT 167.960 309.700 169.990 310.310 ;
        RECT 172.130 309.720 174.160 312.540 ;
        RECT 176.120 310.440 178.110 313.150 ;
        RECT 176.110 309.690 178.140 310.440 ;
        RECT 180.100 310.420 182.100 313.800 ;
        RECT 180.070 309.720 182.100 310.420 ;
        RECT 184.200 310.350 186.110 314.420 ;
        RECT 188.240 310.370 190.190 315.090 ;
        RECT 192.220 310.370 194.210 315.730 ;
        RECT 196.330 316.030 198.290 316.350 ;
        RECT 200.430 316.460 202.370 316.960 ;
        RECT 222.950 316.850 223.380 316.870 ;
        RECT 204.450 316.820 206.410 316.850 ;
        RECT 222.930 316.820 223.390 316.850 ;
        RECT 204.450 316.470 223.390 316.820 ;
        RECT 196.330 310.370 198.280 316.030 ;
        RECT 200.430 310.390 202.360 316.460 ;
        RECT 184.120 309.700 186.150 310.350 ;
        RECT 188.190 309.720 190.220 310.370 ;
        RECT 192.220 309.720 194.250 310.370 ;
        RECT 196.270 309.720 198.300 310.370 ;
        RECT 200.340 309.610 202.370 310.390 ;
        RECT 204.450 310.370 206.410 316.470 ;
        RECT 222.930 316.450 223.390 316.470 ;
        RECT 222.950 316.440 223.380 316.450 ;
        RECT 223.850 316.040 224.280 316.060 ;
        RECT 223.840 316.030 224.290 316.040 ;
        RECT 208.380 315.650 224.290 316.030 ;
        RECT 204.420 309.720 206.450 310.370 ;
        RECT 208.380 310.350 210.340 315.650 ;
        RECT 223.850 315.630 224.280 315.650 ;
        RECT 224.770 315.210 225.220 315.220 ;
        RECT 212.530 314.830 225.220 315.210 ;
        RECT 212.530 310.370 214.510 314.830 ;
        RECT 225.610 314.420 226.030 314.450 ;
        RECT 216.640 314.040 226.030 314.420 ;
        RECT 208.370 309.700 210.400 310.350 ;
        RECT 212.490 309.720 214.520 310.370 ;
        RECT 216.640 310.340 218.620 314.040 ;
        RECT 225.610 314.010 226.030 314.040 ;
        RECT 227.750 311.250 227.950 319.400 ;
        RECT 221.710 311.050 227.950 311.250 ;
        RECT 228.870 311.190 229.070 322.760 ;
        RECT 232.630 322.640 232.950 322.760 ;
        RECT 229.840 321.350 232.650 321.360 ;
        RECT 229.840 321.160 232.950 321.350 ;
        RECT 229.380 311.280 229.700 311.600 ;
        RECT 228.860 311.050 229.070 311.190 ;
        RECT 221.710 310.370 221.910 311.050 ;
        RECT 228.870 310.840 229.070 311.050 ;
        RECT 226.640 310.640 229.070 310.840 ;
        RECT 226.640 310.370 226.840 310.640 ;
        RECT 229.840 310.370 230.050 321.160 ;
        RECT 232.630 321.030 232.950 321.160 ;
        RECT 231.620 319.700 231.930 319.730 ;
        RECT 232.620 319.700 232.940 319.740 ;
        RECT 231.620 319.450 232.940 319.700 ;
        RECT 231.620 314.750 231.920 319.450 ;
        RECT 232.620 319.420 232.940 319.450 ;
        RECT 232.630 317.800 232.950 318.120 ;
        RECT 232.740 316.510 232.930 317.800 ;
        RECT 232.620 316.190 232.940 316.510 ;
        RECT 232.210 314.750 232.530 314.860 ;
        RECT 231.620 314.540 232.530 314.750 ;
        RECT 231.620 314.530 232.380 314.540 ;
        RECT 231.620 313.110 231.920 314.530 ;
        RECT 232.740 313.310 232.930 316.190 ;
        RECT 231.620 312.950 231.980 313.110 ;
        RECT 232.620 312.990 232.940 313.310 ;
        RECT 230.320 311.280 230.640 311.600 ;
        RECT 231.270 311.510 231.590 311.580 ;
        RECT 231.770 311.510 231.980 312.950 ;
        RECT 232.740 311.600 232.930 312.990 ;
        RECT 231.270 311.310 231.980 311.510 ;
        RECT 231.270 311.260 231.590 311.310 ;
        RECT 216.630 309.690 218.660 310.340 ;
        RECT 220.620 309.720 222.650 310.370 ;
        RECT 224.640 310.070 226.840 310.370 ;
        RECT 224.640 309.720 226.670 310.070 ;
        RECT 228.720 309.720 230.750 310.370 ;
        RECT 231.770 310.280 231.980 311.310 ;
        RECT 232.580 311.280 232.930 311.600 ;
        RECT 232.720 311.070 232.930 311.280 ;
        RECT 232.720 311.050 237.740 311.070 ;
        RECT 232.740 310.880 237.740 311.050 ;
        RECT 237.550 310.420 237.740 310.880 ;
        RECT 232.900 310.280 234.930 310.370 ;
        RECT 237.550 310.350 238.580 310.420 ;
        RECT 231.770 310.070 234.930 310.280 ;
        RECT 232.900 309.720 234.930 310.070 ;
        RECT 236.880 309.700 238.910 310.350 ;
        RECT 66.630 306.460 127.730 308.540 ;
        RECT 61.790 72.370 64.620 76.150 ;
        RECT 62.280 71.810 64.360 72.370 ;
        RECT 66.630 47.570 68.710 306.460 ;
        RECT 70.790 301.760 127.730 303.840 ;
        RECT 66.280 43.850 68.930 47.570 ;
        RECT 66.630 43.840 68.710 43.850 ;
        RECT 70.790 18.870 72.870 301.760 ;
        RECT 70.600 15.340 73.270 18.870 ;
        RECT 132.330 9.510 135.670 301.900 ;
        RECT 335.350 246.810 337.440 333.840 ;
        RECT 339.440 275.580 341.530 339.040 ;
        RECT 343.520 304.080 345.610 343.920 ;
        RECT 347.660 332.640 349.750 349.320 ;
        RECT 347.460 329.100 349.890 332.640 ;
        RECT 347.660 328.430 349.750 329.100 ;
        RECT 343.280 300.510 345.790 304.080 ;
        RECT 339.240 271.870 341.760 275.580 ;
        RECT 339.440 271.840 341.530 271.870 ;
        RECT 335.080 243.390 337.440 246.810 ;
        RECT 335.350 242.680 337.440 243.390 ;
      LAYER via2 ;
        RECT 203.190 361.360 203.530 361.700 ;
        RECT 202.120 357.880 202.450 358.230 ;
        RECT 203.210 355.310 203.550 355.670 ;
  END
END sky130_hilas_TopProtectStructure

MACRO sky130_hilas_nFETLarge
  CLASS CORE ;
  FOREIGN sky130_hilas_nFETLarge ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.570 BY 6.030 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    USE ANALOG ;
    ANTENNAGATEAREA 2.642500 ;
    PORT
      LAYER met2 ;
        RECT 0.000 0.330 0.600 0.820 ;
        RECT 0.000 0.000 0.610 0.330 ;
    END
  END GATE
  PIN SOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 1.343400 ;
    PORT
      LAYER met2 ;
        RECT 0.330 5.590 3.390 5.600 ;
        RECT 0.240 5.260 3.390 5.590 ;
        RECT 0.240 2.810 0.560 5.260 ;
        RECT 3.060 5.250 3.370 5.260 ;
        RECT 0.240 2.480 3.400 2.810 ;
        RECT 0.240 1.440 0.560 2.480 ;
        RECT 0.240 1.120 3.400 1.440 ;
        RECT 0.860 1.110 1.170 1.120 ;
        RECT 1.960 1.110 2.270 1.120 ;
        RECT 3.060 1.110 3.370 1.120 ;
    END
  END SOURCE
  PIN DRAIN
    USE ANALOG ;
    ANTENNADIFFAREA 2.723900 ;
    PORT
      LAYER met2 ;
        RECT 1.420 4.880 1.730 4.910 ;
        RECT 2.510 4.880 2.820 4.890 ;
        RECT 1.420 4.580 4.370 4.880 ;
        RECT 2.510 4.560 2.820 4.580 ;
        RECT 3.620 4.540 4.370 4.580 ;
        RECT 3.990 4.410 4.370 4.540 ;
        RECT 4.020 3.540 4.370 4.410 ;
        RECT 1.420 3.210 4.370 3.540 ;
        RECT 4.020 0.770 4.370 3.210 ;
        RECT 1.430 0.760 4.370 0.770 ;
        RECT 1.420 0.450 4.370 0.760 ;
        RECT 1.420 0.440 4.140 0.450 ;
        RECT 1.420 0.430 1.730 0.440 ;
        RECT 2.510 0.430 2.820 0.440 ;
    END
  END DRAIN
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.180 2.450 0.450 2.480 ;
        RECT 0.180 1.920 0.460 2.450 ;
        RECT 0.000 1.620 0.460 1.920 ;
        RECT 0.000 1.600 0.470 1.620 ;
        RECT 0.180 1.170 0.470 1.600 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.880 5.510 1.200 5.550 ;
        RECT 1.970 5.510 2.290 5.550 ;
        RECT 0.880 5.320 1.210 5.510 ;
        RECT 1.970 5.320 2.300 5.510 ;
        RECT 0.880 5.290 1.200 5.320 ;
        RECT 1.970 5.290 2.290 5.320 ;
        RECT 1.430 4.830 1.750 4.870 ;
        RECT 2.600 4.850 2.770 5.890 ;
        RECT 3.150 5.540 3.320 5.890 ;
        RECT 3.070 5.500 3.390 5.540 ;
        RECT 3.070 5.310 3.400 5.500 ;
        RECT 3.070 5.280 3.390 5.310 ;
        RECT 1.430 4.640 1.760 4.830 ;
        RECT 2.520 4.810 2.840 4.850 ;
        RECT 1.430 4.610 1.750 4.640 ;
        RECT 2.520 4.620 2.850 4.810 ;
        RECT 2.520 4.590 2.840 4.620 ;
        RECT 2.600 3.500 2.770 4.590 ;
        RECT 1.430 3.460 1.750 3.500 ;
        RECT 2.520 3.460 2.840 3.500 ;
        RECT 3.150 3.490 3.320 5.280 ;
        RECT 3.700 4.840 3.870 5.890 ;
        RECT 3.630 4.800 3.950 4.840 ;
        RECT 3.630 4.610 3.960 4.800 ;
        RECT 3.630 4.580 3.950 4.610 ;
        RECT 3.700 3.500 3.870 4.580 ;
        RECT 3.620 3.460 3.940 3.500 ;
        RECT 4.250 3.490 4.420 5.890 ;
        RECT 4.800 3.490 4.970 5.890 ;
        RECT 5.350 3.490 5.520 5.890 ;
        RECT 1.430 3.270 1.760 3.460 ;
        RECT 2.520 3.270 2.850 3.460 ;
        RECT 3.620 3.270 3.950 3.460 ;
        RECT 1.430 3.240 1.750 3.270 ;
        RECT 2.520 3.240 2.840 3.270 ;
        RECT 3.620 3.240 3.940 3.270 ;
        RECT 0.950 2.800 1.120 3.180 ;
        RECT 1.500 2.800 1.670 3.180 ;
        RECT 2.050 2.800 2.220 3.180 ;
        RECT 0.870 2.730 1.190 2.770 ;
        RECT 1.970 2.730 2.290 2.770 ;
        RECT 0.870 2.540 1.200 2.730 ;
        RECT 1.970 2.540 2.300 2.730 ;
        RECT 0.870 2.510 1.190 2.540 ;
        RECT 1.970 2.510 2.290 2.540 ;
        RECT 0.240 1.200 0.410 2.420 ;
        RECT 0.870 1.360 1.190 1.400 ;
        RECT 1.970 1.360 2.290 1.400 ;
        RECT 0.870 1.170 1.200 1.360 ;
        RECT 1.970 1.170 2.300 1.360 ;
        RECT 0.870 1.140 1.190 1.170 ;
        RECT 1.970 1.140 2.290 1.170 ;
        RECT 0.190 0.750 0.700 1.010 ;
        RECT 0.190 0.680 0.710 0.750 ;
        RECT 2.600 0.720 2.770 3.180 ;
        RECT 3.150 2.770 3.320 3.180 ;
        RECT 3.070 2.730 3.390 2.770 ;
        RECT 3.070 2.540 3.400 2.730 ;
        RECT 3.070 2.510 3.390 2.540 ;
        RECT 3.150 1.400 3.320 2.510 ;
        RECT 3.070 1.360 3.390 1.400 ;
        RECT 3.070 1.170 3.400 1.360 ;
        RECT 3.070 1.140 3.390 1.170 ;
        RECT 0.200 0.000 0.710 0.680 ;
        RECT 1.430 0.680 1.750 0.720 ;
        RECT 2.520 0.680 2.840 0.720 ;
        RECT 3.150 0.710 3.320 1.140 ;
        RECT 3.700 0.730 3.870 3.180 ;
        RECT 3.620 0.690 3.940 0.730 ;
        RECT 4.250 0.710 4.420 3.110 ;
        RECT 4.800 0.710 4.970 3.110 ;
        RECT 5.350 0.710 5.520 3.110 ;
        RECT 1.430 0.490 1.760 0.680 ;
        RECT 2.520 0.490 2.850 0.680 ;
        RECT 3.620 0.500 3.950 0.690 ;
        RECT 1.430 0.460 1.750 0.490 ;
        RECT 2.520 0.460 2.840 0.490 ;
        RECT 3.620 0.470 3.940 0.500 ;
      LAYER mcon ;
        RECT 0.940 5.330 1.110 5.500 ;
        RECT 2.030 5.330 2.200 5.500 ;
        RECT 3.130 5.320 3.300 5.490 ;
        RECT 1.490 4.650 1.660 4.820 ;
        RECT 2.580 4.630 2.750 4.800 ;
        RECT 3.690 4.620 3.860 4.790 ;
        RECT 1.490 3.280 1.660 3.450 ;
        RECT 2.580 3.280 2.750 3.450 ;
        RECT 3.680 3.280 3.850 3.450 ;
        RECT 0.930 2.550 1.100 2.720 ;
        RECT 2.030 2.550 2.200 2.720 ;
        RECT 0.240 2.250 0.410 2.420 ;
        RECT 0.240 1.890 0.410 2.060 ;
        RECT 0.930 1.180 1.100 1.350 ;
        RECT 2.030 1.180 2.200 1.350 ;
        RECT 3.130 2.550 3.300 2.720 ;
        RECT 3.130 1.180 3.300 1.350 ;
        RECT 0.360 0.540 0.530 0.710 ;
        RECT 1.490 0.500 1.660 0.670 ;
        RECT 2.580 0.500 2.750 0.670 ;
        RECT 3.680 0.510 3.850 0.680 ;
        RECT 0.370 0.070 0.540 0.240 ;
      LAYER met1 ;
        RECT 0.870 5.260 1.190 5.580 ;
        RECT 1.960 5.260 2.280 5.580 ;
        RECT 3.060 5.250 3.380 5.570 ;
        RECT 1.420 4.580 1.740 4.900 ;
        RECT 2.510 4.560 2.830 4.880 ;
        RECT 3.620 4.550 3.940 4.870 ;
        RECT 1.420 3.210 1.740 3.530 ;
        RECT 2.510 3.210 2.830 3.530 ;
        RECT 3.610 3.210 3.930 3.530 ;
        RECT 0.860 2.480 1.180 2.800 ;
        RECT 1.960 2.480 2.280 2.800 ;
        RECT 3.060 2.480 3.380 2.800 ;
        RECT 0.860 1.110 1.180 1.430 ;
        RECT 1.960 1.110 2.280 1.430 ;
        RECT 3.060 1.110 3.380 1.430 ;
        RECT 0.290 0.470 0.610 0.790 ;
        RECT 1.420 0.430 1.740 0.750 ;
        RECT 2.510 0.430 2.830 0.750 ;
        RECT 3.610 0.440 3.930 0.760 ;
        RECT 0.300 0.000 0.620 0.320 ;
      LAYER via ;
        RECT 0.900 5.290 1.160 5.550 ;
        RECT 1.990 5.290 2.250 5.550 ;
        RECT 3.090 5.280 3.350 5.540 ;
        RECT 1.450 4.610 1.710 4.870 ;
        RECT 2.540 4.590 2.800 4.850 ;
        RECT 3.650 4.580 3.910 4.840 ;
        RECT 1.450 3.240 1.710 3.500 ;
        RECT 2.540 3.240 2.800 3.500 ;
        RECT 3.640 3.240 3.900 3.500 ;
        RECT 0.890 2.510 1.150 2.770 ;
        RECT 1.990 2.510 2.250 2.770 ;
        RECT 3.090 2.510 3.350 2.770 ;
        RECT 0.890 1.140 1.150 1.400 ;
        RECT 1.990 1.140 2.250 1.400 ;
        RECT 3.090 1.140 3.350 1.400 ;
        RECT 0.320 0.500 0.580 0.760 ;
        RECT 1.450 0.460 1.710 0.720 ;
        RECT 2.540 0.460 2.800 0.720 ;
        RECT 3.640 0.470 3.900 0.730 ;
        RECT 0.330 0.030 0.590 0.290 ;
  END
END sky130_hilas_nFETLarge

END LIBRARY