magic
tech sky130A
timestamp 1626781805
<< metal1 >>
rect 14 1024 1179 1044
rect 14 471 30 1024
rect 11 455 30 471
rect 11 20 27 455
rect 1156 21 1179 1024
rect 513 20 1179 21
rect 11 7 1179 20
rect 11 6 528 7
<< via1 >>
rect 30 455 1156 1024
rect 27 21 1156 455
rect 27 20 513 21
<< metal2 >>
rect -6 1024 1212 1064
rect -6 455 30 1024
rect -6 20 27 455
rect 1156 21 1212 1024
rect 513 20 1212 21
rect -6 -9 1212 20
<< via2 >>
rect 37 30 1133 1004
<< metal3 >>
rect -25 1004 1232 1087
rect -25 30 37 1004
rect 1133 30 1232 1004
rect -25 -21 1232 30
<< end >>
