magic
tech sky130A
timestamp 1628707374
<< error_p >>
rect 61 98 100 101
rect 61 56 100 59
<< nwell >>
rect 0 0 161 121
<< pmos >>
rect 61 59 100 98
<< pdiff >>
rect 34 87 61 98
rect 34 70 38 87
rect 55 70 61 87
rect 34 59 61 70
rect 100 87 127 98
rect 100 70 106 87
rect 123 70 127 87
rect 100 59 127 70
<< pdiffc >>
rect 38 70 55 87
rect 106 70 123 87
<< poly >>
rect 0 96 26 111
rect 61 98 100 111
rect 11 51 26 96
rect 61 51 100 59
rect 11 36 150 51
rect 135 15 150 36
rect 135 0 161 15
<< locali >>
rect 38 87 55 95
rect 38 62 55 70
rect 106 87 123 95
rect 106 62 123 70
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
