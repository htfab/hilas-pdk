magic
tech sky130A
timestamp 1627742263
<< error_s >>
rect 1135 577 1185 587
rect 1275 577 1325 588
rect 1455 577 1505 588
rect 1072 565 1089 567
rect 1072 546 1089 548
rect 1210 545 1215 550
rect 1245 546 1275 550
rect 1135 535 1185 545
rect 1275 535 1325 546
rect 1455 535 1505 546
rect 1072 531 1089 533
rect 1135 515 1185 526
rect 1072 512 1089 514
rect 1234 509 1239 526
rect 1455 515 1505 526
rect 1185 484 1215 490
rect 1427 484 1455 490
rect 1505 484 1533 490
rect 1135 473 1185 484
rect 1455 473 1505 484
rect 1135 424 1185 435
rect 1455 424 1505 435
rect 1185 418 1215 424
rect 1427 418 1455 424
rect 1505 418 1533 424
rect 1210 399 1215 418
rect 1072 394 1089 396
rect 1234 393 1239 399
rect 1135 382 1185 393
rect 1234 386 1239 387
rect 1234 382 1251 386
rect 1455 382 1505 393
rect 1072 375 1089 377
rect 1135 363 1185 373
rect 1275 362 1325 373
rect 1455 362 1505 373
rect 1072 360 1089 362
rect 1072 341 1089 343
rect 1135 321 1185 331
rect 1275 320 1325 331
rect 1455 320 1505 331
rect 1135 284 1185 294
rect 1275 284 1325 295
rect 1455 284 1505 295
rect 1072 272 1089 274
rect 1072 253 1089 255
rect 1210 252 1215 257
rect 1245 253 1275 257
rect 1135 242 1185 252
rect 1275 242 1325 253
rect 1455 242 1505 253
rect 1072 238 1089 240
rect 1135 222 1185 233
rect 1072 219 1089 221
rect 1234 216 1239 233
rect 1455 222 1505 233
rect 1185 191 1215 197
rect 1427 191 1455 197
rect 1505 191 1533 197
rect 1135 180 1185 191
rect 1455 180 1505 191
rect 1135 131 1185 142
rect 1455 131 1505 142
rect 1185 125 1215 131
rect 1427 125 1455 131
rect 1505 125 1533 131
rect 1210 106 1215 125
rect 1072 101 1089 103
rect 1234 100 1239 106
rect 1135 89 1185 100
rect 1234 93 1239 94
rect 1234 89 1251 93
rect 1455 89 1505 100
rect 1072 82 1089 84
rect 1135 70 1185 80
rect 1275 69 1325 80
rect 1455 69 1505 80
rect 1072 67 1089 69
rect 1072 48 1089 50
rect 1135 28 1185 38
rect 1275 27 1325 38
rect 1455 27 1505 38
<< metal1 >>
rect 1108 603 1133 610
rect 1407 603 1430 610
rect 1542 605 1561 610
rect 1407 5 1430 13
rect 1542 5 1561 12
<< metal2 >>
rect 1055 559 1180 560
rect 1055 543 1249 559
rect 1055 542 1180 543
rect 1614 501 1622 524
rect 1611 384 1622 407
rect 1055 372 1174 374
rect 1055 356 1246 372
rect 1055 258 1107 259
rect 1055 257 1177 258
rect 1055 241 1250 257
rect 1614 208 1622 231
rect 1613 91 1622 114
rect 1055 74 1107 75
rect 1055 57 1253 74
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_2
timestamp 1627742263
transform 1 0 1282 0 1 45
box -232 -40 336 119
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_1
timestamp 1627742263
transform 1 0 1282 0 -1 570
box -232 -40 336 119
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_3
timestamp 1627742263
transform 1 0 1282 0 -1 277
box -232 -40 336 119
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_0
timestamp 1627742263
transform 1 0 1282 0 1 338
box -232 -40 336 119
<< labels >>
rlabel metal2 1107 542 1112 560 0 DRAIN1
port 4 nsew analog default
rlabel metal2 1107 356 1112 374 0 DRAIN2
port 3 nsew analog default
rlabel metal2 1107 241 1112 258 0 DRAIN3
port 2 nsew
rlabel metal2 1107 57 1112 74 0 DRAIN4
port 1 nsew
rlabel metal1 1108 603 1133 610 0 VINJ
port 9 nsew power default
rlabel metal1 1407 603 1430 610 0 DRAIN_MUX
port 10 nsew analog default
rlabel metal1 1407 5 1430 13 0 DRAIN_MUX
port 10 nsew analog default
rlabel metal1 1542 5 1561 12 0 VGND
port 11 nsew ground default
rlabel metal1 1542 605 1561 610 0 VGND
port 11 nsew ground default
rlabel metal2 1613 91 1618 114 0 SELECT4
port 12 nsew
rlabel metal2 1614 208 1622 231 0 SELECT3
port 13 nsew
rlabel metal2 1611 384 1622 407 0 SELECT2
port 14 nsew
rlabel metal2 1614 501 1622 524 0 SELECT1
port 15 nsew
<< end >>
