magic
tech sky130A
timestamp 1607184666
<< error_s >>
rect 609 372 626 373
rect 633 361 634 402
rect 597 349 601 361
rect 633 349 638 361
rect 633 333 634 349
rect 633 301 634 332
rect 633 243 634 272
use sky130_hilas_TACoreBlock2  sky130_hilas_TACoreBlock2_0
timestamp 1607028117
transform 1 0 524 0 1 391
box -61 -192 158 285
<< end >>
