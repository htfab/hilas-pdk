magic
tech sky130A
timestamp 1634057770
<< checkpaint >>
rect -606 1002 838 1018
rect -606 922 907 1002
rect -606 -569 988 922
rect -405 -630 988 -569
<< error_s >>
rect 50 351 77 357
rect 50 309 77 315
rect 50 284 77 290
rect 50 242 77 248
rect 50 201 77 207
rect 50 159 77 165
rect 50 134 77 140
rect 50 92 77 98
<< metal1 >>
rect 96 89 130 661
rect 163 90 190 660
<< metal2 >>
rect 1 322 292 344
rect 0 105 271 128
use sky130_hilas_pFETmirror02  sky130_hilas_pFETmirror02_0
timestamp 1634057728
transform 1 0 225 0 1 0
box 0 0 133 292
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_1
timestamp 1634057729
transform 1 0 24 0 1 241
box 0 0 184 147
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_0
timestamp 1634057729
transform 1 0 24 0 -1 208
box 0 0 184 147
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1634057699
transform 1 0 243 0 1 339
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1634057699
transform 1 0 235 0 1 114
box 0 0 34 33
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1634057708
transform 1 0 178 0 1 237
box 0 0 23 29
<< labels >>
rlabel space 281 322 292 345 0 output2
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
