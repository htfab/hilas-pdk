* Copyright 2020 The Hilas PDK Authors
* 
* This file is part of HILAS.
* 
* HILAS is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published by
* the Free Software Foundation, version 3 of the License.
* 
* HILAS is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
* 
* You should have received a copy of the GNU Lesser General Public License
* along with HILAS.  If not, see <https://www.gnu.org/licenses/>.
* 
* Licensed under the Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
* https://www.gnu.org/licenses/lgpl-3.0.en.html
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
* SPDX-License-Identifier: LGPL-3.0
* 
* 

* NGSPICE file created from sky130_hilas_Trans4small.ext - technology: sky130A

.subckt sky130_hilas_pFETdevice01e a_42_n38# w_n242_n110# $SUB a_n92_n38# a_n160_n84#
X0 a_42_n38# a_n160_n84# a_n92_n38# w_n242_n110# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends

.subckt sky130_hilas_nFET03a m2_150_6# $SUB m2_n222_4# a_n184_n58#
X0 m2_150_6# a_n184_n58# m2_n222_4# $SUB sky130_fd_pr__nfet_01v8 w=350000u l=270000u
.ends

.subckt sky130_hilas_Trans4small NFET_SOURCE1 NFET_GATE1 NFET_SOURCE2 NFET_GATE2 NFET_SOURCE3
+ NFET_GATE3 PFET_SOURCE1 PFET_GATE1 PFET_SOURCE2 PFET_GATE2 PFET_SOURCE3 PFET_GATE3
+ WELL VGND PFET_DRAIN3 PFET_DRAIN2 PFET_DRAIN1 NFET_DRAIN3 NFET_DRAIN2 NFET_DRAIN1
Xsky130_hilas_pFETdevice01e_0 PFET_DRAIN1 WELL VGND PFET_SOURCE1 PFET_GATE1 sky130_hilas_pFETdevice01e
Xsky130_hilas_pFETdevice01e_1 PFET_DRAIN2 WELL VGND PFET_SOURCE2 PFET_GATE2 sky130_hilas_pFETdevice01e
Xsky130_hilas_pFETdevice01e_2 PFET_DRAIN3 WELL VGND PFET_SOURCE3 PFET_GATE3 sky130_hilas_pFETdevice01e
Xsky130_hilas_nFET03a_0 NFET_DRAIN3 VGND NFET_SOURCE3 NFET_GATE3 sky130_hilas_nFET03a
Xsky130_hilas_nFET03a_1 NFET_DRAIN2 VGND NFET_SOURCE2 NFET_GATE2 sky130_hilas_nFET03a
Xsky130_hilas_nFET03a_3 NFET_DRAIN1 VGND NFET_SOURCE1 NFET_GATE1 sky130_hilas_nFET03a
.ends

