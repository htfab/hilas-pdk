magic
tech sky130A
timestamp 1628707300
<< checkpaint >>
rect -626 2929 807 2962
rect -626 2920 809 2929
rect 2410 2920 5324 2962
rect -626 1098 5324 2920
rect -57 994 5324 1098
rect -1 608 5324 994
rect 1134 501 5178 608
rect 1136 310 5178 501
rect 2014 263 5178 310
rect 3033 216 5178 263
rect 3033 -630 4842 216
<< error_s >>
rect 1567 1475 1617 1481
rect 1639 1475 1689 1481
rect 3608 1475 3658 1481
rect 3680 1475 3730 1481
rect 4068 1479 4095 1485
rect 1567 1433 1617 1439
rect 1639 1433 1689 1439
rect 3608 1433 3658 1439
rect 3680 1433 3730 1439
rect 4068 1437 4095 1443
rect 4068 1412 4095 1418
rect 1752 1331 1755 1381
rect 1794 1331 1797 1381
rect 1888 1331 1890 1381
rect 1930 1331 1932 1381
rect 4068 1370 4095 1376
rect 4068 1329 4095 1335
rect 1752 1252 1755 1302
rect 1794 1252 1797 1302
rect 1888 1252 1890 1302
rect 1930 1252 1932 1302
rect 4068 1287 4095 1293
rect 4068 1262 4095 1268
rect 4068 1220 4095 1226
rect 4068 1179 4095 1185
rect 1752 1099 1755 1149
rect 1794 1099 1797 1149
rect 1888 1099 1890 1149
rect 1930 1099 1932 1149
rect 4068 1137 4095 1143
rect 4068 1112 4095 1118
rect 4068 1070 4095 1076
rect 1752 1020 1755 1070
rect 1794 1020 1797 1070
rect 1888 1020 1890 1070
rect 1930 1020 1932 1070
rect 4068 1029 4095 1035
rect 4068 987 4095 993
rect 1567 962 1617 968
rect 1639 962 1689 968
rect 3608 962 3658 968
rect 3680 962 3730 968
rect 4068 962 4095 968
rect 1567 920 1617 926
rect 1639 920 1689 926
rect 3608 920 3658 926
rect 3680 920 3730 926
rect 4068 920 4095 926
<< nwell >>
rect 1500 1502 1831 1503
rect 3797 1502 3931 1503
rect 1520 1471 1552 1501
rect 3747 1471 3779 1501
rect 4182 1485 4310 1503
rect 4182 898 4310 917
<< metal1 >>
rect 1536 1501 1552 1503
rect 1520 1499 1552 1501
rect 1520 1473 1523 1499
rect 1549 1473 1552 1499
rect 1577 1497 1596 1503
rect 1764 1492 1785 1503
rect 1811 1495 1830 1503
rect 1852 1497 1873 1503
rect 1960 1496 1978 1503
rect 2576 1488 2618 1503
rect 2679 1488 2721 1503
rect 3049 1495 3072 1503
rect 3701 1495 3720 1503
rect 3745 1501 3773 1503
rect 3745 1499 3779 1501
rect 3745 1495 3750 1499
rect 2576 1474 2721 1488
rect 1520 1471 1552 1473
rect 3747 1473 3750 1495
rect 3776 1473 3779 1499
rect 4114 1489 4148 1503
rect 4180 1488 4208 1503
rect 3747 1471 3779 1473
rect 3961 946 3993 948
rect 2342 931 2374 933
rect 1765 899 1788 911
rect 2342 905 2345 931
rect 2371 905 2374 931
rect 2342 903 2374 905
rect 2922 931 2954 933
rect 2922 905 2925 931
rect 2951 905 2954 931
rect 3961 920 3964 946
rect 3990 920 3993 946
rect 3961 918 3993 920
rect 3961 915 4004 918
rect 4064 917 4115 918
rect 4064 915 4148 917
rect 3961 912 4148 915
rect 3976 907 4148 912
rect 2922 903 2954 905
rect 3979 904 4148 907
rect 3701 898 3720 903
rect 3745 898 3773 903
rect 3982 902 4148 904
rect 3989 901 4085 902
rect 4114 898 4148 902
rect 4181 898 4208 919
<< via1 >>
rect 1523 1473 1549 1499
rect 3750 1473 3776 1499
rect 2345 905 2371 931
rect 2925 905 2951 931
rect 3964 920 3990 946
<< metal2 >>
rect 1520 1499 1552 1501
rect 1520 1473 1523 1499
rect 1549 1489 1552 1499
rect 3747 1499 3779 1501
rect 3747 1489 3750 1499
rect 1549 1473 3750 1489
rect 3776 1473 3779 1499
rect 3857 1476 3888 1500
rect 1520 1471 3779 1473
rect 1500 1435 1508 1453
rect 3968 1413 3990 1415
rect 3963 1379 3990 1413
rect 3789 1329 3824 1351
rect 3970 1322 3990 1323
rect 2651 1280 3450 1300
rect 3970 1289 3992 1322
rect 3972 1288 3992 1289
rect 3310 1212 3332 1213
rect 2652 1187 3335 1212
rect 3428 1208 3450 1280
rect 3865 1209 3897 1233
rect 4299 1232 4310 1255
rect 2652 1095 3003 1114
rect 2980 1035 3003 1095
rect 3306 1070 3335 1187
rect 3425 1204 3450 1208
rect 3425 1140 3451 1204
rect 4299 1150 4310 1172
rect 3425 1119 3838 1140
rect 3817 1105 3838 1119
rect 3817 1084 4018 1105
rect 3306 1048 3595 1070
rect 3306 1047 3335 1048
rect 2980 1020 3002 1035
rect 3417 1020 4017 1025
rect 2980 1005 4017 1020
rect 2980 1004 4004 1005
rect 2980 998 3456 1004
rect 1500 948 1508 966
rect 3961 946 3993 948
rect 3961 933 3964 946
rect 2342 931 3964 933
rect 2342 905 2345 931
rect 2371 918 2925 931
rect 2371 905 2374 918
rect 2342 903 2374 905
rect 2922 905 2925 918
rect 2951 920 3964 931
rect 3990 920 3993 946
rect 2951 918 3993 920
rect 2951 905 2954 918
rect 2922 903 2954 905
use sky130_hilas_FGBias2x1cell  sky130_hilas_FGBias2x1cell_0
timestamp 1628707287
transform 1 0 3040 0 1 1280
box 0 0 1654 1052
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1628707287
transform 1 0 3663 0 -1 1063
box 0 0 549 1063
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1628707291
transform 1 0 4155 0 1 939
box 0 0 358 746
use sky130_hilas_FGtrans2x1cell  sky130_hilas_FGtrans2x1cell_0
timestamp 1628707287
transform -1 0 2257 0 1 1280
box 0 0 2257 1052
<< labels >>
rlabel metal1 4114 1497 4148 1503 0 VGND
port 11 nsew
rlabel metal1 4180 1497 4208 1503 0 VPWR
port 10 nsew
rlabel metal1 4181 898 4208 904 0 VPWR
port 10 nsew
rlabel metal1 4114 898 4148 904 0 VGND
port 11 nsew
rlabel metal2 3865 1209 3897 1233 0 VIN21
port 9 nsew
rlabel metal2 3857 1476 3888 1500 1 VIN22
port 8 n
rlabel metal1 1765 899 1788 911 0 VIN12
port 18 nsew
rlabel metal1 1764 1492 1785 1503 0 VIN11
port 5 nsew
rlabel metal1 2679 1496 2721 1503 0 VTUN
port 1 nsew
rlabel metal1 2576 1496 2618 1503 0 VTUN
rlabel metal1 1852 1497 1873 1503 0 PROG
port 3 nsew
rlabel metal1 1536 1497 1552 1503 0 VINJ
port 6 nsew
rlabel metal1 3745 1495 3773 1503 0 VINJ
port 6 nsew
rlabel metal2 4299 1232 4310 1255 0 OUTPUT1
port 13 nsew
rlabel metal2 4299 1150 4310 1172 0 OUTPUT2
port 12 nsew
rlabel metal1 1577 1497 1596 1503 0 GATESEL1
port 14 nsew
rlabel metal1 3701 898 3720 903 0 GATESEL2
port 15 nsew
rlabel metal1 3745 898 3773 903 0 VINJ
port 6 nsew
rlabel metal1 3701 1495 3720 1503 0 GATESEL2
port 15 nsew
rlabel metal2 1500 1435 1508 1453 0 DRAIN1
port 16 nsew
rlabel metal2 1500 948 1508 966 0 DRAIN2
port 17 nsew
rlabel metal1 3049 1495 3072 1503 0 GATE1
port 4 nsew
rlabel metal1 1811 1495 1830 1503 0 GATE2
port 19 nsew
rlabel metal1 1960 1496 1978 1503 0 RUN
port 20 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
