magic
tech sky130A
timestamp 1628704274
<< metal1 >>
rect 771 1164 1160 1244
rect 3630 1164 4019 1244
rect 6489 1164 6878 1244
rect 10679 1166 11068 1246
rect 14891 1164 15280 1244
rect 17750 1164 18139 1244
rect 20610 1164 20999 1244
rect 23469 1164 23858 1244
rect 26327 1164 26716 1244
rect 29186 1164 29575 1244
rect 32046 1164 32435 1244
rect 1253 0 1648 77
rect 4113 0 4508 77
rect 6971 0 7366 77
rect 11248 0 11496 77
rect 15373 1 15768 78
rect 18232 0 18627 77
rect 21091 0 21486 77
rect 23950 0 24345 77
rect 26810 0 27205 77
rect 29668 0 30063 77
rect 32527 0 32922 77
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_1
timestamp 1627735001
transform 1 0 3604 0 1 306
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_0
timestamp 1627735001
transform 1 0 745 0 1 306
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_2
timestamp 1627735001
transform 1 0 6463 0 1 306
box -745 -229 2114 858
use sky130_hilas_polyresistorGND  sky130_hilas_polyresistorGND_0
timestamp 1627736296
transform 1 0 11322 0 1 134
box -2749 -57 2798 1032
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_3
timestamp 1627735001
transform 1 0 14865 0 1 306
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_4
timestamp 1627735001
transform 1 0 17724 0 1 306
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_5
timestamp 1627735001
transform 1 0 20583 0 1 306
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_6
timestamp 1627735001
transform 1 0 23442 0 1 306
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_9
timestamp 1627735001
transform 1 0 26301 0 1 306
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_7
timestamp 1627735001
transform 1 0 29160 0 1 306
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_8
timestamp 1627735001
transform 1 0 32019 0 1 306
box -745 -229 2114 858
<< labels >>
rlabel metal1 32046 1164 32435 1244 0 ANALOG00
port 1 nsew
rlabel metal1 29186 1164 29575 1244 0 ANALOG01
port 2 nsew
rlabel metal1 26327 1164 26716 1244 0 ANALOG02
port 3 nsew
rlabel metal1 23469 1164 23858 1244 0 ANALOG03
port 4 nsew
rlabel metal1 20610 1164 20999 1244 0 ANALOG04
port 5 nsew
rlabel metal1 17750 1164 18139 1244 0 ANALOG05
port 6 nsew
rlabel metal1 14891 1164 15280 1244 0 ANALOG06
port 7 nsew
rlabel metal1 10679 1166 11068 1246 0 ANALOG07
port 8 nsew
rlabel metal1 6489 1164 6878 1244 0 ANALOG08
port 9 nsew
rlabel metal1 3630 1164 4019 1244 0 ANALOG09
port 10 nsew
rlabel metal1 771 1164 1160 1244 0 ANALOG10
port 11 nsew
rlabel metal1 32527 0 32922 77 0 PIN1
port 12 nsew
rlabel metal1 29668 0 30063 77 0 PIN2
port 13 nsew
rlabel metal1 26810 0 27205 77 0 PIN3
port 14 nsew
rlabel metal1 23950 0 24345 77 0 PIN4
port 15 nsew
rlabel metal1 21091 0 21486 77 0 PIN5
port 16 nsew
rlabel metal1 18232 0 18627 77 0 PIN6
port 17 nsew
rlabel metal1 15373 1 15768 78 0 PIN7
port 18 nsew
rlabel metal1 6971 0 7366 77 0 PIN8
port 19 nsew
rlabel metal1 4113 0 4508 77 0 PIN9
port 20 nsew
rlabel metal1 1253 0 1648 77 0 PIN10
port 21 nsew
rlabel metal1 11248 0 11496 77 0 VTUN
port 22 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
