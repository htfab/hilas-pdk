magic
tech sky130A
timestamp 1628617052
<< checkpaint >>
rect -589 929 918 937
rect -599 789 918 929
rect -599 780 920 789
rect -599 -360 934 780
rect -584 -507 934 -360
rect -584 -600 925 -507
rect -584 -608 915 -600
<< nwell >>
rect 0 156 308 302
<< nmos >>
rect 48 58 259 118
<< pmos >>
rect 48 199 259 260
<< ndiff >>
rect 19 114 48 118
rect 19 97 25 114
rect 42 97 48 114
rect 19 80 48 97
rect 19 63 25 80
rect 42 63 48 80
rect 19 58 48 63
rect 259 114 288 118
rect 259 97 265 114
rect 282 97 288 114
rect 259 80 288 97
rect 259 63 265 80
rect 282 63 288 80
rect 259 58 288 63
<< pdiff >>
rect 19 254 48 260
rect 19 237 25 254
rect 42 237 48 254
rect 19 220 48 237
rect 19 203 25 220
rect 42 203 48 220
rect 19 199 48 203
rect 259 255 289 260
rect 259 238 265 255
rect 283 238 289 255
rect 259 221 289 238
rect 259 203 265 221
rect 283 203 289 221
rect 259 199 289 203
<< ndiffc >>
rect 25 97 42 114
rect 25 63 42 80
rect 265 97 282 114
rect 265 63 282 80
<< pdiffc >>
rect 25 237 42 254
rect 25 203 42 220
rect 265 238 283 255
rect 265 203 283 221
<< poly >>
rect 48 260 259 273
rect 48 181 259 199
rect 48 180 149 181
rect 81 153 82 180
rect 115 153 116 180
rect 222 133 223 159
rect 256 133 257 159
rect 189 132 259 133
rect 48 118 259 132
rect 48 45 259 58
<< locali >>
rect 17 296 291 302
rect 17 295 76 296
rect 84 295 183 296
rect 193 295 291 296
rect 17 255 291 295
rect 17 254 265 255
rect 17 237 25 254
rect 42 238 265 254
rect 283 238 291 255
rect 42 237 291 238
rect 17 221 291 237
rect 17 220 265 221
rect 17 203 25 220
rect 42 203 265 220
rect 283 203 291 221
rect 17 199 291 203
rect 17 114 149 180
rect 189 137 291 199
rect 17 97 25 114
rect 42 97 265 114
rect 282 97 291 114
rect 17 80 291 97
rect 17 63 25 80
rect 42 63 265 80
rect 282 63 291 80
rect 17 25 291 63
<< metal1 >>
rect 17 254 291 302
rect 17 1 291 63
rect 17 0 290 1
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1628616972
transform 1 0 56 0 1 30
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1628616972
transform 1 0 92 0 1 30
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_3
timestamp 1628616972
transform 1 0 128 0 1 30
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_5
timestamp 1628616972
transform 1 0 164 0 1 30
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_2
timestamp 1628616972
transform 1 0 200 0 1 30
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_4
timestamp 1628616972
transform 1 0 236 0 1 30
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_7
timestamp 1628616972
transform 1 0 272 0 1 30
box 0 0 23 29
use sky130_hilas_poly2li  sky130_hilas_poly2li_2
timestamp 1628617008
transform 0 1 96 -1 0 171
box 0 0 27 33
use sky130_hilas_poly2li  sky130_hilas_poly2li_1
timestamp 1628617008
transform 0 1 62 -1 0 171
box 0 0 27 33
use sky130_hilas_poly2li  sky130_hilas_poly2li_5
timestamp 1628617008
transform 0 1 130 -1 0 171
box 0 0 27 33
use sky130_hilas_poly2li  sky130_hilas_poly2li_4
timestamp 1628617008
transform 0 1 203 -1 0 150
box 0 0 27 33
use sky130_hilas_poly2li  sky130_hilas_poly2li_0
timestamp 1628617008
transform 0 1 237 -1 0 150
box 0 0 27 33
use sky130_hilas_poly2li  sky130_hilas_poly2li_3
timestamp 1628617008
transform 0 1 271 -1 0 150
box 0 0 27 33
use sky130_hilas_li2m1  sky130_hilas_li2m1_9
timestamp 1628616972
transform 1 0 41 0 1 278
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_10
timestamp 1628616972
transform 1 0 77 0 1 278
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_11
timestamp 1628616972
transform 1 0 113 0 1 278
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_12
timestamp 1628616972
transform 1 0 149 0 1 278
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_13
timestamp 1628616972
transform 1 0 185 0 1 278
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_14
timestamp 1628616972
transform 1 0 221 0 1 278
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_15
timestamp 1628616972
transform 1 0 265 0 1 278
box 0 0 23 29
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
