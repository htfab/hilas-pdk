magic
tech sky130A
timestamp 1628616694
<< error_p >>
rect 50 111 79 129
rect 50 79 51 80
rect 78 79 79 80
rect 0 50 18 79
rect 49 78 80 79
rect 50 69 79 78
rect 50 60 60 69
rect 69 60 79 69
rect 50 51 79 60
rect 49 50 80 51
rect 111 50 129 79
rect 50 49 51 50
rect 78 49 79 50
rect 50 0 79 18
<< mvnmos >>
rect 18 79 111 111
rect 18 50 50 79
rect 79 50 111 79
rect 18 18 111 50
<< mvndiff >>
rect 50 73 79 79
rect 50 56 56 73
rect 73 56 79 73
rect 50 50 79 56
<< mvndiffc >>
rect 56 56 73 73
<< poly >>
rect 5 111 124 124
rect 5 18 18 111
rect 111 18 124 111
rect 5 5 124 18
<< locali >>
rect 56 107 73 110
rect 56 73 73 90
rect 56 38 73 56
<< viali >>
rect 56 90 73 107
rect 56 21 73 38
<< metal1 >>
rect 53 107 76 129
rect 53 90 56 107
rect 73 90 76 107
rect 53 38 76 90
rect 53 21 56 38
rect 73 21 76 38
rect 53 0 76 21
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
