VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_pFETdevice01e
  CLASS BLOCK ;
  FOREIGN /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_pFETdevice01e ;
  ORIGIN 1.210 0.550 ;
  SIZE 2.030 BY 0.990 ;
  OBS
      LAYER nwell ;
        RECT -1.210 -0.550 0.820 0.440 ;
      LAYER li1 ;
        RECT -1.040 -0.460 0.770 0.230 ;
      LAYER met1 ;
        RECT -1.100 -0.520 0.750 0.260 ;
      LAYER met2 ;
        RECT -1.210 -0.520 0.740 0.270 ;
  END
END /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_pFETdevice01e
END LIBRARY

