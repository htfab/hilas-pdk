magic
tech sky130A
timestamp 1629137187
<< checkpaint >>
rect -560 1111 939 1204
rect -560 956 948 1111
rect -575 -352 948 956
rect -560 -507 948 -352
rect -560 -600 939 -507
<< psubdiff >>
rect 330 31 331 114
<< locali >>
rect 305 490 324 579
rect 305 25 331 114
<< metal1 >>
rect 0 541 35 604
rect 0 525 262 541
rect 296 550 403 604
rect 296 541 315 550
rect 288 525 315 541
rect 0 524 315 525
rect 341 524 403 550
rect 0 510 403 524
rect 0 509 315 510
rect 0 483 260 509
rect 286 484 315 509
rect 341 484 403 510
rect 286 483 403 484
rect 0 473 403 483
rect 0 419 403 442
rect 0 392 51 419
rect 78 392 106 419
rect 133 392 403 419
rect 0 362 403 392
rect 0 361 106 362
rect 0 334 50 361
rect 77 335 106 361
rect 133 335 403 362
rect 77 334 403 335
rect 0 278 403 334
rect 0 277 106 278
rect 0 250 51 277
rect 78 251 106 277
rect 133 251 403 278
rect 78 250 403 251
rect 0 227 403 250
rect 0 200 51 227
rect 78 225 403 227
rect 78 200 104 225
rect 0 198 104 200
rect 131 198 403 225
rect 0 163 403 198
rect 0 100 403 127
rect 0 74 276 100
rect 302 74 324 100
rect 350 74 403 100
rect 0 59 403 74
rect 0 33 274 59
rect 300 33 323 59
rect 349 33 403 59
rect 0 3 403 33
rect 0 0 36 3
rect 305 1 403 3
rect 304 0 403 1
<< via1 >>
rect 262 525 288 551
rect 315 524 341 550
rect 260 483 286 509
rect 315 484 341 510
rect 51 392 78 419
rect 106 392 133 419
rect 50 334 77 361
rect 106 335 133 362
rect 51 250 78 277
rect 106 251 133 278
rect 51 200 78 227
rect 104 198 131 225
rect 276 74 302 100
rect 324 74 350 100
rect 274 33 300 59
rect 323 33 349 59
<< metal2 >>
rect 36 419 166 604
rect 36 392 51 419
rect 78 392 106 419
rect 133 392 166 419
rect 36 362 166 392
rect 36 361 106 362
rect 36 334 50 361
rect 77 335 106 361
rect 133 335 166 362
rect 77 334 166 335
rect 36 278 166 334
rect 36 277 106 278
rect 36 250 51 277
rect 78 251 106 277
rect 133 251 166 278
rect 78 250 166 251
rect 36 227 166 250
rect 36 200 51 227
rect 78 225 166 227
rect 78 200 104 225
rect 36 198 104 200
rect 131 198 166 225
rect 36 0 166 198
rect 244 551 374 604
rect 244 525 262 551
rect 288 550 374 551
rect 288 525 315 550
rect 244 524 315 525
rect 341 524 374 550
rect 244 510 374 524
rect 244 509 315 510
rect 244 483 260 509
rect 286 484 315 509
rect 341 484 374 510
rect 286 483 374 484
rect 244 462 374 483
rect 244 132 373 462
rect 244 100 374 132
rect 244 74 276 100
rect 302 74 324 100
rect 350 74 374 100
rect 244 59 374 74
rect 244 33 274 59
rect 300 33 323 59
rect 349 33 374 59
rect 244 0 374 33
use sky130_hilas_DecoupVinj00  CapDeco_0
timestamp 1625358249
transform 1 0 -68 0 -1 491
box 68 -113 473 189
use sky130_hilas_DecoupVinj00  CapDeco_1
timestamp 1625358249
transform 1 0 -68 0 1 113
box 68 -113 473 189
<< labels >>
rlabel metal1 14 0 23 63 0 VGND 
port 1 nsew
rlabel metal1 388 0 403 63 0 VGND 
port 1 nsew
rlabel metal2 36 594 166 604 0 VINJ
port 1 nsew
rlabel metal2 244 596 374 604 0 VGND
port 2 nsew
rlabel metal2 36 0 166 12 0 VINJ
port 1 nsew
rlabel metal2 244 0 374 12 0 VGND
port 2 nsew
rlabel metal1 386 256 403 350 0 VINJ
port 1 nsew
rlabel metal1 0 254 17 350 0 VINJ
port 1 nsew
rlabel metal1 14 541 22 604 0 VGND
port 3 nsew
rlabel metal1 393 541 403 604 0 VGND
port 2 nsew
<< end >>
