magic
tech sky130A
timestamp 1632494644
<< nmos >>
rect -18 -34 2 25
rect 88 -34 108 25
<< ndiff >>
rect 116 25 146 33
rect -47 21 -18 25
rect -47 4 -41 21
rect -24 4 -18 21
rect -47 -13 -18 4
rect -47 -30 -41 -13
rect -24 -30 -18 -13
rect -47 -34 -18 -30
rect 2 21 32 25
rect 2 4 9 21
rect 26 4 32 21
rect 2 -13 32 4
rect 2 -30 9 -13
rect 26 -30 32 -13
rect 2 -34 32 -30
rect 59 21 88 25
rect 59 4 65 21
rect 82 4 88 21
rect 59 -13 88 4
rect 59 -30 65 -13
rect 82 -30 88 -13
rect 59 -34 88 -30
rect 108 21 146 25
rect 108 4 122 21
rect 139 4 146 21
rect 108 -13 146 4
rect 108 -30 122 -13
rect 139 -30 146 -13
rect 108 -34 146 -30
rect 116 -42 146 -34
<< ndiffc >>
rect -41 4 -24 21
rect -41 -30 -24 -13
rect 9 4 26 21
rect 9 -30 26 -13
rect 65 4 82 21
rect 65 -30 82 -13
rect 122 4 139 21
rect 122 -30 139 -13
<< psubdiff >>
rect 146 21 175 33
rect 146 4 156 21
rect 173 4 175 21
rect 146 -13 175 4
rect 146 -30 156 -13
rect 173 -30 175 -13
rect 146 -42 175 -30
<< psubdiffcont >>
rect 156 4 173 21
rect 156 -30 173 -13
<< poly >>
rect 43 61 108 66
rect 43 44 51 61
rect 68 44 108 61
rect 43 38 108 44
rect -18 25 2 38
rect 88 25 108 38
rect -18 -43 2 -34
rect -63 -53 2 -43
rect 88 -47 108 -34
rect -63 -70 -55 -53
rect -38 -70 2 -53
rect -63 -75 2 -70
<< polycont >>
rect 51 44 68 61
rect -55 -70 -38 -53
<< locali >>
rect 11 61 32 63
rect 9 44 13 61
rect 30 44 51 61
rect 68 44 76 61
rect 9 21 34 44
rect 122 21 173 29
rect -50 4 -41 21
rect -24 4 -16 21
rect 1 4 9 21
rect 26 4 34 21
rect 56 4 65 21
rect 82 4 90 21
rect 139 4 156 21
rect -50 -13 -16 4
rect 9 -13 26 4
rect 65 -13 82 4
rect 122 -13 139 4
rect 156 -13 173 4
rect -50 -30 -41 -13
rect -24 -30 -16 -13
rect 1 -30 9 -13
rect 26 -30 34 -13
rect 56 -30 65 -13
rect 82 -30 90 -13
rect 139 -30 156 -13
rect 65 -53 82 -30
rect 122 -38 173 -30
rect -64 -70 -55 -53
rect -38 -70 82 -53
<< viali >>
rect 13 44 30 61
rect 139 -13 156 4
<< metal1 >>
rect 10 61 33 67
rect 10 44 13 61
rect 30 44 33 61
rect 10 -76 33 44
rect 136 4 159 53
rect 136 -13 139 4
rect 156 -13 159 4
rect 136 -76 159 -13
<< metal2 >>
rect -54 -2 175 14
rect -108 -72 -96 -51
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1632488964
transform 1 0 -69 0 1 7
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1632488964
transform 1 0 -84 0 1 -61
box -14 -15 20 18
<< end >>
