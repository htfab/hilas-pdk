magic
tech sky130A
timestamp 1628698498
<< metal3 >>
rect -392 333 -161 336
rect -392 -245 31 333
rect -164 -247 31 -245
<< mimcap >>
rect -332 -104 -10 295
rect -332 -118 -288 -104
rect -274 -118 -260 -104
rect -246 -118 -232 -104
rect -218 -118 -204 -104
rect -190 -118 -176 -104
rect -162 -118 -149 -104
rect -135 -118 -121 -104
rect -107 -118 -93 -104
rect -79 -118 -10 -104
rect -332 -205 -10 -118
<< mimcapcontact >>
rect -288 -118 -274 -104
rect -260 -118 -246 -104
rect -232 -118 -218 -104
rect -204 -118 -190 -104
rect -176 -118 -162 -104
rect -149 -118 -135 -104
rect -121 -118 -107 -104
rect -93 -118 -79 -104
<< metal4 >>
rect -354 -104 -53 -90
rect -354 -118 -288 -104
rect -274 -118 -260 -104
rect -246 -118 -232 -104
rect -218 -118 -204 -104
rect -190 -118 -176 -104
rect -162 -118 -149 -104
rect -135 -118 -121 -104
rect -107 -118 -93 -104
rect -79 -118 -53 -104
rect -354 -137 -53 -118
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
