VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_FGBias2x1cell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_FGBias2x1cell ;
  ORIGIN 3.960 3.820 ;
  SIZE 11.530 BY 6.050 ;
  PIN Vtun
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT -3.610 0.440 -3.190 2.230 ;
    END
    PORT
      LAYER met1 ;
        RECT -3.610 -3.820 -3.190 -1.560 ;
    END
  END Vtun
  PIN GND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT -1.130 -0.770 -0.900 2.230 ;
    END
    PORT
      LAYER met1 ;
        RECT -1.130 -3.820 -0.900 -0.940 ;
    END
  END GND
  PIN gate_control
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 0.090 0.940 0.320 2.230 ;
    END
  END gate_control
  PIN Gate_control
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 0.090 -3.820 0.320 -2.630 ;
    END
  END Gate_control
  PIN drain1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -3.960 1.550 5.110 1.730 ;
    END
  END drain1
  PIN drain4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -3.960 -3.300 5.110 -3.150 ;
    END
  END drain4
  PIN Vinj
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 7.050 1.520 7.330 2.230 ;
    END
  END Vinj
  PIN output1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.530 0.490 7.570 0.710 ;
    END
  END output1
  PIN output2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.530 -2.260 7.570 -2.050 ;
    END
  END output2
  OBS
      LAYER li1 ;
        RECT -3.520 -3.490 7.180 1.900 ;
      LAYER met1 ;
        RECT -2.910 0.160 -1.410 2.230 ;
        RECT -3.610 -1.280 -1.410 0.160 ;
        RECT -2.910 -3.820 -1.410 -1.280 ;
        RECT -0.620 0.660 -0.190 2.230 ;
        RECT 0.600 1.240 6.770 2.230 ;
        RECT 0.600 0.660 7.410 1.240 ;
        RECT -0.620 -2.350 7.410 0.660 ;
        RECT -0.620 -3.820 -0.190 -2.350 ;
        RECT 0.600 -3.820 7.410 -2.350 ;
      LAYER met2 ;
        RECT 5.390 1.270 7.570 1.930 ;
        RECT 4.840 0.990 7.570 1.270 ;
        RECT 4.840 0.210 5.250 0.990 ;
        RECT 4.840 -1.770 7.570 0.210 ;
        RECT 4.840 -2.540 5.250 -1.770 ;
        RECT 4.840 -2.870 7.570 -2.540 ;
        RECT 5.390 -3.520 7.570 -2.870 ;
  END
END sky130_hilas_FGBias2x1cell
END LIBRARY

