VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_nfetmirrorpairs2
  CLASS BLOCK ;
  FOREIGN sky130_hilas_nfetmirrorpairs2 ;
  ORIGIN 3.090 1.920 ;
  SIZE 4.670 BY 4.770 ;
  OBS
      LAYER nwell ;
        RECT -0.610 1.120 1.580 2.850 ;
      LAYER li1 ;
        RECT -0.400 2.010 1.360 2.530 ;
        RECT -0.400 1.400 0.310 1.570 ;
        RECT 0.620 1.400 1.320 1.570 ;
        RECT -0.050 1.230 0.310 1.400 ;
        RECT -0.050 0.870 0.600 1.230 ;
        RECT -0.050 0.640 0.220 0.870 ;
        RECT 0.850 0.650 1.100 1.400 ;
        RECT -0.080 0.470 0.250 0.640 ;
        RECT 0.770 0.470 1.100 0.650 ;
        RECT -0.120 -0.200 0.290 0.040 ;
        RECT 0.730 -0.200 1.140 0.040 ;
        RECT -0.120 -0.580 1.140 -0.200 ;
        RECT -0.120 -0.840 0.290 -0.580 ;
        RECT 0.730 -0.830 1.140 -0.580 ;
        RECT -0.090 -1.430 0.250 -1.260 ;
        RECT 0.760 -1.430 1.120 -1.250 ;
        RECT -0.010 -1.920 0.170 -1.430 ;
        RECT 0.840 -1.920 1.030 -1.430 ;
  END
END sky130_hilas_nfetmirrorpairs2
END LIBRARY

