magic
tech sky130A
timestamp 1632251359
<< metal1 >>
rect 39 1045 1204 1065
rect 39 492 55 1045
rect 36 476 55 492
rect 36 41 52 476
rect 1181 42 1204 1045
rect 538 41 1204 42
rect 36 28 1204 41
rect 36 27 553 28
<< via1 >>
rect 55 476 1181 1045
rect 52 42 1181 476
rect 52 41 538 42
<< metal2 >>
rect 19 1045 1237 1085
rect 19 476 55 1045
rect 19 41 52 476
rect 1181 42 1237 1045
rect 538 41 1237 42
rect 19 12 1237 41
<< via2 >>
rect 62 51 1158 1025
<< metal3 >>
rect 0 1025 1257 1108
rect 0 51 62 1025
rect 1158 51 1257 1025
rect 0 0 1257 51
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
