VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_hilas_VinjDiodeProtect01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_VinjDiodeProtect01 ;
  ORIGIN 7.450 2.290 ;
  SIZE 28.590 BY 10.870 ;
  PIN OUTPUT 
    ANTENNADIFFAREA 58.900799 ;
    PORT
      LAYER met1 ;
        RECT 6.900 7.960 7.250 8.120 ;
        RECT 6.890 7.010 7.260 7.960 ;
        RECT 6.540 6.640 9.010 7.010 ;
        RECT 5.100 5.180 9.010 6.640 ;
        RECT -4.610 5.170 9.010 5.180 ;
        RECT -5.280 4.610 9.010 5.170 ;
        RECT -5.280 0.310 18.070 4.610 ;
        RECT -5.280 0.030 9.010 0.310 ;
        RECT 5.100 -1.520 9.010 0.030 ;
        RECT 5.080 -2.290 9.030 -1.520 ;
    END
  END OUTPUT 
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT -7.450 5.090 21.140 6.490 ;
        RECT -6.980 5.080 -6.050 5.090 ;
        RECT -6.730 3.970 -6.560 5.080 ;
    END
    PORT
      LAYER met1 ;
        RECT -7.010 5.840 -4.640 6.470 ;
        RECT 16.330 5.990 20.460 6.390 ;
        RECT 16.330 5.900 20.470 5.990 ;
        RECT -6.980 3.880 -6.030 5.840 ;
        RECT -5.280 5.820 -4.700 5.840 ;
        RECT 19.940 5.000 20.470 5.900 ;
        RECT -6.750 -1.790 -6.030 3.880 ;
      LAYER via ;
        RECT -6.790 5.990 -4.760 6.320 ;
        RECT 16.600 5.990 19.590 6.340 ;
        RECT -6.850 5.130 -6.150 5.750 ;
        RECT 20.030 5.190 20.380 5.950 ;
    END
  END VGND
  PIN VINJ
    ANTENNADIFFAREA 9.088799 ;
    PORT
      LAYER nwell ;
        RECT 7.420 -0.380 19.470 5.560 ;
      LAYER met2 ;
        RECT 18.890 0.190 19.530 3.200 ;
        RECT -7.450 -1.210 21.140 0.190 ;
        RECT 17.990 -1.340 20.620 -1.210 ;
        RECT 17.990 -1.850 20.540 -1.340 ;
        RECT 17.990 -1.920 18.610 -1.850 ;
    END
  END VINJ
  PIN INPUT
    PORT
      LAYER met1 ;
        RECT 0.260 7.990 4.160 8.580 ;
        RECT 0.260 6.640 0.550 7.990 ;
    END
  END INPUT
  OBS
      LAYER li1 ;
        RECT 0.280 6.640 0.530 8.100 ;
        RECT 0.320 6.630 0.490 6.640 ;
        RECT 6.960 6.610 7.210 8.090 ;
        RECT -6.900 5.890 20.480 6.400 ;
        RECT -6.900 3.960 -6.100 5.890 ;
        RECT -5.520 5.440 -5.350 5.520 ;
        RECT 5.720 5.440 5.950 5.530 ;
        RECT -5.520 5.430 5.950 5.440 ;
        RECT -6.900 -0.620 -6.390 3.960 ;
        RECT -5.530 -0.040 5.950 5.430 ;
        RECT -5.600 -0.210 5.950 -0.040 ;
        RECT -5.530 -0.270 -5.340 -0.210 ;
        RECT 5.720 -0.450 5.950 -0.210 ;
        RECT -5.650 -0.620 -3.850 -0.610 ;
        RECT 6.510 -0.620 7.020 5.890 ;
        RECT 7.780 5.000 19.030 5.170 ;
        RECT 7.780 0.130 7.950 5.000 ;
        RECT 8.340 4.670 18.450 4.690 ;
        RECT 8.340 4.630 18.470 4.670 ;
        RECT 8.290 4.460 18.470 4.630 ;
        RECT 8.340 0.440 18.470 4.460 ;
        RECT 18.860 3.240 19.030 5.000 ;
        RECT 8.340 0.360 18.450 0.440 ;
        RECT 7.770 0.060 7.950 0.130 ;
        RECT 18.860 0.060 19.470 3.240 ;
        RECT 7.770 -0.110 19.470 0.060 ;
        RECT 18.930 -0.220 19.470 -0.110 ;
        RECT 19.930 -0.460 20.480 5.890 ;
        RECT 19.920 -0.620 20.480 -0.460 ;
        RECT -6.900 -0.960 20.480 -0.620 ;
        RECT -6.870 -1.130 20.480 -0.960 ;
        RECT -6.870 -1.150 -6.180 -1.130 ;
        RECT -5.670 -1.140 -3.870 -1.130 ;
      LAYER mcon ;
        RECT 0.320 7.580 0.490 7.750 ;
        RECT 0.320 7.220 0.490 7.390 ;
        RECT 0.320 6.850 0.490 7.020 ;
        RECT 7.000 7.900 7.170 8.070 ;
        RECT 7.000 7.540 7.170 7.710 ;
        RECT 7.000 7.180 7.170 7.350 ;
        RECT 7.000 6.820 7.170 6.990 ;
        RECT -6.820 6.230 -4.960 6.240 ;
        RECT -6.820 6.060 -4.950 6.230 ;
        RECT 16.540 6.050 19.700 6.230 ;
        RECT -6.780 3.970 -6.600 5.870 ;
        RECT -6.380 3.960 -6.200 5.870 ;
        RECT -5.190 4.930 5.790 5.100 ;
        RECT -5.190 4.310 5.790 4.480 ;
        RECT -5.180 3.690 5.800 3.860 ;
        RECT -5.160 3.110 5.820 3.280 ;
        RECT -5.150 2.520 5.830 2.690 ;
        RECT -5.150 1.920 5.830 2.090 ;
        RECT -5.200 1.320 5.780 1.490 ;
        RECT -5.190 0.710 5.790 0.880 ;
        RECT -5.200 0.110 5.780 0.280 ;
        RECT 8.540 4.170 17.990 4.340 ;
        RECT 8.530 3.420 17.920 3.590 ;
        RECT 8.560 2.700 17.960 2.870 ;
        RECT 8.570 2.040 17.940 2.210 ;
        RECT 8.560 1.390 18.010 1.560 ;
        RECT 8.570 0.750 17.960 0.920 ;
        RECT 20.110 5.070 20.310 6.000 ;
        RECT 19.040 -0.170 19.390 3.130 ;
      LAYER met1 ;
        RECT 18.840 3.190 19.410 3.200 ;
        RECT 18.840 -0.230 19.460 3.190 ;
        RECT 18.840 -0.240 19.410 -0.230 ;
        RECT 18.010 -1.870 18.570 -1.370 ;
        RECT 18.020 -2.090 18.570 -1.870 ;
      LAYER via ;
        RECT 19.000 -0.100 19.420 3.070 ;
        RECT 18.030 -1.920 18.550 -1.400 ;
  END
END sky130_hilas_VinjDiodeProtect01

MACRO sky130_hilas_TA2Cell_1FG_Strong
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TA2Cell_1FG_Strong ;
  ORIGIN 26.170 -1.350 ;
  SIZE 28.100 BY 6.150 ;
  PIN VTUN
    ANTENNADIFFAREA 5.032200 ;
    PORT
      LAYER nwell ;
        RECT -16.380 6.700 -12.990 7.450 ;
        RECT -16.390 3.130 -12.980 6.700 ;
        RECT -16.380 1.410 -12.990 3.130 ;
      LAYER met1 ;
        RECT -15.410 7.300 -14.990 7.450 ;
        RECT -14.380 7.300 -13.960 7.450 ;
        RECT -15.410 7.160 -13.960 7.300 ;
        RECT -15.410 1.400 -14.990 7.160 ;
        RECT -14.380 1.400 -13.960 7.160 ;
    END
  END VTUN
  PIN PROG
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER met1 ;
        RECT -22.650 4.730 -22.440 7.450 ;
        RECT -22.680 4.220 -22.440 4.730 ;
        RECT -22.650 1.400 -22.440 4.220 ;
    END
  END PROG
  PIN GATE1
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT -10.960 5.060 -8.240 6.710 ;
        RECT -10.960 5.020 -8.250 5.060 ;
        RECT -10.960 3.690 -8.250 3.730 ;
        RECT -10.960 2.040 -8.240 3.690 ;
      LAYER met1 ;
        RECT -10.680 6.240 -10.450 7.450 ;
        RECT -10.680 5.450 -10.420 6.240 ;
        RECT -10.680 3.300 -10.450 5.450 ;
        RECT -10.680 2.510 -10.420 3.300 ;
        RECT -10.680 1.400 -10.450 2.510 ;
    END
  END GATE1
  PIN VIN11
    ANTENNADIFFAREA 0.217200 ;
    PORT
      LAYER met1 ;
        RECT -23.530 7.080 -23.320 7.450 ;
        RECT -23.540 6.790 -23.310 7.080 ;
        RECT -23.530 5.090 -23.320 6.790 ;
        RECT -23.540 4.800 -23.310 5.090 ;
        RECT -23.530 4.660 -23.320 4.800 ;
    END
  END VIN11
  PIN VINJ
    ANTENNADIFFAREA 2.118400 ;
    PORT
      LAYER nwell ;
        RECT -26.170 1.350 -22.860 7.500 ;
        RECT -6.510 7.450 -3.200 7.500 ;
        RECT -6.510 7.440 -1.860 7.450 ;
        RECT -6.510 1.400 -1.350 7.440 ;
        RECT -6.510 1.350 -3.200 1.400 ;
      LAYER met2 ;
        RECT -25.970 7.310 -25.650 7.430 ;
        RECT -3.700 7.310 -3.380 7.430 ;
        RECT -25.970 7.130 -3.380 7.310 ;
        RECT -4.590 4.590 -4.270 4.850 ;
        RECT -4.550 4.570 -3.370 4.590 ;
        RECT -4.550 4.310 -3.330 4.570 ;
        RECT -4.550 4.250 -3.370 4.310 ;
        RECT -4.590 4.240 -3.370 4.250 ;
        RECT -4.590 3.990 -4.270 4.240 ;
    END
    PORT
      LAYER met1 ;
        RECT -3.720 7.430 -3.440 7.450 ;
        RECT -3.720 7.130 -3.380 7.430 ;
        RECT -3.720 6.800 -3.440 7.130 ;
        RECT -3.830 6.200 -3.440 6.800 ;
        RECT -3.720 4.600 -3.440 6.200 ;
        RECT -3.720 4.280 -3.360 4.600 ;
        RECT -3.720 2.650 -3.440 4.280 ;
        RECT -3.830 2.050 -3.440 2.650 ;
        RECT -3.720 1.400 -3.440 2.050 ;
      LAYER via ;
        RECT -3.670 7.150 -3.410 7.410 ;
        RECT -3.620 4.310 -3.360 4.570 ;
    END
  END VINJ
  PIN VIN22
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -1.960 7.430 -1.650 7.440 ;
        RECT -2.530 7.420 -1.650 7.430 ;
        RECT -2.600 7.180 -1.650 7.420 ;
        RECT -1.960 7.110 -1.650 7.180 ;
    END
  END VIN22
  PIN VIN21
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -2.200 4.750 -1.890 4.790 ;
        RECT -2.520 4.740 -1.860 4.750 ;
        RECT -2.520 4.510 -1.420 4.740 ;
        RECT -2.200 4.460 -1.890 4.510 ;
    END
  END VIN21
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.650 1.400 1.930 7.450 ;
      LAYER met1 ;
        RECT 0.630 7.300 0.910 7.450 ;
        RECT 0.640 5.870 0.910 7.300 ;
        RECT 0.640 5.580 0.920 5.870 ;
        RECT 0.640 3.280 0.910 5.580 ;
        RECT 0.640 2.990 0.920 3.280 ;
        RECT 0.640 1.400 0.910 2.990 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT -1.560 1.750 -1.240 1.900 ;
        RECT -17.750 1.600 -1.240 1.750 ;
        RECT -17.750 1.450 -17.430 1.600 ;
        RECT -11.950 1.450 -11.630 1.600 ;
    END
    PORT
      LAYER met1 ;
        RECT -1.560 1.600 -1.240 1.900 ;
        RECT -0.030 1.600 0.310 7.450 ;
        RECT -1.560 1.570 -1.130 1.600 ;
        RECT -0.530 1.570 0.310 1.600 ;
        RECT -1.560 1.540 0.310 1.570 ;
        RECT -1.410 1.490 0.310 1.540 ;
        RECT -1.380 1.460 0.310 1.490 ;
        RECT -1.350 1.440 0.310 1.460 ;
        RECT -1.280 1.430 -0.320 1.440 ;
        RECT -0.030 1.400 0.310 1.440 ;
      LAYER via ;
        RECT -1.530 1.620 -1.270 1.880 ;
    END
  END VGND
  PIN OUTPUT2
    ANTENNADIFFAREA 0.308800 ;
    PORT
      LAYER met2 ;
        RECT -0.990 4.140 -0.680 4.190 ;
        RECT 1.300 4.140 1.610 4.270 ;
        RECT -0.990 3.920 1.930 4.140 ;
        RECT -0.990 3.860 -0.680 3.920 ;
    END
  END OUTPUT2
  PIN OUTPUT1
    ANTENNADIFFAREA 0.308800 ;
    PORT
      LAYER met2 ;
        RECT -0.990 4.970 -0.680 5.030 ;
        RECT 1.310 4.970 1.620 4.990 ;
        RECT -0.990 4.740 1.930 4.970 ;
        RECT -0.990 4.700 -0.680 4.740 ;
        RECT 1.310 4.660 1.620 4.740 ;
    END
  END OUTPUT1
  PIN GATESEL1
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT -25.400 5.990 -25.210 7.450 ;
        RECT -25.430 5.960 -25.210 5.990 ;
        RECT -25.440 5.690 -25.190 5.960 ;
        RECT -25.440 5.680 -25.200 5.690 ;
        RECT -25.430 5.440 -25.200 5.680 ;
        RECT -25.400 3.410 -25.240 5.440 ;
        RECT -25.430 3.170 -25.200 3.410 ;
        RECT -25.440 3.160 -25.200 3.170 ;
        RECT -25.440 2.890 -25.190 3.160 ;
        RECT -25.430 2.860 -25.210 2.890 ;
        RECT -25.400 1.400 -25.210 2.860 ;
    END
  END GATESEL1
  PIN GATESEL2
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT -4.160 5.990 -3.970 7.450 ;
        RECT -4.160 5.960 -3.940 5.990 ;
        RECT -4.180 5.690 -3.930 5.960 ;
        RECT -4.170 5.680 -3.930 5.690 ;
        RECT -4.170 5.440 -3.940 5.680 ;
        RECT -4.130 3.410 -3.970 5.440 ;
        RECT -4.170 3.170 -3.940 3.410 ;
        RECT -4.170 3.160 -3.930 3.170 ;
        RECT -4.180 2.890 -3.930 3.160 ;
        RECT -4.160 2.860 -3.940 2.890 ;
        RECT -4.160 1.400 -3.970 2.860 ;
    END
  END GATESEL2
  PIN DRAIN1
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER met2 ;
        RECT -23.760 6.960 -23.440 6.970 ;
        RECT -24.000 6.950 -23.440 6.960 ;
        RECT -5.680 6.950 -5.370 6.960 ;
        RECT -26.170 6.770 -3.200 6.950 ;
        RECT -24.000 6.630 -23.690 6.770 ;
        RECT -5.680 6.630 -5.370 6.770 ;
    END
  END DRAIN1
  PIN DRAIN2
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER met2 ;
        RECT -24.000 2.080 -23.690 2.220 ;
        RECT -26.170 2.070 -23.690 2.080 ;
        RECT -5.680 2.080 -5.370 2.220 ;
        RECT -5.680 2.070 -3.200 2.080 ;
        RECT -26.170 1.920 -3.200 2.070 ;
        RECT -26.170 1.900 -23.690 1.920 ;
        RECT -24.000 1.890 -23.690 1.900 ;
        RECT -5.680 1.900 -3.200 1.920 ;
        RECT -5.680 1.890 -5.370 1.900 ;
    END
  END DRAIN2
  PIN VIN12
    ANTENNADIFFAREA 0.217200 ;
    PORT
      LAYER met1 ;
        RECT -23.510 4.020 -23.320 4.150 ;
        RECT -23.530 3.730 -23.300 4.020 ;
        RECT -23.510 2.110 -23.320 3.730 ;
        RECT -23.510 1.900 -23.280 2.110 ;
        RECT -23.520 1.820 -23.280 1.900 ;
        RECT -23.520 1.400 -23.290 1.820 ;
    END
  END VIN12
  PIN GATE2
    ANTENNADIFFAREA 0.434600 ;
    PORT
      LAYER met1 ;
        RECT -23.060 6.520 -22.870 7.450 ;
        RECT -23.070 6.230 -22.840 6.520 ;
        RECT -23.060 4.200 -22.870 6.230 ;
        RECT -23.070 3.910 -22.840 4.200 ;
        RECT -23.060 2.620 -22.870 3.910 ;
        RECT -23.080 2.330 -22.850 2.620 ;
        RECT -23.060 1.400 -22.870 2.330 ;
    END
  END GATE2
  PIN RUN
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER met1 ;
        RECT -21.570 2.920 -21.390 7.450 ;
        RECT -21.630 2.580 -21.340 2.920 ;
        RECT -21.570 1.400 -21.390 2.580 ;
    END
  END RUN
  OBS
      LAYER nwell ;
        RECT -21.130 5.060 -18.410 6.710 ;
        RECT -21.130 5.020 -18.420 5.060 ;
        RECT -21.130 3.690 -18.420 3.730 ;
        RECT -21.130 2.040 -18.410 3.690 ;
      LAYER li1 ;
        RECT -2.220 7.400 -2.050 7.450 ;
        RECT -2.220 7.140 -1.660 7.400 ;
        RECT -0.750 7.150 -0.550 7.190 ;
        RECT -2.220 7.120 -2.050 7.140 ;
        RECT -25.770 6.770 -25.570 7.120 ;
        RECT -24.290 6.870 -23.760 7.040 ;
        RECT -23.520 7.020 -23.330 7.050 ;
        RECT -23.520 6.850 -22.460 7.020 ;
        RECT -5.610 6.870 -5.080 7.040 ;
        RECT -23.520 6.820 -23.330 6.850 ;
        RECT -25.780 6.740 -25.570 6.770 ;
        RECT -25.780 6.160 -25.560 6.740 ;
        RECT -25.780 6.150 -25.570 6.160 ;
        RECT -25.400 5.980 -25.210 5.990 ;
        RECT -25.410 5.690 -25.210 5.980 ;
        RECT -25.470 5.360 -25.200 5.690 ;
        RECT -25.010 4.880 -24.840 6.490 ;
        RECT -24.180 5.390 -24.010 6.480 ;
        RECT -23.050 6.460 -22.860 6.490 ;
        RECT -23.590 6.290 -22.860 6.460 ;
        RECT -22.630 6.460 -22.460 6.850 ;
        RECT -3.800 6.770 -3.600 7.120 ;
        RECT -3.800 6.740 -3.590 6.770 ;
        RECT -22.630 6.290 -21.890 6.460 ;
        RECT -23.050 6.260 -22.860 6.290 ;
        RECT -20.830 5.670 -20.600 6.190 ;
        RECT -23.590 5.500 -20.600 5.670 ;
        RECT -24.410 5.350 -24.010 5.390 ;
        RECT -24.420 5.160 -24.010 5.350 ;
        RECT -15.630 5.310 -15.080 5.740 ;
        RECT -14.290 5.310 -13.740 5.740 ;
        RECT -10.660 5.500 -10.430 6.190 ;
        RECT -5.360 5.960 -5.190 6.480 ;
        RECT -5.520 5.700 -5.190 5.960 ;
        RECT -24.410 5.130 -24.010 5.160 ;
        RECT -25.020 4.690 -24.840 4.880 ;
        RECT -24.180 4.790 -24.010 5.130 ;
        RECT -23.520 4.880 -23.330 5.060 ;
        RECT -23.590 4.710 -23.240 4.880 ;
        RECT -22.670 4.300 -22.460 4.730 ;
        RECT -22.240 4.710 -21.900 4.880 ;
        RECT -22.650 4.280 -22.480 4.300 ;
        RECT -25.020 3.970 -24.840 4.160 ;
        RECT -25.470 3.160 -25.200 3.490 ;
        RECT -25.410 2.870 -25.210 3.160 ;
        RECT -25.400 2.860 -25.210 2.870 ;
        RECT -25.780 2.690 -25.570 2.700 ;
        RECT -25.780 2.110 -25.560 2.690 ;
        RECT -25.010 2.360 -24.840 3.970 ;
        RECT -24.180 3.700 -24.010 4.060 ;
        RECT -23.590 3.970 -23.240 4.140 ;
        RECT -23.050 4.120 -22.860 4.170 ;
        RECT -22.150 4.140 -21.980 4.710 ;
        RECT -17.870 4.480 -17.680 4.880 ;
        RECT -11.690 4.480 -11.500 4.880 ;
        RECT -5.360 4.790 -5.190 5.700 ;
        RECT -4.530 4.880 -4.360 6.490 ;
        RECT -3.810 6.160 -3.590 6.740 ;
        RECT -3.800 6.150 -3.590 6.160 ;
        RECT -2.800 6.040 -2.620 6.970 ;
        RECT -0.980 6.890 -0.550 7.150 ;
        RECT -2.070 6.710 -1.740 6.880 ;
        RECT -0.750 6.860 -0.550 6.890 ;
        RECT -1.990 6.570 -1.740 6.710 ;
        RECT -1.990 6.310 -1.510 6.570 ;
        RECT -1.160 6.500 -0.990 6.540 ;
        RECT -0.750 6.500 -0.550 6.530 ;
        RECT -2.920 6.010 -2.600 6.040 ;
        RECT -4.160 5.980 -3.970 5.990 ;
        RECT -4.160 5.690 -3.960 5.980 ;
        RECT -2.920 5.820 -2.590 6.010 ;
        RECT -2.920 5.780 -2.600 5.820 ;
        RECT -4.170 5.360 -3.880 5.690 ;
        RECT -4.530 4.690 -4.350 4.880 ;
        RECT -17.870 4.470 -17.490 4.480 ;
        RECT -21.230 4.290 -17.490 4.470 ;
        RECT -17.870 4.250 -17.490 4.290 ;
        RECT -11.880 4.470 -11.500 4.480 ;
        RECT -11.880 4.290 -8.140 4.470 ;
        RECT -11.880 4.250 -11.500 4.290 ;
        RECT -23.050 4.110 -22.820 4.120 ;
        RECT -22.240 4.110 -21.900 4.140 ;
        RECT -23.050 3.970 -21.900 4.110 ;
        RECT -23.510 3.760 -23.320 3.970 ;
        RECT -23.050 3.940 -22.070 3.970 ;
        RECT -22.910 3.910 -22.070 3.940 ;
        RECT -17.870 3.870 -17.680 4.250 ;
        RECT -24.420 3.660 -24.010 3.700 ;
        RECT -24.430 3.470 -24.010 3.660 ;
        RECT -15.630 3.580 -15.080 4.010 ;
        RECT -14.290 3.580 -13.740 4.010 ;
        RECT -11.690 3.870 -11.500 4.250 ;
        RECT -24.420 3.440 -24.010 3.470 ;
        RECT -24.180 2.370 -24.010 3.440 ;
        RECT -23.590 3.250 -20.660 3.350 ;
        RECT -23.590 3.180 -20.600 3.250 ;
        RECT -21.570 2.860 -21.400 2.920 ;
        RECT -21.590 2.650 -21.380 2.860 ;
        RECT -23.060 2.560 -22.870 2.590 ;
        RECT -21.570 2.580 -21.400 2.650 ;
        RECT -20.830 2.560 -20.600 3.180 ;
        RECT -10.660 2.560 -10.430 3.290 ;
        RECT -5.360 3.200 -5.190 4.060 ;
        RECT -5.520 2.940 -5.190 3.200 ;
        RECT -23.590 2.390 -22.870 2.560 ;
        RECT -23.060 2.360 -22.870 2.390 ;
        RECT -22.700 2.390 -21.890 2.560 ;
        RECT -25.780 2.080 -25.570 2.110 ;
        RECT -25.770 1.730 -25.570 2.080 ;
        RECT -23.490 2.050 -23.300 2.080 ;
        RECT -22.700 2.050 -22.510 2.390 ;
        RECT -5.360 2.370 -5.190 2.940 ;
        RECT -4.530 3.970 -4.350 4.160 ;
        RECT -4.530 2.360 -4.360 3.970 ;
        RECT -4.170 3.160 -3.880 3.490 ;
        RECT -4.160 2.870 -3.960 3.160 ;
        RECT -4.160 2.860 -3.970 2.870 ;
        RECT -3.800 2.690 -3.590 2.700 ;
        RECT -3.810 2.110 -3.590 2.690 ;
        RECT -24.290 1.810 -23.760 1.980 ;
        RECT -23.490 1.870 -22.510 2.050 ;
        RECT -3.800 2.080 -3.590 2.110 ;
        RECT -23.490 1.850 -23.300 1.870 ;
        RECT -5.610 1.810 -5.080 1.980 ;
        RECT -3.800 1.730 -3.600 2.080 ;
        RECT -2.800 1.870 -2.620 5.780 ;
        RECT -1.990 4.930 -1.820 6.310 ;
        RECT -1.160 6.240 -0.550 6.500 ;
        RECT -1.160 6.210 -0.990 6.240 ;
        RECT -0.750 6.200 -0.550 6.240 ;
        RECT -0.160 6.200 0.390 7.190 ;
        RECT 1.210 7.040 1.840 7.210 ;
        RECT 1.210 6.940 1.600 7.040 ;
        RECT 1.210 6.910 1.590 6.940 ;
        RECT 1.210 6.760 1.570 6.910 ;
        RECT 0.860 6.590 1.570 6.760 ;
        RECT 0.860 5.840 1.560 6.150 ;
        RECT -1.160 5.650 -0.990 5.680 ;
        RECT -0.750 5.650 -0.550 5.690 ;
        RECT -1.160 5.390 -0.550 5.650 ;
        RECT -1.160 5.350 -0.990 5.390 ;
        RECT -0.750 5.360 -0.550 5.390 ;
        RECT -0.750 5.000 -0.550 5.030 ;
        RECT -2.190 4.730 -1.870 4.760 ;
        RECT -0.980 4.740 -0.550 5.000 ;
        RECT -2.190 4.540 -1.860 4.730 ;
        RECT -0.750 4.700 -0.550 4.740 ;
        RECT -0.160 4.700 0.390 5.690 ;
        RECT 0.710 5.610 1.560 5.840 ;
        RECT 0.860 5.270 1.560 5.610 ;
        RECT 1.320 4.910 1.640 4.950 ;
        RECT 1.320 4.850 1.650 4.910 ;
        RECT 0.850 4.720 1.650 4.850 ;
        RECT 0.850 4.690 1.640 4.720 ;
        RECT 0.850 4.670 1.550 4.690 ;
        RECT -2.190 4.500 -1.870 4.540 ;
        RECT -2.190 4.420 -2.020 4.500 ;
        RECT -2.240 4.250 -2.020 4.420 ;
        RECT -2.240 4.090 -2.070 4.250 ;
        RECT 1.310 4.190 1.630 4.230 ;
        RECT -0.750 4.150 -0.550 4.190 ;
        RECT -1.710 3.830 -1.520 3.950 ;
        RECT -0.980 3.890 -0.550 4.150 ;
        RECT -0.750 3.860 -0.550 3.890 ;
        RECT -2.070 3.720 -1.520 3.830 ;
        RECT -2.070 3.660 -1.530 3.720 ;
        RECT -1.990 1.880 -1.820 3.660 ;
        RECT -1.160 3.500 -0.990 3.540 ;
        RECT -0.750 3.500 -0.550 3.530 ;
        RECT -1.160 3.240 -0.550 3.500 ;
        RECT -1.160 3.210 -0.990 3.240 ;
        RECT -0.750 3.200 -0.550 3.240 ;
        RECT -0.160 3.200 0.390 4.190 ;
        RECT 0.850 4.010 1.640 4.190 ;
        RECT 1.310 4.000 1.640 4.010 ;
        RECT 1.310 3.970 1.630 4.000 ;
        RECT 0.860 3.250 1.560 3.590 ;
        RECT 0.710 3.020 1.560 3.250 ;
        RECT 0.860 2.710 1.560 3.020 ;
        RECT -1.160 2.650 -0.990 2.680 ;
        RECT -0.750 2.650 -0.550 2.690 ;
        RECT -1.160 2.390 -0.550 2.650 ;
        RECT -1.160 2.350 -0.990 2.390 ;
        RECT -0.750 2.360 -0.550 2.390 ;
        RECT -0.750 2.000 -0.550 2.030 ;
        RECT -0.980 1.740 -0.550 2.000 ;
        RECT -0.750 1.700 -0.550 1.740 ;
        RECT -0.160 1.700 0.390 2.690 ;
        RECT 0.860 2.100 1.570 2.270 ;
        RECT 1.210 1.820 1.570 2.100 ;
        RECT 1.210 1.650 1.840 1.820 ;
      LAYER mcon ;
        RECT -1.890 7.180 -1.720 7.350 ;
        RECT -23.940 6.870 -23.760 7.040 ;
        RECT -23.510 6.850 -23.340 7.020 ;
        RECT -25.750 6.570 -25.580 6.740 ;
        RECT -25.400 5.730 -25.220 5.920 ;
        RECT -23.040 6.290 -22.870 6.460 ;
        RECT -3.790 6.570 -3.620 6.740 ;
        RECT -20.800 5.990 -20.630 6.160 ;
        RECT -10.630 5.990 -10.460 6.160 ;
        RECT -20.800 5.540 -20.630 5.710 ;
        RECT -24.320 5.170 -24.150 5.340 ;
        RECT -15.350 5.390 -15.080 5.660 ;
        RECT -14.290 5.390 -14.020 5.660 ;
        RECT -10.630 5.540 -10.460 5.710 ;
        RECT -5.460 5.740 -5.290 5.910 ;
        RECT -23.510 4.860 -23.340 5.030 ;
        RECT -0.920 6.930 -0.750 7.100 ;
        RECT 0.060 6.610 0.230 6.780 ;
        RECT 1.330 6.950 1.500 7.120 ;
        RECT -1.740 6.350 -1.570 6.520 ;
        RECT -4.150 5.730 -3.970 5.920 ;
        RECT -2.860 5.830 -2.690 6.000 ;
        RECT -17.670 4.280 -17.500 4.450 ;
        RECT -11.870 4.280 -11.700 4.450 ;
        RECT -25.400 2.930 -25.220 3.120 ;
        RECT -23.040 3.970 -22.870 4.140 ;
        RECT -23.500 3.790 -23.330 3.960 ;
        RECT -24.330 3.480 -24.160 3.650 ;
        RECT -15.350 3.660 -15.080 3.930 ;
        RECT -14.290 3.660 -14.020 3.930 ;
        RECT -20.800 3.040 -20.630 3.210 ;
        RECT -20.800 2.590 -20.630 2.760 ;
        RECT -10.630 3.040 -10.460 3.210 ;
        RECT -5.460 2.980 -5.290 3.150 ;
        RECT -10.630 2.590 -10.460 2.760 ;
        RECT -23.050 2.390 -22.880 2.560 ;
        RECT -25.750 2.110 -25.580 2.280 ;
        RECT -4.150 2.930 -3.970 3.120 ;
        RECT -3.790 2.110 -3.620 2.280 ;
        RECT -23.940 1.810 -23.760 1.980 ;
        RECT -23.480 1.880 -23.310 2.050 ;
        RECT -0.970 6.280 -0.800 6.450 ;
        RECT -0.970 5.440 -0.800 5.610 ;
        RECT 0.720 5.640 0.890 5.810 ;
        RECT 0.060 5.110 0.230 5.280 ;
        RECT -0.920 4.790 -0.750 4.960 ;
        RECT -2.130 4.550 -1.960 4.720 ;
        RECT 1.380 4.730 1.550 4.900 ;
        RECT -1.700 3.750 -1.530 3.920 ;
        RECT -0.920 3.930 -0.750 4.100 ;
        RECT 1.370 4.010 1.540 4.180 ;
        RECT 0.060 3.610 0.230 3.780 ;
        RECT -0.970 3.280 -0.800 3.450 ;
        RECT 0.720 3.050 0.890 3.220 ;
        RECT -0.970 2.440 -0.800 2.610 ;
        RECT 0.060 2.110 0.230 2.280 ;
        RECT -0.920 1.790 -0.750 1.960 ;
        RECT 1.290 1.760 1.460 1.930 ;
      LAYER met1 ;
        RECT -25.810 7.430 -25.650 7.450 ;
        RECT -25.970 7.130 -25.650 7.430 ;
        RECT -25.810 6.800 -25.650 7.130 ;
        RECT -25.810 6.250 -25.540 6.800 ;
        RECT -24.000 6.630 -23.690 7.070 ;
        RECT -25.820 6.200 -25.540 6.250 ;
        RECT -25.820 6.110 -25.650 6.200 ;
        RECT -25.810 2.740 -25.650 6.110 ;
        RECT -20.850 5.450 -20.590 6.240 ;
        RECT -24.400 5.100 -24.080 5.420 ;
        RECT -25.050 4.590 -24.810 5.010 ;
        RECT -25.080 4.270 -24.810 4.590 ;
        RECT -25.050 3.840 -24.810 4.270 ;
        RECT -24.410 3.410 -24.090 3.730 ;
        RECT -25.820 2.650 -25.650 2.740 ;
        RECT -25.820 2.600 -25.540 2.650 ;
        RECT -25.810 2.050 -25.540 2.600 ;
        RECT -20.850 2.510 -20.590 3.300 ;
        RECT -25.810 1.400 -25.650 2.050 ;
        RECT -24.000 1.780 -23.690 2.220 ;
        RECT -17.700 1.750 -17.470 7.450 ;
        RECT -11.900 1.750 -11.670 7.450 ;
        RECT -1.970 7.110 -1.650 7.430 ;
        RECT -5.680 6.630 -5.370 7.070 ;
        RECT -0.990 6.860 -0.670 7.180 ;
        RECT 1.260 6.880 1.580 7.200 ;
        RECT -1.820 6.280 -1.500 6.600 ;
        RECT -1.040 6.210 -0.720 6.530 ;
        RECT -5.530 5.670 -5.210 5.990 ;
        RECT -2.930 5.750 -2.610 6.070 ;
        RECT -1.710 5.590 -1.500 5.700 ;
        RECT -1.730 5.270 -1.470 5.590 ;
        RECT -1.040 5.360 -0.720 5.680 ;
        RECT -4.560 4.880 -4.320 5.010 ;
        RECT -4.560 4.560 -4.300 4.880 ;
        RECT -2.200 4.470 -1.880 4.790 ;
        RECT -4.560 3.960 -4.300 4.280 ;
        RECT -1.710 3.980 -1.500 5.270 ;
        RECT -0.990 4.710 -0.670 5.030 ;
        RECT 1.310 4.660 1.630 4.980 ;
        RECT -4.560 3.840 -4.320 3.960 ;
        RECT -1.730 3.690 -1.500 3.980 ;
        RECT -0.990 3.860 -0.670 4.180 ;
        RECT 1.300 3.940 1.620 4.260 ;
        RECT -5.530 2.910 -5.210 3.230 ;
        RECT -1.040 3.210 -0.720 3.530 ;
        RECT -1.040 2.360 -0.720 2.680 ;
        RECT -5.680 1.780 -5.370 2.220 ;
        RECT -17.750 1.450 -17.430 1.750 ;
        RECT -11.950 1.450 -11.630 1.750 ;
        RECT -0.990 1.710 -0.670 2.030 ;
        RECT 1.220 1.690 1.540 2.010 ;
        RECT -17.700 1.400 -17.470 1.450 ;
        RECT -11.900 1.400 -11.670 1.450 ;
      LAYER via ;
        RECT -25.940 7.150 -25.680 7.410 ;
        RECT -23.980 6.660 -23.720 6.920 ;
        RECT -24.370 5.130 -24.110 5.390 ;
        RECT -25.080 4.300 -24.820 4.560 ;
        RECT -24.380 3.440 -24.120 3.700 ;
        RECT -23.980 1.930 -23.720 2.190 ;
        RECT -1.940 7.140 -1.680 7.400 ;
        RECT -5.650 6.660 -5.390 6.920 ;
        RECT -0.960 6.890 -0.700 7.150 ;
        RECT 1.290 6.910 1.550 7.170 ;
        RECT -1.790 6.310 -1.530 6.570 ;
        RECT -1.010 6.240 -0.750 6.500 ;
        RECT -5.500 5.700 -5.240 5.960 ;
        RECT -2.900 5.780 -2.640 6.040 ;
        RECT -1.730 5.300 -1.470 5.560 ;
        RECT -1.010 5.390 -0.750 5.650 ;
        RECT -4.560 4.590 -4.300 4.850 ;
        RECT -2.170 4.500 -1.910 4.760 ;
        RECT -4.560 3.990 -4.300 4.250 ;
        RECT -0.960 4.740 -0.700 5.000 ;
        RECT 1.340 4.690 1.600 4.950 ;
        RECT -0.960 3.890 -0.700 4.150 ;
        RECT 1.330 3.970 1.590 4.230 ;
        RECT -1.010 3.240 -0.750 3.500 ;
        RECT -5.500 2.940 -5.240 3.200 ;
        RECT -1.010 2.390 -0.750 2.650 ;
        RECT -5.650 1.930 -5.390 2.190 ;
        RECT -17.720 1.470 -17.460 1.730 ;
        RECT -11.920 1.470 -11.660 1.730 ;
        RECT -0.960 1.740 -0.700 2.000 ;
        RECT 1.250 1.720 1.510 1.980 ;
      LAYER met2 ;
        RECT -0.990 7.110 -0.680 7.190 ;
        RECT 1.260 7.110 1.570 7.210 ;
        RECT -0.990 6.880 1.570 7.110 ;
        RECT -0.990 6.860 -0.680 6.880 ;
        RECT -1.810 6.570 -1.500 6.610 ;
        RECT -1.990 6.460 -1.270 6.570 ;
        RECT -1.040 6.460 -0.730 6.540 ;
        RECT -1.990 6.320 -0.730 6.460 ;
        RECT -1.810 6.280 -0.730 6.320 ;
        RECT -1.540 6.250 -0.730 6.280 ;
        RECT -1.540 6.210 -1.270 6.250 ;
        RECT -1.040 6.210 -0.730 6.250 ;
        RECT -5.530 5.930 -5.220 6.000 ;
        RECT -2.930 5.930 -2.620 6.070 ;
        RECT -5.530 5.740 -2.620 5.930 ;
        RECT -5.530 5.710 -2.930 5.740 ;
        RECT -5.530 5.670 -5.220 5.710 ;
        RECT -1.470 5.640 -1.270 5.650 ;
        RECT -1.040 5.640 -0.730 5.680 ;
        RECT -1.470 5.560 -0.730 5.640 ;
        RECT -1.760 5.540 -0.730 5.560 ;
        RECT -1.810 5.430 -0.730 5.540 ;
        RECT -24.390 5.410 -24.080 5.430 ;
        RECT -14.660 5.410 -6.670 5.420 ;
        RECT -24.390 5.220 -6.670 5.410 ;
        RECT -1.810 5.300 -1.250 5.430 ;
        RECT -1.040 5.350 -0.730 5.430 ;
        RECT -1.810 5.290 -1.340 5.300 ;
        RECT -24.390 5.100 -24.080 5.220 ;
        RECT -25.110 4.530 -24.790 4.560 ;
        RECT -8.070 4.540 -7.850 4.550 ;
        RECT -14.650 4.530 -7.820 4.540 ;
        RECT -25.110 4.300 -7.820 4.530 ;
        RECT -6.890 4.500 -6.670 5.220 ;
        RECT -14.650 4.290 -7.820 4.300 ;
        RECT -24.400 3.550 -24.090 3.740 ;
        RECT -14.650 3.550 -11.140 3.560 ;
        RECT -24.400 3.410 -11.140 3.550 ;
        RECT -24.370 3.370 -11.140 3.410 ;
        RECT -24.370 3.360 -14.650 3.370 ;
        RECT -11.370 2.770 -11.140 3.370 ;
        RECT -8.110 3.120 -7.820 4.290 ;
        RECT -6.920 4.460 -6.670 4.500 ;
        RECT -6.920 3.820 -6.660 4.460 ;
        RECT -6.920 3.610 -2.790 3.820 ;
        RECT -3.000 3.470 -2.790 3.610 ;
        RECT -1.040 3.470 -0.730 3.540 ;
        RECT -3.000 3.260 -0.730 3.470 ;
        RECT -1.340 3.250 -0.730 3.260 ;
        RECT -5.530 3.170 -5.220 3.240 ;
        RECT -1.040 3.210 -0.730 3.250 ;
        RECT -5.530 3.120 -3.200 3.170 ;
        RECT -8.110 2.960 -3.200 3.120 ;
        RECT -8.110 2.900 -5.220 2.960 ;
        RECT -8.110 2.890 -7.820 2.900 ;
        RECT -11.370 2.620 -11.150 2.770 ;
        RECT -1.040 2.670 -0.730 2.680 ;
        RECT -7.000 2.620 -0.730 2.670 ;
        RECT -11.370 2.460 -0.730 2.620 ;
        RECT -11.370 2.400 -6.610 2.460 ;
        RECT -1.340 2.430 -0.730 2.460 ;
        RECT -1.040 2.350 -0.730 2.430 ;
        RECT -0.990 1.980 -0.680 2.030 ;
        RECT 1.220 1.980 1.530 2.020 ;
        RECT -0.990 1.750 1.720 1.980 ;
        RECT -0.990 1.700 -0.680 1.750 ;
        RECT 1.220 1.690 1.530 1.750 ;
  END
END sky130_hilas_TA2Cell_1FG_Strong

MACRO sky130_hilas_pFETmed
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pFETmed ;
  ORIGIN -1.470 0.220 ;
  SIZE 1.190 BY 2.870 ;
  OBS
      LAYER nwell ;
        RECT 1.470 -0.220 2.660 2.650 ;
      LAYER li1 ;
        RECT 1.710 -0.070 1.880 2.420 ;
        RECT 2.260 -0.080 2.430 2.420 ;
  END
END sky130_hilas_pFETmed

MACRO sky130_hilas_capacitorSize02
  CLASS BLOCK ;
  FOREIGN sky130_hilas_capacitorSize02 ;
  ORIGIN -14.140 0.480 ;
  SIZE 7.970 BY 5.830 ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 21.370 2.140 22.030 2.800 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 14.250 2.720 14.910 2.780 ;
        RECT 15.300 2.720 16.310 2.730 ;
        RECT 14.250 2.220 17.940 2.720 ;
        RECT 14.250 2.210 15.660 2.220 ;
        RECT 14.250 2.120 14.910 2.210 ;
        RECT 17.300 1.100 17.930 2.220 ;
        RECT 17.300 1.090 19.450 1.100 ;
        RECT 15.980 0.790 19.450 1.090 ;
        RECT 15.980 0.620 18.990 0.790 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 14.140 4.800 22.110 4.980 ;
        RECT 14.140 4.370 22.110 4.550 ;
        RECT 14.170 3.370 22.110 3.550 ;
        RECT 14.170 2.940 22.110 3.120 ;
        RECT 14.380 2.600 14.750 2.660 ;
        RECT 14.160 2.320 14.750 2.600 ;
        RECT 14.380 2.260 14.750 2.320 ;
        RECT 21.500 2.620 21.870 2.680 ;
        RECT 21.500 2.340 22.110 2.620 ;
        RECT 21.500 2.280 21.870 2.340 ;
        RECT 14.170 1.790 22.110 1.960 ;
        RECT 14.170 1.370 22.110 1.540 ;
        RECT 14.170 0.390 22.110 0.560 ;
        RECT 14.170 -0.050 22.110 0.120 ;
      LAYER via2 ;
        RECT 14.430 2.320 14.710 2.600 ;
        RECT 21.550 2.340 21.830 2.620 ;
      LAYER met3 ;
        RECT 15.600 5.320 17.910 5.350 ;
        RECT 15.600 2.830 19.830 5.320 ;
        RECT 14.160 2.060 14.950 2.810 ;
        RECT 15.600 2.080 22.070 2.830 ;
        RECT 15.600 -0.460 19.830 2.080 ;
        RECT 17.880 -0.480 19.830 -0.460 ;
      LAYER via3 ;
        RECT 14.350 2.210 14.780 2.690 ;
        RECT 21.470 2.230 21.900 2.710 ;
  END
END sky130_hilas_capacitorSize02

MACRO sky130_hilas_swc4x2cellOverlap
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc4x2cellOverlap ;
  ORIGIN 10.010 -7.230 ;
  SIZE 17.980 BY 6.160 ;
  PIN VERT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met1 ;
        RECT -8.840 12.650 -8.680 13.380 ;
        RECT -8.880 12.630 -8.680 12.650 ;
        RECT -8.890 12.390 -8.660 12.630 ;
        RECT -8.890 12.340 -8.680 12.390 ;
        RECT -8.840 11.280 -8.680 12.340 ;
        RECT -8.890 11.230 -8.680 11.280 ;
        RECT -8.890 10.990 -8.660 11.230 ;
        RECT -8.880 10.970 -8.680 10.990 ;
        RECT -8.840 9.640 -8.680 10.970 ;
        RECT -8.880 9.620 -8.680 9.640 ;
        RECT -8.890 9.380 -8.660 9.620 ;
        RECT -8.890 9.330 -8.680 9.380 ;
        RECT -8.840 8.280 -8.680 9.330 ;
        RECT -8.890 8.230 -8.680 8.280 ;
        RECT -8.890 7.990 -8.660 8.230 ;
        RECT -8.880 7.970 -8.680 7.990 ;
        RECT -8.840 7.240 -8.680 7.970 ;
    END
  END VERT1
  PIN HORIZ1
    USE ANALOG ;
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT -7.850 12.400 -7.540 12.420 ;
        RECT 5.490 12.400 5.800 12.420 ;
        RECT -10.010 12.220 7.970 12.400 ;
        RECT -7.850 12.090 -7.540 12.220 ;
        RECT 5.490 12.090 5.800 12.220 ;
    END
  END HORIZ1
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT -7.850 12.830 -7.540 12.970 ;
        RECT 5.490 12.830 5.800 12.970 ;
        RECT -10.010 12.650 7.960 12.830 ;
        RECT -7.850 12.640 -7.540 12.650 ;
        RECT 5.490 12.640 5.800 12.650 ;
    END
  END DRAIN1
  PIN HORIZ2
    USE ANALOG ;
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT -7.850 11.400 -7.540 11.530 ;
        RECT 5.490 11.400 5.800 11.530 ;
        RECT -10.010 11.220 7.970 11.400 ;
        RECT -7.850 11.200 -7.540 11.220 ;
        RECT 5.490 11.200 5.800 11.220 ;
    END
  END HORIZ2
  PIN DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT -7.850 10.970 -7.540 10.980 ;
        RECT 5.490 10.970 5.800 10.980 ;
        RECT -10.010 10.790 7.970 10.970 ;
        RECT -7.850 10.650 -7.540 10.790 ;
        RECT 5.490 10.650 5.800 10.790 ;
    END
  END DRAIN2
  PIN DRAIN3
    USE ANALOG ;
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT -7.850 9.820 -7.540 9.960 ;
        RECT -10.010 9.810 -7.540 9.820 ;
        RECT 5.490 9.820 5.800 9.960 ;
        RECT 5.490 9.810 7.960 9.820 ;
        RECT -10.010 9.640 7.960 9.810 ;
        RECT -7.850 9.630 -7.540 9.640 ;
        RECT 5.490 9.630 5.800 9.640 ;
    END
  END DRAIN3
  PIN HORIZ3
    USE ANALOG ;
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT -7.850 9.390 -7.540 9.410 ;
        RECT 5.490 9.390 5.800 9.410 ;
        RECT -10.010 9.220 7.960 9.390 ;
        RECT -10.010 9.210 -7.450 9.220 ;
        RECT 5.400 9.210 7.960 9.220 ;
        RECT -7.850 9.080 -7.540 9.210 ;
        RECT 5.490 9.080 5.800 9.210 ;
    END
  END HORIZ3
  PIN HORIZ4
    USE ANALOG ;
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT -7.850 8.410 -7.540 8.530 ;
        RECT 5.490 8.410 5.800 8.530 ;
        RECT -7.850 8.400 5.800 8.410 ;
        RECT -10.010 8.240 7.960 8.400 ;
        RECT -10.010 8.220 -7.450 8.240 ;
        RECT 5.400 8.220 7.960 8.240 ;
        RECT -7.850 8.200 -7.540 8.220 ;
        RECT 5.490 8.200 5.800 8.220 ;
    END
  END HORIZ4
  PIN DRAIN4
    USE ANALOG ;
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT -7.850 7.970 -7.540 7.980 ;
        RECT 5.490 7.970 5.800 7.980 ;
        RECT -10.010 7.800 7.960 7.970 ;
        RECT -10.010 7.790 -7.540 7.800 ;
        RECT -7.850 7.650 -7.540 7.790 ;
        RECT 5.490 7.790 7.960 7.800 ;
        RECT 5.490 7.650 5.800 7.790 ;
    END
  END DRAIN4
  PIN VINJ
    ANTENNADIFFAREA 1.088000 ;
    PORT
      LAYER nwell ;
        RECT -10.010 13.330 -7.450 13.390 ;
        RECT -10.010 7.280 -3.450 13.330 ;
        RECT -10.010 7.230 -7.450 7.280 ;
      LAYER met1 ;
        RECT -9.650 12.680 -9.490 13.380 ;
        RECT -9.650 12.130 -9.380 12.680 ;
        RECT -9.660 12.080 -9.380 12.130 ;
        RECT -9.660 11.990 -9.490 12.080 ;
        RECT -9.650 11.630 -9.490 11.990 ;
        RECT -9.660 11.540 -9.490 11.630 ;
        RECT -9.660 11.490 -9.380 11.540 ;
        RECT -9.650 10.940 -9.380 11.490 ;
        RECT -9.650 9.670 -9.490 10.940 ;
        RECT -9.650 9.120 -9.380 9.670 ;
        RECT -9.660 9.070 -9.380 9.120 ;
        RECT -9.660 8.980 -9.490 9.070 ;
        RECT -9.650 8.630 -9.490 8.980 ;
        RECT -9.660 8.540 -9.490 8.630 ;
        RECT -9.660 8.490 -9.380 8.540 ;
        RECT -9.650 7.940 -9.380 8.490 ;
        RECT -9.650 7.240 -9.490 7.940 ;
    END
    PORT
      LAYER nwell ;
        RECT 5.400 13.330 7.960 13.390 ;
        RECT 1.400 7.280 7.960 13.330 ;
        RECT 5.400 7.230 7.960 7.280 ;
      LAYER met1 ;
        RECT 7.440 12.680 7.600 13.380 ;
        RECT 7.330 12.130 7.600 12.680 ;
        RECT 7.330 12.080 7.610 12.130 ;
        RECT 7.440 11.990 7.610 12.080 ;
        RECT 7.440 11.630 7.600 11.990 ;
        RECT 7.440 11.540 7.610 11.630 ;
        RECT 7.330 11.490 7.610 11.540 ;
        RECT 7.330 10.940 7.600 11.490 ;
        RECT 7.440 9.670 7.600 10.940 ;
        RECT 7.330 9.120 7.600 9.670 ;
        RECT 7.330 9.070 7.610 9.120 ;
        RECT 7.440 8.980 7.610 9.070 ;
        RECT 7.440 8.630 7.600 8.980 ;
        RECT 7.440 8.540 7.610 8.630 ;
        RECT 7.330 8.490 7.610 8.540 ;
        RECT 7.330 7.940 7.600 8.490 ;
        RECT 7.440 7.240 7.600 7.940 ;
    END
  END VINJ
  PIN GATESELECT1
    USE ANALOG ;
    ANTENNAGATEAREA 0.720000 ;
    PORT
      LAYER met1 ;
        RECT -9.240 12.340 -9.050 13.330 ;
        RECT -9.240 12.220 -9.070 12.340 ;
        RECT -9.240 11.400 -9.080 12.220 ;
        RECT -9.240 11.280 -9.070 11.400 ;
        RECT -9.240 10.420 -9.050 11.280 ;
        RECT -9.270 10.190 -9.030 10.420 ;
        RECT -9.240 9.330 -9.050 10.190 ;
        RECT -9.240 9.210 -9.070 9.330 ;
        RECT -9.240 8.400 -9.080 9.210 ;
        RECT -9.240 8.280 -9.070 8.400 ;
        RECT -9.240 7.290 -9.050 8.280 ;
    END
  END GATESELECT1
  PIN VERT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met1 ;
        RECT 6.630 12.650 6.790 13.380 ;
        RECT 6.630 12.630 6.830 12.650 ;
        RECT 6.610 12.390 6.840 12.630 ;
        RECT 6.630 12.340 6.840 12.390 ;
        RECT 6.630 11.280 6.790 12.340 ;
        RECT 6.630 11.230 6.840 11.280 ;
        RECT 6.610 10.990 6.840 11.230 ;
        RECT 6.630 10.970 6.830 10.990 ;
        RECT 6.630 9.640 6.790 10.970 ;
        RECT 6.630 9.620 6.830 9.640 ;
        RECT 6.610 9.380 6.840 9.620 ;
        RECT 6.630 9.330 6.840 9.380 ;
        RECT 6.630 8.280 6.790 9.330 ;
        RECT 6.630 8.230 6.840 8.280 ;
        RECT 6.610 7.990 6.840 8.230 ;
        RECT 6.630 7.970 6.830 7.990 ;
        RECT 6.630 7.240 6.790 7.970 ;
    END
  END VERT2
  PIN GATESELECT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.720000 ;
    PORT
      LAYER met1 ;
        RECT 7.000 12.340 7.190 13.330 ;
        RECT 7.020 12.220 7.190 12.340 ;
        RECT 7.030 11.400 7.190 12.220 ;
        RECT 7.020 11.280 7.190 11.400 ;
        RECT 7.000 10.420 7.190 11.280 ;
        RECT 6.980 10.190 7.220 10.420 ;
        RECT 7.000 9.330 7.190 10.190 ;
        RECT 7.020 9.210 7.190 9.330 ;
        RECT 7.030 8.400 7.190 9.210 ;
        RECT 7.020 8.280 7.190 8.400 ;
        RECT 7.000 7.290 7.190 8.280 ;
    END
  END GATESELECT2
  PIN GATE2
    USE ANALOG ;
    ANTENNADIFFAREA 1.345600 ;
    PORT
      LAYER met1 ;
        RECT 3.280 12.100 3.520 13.330 ;
        RECT 3.280 11.880 3.530 12.100 ;
        RECT 3.280 10.630 3.520 11.880 ;
        RECT 3.280 10.410 3.530 10.630 ;
        RECT 3.280 9.160 3.520 10.410 ;
        RECT 3.280 8.940 3.530 9.160 ;
        RECT 3.280 7.690 3.520 8.940 ;
        RECT 3.280 7.470 3.530 7.690 ;
        RECT 3.280 7.280 3.520 7.470 ;
    END
  END GATE2
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 1.345600 ;
    PORT
      LAYER met1 ;
        RECT -5.570 12.100 -5.320 13.330 ;
        RECT -5.580 11.880 -5.320 12.100 ;
        RECT -5.570 10.630 -5.320 11.880 ;
        RECT -5.580 10.410 -5.320 10.630 ;
        RECT -5.570 9.160 -5.320 10.410 ;
        RECT -5.580 8.940 -5.320 9.160 ;
        RECT -5.570 7.690 -5.320 8.940 ;
        RECT -5.580 7.470 -5.320 7.690 ;
        RECT -5.570 7.280 -5.320 7.470 ;
    END
  END GATE1
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 0.336400 ;
    PORT
      LAYER met1 ;
        RECT -1.960 7.280 -1.660 13.330 ;
    END
    PORT
      LAYER met1 ;
        RECT -0.380 7.280 -0.080 13.330 ;
    END
  END VTUN
  OBS
      LAYER li1 ;
        RECT -9.610 12.650 -9.410 13.000 ;
        RECT -7.870 12.920 -7.550 12.930 ;
        RECT -8.130 12.750 -7.550 12.920 ;
        RECT -7.880 12.700 -7.550 12.750 ;
        RECT -7.870 12.670 -7.550 12.700 ;
        RECT -9.620 12.620 -9.410 12.650 ;
        RECT -9.620 12.030 -9.400 12.620 ;
        RECT -8.880 12.030 -8.680 12.630 ;
        RECT -7.870 12.340 -7.550 12.380 ;
        RECT -7.880 12.300 -7.550 12.340 ;
        RECT -8.130 12.130 -7.550 12.300 ;
        RECT -7.870 12.120 -7.550 12.130 ;
        RECT -7.110 12.020 -3.800 13.000 ;
        RECT -1.890 12.120 -1.720 13.010 ;
        RECT -0.330 12.120 -0.160 13.010 ;
        RECT 1.750 12.020 5.060 13.000 ;
        RECT 5.500 12.920 5.820 12.930 ;
        RECT 5.500 12.750 6.080 12.920 ;
        RECT 5.500 12.700 5.830 12.750 ;
        RECT 5.500 12.670 5.820 12.700 ;
        RECT 7.360 12.650 7.560 13.000 ;
        RECT 5.500 12.340 5.820 12.380 ;
        RECT 5.500 12.300 5.830 12.340 ;
        RECT 5.500 12.130 6.080 12.300 ;
        RECT 5.500 12.120 5.820 12.130 ;
        RECT 6.630 12.030 6.830 12.630 ;
        RECT 7.360 12.620 7.570 12.650 ;
        RECT 7.350 12.030 7.570 12.620 ;
        RECT -9.620 11.000 -9.400 11.590 ;
        RECT -9.620 10.970 -9.410 11.000 ;
        RECT -8.880 10.990 -8.680 11.590 ;
        RECT -7.870 11.490 -7.550 11.500 ;
        RECT -8.130 11.320 -7.550 11.490 ;
        RECT -7.880 11.280 -7.550 11.320 ;
        RECT -7.870 11.240 -7.550 11.280 ;
        RECT -9.610 10.620 -9.410 10.970 ;
        RECT -7.870 10.920 -7.550 10.950 ;
        RECT -7.880 10.870 -7.550 10.920 ;
        RECT -8.130 10.700 -7.550 10.870 ;
        RECT -7.870 10.690 -7.550 10.700 ;
        RECT -7.110 10.550 -3.800 11.530 ;
        RECT -1.890 10.600 -1.720 11.490 ;
        RECT -0.330 10.600 -0.160 11.490 ;
        RECT 1.750 10.550 5.060 11.530 ;
        RECT 5.500 11.490 5.820 11.500 ;
        RECT 5.500 11.320 6.080 11.490 ;
        RECT 5.500 11.280 5.830 11.320 ;
        RECT 5.500 11.240 5.820 11.280 ;
        RECT 6.630 10.990 6.830 11.590 ;
        RECT 7.350 11.000 7.570 11.590 ;
        RECT 7.360 10.970 7.570 11.000 ;
        RECT 5.500 10.920 5.820 10.950 ;
        RECT 5.500 10.870 5.830 10.920 ;
        RECT 5.500 10.700 6.080 10.870 ;
        RECT 5.500 10.690 5.820 10.700 ;
        RECT 7.360 10.620 7.560 10.970 ;
        RECT -9.240 10.220 -8.800 10.390 ;
        RECT 6.750 10.220 7.190 10.390 ;
        RECT -9.610 9.640 -9.410 9.990 ;
        RECT -7.870 9.910 -7.550 9.920 ;
        RECT -8.130 9.740 -7.550 9.910 ;
        RECT -7.880 9.690 -7.550 9.740 ;
        RECT -7.870 9.660 -7.550 9.690 ;
        RECT -9.620 9.610 -9.410 9.640 ;
        RECT -9.620 9.020 -9.400 9.610 ;
        RECT -8.880 9.020 -8.680 9.620 ;
        RECT -7.870 9.330 -7.550 9.370 ;
        RECT -7.880 9.290 -7.550 9.330 ;
        RECT -8.130 9.120 -7.550 9.290 ;
        RECT -7.870 9.110 -7.550 9.120 ;
        RECT -7.110 9.080 -3.800 10.060 ;
        RECT -1.890 9.150 -1.720 10.040 ;
        RECT -0.330 9.150 -0.160 10.040 ;
        RECT 1.750 9.080 5.060 10.060 ;
        RECT 5.500 9.910 5.820 9.920 ;
        RECT 5.500 9.740 6.080 9.910 ;
        RECT 5.500 9.690 5.830 9.740 ;
        RECT 5.500 9.660 5.820 9.690 ;
        RECT 7.360 9.640 7.560 9.990 ;
        RECT 5.500 9.330 5.820 9.370 ;
        RECT 5.500 9.290 5.830 9.330 ;
        RECT 5.500 9.120 6.080 9.290 ;
        RECT 5.500 9.110 5.820 9.120 ;
        RECT 6.630 9.020 6.830 9.620 ;
        RECT 7.360 9.610 7.570 9.640 ;
        RECT 7.350 9.020 7.570 9.610 ;
        RECT -9.620 8.000 -9.400 8.590 ;
        RECT -9.620 7.970 -9.410 8.000 ;
        RECT -8.880 7.990 -8.680 8.590 ;
        RECT -7.870 8.490 -7.550 8.500 ;
        RECT -8.130 8.320 -7.550 8.490 ;
        RECT -7.880 8.280 -7.550 8.320 ;
        RECT -7.870 8.240 -7.550 8.280 ;
        RECT -9.610 7.620 -9.410 7.970 ;
        RECT -7.870 7.920 -7.550 7.950 ;
        RECT -7.880 7.870 -7.550 7.920 ;
        RECT -8.130 7.700 -7.550 7.870 ;
        RECT -7.870 7.690 -7.550 7.700 ;
        RECT -7.110 7.610 -3.800 8.590 ;
        RECT -1.890 7.610 -1.720 8.500 ;
        RECT -0.330 7.610 -0.160 8.500 ;
        RECT 1.750 7.610 5.060 8.590 ;
        RECT 5.500 8.490 5.820 8.500 ;
        RECT 5.500 8.320 6.080 8.490 ;
        RECT 5.500 8.280 5.830 8.320 ;
        RECT 5.500 8.240 5.820 8.280 ;
        RECT 6.630 7.990 6.830 8.590 ;
        RECT 7.350 8.000 7.570 8.590 ;
        RECT 7.360 7.970 7.570 8.000 ;
        RECT 5.500 7.920 5.820 7.950 ;
        RECT 5.500 7.870 5.830 7.920 ;
        RECT 5.500 7.700 6.080 7.870 ;
        RECT 5.500 7.690 5.820 7.700 ;
        RECT 7.360 7.620 7.560 7.970 ;
      LAYER mcon ;
        RECT -7.780 12.710 -7.610 12.880 ;
        RECT -5.540 12.770 -5.370 12.940 ;
        RECT -9.590 12.450 -9.420 12.620 ;
        RECT -8.860 12.420 -8.690 12.590 ;
        RECT -7.780 12.160 -7.610 12.330 ;
        RECT -5.540 12.080 -5.370 12.250 ;
        RECT -1.890 12.810 -1.720 12.980 ;
        RECT -0.330 12.810 -0.160 12.980 ;
        RECT 3.320 12.770 3.490 12.940 ;
        RECT 5.560 12.710 5.730 12.880 ;
        RECT 6.640 12.420 6.810 12.590 ;
        RECT 3.320 12.080 3.490 12.250 ;
        RECT 5.560 12.160 5.730 12.330 ;
        RECT 7.370 12.450 7.540 12.620 ;
        RECT -9.590 11.000 -9.420 11.170 ;
        RECT -7.780 11.290 -7.610 11.460 ;
        RECT -5.540 11.300 -5.370 11.470 ;
        RECT -8.860 11.030 -8.690 11.200 ;
        RECT -7.780 10.740 -7.610 10.910 ;
        RECT -5.540 10.610 -5.370 10.780 ;
        RECT -1.890 11.290 -1.720 11.460 ;
        RECT -0.330 11.290 -0.160 11.460 ;
        RECT 3.320 11.300 3.490 11.470 ;
        RECT 5.560 11.290 5.730 11.460 ;
        RECT 6.640 11.030 6.810 11.200 ;
        RECT 7.370 11.000 7.540 11.170 ;
        RECT 3.320 10.610 3.490 10.780 ;
        RECT 5.560 10.740 5.730 10.910 ;
        RECT 7.010 10.220 7.190 10.390 ;
        RECT -7.780 9.700 -7.610 9.870 ;
        RECT -5.540 9.830 -5.370 10.000 ;
        RECT -9.590 9.440 -9.420 9.610 ;
        RECT -8.860 9.410 -8.690 9.580 ;
        RECT -7.780 9.150 -7.610 9.320 ;
        RECT -5.540 9.140 -5.370 9.310 ;
        RECT -1.890 9.840 -1.720 10.010 ;
        RECT -0.330 9.840 -0.160 10.010 ;
        RECT 3.320 9.830 3.490 10.000 ;
        RECT 5.560 9.700 5.730 9.870 ;
        RECT 6.640 9.410 6.810 9.580 ;
        RECT 3.320 9.140 3.490 9.310 ;
        RECT 5.560 9.150 5.730 9.320 ;
        RECT 7.370 9.440 7.540 9.610 ;
        RECT -9.590 8.000 -9.420 8.170 ;
        RECT -7.780 8.290 -7.610 8.460 ;
        RECT -5.540 8.360 -5.370 8.530 ;
        RECT -8.860 8.030 -8.690 8.200 ;
        RECT -7.780 7.740 -7.610 7.910 ;
        RECT -5.540 7.670 -5.370 7.840 ;
        RECT -1.890 8.300 -1.720 8.470 ;
        RECT -0.330 8.300 -0.160 8.470 ;
        RECT 3.320 8.360 3.490 8.530 ;
        RECT 5.560 8.290 5.730 8.460 ;
        RECT 6.640 8.030 6.810 8.200 ;
        RECT 7.370 8.000 7.540 8.170 ;
        RECT 3.320 7.670 3.490 7.840 ;
        RECT 5.560 7.740 5.730 7.910 ;
      LAYER met1 ;
        RECT -7.860 12.640 -7.540 12.960 ;
        RECT 5.490 12.640 5.810 12.960 ;
        RECT -7.860 12.090 -7.540 12.410 ;
        RECT 5.490 12.090 5.810 12.410 ;
        RECT -7.860 11.210 -7.540 11.530 ;
        RECT 5.490 11.210 5.810 11.530 ;
        RECT -7.860 10.660 -7.540 10.980 ;
        RECT 5.490 10.660 5.810 10.980 ;
        RECT -7.860 9.630 -7.540 9.950 ;
        RECT 5.490 9.630 5.810 9.950 ;
        RECT -7.860 9.080 -7.540 9.400 ;
        RECT 5.490 9.080 5.810 9.400 ;
        RECT -7.860 8.210 -7.540 8.530 ;
        RECT 5.490 8.210 5.810 8.530 ;
        RECT -7.860 7.660 -7.540 7.980 ;
        RECT 5.490 7.660 5.810 7.980 ;
      LAYER via ;
        RECT -7.830 12.670 -7.570 12.930 ;
        RECT 5.520 12.670 5.780 12.930 ;
        RECT -7.830 12.120 -7.570 12.380 ;
        RECT 5.520 12.120 5.780 12.380 ;
        RECT -7.830 11.240 -7.570 11.500 ;
        RECT 5.520 11.240 5.780 11.500 ;
        RECT -7.830 10.690 -7.570 10.950 ;
        RECT 5.520 10.690 5.780 10.950 ;
        RECT -7.830 9.660 -7.570 9.920 ;
        RECT 5.520 9.660 5.780 9.920 ;
        RECT -7.830 9.110 -7.570 9.370 ;
        RECT 5.520 9.110 5.780 9.370 ;
        RECT -7.830 8.240 -7.570 8.500 ;
        RECT 5.520 8.240 5.780 8.500 ;
        RECT -7.830 7.690 -7.570 7.950 ;
        RECT 5.520 7.690 5.780 7.950 ;
  END
END sky130_hilas_swc4x2cellOverlap

MACRO sky130_hilas_TopLevelTextStructure
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TopLevelTextStructure ;
  ORIGIN -2.180 7.930 ;
  SIZE 130.250 BY 75.780 ;
  PIN DIG24 
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 59.800 22.940 60.110 22.960 ;
        RECT 67.600 22.940 67.740 22.950 ;
        RECT 57.640 22.760 67.750 22.940 ;
        RECT 59.800 22.750 67.750 22.760 ;
        RECT 59.800 22.630 60.110 22.750 ;
        RECT 67.600 22.610 67.750 22.750 ;
        RECT 67.600 22.520 68.810 22.610 ;
        RECT 67.600 22.460 68.940 22.520 ;
        RECT 67.600 22.450 71.210 22.460 ;
        RECT 75.910 22.450 76.230 22.500 ;
        RECT 67.600 22.410 76.230 22.450 ;
        RECT 68.630 22.300 76.230 22.410 ;
        RECT 68.630 22.190 68.940 22.300 ;
        RECT 71.130 22.290 76.230 22.300 ;
        RECT 75.910 22.240 76.230 22.290 ;
        RECT 75.890 12.830 132.430 13.330 ;
        RECT 130.420 -7.170 132.430 12.830 ;
        RECT 130.390 -7.750 132.430 -7.170 ;
        RECT 130.390 -7.820 132.420 -7.750 ;
    END
  END DIG24 
  PIN DIG23
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 59.800 21.850 60.110 21.980 ;
        RECT 57.640 21.670 68.910 21.850 ;
        RECT 59.800 21.650 60.110 21.670 ;
        RECT 68.630 21.640 68.910 21.670 ;
        RECT 68.630 21.530 68.940 21.640 ;
        RECT 68.630 21.520 71.210 21.530 ;
        RECT 75.390 21.520 75.710 21.570 ;
        RECT 68.630 21.370 75.710 21.520 ;
        RECT 68.630 21.310 68.940 21.370 ;
        RECT 71.130 21.360 75.710 21.370 ;
        RECT 75.390 21.310 75.710 21.360 ;
        RECT 126.330 12.430 128.340 12.450 ;
        RECT 75.350 11.930 128.340 12.430 ;
        RECT 126.330 -7.190 128.340 11.930 ;
        RECT 126.330 -7.840 128.370 -7.190 ;
        RECT 126.330 -7.920 128.340 -7.840 ;
    END
  END DIG23
  PIN DIG22
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 68.630 19.720 68.940 19.750 ;
        RECT 67.240 19.690 68.940 19.720 ;
        RECT 67.240 19.680 71.210 19.690 ;
        RECT 74.920 19.680 75.240 19.730 ;
        RECT 67.240 19.560 75.240 19.680 ;
        RECT 67.240 19.550 67.700 19.560 ;
        RECT 68.630 19.530 75.240 19.560 ;
        RECT 68.630 19.420 68.940 19.530 ;
        RECT 71.130 19.520 75.240 19.530 ;
        RECT 74.920 19.470 75.240 19.520 ;
        RECT 74.880 11.510 124.150 11.530 ;
        RECT 74.880 11.030 124.260 11.510 ;
        RECT 122.250 -7.170 124.260 11.030 ;
        RECT 122.250 -7.820 124.320 -7.170 ;
        RECT 122.250 -7.860 124.260 -7.820 ;
    END
  END DIG22
  PIN DIG21
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 68.630 18.760 68.940 18.870 ;
        RECT 68.630 18.750 71.210 18.760 ;
        RECT 74.420 18.750 74.740 18.800 ;
        RECT 67.700 18.740 74.740 18.750 ;
        RECT 60.080 18.730 74.740 18.740 ;
        RECT 59.800 18.600 74.740 18.730 ;
        RECT 57.640 18.570 68.940 18.600 ;
        RECT 71.130 18.590 74.740 18.600 ;
        RECT 57.640 18.420 60.200 18.570 ;
        RECT 68.630 18.540 68.940 18.570 ;
        RECT 74.420 18.540 74.740 18.590 ;
        RECT 59.800 18.400 60.110 18.420 ;
        RECT 74.400 10.620 120.190 10.630 ;
        RECT 74.400 10.130 120.400 10.620 ;
        RECT 118.390 -7.170 120.400 10.130 ;
        RECT 118.330 -7.690 120.400 -7.170 ;
        RECT 118.330 -7.820 120.360 -7.690 ;
    END
  END DIG21
  PIN DIG29
    ANTENNAGATEAREA 3.650400 ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.260 110.350 0.580 ;
        RECT 110.140 -1.030 110.330 0.260 ;
        RECT 110.020 -1.350 110.340 -1.030 ;
        RECT 110.140 -4.230 110.330 -1.350 ;
        RECT 110.020 -4.550 110.340 -4.230 ;
        RECT 110.140 -5.940 110.330 -4.550 ;
        RECT 109.980 -6.260 110.330 -5.940 ;
        RECT 110.120 -6.470 110.330 -6.260 ;
        RECT 110.120 -6.490 115.140 -6.470 ;
        RECT 110.140 -6.660 115.140 -6.490 ;
        RECT 114.950 -7.120 115.140 -6.660 ;
        RECT 114.950 -7.190 115.980 -7.120 ;
        RECT 114.280 -7.840 116.310 -7.190 ;
    END
  END DIG29
  PIN DIG28
    ANTENNAGATEAREA 2.281500 ;
    PORT
      LAYER met2 ;
        RECT 109.020 2.160 109.330 2.190 ;
        RECT 110.020 2.160 110.340 2.200 ;
        RECT 109.020 1.910 110.340 2.160 ;
        RECT 109.020 -2.790 109.320 1.910 ;
        RECT 110.020 1.880 110.340 1.910 ;
        RECT 109.610 -2.790 109.930 -2.680 ;
        RECT 109.020 -3.000 109.930 -2.790 ;
        RECT 109.020 -3.010 109.780 -3.000 ;
        RECT 109.020 -4.430 109.320 -3.010 ;
        RECT 109.020 -4.590 109.380 -4.430 ;
        RECT 108.670 -6.030 108.990 -5.960 ;
        RECT 109.170 -6.030 109.380 -4.590 ;
        RECT 108.670 -6.230 109.380 -6.030 ;
        RECT 108.670 -6.280 108.990 -6.230 ;
        RECT 109.170 -7.260 109.380 -6.230 ;
        RECT 110.300 -7.260 112.330 -7.170 ;
        RECT 109.170 -7.470 112.330 -7.260 ;
        RECT 110.300 -7.820 112.330 -7.470 ;
    END
  END DIG28
  PIN DIG27
    ANTENNAGATEAREA 0.608400 ;
    PORT
      LAYER met2 ;
        RECT 107.240 3.810 110.050 3.820 ;
        RECT 107.240 3.620 110.350 3.810 ;
        RECT 107.240 -7.170 107.450 3.620 ;
        RECT 110.030 3.490 110.350 3.620 ;
        RECT 106.120 -7.820 108.150 -7.170 ;
    END
  END DIG27
  PIN DIG26
    ANTENNAGATEAREA 0.456300 ;
    PORT
      LAYER met2 ;
        RECT 106.270 5.370 106.470 5.380 ;
        RECT 110.030 5.370 110.350 5.420 ;
        RECT 106.270 5.220 110.350 5.370 ;
        RECT 106.270 -6.350 106.470 5.220 ;
        RECT 110.030 5.100 110.350 5.220 ;
        RECT 106.260 -6.490 106.470 -6.350 ;
        RECT 106.270 -6.700 106.470 -6.490 ;
        RECT 104.040 -6.900 106.470 -6.700 ;
        RECT 104.040 -7.170 104.240 -6.900 ;
        RECT 102.040 -7.470 104.240 -7.170 ;
        RECT 102.040 -7.820 104.070 -7.470 ;
    END
  END DIG26
  PIN DIG25
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER met2 ;
        RECT 105.120 1.770 105.380 2.090 ;
        RECT 105.150 -6.290 105.350 1.770 ;
        RECT 99.110 -6.490 105.350 -6.290 ;
        RECT 99.110 -7.170 99.310 -6.490 ;
        RECT 98.020 -7.820 100.050 -7.170 ;
    END
  END DIG25
  PIN DIG20
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT 103.020 39.410 103.420 39.420 ;
        RECT 103.000 39.350 103.440 39.410 ;
        RECT 103.000 39.170 106.850 39.350 ;
        RECT 107.730 39.170 108.050 39.260 ;
        RECT 103.000 39.150 108.050 39.170 ;
        RECT 103.020 39.140 103.420 39.150 ;
        RECT 106.500 38.970 108.050 39.150 ;
        RECT 103.010 -3.120 103.430 -3.090 ;
        RECT 94.040 -3.500 103.430 -3.120 ;
        RECT 94.040 -7.200 96.020 -3.500 ;
        RECT 103.010 -3.530 103.430 -3.500 ;
        RECT 94.030 -7.850 96.060 -7.200 ;
    END
  END DIG20
  PIN DIG19
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT 102.200 40.110 102.590 40.130 ;
        RECT 102.190 40.000 102.600 40.110 ;
        RECT 102.190 39.900 106.850 40.000 ;
        RECT 102.190 39.800 108.050 39.900 ;
        RECT 102.190 39.700 102.600 39.800 ;
        RECT 106.620 39.700 108.050 39.800 ;
        RECT 102.200 39.680 102.590 39.700 ;
        RECT 107.730 39.610 108.050 39.700 ;
        RECT 102.170 -2.330 102.620 -2.320 ;
        RECT 89.930 -2.710 102.620 -2.330 ;
        RECT 89.930 -7.170 91.910 -2.710 ;
        RECT 89.890 -7.820 91.920 -7.170 ;
    END
  END DIG19
  PIN DIG18
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT 101.280 42.370 101.640 42.470 ;
        RECT 107.730 42.370 108.050 42.460 ;
        RECT 101.280 42.170 108.050 42.370 ;
        RECT 101.280 42.050 101.640 42.170 ;
        RECT 101.250 -1.500 101.680 -1.480 ;
        RECT 101.240 -1.510 101.690 -1.500 ;
        RECT 85.780 -1.890 101.690 -1.510 ;
        RECT 85.780 -7.190 87.740 -1.890 ;
        RECT 101.250 -1.910 101.680 -1.890 ;
        RECT 85.770 -7.840 87.800 -7.190 ;
    END
  END DIG18
  PIN DIG17
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT 100.270 43.020 100.730 43.150 ;
        RECT 106.580 43.020 108.050 43.100 ;
        RECT 100.270 42.900 108.050 43.020 ;
        RECT 100.270 42.820 106.850 42.900 ;
        RECT 100.270 42.700 100.730 42.820 ;
        RECT 107.730 42.810 108.050 42.900 ;
        RECT 100.350 -0.690 100.780 -0.670 ;
        RECT 81.850 -0.720 83.810 -0.690 ;
        RECT 100.330 -0.720 100.790 -0.690 ;
        RECT 81.850 -1.070 100.790 -0.720 ;
        RECT 81.850 -7.170 83.810 -1.070 ;
        RECT 100.330 -1.090 100.790 -1.070 ;
        RECT 100.350 -1.100 100.780 -1.090 ;
        RECT 81.820 -7.820 83.850 -7.170 ;
    END
  END DIG17
  PIN DIG16
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 40.870 49.380 41.330 49.450 ;
        RECT 40.480 49.210 41.330 49.380 ;
        RECT 39.510 48.650 39.900 48.740 ;
        RECT 40.480 48.650 40.650 49.210 ;
        RECT 40.870 49.130 41.330 49.210 ;
        RECT 39.510 48.480 40.660 48.650 ;
        RECT 39.490 -0.230 39.910 -0.220 ;
        RECT 39.490 -0.480 79.760 -0.230 ;
        RECT 39.490 -0.560 79.770 -0.480 ;
        RECT 39.490 -0.570 39.910 -0.560 ;
        RECT 73.730 -0.580 79.770 -0.560 ;
        RECT 77.830 -1.080 79.770 -0.580 ;
        RECT 77.830 -7.150 79.760 -1.080 ;
        RECT 77.740 -7.930 79.770 -7.150 ;
    END
  END DIG16
  PIN DIG15
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 40.870 47.550 41.330 47.700 ;
        RECT 40.480 47.380 41.330 47.550 ;
        RECT 38.910 47.110 39.240 47.120 ;
        RECT 38.890 47.010 39.260 47.110 ;
        RECT 40.480 47.010 40.650 47.380 ;
        RECT 38.890 46.840 40.650 47.010 ;
        RECT 38.890 46.730 39.260 46.840 ;
        RECT 40.480 46.830 40.650 46.840 ;
        RECT 38.890 -0.850 39.270 -0.840 ;
        RECT 38.890 -1.180 75.690 -0.850 ;
        RECT 38.890 -1.190 39.270 -1.180 ;
        RECT 69.620 -1.190 75.690 -1.180 ;
        RECT 73.730 -1.510 75.690 -1.190 ;
        RECT 73.730 -7.170 75.680 -1.510 ;
        RECT 73.670 -7.820 75.700 -7.170 ;
    END
  END DIG15
  PIN DIG14
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 40.870 45.820 41.330 45.950 ;
        RECT 40.440 45.650 41.330 45.820 ;
        RECT 38.310 45.530 38.700 45.630 ;
        RECT 40.440 45.530 40.610 45.650 ;
        RECT 40.870 45.630 41.330 45.650 ;
        RECT 38.310 45.360 40.610 45.530 ;
        RECT 38.310 45.260 38.700 45.360 ;
        RECT 38.250 -1.480 38.670 -1.470 ;
        RECT 38.250 -1.810 71.610 -1.480 ;
        RECT 38.250 -1.820 38.670 -1.810 ;
        RECT 69.620 -7.170 71.610 -1.810 ;
        RECT 69.620 -7.820 71.650 -7.170 ;
    END
  END DIG14
  PIN DIG13
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 40.870 44.100 41.330 44.200 ;
        RECT 37.670 43.930 38.060 44.020 ;
        RECT 40.610 43.930 41.330 44.100 ;
        RECT 37.670 43.880 41.330 43.930 ;
        RECT 37.670 43.760 41.240 43.880 ;
        RECT 37.670 43.670 38.060 43.760 ;
        RECT 40.610 43.740 40.780 43.760 ;
        RECT 37.660 -2.120 38.060 -2.100 ;
        RECT 37.660 -2.450 67.600 -2.120 ;
        RECT 37.660 -2.460 38.060 -2.450 ;
        RECT 65.640 -7.170 67.590 -2.450 ;
        RECT 65.590 -7.820 67.620 -7.170 ;
    END
  END DIG13
  PIN DIG12
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 37.030 43.360 37.420 43.470 ;
        RECT 40.870 43.360 41.330 43.410 ;
        RECT 37.030 43.190 41.330 43.360 ;
        RECT 37.030 43.090 37.420 43.190 ;
        RECT 40.870 43.090 41.330 43.190 ;
        RECT 37.000 -2.790 37.410 -2.780 ;
        RECT 36.990 -3.120 63.510 -2.790 ;
        RECT 37.000 -3.140 37.410 -3.120 ;
        RECT 61.600 -7.190 63.510 -3.120 ;
        RECT 61.520 -7.840 63.550 -7.190 ;
    END
  END DIG12
  PIN DIG11
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 36.420 41.790 36.810 41.890 ;
        RECT 36.420 41.660 41.240 41.790 ;
        RECT 36.420 41.620 41.330 41.660 ;
        RECT 36.420 41.520 36.810 41.620 ;
        RECT 40.690 41.460 41.330 41.620 ;
        RECT 40.870 41.340 41.330 41.460 ;
        RECT 36.420 -3.410 36.830 -3.400 ;
        RECT 36.420 -3.430 59.490 -3.410 ;
        RECT 36.420 -3.740 59.500 -3.430 ;
        RECT 36.420 -3.750 36.830 -3.740 ;
        RECT 57.500 -7.120 59.500 -3.740 ;
        RECT 57.470 -7.820 59.500 -7.120 ;
    END
  END DIG11
  PIN DIG10
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 35.790 40.260 36.210 40.350 ;
        RECT 35.790 40.090 40.690 40.260 ;
        RECT 35.790 40.000 36.210 40.090 ;
        RECT 40.520 39.910 40.690 40.090 ;
        RECT 40.520 39.740 41.330 39.910 ;
        RECT 40.870 39.590 41.330 39.740 ;
        RECT 35.820 -4.060 36.210 -4.050 ;
        RECT 35.820 -4.380 55.510 -4.060 ;
        RECT 35.920 -4.390 55.510 -4.380 ;
        RECT 53.520 -7.100 55.510 -4.390 ;
        RECT 53.510 -7.850 55.540 -7.100 ;
    END
  END DIG10
  PIN DIG09
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 35.230 38.690 35.620 38.780 ;
        RECT 35.230 38.520 40.600 38.690 ;
        RECT 35.230 38.430 35.620 38.520 ;
        RECT 40.440 38.410 40.600 38.520 ;
        RECT 40.440 38.110 40.610 38.410 ;
        RECT 40.870 38.110 41.330 38.160 ;
        RECT 40.440 37.940 41.330 38.110 ;
        RECT 40.870 37.840 41.330 37.940 ;
        RECT 35.240 -4.670 35.630 -4.620 ;
        RECT 35.240 -4.950 51.600 -4.670 ;
        RECT 35.500 -5.000 51.600 -4.950 ;
        RECT 49.530 -7.820 51.560 -5.000 ;
    END
  END DIG09
  PIN DIG08
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 34.620 33.220 34.990 33.340 ;
        RECT 40.870 33.220 41.330 33.280 ;
        RECT 34.620 33.050 41.330 33.220 ;
        RECT 34.620 32.940 34.990 33.050 ;
        RECT 40.870 32.960 41.330 33.050 ;
        RECT 34.660 -5.640 47.400 -5.310 ;
        RECT 45.350 -6.940 47.380 -5.640 ;
        RECT 45.350 -7.230 47.390 -6.940 ;
        RECT 45.360 -7.840 47.390 -7.230 ;
    END
  END DIG08
  PIN DIG07
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 33.980 31.630 34.370 31.720 ;
        RECT 33.980 31.530 40.940 31.630 ;
        RECT 33.980 31.460 41.330 31.530 ;
        RECT 33.980 31.370 34.370 31.460 ;
        RECT 40.650 31.340 41.330 31.460 ;
        RECT 40.870 31.210 41.330 31.340 ;
        RECT 41.270 -5.940 43.290 -5.920 ;
        RECT 34.110 -5.950 43.320 -5.940 ;
        RECT 34.010 -6.270 43.320 -5.950 ;
        RECT 34.010 -6.280 34.400 -6.270 ;
        RECT 41.240 -7.820 43.320 -6.270 ;
    END
  END DIG07
  PIN DIG06
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 33.360 30.080 33.750 30.160 ;
        RECT 33.360 29.910 40.540 30.080 ;
        RECT 33.360 29.830 33.750 29.910 ;
        RECT 40.390 29.840 40.540 29.910 ;
        RECT 40.390 29.730 40.560 29.840 ;
        RECT 40.870 29.730 41.330 29.780 ;
        RECT 40.390 29.560 41.330 29.730 ;
        RECT 40.870 29.460 41.330 29.560 ;
        RECT 33.370 -6.930 39.350 -6.590 ;
        RECT 37.320 -7.190 39.360 -6.930 ;
        RECT 37.310 -7.850 39.360 -7.190 ;
    END
  END DIG06
  PIN DIG05
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 32.750 28.600 33.170 28.690 ;
        RECT 32.750 28.430 40.560 28.600 ;
        RECT 32.750 28.330 33.170 28.430 ;
        RECT 40.390 27.940 40.560 28.430 ;
        RECT 40.870 27.940 41.330 28.030 ;
        RECT 40.390 27.770 41.330 27.940 ;
        RECT 40.870 27.710 41.330 27.770 ;
        RECT 32.760 -7.180 33.310 -7.160 ;
        RECT 32.760 -7.610 35.310 -7.180 ;
        RECT 33.280 -7.840 35.310 -7.610 ;
    END
  END DIG05
  PIN DIG04
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 40.830 24.140 41.290 24.220 ;
        RECT 40.580 23.900 41.290 24.140 ;
        RECT 40.580 23.870 40.960 23.900 ;
        RECT 40.580 23.650 40.860 23.870 ;
        RECT 32.110 23.430 32.520 23.530 ;
        RECT 40.580 23.430 40.850 23.650 ;
        RECT 32.110 23.260 40.850 23.430 ;
        RECT 32.110 23.170 32.520 23.260 ;
        RECT 40.580 23.250 40.750 23.260 ;
        RECT 31.260 -7.160 31.910 -7.150 ;
        RECT 29.230 -7.790 31.910 -7.160 ;
        RECT 29.230 -7.820 31.260 -7.790 ;
    END
  END DIG04
  PIN DIG03
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 40.830 22.380 41.290 22.470 ;
        RECT 40.520 22.210 41.290 22.380 ;
        RECT 31.450 21.860 31.840 21.970 ;
        RECT 40.520 21.920 40.690 22.210 ;
        RECT 40.830 22.150 41.290 22.210 ;
        RECT 40.520 21.860 40.680 21.920 ;
        RECT 31.450 21.700 40.680 21.860 ;
        RECT 31.450 21.690 40.330 21.700 ;
        RECT 31.450 21.590 31.840 21.690 ;
        RECT 31.430 -6.530 31.920 -6.330 ;
        RECT 25.820 -6.550 31.920 -6.530 ;
        RECT 25.250 -6.830 31.920 -6.550 ;
        RECT 25.250 -6.930 31.830 -6.830 ;
        RECT 25.250 -7.160 27.230 -6.930 ;
        RECT 25.230 -7.820 27.260 -7.160 ;
    END
  END DIG03
  PIN DIG02
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 40.830 20.570 41.290 20.720 ;
        RECT 40.440 20.400 41.290 20.570 ;
        RECT 40.440 20.360 40.610 20.400 ;
        RECT 30.840 20.320 31.210 20.330 ;
        RECT 40.440 20.320 40.600 20.360 ;
        RECT 30.840 20.150 40.600 20.320 ;
        RECT 30.840 19.940 31.210 20.150 ;
        RECT 30.750 -5.720 31.290 -5.650 ;
        RECT 21.320 -6.150 31.290 -5.720 ;
        RECT 21.320 -7.160 23.300 -6.150 ;
        RECT 21.270 -7.820 23.300 -7.160 ;
    END
  END DIG02
  PIN DIG01
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 30.150 18.780 30.540 18.880 ;
        RECT 40.830 18.850 41.290 18.970 ;
        RECT 40.350 18.780 41.290 18.850 ;
        RECT 30.150 18.680 41.290 18.780 ;
        RECT 30.150 18.610 40.640 18.680 ;
        RECT 40.830 18.650 41.290 18.680 ;
        RECT 30.150 18.510 30.540 18.610 ;
        RECT 40.470 18.590 40.640 18.610 ;
        RECT 30.100 -4.880 30.640 -4.840 ;
        RECT 17.270 -4.920 30.640 -4.880 ;
        RECT 17.220 -5.310 30.640 -4.920 ;
        RECT 17.220 -7.190 19.230 -5.310 ;
        RECT 30.100 -5.340 30.640 -5.310 ;
        RECT 17.200 -7.850 19.230 -7.190 ;
    END
  END DIG01
  PIN CAP2    
    ANTENNAGATEAREA 6.526000 ;
    ANTENNADIFFAREA 0.336400 ;
    PORT
      LAYER met2 ;
        RECT 27.340 51.290 27.660 51.300 ;
        RECT 91.770 51.290 92.300 51.320 ;
        RECT 27.340 51.060 92.300 51.290 ;
        RECT 27.340 51.000 27.660 51.060 ;
        RECT 91.770 50.710 92.300 51.060 ;
        RECT 91.620 14.820 92.220 14.870 ;
        RECT 118.030 14.820 120.130 15.760 ;
        RECT 91.620 14.350 120.130 14.820 ;
        RECT 91.620 14.310 92.220 14.350 ;
        RECT 118.030 13.680 120.130 14.350 ;
        RECT 118.050 13.670 118.820 13.680 ;
        RECT 67.370 10.620 67.970 11.110 ;
        RECT 67.360 10.290 67.970 10.620 ;
        RECT 67.250 6.470 67.770 6.490 ;
        RECT 91.740 6.470 92.300 6.480 ;
        RECT 67.250 6.010 92.390 6.470 ;
        RECT 67.250 5.960 67.780 6.010 ;
        RECT 67.250 5.910 67.770 5.960 ;
    END
  END CAP2    
  PIN GENERALGATE01   
    ANTENNAGATEAREA 8.556000 ;
    ANTENNADIFFAREA 0.859400 ;
    PORT
      LAYER nwell ;
        RECT 28.530 61.660 31.240 61.700 ;
        RECT 28.520 60.010 31.240 61.660 ;
      LAYER met3 ;
        RECT 79.410 46.940 79.860 47.690 ;
        RECT 79.410 40.780 79.780 46.940 ;
        RECT 79.410 40.450 79.900 40.780 ;
        RECT 79.460 40.290 79.900 40.450 ;
    END
  END GENERALGATE01   
  PIN GATEANDCAP1    
    ANTENNAGATEAREA 22.864000 ;
    ANTENNADIFFAREA 1.740800 ;
    PORT
      LAYER nwell ;
        RECT 28.530 58.670 31.240 58.710 ;
        RECT 28.520 56.010 31.240 58.670 ;
      LAYER met2 ;
        RECT 30.590 52.210 30.960 52.270 ;
        RECT 93.790 52.210 94.330 52.230 ;
        RECT 30.590 51.980 94.330 52.210 ;
        RECT 30.590 51.920 30.960 51.980 ;
        RECT 93.790 51.670 94.330 51.980 ;
        RECT 18.720 46.330 19.040 46.380 ;
        RECT 19.450 46.330 19.760 46.430 ;
        RECT 18.720 46.160 19.760 46.330 ;
        RECT 18.720 46.120 19.040 46.160 ;
        RECT 19.450 46.100 19.760 46.160 ;
        RECT 18.690 45.410 19.010 45.460 ;
        RECT 19.430 45.410 19.740 45.510 ;
        RECT 18.690 45.240 19.740 45.410 ;
        RECT 18.690 45.200 19.010 45.240 ;
        RECT 19.430 45.180 19.740 45.240 ;
        RECT 18.700 44.490 19.020 44.540 ;
        RECT 19.410 44.490 19.720 44.520 ;
        RECT 18.700 44.320 19.720 44.490 ;
        RECT 18.700 44.280 19.020 44.320 ;
        RECT 19.410 44.190 19.720 44.320 ;
        RECT 18.050 43.480 18.370 43.520 ;
        RECT 19.670 43.490 19.990 43.550 ;
        RECT 19.360 43.480 19.990 43.490 ;
        RECT 18.050 43.300 19.990 43.480 ;
        RECT 18.050 43.290 19.480 43.300 ;
        RECT 18.050 43.260 18.370 43.290 ;
        RECT 19.670 43.230 19.990 43.300 ;
        RECT 18.010 42.520 18.330 42.560 ;
        RECT 18.010 42.500 19.480 42.520 ;
        RECT 19.670 42.500 19.990 42.560 ;
        RECT 18.010 42.330 19.990 42.500 ;
        RECT 18.010 42.300 18.330 42.330 ;
        RECT 19.360 42.310 19.990 42.330 ;
        RECT 19.670 42.240 19.990 42.310 ;
        RECT 18.050 41.560 18.370 41.600 ;
        RECT 18.050 41.510 19.480 41.560 ;
        RECT 19.670 41.510 19.990 41.570 ;
        RECT 18.050 41.370 19.990 41.510 ;
        RECT 18.050 41.340 18.370 41.370 ;
        RECT 19.360 41.320 19.990 41.370 ;
        RECT 19.670 41.250 19.990 41.320 ;
        RECT 18.010 26.530 18.320 26.550 ;
        RECT 18.670 26.530 18.980 26.550 ;
        RECT 18.010 26.060 25.330 26.530 ;
        RECT 18.010 26.040 18.320 26.060 ;
        RECT 18.670 26.040 18.980 26.060 ;
        RECT 24.860 25.380 25.330 26.060 ;
        RECT 117.630 25.380 118.530 26.350 ;
        RECT 16.680 25.250 16.940 25.320 ;
        RECT 18.730 25.250 19.050 25.270 ;
        RECT 20.490 25.250 20.820 25.290 ;
        RECT 16.680 25.060 20.820 25.250 ;
        RECT 16.680 25.000 16.940 25.060 ;
        RECT 18.730 25.010 19.050 25.060 ;
        RECT 20.490 25.020 20.820 25.060 ;
        RECT 24.860 24.910 118.530 25.380 ;
        RECT 16.130 24.850 16.450 24.890 ;
        RECT 18.070 24.850 18.390 24.910 ;
        RECT 20.990 24.850 21.310 24.890 ;
        RECT 16.130 24.660 21.310 24.850 ;
        RECT 93.790 24.790 94.360 24.910 ;
        RECT 16.130 24.630 16.450 24.660 ;
        RECT 18.070 24.650 18.390 24.660 ;
        RECT 20.990 24.630 21.310 24.660 ;
        RECT 117.630 24.260 118.530 24.910 ;
        RECT 17.150 22.500 17.470 22.520 ;
        RECT 16.930 22.280 17.470 22.500 ;
        RECT 17.150 22.260 17.470 22.280 ;
        RECT 19.900 21.920 20.220 22.040 ;
        RECT 16.930 21.720 20.220 21.920 ;
        RECT 16.930 21.710 19.910 21.720 ;
        RECT 16.930 21.500 19.910 21.520 ;
        RECT 16.930 21.310 20.230 21.500 ;
        RECT 19.910 21.180 20.230 21.310 ;
        RECT 16.160 20.980 16.450 20.990 ;
        RECT 16.150 20.960 16.470 20.980 ;
        RECT 17.150 20.960 17.470 20.970 ;
        RECT 16.150 20.740 17.470 20.960 ;
        RECT 16.150 20.720 16.470 20.740 ;
        RECT 16.160 20.700 16.450 20.720 ;
        RECT 17.150 20.710 17.470 20.740 ;
        RECT 18.830 13.830 19.440 14.160 ;
        RECT 18.840 13.340 19.440 13.830 ;
        RECT 57.560 10.590 58.160 11.080 ;
        RECT 57.550 10.260 58.160 10.590 ;
        RECT 57.370 7.860 94.450 8.320 ;
        RECT 57.440 7.760 57.960 7.860 ;
        RECT 93.800 7.800 94.360 7.860 ;
        RECT 18.870 6.590 19.480 6.610 ;
        RECT 18.870 6.280 21.220 6.590 ;
        RECT 18.880 6.250 21.220 6.280 ;
        RECT 18.880 6.010 21.260 6.250 ;
        RECT 18.880 5.990 21.220 6.010 ;
        RECT 18.880 5.790 19.480 5.990 ;
        RECT 20.250 5.920 20.910 5.990 ;
        RECT 20.280 5.910 20.880 5.920 ;
    END
  END GATEANDCAP1    
  PIN GENERALGATE02
    ANTENNAGATEAREA 8.556000 ;
    ANTENNADIFFAREA 0.974100 ;
    PORT
      LAYER met3 ;
        RECT 80.450 46.930 80.900 47.680 ;
        RECT 80.530 44.290 80.900 46.930 ;
        RECT 80.530 43.690 80.970 44.290 ;
        RECT 80.530 38.580 80.900 43.690 ;
        RECT 80.520 37.710 80.990 38.580 ;
    END
  END GENERALGATE02
  PIN OUTPUTTA1    
    ANTENNAGATEAREA 0.477400 ;
    PORT
      LAYER met2 ;
        RECT 8.730 57.790 9.040 58.020 ;
        RECT 5.640 57.690 9.040 57.790 ;
        RECT 5.640 57.560 9.020 57.690 ;
        RECT 5.640 57.530 5.960 57.560 ;
        RECT 115.050 55.250 115.820 55.400 ;
        RECT 5.560 54.830 115.820 55.250 ;
        RECT 115.050 54.690 115.820 54.830 ;
        RECT 114.860 35.490 115.640 35.640 ;
        RECT 117.600 35.490 118.500 36.410 ;
        RECT 114.860 35.020 118.500 35.490 ;
        RECT 114.860 34.870 115.640 35.020 ;
        RECT 117.600 34.320 118.500 35.020 ;
    END
  END OUTPUTTA1    
  PIN GATENFET1   
    ANTENNADIFFAREA 0.849600 ;
    PORT
      LAYER met2 ;
        RECT 110.000 43.100 110.320 43.140 ;
        RECT 111.010 43.100 111.330 43.130 ;
        RECT 109.950 42.900 113.720 43.100 ;
        RECT 110.000 42.880 110.320 42.900 ;
        RECT 111.010 42.870 111.330 42.900 ;
        RECT 112.000 42.820 113.710 42.900 ;
        RECT 110.000 42.370 110.320 42.390 ;
        RECT 111.010 42.370 111.330 42.400 ;
        RECT 113.510 42.370 113.710 42.820 ;
        RECT 109.950 42.170 113.710 42.370 ;
        RECT 110.000 42.130 110.320 42.170 ;
        RECT 111.010 42.140 111.330 42.170 ;
        RECT 113.510 41.120 113.710 42.170 ;
        RECT 117.600 41.120 118.500 41.790 ;
        RECT 113.510 40.690 118.500 41.120 ;
        RECT 113.510 40.000 113.710 40.690 ;
        RECT 110.000 39.900 110.320 39.940 ;
        RECT 111.010 39.900 111.330 39.930 ;
        RECT 112.000 39.900 113.710 40.000 ;
        RECT 109.950 39.700 113.710 39.900 ;
        RECT 117.600 39.700 118.500 40.690 ;
        RECT 110.000 39.680 110.320 39.700 ;
        RECT 111.010 39.670 111.330 39.700 ;
        RECT 113.510 39.350 113.710 39.700 ;
        RECT 110.000 39.170 110.320 39.190 ;
        RECT 111.010 39.170 111.330 39.200 ;
        RECT 112.000 39.170 113.710 39.350 ;
        RECT 109.950 39.030 113.710 39.170 ;
        RECT 109.950 38.970 113.700 39.030 ;
        RECT 110.000 38.930 110.320 38.970 ;
        RECT 111.010 38.940 111.330 38.970 ;
    END
  END GATENFET1   
  PIN DACOUTPUT  
    ANTENNADIFFAREA 3.264300 ;
    PORT
      LAYER met2 ;
        RECT 118.130 46.520 118.490 46.530 ;
        RECT 104.280 46.340 104.580 46.360 ;
        RECT 117.570 46.340 118.490 46.520 ;
        RECT 104.270 46.240 118.490 46.340 ;
        RECT 104.270 45.920 118.530 46.240 ;
        RECT 104.280 45.900 104.580 45.920 ;
        RECT 117.570 45.580 118.530 45.920 ;
        RECT 117.630 44.150 118.530 45.580 ;
    END
  END DACOUTPUT  
  PIN DRAINOUT
    ANTENNADIFFAREA 2.539200 ;
    PORT
      LAYER met2 ;
        RECT 89.290 48.650 89.720 48.670 ;
        RECT 117.640 48.650 118.500 50.630 ;
        RECT 89.290 48.530 118.500 48.650 ;
        RECT 89.290 48.280 118.390 48.530 ;
        RECT 89.290 48.250 89.700 48.280 ;
        RECT 51.630 26.390 51.940 26.410 ;
        RECT 89.270 26.390 89.720 26.420 ;
        RECT 51.630 25.980 89.720 26.390 ;
        RECT 51.630 25.960 51.940 25.980 ;
        RECT 89.270 25.960 89.720 25.980 ;
    END
  END DRAINOUT
  PIN ROWTERM2
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT 88.410 53.720 88.830 53.740 ;
        RECT 117.640 53.720 118.500 55.020 ;
        RECT 88.410 53.350 118.500 53.720 ;
        RECT 88.410 53.330 88.830 53.350 ;
        RECT 117.640 52.920 118.500 53.350 ;
        RECT 88.350 31.500 88.790 31.620 ;
        RECT 88.220 31.320 88.790 31.500 ;
        RECT 59.770 31.160 60.080 31.290 ;
        RECT 75.260 31.160 75.570 31.290 ;
        RECT 88.340 31.220 88.790 31.320 ;
        RECT 88.340 31.160 88.740 31.220 ;
        RECT 57.610 30.980 88.740 31.160 ;
        RECT 59.770 30.960 60.080 30.980 ;
        RECT 75.260 30.960 75.570 30.980 ;
    END
  END ROWTERM2
  PIN COLUMN2
    ANTENNAGATEAREA 1.620000 ;
    ANTENNADIFFAREA 0.640800 ;
    PORT
      LAYER met2 ;
        RECT 87.630 58.430 88.070 58.450 ;
        RECT 117.670 58.430 118.530 59.110 ;
        RECT 87.630 58.060 118.530 58.430 ;
        RECT 87.630 58.040 88.070 58.060 ;
        RECT 117.670 57.010 118.530 58.060 ;
        RECT 46.840 50.270 47.160 50.280 ;
        RECT 46.830 50.260 47.160 50.270 ;
        RECT 47.870 50.260 48.190 50.310 ;
        RECT 46.830 50.060 52.150 50.260 ;
        RECT 46.830 50.010 47.160 50.060 ;
        RECT 47.870 50.050 48.190 50.060 ;
        RECT 46.840 49.990 47.160 50.010 ;
        RECT 51.950 49.560 52.150 50.060 ;
        RECT 77.970 49.560 78.280 49.620 ;
        RECT 51.950 49.360 78.280 49.560 ;
        RECT 77.970 49.300 78.280 49.360 ;
        RECT 87.610 33.870 88.040 33.950 ;
        RECT 76.350 33.610 88.040 33.870 ;
        RECT 76.350 33.600 76.670 33.610 ;
        RECT 87.610 33.540 88.040 33.610 ;
    END
  END COLUMN2
  PIN COLUMN1
    ANTENNAGATEAREA 1.620000 ;
    ANTENNADIFFAREA 0.640800 ;
    PORT
      LAYER met2 ;
        RECT 86.800 61.890 87.260 61.910 ;
        RECT 117.670 61.890 118.530 63.240 ;
        RECT 86.800 61.520 118.530 61.890 ;
        RECT 86.800 61.500 87.260 61.520 ;
        RECT 117.670 61.140 118.530 61.520 ;
        RECT 56.900 49.090 57.220 49.140 ;
        RECT 51.900 48.890 57.270 49.090 ;
        RECT 46.840 48.520 47.160 48.530 ;
        RECT 46.830 48.510 47.160 48.520 ;
        RECT 47.870 48.510 48.190 48.560 ;
        RECT 51.900 48.510 52.100 48.890 ;
        RECT 56.900 48.880 57.220 48.890 ;
        RECT 46.830 48.310 52.100 48.510 ;
        RECT 46.830 48.260 47.160 48.310 ;
        RECT 47.870 48.300 48.190 48.310 ;
        RECT 46.840 48.240 47.160 48.260 ;
        RECT 59.010 34.470 59.330 34.480 ;
        RECT 86.820 34.470 87.280 34.540 ;
        RECT 59.010 34.190 87.280 34.470 ;
        RECT 59.010 34.140 59.330 34.190 ;
        RECT 86.820 34.130 87.280 34.190 ;
    END
  END COLUMN1
  PIN GATE2
    ANTENNADIFFAREA 6.691500 ;
    PORT
      LAYER nwell ;
        RECT 71.400 44.420 74.120 46.070 ;
        RECT 71.400 44.380 74.110 44.420 ;
        RECT 71.400 43.050 74.110 43.090 ;
        RECT 71.400 41.400 74.120 43.050 ;
        RECT 71.400 38.390 74.120 40.040 ;
        RECT 71.400 38.350 74.110 38.390 ;
        RECT 71.400 37.020 74.110 37.060 ;
        RECT 71.400 35.370 74.120 37.020 ;
        RECT 71.410 26.760 73.640 33.250 ;
      LAYER met2 ;
        RECT 71.660 50.130 71.940 50.150 ;
        RECT 71.640 50.100 71.960 50.130 ;
        RECT 103.780 50.100 105.120 50.640 ;
        RECT 71.640 49.890 105.120 50.100 ;
        RECT 71.640 49.870 71.960 49.890 ;
        RECT 71.660 49.850 71.940 49.870 ;
        RECT 103.780 49.360 105.120 49.890 ;
    END
  END GATE2
  PIN DRAININJECT
    ANTENNADIFFAREA 0.113400 ;
    PORT
      LAYER met2 ;
        RECT 47.180 60.000 47.630 60.020 ;
        RECT 47.170 59.940 47.650 60.000 ;
        RECT 24.780 59.800 47.650 59.940 ;
        RECT 24.760 59.640 47.650 59.800 ;
        RECT 24.760 59.480 25.080 59.640 ;
        RECT 47.170 59.580 47.650 59.640 ;
        RECT 47.180 59.560 47.630 59.580 ;
        RECT 24.760 59.470 25.070 59.480 ;
    END
  END DRAININJECT
  PIN VTUN
    ANTENNADIFFAREA 17.387499 ;
    PORT
      LAYER nwell ;
        RECT 33.720 59.960 35.940 61.650 ;
        RECT 65.980 46.060 69.370 46.810 ;
        RECT 65.970 42.490 69.380 46.060 ;
        RECT 65.970 41.150 69.370 42.490 ;
        RECT 65.980 40.030 69.370 41.150 ;
        RECT 65.980 36.460 69.380 40.030 ;
        RECT 65.990 34.740 69.370 36.460 ;
        RECT 65.950 26.760 69.390 33.250 ;
        RECT 65.980 17.430 67.710 23.930 ;
      LAYER met2 ;
        RECT 43.330 59.240 43.780 59.260 ;
        RECT 43.320 59.230 43.800 59.240 ;
        RECT 66.940 59.230 68.360 59.270 ;
        RECT 43.320 58.830 68.410 59.230 ;
        RECT 43.320 58.820 43.800 58.830 ;
        RECT 43.330 58.800 43.780 58.820 ;
        RECT 66.940 58.790 68.360 58.830 ;
    END
  END VTUN
  PIN VREFCHAR
    ANTENNAGATEAREA 6.711000 ;
    PORT
      LAYER met2 ;
        RECT 2.950 62.460 3.630 63.680 ;
        RECT 4.180 62.460 4.630 62.560 ;
        RECT 2.950 62.230 4.630 62.460 ;
        RECT 2.950 61.360 3.630 62.230 ;
        RECT 4.180 62.130 4.630 62.230 ;
        RECT 9.150 59.710 9.470 60.030 ;
        RECT 4.280 58.660 4.710 59.130 ;
        RECT 9.170 58.670 9.440 59.710 ;
        RECT 6.650 58.660 9.440 58.670 ;
        RECT 4.280 58.650 9.440 58.660 ;
        RECT 4.370 58.440 9.440 58.650 ;
        RECT 4.370 58.430 8.920 58.440 ;
        RECT 73.110 10.610 73.710 11.100 ;
        RECT 73.100 10.280 73.710 10.610 ;
        RECT 4.110 0.400 4.610 0.510 ;
        RECT 73.080 0.430 73.470 0.440 ;
        RECT 73.070 0.400 73.470 0.430 ;
        RECT 4.110 0.120 73.470 0.400 ;
        RECT 4.110 0.040 4.610 0.120 ;
        RECT 73.070 0.100 73.470 0.120 ;
        RECT 73.080 0.090 73.470 0.100 ;
    END
  END VREFCHAR
  PIN CHAROUTPUT
    ANTENNADIFFAREA 0.359600 ;
    PORT
      LAYER met2 ;
        RECT 2.950 58.270 3.630 59.150 ;
        RECT 2.950 58.240 6.610 58.270 ;
        RECT 2.950 57.980 6.910 58.240 ;
        RECT 2.950 57.950 6.610 57.980 ;
        RECT 2.950 56.830 3.630 57.950 ;
    END
  END CHAROUTPUT
  PIN LARGECAPACITOR
    ANTENNADIFFAREA 6.079600 ;
    PORT
      LAYER nwell ;
        RECT 11.700 57.080 21.390 61.680 ;
        RECT 11.100 55.690 21.390 57.080 ;
      LAYER met2 ;
        RECT 2.500 54.010 3.180 54.680 ;
        RECT 11.420 54.010 11.890 54.030 ;
        RECT 2.500 53.430 11.890 54.010 ;
        RECT 2.500 53.190 3.220 53.430 ;
        RECT 11.420 53.410 11.890 53.430 ;
        RECT 2.500 52.360 3.180 53.190 ;
    END
  END LARGECAPACITOR
  PIN DRAIN6N
    ANTENNADIFFAREA 4.231200 ;
    PORT
      LAYER met2 ;
        RECT 16.620 13.720 16.930 13.730 ;
        RECT 17.710 13.720 18.020 13.730 ;
        RECT 15.300 13.710 18.020 13.720 ;
        RECT 15.070 13.400 18.020 13.710 ;
        RECT 15.070 13.390 18.010 13.400 ;
        RECT 15.070 10.950 15.420 13.390 ;
        RECT 15.070 10.620 18.020 10.950 ;
        RECT 15.070 9.750 15.420 10.620 ;
        RECT 15.070 9.620 15.450 9.750 ;
        RECT 13.790 9.600 14.160 9.610 ;
        RECT 15.070 9.600 15.820 9.620 ;
        RECT 12.470 9.580 15.820 9.600 ;
        RECT 16.620 9.580 16.930 9.600 ;
        RECT 2.900 8.780 4.170 9.480 ;
        RECT 12.470 9.280 18.020 9.580 ;
        RECT 12.470 9.220 15.080 9.280 ;
        RECT 16.620 9.270 16.930 9.280 ;
        RECT 17.710 9.250 18.020 9.280 ;
        RECT 12.470 8.780 12.850 9.220 ;
        RECT 13.790 9.200 14.160 9.220 ;
        RECT 2.900 8.400 12.850 8.780 ;
        RECT 2.900 7.600 4.170 8.400 ;
    END
  END DRAIN6N
  PIN DRAIN6P
    ANTENNADIFFAREA 4.317200 ;
    PORT
      LAYER met2 ;
        RECT 16.660 6.170 16.970 6.180 ;
        RECT 17.750 6.170 18.060 6.180 ;
        RECT 15.340 6.160 18.060 6.170 ;
        RECT 15.110 5.850 18.060 6.160 ;
        RECT 15.110 5.840 18.050 5.850 ;
        RECT 2.900 3.550 4.170 4.460 ;
        RECT 2.900 3.170 12.870 3.550 ;
        RECT 2.900 2.580 4.170 3.170 ;
        RECT 12.490 2.320 12.870 3.170 ;
        RECT 15.110 3.400 15.460 5.840 ;
        RECT 15.110 3.070 18.060 3.400 ;
        RECT 13.790 2.320 14.160 2.330 ;
        RECT 15.110 2.320 15.460 3.070 ;
        RECT 12.490 2.200 15.460 2.320 ;
        RECT 12.490 2.070 15.490 2.200 ;
        RECT 12.490 2.030 15.860 2.070 ;
        RECT 16.660 2.030 16.970 2.050 ;
        RECT 12.490 1.940 18.060 2.030 ;
        RECT 13.790 1.920 14.160 1.940 ;
        RECT 15.110 1.730 18.060 1.940 ;
        RECT 16.660 1.720 16.970 1.730 ;
        RECT 17.750 1.700 18.060 1.730 ;
    END
  END DRAIN6P
  PIN DRAIN5P
    ANTENNADIFFAREA 0.727900 ;
    PORT
      LAYER met2 ;
        RECT 12.060 19.230 12.470 19.250 ;
        RECT 13.830 19.230 15.820 19.250 ;
        RECT 12.060 19.190 15.820 19.230 ;
        RECT 18.800 19.190 19.110 19.240 ;
        RECT 12.060 18.970 19.110 19.190 ;
        RECT 12.060 18.860 14.210 18.970 ;
        RECT 18.800 18.910 19.110 18.970 ;
        RECT 12.060 18.840 12.470 18.860 ;
        RECT 13.830 18.840 14.200 18.860 ;
        RECT 2.840 12.990 4.110 13.770 ;
        RECT 12.070 12.990 12.480 13.010 ;
        RECT 2.840 12.620 12.480 12.990 ;
        RECT 2.840 11.890 4.110 12.620 ;
        RECT 12.070 12.600 12.480 12.620 ;
    END
  END DRAIN5P
  PIN DARIN4P
    ANTENNADIFFAREA 0.727900 ;
    PORT
      LAYER met2 ;
        RECT 2.900 22.240 4.170 23.010 ;
        RECT 2.900 21.870 8.890 22.240 ;
        RECT 2.900 21.130 4.170 21.870 ;
        RECT 8.520 20.210 8.890 21.870 ;
        RECT 8.520 20.030 14.470 20.210 ;
        RECT 8.520 19.960 14.540 20.030 ;
        RECT 15.930 19.960 17.200 19.970 ;
        RECT 17.630 19.960 17.940 20.020 ;
        RECT 8.520 19.840 17.940 19.960 ;
        RECT 13.830 19.800 17.940 19.840 ;
        RECT 14.190 19.750 17.940 19.800 ;
        RECT 17.630 19.690 17.940 19.750 ;
    END
  END DARIN4P
  PIN DRAIN5N
    ANTENNADIFFAREA 0.688800 ;
    PORT
      LAYER met2 ;
        RECT 6.830 23.890 7.600 24.080 ;
        RECT 13.830 23.890 14.220 23.910 ;
        RECT 6.830 23.850 14.220 23.890 ;
        RECT 17.600 23.850 17.910 23.900 ;
        RECT 6.830 23.640 17.910 23.850 ;
        RECT 6.830 23.520 14.210 23.640 ;
        RECT 17.600 23.570 17.910 23.640 ;
        RECT 6.830 23.340 7.600 23.520 ;
        RECT 13.830 23.500 14.200 23.520 ;
        RECT 2.900 18.100 4.170 18.920 ;
        RECT 6.830 18.100 7.630 18.240 ;
        RECT 2.900 17.600 7.630 18.100 ;
        RECT 2.900 17.040 4.170 17.600 ;
        RECT 6.830 17.470 7.630 17.600 ;
    END
  END DRAIN5N
  PIN DRAIN4N
    ANTENNADIFFAREA 0.688800 ;
    PORT
      LAYER met2 ;
        RECT 2.840 26.270 4.110 27.110 ;
        RECT 2.840 25.900 12.540 26.270 ;
        RECT 2.840 25.230 4.110 25.900 ;
        RECT 12.170 24.550 12.540 25.900 ;
        RECT 12.170 24.540 14.200 24.550 ;
        RECT 12.170 24.360 14.420 24.540 ;
        RECT 12.170 24.300 15.820 24.360 ;
        RECT 18.820 24.300 19.130 24.340 ;
        RECT 12.170 24.180 19.130 24.300 ;
        RECT 13.830 24.140 19.130 24.180 ;
        RECT 14.200 24.080 19.130 24.140 ;
        RECT 18.820 24.010 19.130 24.080 ;
    END
  END DRAIN4N
  PIN DRAIN3P
    ANTENNADIFFAREA 0.117600 ;
    PORT
      LAYER met2 ;
        RECT 13.830 41.930 19.480 41.980 ;
        RECT 19.700 41.930 20.010 42.040 ;
        RECT 13.830 41.790 20.010 41.930 ;
        RECT 2.900 30.420 4.170 31.330 ;
        RECT 13.830 30.420 14.200 41.790 ;
        RECT 19.360 41.740 20.010 41.790 ;
        RECT 19.700 41.710 20.010 41.740 ;
        RECT 2.900 30.050 14.200 30.420 ;
        RECT 2.900 29.450 4.170 30.050 ;
    END
  END DRAIN3P
  PIN DRAIN2P
    ANTENNADIFFAREA 0.235200 ;
    PORT
      LAYER met2 ;
        RECT 19.700 43.910 20.010 44.020 ;
        RECT 19.360 43.900 20.010 43.910 ;
        RECT 12.990 43.880 20.010 43.900 ;
        RECT 12.700 43.720 20.010 43.880 ;
        RECT 12.700 43.710 19.480 43.720 ;
        RECT 12.700 43.530 14.200 43.710 ;
        RECT 19.700 43.690 20.010 43.720 ;
        RECT 12.700 42.940 13.360 43.530 ;
        RECT 13.830 43.490 14.200 43.530 ;
        RECT 12.700 42.920 19.480 42.940 ;
        RECT 19.700 42.920 20.010 43.030 ;
        RECT 12.700 42.750 20.010 42.920 ;
        RECT 12.700 42.570 14.200 42.750 ;
        RECT 19.360 42.730 20.010 42.750 ;
        RECT 19.700 42.700 20.010 42.730 ;
        RECT 12.700 42.560 13.370 42.570 ;
        RECT 12.700 42.520 13.360 42.560 ;
        RECT 13.830 42.530 14.200 42.570 ;
        RECT 2.840 35.260 4.110 36.150 ;
        RECT 12.700 35.260 13.070 42.520 ;
        RECT 2.840 34.890 13.070 35.260 ;
        RECT 2.840 34.270 4.110 34.890 ;
    END
  END DRAIN2P
  PIN DRAIN3N
    ANTENNADIFFAREA 0.390600 ;
    PORT
      LAYER met2 ;
        RECT 13.830 46.970 14.200 46.980 ;
        RECT 12.040 46.740 14.200 46.970 ;
        RECT 19.880 46.840 20.190 46.930 ;
        RECT 19.290 46.740 20.190 46.840 ;
        RECT 12.040 46.670 20.190 46.740 ;
        RECT 12.040 46.610 19.460 46.670 ;
        RECT 12.040 45.910 12.660 46.610 ;
        RECT 13.830 46.570 19.460 46.610 ;
        RECT 19.880 46.600 20.190 46.670 ;
        RECT 13.830 45.910 14.200 45.950 ;
        RECT 11.510 45.820 14.200 45.910 ;
        RECT 19.890 45.850 20.200 45.940 ;
        RECT 19.360 45.820 20.200 45.850 ;
        RECT 11.510 45.680 20.200 45.820 ;
        RECT 11.510 45.650 19.460 45.680 ;
        RECT 11.510 45.540 14.200 45.650 ;
        RECT 19.890 45.610 20.200 45.680 ;
        RECT 11.510 45.430 12.660 45.540 ;
        RECT 11.510 44.980 12.620 45.430 ;
        RECT 13.830 44.980 14.200 45.020 ;
        RECT 11.510 44.900 14.200 44.980 ;
        RECT 11.510 44.870 19.460 44.900 ;
        RECT 11.510 44.860 19.500 44.870 ;
        RECT 19.890 44.860 20.200 44.950 ;
        RECT 11.510 44.730 20.200 44.860 ;
        RECT 11.510 44.610 14.200 44.730 ;
        RECT 19.360 44.690 20.200 44.730 ;
        RECT 19.890 44.620 20.200 44.690 ;
        RECT 11.510 44.570 12.410 44.610 ;
        RECT 2.900 40.020 4.170 40.900 ;
        RECT 11.510 40.020 11.880 44.570 ;
        RECT 2.900 39.650 11.880 40.020 ;
        RECT 2.900 39.020 4.170 39.650 ;
    END
  END DRAIN3N
  PIN SOURCEN
    ANTENNADIFFAREA 5.999400 ;
    PORT
      LAYER met2 ;
        RECT 22.480 48.050 22.770 48.070 ;
        RECT 10.030 47.650 22.790 48.050 ;
        RECT 2.470 44.960 3.740 45.830 ;
        RECT 10.030 44.960 10.430 47.650 ;
        RECT 22.480 47.640 22.770 47.650 ;
        RECT 20.970 46.850 21.280 46.940 ;
        RECT 20.970 46.750 21.430 46.850 ;
        RECT 22.490 46.750 22.810 46.800 ;
        RECT 20.970 46.610 22.870 46.750 ;
        RECT 21.270 46.580 22.870 46.610 ;
        RECT 22.490 46.540 22.810 46.580 ;
        RECT 20.980 45.860 21.290 45.950 ;
        RECT 20.980 45.830 21.440 45.860 ;
        RECT 22.490 45.830 22.810 45.880 ;
        RECT 20.980 45.660 22.870 45.830 ;
        RECT 20.980 45.620 21.290 45.660 ;
        RECT 22.490 45.620 22.810 45.660 ;
        RECT 2.470 44.560 10.430 44.960 ;
        RECT 20.980 44.910 21.290 44.960 ;
        RECT 22.460 44.910 22.780 44.960 ;
        RECT 20.980 44.740 22.870 44.910 ;
        RECT 20.980 44.700 21.440 44.740 ;
        RECT 22.460 44.700 22.780 44.740 ;
        RECT 20.980 44.630 21.290 44.700 ;
        RECT 2.470 43.950 3.740 44.560 ;
        RECT 19.470 24.270 19.780 24.340 ;
        RECT 22.470 24.290 22.770 24.310 ;
        RECT 22.460 24.270 22.780 24.290 ;
        RECT 19.470 24.060 22.780 24.270 ;
        RECT 19.470 24.010 19.780 24.060 ;
        RECT 20.240 24.050 22.780 24.060 ;
        RECT 18.300 23.830 18.610 23.900 ;
        RECT 20.240 23.830 20.460 24.050 ;
        RECT 22.460 24.030 22.780 24.050 ;
        RECT 22.470 24.010 22.770 24.030 ;
        RECT 18.300 23.610 20.460 23.830 ;
        RECT 18.300 23.570 18.610 23.610 ;
        RECT 16.070 13.040 16.380 13.050 ;
        RECT 17.170 13.040 17.480 13.050 ;
        RECT 18.270 13.040 18.580 13.050 ;
        RECT 16.040 12.720 19.200 13.040 ;
        RECT 18.880 11.680 19.200 12.720 ;
        RECT 16.040 11.350 19.200 11.680 ;
        RECT 16.070 8.900 16.380 8.910 ;
        RECT 18.880 8.900 19.200 11.350 ;
        RECT 22.460 8.900 22.740 8.910 ;
        RECT 16.050 8.570 22.760 8.900 ;
        RECT 16.050 8.560 19.110 8.570 ;
        RECT 22.460 8.550 22.740 8.570 ;
    END
  END SOURCEN
  PIN SOURCEP
    ANTENNADIFFAREA 6.113200 ;
    PORT
      LAYER met2 ;
        RECT 2.180 48.860 3.450 50.320 ;
        RECT 13.530 48.860 13.830 48.870 ;
        RECT 23.120 48.860 23.410 48.880 ;
        RECT 2.180 48.470 23.440 48.860 ;
        RECT 2.180 48.440 3.450 48.470 ;
        RECT 23.120 48.450 23.410 48.470 ;
        RECT 21.000 43.840 21.310 43.920 ;
        RECT 23.100 43.840 23.420 43.870 ;
        RECT 21.000 43.640 23.520 43.840 ;
        RECT 21.000 43.590 21.310 43.640 ;
        RECT 23.100 43.610 23.420 43.640 ;
        RECT 21.000 42.880 21.310 42.930 ;
        RECT 23.110 42.880 23.430 42.910 ;
        RECT 21.000 42.680 23.520 42.880 ;
        RECT 21.000 42.600 21.310 42.680 ;
        RECT 23.110 42.650 23.430 42.680 ;
        RECT 21.000 41.920 21.310 41.940 ;
        RECT 23.100 41.920 23.420 41.950 ;
        RECT 21.000 41.720 23.520 41.920 ;
        RECT 21.000 41.610 21.310 41.720 ;
        RECT 23.100 41.690 23.420 41.720 ;
        RECT 18.320 19.940 18.630 20.010 ;
        RECT 23.110 19.960 23.400 19.980 ;
        RECT 18.320 19.930 20.460 19.940 ;
        RECT 23.100 19.930 23.420 19.960 ;
        RECT 18.320 19.730 23.420 19.930 ;
        RECT 18.320 19.680 18.630 19.730 ;
        RECT 20.250 19.720 23.420 19.730 ;
        RECT 19.510 19.110 19.820 19.180 ;
        RECT 20.250 19.110 20.460 19.720 ;
        RECT 23.100 19.700 23.420 19.720 ;
        RECT 23.110 19.680 23.400 19.700 ;
        RECT 19.510 18.900 20.460 19.110 ;
        RECT 19.510 18.850 19.820 18.900 ;
        RECT 16.110 5.490 16.420 5.500 ;
        RECT 17.210 5.490 17.520 5.500 ;
        RECT 18.310 5.490 18.620 5.500 ;
        RECT 16.080 5.170 19.240 5.490 ;
        RECT 18.920 4.130 19.240 5.170 ;
        RECT 16.080 3.800 19.240 4.130 ;
        RECT 16.110 1.350 16.420 1.360 ;
        RECT 18.920 1.350 19.240 3.800 ;
        RECT 23.040 1.350 23.350 1.370 ;
        RECT 16.090 1.010 23.350 1.350 ;
        RECT 23.040 0.990 23.350 1.010 ;
    END
  END SOURCEP
  PIN GATE1
    ANTENNADIFFAREA 0.434600 ;
    PORT
      LAYER met2 ;
        RECT 59.240 50.710 59.560 50.750 ;
        RECT 74.890 50.710 76.170 50.810 ;
        RECT 59.240 50.500 76.170 50.710 ;
        RECT 59.240 50.470 59.560 50.500 ;
    END
  END GATE1
  PIN VINJ
    ANTENNADIFFAREA 1.929800 ;
    PORT
      LAYER nwell ;
        RECT 6.090 58.170 8.830 61.670 ;
        RECT 22.970 55.670 26.970 61.660 ;
      LAYER met2 ;
        RECT 2.800 60.260 5.280 60.270 ;
        RECT 6.590 60.260 6.910 60.460 ;
        RECT 7.320 60.260 7.630 60.470 ;
        RECT 8.000 60.260 8.320 60.470 ;
        RECT 8.660 60.260 23.310 60.390 ;
        RECT 2.800 60.180 23.310 60.260 ;
        RECT 2.800 60.010 8.800 60.180 ;
        RECT 22.730 60.170 23.480 60.180 ;
        RECT 2.800 59.870 8.660 60.010 ;
        RECT 5.070 59.500 8.660 59.870 ;
        RECT 22.730 59.870 24.350 60.170 ;
        RECT 22.730 59.730 22.970 59.870 ;
        RECT 24.050 59.810 24.350 59.870 ;
        RECT 6.590 59.330 6.910 59.500 ;
        RECT 7.320 59.300 7.630 59.500 ;
        RECT 8.020 59.350 8.340 59.500 ;
        RECT 22.710 59.400 23.020 59.730 ;
        RECT 24.050 59.490 24.380 59.810 ;
        RECT 24.070 59.480 24.380 59.490 ;
    END
    PORT
      LAYER met2 ;
        RECT 2.500 51.860 3.010 51.980 ;
        RECT 2.500 51.570 5.600 51.860 ;
        RECT 3.010 51.560 5.600 51.570 ;
    END
    PORT
      LAYER nwell ;
        RECT 47.070 36.590 49.570 50.700 ;
        RECT 56.190 43.730 59.500 46.860 ;
        RECT 52.090 40.830 59.500 43.730 ;
        RECT 75.850 46.810 79.160 46.860 ;
        RECT 75.850 46.800 80.500 46.810 ;
        RECT 52.090 37.140 59.510 40.830 ;
        RECT 56.200 34.680 59.510 37.140 ;
        RECT 75.850 34.730 81.010 46.800 ;
        RECT 75.850 34.680 79.160 34.730 ;
        RECT 47.070 26.460 49.570 33.460 ;
        RECT 52.070 26.670 55.490 33.260 ;
        RECT 57.610 26.760 60.170 33.260 ;
        RECT 75.170 26.760 77.730 33.260 ;
        RECT 47.030 17.400 49.530 24.400 ;
        RECT 52.100 23.590 55.520 23.990 ;
        RECT 57.640 23.660 60.200 23.930 ;
        RECT 57.240 23.590 60.200 23.660 ;
        RECT 52.100 17.590 60.200 23.590 ;
        RECT 52.100 17.400 55.520 17.590 ;
        RECT 57.640 17.430 60.200 17.590 ;
      LAYER met2 ;
        RECT 48.840 57.620 49.340 57.650 ;
        RECT 54.560 57.620 55.060 57.650 ;
        RECT 48.840 57.210 79.000 57.620 ;
        RECT 48.990 57.180 79.000 57.210 ;
        RECT 56.390 46.670 56.710 46.790 ;
        RECT 78.660 46.670 78.980 46.790 ;
        RECT 56.390 46.490 78.980 46.670 ;
        RECT 77.770 43.950 78.090 44.210 ;
        RECT 77.810 43.930 78.990 43.950 ;
        RECT 77.810 43.670 79.030 43.930 ;
        RECT 77.810 43.610 78.990 43.670 ;
        RECT 77.770 43.600 78.990 43.610 ;
        RECT 77.770 43.350 78.090 43.600 ;
        RECT 56.440 40.610 56.760 40.730 ;
        RECT 78.640 40.610 78.960 40.730 ;
        RECT 56.440 40.430 78.960 40.610 ;
        RECT 77.770 37.920 78.090 38.180 ;
        RECT 77.810 37.900 78.990 37.920 ;
        RECT 77.810 37.640 79.030 37.900 ;
        RECT 77.810 37.580 78.990 37.640 ;
        RECT 77.770 37.570 78.990 37.580 ;
        RECT 77.770 37.320 78.090 37.570 ;
        RECT 57.810 32.980 77.550 33.160 ;
        RECT 57.810 32.840 58.230 32.980 ;
        RECT 77.210 32.850 77.550 32.980 ;
        RECT 48.920 17.050 49.250 17.070 ;
        RECT 48.910 16.970 49.260 17.050 ;
        RECT 54.660 16.970 54.980 17.030 ;
        RECT 48.910 16.810 54.980 16.970 ;
        RECT 48.910 16.740 49.260 16.810 ;
        RECT 54.660 16.760 54.980 16.810 ;
        RECT 48.300 15.970 48.740 15.980 ;
        RECT 2.980 15.960 48.740 15.970 ;
        RECT 2.980 15.550 48.760 15.960 ;
        RECT 41.450 15.540 41.930 15.550 ;
        RECT 48.280 15.540 48.760 15.550 ;
        RECT 48.300 15.530 48.740 15.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.380 57.140 57.110 64.010 ;
        RECT 56.540 46.790 56.710 57.140 ;
        RECT 56.390 46.490 56.710 46.790 ;
        RECT 56.550 46.160 56.710 46.490 ;
        RECT 56.550 45.610 56.820 46.160 ;
        RECT 56.540 45.560 56.820 45.610 ;
        RECT 56.540 45.470 56.710 45.560 ;
        RECT 56.550 42.100 56.710 45.470 ;
        RECT 56.540 42.010 56.710 42.100 ;
        RECT 56.540 41.960 56.820 42.010 ;
        RECT 56.550 41.410 56.820 41.960 ;
        RECT 56.550 40.780 56.710 41.410 ;
        RECT 56.440 40.730 56.720 40.780 ;
        RECT 56.440 40.450 56.760 40.730 ;
        RECT 56.440 40.130 56.720 40.450 ;
        RECT 56.440 39.530 56.830 40.130 ;
        RECT 56.440 35.980 56.720 39.530 ;
        RECT 56.440 35.380 56.830 35.980 ;
        RECT 56.440 33.900 56.720 35.380 ;
        RECT 56.440 33.620 58.160 33.900 ;
        RECT 57.960 33.390 58.160 33.620 ;
        RECT 57.970 33.130 58.130 33.390 ;
        RECT 57.820 32.990 58.130 33.130 ;
        RECT 57.810 32.840 58.130 32.990 ;
        RECT 57.970 32.550 58.130 32.840 ;
        RECT 57.970 32.000 58.240 32.550 ;
        RECT 57.960 31.950 58.240 32.000 ;
        RECT 57.960 31.860 58.130 31.950 ;
        RECT 57.970 31.390 58.130 31.860 ;
        RECT 57.960 31.300 58.130 31.390 ;
        RECT 57.960 31.250 58.240 31.300 ;
        RECT 57.970 30.700 58.240 31.250 ;
        RECT 57.970 29.310 58.130 30.700 ;
        RECT 57.970 28.760 58.240 29.310 ;
        RECT 57.960 28.710 58.240 28.760 ;
        RECT 57.960 28.620 58.130 28.710 ;
        RECT 57.970 28.160 58.130 28.620 ;
        RECT 57.960 28.070 58.130 28.160 ;
        RECT 57.960 28.020 58.240 28.070 ;
        RECT 57.970 27.470 58.240 28.020 ;
        RECT 57.970 26.770 58.160 27.470 ;
        RECT 58.000 23.220 58.160 26.770 ;
        RECT 58.000 22.670 58.270 23.220 ;
        RECT 57.990 22.620 58.270 22.670 ;
        RECT 57.990 22.530 58.160 22.620 ;
        RECT 58.000 22.080 58.160 22.530 ;
        RECT 57.990 21.990 58.160 22.080 ;
        RECT 57.990 21.940 58.270 21.990 ;
        RECT 58.000 21.390 58.270 21.940 ;
        RECT 58.000 19.980 58.160 21.390 ;
        RECT 58.000 19.430 58.270 19.980 ;
        RECT 57.990 19.380 58.270 19.430 ;
        RECT 57.990 19.290 58.160 19.380 ;
        RECT 58.000 18.830 58.160 19.290 ;
        RECT 57.990 18.740 58.160 18.830 ;
        RECT 57.990 18.690 58.270 18.740 ;
        RECT 58.000 18.140 58.270 18.690 ;
        RECT 58.000 17.440 58.160 18.140 ;
      LAYER via ;
        RECT 56.410 57.180 56.850 57.620 ;
        RECT 56.420 46.510 56.680 46.770 ;
        RECT 56.470 40.460 56.730 40.720 ;
        RECT 57.850 32.860 58.110 33.120 ;
    END
  END VINJ
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 7.300 56.620 7.610 56.830 ;
        RECT 8.730 56.620 9.040 56.850 ;
        RECT 4.950 56.460 9.870 56.620 ;
        RECT 3.140 56.290 9.870 56.460 ;
        RECT 3.140 56.240 9.880 56.290 ;
        RECT 3.140 56.130 9.900 56.240 ;
        RECT 3.140 56.060 5.410 56.130 ;
        RECT 3.140 55.860 3.540 56.060 ;
        RECT 6.510 55.920 6.820 56.130 ;
        RECT 7.440 55.920 7.750 56.130 ;
        RECT 8.140 55.920 8.450 56.130 ;
        RECT 8.880 55.950 9.900 56.130 ;
        RECT 21.990 55.950 22.300 56.070 ;
        RECT 31.850 55.950 32.160 56.090 ;
        RECT 8.880 55.920 32.160 55.950 ;
        RECT 2.790 55.460 3.540 55.860 ;
        RECT 8.900 55.760 32.160 55.920 ;
        RECT 8.900 55.740 32.130 55.760 ;
    END
    PORT
      LAYER met2 ;
        RECT 44.420 56.610 44.920 56.630 ;
        RECT 50.160 56.610 50.600 56.660 ;
        RECT 64.530 56.610 65.030 56.630 ;
        RECT 44.420 56.190 70.930 56.610 ;
        RECT 44.570 56.170 70.930 56.190 ;
        RECT 50.160 56.160 50.600 56.170 ;
        RECT 70.330 56.150 70.830 56.170 ;
        RECT 2.460 51.060 2.970 51.080 ;
        RECT 22.100 51.060 22.500 51.070 ;
        RECT 2.460 50.710 22.500 51.060 ;
        RECT 2.460 50.670 2.970 50.710 ;
        RECT 22.100 50.680 22.500 50.710 ;
        RECT 80.800 41.110 81.120 41.260 ;
        RECT 64.610 40.960 81.120 41.110 ;
        RECT 64.610 40.810 64.930 40.960 ;
        RECT 70.410 40.810 70.730 40.960 ;
        RECT 64.680 37.620 65.000 37.670 ;
        RECT 64.680 37.370 70.700 37.620 ;
        RECT 70.380 37.300 70.700 37.370 ;
        RECT 70.380 35.080 70.700 35.090 ;
        RECT 80.820 35.080 81.150 35.220 ;
        RECT 70.380 34.920 81.150 35.080 ;
        RECT 70.380 34.910 71.070 34.920 ;
        RECT 70.380 34.790 70.700 34.910 ;
        RECT 60.680 28.540 61.000 28.600 ;
        RECT 64.610 28.540 64.930 28.550 ;
        RECT 70.410 28.540 70.730 28.550 ;
        RECT 74.340 28.540 74.660 28.600 ;
        RECT 60.680 28.360 74.660 28.540 ;
        RECT 60.680 28.310 61.000 28.360 ;
        RECT 64.610 28.290 64.930 28.360 ;
        RECT 70.410 28.290 70.730 28.360 ;
        RECT 74.340 28.310 74.660 28.360 ;
        RECT 19.980 23.110 20.300 23.170 ;
        RECT 21.850 23.140 22.140 23.160 ;
        RECT 19.980 23.100 20.460 23.110 ;
        RECT 21.840 23.100 22.160 23.140 ;
        RECT 19.980 22.910 22.160 23.100 ;
        RECT 19.980 22.900 20.460 22.910 ;
        RECT 19.980 22.850 20.300 22.900 ;
        RECT 21.840 22.880 22.160 22.910 ;
        RECT 21.850 22.860 22.140 22.880 ;
        RECT 70.760 19.200 71.090 19.290 ;
        RECT 60.830 19.130 61.150 19.190 ;
        RECT 64.410 19.130 71.090 19.200 ;
        RECT 60.830 19.030 71.090 19.130 ;
        RECT 60.830 18.960 65.180 19.030 ;
        RECT 70.760 19.000 71.090 19.030 ;
        RECT 60.830 18.910 61.150 18.960 ;
        RECT 64.850 18.900 65.180 18.960 ;
        RECT 44.490 16.350 44.820 16.590 ;
        RECT 50.350 16.480 50.650 16.490 ;
        RECT 50.340 16.350 50.660 16.480 ;
        RECT 60.880 16.350 61.160 16.650 ;
        RECT 64.910 16.350 65.210 16.630 ;
        RECT 44.490 16.330 65.210 16.350 ;
        RECT 44.490 16.300 65.200 16.330 ;
        RECT 44.490 16.190 65.140 16.300 ;
        RECT 73.750 15.880 74.050 15.900 ;
        RECT 70.320 15.540 74.060 15.880 ;
        RECT 70.340 15.530 70.650 15.540 ;
        RECT 2.960 14.580 44.940 15.000 ;
        RECT 26.010 14.080 26.840 14.580 ;
        RECT 73.150 13.090 73.470 15.540 ;
        RECT 73.750 15.520 74.060 15.540 ;
        RECT 70.310 12.760 73.470 13.090 ;
        RECT 19.600 12.560 19.890 12.580 ;
        RECT 21.830 12.560 22.140 12.580 ;
        RECT 19.590 12.200 22.140 12.560 ;
        RECT 19.600 12.180 19.890 12.200 ;
        RECT 21.830 12.180 22.140 12.200 ;
        RECT 73.150 11.720 73.470 12.760 ;
        RECT 70.310 11.400 73.470 11.720 ;
        RECT 70.340 11.390 70.650 11.400 ;
        RECT 71.440 11.390 71.750 11.400 ;
        RECT 72.540 11.390 72.850 11.400 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.530 63.860 62.510 64.010 ;
        RECT 61.540 56.610 62.510 63.860 ;
        RECT 61.520 56.140 62.530 56.610 ;
      LAYER via ;
        RECT 61.550 56.180 62.500 56.590 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 19.360 44.180 21.390 44.190 ;
        RECT 19.360 41.090 21.930 44.180 ;
        RECT 41.430 36.590 43.200 50.700 ;
        RECT 83.010 34.730 84.290 46.810 ;
        RECT 107.560 37.830 110.320 44.240 ;
        RECT 41.430 26.460 43.200 33.460 ;
        RECT 17.530 21.260 19.900 21.460 ;
        RECT 17.530 19.290 20.460 21.260 ;
        RECT 17.530 18.590 19.900 19.290 ;
        RECT 41.390 17.400 43.160 24.400 ;
        RECT 59.410 16.150 67.250 16.160 ;
        RECT 57.400 16.130 67.250 16.150 ;
        RECT 49.600 10.460 67.250 16.130 ;
        RECT 49.600 10.430 57.440 10.460 ;
        RECT 104.390 9.810 110.040 9.980 ;
        RECT 14.840 0.740 18.760 6.440 ;
        RECT 104.390 -6.120 111.390 9.810 ;
        RECT 110.030 -6.130 111.390 -6.120 ;
      LAYER met2 ;
        RECT 41.670 53.400 41.970 53.460 ;
        RECT 82.990 53.400 83.290 53.430 ;
        RECT 41.670 53.170 83.360 53.400 ;
        RECT 41.670 53.140 41.970 53.170 ;
        RECT 82.990 53.090 83.290 53.170 ;
        RECT 83.200 47.630 83.670 47.690 ;
        RECT 108.100 47.640 108.390 47.650 ;
        RECT 108.100 47.630 108.400 47.640 ;
        RECT 118.630 47.630 119.080 47.650 ;
        RECT 83.200 47.200 119.090 47.630 ;
        RECT 108.100 47.190 108.400 47.200 ;
        RECT 108.100 47.170 108.390 47.190 ;
        RECT 19.960 20.500 20.280 20.550 ;
        RECT 21.420 20.500 21.740 20.550 ;
        RECT 19.960 20.290 21.740 20.500 ;
        RECT 19.960 20.230 20.280 20.290 ;
        RECT 21.420 20.250 21.740 20.290 ;
        RECT 97.860 17.310 98.420 17.380 ;
        RECT 110.580 17.310 111.260 17.370 ;
        RECT 118.110 17.310 118.770 17.950 ;
        RECT 97.860 16.900 118.770 17.310 ;
        RECT 97.860 16.850 98.420 16.900 ;
        RECT 110.580 16.840 111.260 16.900 ;
        RECT 118.110 16.800 118.770 16.900 ;
        RECT 60.110 15.170 60.420 15.200 ;
        RECT 61.200 15.170 61.510 15.180 ;
        RECT 65.150 15.170 65.460 15.180 ;
        RECT 66.240 15.170 66.550 15.200 ;
        RECT 50.300 15.140 50.610 15.170 ;
        RECT 51.390 15.140 51.700 15.150 ;
        RECT 55.340 15.140 55.650 15.150 ;
        RECT 56.430 15.140 56.740 15.170 ;
        RECT 50.300 14.840 53.250 15.140 ;
        RECT 51.390 14.820 51.700 14.840 ;
        RECT 52.500 14.800 53.250 14.840 ;
        RECT 52.870 14.670 53.250 14.800 ;
        RECT 52.900 13.800 53.250 14.670 ;
        RECT 50.300 13.470 53.250 13.800 ;
        RECT 52.900 11.030 53.250 13.470 ;
        RECT 50.310 11.020 53.250 11.030 ;
        RECT 50.300 10.710 53.250 11.020 ;
        RECT 53.790 14.840 56.740 15.140 ;
        RECT 60.110 14.870 63.060 15.170 ;
        RECT 61.200 14.850 61.510 14.870 ;
        RECT 53.790 14.800 54.540 14.840 ;
        RECT 55.340 14.820 55.650 14.840 ;
        RECT 62.310 14.830 63.060 14.870 ;
        RECT 53.790 14.670 54.170 14.800 ;
        RECT 62.680 14.700 63.060 14.830 ;
        RECT 53.790 13.800 54.140 14.670 ;
        RECT 62.710 13.830 63.060 14.700 ;
        RECT 53.790 13.470 56.740 13.800 ;
        RECT 60.110 13.500 63.060 13.830 ;
        RECT 53.790 11.030 54.140 13.470 ;
        RECT 62.710 11.060 63.060 13.500 ;
        RECT 60.120 11.050 63.060 11.060 ;
        RECT 53.790 11.020 56.730 11.030 ;
        RECT 53.790 10.710 56.740 11.020 ;
        RECT 60.110 10.740 63.060 11.050 ;
        RECT 63.600 14.870 66.550 15.170 ;
        RECT 63.600 14.830 64.350 14.870 ;
        RECT 65.150 14.850 65.460 14.870 ;
        RECT 63.600 14.700 63.980 14.830 ;
        RECT 63.600 13.830 63.950 14.700 ;
        RECT 63.600 13.500 66.550 13.830 ;
        RECT 63.600 11.060 63.950 13.500 ;
        RECT 63.600 11.050 66.540 11.060 ;
        RECT 63.600 10.740 66.550 11.050 ;
        RECT 60.110 10.730 62.830 10.740 ;
        RECT 63.830 10.730 66.550 10.740 ;
        RECT 60.110 10.720 60.420 10.730 ;
        RECT 61.200 10.720 61.510 10.730 ;
        RECT 65.150 10.720 65.460 10.730 ;
        RECT 66.240 10.720 66.550 10.730 ;
        RECT 50.300 10.700 53.020 10.710 ;
        RECT 54.020 10.700 56.740 10.710 ;
        RECT 50.300 10.690 50.610 10.700 ;
        RECT 51.390 10.690 51.700 10.700 ;
        RECT 55.340 10.690 55.650 10.700 ;
        RECT 56.430 10.690 56.740 10.700 ;
        RECT 52.990 10.020 63.890 10.050 ;
        RECT 52.980 9.770 63.890 10.020 ;
        RECT 52.980 9.740 53.320 9.770 ;
        RECT 53.720 9.760 54.060 9.770 ;
        RECT 62.790 9.740 63.130 9.770 ;
        RECT 110.040 7.320 110.330 7.380 ;
        RECT 15.040 7.220 15.390 7.250 ;
        RECT 21.420 7.240 21.750 7.280 ;
        RECT 21.410 7.220 21.760 7.240 ;
        RECT 15.040 6.960 25.070 7.220 ;
        RECT 109.870 7.010 110.330 7.320 ;
        RECT 110.040 6.970 110.330 7.010 ;
        RECT 15.080 6.930 25.070 6.960 ;
        RECT 21.420 6.910 21.750 6.930 ;
        RECT 24.770 4.850 25.060 6.930 ;
        RECT 110.050 6.650 110.330 6.970 ;
        RECT 109.870 6.340 110.330 6.650 ;
        RECT 110.050 6.220 110.330 6.340 ;
        RECT 41.190 4.850 41.510 4.870 ;
        RECT 97.190 4.850 98.350 4.880 ;
        RECT 24.580 3.730 98.350 4.850 ;
        RECT 41.190 3.710 41.510 3.730 ;
        RECT 52.560 3.650 54.480 3.730 ;
        RECT 62.370 3.620 64.300 3.730 ;
        RECT 97.190 3.700 98.350 3.730 ;
    END
    PORT
      LAYER met1 ;
        RECT 53.020 16.170 53.280 16.240 ;
        RECT 53.760 16.170 54.020 16.240 ;
        RECT 53.020 15.140 54.020 16.170 ;
        RECT 52.780 15.130 53.280 15.140 ;
        RECT 52.500 14.820 53.280 15.130 ;
        RECT 52.500 14.810 52.820 14.820 ;
        RECT 53.020 13.800 53.280 14.820 ;
        RECT 52.780 13.790 53.280 13.800 ;
        RECT 52.490 13.480 53.280 13.790 ;
        RECT 52.490 13.470 52.810 13.480 ;
        RECT 53.020 11.030 53.280 13.480 ;
        RECT 52.780 11.020 53.280 11.030 ;
        RECT 52.490 10.710 53.280 11.020 ;
        RECT 52.490 10.700 52.810 10.710 ;
        RECT 53.020 10.050 53.280 10.710 ;
        RECT 53.760 15.130 54.260 15.140 ;
        RECT 53.760 14.820 54.540 15.130 ;
        RECT 53.760 13.790 54.020 14.820 ;
        RECT 54.220 14.810 54.540 14.820 ;
        RECT 53.760 13.470 54.550 13.790 ;
        RECT 53.760 11.020 54.020 13.470 ;
        RECT 53.760 10.700 54.550 11.020 ;
        RECT 53.760 10.070 54.020 10.700 ;
        RECT 53.010 9.710 53.290 10.050 ;
        RECT 53.750 9.730 54.030 10.070 ;
        RECT 53.020 8.300 53.280 9.710 ;
        RECT 53.760 8.300 54.020 9.730 ;
        RECT 53.020 4.870 54.020 8.300 ;
        RECT 52.540 4.830 54.470 4.870 ;
        RECT 52.000 3.640 54.470 4.830 ;
        RECT 52.000 -7.850 52.940 3.640 ;
      LAYER via ;
        RECT 52.530 14.840 52.790 15.100 ;
        RECT 52.520 13.500 52.780 13.760 ;
        RECT 52.520 10.730 52.780 10.990 ;
        RECT 54.250 14.840 54.510 15.100 ;
        RECT 54.260 13.500 54.520 13.760 ;
        RECT 54.260 10.730 54.520 10.990 ;
        RECT 53.010 9.740 53.290 10.020 ;
        RECT 53.750 9.760 54.030 10.040 ;
        RECT 53.330 4.790 54.450 4.810 ;
        RECT 52.590 3.690 54.450 4.790 ;
        RECT 52.590 3.670 53.710 3.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 62.830 16.090 63.090 16.270 ;
        RECT 63.570 16.090 63.830 16.270 ;
        RECT 62.830 15.160 63.830 16.090 ;
        RECT 62.310 14.840 63.090 15.160 ;
        RECT 62.830 13.820 63.090 14.840 ;
        RECT 62.300 13.500 63.090 13.820 ;
        RECT 62.830 11.050 63.090 13.500 ;
        RECT 62.300 10.730 63.090 11.050 ;
        RECT 62.830 10.050 63.090 10.730 ;
        RECT 63.570 14.840 64.350 15.160 ;
        RECT 63.570 13.810 63.830 14.840 ;
        RECT 64.040 13.810 64.360 13.820 ;
        RECT 63.570 13.500 64.360 13.810 ;
        RECT 63.570 13.490 64.070 13.500 ;
        RECT 63.570 11.050 63.830 13.490 ;
        RECT 63.570 10.730 64.360 11.050 ;
        RECT 62.820 9.710 63.100 10.050 ;
        RECT 62.830 8.530 63.090 9.710 ;
        RECT 63.570 8.530 63.830 10.730 ;
        RECT 62.830 4.930 63.830 8.530 ;
        RECT 62.830 4.890 64.850 4.930 ;
        RECT 62.350 3.610 64.850 4.890 ;
        RECT 63.960 -6.390 64.850 3.610 ;
        RECT 63.960 -7.120 64.880 -6.390 ;
        RECT 63.930 -7.850 64.850 -7.120 ;
      LAYER via ;
        RECT 62.340 14.870 62.600 15.130 ;
        RECT 62.330 13.530 62.590 13.790 ;
        RECT 62.330 10.760 62.590 11.020 ;
        RECT 64.060 14.870 64.320 15.130 ;
        RECT 64.070 13.530 64.330 13.790 ;
        RECT 64.070 10.760 64.330 11.020 ;
        RECT 62.820 9.740 63.100 10.020 ;
        RECT 62.400 3.640 64.260 4.830 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 61.230 44.420 63.950 46.070 ;
        RECT 61.230 44.380 63.940 44.420 ;
        RECT 61.230 43.050 63.940 43.090 ;
        RECT 61.230 41.400 63.950 43.050 ;
        RECT 61.240 38.390 63.960 40.040 ;
        RECT 61.250 38.350 63.960 38.390 ;
        RECT 61.250 37.020 63.960 37.060 ;
        RECT 61.240 35.370 63.960 37.020 ;
        RECT 61.700 26.760 63.930 33.250 ;
        RECT 61.730 17.430 63.960 23.920 ;
      LAYER li1 ;
        RECT 6.050 61.390 6.220 61.550 ;
        RECT 7.450 61.390 7.620 61.550 ;
        RECT 6.050 61.250 6.290 61.390 ;
        RECT 6.050 61.220 7.090 61.250 ;
        RECT 7.450 61.240 7.660 61.390 ;
        RECT 9.290 61.280 9.960 61.450 ;
        RECT 7.450 61.220 8.500 61.240 ;
        RECT 6.090 61.070 7.090 61.220 ;
        RECT 7.490 61.070 8.500 61.220 ;
        RECT 9.290 60.490 9.960 60.660 ;
        RECT 7.300 60.390 7.620 60.430 ;
        RECT 6.420 60.220 8.500 60.390 ;
        RECT 23.310 60.350 26.620 61.330 ;
        RECT 30.710 60.530 30.940 61.220 ;
        RECT 35.410 60.480 35.640 61.170 ;
        RECT 7.290 60.200 7.620 60.220 ;
        RECT 7.300 60.170 7.620 60.200 ;
        RECT 6.600 59.810 8.420 59.980 ;
        RECT 7.300 59.570 7.620 59.590 ;
        RECT 6.420 59.400 8.500 59.570 ;
        RECT 9.210 59.560 9.420 59.990 ;
        RECT 23.420 59.690 23.590 60.040 ;
        RECT 24.140 59.770 24.310 59.800 ;
        RECT 24.050 59.730 24.370 59.770 ;
        RECT 24.820 59.760 24.990 59.800 ;
        RECT 22.690 59.650 23.590 59.690 ;
        RECT 9.230 59.540 9.400 59.560 ;
        RECT 22.680 59.460 23.590 59.650 ;
        RECT 24.040 59.540 24.370 59.730 ;
        RECT 24.740 59.720 25.060 59.760 ;
        RECT 24.050 59.510 24.370 59.540 ;
        RECT 24.730 59.530 25.060 59.720 ;
        RECT 24.140 59.470 24.310 59.510 ;
        RECT 24.740 59.500 25.060 59.530 ;
        RECT 24.820 59.470 24.990 59.500 ;
        RECT 22.690 59.430 23.590 59.460 ;
        RECT 31.920 59.450 32.090 59.470 ;
        RECT 7.290 59.360 7.620 59.400 ;
        RECT 7.300 59.330 7.620 59.360 ;
        RECT 9.290 59.060 9.960 59.230 ;
        RECT 6.420 58.560 7.090 58.730 ;
        RECT 7.820 58.560 8.500 58.730 ;
        RECT 8.800 58.440 8.990 58.500 ;
        RECT 8.800 58.270 9.970 58.440 ;
        RECT 8.730 57.990 8.900 58.020 ;
        RECT 8.730 57.960 9.060 57.990 ;
        RECT 8.730 57.770 9.070 57.960 ;
        RECT 8.730 57.730 9.060 57.770 ;
        RECT 8.730 57.690 8.900 57.730 ;
        RECT 7.480 57.610 7.650 57.670 ;
        RECT 9.300 57.660 9.970 57.830 ;
        RECT 6.420 57.440 7.090 57.610 ;
        RECT 7.480 57.440 8.500 57.610 ;
        RECT 7.480 57.340 7.650 57.440 ;
        RECT 7.280 56.770 7.600 56.790 ;
        RECT 8.710 56.770 9.030 56.810 ;
        RECT 6.410 56.600 9.990 56.770 ;
        RECT 7.270 56.560 7.600 56.600 ;
        RECT 8.700 56.580 9.030 56.600 ;
        RECT 7.280 56.530 7.600 56.560 ;
        RECT 8.710 56.550 9.030 56.580 ;
        RECT 6.490 56.170 6.810 56.210 ;
        RECT 7.420 56.170 7.740 56.210 ;
        RECT 8.120 56.170 8.440 56.210 ;
        RECT 8.860 56.170 9.180 56.210 ;
        RECT 6.480 56.100 6.810 56.170 ;
        RECT 7.410 56.100 7.740 56.170 ;
        RECT 8.110 56.100 8.440 56.170 ;
        RECT 8.850 56.150 9.180 56.170 ;
        RECT 9.570 56.160 9.890 56.200 ;
        RECT 9.560 56.150 9.890 56.160 ;
        RECT 8.850 56.100 9.890 56.150 ;
        RECT 6.460 55.930 9.890 56.100 ;
        RECT 11.560 55.990 11.730 56.660 ;
        RECT 22.050 56.570 22.220 59.220 ;
        RECT 23.420 59.030 23.590 59.430 ;
        RECT 29.030 59.280 32.090 59.450 ;
        RECT 31.920 58.630 32.090 59.280 ;
        RECT 23.310 57.550 26.620 58.530 ;
        RECT 31.920 58.460 33.190 58.630 ;
        RECT 30.710 57.540 30.940 58.230 ;
        RECT 22.050 56.030 22.230 56.570 ;
        RECT 21.970 55.990 22.290 56.030 ;
        RECT 23.310 56.000 26.620 56.980 ;
        RECT 30.710 56.530 30.940 57.220 ;
        RECT 31.920 56.050 32.090 58.460 ;
        RECT 34.660 56.810 34.830 57.700 ;
        RECT 31.830 56.010 32.150 56.050 ;
        RECT 9.040 55.920 9.890 55.930 ;
        RECT 21.960 55.800 22.290 55.990 ;
        RECT 31.820 55.820 32.150 56.010 ;
        RECT 21.970 55.770 22.290 55.800 ;
        RECT 31.830 55.790 32.150 55.820 ;
        RECT 22.000 52.210 23.520 52.220 ;
        RECT 22.000 51.420 23.550 52.210 ;
        RECT 43.090 50.160 43.440 50.260 ;
        RECT 46.850 50.250 47.140 50.270 ;
        RECT 46.680 50.210 47.140 50.250 ;
        RECT 45.700 50.190 47.140 50.210 ;
        RECT 44.750 50.160 45.210 50.190 ;
        RECT 41.680 49.990 42.440 50.160 ;
        RECT 42.690 49.990 43.860 50.160 ;
        RECT 44.100 50.020 45.210 50.160 ;
        RECT 45.660 50.030 47.140 50.190 ;
        RECT 45.660 50.020 46.850 50.030 ;
        RECT 44.100 49.990 44.920 50.020 ;
        RECT 41.680 49.980 41.910 49.990 ;
        RECT 41.640 49.540 41.910 49.980 ;
        RECT 44.660 49.850 44.920 49.990 ;
        RECT 43.120 49.540 43.450 49.800 ;
        RECT 44.660 49.680 45.840 49.850 ;
        RECT 44.660 49.540 44.920 49.680 ;
        RECT 41.090 49.400 41.260 49.460 ;
        RECT 41.060 49.180 41.280 49.400 ;
        RECT 41.610 49.360 41.940 49.540 ;
        RECT 42.190 49.370 44.350 49.540 ;
        RECT 44.590 49.370 44.920 49.540 ;
        RECT 44.750 49.320 44.920 49.370 ;
        RECT 45.210 49.180 45.420 49.510 ;
        RECT 45.660 49.240 45.840 49.680 ;
        RECT 47.470 49.580 47.640 50.340 ;
        RECT 47.840 50.190 48.290 50.340 ;
        RECT 47.840 50.020 48.440 50.190 ;
        RECT 48.900 50.010 49.230 50.180 ;
        RECT 47.260 49.570 47.640 49.580 ;
        RECT 47.260 49.510 47.730 49.570 ;
        RECT 48.980 49.550 49.160 50.010 ;
        RECT 46.390 49.400 47.730 49.510 ;
        RECT 46.390 49.340 47.650 49.400 ;
        RECT 48.200 49.380 49.160 49.550 ;
        RECT 47.260 49.290 47.650 49.340 ;
        RECT 41.090 49.130 41.260 49.180 ;
        RECT 43.090 48.410 43.440 48.510 ;
        RECT 46.850 48.500 47.140 48.520 ;
        RECT 46.680 48.460 47.140 48.500 ;
        RECT 45.700 48.440 47.140 48.460 ;
        RECT 44.750 48.410 45.210 48.440 ;
        RECT 41.680 48.240 42.440 48.410 ;
        RECT 42.690 48.240 43.860 48.410 ;
        RECT 44.100 48.270 45.210 48.410 ;
        RECT 45.660 48.280 47.140 48.440 ;
        RECT 45.660 48.270 46.850 48.280 ;
        RECT 44.100 48.240 44.920 48.270 ;
        RECT 41.680 48.230 41.910 48.240 ;
        RECT 41.640 47.790 41.910 48.230 ;
        RECT 44.660 48.100 44.920 48.240 ;
        RECT 43.120 47.790 43.450 48.050 ;
        RECT 44.660 47.930 45.840 48.100 ;
        RECT 44.660 47.790 44.920 47.930 ;
        RECT 41.090 47.650 41.260 47.710 ;
        RECT 41.060 47.430 41.280 47.650 ;
        RECT 41.610 47.610 41.940 47.790 ;
        RECT 42.190 47.620 44.350 47.790 ;
        RECT 44.590 47.620 44.920 47.790 ;
        RECT 44.750 47.570 44.920 47.620 ;
        RECT 45.210 47.430 45.420 47.760 ;
        RECT 45.660 47.490 45.840 47.930 ;
        RECT 47.470 47.830 47.640 48.590 ;
        RECT 47.840 48.440 48.290 48.590 ;
        RECT 47.840 48.270 48.440 48.440 ;
        RECT 48.900 48.260 49.230 48.430 ;
        RECT 69.970 48.260 70.640 49.130 ;
        RECT 82.250 48.280 84.350 49.130 ;
        RECT 47.260 47.820 47.640 47.830 ;
        RECT 47.260 47.760 47.730 47.820 ;
        RECT 48.980 47.800 49.160 48.260 ;
        RECT 46.390 47.650 47.730 47.760 ;
        RECT 46.390 47.590 47.650 47.650 ;
        RECT 48.200 47.630 49.160 47.800 ;
        RECT 47.260 47.540 47.650 47.590 ;
        RECT 41.090 47.380 41.260 47.430 ;
        RECT 20.200 46.890 20.400 46.930 ;
        RECT 19.890 46.630 20.400 46.890 ;
        RECT 20.200 46.600 20.400 46.630 ;
        RECT 20.790 46.900 20.990 46.930 ;
        RECT 20.790 46.860 21.300 46.900 ;
        RECT 20.790 46.670 21.310 46.860 ;
        RECT 20.790 46.640 21.300 46.670 ;
        RECT 43.090 46.660 43.440 46.760 ;
        RECT 46.850 46.750 47.140 46.770 ;
        RECT 46.680 46.710 47.140 46.750 ;
        RECT 45.700 46.690 47.140 46.710 ;
        RECT 44.750 46.660 45.210 46.690 ;
        RECT 20.790 46.600 20.990 46.640 ;
        RECT 41.680 46.490 42.440 46.660 ;
        RECT 42.690 46.490 43.860 46.660 ;
        RECT 44.100 46.520 45.210 46.660 ;
        RECT 45.660 46.530 47.140 46.690 ;
        RECT 45.660 46.520 46.850 46.530 ;
        RECT 44.100 46.490 44.920 46.520 ;
        RECT 41.680 46.480 41.910 46.490 ;
        RECT 19.620 46.390 19.980 46.460 ;
        RECT 19.460 46.290 19.980 46.390 ;
        RECT 21.490 46.350 21.660 46.400 ;
        RECT 21.480 46.320 21.660 46.350 ;
        RECT 21.480 46.310 21.910 46.320 ;
        RECT 19.460 46.210 19.830 46.290 ;
        RECT 19.460 46.160 19.790 46.210 ;
        RECT 19.460 46.130 19.780 46.160 ;
        RECT 21.480 46.080 22.070 46.310 ;
        RECT 21.480 46.070 21.910 46.080 ;
        RECT 21.480 46.040 21.670 46.070 ;
        RECT 41.640 46.040 41.910 46.480 ;
        RECT 44.660 46.350 44.920 46.490 ;
        RECT 43.120 46.040 43.450 46.300 ;
        RECT 44.660 46.180 45.840 46.350 ;
        RECT 44.660 46.040 44.920 46.180 ;
        RECT 21.490 46.010 21.670 46.040 ;
        RECT 20.210 45.900 20.410 45.940 ;
        RECT 19.900 45.640 20.410 45.900 ;
        RECT 20.210 45.610 20.410 45.640 ;
        RECT 20.800 45.910 21.000 45.940 ;
        RECT 20.800 45.870 21.310 45.910 ;
        RECT 41.090 45.900 41.260 45.960 ;
        RECT 20.800 45.680 21.320 45.870 ;
        RECT 41.060 45.680 41.280 45.900 ;
        RECT 41.610 45.860 41.940 46.040 ;
        RECT 42.190 45.870 44.350 46.040 ;
        RECT 44.590 45.870 44.920 46.040 ;
        RECT 44.750 45.820 44.920 45.870 ;
        RECT 45.210 45.680 45.420 46.010 ;
        RECT 45.660 45.740 45.840 46.180 ;
        RECT 47.470 46.080 47.640 46.840 ;
        RECT 47.840 46.690 48.290 46.840 ;
        RECT 80.140 46.760 80.310 46.810 ;
        RECT 47.840 46.520 48.440 46.690 ;
        RECT 48.900 46.510 49.230 46.680 ;
        RECT 47.260 46.070 47.640 46.080 ;
        RECT 47.260 46.010 47.730 46.070 ;
        RECT 48.980 46.050 49.160 46.510 ;
        RECT 80.140 46.500 80.700 46.760 ;
        RECT 81.610 46.510 81.810 46.550 ;
        RECT 80.140 46.480 80.310 46.500 ;
        RECT 56.590 46.130 56.790 46.480 ;
        RECT 58.070 46.230 58.600 46.400 ;
        RECT 58.840 46.380 59.030 46.410 ;
        RECT 58.840 46.210 59.900 46.380 ;
        RECT 76.750 46.230 77.280 46.400 ;
        RECT 58.840 46.180 59.030 46.210 ;
        RECT 46.390 45.900 47.730 46.010 ;
        RECT 46.390 45.840 47.650 45.900 ;
        RECT 48.200 45.880 49.160 46.050 ;
        RECT 56.580 46.100 56.790 46.130 ;
        RECT 47.260 45.790 47.650 45.840 ;
        RECT 20.800 45.650 21.310 45.680 ;
        RECT 20.800 45.610 21.000 45.650 ;
        RECT 41.090 45.630 41.260 45.680 ;
        RECT 56.580 45.520 56.800 46.100 ;
        RECT 56.580 45.510 56.790 45.520 ;
        RECT 19.440 45.300 19.990 45.470 ;
        RECT 56.960 45.340 57.150 45.350 ;
        RECT 19.440 45.240 19.770 45.300 ;
        RECT 19.440 45.210 19.760 45.240 ;
        RECT 20.210 44.910 20.410 44.950 ;
        RECT 19.900 44.650 20.410 44.910 ;
        RECT 20.210 44.620 20.410 44.650 ;
        RECT 20.800 44.920 21.000 44.950 ;
        RECT 20.800 44.880 21.310 44.920 ;
        RECT 43.090 44.910 43.440 45.010 ;
        RECT 46.850 45.000 47.140 45.020 ;
        RECT 46.680 44.960 47.140 45.000 ;
        RECT 45.700 44.940 47.140 44.960 ;
        RECT 44.750 44.910 45.210 44.940 ;
        RECT 20.800 44.690 21.320 44.880 ;
        RECT 41.680 44.740 42.440 44.910 ;
        RECT 42.690 44.740 43.860 44.910 ;
        RECT 44.100 44.770 45.210 44.910 ;
        RECT 45.660 44.780 47.140 44.940 ;
        RECT 45.660 44.770 46.850 44.780 ;
        RECT 44.100 44.740 44.920 44.770 ;
        RECT 41.680 44.730 41.910 44.740 ;
        RECT 20.800 44.660 21.310 44.690 ;
        RECT 20.800 44.620 21.000 44.660 ;
        RECT 19.420 44.310 19.990 44.480 ;
        RECT 19.420 44.250 19.750 44.310 ;
        RECT 41.640 44.290 41.910 44.730 ;
        RECT 44.660 44.600 44.920 44.740 ;
        RECT 43.120 44.290 43.450 44.550 ;
        RECT 44.660 44.430 45.840 44.600 ;
        RECT 44.660 44.290 44.920 44.430 ;
        RECT 19.420 44.220 19.740 44.250 ;
        RECT 41.090 44.150 41.260 44.210 ;
        RECT 19.710 43.940 20.030 43.980 ;
        RECT 19.710 43.920 20.040 43.940 ;
        RECT 41.060 43.930 41.280 44.150 ;
        RECT 41.610 44.110 41.940 44.290 ;
        RECT 42.190 44.120 44.350 44.290 ;
        RECT 44.590 44.120 44.920 44.290 ;
        RECT 44.750 44.070 44.920 44.120 ;
        RECT 45.210 43.930 45.420 44.260 ;
        RECT 45.660 43.990 45.840 44.430 ;
        RECT 47.470 44.330 47.640 45.090 ;
        RECT 47.840 44.940 48.290 45.090 ;
        RECT 56.950 45.050 57.150 45.340 ;
        RECT 47.840 44.770 48.440 44.940 ;
        RECT 48.900 44.760 49.230 44.930 ;
        RECT 47.260 44.320 47.640 44.330 ;
        RECT 47.260 44.260 47.730 44.320 ;
        RECT 48.980 44.300 49.160 44.760 ;
        RECT 56.890 44.720 57.160 45.050 ;
        RECT 46.390 44.150 47.730 44.260 ;
        RECT 46.390 44.090 47.650 44.150 ;
        RECT 48.200 44.130 49.160 44.300 ;
        RECT 57.350 44.240 57.520 45.850 ;
        RECT 58.180 44.750 58.350 45.840 ;
        RECT 59.310 45.820 59.500 45.850 ;
        RECT 58.770 45.650 59.500 45.820 ;
        RECT 59.730 45.820 59.900 46.210 ;
        RECT 78.560 46.130 78.760 46.480 ;
        RECT 78.560 46.100 78.770 46.130 ;
        RECT 59.730 45.650 60.470 45.820 ;
        RECT 59.310 45.620 59.500 45.650 ;
        RECT 61.530 45.030 61.760 45.550 ;
        RECT 58.770 44.860 61.760 45.030 ;
        RECT 57.950 44.710 58.350 44.750 ;
        RECT 57.940 44.520 58.350 44.710 ;
        RECT 66.730 44.670 67.280 45.100 ;
        RECT 68.070 44.670 68.620 45.100 ;
        RECT 71.700 44.860 71.930 45.550 ;
        RECT 77.000 45.320 77.170 45.840 ;
        RECT 76.840 45.060 77.170 45.320 ;
        RECT 57.950 44.490 58.350 44.520 ;
        RECT 47.260 44.040 47.650 44.090 ;
        RECT 57.340 44.050 57.520 44.240 ;
        RECT 58.180 44.150 58.350 44.490 ;
        RECT 58.840 44.240 59.030 44.420 ;
        RECT 58.770 44.070 59.120 44.240 ;
        RECT 19.710 43.720 20.330 43.920 ;
        RECT 20.160 43.590 20.330 43.720 ;
        RECT 20.840 43.880 21.010 43.920 ;
        RECT 41.090 43.880 41.260 43.930 ;
        RECT 20.840 43.840 21.330 43.880 ;
        RECT 20.840 43.650 21.340 43.840 ;
        RECT 59.690 43.660 59.900 44.090 ;
        RECT 60.120 44.070 60.460 44.240 ;
        RECT 20.840 43.620 21.330 43.650 ;
        RECT 59.710 43.640 59.880 43.660 ;
        RECT 20.840 43.590 21.010 43.620 ;
        RECT 19.520 43.480 19.950 43.500 ;
        RECT 19.500 43.310 19.950 43.480 ;
        RECT 41.090 43.360 41.260 43.410 ;
        RECT 19.520 43.290 19.950 43.310 ;
        RECT 41.060 43.140 41.280 43.360 ;
        RECT 41.090 43.080 41.260 43.140 ;
        RECT 41.610 43.000 41.940 43.180 ;
        RECT 44.750 43.170 44.920 43.220 ;
        RECT 42.190 43.000 44.350 43.170 ;
        RECT 44.590 43.000 44.920 43.170 ;
        RECT 45.210 43.030 45.420 43.360 ;
        RECT 19.710 42.950 20.030 42.990 ;
        RECT 19.710 42.930 20.040 42.950 ;
        RECT 19.710 42.730 20.330 42.930 ;
        RECT 20.160 42.600 20.330 42.730 ;
        RECT 20.840 42.890 21.010 42.930 ;
        RECT 20.840 42.850 21.330 42.890 ;
        RECT 20.840 42.660 21.340 42.850 ;
        RECT 20.840 42.630 21.330 42.660 ;
        RECT 20.840 42.600 21.010 42.630 ;
        RECT 41.640 42.560 41.910 43.000 ;
        RECT 43.120 42.740 43.450 43.000 ;
        RECT 44.660 42.860 44.920 43.000 ;
        RECT 45.660 42.860 45.840 43.300 ;
        RECT 47.260 43.200 47.650 43.250 ;
        RECT 46.390 43.140 47.650 43.200 ;
        RECT 46.390 43.030 47.730 43.140 ;
        RECT 47.260 42.970 47.730 43.030 ;
        RECT 48.200 42.990 49.160 43.160 ;
        RECT 47.260 42.960 47.640 42.970 ;
        RECT 41.680 42.550 41.910 42.560 ;
        RECT 44.660 42.690 45.840 42.860 ;
        RECT 44.660 42.550 44.920 42.690 ;
        RECT 19.520 42.490 19.950 42.510 ;
        RECT 19.500 42.320 19.950 42.490 ;
        RECT 41.680 42.380 42.440 42.550 ;
        RECT 42.690 42.380 43.860 42.550 ;
        RECT 44.100 42.520 44.920 42.550 ;
        RECT 44.100 42.380 45.210 42.520 ;
        RECT 21.450 42.360 21.680 42.370 ;
        RECT 19.520 42.300 19.950 42.320 ;
        RECT 21.370 42.190 21.700 42.360 ;
        RECT 43.090 42.280 43.440 42.380 ;
        RECT 44.750 42.350 45.210 42.380 ;
        RECT 45.660 42.510 46.850 42.520 ;
        RECT 45.660 42.350 47.140 42.510 ;
        RECT 45.700 42.330 47.140 42.350 ;
        RECT 46.680 42.290 47.140 42.330 ;
        RECT 46.850 42.270 47.140 42.290 ;
        RECT 47.470 42.200 47.640 42.960 ;
        RECT 48.980 42.530 49.160 42.990 ;
        RECT 50.150 42.980 50.320 43.400 ;
        RECT 50.960 43.280 51.200 43.310 ;
        RECT 50.630 43.110 51.200 43.280 ;
        RECT 51.440 43.110 52.780 43.280 ;
        RECT 53.230 43.110 54.190 43.280 ;
        RECT 50.960 43.070 51.200 43.110 ;
        RECT 53.740 43.100 53.910 43.110 ;
        RECT 50.080 42.760 50.250 42.800 ;
        RECT 50.020 42.590 50.250 42.760 ;
        RECT 47.840 42.350 48.440 42.520 ;
        RECT 48.900 42.360 49.230 42.530 ;
        RECT 47.840 42.200 48.290 42.350 ;
        RECT 50.080 42.240 50.250 42.590 ;
        RECT 50.420 42.660 50.610 42.680 ;
        RECT 53.370 42.660 53.710 42.840 ;
        RECT 50.420 42.490 50.980 42.660 ;
        RECT 51.440 42.490 54.190 42.660 ;
        RECT 50.420 42.450 50.610 42.490 ;
        RECT 54.720 42.420 54.890 43.350 ;
        RECT 55.120 42.510 55.290 43.400 ;
        RECT 57.340 43.330 57.520 43.520 ;
        RECT 56.890 42.520 57.160 42.850 ;
        RECT 56.950 42.230 57.150 42.520 ;
        RECT 56.960 42.220 57.150 42.230 ;
        RECT 21.450 42.180 21.680 42.190 ;
        RECT 56.580 42.050 56.790 42.060 ;
        RECT 19.710 41.960 20.030 42.000 ;
        RECT 19.710 41.940 20.040 41.960 ;
        RECT 19.710 41.740 20.330 41.940 ;
        RECT 20.160 41.610 20.330 41.740 ;
        RECT 20.840 41.900 21.010 41.940 ;
        RECT 20.840 41.860 21.330 41.900 ;
        RECT 20.840 41.670 21.340 41.860 ;
        RECT 20.840 41.640 21.330 41.670 ;
        RECT 20.840 41.610 21.010 41.640 ;
        RECT 41.090 41.610 41.260 41.660 ;
        RECT 19.520 41.500 19.950 41.520 ;
        RECT 19.500 41.330 19.950 41.500 ;
        RECT 41.060 41.390 41.280 41.610 ;
        RECT 41.090 41.330 41.260 41.390 ;
        RECT 19.520 41.310 19.950 41.330 ;
        RECT 41.610 41.250 41.940 41.430 ;
        RECT 44.750 41.420 44.920 41.470 ;
        RECT 42.190 41.250 44.350 41.420 ;
        RECT 44.590 41.250 44.920 41.420 ;
        RECT 45.210 41.280 45.420 41.610 ;
        RECT 41.640 40.810 41.910 41.250 ;
        RECT 43.120 40.990 43.450 41.250 ;
        RECT 44.660 41.110 44.920 41.250 ;
        RECT 45.660 41.110 45.840 41.550 ;
        RECT 47.260 41.450 47.650 41.500 ;
        RECT 50.080 41.480 50.250 41.830 ;
        RECT 46.390 41.390 47.650 41.450 ;
        RECT 46.390 41.280 47.730 41.390 ;
        RECT 47.260 41.220 47.730 41.280 ;
        RECT 48.200 41.240 49.160 41.410 ;
        RECT 50.020 41.310 50.250 41.480 ;
        RECT 50.420 41.580 50.610 41.620 ;
        RECT 50.420 41.410 50.980 41.580 ;
        RECT 51.440 41.410 54.190 41.580 ;
        RECT 50.420 41.390 50.610 41.410 ;
        RECT 50.080 41.270 50.250 41.310 ;
        RECT 47.260 41.210 47.640 41.220 ;
        RECT 41.680 40.800 41.910 40.810 ;
        RECT 44.660 40.940 45.840 41.110 ;
        RECT 44.660 40.800 44.920 40.940 ;
        RECT 41.680 40.630 42.440 40.800 ;
        RECT 42.690 40.630 43.860 40.800 ;
        RECT 44.100 40.770 44.920 40.800 ;
        RECT 44.100 40.630 45.210 40.770 ;
        RECT 43.090 40.530 43.440 40.630 ;
        RECT 44.750 40.600 45.210 40.630 ;
        RECT 45.660 40.760 46.850 40.770 ;
        RECT 45.660 40.600 47.140 40.760 ;
        RECT 45.700 40.580 47.140 40.600 ;
        RECT 46.680 40.540 47.140 40.580 ;
        RECT 46.850 40.520 47.140 40.540 ;
        RECT 47.470 40.450 47.640 41.210 ;
        RECT 48.980 40.780 49.160 41.240 ;
        RECT 53.370 41.230 53.710 41.410 ;
        RECT 47.840 40.600 48.440 40.770 ;
        RECT 48.900 40.610 49.230 40.780 ;
        RECT 50.150 40.670 50.320 41.090 ;
        RECT 50.960 40.960 51.200 41.000 ;
        RECT 53.740 40.960 53.910 40.970 ;
        RECT 50.630 40.790 51.200 40.960 ;
        RECT 51.440 40.790 52.780 40.960 ;
        RECT 53.230 40.790 54.190 40.960 ;
        RECT 50.960 40.760 51.200 40.790 ;
        RECT 54.720 40.720 54.890 41.650 ;
        RECT 55.120 40.670 55.290 41.560 ;
        RECT 56.580 41.470 56.800 42.050 ;
        RECT 57.350 41.720 57.520 43.330 ;
        RECT 58.180 43.060 58.350 43.420 ;
        RECT 58.770 43.330 59.120 43.500 ;
        RECT 59.310 43.480 59.500 43.530 ;
        RECT 60.210 43.500 60.380 44.070 ;
        RECT 64.490 43.840 64.680 44.240 ;
        RECT 70.670 43.840 70.860 44.240 ;
        RECT 77.000 44.150 77.170 45.060 ;
        RECT 77.830 44.240 78.000 45.850 ;
        RECT 78.550 45.520 78.770 46.100 ;
        RECT 78.560 45.510 78.770 45.520 ;
        RECT 79.560 45.400 79.740 46.330 ;
        RECT 81.380 46.250 81.810 46.510 ;
        RECT 80.290 46.070 80.620 46.240 ;
        RECT 81.610 46.220 81.810 46.250 ;
        RECT 80.370 45.930 80.620 46.070 ;
        RECT 80.370 45.670 80.850 45.930 ;
        RECT 81.200 45.860 81.370 45.900 ;
        RECT 81.610 45.860 81.810 45.890 ;
        RECT 79.440 45.370 79.760 45.400 ;
        RECT 78.200 45.340 78.390 45.350 ;
        RECT 78.200 45.050 78.400 45.340 ;
        RECT 79.440 45.180 79.770 45.370 ;
        RECT 79.440 45.140 79.760 45.180 ;
        RECT 78.190 44.720 78.480 45.050 ;
        RECT 77.830 44.050 78.010 44.240 ;
        RECT 64.490 43.830 64.870 43.840 ;
        RECT 61.130 43.650 64.870 43.830 ;
        RECT 64.490 43.610 64.870 43.650 ;
        RECT 70.480 43.830 70.860 43.840 ;
        RECT 70.480 43.650 74.220 43.830 ;
        RECT 70.480 43.610 70.860 43.650 ;
        RECT 59.310 43.470 59.540 43.480 ;
        RECT 60.120 43.470 60.460 43.500 ;
        RECT 59.310 43.330 60.460 43.470 ;
        RECT 58.850 43.120 59.040 43.330 ;
        RECT 59.310 43.300 60.290 43.330 ;
        RECT 59.450 43.270 60.290 43.300 ;
        RECT 64.490 43.230 64.680 43.610 ;
        RECT 57.940 43.020 58.350 43.060 ;
        RECT 57.930 42.830 58.350 43.020 ;
        RECT 66.730 42.940 67.280 43.370 ;
        RECT 68.070 42.940 68.620 43.370 ;
        RECT 70.670 43.230 70.860 43.610 ;
        RECT 57.940 42.800 58.350 42.830 ;
        RECT 58.180 41.730 58.350 42.800 ;
        RECT 58.770 42.610 61.700 42.710 ;
        RECT 58.770 42.540 61.760 42.610 ;
        RECT 60.790 42.220 60.960 42.280 ;
        RECT 60.770 42.010 60.980 42.220 ;
        RECT 59.300 41.920 59.490 41.950 ;
        RECT 60.790 41.940 60.960 42.010 ;
        RECT 61.530 41.920 61.760 42.540 ;
        RECT 71.700 41.920 71.930 42.650 ;
        RECT 77.000 42.560 77.170 43.420 ;
        RECT 76.840 42.300 77.170 42.560 ;
        RECT 58.770 41.750 59.490 41.920 ;
        RECT 59.300 41.720 59.490 41.750 ;
        RECT 59.660 41.750 60.470 41.920 ;
        RECT 56.580 41.440 56.790 41.470 ;
        RECT 56.590 41.090 56.790 41.440 ;
        RECT 58.870 41.410 59.060 41.440 ;
        RECT 59.660 41.410 59.850 41.750 ;
        RECT 77.000 41.730 77.170 42.300 ;
        RECT 77.830 43.330 78.010 43.520 ;
        RECT 77.830 41.720 78.000 43.330 ;
        RECT 78.190 42.520 78.480 42.850 ;
        RECT 78.200 42.230 78.400 42.520 ;
        RECT 78.200 42.220 78.390 42.230 ;
        RECT 78.560 42.050 78.770 42.060 ;
        RECT 78.550 41.470 78.770 42.050 ;
        RECT 58.070 41.170 58.600 41.340 ;
        RECT 58.870 41.230 59.850 41.410 ;
        RECT 78.560 41.440 78.770 41.470 ;
        RECT 58.870 41.210 59.060 41.230 ;
        RECT 76.750 41.170 77.280 41.340 ;
        RECT 78.560 41.090 78.760 41.440 ;
        RECT 79.560 41.230 79.740 45.140 ;
        RECT 80.370 44.290 80.540 45.670 ;
        RECT 81.200 45.600 81.810 45.860 ;
        RECT 81.200 45.570 81.370 45.600 ;
        RECT 81.610 45.560 81.810 45.600 ;
        RECT 82.200 45.560 82.750 46.550 ;
        RECT 83.570 46.400 84.200 46.570 ;
        RECT 83.570 46.300 83.960 46.400 ;
        RECT 83.570 46.270 83.950 46.300 ;
        RECT 83.570 46.120 83.930 46.270 ;
        RECT 83.220 45.950 83.930 46.120 ;
        RECT 83.220 45.200 83.920 45.510 ;
        RECT 81.200 45.010 81.370 45.040 ;
        RECT 81.610 45.010 81.810 45.050 ;
        RECT 81.200 44.750 81.810 45.010 ;
        RECT 81.200 44.710 81.370 44.750 ;
        RECT 81.610 44.720 81.810 44.750 ;
        RECT 81.610 44.360 81.810 44.390 ;
        RECT 80.170 44.090 80.490 44.120 ;
        RECT 81.380 44.100 81.810 44.360 ;
        RECT 80.170 43.900 80.500 44.090 ;
        RECT 81.610 44.060 81.810 44.100 ;
        RECT 82.200 44.060 82.750 45.050 ;
        RECT 83.070 44.970 83.920 45.200 ;
        RECT 83.220 44.630 83.920 44.970 ;
        RECT 83.680 44.270 84.000 44.310 ;
        RECT 83.680 44.210 84.010 44.270 ;
        RECT 83.210 44.080 84.010 44.210 ;
        RECT 83.210 44.050 84.000 44.080 ;
        RECT 83.210 44.030 83.910 44.050 ;
        RECT 109.090 44.020 109.410 44.050 ;
        RECT 110.660 44.020 110.980 44.050 ;
        RECT 80.170 43.860 80.490 43.900 ;
        RECT 80.170 43.780 80.340 43.860 ;
        RECT 80.120 43.610 80.340 43.780 ;
        RECT 107.870 43.680 108.040 43.960 ;
        RECT 109.090 43.830 109.420 44.020 ;
        RECT 110.100 43.880 110.290 43.900 ;
        RECT 109.090 43.790 109.410 43.830 ;
        RECT 107.870 43.640 108.080 43.680 ;
        RECT 107.870 43.620 108.100 43.640 ;
        RECT 109.220 43.630 109.390 43.790 ;
        RECT 109.830 43.710 110.290 43.880 ;
        RECT 110.660 43.830 110.990 44.020 ;
        RECT 111.230 43.880 111.420 43.910 ;
        RECT 110.660 43.790 110.980 43.830 ;
        RECT 110.080 43.700 110.290 43.710 ;
        RECT 110.100 43.670 110.290 43.700 ;
        RECT 110.720 43.630 110.890 43.790 ;
        RECT 111.230 43.710 111.670 43.880 ;
        RECT 111.230 43.680 111.420 43.710 ;
        RECT 80.120 43.450 80.290 43.610 ;
        RECT 107.870 43.600 108.130 43.620 ;
        RECT 83.670 43.550 83.990 43.590 ;
        RECT 107.870 43.550 108.210 43.600 ;
        RECT 81.610 43.510 81.810 43.550 ;
        RECT 80.650 43.190 80.840 43.310 ;
        RECT 81.380 43.250 81.810 43.510 ;
        RECT 81.610 43.220 81.810 43.250 ;
        RECT 80.290 43.080 80.840 43.190 ;
        RECT 80.290 43.020 80.830 43.080 ;
        RECT 80.370 41.240 80.540 43.020 ;
        RECT 81.200 42.860 81.370 42.900 ;
        RECT 81.610 42.860 81.810 42.890 ;
        RECT 81.200 42.600 81.810 42.860 ;
        RECT 81.200 42.570 81.370 42.600 ;
        RECT 81.610 42.560 81.810 42.600 ;
        RECT 82.200 42.560 82.750 43.550 ;
        RECT 83.210 43.370 84.000 43.550 ;
        RECT 107.870 43.490 108.360 43.550 ;
        RECT 107.870 43.460 108.380 43.490 ;
        RECT 107.910 43.430 108.380 43.460 ;
        RECT 108.040 43.380 108.380 43.430 ;
        RECT 108.160 43.370 108.380 43.380 ;
        RECT 83.670 43.360 84.000 43.370 ;
        RECT 83.670 43.330 83.990 43.360 ;
        RECT 108.170 43.340 108.380 43.370 ;
        RECT 108.190 43.260 108.380 43.340 ;
        RECT 109.550 43.260 109.880 43.380 ;
        RECT 111.950 43.290 112.120 43.970 ;
        RECT 107.700 43.210 107.870 43.230 ;
        RECT 83.220 42.610 83.920 42.950 ;
        RECT 107.680 42.780 107.890 43.210 ;
        RECT 108.190 43.090 108.710 43.260 ;
        RECT 108.190 43.060 108.380 43.090 ;
        RECT 109.060 43.080 110.960 43.260 ;
        RECT 111.690 43.250 112.120 43.290 ;
        RECT 111.340 43.090 112.120 43.250 ;
        RECT 111.340 43.080 111.880 43.090 ;
        RECT 111.690 43.060 111.880 43.080 ;
        RECT 83.070 42.380 83.920 42.610 ;
        RECT 83.220 42.070 83.920 42.380 ;
        RECT 107.680 42.060 107.890 42.490 ;
        RECT 108.190 42.180 108.380 42.210 ;
        RECT 111.690 42.190 111.880 42.210 ;
        RECT 81.200 42.010 81.370 42.040 ;
        RECT 81.610 42.010 81.810 42.050 ;
        RECT 81.200 41.750 81.810 42.010 ;
        RECT 81.200 41.710 81.370 41.750 ;
        RECT 81.610 41.720 81.810 41.750 ;
        RECT 81.610 41.360 81.810 41.390 ;
        RECT 81.380 41.100 81.810 41.360 ;
        RECT 81.610 41.060 81.810 41.100 ;
        RECT 82.200 41.060 82.750 42.050 ;
        RECT 107.700 42.040 107.870 42.060 ;
        RECT 108.190 42.010 108.710 42.180 ;
        RECT 109.060 42.010 110.960 42.190 ;
        RECT 111.340 42.180 111.880 42.190 ;
        RECT 111.340 42.020 112.120 42.180 ;
        RECT 108.190 41.930 108.380 42.010 ;
        RECT 108.170 41.900 108.380 41.930 ;
        RECT 108.160 41.890 108.380 41.900 ;
        RECT 109.550 41.890 109.880 42.010 ;
        RECT 111.690 41.980 112.120 42.020 ;
        RECT 108.040 41.840 108.380 41.890 ;
        RECT 107.910 41.810 108.380 41.840 ;
        RECT 107.870 41.780 108.380 41.810 ;
        RECT 107.870 41.720 108.360 41.780 ;
        RECT 107.870 41.670 108.210 41.720 ;
        RECT 107.870 41.650 108.130 41.670 ;
        RECT 107.870 41.630 108.100 41.650 ;
        RECT 83.220 41.460 83.930 41.630 ;
        RECT 83.570 41.180 83.930 41.460 ;
        RECT 107.870 41.590 108.080 41.630 ;
        RECT 107.870 41.310 108.040 41.590 ;
        RECT 109.220 41.480 109.390 41.640 ;
        RECT 110.100 41.570 110.290 41.600 ;
        RECT 110.080 41.560 110.290 41.570 ;
        RECT 109.090 41.440 109.410 41.480 ;
        RECT 109.090 41.250 109.420 41.440 ;
        RECT 109.830 41.390 110.290 41.560 ;
        RECT 110.720 41.480 110.890 41.640 ;
        RECT 111.230 41.560 111.420 41.590 ;
        RECT 110.100 41.370 110.290 41.390 ;
        RECT 110.660 41.440 110.980 41.480 ;
        RECT 110.660 41.250 110.990 41.440 ;
        RECT 111.230 41.390 111.670 41.560 ;
        RECT 111.230 41.360 111.420 41.390 ;
        RECT 111.950 41.300 112.120 41.980 ;
        RECT 109.090 41.220 109.410 41.250 ;
        RECT 110.660 41.220 110.980 41.250 ;
        RECT 83.570 41.010 84.200 41.180 ;
        RECT 109.090 40.820 109.410 40.850 ;
        RECT 110.660 40.820 110.980 40.850 ;
        RECT 80.140 40.730 80.310 40.780 ;
        RECT 47.840 40.450 48.290 40.600 ;
        RECT 41.090 39.860 41.260 39.910 ;
        RECT 41.060 39.640 41.280 39.860 ;
        RECT 41.090 39.580 41.260 39.640 ;
        RECT 41.610 39.500 41.940 39.680 ;
        RECT 44.750 39.670 44.920 39.720 ;
        RECT 42.190 39.500 44.350 39.670 ;
        RECT 44.590 39.500 44.920 39.670 ;
        RECT 45.210 39.530 45.420 39.860 ;
        RECT 41.640 39.060 41.910 39.500 ;
        RECT 43.120 39.240 43.450 39.500 ;
        RECT 44.660 39.360 44.920 39.500 ;
        RECT 45.660 39.360 45.840 39.800 ;
        RECT 50.150 39.780 50.320 40.200 ;
        RECT 50.960 40.080 51.200 40.110 ;
        RECT 50.630 39.910 51.200 40.080 ;
        RECT 51.440 39.910 52.780 40.080 ;
        RECT 53.230 39.910 54.190 40.080 ;
        RECT 50.960 39.870 51.200 39.910 ;
        RECT 53.740 39.900 53.910 39.910 ;
        RECT 47.260 39.700 47.650 39.750 ;
        RECT 46.390 39.640 47.650 39.700 ;
        RECT 46.390 39.530 47.730 39.640 ;
        RECT 47.260 39.470 47.730 39.530 ;
        RECT 48.200 39.490 49.160 39.660 ;
        RECT 50.080 39.560 50.250 39.600 ;
        RECT 47.260 39.460 47.640 39.470 ;
        RECT 41.680 39.050 41.910 39.060 ;
        RECT 44.660 39.190 45.840 39.360 ;
        RECT 44.660 39.050 44.920 39.190 ;
        RECT 41.680 38.880 42.440 39.050 ;
        RECT 42.690 38.880 43.860 39.050 ;
        RECT 44.100 39.020 44.920 39.050 ;
        RECT 44.100 38.880 45.210 39.020 ;
        RECT 43.090 38.780 43.440 38.880 ;
        RECT 44.750 38.850 45.210 38.880 ;
        RECT 45.660 39.010 46.850 39.020 ;
        RECT 45.660 38.850 47.140 39.010 ;
        RECT 45.700 38.830 47.140 38.850 ;
        RECT 46.680 38.790 47.140 38.830 ;
        RECT 46.850 38.770 47.140 38.790 ;
        RECT 47.470 38.700 47.640 39.460 ;
        RECT 48.980 39.030 49.160 39.490 ;
        RECT 50.020 39.390 50.250 39.560 ;
        RECT 50.080 39.040 50.250 39.390 ;
        RECT 50.420 39.460 50.610 39.480 ;
        RECT 53.370 39.460 53.710 39.640 ;
        RECT 50.420 39.290 50.980 39.460 ;
        RECT 51.440 39.290 54.190 39.460 ;
        RECT 50.420 39.250 50.610 39.290 ;
        RECT 54.720 39.220 54.890 40.150 ;
        RECT 55.120 39.310 55.290 40.200 ;
        RECT 56.600 40.100 56.800 40.450 ;
        RECT 58.080 40.200 58.610 40.370 ;
        RECT 56.590 40.070 56.800 40.100 ;
        RECT 56.590 39.490 56.810 40.070 ;
        RECT 56.590 39.480 56.800 39.490 ;
        RECT 56.970 39.310 57.160 39.320 ;
        RECT 47.840 38.850 48.440 39.020 ;
        RECT 48.900 38.860 49.230 39.030 ;
        RECT 56.960 39.020 57.160 39.310 ;
        RECT 47.840 38.700 48.290 38.850 ;
        RECT 56.880 38.690 57.170 39.020 ;
        RECT 50.080 38.280 50.250 38.630 ;
        RECT 41.090 38.110 41.260 38.160 ;
        RECT 50.020 38.110 50.250 38.280 ;
        RECT 50.420 38.380 50.610 38.420 ;
        RECT 50.420 38.210 50.980 38.380 ;
        RECT 51.440 38.210 54.190 38.380 ;
        RECT 50.420 38.190 50.610 38.210 ;
        RECT 41.060 37.890 41.280 38.110 ;
        RECT 41.090 37.830 41.260 37.890 ;
        RECT 41.610 37.750 41.940 37.930 ;
        RECT 44.750 37.920 44.920 37.970 ;
        RECT 42.190 37.750 44.350 37.920 ;
        RECT 44.590 37.750 44.920 37.920 ;
        RECT 45.210 37.780 45.420 38.110 ;
        RECT 50.080 38.070 50.250 38.110 ;
        RECT 41.640 37.310 41.910 37.750 ;
        RECT 43.120 37.490 43.450 37.750 ;
        RECT 44.660 37.610 44.920 37.750 ;
        RECT 45.660 37.610 45.840 38.050 ;
        RECT 53.370 38.030 53.710 38.210 ;
        RECT 47.260 37.950 47.650 38.000 ;
        RECT 46.390 37.890 47.650 37.950 ;
        RECT 46.390 37.780 47.730 37.890 ;
        RECT 47.260 37.720 47.730 37.780 ;
        RECT 48.200 37.740 49.160 37.910 ;
        RECT 47.260 37.710 47.640 37.720 ;
        RECT 41.680 37.300 41.910 37.310 ;
        RECT 44.660 37.440 45.840 37.610 ;
        RECT 44.660 37.300 44.920 37.440 ;
        RECT 41.680 37.130 42.440 37.300 ;
        RECT 42.690 37.130 43.860 37.300 ;
        RECT 44.100 37.270 44.920 37.300 ;
        RECT 44.100 37.130 45.210 37.270 ;
        RECT 43.090 37.030 43.440 37.130 ;
        RECT 44.750 37.100 45.210 37.130 ;
        RECT 45.660 37.260 46.850 37.270 ;
        RECT 45.660 37.100 47.140 37.260 ;
        RECT 45.700 37.080 47.140 37.100 ;
        RECT 46.680 37.040 47.140 37.080 ;
        RECT 46.850 37.020 47.140 37.040 ;
        RECT 47.470 36.950 47.640 37.710 ;
        RECT 48.980 37.280 49.160 37.740 ;
        RECT 50.150 37.470 50.320 37.890 ;
        RECT 50.960 37.760 51.200 37.800 ;
        RECT 53.740 37.760 53.910 37.770 ;
        RECT 50.630 37.590 51.200 37.760 ;
        RECT 51.440 37.590 52.780 37.760 ;
        RECT 53.230 37.590 54.190 37.760 ;
        RECT 50.960 37.560 51.200 37.590 ;
        RECT 54.720 37.520 54.890 38.450 ;
        RECT 55.120 37.470 55.290 38.360 ;
        RECT 57.360 38.210 57.530 39.820 ;
        RECT 57.350 38.020 57.530 38.210 ;
        RECT 58.190 39.290 58.360 39.810 ;
        RECT 60.800 39.770 65.860 40.600 ;
        RECT 80.140 40.470 80.700 40.730 ;
        RECT 81.610 40.480 81.810 40.520 ;
        RECT 80.140 40.450 80.310 40.470 ;
        RECT 76.750 40.200 77.280 40.370 ;
        RECT 78.560 40.100 78.760 40.450 ;
        RECT 78.560 40.070 78.770 40.100 ;
        RECT 65.310 39.690 65.790 39.770 ;
        RECT 58.190 39.030 58.520 39.290 ;
        RECT 58.190 38.120 58.360 39.030 ;
        RECT 63.430 38.830 63.660 39.520 ;
        RECT 65.310 39.440 65.780 39.690 ;
        RECT 66.740 38.640 67.290 39.070 ;
        RECT 68.070 38.640 68.620 39.070 ;
        RECT 71.700 38.830 71.930 39.520 ;
        RECT 77.000 39.290 77.170 39.810 ;
        RECT 76.840 39.030 77.170 39.290 ;
        RECT 64.500 37.800 64.890 38.210 ;
        RECT 61.140 37.620 64.890 37.800 ;
        RECT 57.350 37.300 57.530 37.490 ;
        RECT 47.840 37.100 48.440 37.270 ;
        RECT 48.900 37.110 49.230 37.280 ;
        RECT 47.840 36.950 48.290 37.100 ;
        RECT 56.880 36.490 57.170 36.820 ;
        RECT 56.960 36.200 57.160 36.490 ;
        RECT 56.970 36.190 57.160 36.200 ;
        RECT 56.590 36.020 56.800 36.030 ;
        RECT 56.590 35.440 56.810 36.020 ;
        RECT 57.360 35.690 57.530 37.300 ;
        RECT 58.190 36.530 58.360 37.390 ;
        RECT 64.500 37.200 64.890 37.620 ;
        RECT 70.440 37.800 70.860 38.210 ;
        RECT 77.000 38.120 77.170 39.030 ;
        RECT 77.830 38.210 78.000 39.820 ;
        RECT 78.550 39.490 78.770 40.070 ;
        RECT 78.560 39.480 78.770 39.490 ;
        RECT 79.560 39.370 79.740 40.300 ;
        RECT 81.380 40.220 81.810 40.480 ;
        RECT 80.290 40.040 80.620 40.210 ;
        RECT 81.610 40.190 81.810 40.220 ;
        RECT 80.370 39.900 80.620 40.040 ;
        RECT 80.370 39.640 80.850 39.900 ;
        RECT 81.200 39.830 81.370 39.870 ;
        RECT 81.610 39.830 81.810 39.860 ;
        RECT 79.440 39.340 79.760 39.370 ;
        RECT 78.200 39.310 78.390 39.320 ;
        RECT 78.200 39.020 78.400 39.310 ;
        RECT 79.440 39.150 79.770 39.340 ;
        RECT 79.440 39.110 79.760 39.150 ;
        RECT 78.190 38.690 78.480 39.020 ;
        RECT 77.830 38.020 78.010 38.210 ;
        RECT 70.440 37.620 74.220 37.800 ;
        RECT 66.740 36.910 67.290 37.340 ;
        RECT 68.070 36.910 68.620 37.340 ;
        RECT 70.440 37.200 70.860 37.620 ;
        RECT 58.190 36.270 58.520 36.530 ;
        RECT 58.190 35.700 58.360 36.270 ;
        RECT 63.430 35.890 63.660 36.620 ;
        RECT 65.470 35.760 65.810 36.010 ;
        RECT 71.700 35.890 71.930 36.620 ;
        RECT 77.000 36.530 77.170 37.390 ;
        RECT 76.840 36.270 77.170 36.530 ;
        RECT 65.470 35.680 65.820 35.760 ;
        RECT 77.000 35.700 77.170 36.270 ;
        RECT 77.830 37.300 78.010 37.490 ;
        RECT 77.830 35.690 78.000 37.300 ;
        RECT 78.190 36.490 78.480 36.820 ;
        RECT 78.200 36.200 78.400 36.490 ;
        RECT 78.200 36.190 78.390 36.200 ;
        RECT 78.560 36.020 78.770 36.030 ;
        RECT 56.590 35.410 56.800 35.440 ;
        RECT 56.600 35.060 56.800 35.410 ;
        RECT 58.080 35.140 58.610 35.310 ;
        RECT 60.770 34.830 65.820 35.680 ;
        RECT 78.550 35.440 78.770 36.020 ;
        RECT 78.560 35.410 78.770 35.440 ;
        RECT 76.750 35.140 77.280 35.310 ;
        RECT 78.560 35.060 78.760 35.410 ;
        RECT 79.560 35.200 79.740 39.110 ;
        RECT 80.370 38.260 80.540 39.640 ;
        RECT 81.200 39.570 81.810 39.830 ;
        RECT 81.200 39.540 81.370 39.570 ;
        RECT 81.610 39.530 81.810 39.570 ;
        RECT 82.200 39.530 82.750 40.520 ;
        RECT 83.570 40.370 84.200 40.540 ;
        RECT 107.870 40.480 108.040 40.760 ;
        RECT 109.090 40.630 109.420 40.820 ;
        RECT 110.100 40.680 110.290 40.700 ;
        RECT 109.090 40.590 109.410 40.630 ;
        RECT 107.870 40.440 108.080 40.480 ;
        RECT 107.870 40.420 108.100 40.440 ;
        RECT 109.220 40.430 109.390 40.590 ;
        RECT 109.830 40.510 110.290 40.680 ;
        RECT 110.660 40.630 110.990 40.820 ;
        RECT 111.230 40.680 111.420 40.710 ;
        RECT 110.660 40.590 110.980 40.630 ;
        RECT 110.080 40.500 110.290 40.510 ;
        RECT 110.100 40.470 110.290 40.500 ;
        RECT 110.720 40.430 110.890 40.590 ;
        RECT 111.230 40.510 111.670 40.680 ;
        RECT 111.230 40.480 111.420 40.510 ;
        RECT 107.870 40.400 108.130 40.420 ;
        RECT 83.570 40.270 83.960 40.370 ;
        RECT 107.870 40.350 108.210 40.400 ;
        RECT 107.870 40.290 108.360 40.350 ;
        RECT 83.570 40.240 83.950 40.270 ;
        RECT 107.870 40.260 108.380 40.290 ;
        RECT 83.570 40.090 83.930 40.240 ;
        RECT 107.910 40.230 108.380 40.260 ;
        RECT 108.040 40.180 108.380 40.230 ;
        RECT 108.160 40.170 108.380 40.180 ;
        RECT 108.170 40.140 108.380 40.170 ;
        RECT 83.220 39.920 83.930 40.090 ;
        RECT 108.190 40.060 108.380 40.140 ;
        RECT 109.550 40.060 109.880 40.180 ;
        RECT 111.950 40.090 112.120 40.770 ;
        RECT 107.700 40.010 107.870 40.030 ;
        RECT 107.680 39.580 107.890 40.010 ;
        RECT 108.190 39.890 108.710 40.060 ;
        RECT 108.190 39.860 108.380 39.890 ;
        RECT 109.060 39.880 110.960 40.060 ;
        RECT 111.690 40.050 112.120 40.090 ;
        RECT 111.340 39.890 112.120 40.050 ;
        RECT 111.340 39.880 111.880 39.890 ;
        RECT 111.690 39.860 111.880 39.880 ;
        RECT 83.220 39.170 83.920 39.480 ;
        RECT 81.200 38.980 81.370 39.010 ;
        RECT 81.610 38.980 81.810 39.020 ;
        RECT 81.200 38.720 81.810 38.980 ;
        RECT 81.200 38.680 81.370 38.720 ;
        RECT 81.610 38.690 81.810 38.720 ;
        RECT 81.610 38.330 81.810 38.360 ;
        RECT 80.170 38.060 80.490 38.090 ;
        RECT 81.380 38.070 81.810 38.330 ;
        RECT 80.170 37.870 80.500 38.060 ;
        RECT 81.610 38.030 81.810 38.070 ;
        RECT 82.200 38.030 82.750 39.020 ;
        RECT 83.070 38.940 83.920 39.170 ;
        RECT 83.220 38.600 83.920 38.940 ;
        RECT 107.680 38.860 107.890 39.290 ;
        RECT 108.190 38.980 108.380 39.010 ;
        RECT 111.690 38.990 111.880 39.010 ;
        RECT 107.700 38.840 107.870 38.860 ;
        RECT 108.190 38.810 108.710 38.980 ;
        RECT 109.060 38.810 110.960 38.990 ;
        RECT 111.340 38.980 111.880 38.990 ;
        RECT 111.340 38.820 112.120 38.980 ;
        RECT 108.190 38.730 108.380 38.810 ;
        RECT 108.170 38.700 108.380 38.730 ;
        RECT 108.160 38.690 108.380 38.700 ;
        RECT 109.550 38.690 109.880 38.810 ;
        RECT 111.690 38.780 112.120 38.820 ;
        RECT 108.040 38.640 108.380 38.690 ;
        RECT 107.910 38.610 108.380 38.640 ;
        RECT 107.870 38.580 108.380 38.610 ;
        RECT 107.870 38.520 108.360 38.580 ;
        RECT 107.870 38.470 108.210 38.520 ;
        RECT 107.870 38.450 108.130 38.470 ;
        RECT 107.870 38.430 108.100 38.450 ;
        RECT 107.870 38.390 108.080 38.430 ;
        RECT 83.680 38.240 84.000 38.280 ;
        RECT 83.680 38.180 84.010 38.240 ;
        RECT 83.210 38.050 84.010 38.180 ;
        RECT 107.870 38.110 108.040 38.390 ;
        RECT 109.220 38.280 109.390 38.440 ;
        RECT 110.100 38.370 110.290 38.400 ;
        RECT 110.080 38.360 110.290 38.370 ;
        RECT 109.090 38.240 109.410 38.280 ;
        RECT 109.090 38.050 109.420 38.240 ;
        RECT 109.830 38.190 110.290 38.360 ;
        RECT 110.720 38.280 110.890 38.440 ;
        RECT 111.230 38.360 111.420 38.390 ;
        RECT 110.100 38.170 110.290 38.190 ;
        RECT 110.660 38.240 110.980 38.280 ;
        RECT 110.660 38.050 110.990 38.240 ;
        RECT 111.230 38.190 111.670 38.360 ;
        RECT 111.230 38.160 111.420 38.190 ;
        RECT 111.950 38.100 112.120 38.780 ;
        RECT 83.210 38.020 84.000 38.050 ;
        RECT 109.090 38.020 109.410 38.050 ;
        RECT 110.660 38.020 110.980 38.050 ;
        RECT 83.210 38.000 83.910 38.020 ;
        RECT 80.170 37.830 80.490 37.870 ;
        RECT 80.170 37.750 80.340 37.830 ;
        RECT 80.120 37.580 80.340 37.750 ;
        RECT 80.120 37.420 80.290 37.580 ;
        RECT 83.670 37.520 83.990 37.560 ;
        RECT 81.610 37.480 81.810 37.520 ;
        RECT 80.650 37.160 80.840 37.280 ;
        RECT 81.380 37.220 81.810 37.480 ;
        RECT 81.610 37.190 81.810 37.220 ;
        RECT 80.290 37.050 80.840 37.160 ;
        RECT 80.290 36.990 80.830 37.050 ;
        RECT 80.370 35.210 80.540 36.990 ;
        RECT 81.200 36.830 81.370 36.870 ;
        RECT 81.610 36.830 81.810 36.860 ;
        RECT 81.200 36.570 81.810 36.830 ;
        RECT 81.200 36.540 81.370 36.570 ;
        RECT 81.610 36.530 81.810 36.570 ;
        RECT 82.200 36.530 82.750 37.520 ;
        RECT 83.210 37.340 84.000 37.520 ;
        RECT 83.670 37.330 84.000 37.340 ;
        RECT 83.670 37.300 83.990 37.330 ;
        RECT 83.220 36.580 83.920 36.920 ;
        RECT 83.070 36.350 83.920 36.580 ;
        RECT 83.220 36.040 83.920 36.350 ;
        RECT 81.200 35.980 81.370 36.010 ;
        RECT 81.610 35.980 81.810 36.020 ;
        RECT 81.200 35.720 81.810 35.980 ;
        RECT 81.200 35.680 81.370 35.720 ;
        RECT 81.610 35.690 81.810 35.720 ;
        RECT 81.610 35.330 81.810 35.360 ;
        RECT 81.380 35.070 81.810 35.330 ;
        RECT 81.610 35.030 81.810 35.070 ;
        RECT 82.200 35.030 82.750 36.020 ;
        RECT 83.220 35.430 83.930 35.600 ;
        RECT 83.570 35.150 83.930 35.430 ;
        RECT 83.570 34.980 84.200 35.150 ;
        RECT 41.090 33.230 41.260 33.280 ;
        RECT 41.060 33.010 41.280 33.230 ;
        RECT 41.090 32.950 41.260 33.010 ;
        RECT 41.610 32.870 41.940 33.050 ;
        RECT 44.750 33.040 44.920 33.090 ;
        RECT 42.190 32.870 44.350 33.040 ;
        RECT 44.590 32.870 44.920 33.040 ;
        RECT 45.210 32.900 45.420 33.230 ;
        RECT 41.640 32.430 41.910 32.870 ;
        RECT 43.120 32.610 43.450 32.870 ;
        RECT 44.660 32.730 44.920 32.870 ;
        RECT 45.660 32.730 45.840 33.170 ;
        RECT 47.260 33.070 47.650 33.120 ;
        RECT 46.390 33.010 47.650 33.070 ;
        RECT 46.390 32.900 47.730 33.010 ;
        RECT 47.260 32.840 47.730 32.900 ;
        RECT 48.200 32.860 49.160 33.030 ;
        RECT 47.260 32.830 47.640 32.840 ;
        RECT 41.680 32.420 41.910 32.430 ;
        RECT 44.660 32.560 45.840 32.730 ;
        RECT 44.660 32.420 44.920 32.560 ;
        RECT 41.680 32.250 42.440 32.420 ;
        RECT 42.690 32.250 43.860 32.420 ;
        RECT 44.100 32.390 44.920 32.420 ;
        RECT 44.100 32.250 45.210 32.390 ;
        RECT 43.090 32.150 43.440 32.250 ;
        RECT 44.750 32.220 45.210 32.250 ;
        RECT 45.660 32.380 46.850 32.390 ;
        RECT 45.660 32.220 47.140 32.380 ;
        RECT 45.700 32.200 47.140 32.220 ;
        RECT 46.680 32.160 47.140 32.200 ;
        RECT 46.850 32.140 47.140 32.160 ;
        RECT 47.470 32.070 47.640 32.830 ;
        RECT 48.980 32.400 49.160 32.860 ;
        RECT 50.130 32.510 50.300 32.930 ;
        RECT 50.940 32.810 51.180 32.840 ;
        RECT 50.610 32.640 51.180 32.810 ;
        RECT 51.420 32.640 52.760 32.810 ;
        RECT 53.210 32.640 54.170 32.810 ;
        RECT 50.940 32.600 51.180 32.640 ;
        RECT 53.720 32.630 53.890 32.640 ;
        RECT 47.840 32.220 48.440 32.390 ;
        RECT 48.900 32.230 49.230 32.400 ;
        RECT 50.060 32.290 50.230 32.330 ;
        RECT 47.840 32.070 48.290 32.220 ;
        RECT 50.000 32.120 50.230 32.290 ;
        RECT 50.060 31.770 50.230 32.120 ;
        RECT 50.400 32.190 50.590 32.210 ;
        RECT 53.350 32.190 53.690 32.370 ;
        RECT 50.400 32.020 50.960 32.190 ;
        RECT 51.420 32.020 54.170 32.190 ;
        RECT 50.400 31.980 50.590 32.020 ;
        RECT 54.700 31.950 54.870 32.880 ;
        RECT 55.100 32.040 55.270 32.930 ;
        RECT 58.010 32.520 58.210 32.870 ;
        RECT 59.750 32.790 60.070 32.800 ;
        RECT 59.490 32.620 60.070 32.790 ;
        RECT 59.740 32.570 60.070 32.620 ;
        RECT 59.750 32.540 60.070 32.570 ;
        RECT 75.270 32.790 75.590 32.800 ;
        RECT 75.270 32.620 75.850 32.790 ;
        RECT 75.270 32.570 75.600 32.620 ;
        RECT 75.270 32.540 75.590 32.570 ;
        RECT 58.000 32.490 58.210 32.520 ;
        RECT 77.130 32.520 77.330 32.870 ;
        RECT 58.000 31.900 58.220 32.490 ;
        RECT 58.740 31.900 58.940 32.500 ;
        RECT 59.750 32.210 60.070 32.250 ;
        RECT 59.740 32.170 60.070 32.210 ;
        RECT 59.490 32.000 60.070 32.170 ;
        RECT 59.750 31.990 60.070 32.000 ;
        RECT 75.270 32.210 75.590 32.250 ;
        RECT 75.270 32.170 75.600 32.210 ;
        RECT 75.270 32.000 75.850 32.170 ;
        RECT 75.270 31.990 75.590 32.000 ;
        RECT 76.400 31.900 76.600 32.500 ;
        RECT 77.130 32.490 77.340 32.520 ;
        RECT 77.120 31.900 77.340 32.490 ;
        RECT 41.090 31.480 41.260 31.530 ;
        RECT 41.060 31.260 41.280 31.480 ;
        RECT 41.090 31.200 41.260 31.260 ;
        RECT 41.610 31.120 41.940 31.300 ;
        RECT 44.750 31.290 44.920 31.340 ;
        RECT 42.190 31.120 44.350 31.290 ;
        RECT 44.590 31.120 44.920 31.290 ;
        RECT 45.210 31.150 45.420 31.480 ;
        RECT 41.640 30.680 41.910 31.120 ;
        RECT 43.120 30.860 43.450 31.120 ;
        RECT 44.660 30.980 44.920 31.120 ;
        RECT 45.660 30.980 45.840 31.420 ;
        RECT 47.260 31.320 47.650 31.370 ;
        RECT 46.390 31.260 47.650 31.320 ;
        RECT 46.390 31.150 47.730 31.260 ;
        RECT 47.260 31.090 47.730 31.150 ;
        RECT 48.200 31.110 49.160 31.280 ;
        RECT 47.260 31.080 47.640 31.090 ;
        RECT 41.680 30.670 41.910 30.680 ;
        RECT 44.660 30.810 45.840 30.980 ;
        RECT 44.660 30.670 44.920 30.810 ;
        RECT 41.680 30.500 42.440 30.670 ;
        RECT 42.690 30.500 43.860 30.670 ;
        RECT 44.100 30.640 44.920 30.670 ;
        RECT 44.100 30.500 45.210 30.640 ;
        RECT 43.090 30.400 43.440 30.500 ;
        RECT 44.750 30.470 45.210 30.500 ;
        RECT 45.660 30.630 46.850 30.640 ;
        RECT 45.660 30.470 47.140 30.630 ;
        RECT 45.700 30.450 47.140 30.470 ;
        RECT 46.680 30.410 47.140 30.450 ;
        RECT 46.850 30.390 47.140 30.410 ;
        RECT 47.470 30.320 47.640 31.080 ;
        RECT 48.980 30.650 49.160 31.110 ;
        RECT 50.060 31.010 50.230 31.360 ;
        RECT 50.000 30.840 50.230 31.010 ;
        RECT 50.400 31.110 50.590 31.150 ;
        RECT 50.400 30.940 50.960 31.110 ;
        RECT 51.420 30.940 54.170 31.110 ;
        RECT 50.400 30.920 50.590 30.940 ;
        RECT 50.060 30.800 50.230 30.840 ;
        RECT 53.350 30.760 53.690 30.940 ;
        RECT 47.840 30.470 48.440 30.640 ;
        RECT 48.900 30.480 49.230 30.650 ;
        RECT 47.840 30.320 48.290 30.470 ;
        RECT 50.130 30.200 50.300 30.620 ;
        RECT 50.940 30.490 51.180 30.530 ;
        RECT 53.720 30.490 53.890 30.500 ;
        RECT 50.610 30.320 51.180 30.490 ;
        RECT 51.420 30.320 52.760 30.490 ;
        RECT 53.210 30.320 54.170 30.490 ;
        RECT 50.940 30.290 51.180 30.320 ;
        RECT 54.700 30.250 54.870 31.180 ;
        RECT 55.100 30.200 55.270 31.090 ;
        RECT 58.000 30.760 58.220 31.350 ;
        RECT 58.000 30.730 58.210 30.760 ;
        RECT 58.740 30.750 58.940 31.350 ;
        RECT 60.750 31.270 60.920 31.800 ;
        RECT 64.690 31.280 64.860 31.810 ;
        RECT 70.480 31.280 70.650 31.810 ;
        RECT 74.420 31.270 74.590 31.800 ;
        RECT 59.750 31.250 60.070 31.260 ;
        RECT 59.490 31.080 60.070 31.250 ;
        RECT 59.740 31.040 60.070 31.080 ;
        RECT 59.750 31.000 60.070 31.040 ;
        RECT 75.270 31.250 75.590 31.260 ;
        RECT 75.270 31.080 75.850 31.250 ;
        RECT 75.270 31.040 75.600 31.080 ;
        RECT 75.270 31.000 75.590 31.040 ;
        RECT 76.400 30.750 76.600 31.350 ;
        RECT 77.120 30.760 77.340 31.350 ;
        RECT 58.010 30.380 58.210 30.730 ;
        RECT 77.130 30.730 77.340 30.760 ;
        RECT 59.750 30.680 60.070 30.710 ;
        RECT 59.740 30.630 60.070 30.680 ;
        RECT 59.490 30.460 60.070 30.630 ;
        RECT 75.270 30.680 75.590 30.710 ;
        RECT 75.270 30.630 75.600 30.680 ;
        RECT 59.750 30.450 60.070 30.460 ;
        RECT 58.380 29.920 58.820 30.090 ;
        RECT 41.090 29.730 41.260 29.780 ;
        RECT 41.060 29.510 41.280 29.730 ;
        RECT 41.090 29.450 41.260 29.510 ;
        RECT 41.610 29.370 41.940 29.550 ;
        RECT 44.750 29.540 44.920 29.590 ;
        RECT 42.190 29.370 44.350 29.540 ;
        RECT 44.590 29.370 44.920 29.540 ;
        RECT 45.210 29.400 45.420 29.730 ;
        RECT 41.640 28.930 41.910 29.370 ;
        RECT 43.120 29.110 43.450 29.370 ;
        RECT 44.660 29.230 44.920 29.370 ;
        RECT 45.660 29.230 45.840 29.670 ;
        RECT 47.260 29.570 47.650 29.620 ;
        RECT 46.390 29.510 47.650 29.570 ;
        RECT 46.390 29.400 47.730 29.510 ;
        RECT 47.260 29.340 47.730 29.400 ;
        RECT 48.200 29.360 49.160 29.530 ;
        RECT 47.260 29.330 47.640 29.340 ;
        RECT 41.680 28.920 41.910 28.930 ;
        RECT 44.660 29.060 45.840 29.230 ;
        RECT 44.660 28.920 44.920 29.060 ;
        RECT 41.680 28.750 42.440 28.920 ;
        RECT 42.690 28.750 43.860 28.920 ;
        RECT 44.100 28.890 44.920 28.920 ;
        RECT 44.100 28.750 45.210 28.890 ;
        RECT 43.090 28.650 43.440 28.750 ;
        RECT 44.750 28.720 45.210 28.750 ;
        RECT 45.660 28.880 46.850 28.890 ;
        RECT 45.660 28.720 47.140 28.880 ;
        RECT 45.700 28.700 47.140 28.720 ;
        RECT 46.680 28.660 47.140 28.700 ;
        RECT 46.850 28.640 47.140 28.660 ;
        RECT 47.470 28.570 47.640 29.330 ;
        RECT 48.980 28.900 49.160 29.360 ;
        RECT 50.130 29.310 50.300 29.730 ;
        RECT 50.940 29.610 51.180 29.640 ;
        RECT 50.610 29.440 51.180 29.610 ;
        RECT 51.420 29.440 52.760 29.610 ;
        RECT 53.210 29.440 54.170 29.610 ;
        RECT 50.940 29.400 51.180 29.440 ;
        RECT 53.720 29.430 53.890 29.440 ;
        RECT 50.060 29.090 50.230 29.130 ;
        RECT 50.000 28.920 50.230 29.090 ;
        RECT 47.840 28.720 48.440 28.890 ;
        RECT 48.900 28.730 49.230 28.900 ;
        RECT 47.840 28.570 48.290 28.720 ;
        RECT 50.060 28.570 50.230 28.920 ;
        RECT 50.400 28.990 50.590 29.010 ;
        RECT 53.350 28.990 53.690 29.170 ;
        RECT 50.400 28.820 50.960 28.990 ;
        RECT 51.420 28.820 54.170 28.990 ;
        RECT 50.400 28.780 50.590 28.820 ;
        RECT 54.700 28.750 54.870 29.680 ;
        RECT 55.100 28.840 55.270 29.730 ;
        RECT 58.010 29.280 58.210 29.630 ;
        RECT 59.750 29.550 60.070 29.560 ;
        RECT 59.490 29.380 60.070 29.550 ;
        RECT 60.750 29.430 60.920 30.440 ;
        RECT 62.680 29.710 63.230 30.140 ;
        RECT 64.680 29.570 64.850 30.580 ;
        RECT 66.710 29.780 67.260 30.210 ;
        RECT 68.080 29.780 68.630 30.210 ;
        RECT 70.490 29.570 70.660 30.580 ;
        RECT 75.270 30.460 75.850 30.630 ;
        RECT 75.270 30.450 75.590 30.460 ;
        RECT 72.110 29.710 72.660 30.140 ;
        RECT 74.420 29.430 74.590 30.440 ;
        RECT 77.130 30.380 77.330 30.730 ;
        RECT 76.520 29.920 76.960 30.090 ;
        RECT 75.270 29.550 75.590 29.560 ;
        RECT 59.740 29.330 60.070 29.380 ;
        RECT 59.750 29.300 60.070 29.330 ;
        RECT 75.270 29.380 75.850 29.550 ;
        RECT 75.270 29.330 75.600 29.380 ;
        RECT 75.270 29.300 75.590 29.330 ;
        RECT 58.000 29.250 58.210 29.280 ;
        RECT 77.130 29.280 77.330 29.630 ;
        RECT 58.000 28.660 58.220 29.250 ;
        RECT 58.740 28.660 58.940 29.260 ;
        RECT 59.750 28.970 60.070 29.010 ;
        RECT 59.740 28.930 60.070 28.970 ;
        RECT 59.490 28.760 60.070 28.930 ;
        RECT 59.750 28.750 60.070 28.760 ;
        RECT 75.270 28.970 75.590 29.010 ;
        RECT 75.270 28.930 75.600 28.970 ;
        RECT 75.270 28.760 75.850 28.930 ;
        RECT 75.270 28.750 75.590 28.760 ;
        RECT 76.400 28.660 76.600 29.260 ;
        RECT 77.130 29.250 77.340 29.280 ;
        RECT 77.120 28.660 77.340 29.250 ;
        RECT 41.090 27.980 41.260 28.030 ;
        RECT 41.060 27.760 41.280 27.980 ;
        RECT 41.090 27.700 41.260 27.760 ;
        RECT 41.610 27.620 41.940 27.800 ;
        RECT 44.750 27.790 44.920 27.840 ;
        RECT 42.190 27.620 44.350 27.790 ;
        RECT 44.590 27.620 44.920 27.790 ;
        RECT 45.210 27.650 45.420 27.980 ;
        RECT 41.640 27.180 41.910 27.620 ;
        RECT 43.120 27.360 43.450 27.620 ;
        RECT 44.660 27.480 44.920 27.620 ;
        RECT 45.660 27.480 45.840 27.920 ;
        RECT 47.260 27.820 47.650 27.870 ;
        RECT 46.390 27.760 47.650 27.820 ;
        RECT 50.060 27.810 50.230 28.160 ;
        RECT 46.390 27.650 47.730 27.760 ;
        RECT 47.260 27.590 47.730 27.650 ;
        RECT 48.200 27.610 49.160 27.780 ;
        RECT 50.000 27.640 50.230 27.810 ;
        RECT 50.400 27.910 50.590 27.950 ;
        RECT 50.400 27.740 50.960 27.910 ;
        RECT 51.420 27.740 54.170 27.910 ;
        RECT 50.400 27.720 50.590 27.740 ;
        RECT 47.260 27.580 47.640 27.590 ;
        RECT 41.680 27.170 41.910 27.180 ;
        RECT 44.660 27.310 45.840 27.480 ;
        RECT 44.660 27.170 44.920 27.310 ;
        RECT 41.680 27.000 42.440 27.170 ;
        RECT 42.690 27.000 43.860 27.170 ;
        RECT 44.100 27.140 44.920 27.170 ;
        RECT 44.100 27.000 45.210 27.140 ;
        RECT 43.090 26.900 43.440 27.000 ;
        RECT 44.750 26.970 45.210 27.000 ;
        RECT 45.660 27.130 46.850 27.140 ;
        RECT 45.660 26.970 47.140 27.130 ;
        RECT 45.700 26.950 47.140 26.970 ;
        RECT 46.680 26.910 47.140 26.950 ;
        RECT 46.850 26.890 47.140 26.910 ;
        RECT 47.470 26.820 47.640 27.580 ;
        RECT 48.980 27.150 49.160 27.610 ;
        RECT 50.060 27.600 50.230 27.640 ;
        RECT 53.350 27.560 53.690 27.740 ;
        RECT 47.840 26.970 48.440 27.140 ;
        RECT 48.900 26.980 49.230 27.150 ;
        RECT 50.130 27.000 50.300 27.420 ;
        RECT 50.940 27.290 51.180 27.330 ;
        RECT 53.720 27.290 53.890 27.300 ;
        RECT 50.610 27.120 51.180 27.290 ;
        RECT 51.420 27.120 52.760 27.290 ;
        RECT 53.210 27.120 54.170 27.290 ;
        RECT 50.940 27.090 51.180 27.120 ;
        RECT 54.700 27.050 54.870 27.980 ;
        RECT 55.100 27.000 55.270 27.890 ;
        RECT 58.000 27.530 58.220 28.120 ;
        RECT 58.000 27.500 58.210 27.530 ;
        RECT 58.740 27.520 58.940 28.120 ;
        RECT 59.750 28.020 60.070 28.030 ;
        RECT 59.490 27.850 60.070 28.020 ;
        RECT 59.740 27.810 60.070 27.850 ;
        RECT 59.750 27.770 60.070 27.810 ;
        RECT 75.270 28.020 75.590 28.030 ;
        RECT 75.270 27.850 75.850 28.020 ;
        RECT 75.270 27.810 75.600 27.850 ;
        RECT 75.270 27.770 75.590 27.810 ;
        RECT 76.400 27.520 76.600 28.120 ;
        RECT 77.120 27.530 77.340 28.120 ;
        RECT 58.010 27.150 58.210 27.500 ;
        RECT 77.130 27.500 77.340 27.530 ;
        RECT 59.750 27.450 60.070 27.480 ;
        RECT 59.740 27.400 60.070 27.450 ;
        RECT 59.490 27.230 60.070 27.400 ;
        RECT 59.750 27.220 60.070 27.230 ;
        RECT 75.270 27.450 75.590 27.480 ;
        RECT 75.270 27.400 75.600 27.450 ;
        RECT 75.270 27.230 75.850 27.400 ;
        RECT 75.270 27.220 75.590 27.230 ;
        RECT 77.130 27.150 77.330 27.500 ;
        RECT 47.840 26.820 48.290 26.970 ;
        RECT 17.760 23.870 17.930 24.360 ;
        RECT 17.610 23.840 17.930 23.870 ;
        RECT 18.310 23.870 18.480 24.360 ;
        RECT 18.950 24.310 19.120 24.360 ;
        RECT 19.500 24.310 19.670 24.360 ;
        RECT 18.830 24.280 19.150 24.310 ;
        RECT 19.480 24.280 19.800 24.310 ;
        RECT 18.830 24.090 19.160 24.280 ;
        RECT 19.480 24.090 19.810 24.280 ;
        RECT 41.050 24.170 41.220 24.220 ;
        RECT 18.830 24.050 19.150 24.090 ;
        RECT 19.480 24.050 19.800 24.090 ;
        RECT 18.310 23.840 18.630 23.870 ;
        RECT 17.610 23.650 17.940 23.840 ;
        RECT 18.310 23.650 18.640 23.840 ;
        RECT 17.610 23.610 17.930 23.650 ;
        RECT 17.220 22.150 17.390 22.170 ;
        RECT 17.200 21.720 17.410 22.150 ;
        RECT 17.760 21.960 17.930 23.610 ;
        RECT 18.310 23.610 18.630 23.650 ;
        RECT 18.310 21.960 18.480 23.610 ;
        RECT 18.950 21.960 19.120 24.050 ;
        RECT 19.500 21.960 19.670 24.050 ;
        RECT 41.020 23.950 41.240 24.170 ;
        RECT 41.050 23.890 41.220 23.950 ;
        RECT 41.570 23.810 41.900 23.990 ;
        RECT 44.710 23.980 44.880 24.030 ;
        RECT 42.150 23.810 44.310 23.980 ;
        RECT 44.550 23.810 44.880 23.980 ;
        RECT 45.170 23.840 45.380 24.170 ;
        RECT 20.050 22.600 20.220 23.450 ;
        RECT 41.600 23.370 41.870 23.810 ;
        RECT 43.080 23.550 43.410 23.810 ;
        RECT 44.620 23.670 44.880 23.810 ;
        RECT 45.620 23.670 45.800 24.110 ;
        RECT 47.220 24.010 47.610 24.060 ;
        RECT 46.350 23.950 47.610 24.010 ;
        RECT 46.350 23.840 47.690 23.950 ;
        RECT 47.220 23.780 47.690 23.840 ;
        RECT 48.160 23.800 49.120 23.970 ;
        RECT 47.220 23.770 47.600 23.780 ;
        RECT 41.640 23.360 41.870 23.370 ;
        RECT 44.620 23.500 45.800 23.670 ;
        RECT 44.620 23.360 44.880 23.500 ;
        RECT 41.640 23.190 42.400 23.360 ;
        RECT 42.650 23.190 43.820 23.360 ;
        RECT 44.060 23.330 44.880 23.360 ;
        RECT 44.060 23.190 45.170 23.330 ;
        RECT 43.050 23.090 43.400 23.190 ;
        RECT 44.710 23.160 45.170 23.190 ;
        RECT 45.620 23.320 46.810 23.330 ;
        RECT 45.620 23.160 47.100 23.320 ;
        RECT 45.660 23.140 47.100 23.160 ;
        RECT 46.640 23.100 47.100 23.140 ;
        RECT 46.810 23.080 47.100 23.100 ;
        RECT 47.430 23.010 47.600 23.770 ;
        RECT 48.940 23.340 49.120 23.800 ;
        RECT 47.800 23.160 48.400 23.330 ;
        RECT 48.860 23.170 49.190 23.340 ;
        RECT 50.160 23.240 50.330 23.660 ;
        RECT 50.970 23.540 51.210 23.570 ;
        RECT 50.640 23.370 51.210 23.540 ;
        RECT 51.450 23.370 52.790 23.540 ;
        RECT 53.240 23.370 54.200 23.540 ;
        RECT 50.970 23.330 51.210 23.370 ;
        RECT 53.750 23.360 53.920 23.370 ;
        RECT 47.800 23.010 48.250 23.160 ;
        RECT 50.090 23.020 50.260 23.060 ;
        RECT 50.030 22.850 50.260 23.020 ;
        RECT 50.090 22.500 50.260 22.850 ;
        RECT 50.430 22.920 50.620 22.940 ;
        RECT 53.380 22.920 53.720 23.100 ;
        RECT 50.430 22.750 50.990 22.920 ;
        RECT 51.450 22.750 54.200 22.920 ;
        RECT 50.430 22.710 50.620 22.750 ;
        RECT 54.730 22.680 54.900 23.610 ;
        RECT 55.130 22.770 55.300 23.660 ;
        RECT 58.040 23.190 58.240 23.540 ;
        RECT 59.780 23.460 60.100 23.470 ;
        RECT 59.520 23.290 60.100 23.460 ;
        RECT 59.770 23.240 60.100 23.290 ;
        RECT 59.780 23.210 60.100 23.240 ;
        RECT 58.030 23.160 58.240 23.190 ;
        RECT 58.030 22.570 58.250 23.160 ;
        RECT 58.770 22.570 58.970 23.170 ;
        RECT 68.490 23.140 68.810 23.170 ;
        RECT 68.490 22.970 70.280 23.140 ;
        RECT 68.490 22.950 68.820 22.970 ;
        RECT 59.780 22.880 60.100 22.920 ;
        RECT 68.490 22.910 68.810 22.950 ;
        RECT 59.770 22.840 60.100 22.880 ;
        RECT 59.520 22.670 60.100 22.840 ;
        RECT 70.110 22.740 70.280 22.970 ;
        RECT 59.780 22.660 60.100 22.670 ;
        RECT 68.960 22.490 69.300 22.740 ;
        RECT 69.470 22.570 69.800 22.740 ;
        RECT 70.020 22.570 70.360 22.740 ;
        RECT 41.050 22.420 41.220 22.470 ;
        RECT 41.020 22.200 41.240 22.420 ;
        RECT 41.050 22.140 41.220 22.200 ;
        RECT 41.570 22.060 41.900 22.240 ;
        RECT 44.710 22.230 44.880 22.280 ;
        RECT 42.150 22.060 44.310 22.230 ;
        RECT 44.550 22.060 44.880 22.230 ;
        RECT 45.170 22.090 45.380 22.420 ;
        RECT 19.940 21.970 20.370 21.990 ;
        RECT 19.940 21.800 20.390 21.970 ;
        RECT 19.940 21.780 20.370 21.800 ;
        RECT 41.600 21.620 41.870 22.060 ;
        RECT 43.080 21.800 43.410 22.060 ;
        RECT 44.620 21.920 44.880 22.060 ;
        RECT 45.620 21.920 45.800 22.360 ;
        RECT 47.220 22.260 47.610 22.310 ;
        RECT 46.350 22.200 47.610 22.260 ;
        RECT 46.350 22.090 47.690 22.200 ;
        RECT 47.220 22.030 47.690 22.090 ;
        RECT 48.160 22.050 49.120 22.220 ;
        RECT 47.220 22.020 47.600 22.030 ;
        RECT 41.640 21.610 41.870 21.620 ;
        RECT 44.620 21.750 45.800 21.920 ;
        RECT 44.620 21.610 44.880 21.750 ;
        RECT 17.210 21.080 17.420 21.510 ;
        RECT 19.950 21.430 20.380 21.450 ;
        RECT 41.640 21.440 42.400 21.610 ;
        RECT 42.650 21.440 43.820 21.610 ;
        RECT 44.060 21.580 44.880 21.610 ;
        RECT 44.060 21.440 45.170 21.580 ;
        RECT 17.230 21.060 17.400 21.080 ;
        RECT 17.770 19.990 17.940 21.310 ;
        RECT 17.640 19.960 17.960 19.990 ;
        RECT 18.320 19.980 18.490 21.320 ;
        RECT 17.640 19.770 17.970 19.960 ;
        RECT 18.320 19.950 18.650 19.980 ;
        RECT 17.640 19.730 17.960 19.770 ;
        RECT 18.320 19.760 18.660 19.950 ;
        RECT 17.770 18.820 17.940 19.730 ;
        RECT 18.320 19.720 18.650 19.760 ;
        RECT 18.320 18.820 18.490 19.720 ;
        RECT 18.950 19.210 19.120 21.310 ;
        RECT 18.810 19.180 19.130 19.210 ;
        RECT 18.810 18.990 19.140 19.180 ;
        RECT 19.500 19.150 19.670 21.320 ;
        RECT 19.950 21.260 20.400 21.430 ;
        RECT 43.050 21.340 43.400 21.440 ;
        RECT 44.710 21.410 45.170 21.440 ;
        RECT 45.620 21.570 46.810 21.580 ;
        RECT 45.620 21.410 47.100 21.570 ;
        RECT 45.660 21.390 47.100 21.410 ;
        RECT 46.640 21.350 47.100 21.390 ;
        RECT 46.810 21.330 47.100 21.350 ;
        RECT 47.430 21.260 47.600 22.020 ;
        RECT 48.940 21.590 49.120 22.050 ;
        RECT 50.090 21.740 50.260 22.090 ;
        RECT 47.800 21.410 48.400 21.580 ;
        RECT 48.860 21.420 49.190 21.590 ;
        RECT 50.030 21.570 50.260 21.740 ;
        RECT 50.430 21.840 50.620 21.880 ;
        RECT 50.430 21.670 50.990 21.840 ;
        RECT 51.450 21.670 54.200 21.840 ;
        RECT 50.430 21.650 50.620 21.670 ;
        RECT 50.090 21.530 50.260 21.570 ;
        RECT 53.380 21.490 53.720 21.670 ;
        RECT 47.800 21.260 48.250 21.410 ;
        RECT 19.950 21.240 20.380 21.260 ;
        RECT 50.160 20.930 50.330 21.350 ;
        RECT 50.970 21.220 51.210 21.260 ;
        RECT 53.750 21.220 53.920 21.230 ;
        RECT 50.640 21.050 51.210 21.220 ;
        RECT 51.450 21.050 52.790 21.220 ;
        RECT 53.240 21.050 54.200 21.220 ;
        RECT 50.970 21.020 51.210 21.050 ;
        RECT 54.730 20.980 54.900 21.910 ;
        RECT 55.130 20.930 55.300 21.820 ;
        RECT 58.030 21.450 58.250 22.040 ;
        RECT 58.030 21.420 58.240 21.450 ;
        RECT 58.770 21.440 58.970 22.040 ;
        RECT 59.780 21.940 60.100 21.950 ;
        RECT 59.520 21.770 60.100 21.940 ;
        RECT 60.910 21.880 61.080 22.410 ;
        RECT 64.930 21.910 65.100 22.440 ;
        RECT 68.640 22.230 69.300 22.490 ;
        RECT 69.550 22.400 69.720 22.570 ;
        RECT 70.110 22.400 70.280 22.570 ;
        RECT 69.470 22.230 69.800 22.400 ;
        RECT 70.020 22.230 70.360 22.400 ;
        RECT 69.550 22.000 69.800 22.230 ;
        RECT 70.680 22.150 71.190 22.820 ;
        RECT 59.770 21.730 60.100 21.770 ;
        RECT 59.780 21.690 60.100 21.730 ;
        RECT 69.550 21.830 70.220 22.000 ;
        RECT 69.550 21.600 69.800 21.830 ;
        RECT 58.040 21.070 58.240 21.420 ;
        RECT 59.780 21.370 60.100 21.400 ;
        RECT 59.770 21.320 60.100 21.370 ;
        RECT 68.640 21.340 69.300 21.600 ;
        RECT 69.470 21.430 69.800 21.600 ;
        RECT 70.020 21.430 70.360 21.600 ;
        RECT 59.520 21.150 60.100 21.320 ;
        RECT 59.780 21.140 60.100 21.150 ;
        RECT 20.040 20.050 20.210 20.720 ;
        RECT 41.050 20.670 41.220 20.720 ;
        RECT 41.020 20.450 41.240 20.670 ;
        RECT 41.050 20.390 41.220 20.450 ;
        RECT 41.570 20.310 41.900 20.490 ;
        RECT 44.710 20.480 44.880 20.530 ;
        RECT 42.150 20.310 44.310 20.480 ;
        RECT 44.550 20.310 44.880 20.480 ;
        RECT 45.170 20.340 45.380 20.670 ;
        RECT 58.410 20.610 58.850 20.780 ;
        RECT 41.600 19.870 41.870 20.310 ;
        RECT 43.080 20.050 43.410 20.310 ;
        RECT 44.620 20.170 44.880 20.310 ;
        RECT 45.620 20.170 45.800 20.610 ;
        RECT 47.220 20.510 47.610 20.560 ;
        RECT 46.350 20.450 47.610 20.510 ;
        RECT 46.350 20.340 47.690 20.450 ;
        RECT 47.220 20.280 47.690 20.340 ;
        RECT 48.160 20.300 49.120 20.470 ;
        RECT 47.220 20.270 47.600 20.280 ;
        RECT 41.640 19.860 41.870 19.870 ;
        RECT 44.620 20.000 45.800 20.170 ;
        RECT 44.620 19.860 44.880 20.000 ;
        RECT 41.640 19.690 42.400 19.860 ;
        RECT 42.650 19.690 43.820 19.860 ;
        RECT 44.060 19.830 44.880 19.860 ;
        RECT 44.060 19.690 45.170 19.830 ;
        RECT 43.050 19.590 43.400 19.690 ;
        RECT 44.710 19.660 45.170 19.690 ;
        RECT 45.620 19.820 46.810 19.830 ;
        RECT 45.620 19.660 47.100 19.820 ;
        RECT 45.660 19.640 47.100 19.660 ;
        RECT 46.640 19.600 47.100 19.640 ;
        RECT 46.810 19.580 47.100 19.600 ;
        RECT 47.430 19.510 47.600 20.270 ;
        RECT 48.940 19.840 49.120 20.300 ;
        RECT 50.160 20.040 50.330 20.460 ;
        RECT 50.970 20.340 51.210 20.370 ;
        RECT 50.640 20.170 51.210 20.340 ;
        RECT 51.450 20.170 52.790 20.340 ;
        RECT 53.240 20.170 54.200 20.340 ;
        RECT 50.970 20.130 51.210 20.170 ;
        RECT 53.750 20.160 53.920 20.170 ;
        RECT 47.800 19.660 48.400 19.830 ;
        RECT 48.860 19.670 49.190 19.840 ;
        RECT 50.090 19.820 50.260 19.860 ;
        RECT 47.800 19.510 48.250 19.660 ;
        RECT 50.030 19.650 50.260 19.820 ;
        RECT 50.090 19.300 50.260 19.650 ;
        RECT 50.430 19.720 50.620 19.740 ;
        RECT 53.380 19.720 53.720 19.900 ;
        RECT 50.430 19.550 50.990 19.720 ;
        RECT 51.450 19.550 54.200 19.720 ;
        RECT 50.430 19.510 50.620 19.550 ;
        RECT 54.730 19.480 54.900 20.410 ;
        RECT 55.130 19.570 55.300 20.460 ;
        RECT 58.040 19.950 58.240 20.300 ;
        RECT 59.780 20.220 60.100 20.230 ;
        RECT 59.520 20.050 60.100 20.220 ;
        RECT 59.770 20.000 60.100 20.050 ;
        RECT 60.900 20.020 61.070 21.210 ;
        RECT 62.710 20.340 63.260 20.770 ;
        RECT 59.780 19.970 60.100 20.000 ;
        RECT 64.920 19.980 65.090 21.150 ;
        RECT 68.960 21.090 69.300 21.340 ;
        RECT 69.550 21.260 69.720 21.430 ;
        RECT 70.110 21.260 70.280 21.430 ;
        RECT 69.470 21.090 69.800 21.260 ;
        RECT 70.020 21.090 70.360 21.260 ;
        RECT 68.490 20.880 68.810 20.920 ;
        RECT 68.490 20.860 68.820 20.880 ;
        RECT 70.110 20.860 70.280 21.090 ;
        RECT 70.680 21.010 71.190 21.680 ;
        RECT 66.740 20.410 67.290 20.840 ;
        RECT 68.490 20.690 70.280 20.860 ;
        RECT 68.490 20.660 68.810 20.690 ;
        RECT 68.490 20.370 68.810 20.400 ;
        RECT 68.490 20.200 70.280 20.370 ;
        RECT 68.490 20.180 68.820 20.200 ;
        RECT 68.490 20.140 68.810 20.180 ;
        RECT 70.110 19.970 70.280 20.200 ;
        RECT 58.030 19.920 58.240 19.950 ;
        RECT 58.030 19.330 58.250 19.920 ;
        RECT 58.770 19.330 58.970 19.930 ;
        RECT 68.960 19.720 69.300 19.970 ;
        RECT 69.470 19.800 69.800 19.970 ;
        RECT 70.020 19.800 70.360 19.970 ;
        RECT 59.780 19.640 60.100 19.680 ;
        RECT 59.770 19.600 60.100 19.640 ;
        RECT 59.520 19.430 60.100 19.600 ;
        RECT 68.640 19.460 69.300 19.720 ;
        RECT 69.550 19.630 69.720 19.800 ;
        RECT 70.110 19.630 70.280 19.800 ;
        RECT 69.470 19.460 69.800 19.630 ;
        RECT 70.020 19.460 70.360 19.630 ;
        RECT 59.780 19.420 60.100 19.430 ;
        RECT 69.550 19.230 69.800 19.460 ;
        RECT 70.680 19.380 71.190 20.050 ;
        RECT 19.500 19.120 19.840 19.150 ;
        RECT 18.810 18.950 19.130 18.990 ;
        RECT 18.950 18.820 19.120 18.950 ;
        RECT 19.500 18.930 19.850 19.120 ;
        RECT 69.550 19.060 70.220 19.230 ;
        RECT 19.500 18.890 19.840 18.930 ;
        RECT 41.050 18.920 41.220 18.970 ;
        RECT 19.500 18.820 19.670 18.890 ;
        RECT 41.020 18.700 41.240 18.920 ;
        RECT 41.050 18.640 41.220 18.700 ;
        RECT 41.570 18.560 41.900 18.740 ;
        RECT 44.710 18.730 44.880 18.780 ;
        RECT 42.150 18.560 44.310 18.730 ;
        RECT 44.550 18.560 44.880 18.730 ;
        RECT 45.170 18.590 45.380 18.920 ;
        RECT 41.600 18.120 41.870 18.560 ;
        RECT 43.080 18.300 43.410 18.560 ;
        RECT 44.620 18.420 44.880 18.560 ;
        RECT 45.620 18.420 45.800 18.860 ;
        RECT 47.220 18.760 47.610 18.810 ;
        RECT 46.350 18.700 47.610 18.760 ;
        RECT 46.350 18.590 47.690 18.700 ;
        RECT 47.220 18.530 47.690 18.590 ;
        RECT 48.160 18.550 49.120 18.720 ;
        RECT 47.220 18.520 47.600 18.530 ;
        RECT 41.640 18.110 41.870 18.120 ;
        RECT 44.620 18.250 45.800 18.420 ;
        RECT 44.620 18.110 44.880 18.250 ;
        RECT 41.640 17.940 42.400 18.110 ;
        RECT 42.650 17.940 43.820 18.110 ;
        RECT 44.060 18.080 44.880 18.110 ;
        RECT 44.060 17.940 45.170 18.080 ;
        RECT 43.050 17.840 43.400 17.940 ;
        RECT 44.710 17.910 45.170 17.940 ;
        RECT 45.620 18.070 46.810 18.080 ;
        RECT 45.620 17.910 47.100 18.070 ;
        RECT 45.660 17.890 47.100 17.910 ;
        RECT 46.640 17.850 47.100 17.890 ;
        RECT 46.810 17.830 47.100 17.850 ;
        RECT 47.430 17.760 47.600 18.520 ;
        RECT 48.940 18.090 49.120 18.550 ;
        RECT 50.090 18.540 50.260 18.890 ;
        RECT 69.550 18.830 69.800 19.060 ;
        RECT 57.050 18.730 57.370 18.770 ;
        RECT 50.030 18.370 50.260 18.540 ;
        RECT 50.430 18.640 50.620 18.680 ;
        RECT 50.430 18.470 50.990 18.640 ;
        RECT 51.450 18.470 54.200 18.640 ;
        RECT 50.430 18.450 50.620 18.470 ;
        RECT 50.090 18.330 50.260 18.370 ;
        RECT 53.380 18.290 53.720 18.470 ;
        RECT 47.800 17.910 48.400 18.080 ;
        RECT 48.860 17.920 49.190 18.090 ;
        RECT 47.800 17.760 48.250 17.910 ;
        RECT 50.160 17.730 50.330 18.150 ;
        RECT 50.970 18.020 51.210 18.060 ;
        RECT 53.750 18.020 53.920 18.030 ;
        RECT 50.640 17.850 51.210 18.020 ;
        RECT 51.450 17.850 52.790 18.020 ;
        RECT 53.240 17.850 54.200 18.020 ;
        RECT 50.970 17.820 51.210 17.850 ;
        RECT 54.730 17.780 54.900 18.710 ;
        RECT 55.130 17.730 55.300 18.620 ;
        RECT 57.050 18.540 57.380 18.730 ;
        RECT 57.050 18.510 57.370 18.540 ;
        RECT 57.100 17.810 57.280 18.510 ;
        RECT 58.030 18.200 58.250 18.790 ;
        RECT 58.030 18.170 58.240 18.200 ;
        RECT 58.770 18.190 58.970 18.790 ;
        RECT 59.780 18.690 60.100 18.700 ;
        RECT 59.520 18.520 60.100 18.690 ;
        RECT 68.640 18.570 69.300 18.830 ;
        RECT 69.470 18.660 69.800 18.830 ;
        RECT 70.020 18.660 70.360 18.830 ;
        RECT 59.770 18.480 60.100 18.520 ;
        RECT 59.780 18.440 60.100 18.480 ;
        RECT 68.960 18.320 69.300 18.570 ;
        RECT 69.550 18.490 69.720 18.660 ;
        RECT 70.110 18.490 70.280 18.660 ;
        RECT 69.470 18.320 69.800 18.490 ;
        RECT 70.020 18.320 70.360 18.490 ;
        RECT 58.040 17.820 58.240 18.170 ;
        RECT 59.780 18.120 60.100 18.150 ;
        RECT 59.770 18.070 60.100 18.120 ;
        RECT 59.520 17.900 60.100 18.070 ;
        RECT 59.780 17.890 60.100 17.900 ;
        RECT 68.490 18.110 68.810 18.150 ;
        RECT 68.490 18.090 68.820 18.110 ;
        RECT 70.110 18.090 70.280 18.320 ;
        RECT 70.680 18.240 71.190 18.910 ;
        RECT 68.490 17.920 70.280 18.090 ;
        RECT 68.490 17.890 68.810 17.920 ;
        RECT 57.100 17.770 57.420 17.810 ;
        RECT 57.100 17.580 57.430 17.770 ;
        RECT 57.100 17.550 57.420 17.580 ;
        RECT 49.840 15.810 50.010 15.900 ;
        RECT 49.760 15.770 50.080 15.810 ;
        RECT 49.760 15.580 50.090 15.770 ;
        RECT 49.760 15.550 50.080 15.580 ;
        RECT 15.570 13.690 15.740 13.760 ;
        RECT 15.500 13.660 15.820 13.690 ;
        RECT 15.490 13.470 15.820 13.660 ;
        RECT 15.500 13.430 15.820 13.470 ;
        RECT 15.570 10.920 15.740 13.430 ;
        RECT 16.120 13.020 16.290 13.760 ;
        RECT 16.670 13.700 16.840 13.760 ;
        RECT 16.600 13.670 16.920 13.700 ;
        RECT 16.590 13.480 16.920 13.670 ;
        RECT 16.600 13.440 16.920 13.480 ;
        RECT 16.050 12.990 16.370 13.020 ;
        RECT 16.040 12.800 16.370 12.990 ;
        RECT 16.050 12.760 16.370 12.800 ;
        RECT 16.120 11.650 16.290 12.760 ;
        RECT 16.050 11.620 16.370 11.650 ;
        RECT 16.040 11.430 16.370 11.620 ;
        RECT 16.050 11.390 16.370 11.430 ;
        RECT 15.500 10.890 15.820 10.920 ;
        RECT 15.490 10.700 15.820 10.890 ;
        RECT 15.500 10.660 15.820 10.700 ;
        RECT 15.570 9.580 15.740 10.660 ;
        RECT 15.490 9.550 15.810 9.580 ;
        RECT 15.480 9.360 15.810 9.550 ;
        RECT 15.490 9.320 15.810 9.360 ;
        RECT 15.570 8.580 15.740 9.320 ;
        RECT 16.120 8.880 16.290 11.390 ;
        RECT 16.670 10.920 16.840 13.440 ;
        RECT 17.220 13.020 17.390 13.760 ;
        RECT 17.770 13.700 17.940 13.760 ;
        RECT 17.690 13.670 18.010 13.700 ;
        RECT 17.680 13.480 18.010 13.670 ;
        RECT 17.690 13.440 18.010 13.480 ;
        RECT 17.150 12.990 17.470 13.020 ;
        RECT 17.140 12.800 17.470 12.990 ;
        RECT 17.150 12.760 17.470 12.800 ;
        RECT 17.220 11.650 17.390 12.760 ;
        RECT 17.150 11.620 17.470 11.650 ;
        RECT 17.140 11.430 17.470 11.620 ;
        RECT 17.150 11.390 17.470 11.430 ;
        RECT 16.600 10.890 16.920 10.920 ;
        RECT 16.590 10.700 16.920 10.890 ;
        RECT 16.600 10.660 16.920 10.700 ;
        RECT 16.670 9.570 16.840 10.660 ;
        RECT 16.600 9.540 16.920 9.570 ;
        RECT 16.590 9.350 16.920 9.540 ;
        RECT 16.600 9.310 16.920 9.350 ;
        RECT 16.050 8.850 16.370 8.880 ;
        RECT 16.040 8.660 16.370 8.850 ;
        RECT 16.050 8.620 16.370 8.660 ;
        RECT 16.120 8.580 16.290 8.620 ;
        RECT 16.670 8.580 16.840 9.310 ;
        RECT 17.220 8.870 17.390 11.390 ;
        RECT 17.770 10.920 17.940 13.440 ;
        RECT 18.320 13.020 18.490 13.760 ;
        RECT 18.730 13.480 19.240 14.160 ;
        RECT 26.000 13.660 26.760 14.080 ;
        RECT 18.730 13.410 19.250 13.480 ;
        RECT 18.740 13.150 19.250 13.410 ;
        RECT 18.250 12.990 18.570 13.020 ;
        RECT 18.240 12.800 18.570 12.990 ;
        RECT 18.250 12.760 18.570 12.800 ;
        RECT 18.320 11.650 18.490 12.760 ;
        RECT 19.030 11.740 19.200 12.960 ;
        RECT 26.020 12.870 26.760 13.660 ;
        RECT 49.840 13.030 50.010 15.550 ;
        RECT 50.390 15.130 50.560 15.900 ;
        RECT 50.940 15.810 51.110 15.900 ;
        RECT 50.850 15.770 51.170 15.810 ;
        RECT 50.850 15.580 51.180 15.770 ;
        RECT 50.850 15.550 51.170 15.580 ;
        RECT 50.310 15.090 50.630 15.130 ;
        RECT 50.310 14.900 50.640 15.090 ;
        RECT 50.310 14.870 50.630 14.900 ;
        RECT 50.390 13.760 50.560 14.870 ;
        RECT 50.310 13.720 50.630 13.760 ;
        RECT 50.310 13.530 50.640 13.720 ;
        RECT 50.310 13.500 50.630 13.530 ;
        RECT 49.750 12.990 50.070 13.030 ;
        RECT 49.750 12.800 50.080 12.990 ;
        RECT 49.750 12.770 50.070 12.800 ;
        RECT 49.840 11.660 50.010 12.770 ;
        RECT 18.250 11.620 18.570 11.650 ;
        RECT 18.240 11.430 18.570 11.620 ;
        RECT 18.250 11.390 18.570 11.430 ;
        RECT 49.750 11.620 50.070 11.660 ;
        RECT 49.750 11.430 50.080 11.620 ;
        RECT 49.750 11.400 50.070 11.430 ;
        RECT 17.690 10.890 18.010 10.920 ;
        RECT 17.680 10.700 18.010 10.890 ;
        RECT 17.690 10.660 18.010 10.700 ;
        RECT 17.770 9.550 17.940 10.660 ;
        RECT 17.690 9.520 18.010 9.550 ;
        RECT 17.680 9.330 18.010 9.520 ;
        RECT 17.690 9.290 18.010 9.330 ;
        RECT 17.150 8.840 17.470 8.870 ;
        RECT 17.140 8.650 17.470 8.840 ;
        RECT 17.150 8.610 17.470 8.650 ;
        RECT 17.220 8.580 17.390 8.610 ;
        RECT 17.770 8.580 17.940 9.290 ;
        RECT 18.320 8.870 18.490 11.390 ;
        RECT 49.070 11.190 49.580 11.270 ;
        RECT 49.070 10.940 49.590 11.190 ;
        RECT 49.080 10.260 49.590 10.940 ;
        RECT 49.840 10.580 50.010 11.400 ;
        RECT 50.390 10.980 50.560 13.500 ;
        RECT 50.940 13.030 51.110 15.550 ;
        RECT 51.490 15.110 51.660 15.900 ;
        RECT 52.040 15.800 52.210 15.900 ;
        RECT 51.950 15.760 52.270 15.800 ;
        RECT 51.950 15.570 52.280 15.760 ;
        RECT 51.950 15.540 52.270 15.570 ;
        RECT 51.400 15.070 51.720 15.110 ;
        RECT 51.400 14.880 51.730 15.070 ;
        RECT 51.400 14.850 51.720 14.880 ;
        RECT 51.490 13.760 51.660 14.850 ;
        RECT 51.400 13.720 51.720 13.760 ;
        RECT 51.400 13.530 51.730 13.720 ;
        RECT 51.400 13.500 51.720 13.530 ;
        RECT 50.850 12.990 51.170 13.030 ;
        RECT 50.850 12.800 51.180 12.990 ;
        RECT 50.850 12.770 51.170 12.800 ;
        RECT 50.940 11.660 51.110 12.770 ;
        RECT 50.850 11.620 51.170 11.660 ;
        RECT 50.850 11.430 51.180 11.620 ;
        RECT 50.850 11.400 51.170 11.430 ;
        RECT 50.310 10.940 50.630 10.980 ;
        RECT 50.310 10.750 50.640 10.940 ;
        RECT 50.310 10.720 50.630 10.750 ;
        RECT 50.390 10.570 50.560 10.720 ;
        RECT 50.940 10.570 51.110 11.400 ;
        RECT 51.490 10.980 51.660 13.500 ;
        RECT 52.040 13.030 52.210 15.540 ;
        RECT 52.590 15.100 52.760 15.900 ;
        RECT 53.130 15.170 53.300 15.930 ;
        RECT 53.740 15.170 53.910 15.930 ;
        RECT 54.280 15.100 54.450 15.900 ;
        RECT 54.830 15.800 55.000 15.900 ;
        RECT 54.770 15.760 55.090 15.800 ;
        RECT 54.760 15.570 55.090 15.760 ;
        RECT 54.770 15.540 55.090 15.570 ;
        RECT 52.510 15.060 52.830 15.100 ;
        RECT 54.210 15.060 54.530 15.100 ;
        RECT 52.510 14.870 52.840 15.060 ;
        RECT 54.200 14.870 54.530 15.060 ;
        RECT 52.510 14.840 52.830 14.870 ;
        RECT 54.210 14.840 54.530 14.870 ;
        RECT 52.590 13.760 52.760 14.840 ;
        RECT 54.280 13.760 54.450 14.840 ;
        RECT 52.500 13.720 52.820 13.760 ;
        RECT 54.220 13.720 54.540 13.760 ;
        RECT 52.500 13.530 52.830 13.720 ;
        RECT 54.210 13.530 54.540 13.720 ;
        RECT 52.500 13.500 52.820 13.530 ;
        RECT 54.220 13.500 54.540 13.530 ;
        RECT 51.950 12.990 52.270 13.030 ;
        RECT 51.950 12.800 52.280 12.990 ;
        RECT 51.950 12.770 52.270 12.800 ;
        RECT 52.040 11.660 52.210 12.770 ;
        RECT 51.950 11.620 52.270 11.660 ;
        RECT 51.950 11.430 52.280 11.620 ;
        RECT 51.950 11.400 52.270 11.430 ;
        RECT 51.400 10.940 51.720 10.980 ;
        RECT 51.400 10.750 51.730 10.940 ;
        RECT 51.400 10.720 51.720 10.750 ;
        RECT 51.490 10.570 51.660 10.720 ;
        RECT 52.040 10.570 52.210 11.400 ;
        RECT 52.590 10.990 52.760 13.500 ;
        RECT 54.280 10.990 54.450 13.500 ;
        RECT 54.830 13.030 55.000 15.540 ;
        RECT 55.380 15.110 55.550 15.900 ;
        RECT 55.930 15.810 56.100 15.900 ;
        RECT 55.870 15.770 56.190 15.810 ;
        RECT 55.860 15.580 56.190 15.770 ;
        RECT 55.870 15.550 56.190 15.580 ;
        RECT 55.320 15.070 55.640 15.110 ;
        RECT 55.310 14.880 55.640 15.070 ;
        RECT 55.320 14.850 55.640 14.880 ;
        RECT 55.380 13.760 55.550 14.850 ;
        RECT 55.320 13.720 55.640 13.760 ;
        RECT 55.310 13.530 55.640 13.720 ;
        RECT 55.320 13.500 55.640 13.530 ;
        RECT 54.770 12.990 55.090 13.030 ;
        RECT 54.760 12.800 55.090 12.990 ;
        RECT 54.770 12.770 55.090 12.800 ;
        RECT 54.830 11.660 55.000 12.770 ;
        RECT 54.770 11.620 55.090 11.660 ;
        RECT 54.760 11.430 55.090 11.620 ;
        RECT 54.770 11.400 55.090 11.430 ;
        RECT 52.500 10.950 52.820 10.990 ;
        RECT 54.220 10.950 54.540 10.990 ;
        RECT 52.500 10.760 52.830 10.950 ;
        RECT 54.210 10.760 54.540 10.950 ;
        RECT 52.500 10.730 52.820 10.760 ;
        RECT 54.220 10.730 54.540 10.760 ;
        RECT 52.590 10.570 52.760 10.730 ;
        RECT 54.280 10.570 54.450 10.730 ;
        RECT 54.830 10.570 55.000 11.400 ;
        RECT 55.380 10.980 55.550 13.500 ;
        RECT 55.930 13.030 56.100 15.550 ;
        RECT 56.480 15.130 56.650 15.900 ;
        RECT 57.030 15.810 57.200 15.900 ;
        RECT 59.650 15.840 59.820 15.930 ;
        RECT 56.960 15.770 57.280 15.810 ;
        RECT 56.950 15.580 57.280 15.770 ;
        RECT 59.570 15.800 59.890 15.840 ;
        RECT 59.570 15.610 59.900 15.800 ;
        RECT 59.570 15.580 59.890 15.610 ;
        RECT 56.960 15.550 57.280 15.580 ;
        RECT 56.410 15.090 56.730 15.130 ;
        RECT 56.400 14.900 56.730 15.090 ;
        RECT 56.410 14.870 56.730 14.900 ;
        RECT 56.480 13.760 56.650 14.870 ;
        RECT 56.410 13.720 56.730 13.760 ;
        RECT 56.400 13.530 56.730 13.720 ;
        RECT 56.410 13.500 56.730 13.530 ;
        RECT 55.870 12.990 56.190 13.030 ;
        RECT 55.860 12.800 56.190 12.990 ;
        RECT 55.870 12.770 56.190 12.800 ;
        RECT 55.930 11.660 56.100 12.770 ;
        RECT 55.870 11.620 56.190 11.660 ;
        RECT 55.860 11.430 56.190 11.620 ;
        RECT 55.870 11.400 56.190 11.430 ;
        RECT 55.320 10.940 55.640 10.980 ;
        RECT 55.310 10.750 55.640 10.940 ;
        RECT 55.320 10.720 55.640 10.750 ;
        RECT 55.380 10.570 55.550 10.720 ;
        RECT 55.930 10.570 56.100 11.400 ;
        RECT 56.480 10.980 56.650 13.500 ;
        RECT 57.030 13.030 57.200 15.550 ;
        RECT 59.650 13.060 59.820 15.580 ;
        RECT 60.200 15.160 60.370 15.930 ;
        RECT 60.750 15.840 60.920 15.930 ;
        RECT 60.660 15.800 60.980 15.840 ;
        RECT 60.660 15.610 60.990 15.800 ;
        RECT 60.660 15.580 60.980 15.610 ;
        RECT 60.120 15.120 60.440 15.160 ;
        RECT 60.120 14.930 60.450 15.120 ;
        RECT 60.120 14.900 60.440 14.930 ;
        RECT 60.200 13.790 60.370 14.900 ;
        RECT 60.120 13.750 60.440 13.790 ;
        RECT 60.120 13.560 60.450 13.750 ;
        RECT 60.120 13.530 60.440 13.560 ;
        RECT 56.970 12.990 57.290 13.030 ;
        RECT 56.960 12.800 57.290 12.990 ;
        RECT 59.560 13.020 59.880 13.060 ;
        RECT 59.560 12.830 59.890 13.020 ;
        RECT 59.560 12.800 59.880 12.830 ;
        RECT 56.970 12.770 57.290 12.800 ;
        RECT 57.030 11.660 57.200 12.770 ;
        RECT 59.650 11.690 59.820 12.800 ;
        RECT 56.970 11.620 57.290 11.660 ;
        RECT 56.960 11.430 57.290 11.620 ;
        RECT 59.560 11.650 59.880 11.690 ;
        RECT 59.560 11.460 59.890 11.650 ;
        RECT 59.560 11.430 59.880 11.460 ;
        RECT 56.970 11.400 57.290 11.430 ;
        RECT 56.410 10.940 56.730 10.980 ;
        RECT 56.400 10.750 56.730 10.940 ;
        RECT 56.410 10.720 56.730 10.750 ;
        RECT 56.480 10.570 56.650 10.720 ;
        RECT 57.030 10.580 57.200 11.400 ;
        RECT 57.460 11.190 57.970 11.270 ;
        RECT 57.450 10.940 57.970 11.190 ;
        RECT 58.880 11.220 59.390 11.300 ;
        RECT 58.880 10.970 59.400 11.220 ;
        RECT 57.450 10.260 57.960 10.940 ;
        RECT 58.890 10.290 59.400 10.970 ;
        RECT 59.650 10.610 59.820 11.430 ;
        RECT 60.200 11.010 60.370 13.530 ;
        RECT 60.750 13.060 60.920 15.580 ;
        RECT 61.300 15.140 61.470 15.930 ;
        RECT 61.850 15.830 62.020 15.930 ;
        RECT 61.760 15.790 62.080 15.830 ;
        RECT 61.760 15.600 62.090 15.790 ;
        RECT 61.760 15.570 62.080 15.600 ;
        RECT 61.210 15.100 61.530 15.140 ;
        RECT 61.210 14.910 61.540 15.100 ;
        RECT 61.210 14.880 61.530 14.910 ;
        RECT 61.300 13.790 61.470 14.880 ;
        RECT 61.210 13.750 61.530 13.790 ;
        RECT 61.210 13.560 61.540 13.750 ;
        RECT 61.210 13.530 61.530 13.560 ;
        RECT 60.660 13.020 60.980 13.060 ;
        RECT 60.660 12.830 60.990 13.020 ;
        RECT 60.660 12.800 60.980 12.830 ;
        RECT 60.750 11.690 60.920 12.800 ;
        RECT 60.660 11.650 60.980 11.690 ;
        RECT 60.660 11.460 60.990 11.650 ;
        RECT 60.660 11.430 60.980 11.460 ;
        RECT 60.120 10.970 60.440 11.010 ;
        RECT 60.120 10.780 60.450 10.970 ;
        RECT 60.120 10.750 60.440 10.780 ;
        RECT 60.200 10.600 60.370 10.750 ;
        RECT 60.750 10.600 60.920 11.430 ;
        RECT 61.300 11.010 61.470 13.530 ;
        RECT 61.850 13.060 62.020 15.570 ;
        RECT 62.400 15.130 62.570 15.930 ;
        RECT 62.940 15.200 63.110 15.960 ;
        RECT 63.550 15.200 63.720 15.960 ;
        RECT 64.090 15.130 64.260 15.930 ;
        RECT 64.640 15.830 64.810 15.930 ;
        RECT 64.580 15.790 64.900 15.830 ;
        RECT 64.570 15.600 64.900 15.790 ;
        RECT 64.580 15.570 64.900 15.600 ;
        RECT 62.320 15.090 62.640 15.130 ;
        RECT 64.020 15.090 64.340 15.130 ;
        RECT 62.320 14.900 62.650 15.090 ;
        RECT 64.010 14.900 64.340 15.090 ;
        RECT 62.320 14.870 62.640 14.900 ;
        RECT 64.020 14.870 64.340 14.900 ;
        RECT 62.400 13.790 62.570 14.870 ;
        RECT 64.090 13.790 64.260 14.870 ;
        RECT 62.310 13.750 62.630 13.790 ;
        RECT 64.030 13.750 64.350 13.790 ;
        RECT 62.310 13.560 62.640 13.750 ;
        RECT 64.020 13.560 64.350 13.750 ;
        RECT 62.310 13.530 62.630 13.560 ;
        RECT 64.030 13.530 64.350 13.560 ;
        RECT 61.760 13.020 62.080 13.060 ;
        RECT 61.760 12.830 62.090 13.020 ;
        RECT 61.760 12.800 62.080 12.830 ;
        RECT 61.850 11.690 62.020 12.800 ;
        RECT 61.760 11.650 62.080 11.690 ;
        RECT 61.760 11.460 62.090 11.650 ;
        RECT 61.760 11.430 62.080 11.460 ;
        RECT 61.210 10.970 61.530 11.010 ;
        RECT 61.210 10.780 61.540 10.970 ;
        RECT 61.210 10.750 61.530 10.780 ;
        RECT 61.300 10.600 61.470 10.750 ;
        RECT 61.850 10.600 62.020 11.430 ;
        RECT 62.400 11.020 62.570 13.530 ;
        RECT 64.090 11.020 64.260 13.530 ;
        RECT 64.640 13.060 64.810 15.570 ;
        RECT 65.190 15.140 65.360 15.930 ;
        RECT 65.740 15.840 65.910 15.930 ;
        RECT 65.680 15.800 66.000 15.840 ;
        RECT 65.670 15.610 66.000 15.800 ;
        RECT 65.680 15.580 66.000 15.610 ;
        RECT 65.130 15.100 65.450 15.140 ;
        RECT 65.120 14.910 65.450 15.100 ;
        RECT 65.130 14.880 65.450 14.910 ;
        RECT 65.190 13.790 65.360 14.880 ;
        RECT 65.130 13.750 65.450 13.790 ;
        RECT 65.120 13.560 65.450 13.750 ;
        RECT 65.130 13.530 65.450 13.560 ;
        RECT 64.580 13.020 64.900 13.060 ;
        RECT 64.570 12.830 64.900 13.020 ;
        RECT 64.580 12.800 64.900 12.830 ;
        RECT 64.640 11.690 64.810 12.800 ;
        RECT 64.580 11.650 64.900 11.690 ;
        RECT 64.570 11.460 64.900 11.650 ;
        RECT 64.580 11.430 64.900 11.460 ;
        RECT 62.310 10.980 62.630 11.020 ;
        RECT 64.030 10.980 64.350 11.020 ;
        RECT 62.310 10.790 62.640 10.980 ;
        RECT 64.020 10.790 64.350 10.980 ;
        RECT 62.310 10.760 62.630 10.790 ;
        RECT 64.030 10.760 64.350 10.790 ;
        RECT 62.400 10.600 62.570 10.760 ;
        RECT 64.090 10.600 64.260 10.760 ;
        RECT 64.640 10.600 64.810 11.430 ;
        RECT 65.190 11.010 65.360 13.530 ;
        RECT 65.740 13.060 65.910 15.580 ;
        RECT 66.290 15.160 66.460 15.930 ;
        RECT 66.840 15.840 67.010 15.930 ;
        RECT 66.770 15.800 67.090 15.840 ;
        RECT 66.760 15.610 67.090 15.800 ;
        RECT 66.770 15.580 67.090 15.610 ;
        RECT 66.220 15.120 66.540 15.160 ;
        RECT 66.210 14.930 66.540 15.120 ;
        RECT 66.220 14.900 66.540 14.930 ;
        RECT 66.290 13.790 66.460 14.900 ;
        RECT 66.220 13.750 66.540 13.790 ;
        RECT 66.210 13.560 66.540 13.750 ;
        RECT 66.220 13.530 66.540 13.560 ;
        RECT 65.680 13.020 66.000 13.060 ;
        RECT 65.670 12.830 66.000 13.020 ;
        RECT 65.680 12.800 66.000 12.830 ;
        RECT 65.740 11.690 65.910 12.800 ;
        RECT 65.680 11.650 66.000 11.690 ;
        RECT 65.670 11.460 66.000 11.650 ;
        RECT 65.680 11.430 66.000 11.460 ;
        RECT 65.130 10.970 65.450 11.010 ;
        RECT 65.120 10.780 65.450 10.970 ;
        RECT 65.130 10.750 65.450 10.780 ;
        RECT 65.190 10.600 65.360 10.750 ;
        RECT 65.740 10.600 65.910 11.430 ;
        RECT 66.290 11.010 66.460 13.530 ;
        RECT 66.840 13.060 67.010 15.580 ;
        RECT 69.840 15.120 70.010 15.860 ;
        RECT 70.390 15.820 70.560 15.860 ;
        RECT 70.320 15.780 70.640 15.820 ;
        RECT 70.310 15.590 70.640 15.780 ;
        RECT 70.320 15.560 70.640 15.590 ;
        RECT 69.760 15.080 70.080 15.120 ;
        RECT 69.750 14.890 70.080 15.080 ;
        RECT 69.760 14.860 70.080 14.890 ;
        RECT 69.840 13.780 70.010 14.860 ;
        RECT 69.770 13.740 70.090 13.780 ;
        RECT 69.760 13.550 70.090 13.740 ;
        RECT 69.770 13.520 70.090 13.550 ;
        RECT 66.780 13.020 67.100 13.060 ;
        RECT 66.770 12.830 67.100 13.020 ;
        RECT 66.780 12.800 67.100 12.830 ;
        RECT 66.840 11.690 67.010 12.800 ;
        RECT 66.780 11.650 67.100 11.690 ;
        RECT 66.770 11.460 67.100 11.650 ;
        RECT 66.780 11.430 67.100 11.460 ;
        RECT 66.220 10.970 66.540 11.010 ;
        RECT 66.210 10.780 66.540 10.970 ;
        RECT 66.220 10.750 66.540 10.780 ;
        RECT 66.290 10.600 66.460 10.750 ;
        RECT 66.840 10.610 67.010 11.430 ;
        RECT 67.270 11.220 67.780 11.300 ;
        RECT 67.260 10.970 67.780 11.220 ;
        RECT 69.840 11.010 70.010 13.520 ;
        RECT 70.390 13.050 70.560 15.560 ;
        RECT 70.940 15.130 71.110 15.860 ;
        RECT 71.490 15.830 71.660 15.860 ;
        RECT 71.420 15.790 71.740 15.830 ;
        RECT 71.410 15.600 71.740 15.790 ;
        RECT 71.420 15.570 71.740 15.600 ;
        RECT 70.870 15.090 71.190 15.130 ;
        RECT 70.860 14.900 71.190 15.090 ;
        RECT 70.870 14.870 71.190 14.900 ;
        RECT 70.940 13.780 71.110 14.870 ;
        RECT 70.870 13.740 71.190 13.780 ;
        RECT 70.860 13.550 71.190 13.740 ;
        RECT 70.870 13.520 71.190 13.550 ;
        RECT 70.320 13.010 70.640 13.050 ;
        RECT 70.310 12.820 70.640 13.010 ;
        RECT 70.320 12.790 70.640 12.820 ;
        RECT 70.390 11.680 70.560 12.790 ;
        RECT 70.320 11.640 70.640 11.680 ;
        RECT 70.310 11.450 70.640 11.640 ;
        RECT 70.320 11.420 70.640 11.450 ;
        RECT 69.770 10.970 70.090 11.010 ;
        RECT 67.260 10.290 67.770 10.970 ;
        RECT 69.760 10.780 70.090 10.970 ;
        RECT 69.770 10.750 70.090 10.780 ;
        RECT 69.840 10.680 70.010 10.750 ;
        RECT 70.390 10.680 70.560 11.420 ;
        RECT 70.940 11.000 71.110 13.520 ;
        RECT 71.490 13.050 71.660 15.570 ;
        RECT 72.040 15.150 72.210 15.860 ;
        RECT 72.590 15.830 72.760 15.860 ;
        RECT 72.510 15.790 72.830 15.830 ;
        RECT 72.500 15.600 72.830 15.790 ;
        RECT 72.510 15.570 72.830 15.600 ;
        RECT 71.960 15.110 72.280 15.150 ;
        RECT 71.950 14.920 72.280 15.110 ;
        RECT 71.960 14.890 72.280 14.920 ;
        RECT 72.040 13.780 72.210 14.890 ;
        RECT 71.960 13.740 72.280 13.780 ;
        RECT 71.950 13.550 72.280 13.740 ;
        RECT 71.960 13.520 72.280 13.550 ;
        RECT 71.420 13.010 71.740 13.050 ;
        RECT 71.410 12.820 71.740 13.010 ;
        RECT 71.420 12.790 71.740 12.820 ;
        RECT 71.490 11.680 71.660 12.790 ;
        RECT 71.420 11.640 71.740 11.680 ;
        RECT 71.410 11.450 71.740 11.640 ;
        RECT 71.420 11.420 71.740 11.450 ;
        RECT 70.870 10.960 71.190 11.000 ;
        RECT 70.860 10.770 71.190 10.960 ;
        RECT 70.870 10.740 71.190 10.770 ;
        RECT 70.940 10.680 71.110 10.740 ;
        RECT 71.490 10.680 71.660 11.420 ;
        RECT 72.040 11.000 72.210 13.520 ;
        RECT 72.590 13.050 72.760 15.570 ;
        RECT 72.520 13.010 72.840 13.050 ;
        RECT 72.510 12.820 72.840 13.010 ;
        RECT 72.520 12.790 72.840 12.820 ;
        RECT 72.590 11.680 72.760 12.790 ;
        RECT 72.520 11.640 72.840 11.680 ;
        RECT 72.510 11.450 72.840 11.640 ;
        RECT 73.300 11.480 73.470 12.700 ;
        RECT 72.520 11.420 72.840 11.450 ;
        RECT 71.960 10.960 72.280 11.000 ;
        RECT 71.950 10.770 72.280 10.960 ;
        RECT 71.960 10.740 72.280 10.770 ;
        RECT 72.040 10.680 72.210 10.740 ;
        RECT 72.590 10.680 72.760 11.420 ;
        RECT 73.010 11.030 73.520 11.290 ;
        RECT 73.000 10.960 73.520 11.030 ;
        RECT 73.000 10.280 73.510 10.960 ;
        RECT 18.240 8.840 18.560 8.870 ;
        RECT 18.230 8.650 18.560 8.840 ;
        RECT 18.240 8.610 18.560 8.650 ;
        RECT 18.320 8.580 18.490 8.610 ;
        RECT 104.390 7.990 104.620 8.000 ;
        RECT 104.370 7.820 109.030 7.990 ;
        RECT 104.390 7.810 104.620 7.820 ;
        RECT 109.930 7.340 110.120 7.350 ;
        RECT 105.590 7.300 109.390 7.310 ;
        RECT 109.900 7.300 110.160 7.340 ;
        RECT 105.590 7.140 110.160 7.300 ;
        RECT 109.160 7.130 110.160 7.140 ;
        RECT 109.160 6.670 109.390 7.130 ;
        RECT 109.900 7.020 110.160 7.130 ;
        RECT 109.930 6.670 110.120 6.680 ;
        RECT 15.600 6.140 15.770 6.300 ;
        RECT 15.540 6.110 15.860 6.140 ;
        RECT 15.530 5.920 15.860 6.110 ;
        RECT 15.540 5.880 15.860 5.920 ;
        RECT 15.600 3.370 15.770 5.880 ;
        RECT 16.150 5.470 16.320 6.300 ;
        RECT 16.700 6.150 16.870 6.300 ;
        RECT 16.640 6.120 16.960 6.150 ;
        RECT 16.630 5.930 16.960 6.120 ;
        RECT 16.640 5.890 16.960 5.930 ;
        RECT 16.090 5.440 16.410 5.470 ;
        RECT 16.080 5.250 16.410 5.440 ;
        RECT 16.090 5.210 16.410 5.250 ;
        RECT 16.150 4.100 16.320 5.210 ;
        RECT 16.090 4.070 16.410 4.100 ;
        RECT 16.080 3.880 16.410 4.070 ;
        RECT 16.090 3.840 16.410 3.880 ;
        RECT 15.540 3.340 15.860 3.370 ;
        RECT 15.530 3.150 15.860 3.340 ;
        RECT 15.540 3.110 15.860 3.150 ;
        RECT 15.600 2.030 15.770 3.110 ;
        RECT 15.530 2.000 15.850 2.030 ;
        RECT 15.520 1.810 15.850 2.000 ;
        RECT 15.530 1.770 15.850 1.810 ;
        RECT 15.060 0.940 15.230 1.700 ;
        RECT 15.600 0.970 15.770 1.770 ;
        RECT 16.150 1.330 16.320 3.840 ;
        RECT 16.700 3.370 16.870 5.890 ;
        RECT 17.250 5.470 17.420 6.300 ;
        RECT 17.800 6.150 17.970 6.300 ;
        RECT 17.730 6.120 18.050 6.150 ;
        RECT 17.720 5.930 18.050 6.120 ;
        RECT 17.730 5.890 18.050 5.930 ;
        RECT 17.190 5.440 17.510 5.470 ;
        RECT 17.180 5.250 17.510 5.440 ;
        RECT 17.190 5.210 17.510 5.250 ;
        RECT 17.250 4.100 17.420 5.210 ;
        RECT 17.190 4.070 17.510 4.100 ;
        RECT 17.180 3.880 17.510 4.070 ;
        RECT 17.190 3.840 17.510 3.880 ;
        RECT 16.640 3.340 16.960 3.370 ;
        RECT 16.630 3.150 16.960 3.340 ;
        RECT 16.640 3.110 16.960 3.150 ;
        RECT 16.700 2.020 16.870 3.110 ;
        RECT 16.640 1.990 16.960 2.020 ;
        RECT 16.630 1.800 16.960 1.990 ;
        RECT 16.640 1.760 16.960 1.800 ;
        RECT 16.090 1.300 16.410 1.330 ;
        RECT 16.080 1.110 16.410 1.300 ;
        RECT 16.090 1.070 16.410 1.110 ;
        RECT 16.150 0.970 16.320 1.070 ;
        RECT 16.700 0.970 16.870 1.760 ;
        RECT 17.250 1.320 17.420 3.840 ;
        RECT 17.800 3.370 17.970 5.890 ;
        RECT 18.350 5.470 18.520 6.290 ;
        RECT 18.770 5.930 19.280 6.610 ;
        RECT 109.160 6.460 110.170 6.670 ;
        RECT 104.390 6.380 104.620 6.390 ;
        RECT 104.370 6.210 108.850 6.380 ;
        RECT 104.390 6.200 104.620 6.210 ;
        RECT 18.770 5.680 19.290 5.930 ;
        RECT 109.160 5.700 109.390 6.460 ;
        RECT 109.900 6.350 110.160 6.460 ;
        RECT 18.780 5.600 19.290 5.680 ;
        RECT 105.610 5.530 109.390 5.700 ;
        RECT 18.290 5.440 18.610 5.470 ;
        RECT 18.280 5.250 18.610 5.440 ;
        RECT 18.290 5.210 18.610 5.250 ;
        RECT 18.350 4.100 18.520 5.210 ;
        RECT 20.350 4.970 22.740 5.340 ;
        RECT 18.290 4.070 18.610 4.100 ;
        RECT 18.280 3.880 18.610 4.070 ;
        RECT 18.290 3.840 18.610 3.880 ;
        RECT 17.730 3.340 18.050 3.370 ;
        RECT 17.720 3.150 18.050 3.340 ;
        RECT 17.730 3.110 18.050 3.150 ;
        RECT 17.800 2.000 17.970 3.110 ;
        RECT 17.730 1.970 18.050 2.000 ;
        RECT 17.720 1.780 18.050 1.970 ;
        RECT 17.730 1.740 18.050 1.780 ;
        RECT 17.190 1.290 17.510 1.320 ;
        RECT 17.180 1.100 17.510 1.290 ;
        RECT 17.190 1.060 17.510 1.100 ;
        RECT 17.250 0.970 17.420 1.060 ;
        RECT 17.800 0.970 17.970 1.740 ;
        RECT 18.350 1.320 18.520 3.840 ;
        RECT 20.400 1.710 22.740 4.970 ;
        RECT 104.390 4.780 104.620 4.790 ;
        RECT 104.370 4.610 108.870 4.780 ;
        RECT 104.390 4.600 104.620 4.610 ;
        RECT 105.610 4.600 105.940 4.610 ;
        RECT 106.570 4.600 106.900 4.610 ;
        RECT 107.530 4.600 107.860 4.610 ;
        RECT 108.490 4.600 108.820 4.610 ;
        RECT 109.160 4.090 109.390 5.530 ;
        RECT 109.880 5.340 110.310 5.360 ;
        RECT 109.860 5.170 110.310 5.340 ;
        RECT 109.880 5.150 110.310 5.170 ;
        RECT 105.610 3.920 109.390 4.090 ;
        RECT 105.670 3.640 106.100 3.660 ;
        RECT 105.650 3.470 106.100 3.640 ;
        RECT 105.670 3.450 106.100 3.470 ;
        RECT 104.390 3.160 104.620 3.170 ;
        RECT 104.370 2.990 108.870 3.160 ;
        RECT 104.390 2.980 104.620 2.990 ;
        RECT 109.160 2.490 109.390 3.920 ;
        RECT 109.880 3.730 110.310 3.750 ;
        RECT 109.860 3.560 110.310 3.730 ;
        RECT 109.880 3.540 110.310 3.560 ;
        RECT 105.620 2.480 109.390 2.490 ;
        RECT 105.610 2.320 109.390 2.480 ;
        RECT 105.610 2.310 105.940 2.320 ;
        RECT 107.530 2.310 107.860 2.320 ;
        RECT 108.490 2.310 108.820 2.320 ;
        RECT 106.670 2.000 107.100 2.020 ;
        RECT 106.670 1.830 107.120 2.000 ;
        RECT 106.670 1.810 107.100 1.830 ;
        RECT 20.400 1.700 22.730 1.710 ;
        RECT 104.390 1.560 104.620 1.570 ;
        RECT 104.370 1.390 108.820 1.560 ;
        RECT 104.390 1.380 104.620 1.390 ;
        RECT 105.610 1.380 105.940 1.390 ;
        RECT 106.570 1.380 106.900 1.390 ;
        RECT 107.530 1.380 107.860 1.390 ;
        RECT 108.490 1.380 108.820 1.390 ;
        RECT 18.280 1.290 18.600 1.320 ;
        RECT 18.270 1.100 18.600 1.290 ;
        RECT 18.280 1.060 18.600 1.100 ;
        RECT 18.350 0.970 18.520 1.060 ;
        RECT 109.160 0.870 109.390 2.320 ;
        RECT 109.870 2.120 110.300 2.140 ;
        RECT 109.850 1.950 110.300 2.120 ;
        RECT 109.870 1.930 110.300 1.950 ;
        RECT 105.600 0.700 109.390 0.870 ;
        RECT 107.580 0.420 108.010 0.440 ;
        RECT 107.560 0.250 108.010 0.420 ;
        RECT 107.580 0.230 108.010 0.250 ;
        RECT 104.390 -0.060 104.620 -0.050 ;
        RECT 104.370 -0.230 108.870 -0.060 ;
        RECT 104.390 -0.240 104.620 -0.230 ;
        RECT 105.610 -0.750 105.940 -0.740 ;
        RECT 106.570 -0.750 106.900 -0.740 ;
        RECT 107.530 -0.750 107.860 -0.740 ;
        RECT 108.490 -0.750 108.820 -0.740 ;
        RECT 109.160 -0.750 109.390 0.700 ;
        RECT 109.880 0.500 110.310 0.520 ;
        RECT 109.860 0.330 110.310 0.500 ;
        RECT 109.880 0.310 110.310 0.330 ;
        RECT 105.600 -0.920 109.390 -0.750 ;
        RECT 104.390 -1.660 104.620 -1.650 ;
        RECT 104.370 -1.670 108.790 -1.660 ;
        RECT 104.370 -1.830 108.820 -1.670 ;
        RECT 104.390 -1.840 104.620 -1.830 ;
        RECT 105.610 -1.840 105.940 -1.830 ;
        RECT 106.570 -1.840 106.900 -1.830 ;
        RECT 107.530 -1.840 107.860 -1.830 ;
        RECT 108.490 -1.840 108.820 -1.830 ;
        RECT 109.160 -2.340 109.390 -0.920 ;
        RECT 109.870 -1.110 110.300 -1.090 ;
        RECT 109.850 -1.280 110.300 -1.110 ;
        RECT 109.870 -1.300 110.300 -1.280 ;
        RECT 105.600 -2.510 109.400 -2.340 ;
        RECT 105.610 -2.520 105.940 -2.510 ;
        RECT 106.570 -2.520 106.900 -2.510 ;
        RECT 107.530 -2.520 107.860 -2.510 ;
        RECT 108.490 -2.520 108.820 -2.510 ;
        RECT 104.390 -3.290 104.620 -3.270 ;
        RECT 105.610 -3.290 105.940 -3.280 ;
        RECT 106.570 -3.290 106.900 -3.280 ;
        RECT 107.530 -3.290 107.860 -3.280 ;
        RECT 108.490 -3.290 108.820 -3.280 ;
        RECT 104.370 -3.460 108.830 -3.290 ;
        RECT 109.160 -3.950 109.390 -2.510 ;
        RECT 109.670 -3.150 109.880 -2.720 ;
        RECT 109.690 -3.170 109.860 -3.150 ;
        RECT 105.600 -4.120 109.390 -3.950 ;
        RECT 105.610 -4.130 105.940 -4.120 ;
        RECT 106.570 -4.130 106.900 -4.120 ;
        RECT 107.530 -4.130 107.860 -4.120 ;
        RECT 108.490 -4.130 108.820 -4.120 ;
        RECT 109.870 -4.310 110.300 -4.290 ;
        RECT 109.850 -4.480 110.300 -4.310 ;
        RECT 109.870 -4.500 110.300 -4.480 ;
        RECT 110.580 -5.290 110.950 9.580 ;
        RECT 110.580 -5.540 110.960 -5.290 ;
        RECT 106.630 -6.020 107.060 -6.000 ;
        RECT 107.570 -6.020 108.000 -6.000 ;
        RECT 109.830 -6.020 110.260 -6.000 ;
        RECT 106.610 -6.190 107.060 -6.020 ;
        RECT 107.550 -6.190 108.000 -6.020 ;
        RECT 108.520 -6.040 108.950 -6.020 ;
        RECT 106.630 -6.210 107.060 -6.190 ;
        RECT 107.570 -6.210 108.000 -6.190 ;
        RECT 108.500 -6.210 108.950 -6.040 ;
        RECT 109.810 -6.190 110.260 -6.020 ;
        RECT 109.830 -6.210 110.260 -6.190 ;
        RECT 108.520 -6.230 108.950 -6.210 ;
      LAYER mcon ;
        RECT 6.670 61.070 6.840 61.240 ;
        RECT 9.540 61.280 9.710 61.450 ;
        RECT 8.080 61.070 8.250 61.240 ;
        RECT 24.880 61.100 25.050 61.270 ;
        RECT 9.540 60.490 9.710 60.660 ;
        RECT 24.880 60.410 25.050 60.580 ;
        RECT 30.740 61.010 30.910 61.180 ;
        RECT 30.740 60.560 30.910 60.730 ;
        RECT 35.440 60.960 35.610 61.130 ;
        RECT 35.440 60.510 35.610 60.680 ;
        RECT 6.670 60.220 6.840 60.390 ;
        RECT 7.390 60.210 7.560 60.380 ;
        RECT 8.080 60.220 8.250 60.390 ;
        RECT 6.850 59.810 7.020 59.980 ;
        RECT 7.910 59.810 8.080 59.980 ;
        RECT 6.670 59.400 6.840 59.570 ;
        RECT 7.390 59.370 7.560 59.540 ;
        RECT 8.080 59.400 8.250 59.570 ;
        RECT 22.780 59.470 22.950 59.640 ;
        RECT 24.140 59.550 24.310 59.720 ;
        RECT 24.830 59.540 25.000 59.710 ;
        RECT 9.540 59.060 9.710 59.230 ;
        RECT 6.670 58.560 6.840 58.730 ;
        RECT 8.080 58.560 8.250 58.730 ;
        RECT 8.810 58.300 8.980 58.470 ;
        RECT 8.800 57.780 8.970 57.950 ;
        RECT 9.550 57.660 9.720 57.830 ;
        RECT 6.670 57.440 6.840 57.610 ;
        RECT 8.080 57.440 8.250 57.610 ;
        RECT 7.370 56.570 7.540 56.740 ;
        RECT 8.800 56.590 8.970 56.760 ;
        RECT 11.560 56.240 11.730 56.410 ;
        RECT 6.580 55.990 6.750 56.160 ;
        RECT 7.510 55.990 7.680 56.160 ;
        RECT 8.210 55.990 8.380 56.160 ;
        RECT 8.950 55.990 9.120 56.160 ;
        RECT 9.660 55.980 9.830 56.150 ;
        RECT 24.880 58.300 25.050 58.470 ;
        RECT 24.880 57.610 25.050 57.780 ;
        RECT 30.740 58.020 30.910 58.190 ;
        RECT 30.740 57.570 30.910 57.740 ;
        RECT 30.740 57.010 30.910 57.180 ;
        RECT 24.880 56.750 25.050 56.920 ;
        RECT 30.740 56.560 30.910 56.730 ;
        RECT 24.880 56.060 25.050 56.230 ;
        RECT 34.660 57.500 34.830 57.670 ;
        RECT 22.060 55.810 22.230 55.980 ;
        RECT 31.920 55.830 32.090 56.000 ;
        RECT 22.070 51.450 22.500 52.190 ;
        RECT 43.170 50.030 43.380 50.240 ;
        RECT 46.910 50.050 47.080 50.220 ;
        RECT 41.700 49.660 41.870 49.830 ;
        RECT 47.950 50.090 48.120 50.260 ;
        RECT 48.990 49.750 49.160 49.920 ;
        RECT 48.990 49.390 49.160 49.560 ;
        RECT 43.170 48.280 43.380 48.490 ;
        RECT 46.910 48.300 47.080 48.470 ;
        RECT 41.700 47.910 41.870 48.080 ;
        RECT 47.950 48.340 48.120 48.510 ;
        RECT 70.360 48.290 70.620 49.110 ;
        RECT 82.310 48.320 82.630 49.110 ;
        RECT 48.990 48.000 49.160 48.170 ;
        RECT 48.990 47.640 49.160 47.810 ;
        RECT 19.950 46.670 20.120 46.840 ;
        RECT 21.040 46.680 21.210 46.850 ;
        RECT 43.170 46.530 43.380 46.740 ;
        RECT 46.910 46.550 47.080 46.720 ;
        RECT 19.520 46.170 19.690 46.340 ;
        RECT 21.890 46.110 22.060 46.280 ;
        RECT 41.700 46.160 41.870 46.330 ;
        RECT 19.960 45.680 20.130 45.850 ;
        RECT 21.050 45.690 21.220 45.860 ;
        RECT 47.950 46.590 48.120 46.760 ;
        RECT 80.470 46.540 80.640 46.710 ;
        RECT 48.990 46.250 49.160 46.420 ;
        RECT 58.420 46.230 58.600 46.400 ;
        RECT 58.850 46.210 59.020 46.380 ;
        RECT 48.990 45.890 49.160 46.060 ;
        RECT 56.610 45.930 56.780 46.100 ;
        RECT 19.500 45.250 19.670 45.420 ;
        RECT 56.960 45.090 57.140 45.280 ;
        RECT 19.960 44.690 20.130 44.860 ;
        RECT 21.050 44.700 21.220 44.870 ;
        RECT 43.170 44.780 43.380 44.990 ;
        RECT 46.910 44.800 47.080 44.970 ;
        RECT 19.480 44.260 19.650 44.430 ;
        RECT 41.700 44.410 41.870 44.580 ;
        RECT 47.950 44.840 48.120 45.010 ;
        RECT 48.990 44.500 49.160 44.670 ;
        RECT 48.990 44.140 49.160 44.310 ;
        RECT 59.320 45.650 59.490 45.820 ;
        RECT 78.570 45.930 78.740 46.100 ;
        RECT 61.560 45.350 61.730 45.520 ;
        RECT 71.730 45.350 71.900 45.520 ;
        RECT 61.560 44.900 61.730 45.070 ;
        RECT 58.040 44.530 58.210 44.700 ;
        RECT 67.010 44.750 67.280 45.020 ;
        RECT 68.070 44.750 68.340 45.020 ;
        RECT 71.730 44.900 71.900 45.070 ;
        RECT 76.900 45.100 77.070 45.270 ;
        RECT 58.850 44.220 59.020 44.390 ;
        RECT 19.770 43.760 19.940 43.930 ;
        RECT 21.070 43.660 21.240 43.830 ;
        RECT 19.770 42.770 19.940 42.940 ;
        RECT 21.070 42.670 21.240 42.840 ;
        RECT 41.700 42.710 41.870 42.880 ;
        RECT 50.150 43.230 50.320 43.400 ;
        RECT 48.990 42.980 49.160 43.150 ;
        RECT 50.990 43.110 51.160 43.280 ;
        RECT 51.740 43.110 51.910 43.280 ;
        RECT 21.480 42.190 21.650 42.360 ;
        RECT 43.170 42.300 43.380 42.510 ;
        RECT 46.910 42.320 47.080 42.490 ;
        RECT 48.990 42.620 49.160 42.790 ;
        RECT 47.950 42.280 48.120 42.450 ;
        RECT 54.720 42.780 54.890 42.950 ;
        RECT 50.430 42.480 50.600 42.650 ;
        RECT 55.120 43.230 55.290 43.400 ;
        RECT 81.440 46.290 81.610 46.460 ;
        RECT 82.420 45.970 82.590 46.140 ;
        RECT 83.690 46.310 83.860 46.480 ;
        RECT 80.620 45.710 80.790 45.880 ;
        RECT 78.210 45.090 78.390 45.280 ;
        RECT 79.500 45.190 79.670 45.360 ;
        RECT 64.690 43.640 64.860 43.810 ;
        RECT 70.490 43.640 70.660 43.810 ;
        RECT 55.120 42.870 55.290 43.040 ;
        RECT 56.960 42.290 57.140 42.480 ;
        RECT 19.770 41.780 19.940 41.950 ;
        RECT 21.070 41.680 21.240 41.850 ;
        RECT 41.700 40.960 41.870 41.130 ;
        RECT 48.990 41.230 49.160 41.400 ;
        RECT 50.430 41.420 50.600 41.590 ;
        RECT 59.320 43.330 59.490 43.500 ;
        RECT 58.860 43.150 59.030 43.320 ;
        RECT 58.030 42.840 58.200 43.010 ;
        RECT 67.010 43.020 67.280 43.290 ;
        RECT 68.070 43.020 68.340 43.290 ;
        RECT 61.560 42.400 61.730 42.570 ;
        RECT 61.560 41.950 61.730 42.120 ;
        RECT 71.730 42.400 71.900 42.570 ;
        RECT 76.900 42.340 77.070 42.510 ;
        RECT 71.730 41.950 71.900 42.120 ;
        RECT 59.310 41.750 59.480 41.920 ;
        RECT 43.170 40.550 43.380 40.760 ;
        RECT 46.910 40.570 47.080 40.740 ;
        RECT 54.720 41.120 54.890 41.290 ;
        RECT 48.990 40.870 49.160 41.040 ;
        RECT 47.950 40.530 48.120 40.700 ;
        RECT 50.990 40.790 51.160 40.960 ;
        RECT 51.740 40.790 51.910 40.960 ;
        RECT 53.740 40.800 53.910 40.970 ;
        RECT 55.120 41.390 55.290 41.560 ;
        RECT 56.610 41.470 56.780 41.640 ;
        RECT 55.120 41.030 55.290 41.200 ;
        RECT 78.210 42.290 78.390 42.480 ;
        RECT 78.570 41.470 78.740 41.640 ;
        RECT 58.420 41.170 58.600 41.340 ;
        RECT 58.880 41.240 59.050 41.410 ;
        RECT 81.390 45.640 81.560 45.810 ;
        RECT 81.390 44.800 81.560 44.970 ;
        RECT 83.080 45.000 83.250 45.170 ;
        RECT 82.420 44.470 82.590 44.640 ;
        RECT 81.440 44.150 81.610 44.320 ;
        RECT 80.230 43.910 80.400 44.080 ;
        RECT 83.740 44.090 83.910 44.260 ;
        RECT 109.150 43.840 109.320 44.010 ;
        RECT 110.110 43.700 110.280 43.870 ;
        RECT 110.720 43.840 110.890 44.010 ;
        RECT 111.240 43.710 111.410 43.880 ;
        RECT 80.660 43.110 80.830 43.280 ;
        RECT 81.440 43.290 81.610 43.460 ;
        RECT 83.730 43.370 83.900 43.540 ;
        RECT 82.420 42.970 82.590 43.140 ;
        RECT 81.390 42.640 81.560 42.810 ;
        RECT 107.700 43.060 107.870 43.230 ;
        RECT 108.200 43.090 108.370 43.260 ;
        RECT 111.700 43.090 111.870 43.260 ;
        RECT 83.080 42.410 83.250 42.580 ;
        RECT 81.390 41.800 81.560 41.970 ;
        RECT 108.200 42.010 108.370 42.180 ;
        RECT 111.700 42.010 111.870 42.180 ;
        RECT 82.420 41.470 82.590 41.640 ;
        RECT 81.440 41.150 81.610 41.320 ;
        RECT 83.650 41.120 83.820 41.290 ;
        RECT 109.150 41.260 109.320 41.430 ;
        RECT 110.110 41.400 110.280 41.570 ;
        RECT 110.720 41.260 110.890 41.430 ;
        RECT 111.240 41.390 111.410 41.560 ;
        RECT 50.150 40.030 50.320 40.200 ;
        RECT 41.700 39.210 41.870 39.380 ;
        RECT 50.990 39.910 51.160 40.080 ;
        RECT 51.740 39.910 51.910 40.080 ;
        RECT 48.990 39.480 49.160 39.650 ;
        RECT 43.170 38.800 43.380 39.010 ;
        RECT 46.910 38.820 47.080 38.990 ;
        RECT 48.990 39.120 49.160 39.290 ;
        RECT 54.720 39.580 54.890 39.750 ;
        RECT 50.430 39.280 50.600 39.450 ;
        RECT 55.120 40.030 55.290 40.200 ;
        RECT 58.430 40.200 58.610 40.370 ;
        RECT 55.120 39.670 55.290 39.840 ;
        RECT 56.620 39.900 56.790 40.070 ;
        RECT 56.970 39.060 57.150 39.250 ;
        RECT 47.950 38.780 48.120 38.950 ;
        RECT 50.430 38.220 50.600 38.390 ;
        RECT 41.700 37.460 41.870 37.630 ;
        RECT 54.720 37.920 54.890 38.090 ;
        RECT 48.990 37.730 49.160 37.900 ;
        RECT 43.170 37.050 43.380 37.260 ;
        RECT 46.910 37.070 47.080 37.240 ;
        RECT 48.990 37.370 49.160 37.540 ;
        RECT 50.990 37.590 51.160 37.760 ;
        RECT 51.740 37.590 51.910 37.760 ;
        RECT 53.740 37.600 53.910 37.770 ;
        RECT 55.120 38.190 55.290 38.360 ;
        RECT 80.470 40.510 80.640 40.680 ;
        RECT 78.570 39.900 78.740 40.070 ;
        RECT 63.460 39.320 63.630 39.490 ;
        RECT 65.550 39.480 65.720 39.650 ;
        RECT 58.290 39.070 58.460 39.240 ;
        RECT 71.730 39.320 71.900 39.490 ;
        RECT 63.460 38.870 63.630 39.040 ;
        RECT 67.020 38.720 67.290 38.990 ;
        RECT 68.070 38.720 68.340 38.990 ;
        RECT 71.730 38.870 71.900 39.040 ;
        RECT 76.900 39.070 77.070 39.240 ;
        RECT 55.120 37.830 55.290 38.000 ;
        RECT 64.700 37.970 64.870 38.140 ;
        RECT 64.700 37.610 64.870 37.780 ;
        RECT 47.950 37.030 48.120 37.200 ;
        RECT 56.970 36.260 57.150 36.450 ;
        RECT 64.710 37.250 64.880 37.420 ;
        RECT 70.490 37.970 70.660 38.140 ;
        RECT 81.440 40.260 81.610 40.430 ;
        RECT 82.420 39.940 82.590 40.110 ;
        RECT 83.690 40.280 83.860 40.450 ;
        RECT 109.150 40.640 109.320 40.810 ;
        RECT 110.110 40.500 110.280 40.670 ;
        RECT 110.720 40.640 110.890 40.810 ;
        RECT 111.240 40.510 111.410 40.680 ;
        RECT 80.620 39.680 80.790 39.850 ;
        RECT 78.210 39.060 78.390 39.250 ;
        RECT 79.500 39.160 79.670 39.330 ;
        RECT 70.490 37.610 70.660 37.780 ;
        RECT 67.020 36.990 67.290 37.260 ;
        RECT 68.070 36.990 68.340 37.260 ;
        RECT 70.490 37.250 70.660 37.420 ;
        RECT 58.290 36.310 58.460 36.480 ;
        RECT 63.460 36.370 63.630 36.540 ;
        RECT 63.460 35.920 63.630 36.090 ;
        RECT 71.730 36.370 71.900 36.540 ;
        RECT 76.900 36.310 77.070 36.480 ;
        RECT 65.580 35.790 65.750 35.960 ;
        RECT 71.730 35.920 71.900 36.090 ;
        RECT 78.210 36.260 78.390 36.450 ;
        RECT 56.620 35.440 56.790 35.610 ;
        RECT 58.430 35.140 58.610 35.310 ;
        RECT 78.570 35.440 78.740 35.610 ;
        RECT 81.390 39.610 81.560 39.780 ;
        RECT 107.700 39.860 107.870 40.030 ;
        RECT 108.200 39.890 108.370 40.060 ;
        RECT 111.700 39.890 111.870 40.060 ;
        RECT 81.390 38.770 81.560 38.940 ;
        RECT 83.080 38.970 83.250 39.140 ;
        RECT 82.420 38.440 82.590 38.610 ;
        RECT 108.200 38.810 108.370 38.980 ;
        RECT 111.700 38.810 111.870 38.980 ;
        RECT 81.440 38.120 81.610 38.290 ;
        RECT 80.230 37.880 80.400 38.050 ;
        RECT 83.740 38.060 83.910 38.230 ;
        RECT 109.150 38.060 109.320 38.230 ;
        RECT 110.110 38.200 110.280 38.370 ;
        RECT 110.720 38.060 110.890 38.230 ;
        RECT 111.240 38.190 111.410 38.360 ;
        RECT 80.660 37.080 80.830 37.250 ;
        RECT 81.440 37.260 81.610 37.430 ;
        RECT 83.730 37.340 83.900 37.510 ;
        RECT 82.420 36.940 82.590 37.110 ;
        RECT 81.390 36.610 81.560 36.780 ;
        RECT 83.080 36.380 83.250 36.550 ;
        RECT 81.390 35.770 81.560 35.940 ;
        RECT 82.420 35.440 82.590 35.610 ;
        RECT 81.440 35.120 81.610 35.290 ;
        RECT 83.650 35.090 83.820 35.260 ;
        RECT 41.700 32.580 41.870 32.750 ;
        RECT 48.990 32.850 49.160 33.020 ;
        RECT 43.170 32.170 43.380 32.380 ;
        RECT 46.910 32.190 47.080 32.360 ;
        RECT 48.990 32.490 49.160 32.660 ;
        RECT 50.130 32.760 50.300 32.930 ;
        RECT 50.970 32.640 51.140 32.810 ;
        RECT 51.720 32.640 51.890 32.810 ;
        RECT 47.950 32.150 48.120 32.320 ;
        RECT 54.700 32.310 54.870 32.480 ;
        RECT 50.410 32.010 50.580 32.180 ;
        RECT 55.100 32.760 55.270 32.930 ;
        RECT 55.100 32.400 55.270 32.570 ;
        RECT 59.840 32.580 60.010 32.750 ;
        RECT 75.330 32.580 75.500 32.750 ;
        RECT 58.030 32.320 58.200 32.490 ;
        RECT 58.760 32.290 58.930 32.460 ;
        RECT 76.410 32.290 76.580 32.460 ;
        RECT 59.840 32.030 60.010 32.200 ;
        RECT 75.330 32.030 75.500 32.200 ;
        RECT 77.140 32.320 77.310 32.490 ;
        RECT 60.750 31.630 60.920 31.800 ;
        RECT 41.700 30.830 41.870 31.000 ;
        RECT 48.990 31.100 49.160 31.270 ;
        RECT 43.170 30.420 43.380 30.630 ;
        RECT 46.910 30.440 47.080 30.610 ;
        RECT 48.990 30.740 49.160 30.910 ;
        RECT 50.410 30.950 50.580 31.120 ;
        RECT 54.700 30.650 54.870 30.820 ;
        RECT 47.950 30.400 48.120 30.570 ;
        RECT 50.970 30.320 51.140 30.490 ;
        RECT 51.720 30.320 51.890 30.490 ;
        RECT 53.720 30.330 53.890 30.500 ;
        RECT 55.100 30.920 55.270 31.090 ;
        RECT 58.030 30.760 58.200 30.930 ;
        RECT 64.690 31.640 64.860 31.810 ;
        RECT 70.480 31.640 70.650 31.810 ;
        RECT 74.420 31.630 74.590 31.800 ;
        RECT 59.840 31.050 60.010 31.220 ;
        RECT 75.330 31.050 75.500 31.220 ;
        RECT 58.760 30.790 58.930 30.960 ;
        RECT 76.410 30.790 76.580 30.960 ;
        RECT 77.140 30.760 77.310 30.930 ;
        RECT 55.100 30.560 55.270 30.730 ;
        RECT 59.840 30.500 60.010 30.670 ;
        RECT 60.750 30.040 60.920 30.210 ;
        RECT 64.680 30.180 64.850 30.350 ;
        RECT 75.330 30.500 75.500 30.670 ;
        RECT 41.700 29.080 41.870 29.250 ;
        RECT 50.130 29.560 50.300 29.730 ;
        RECT 48.990 29.350 49.160 29.520 ;
        RECT 43.170 28.670 43.380 28.880 ;
        RECT 46.910 28.690 47.080 28.860 ;
        RECT 50.970 29.440 51.140 29.610 ;
        RECT 51.720 29.440 51.890 29.610 ;
        RECT 48.990 28.990 49.160 29.160 ;
        RECT 47.950 28.650 48.120 28.820 ;
        RECT 54.700 29.110 54.870 29.280 ;
        RECT 50.410 28.810 50.580 28.980 ;
        RECT 55.100 29.560 55.270 29.730 ;
        RECT 60.750 29.680 60.920 29.850 ;
        RECT 62.960 29.790 63.230 30.060 ;
        RECT 64.680 29.820 64.850 29.990 ;
        RECT 55.100 29.200 55.270 29.370 ;
        RECT 59.840 29.340 60.010 29.510 ;
        RECT 66.990 29.860 67.260 30.130 ;
        RECT 68.080 29.860 68.350 30.130 ;
        RECT 70.490 30.180 70.660 30.350 ;
        RECT 70.490 29.820 70.660 29.990 ;
        RECT 72.110 29.790 72.380 30.060 ;
        RECT 74.420 30.040 74.590 30.210 ;
        RECT 76.780 29.920 76.960 30.090 ;
        RECT 74.420 29.680 74.590 29.850 ;
        RECT 75.330 29.340 75.500 29.510 ;
        RECT 58.030 29.080 58.200 29.250 ;
        RECT 58.760 29.050 58.930 29.220 ;
        RECT 76.410 29.050 76.580 29.220 ;
        RECT 59.840 28.790 60.010 28.960 ;
        RECT 75.330 28.790 75.500 28.960 ;
        RECT 77.140 29.080 77.310 29.250 ;
        RECT 41.700 27.330 41.870 27.500 ;
        RECT 48.990 27.600 49.160 27.770 ;
        RECT 50.410 27.750 50.580 27.920 ;
        RECT 43.170 26.920 43.380 27.130 ;
        RECT 46.910 26.940 47.080 27.110 ;
        RECT 54.700 27.450 54.870 27.620 ;
        RECT 48.990 27.240 49.160 27.410 ;
        RECT 47.950 26.900 48.120 27.070 ;
        RECT 50.970 27.120 51.140 27.290 ;
        RECT 51.720 27.120 51.890 27.290 ;
        RECT 53.720 27.130 53.890 27.300 ;
        RECT 55.100 27.720 55.270 27.890 ;
        RECT 55.100 27.360 55.270 27.530 ;
        RECT 58.030 27.530 58.200 27.700 ;
        RECT 59.840 27.820 60.010 27.990 ;
        RECT 75.330 27.820 75.500 27.990 ;
        RECT 58.760 27.560 58.930 27.730 ;
        RECT 76.410 27.560 76.580 27.730 ;
        RECT 77.140 27.530 77.310 27.700 ;
        RECT 59.840 27.270 60.010 27.440 ;
        RECT 75.330 27.270 75.500 27.440 ;
        RECT 18.890 24.100 19.060 24.270 ;
        RECT 19.540 24.100 19.710 24.270 ;
        RECT 17.670 23.660 17.840 23.830 ;
        RECT 18.370 23.660 18.540 23.830 ;
        RECT 17.220 22.000 17.390 22.170 ;
        RECT 41.660 23.520 41.830 23.690 ;
        RECT 48.950 23.790 49.120 23.960 ;
        RECT 20.050 23.280 20.220 23.450 ;
        RECT 43.130 23.110 43.340 23.320 ;
        RECT 46.870 23.130 47.040 23.300 ;
        RECT 48.950 23.430 49.120 23.600 ;
        RECT 50.160 23.490 50.330 23.660 ;
        RECT 47.910 23.090 48.080 23.260 ;
        RECT 51.000 23.370 51.170 23.540 ;
        RECT 51.750 23.370 51.920 23.540 ;
        RECT 54.730 23.040 54.900 23.210 ;
        RECT 50.440 22.740 50.610 22.910 ;
        RECT 55.130 23.490 55.300 23.660 ;
        RECT 55.130 23.130 55.300 23.300 ;
        RECT 59.870 23.250 60.040 23.420 ;
        RECT 58.060 22.990 58.230 23.160 ;
        RECT 58.790 22.960 58.960 23.130 ;
        RECT 68.550 22.960 68.720 23.130 ;
        RECT 59.870 22.700 60.040 22.870 ;
        RECT 20.220 21.800 20.390 21.970 ;
        RECT 41.660 21.770 41.830 21.940 ;
        RECT 60.910 22.240 61.080 22.410 ;
        RECT 48.950 22.040 49.120 22.210 ;
        RECT 17.700 19.780 17.870 19.950 ;
        RECT 18.390 19.770 18.560 19.940 ;
        RECT 18.870 19.000 19.040 19.170 ;
        RECT 20.230 21.260 20.400 21.430 ;
        RECT 43.130 21.360 43.340 21.570 ;
        RECT 46.870 21.380 47.040 21.550 ;
        RECT 48.950 21.680 49.120 21.850 ;
        RECT 47.910 21.340 48.080 21.510 ;
        RECT 50.440 21.680 50.610 21.850 ;
        RECT 54.730 21.380 54.900 21.550 ;
        RECT 51.000 21.050 51.170 21.220 ;
        RECT 51.750 21.050 51.920 21.220 ;
        RECT 53.750 21.060 53.920 21.230 ;
        RECT 55.130 21.650 55.300 21.820 ;
        RECT 55.130 21.290 55.300 21.460 ;
        RECT 58.060 21.450 58.230 21.620 ;
        RECT 59.870 21.740 60.040 21.910 ;
        RECT 64.930 22.270 65.100 22.440 ;
        RECT 68.700 22.280 68.870 22.450 ;
        RECT 70.850 22.400 71.020 22.570 ;
        RECT 69.590 21.830 69.760 22.000 ;
        RECT 58.790 21.480 58.960 21.650 ;
        RECT 59.870 21.190 60.040 21.360 ;
        RECT 68.700 21.380 68.870 21.550 ;
        RECT 60.900 21.040 61.070 21.210 ;
        RECT 20.040 20.300 20.210 20.470 ;
        RECT 41.660 20.020 41.830 20.190 ;
        RECT 64.920 20.980 65.090 21.150 ;
        RECT 70.850 21.260 71.020 21.430 ;
        RECT 48.950 20.290 49.120 20.460 ;
        RECT 43.130 19.610 43.340 19.820 ;
        RECT 46.870 19.630 47.040 19.800 ;
        RECT 48.950 19.930 49.120 20.100 ;
        RECT 50.160 20.290 50.330 20.460 ;
        RECT 51.000 20.170 51.170 20.340 ;
        RECT 51.750 20.170 51.920 20.340 ;
        RECT 47.910 19.590 48.080 19.760 ;
        RECT 54.730 19.840 54.900 20.010 ;
        RECT 50.440 19.540 50.610 19.710 ;
        RECT 55.130 20.290 55.300 20.460 ;
        RECT 60.900 20.380 61.070 20.550 ;
        RECT 55.130 19.930 55.300 20.100 ;
        RECT 59.870 20.010 60.040 20.180 ;
        RECT 62.990 20.420 63.260 20.690 ;
        RECT 64.920 20.340 65.090 20.510 ;
        RECT 67.020 20.490 67.290 20.760 ;
        RECT 68.550 20.700 68.720 20.870 ;
        RECT 68.550 20.190 68.720 20.360 ;
        RECT 58.060 19.750 58.230 19.920 ;
        RECT 58.790 19.720 58.960 19.890 ;
        RECT 59.870 19.460 60.040 19.630 ;
        RECT 68.700 19.510 68.870 19.680 ;
        RECT 70.850 19.630 71.020 19.800 ;
        RECT 19.580 18.940 19.750 19.110 ;
        RECT 69.590 19.060 69.760 19.230 ;
        RECT 41.660 18.270 41.830 18.440 ;
        RECT 48.950 18.540 49.120 18.710 ;
        RECT 43.130 17.860 43.340 18.070 ;
        RECT 46.870 17.880 47.040 18.050 ;
        RECT 50.440 18.480 50.610 18.650 ;
        RECT 48.950 18.180 49.120 18.350 ;
        RECT 54.730 18.180 54.900 18.350 ;
        RECT 47.910 17.840 48.080 18.010 ;
        RECT 51.000 17.850 51.170 18.020 ;
        RECT 51.750 17.850 51.920 18.020 ;
        RECT 53.750 17.860 53.920 18.030 ;
        RECT 55.130 18.450 55.300 18.620 ;
        RECT 57.110 18.550 57.280 18.720 ;
        RECT 55.130 18.090 55.300 18.260 ;
        RECT 58.060 18.200 58.230 18.370 ;
        RECT 59.870 18.490 60.040 18.660 ;
        RECT 68.700 18.610 68.870 18.780 ;
        RECT 58.790 18.230 58.960 18.400 ;
        RECT 70.850 18.490 71.020 18.660 ;
        RECT 59.870 17.940 60.040 18.110 ;
        RECT 68.550 17.930 68.720 18.100 ;
        RECT 57.160 17.590 57.330 17.760 ;
        RECT 49.820 15.590 49.990 15.760 ;
        RECT 18.900 13.920 19.070 14.090 ;
        RECT 15.590 13.480 15.760 13.650 ;
        RECT 16.690 13.490 16.860 13.660 ;
        RECT 16.140 12.810 16.310 12.980 ;
        RECT 16.140 11.440 16.310 11.610 ;
        RECT 15.590 10.710 15.760 10.880 ;
        RECT 15.580 9.370 15.750 9.540 ;
        RECT 17.780 13.490 17.950 13.660 ;
        RECT 17.240 12.810 17.410 12.980 ;
        RECT 17.240 11.440 17.410 11.610 ;
        RECT 16.690 10.710 16.860 10.880 ;
        RECT 16.690 9.360 16.860 9.530 ;
        RECT 16.140 8.670 16.310 8.840 ;
        RECT 26.220 13.740 26.390 14.080 ;
        RECT 26.590 13.740 26.760 14.080 ;
        RECT 18.910 13.450 19.080 13.620 ;
        RECT 18.340 12.810 18.510 12.980 ;
        RECT 19.030 12.790 19.200 12.960 ;
        RECT 50.910 15.590 51.080 15.760 ;
        RECT 50.370 14.910 50.540 15.080 ;
        RECT 50.370 13.540 50.540 13.710 ;
        RECT 49.810 12.810 49.980 12.980 ;
        RECT 19.030 12.100 19.200 12.270 ;
        RECT 18.340 11.440 18.510 11.610 ;
        RECT 49.810 11.440 49.980 11.610 ;
        RECT 17.780 10.710 17.950 10.880 ;
        RECT 17.780 9.340 17.950 9.510 ;
        RECT 17.240 8.660 17.410 8.830 ;
        RECT 49.240 10.800 49.410 10.970 ;
        RECT 52.010 15.580 52.180 15.750 ;
        RECT 51.460 14.890 51.630 15.060 ;
        RECT 51.460 13.540 51.630 13.710 ;
        RECT 50.910 12.810 51.080 12.980 ;
        RECT 50.910 11.440 51.080 11.610 ;
        RECT 50.370 10.760 50.540 10.930 ;
        RECT 53.130 15.760 53.300 15.930 ;
        RECT 53.130 15.400 53.300 15.570 ;
        RECT 53.740 15.760 53.910 15.930 ;
        RECT 53.740 15.400 53.910 15.570 ;
        RECT 54.860 15.580 55.030 15.750 ;
        RECT 52.570 14.880 52.740 15.050 ;
        RECT 54.300 14.880 54.470 15.050 ;
        RECT 52.560 13.540 52.730 13.710 ;
        RECT 54.310 13.540 54.480 13.710 ;
        RECT 52.010 12.810 52.180 12.980 ;
        RECT 52.010 11.440 52.180 11.610 ;
        RECT 51.460 10.760 51.630 10.930 ;
        RECT 55.960 15.590 56.130 15.760 ;
        RECT 55.410 14.890 55.580 15.060 ;
        RECT 55.410 13.540 55.580 13.710 ;
        RECT 54.860 12.810 55.030 12.980 ;
        RECT 54.860 11.440 55.030 11.610 ;
        RECT 52.560 10.770 52.730 10.940 ;
        RECT 54.310 10.770 54.480 10.940 ;
        RECT 57.050 15.590 57.220 15.760 ;
        RECT 59.630 15.620 59.800 15.790 ;
        RECT 56.500 14.910 56.670 15.080 ;
        RECT 56.500 13.540 56.670 13.710 ;
        RECT 55.960 12.810 56.130 12.980 ;
        RECT 55.960 11.440 56.130 11.610 ;
        RECT 55.410 10.760 55.580 10.930 ;
        RECT 60.720 15.620 60.890 15.790 ;
        RECT 60.180 14.940 60.350 15.110 ;
        RECT 60.180 13.570 60.350 13.740 ;
        RECT 57.060 12.810 57.230 12.980 ;
        RECT 59.620 12.840 59.790 13.010 ;
        RECT 57.060 11.440 57.230 11.610 ;
        RECT 59.620 11.470 59.790 11.640 ;
        RECT 56.500 10.760 56.670 10.930 ;
        RECT 57.630 10.800 57.800 10.970 ;
        RECT 49.250 10.330 49.420 10.500 ;
        RECT 57.620 10.330 57.790 10.500 ;
        RECT 59.050 10.830 59.220 11.000 ;
        RECT 61.820 15.610 61.990 15.780 ;
        RECT 61.270 14.920 61.440 15.090 ;
        RECT 61.270 13.570 61.440 13.740 ;
        RECT 60.720 12.840 60.890 13.010 ;
        RECT 60.720 11.470 60.890 11.640 ;
        RECT 60.180 10.790 60.350 10.960 ;
        RECT 62.940 15.790 63.110 15.960 ;
        RECT 62.940 15.430 63.110 15.600 ;
        RECT 63.550 15.790 63.720 15.960 ;
        RECT 63.550 15.430 63.720 15.600 ;
        RECT 64.670 15.610 64.840 15.780 ;
        RECT 62.380 14.910 62.550 15.080 ;
        RECT 64.110 14.910 64.280 15.080 ;
        RECT 62.370 13.570 62.540 13.740 ;
        RECT 64.120 13.570 64.290 13.740 ;
        RECT 61.820 12.840 61.990 13.010 ;
        RECT 61.820 11.470 61.990 11.640 ;
        RECT 61.270 10.790 61.440 10.960 ;
        RECT 65.770 15.620 65.940 15.790 ;
        RECT 65.220 14.920 65.390 15.090 ;
        RECT 65.220 13.570 65.390 13.740 ;
        RECT 64.670 12.840 64.840 13.010 ;
        RECT 64.670 11.470 64.840 11.640 ;
        RECT 62.370 10.800 62.540 10.970 ;
        RECT 64.120 10.800 64.290 10.970 ;
        RECT 66.860 15.620 67.030 15.790 ;
        RECT 66.310 14.940 66.480 15.110 ;
        RECT 66.310 13.570 66.480 13.740 ;
        RECT 65.770 12.840 65.940 13.010 ;
        RECT 65.770 11.470 65.940 11.640 ;
        RECT 65.220 10.790 65.390 10.960 ;
        RECT 70.410 15.600 70.580 15.770 ;
        RECT 69.850 14.900 70.020 15.070 ;
        RECT 69.860 13.560 70.030 13.730 ;
        RECT 66.870 12.840 67.040 13.010 ;
        RECT 66.870 11.470 67.040 11.640 ;
        RECT 66.310 10.790 66.480 10.960 ;
        RECT 71.510 15.610 71.680 15.780 ;
        RECT 70.960 14.910 71.130 15.080 ;
        RECT 70.960 13.560 71.130 13.730 ;
        RECT 70.410 12.830 70.580 13.000 ;
        RECT 70.410 11.460 70.580 11.630 ;
        RECT 67.440 10.830 67.610 11.000 ;
        RECT 59.060 10.360 59.230 10.530 ;
        RECT 69.860 10.790 70.030 10.960 ;
        RECT 72.600 15.610 72.770 15.780 ;
        RECT 72.050 14.930 72.220 15.100 ;
        RECT 72.050 13.560 72.220 13.730 ;
        RECT 71.510 12.830 71.680 13.000 ;
        RECT 71.510 11.460 71.680 11.630 ;
        RECT 70.960 10.780 71.130 10.950 ;
        RECT 72.610 12.830 72.780 13.000 ;
        RECT 73.300 12.530 73.470 12.700 ;
        RECT 73.300 12.170 73.470 12.340 ;
        RECT 72.610 11.460 72.780 11.630 ;
        RECT 72.050 10.780 72.220 10.950 ;
        RECT 73.180 10.820 73.350 10.990 ;
        RECT 67.430 10.360 67.600 10.530 ;
        RECT 73.170 10.350 73.340 10.520 ;
        RECT 18.330 8.660 18.500 8.830 ;
        RECT 104.420 7.820 104.590 7.990 ;
        RECT 109.940 7.080 110.110 7.250 ;
        RECT 18.940 6.370 19.110 6.540 ;
        RECT 15.630 5.930 15.800 6.100 ;
        RECT 16.730 5.940 16.900 6.110 ;
        RECT 16.180 5.260 16.350 5.430 ;
        RECT 16.180 3.890 16.350 4.060 ;
        RECT 15.630 3.160 15.800 3.330 ;
        RECT 15.620 1.820 15.790 1.990 ;
        RECT 15.060 1.300 15.230 1.470 ;
        RECT 17.820 5.940 17.990 6.110 ;
        RECT 17.280 5.260 17.450 5.430 ;
        RECT 17.280 3.890 17.450 4.060 ;
        RECT 16.730 3.160 16.900 3.330 ;
        RECT 16.730 1.810 16.900 1.980 ;
        RECT 16.180 1.120 16.350 1.290 ;
        RECT 104.420 6.210 104.590 6.380 ;
        RECT 18.950 5.900 19.120 6.070 ;
        RECT 109.940 6.410 110.110 6.580 ;
        RECT 18.380 5.260 18.550 5.430 ;
        RECT 18.380 3.890 18.550 4.060 ;
        RECT 17.820 3.160 17.990 3.330 ;
        RECT 17.820 1.790 17.990 1.960 ;
        RECT 17.280 1.110 17.450 1.280 ;
        RECT 20.410 1.770 20.580 5.290 ;
        RECT 20.770 1.770 20.940 5.290 ;
        RECT 21.130 1.770 21.300 5.290 ;
        RECT 21.820 1.770 21.990 5.290 ;
        RECT 22.180 1.770 22.350 5.290 ;
        RECT 22.540 1.770 22.710 5.290 ;
        RECT 104.420 4.610 104.590 4.780 ;
        RECT 104.420 2.990 104.590 3.160 ;
        RECT 106.950 1.830 107.120 2.000 ;
        RECT 104.420 1.390 104.590 1.560 ;
        RECT 18.370 1.110 18.540 1.280 ;
        RECT 104.420 -0.230 104.590 -0.060 ;
        RECT 104.420 -1.830 104.590 -1.660 ;
        RECT 104.420 -3.450 104.590 -3.280 ;
        RECT 110.780 -5.440 110.950 9.510 ;
      LAYER met1 ;
        RECT 82.330 66.110 82.670 66.250 ;
        RECT 90.210 66.110 90.930 67.850 ;
        RECT 82.330 65.390 90.930 66.110 ;
        RECT 30.260 62.940 31.600 63.390 ;
        RECT 4.160 62.100 4.660 62.580 ;
        RECT 30.260 62.520 43.780 62.940 ;
        RECT 45.570 62.850 48.760 63.970 ;
        RECT 30.260 62.380 31.600 62.520 ;
        RECT 4.260 59.140 4.650 62.100 ;
        RECT 24.850 61.780 27.620 62.020 ;
        RECT 6.630 61.320 6.890 61.520 ;
        RECT 9.490 61.480 9.750 61.570 ;
        RECT 6.570 61.010 6.950 61.320 ;
        RECT 7.980 61.010 9.010 61.320 ;
        RECT 9.480 61.250 9.770 61.480 ;
        RECT 6.620 60.220 6.880 60.490 ;
        RECT 7.310 60.220 7.630 60.460 ;
        RECT 8.030 60.220 8.290 60.500 ;
        RECT 6.580 59.560 8.330 60.220 ;
        RECT 6.620 59.300 6.880 59.560 ;
        RECT 7.310 59.300 7.630 59.560 ;
        RECT 8.050 59.320 8.310 59.560 ;
        RECT 4.260 58.650 4.730 59.140 ;
        RECT 4.260 58.640 4.710 58.650 ;
        RECT 4.260 0.530 4.650 58.640 ;
        RECT 6.640 58.270 6.870 58.790 ;
        RECT 6.620 57.950 6.880 58.270 ;
        RECT 5.670 57.500 5.930 57.820 ;
        RECT 5.680 55.280 5.920 57.500 ;
        RECT 6.640 57.380 6.870 57.950 ;
        RECT 8.050 57.380 8.280 58.790 ;
        RECT 8.770 58.240 9.010 61.010 ;
        RECT 24.850 60.690 25.090 61.780 ;
        RECT 9.430 60.560 9.820 60.690 ;
        RECT 9.430 60.270 9.850 60.560 ;
        RECT 24.850 60.430 25.080 60.690 ;
        RECT 9.150 59.710 9.470 60.030 ;
        RECT 9.200 59.480 9.430 59.710 ;
        RECT 9.620 59.330 9.850 60.270 ;
        RECT 24.840 60.210 25.080 60.430 ;
        RECT 22.700 59.400 23.020 59.720 ;
        RECT 24.060 59.480 24.380 59.800 ;
        RECT 24.750 59.470 25.070 59.790 ;
        RECT 9.490 59.260 9.850 59.330 ;
        RECT 9.430 59.150 9.850 59.260 ;
        RECT 9.430 59.030 9.820 59.150 ;
        RECT 8.730 57.700 9.050 58.020 ;
        RECT 9.490 57.860 9.760 59.030 ;
        RECT 24.850 57.890 25.090 58.530 ;
        RECT 9.490 57.630 9.820 57.860 ;
        RECT 24.850 57.630 25.080 57.890 ;
        RECT 24.840 56.980 25.080 57.630 ;
        RECT 7.290 56.500 7.610 56.820 ;
        RECT 8.720 56.520 9.040 56.840 ;
        RECT 6.500 55.920 6.820 56.240 ;
        RECT 7.430 55.920 7.750 56.240 ;
        RECT 8.130 55.920 8.450 56.240 ;
        RECT 8.870 55.920 9.190 56.240 ;
        RECT 9.580 55.910 9.900 56.230 ;
        RECT 5.590 54.800 6.010 55.280 ;
        RECT 11.480 54.040 11.770 56.730 ;
        RECT 24.840 56.340 25.090 56.980 ;
        RECT 21.980 55.740 22.300 56.060 ;
        RECT 11.460 53.370 11.870 54.040 ;
        RECT 24.840 52.680 25.080 56.340 ;
        RECT 24.790 52.340 25.130 52.680 ;
        RECT 22.040 52.240 22.530 52.250 ;
        RECT 18.110 43.550 18.340 47.030 ;
        RECT 18.780 46.410 19.000 47.030 ;
        RECT 19.880 46.600 20.200 46.920 ;
        RECT 20.970 46.610 21.290 46.930 ;
        RECT 18.750 46.090 19.010 46.410 ;
        RECT 19.450 46.100 19.770 46.420 ;
        RECT 18.780 45.490 19.000 46.090 ;
        RECT 19.890 45.610 20.210 45.930 ;
        RECT 20.980 45.620 21.300 45.940 ;
        RECT 18.720 45.170 19.000 45.490 ;
        RECT 19.430 45.180 19.750 45.500 ;
        RECT 18.780 44.570 19.000 45.170 ;
        RECT 19.890 44.620 20.210 44.940 ;
        RECT 20.980 44.630 21.300 44.950 ;
        RECT 18.730 44.250 19.000 44.570 ;
        RECT 18.080 43.230 18.340 43.550 ;
        RECT 18.110 42.590 18.340 43.230 ;
        RECT 18.040 42.270 18.340 42.590 ;
        RECT 18.110 41.630 18.340 42.270 ;
        RECT 18.080 41.310 18.340 41.630 ;
        RECT 18.110 26.560 18.340 41.310 ;
        RECT 18.780 26.560 19.000 44.250 ;
        RECT 19.410 44.190 19.730 44.510 ;
        RECT 19.700 43.690 20.020 44.010 ;
        RECT 21.000 43.590 21.320 43.910 ;
        RECT 19.670 43.510 19.990 43.550 ;
        RECT 19.440 43.280 19.990 43.510 ;
        RECT 19.670 43.230 19.990 43.280 ;
        RECT 19.700 42.700 20.020 43.020 ;
        RECT 21.000 42.600 21.320 42.920 ;
        RECT 19.670 42.520 19.990 42.560 ;
        RECT 19.440 42.290 19.990 42.520 ;
        RECT 21.470 42.390 21.690 51.300 ;
        RECT 22.030 51.090 22.540 52.240 ;
        RECT 27.380 51.310 27.620 61.780 ;
        RECT 30.690 61.450 33.720 61.720 ;
        RECT 30.690 60.470 30.960 61.450 ;
        RECT 30.700 58.260 30.960 58.280 ;
        RECT 30.660 52.280 30.970 58.260 ;
        RECT 31.840 55.760 32.160 56.080 ;
        RECT 30.580 51.910 30.970 52.280 ;
        RECT 33.450 51.770 33.720 61.450 ;
        RECT 35.400 60.430 35.660 62.520 ;
        RECT 43.360 59.270 43.780 62.520 ;
        RECT 47.170 60.030 47.590 62.850 ;
        RECT 74.160 62.840 77.350 63.960 ;
        RECT 47.170 59.550 47.640 60.030 ;
        RECT 43.320 58.790 43.800 59.270 ;
        RECT 66.930 58.770 68.400 59.300 ;
        RECT 34.630 57.720 34.860 57.890 ;
        RECT 34.620 55.850 34.870 57.720 ;
        RECT 48.870 57.180 49.310 57.680 ;
        RECT 54.590 57.180 55.030 57.680 ;
        RECT 44.450 56.160 44.890 56.660 ;
        RECT 34.620 55.670 34.880 55.850 ;
        RECT 34.620 52.770 34.870 55.670 ;
        RECT 41.660 53.420 41.980 53.470 ;
        RECT 41.570 53.130 41.980 53.420 ;
        RECT 34.580 52.410 34.910 52.770 ;
        RECT 33.410 51.460 33.750 51.770 ;
        RECT 21.980 50.990 22.540 51.090 ;
        RECT 27.330 50.990 27.670 51.310 ;
        RECT 21.870 50.590 22.540 50.990 ;
        RECT 41.570 50.700 41.810 53.130 ;
        RECT 44.510 50.700 44.820 56.160 ;
        RECT 21.870 50.560 22.530 50.590 ;
        RECT 21.870 46.340 22.090 50.560 ;
        RECT 41.570 49.630 41.910 50.700 ;
        RECT 43.090 49.990 43.440 50.280 ;
        RECT 43.090 49.970 43.290 49.990 ;
        RECT 40.930 49.130 41.340 49.460 ;
        RECT 23.090 48.440 23.440 48.900 ;
        RECT 39.520 48.460 39.890 48.770 ;
        RECT 22.490 48.080 22.740 48.200 ;
        RECT 22.460 47.620 22.780 48.080 ;
        RECT 21.860 46.050 22.090 46.340 ;
        RECT 19.670 42.240 19.990 42.290 ;
        RECT 21.420 42.160 21.710 42.390 ;
        RECT 19.700 41.710 20.020 42.030 ;
        RECT 21.000 41.610 21.320 41.930 ;
        RECT 19.670 41.530 19.990 41.570 ;
        RECT 19.440 41.300 19.990 41.530 ;
        RECT 19.670 41.250 19.990 41.300 ;
        RECT 18.000 26.030 18.340 26.560 ;
        RECT 18.660 26.030 19.000 26.560 ;
        RECT 16.690 25.290 16.920 25.360 ;
        RECT 16.650 25.030 16.970 25.290 ;
        RECT 16.200 24.920 16.430 24.960 ;
        RECT 16.160 24.600 16.430 24.920 ;
        RECT 6.850 23.360 7.570 24.060 ;
        RECT 6.860 18.210 7.520 23.360 ;
        RECT 16.200 21.080 16.430 24.600 ;
        RECT 16.690 22.560 16.920 25.030 ;
        RECT 18.110 24.940 18.340 26.030 ;
        RECT 18.780 25.300 19.000 26.030 ;
        RECT 20.540 25.320 20.810 25.360 ;
        RECT 18.760 24.980 19.020 25.300 ;
        RECT 20.520 24.990 20.810 25.320 ;
        RECT 18.100 24.620 18.360 24.940 ;
        RECT 18.820 24.020 19.140 24.340 ;
        RECT 19.470 24.020 19.790 24.340 ;
        RECT 17.600 23.580 17.920 23.900 ;
        RECT 18.300 23.580 18.620 23.900 ;
        RECT 19.990 22.570 20.280 23.480 ;
        RECT 16.690 22.550 17.420 22.560 ;
        RECT 16.690 22.230 17.440 22.550 ;
        RECT 16.690 22.190 17.420 22.230 ;
        RECT 16.200 21.010 16.460 21.080 ;
        RECT 16.180 21.000 16.460 21.010 ;
        RECT 16.150 20.690 16.470 21.000 ;
        RECT 12.050 18.830 12.480 19.260 ;
        RECT 6.860 17.490 7.600 18.210 ;
        RECT 12.100 13.020 12.470 18.830 ;
        RECT 16.690 14.690 16.920 22.190 ;
        RECT 17.190 21.940 17.420 22.190 ;
        RECT 19.900 22.000 20.220 22.040 ;
        RECT 20.540 22.020 20.810 24.990 ;
        RECT 20.420 22.000 20.810 22.020 ;
        RECT 17.190 21.720 17.410 21.940 ;
        RECT 19.900 21.770 20.810 22.000 ;
        RECT 21.020 24.920 21.260 24.960 ;
        RECT 21.020 24.600 21.280 24.920 ;
        RECT 19.900 21.720 20.220 21.770 ;
        RECT 17.210 21.290 17.430 21.510 ;
        RECT 17.200 21.000 17.430 21.290 ;
        RECT 19.910 21.460 20.230 21.500 ;
        RECT 21.020 21.460 21.260 24.600 ;
        RECT 19.910 21.230 21.260 21.460 ;
        RECT 19.910 21.180 20.230 21.230 ;
        RECT 17.180 20.680 17.440 21.000 ;
        RECT 19.980 20.550 20.250 20.730 ;
        RECT 19.960 20.230 20.280 20.550 ;
        RECT 19.980 20.060 20.250 20.230 ;
        RECT 17.630 19.700 17.950 20.020 ;
        RECT 18.320 19.690 18.640 20.010 ;
        RECT 18.800 18.920 19.120 19.240 ;
        RECT 19.510 18.860 19.830 19.180 ;
        RECT 16.690 14.460 19.140 14.690 ;
        RECT 18.820 13.840 19.140 14.460 ;
        RECT 15.510 13.400 15.830 13.720 ;
        RECT 16.610 13.410 16.930 13.730 ;
        RECT 17.700 13.410 18.020 13.730 ;
        RECT 18.830 13.370 19.150 13.690 ;
        RECT 12.060 12.590 12.490 13.020 ;
        RECT 16.060 12.730 16.380 13.050 ;
        RECT 17.160 12.730 17.480 13.050 ;
        RECT 18.260 12.730 18.580 13.050 ;
        RECT 18.970 12.560 19.260 12.990 ;
        RECT 19.580 12.560 19.910 12.590 ;
        RECT 18.970 12.540 19.910 12.560 ;
        RECT 18.980 12.240 19.910 12.540 ;
        RECT 18.980 11.710 19.260 12.240 ;
        RECT 19.580 12.170 19.910 12.240 ;
        RECT 18.990 11.680 19.260 11.710 ;
        RECT 16.060 11.360 16.380 11.680 ;
        RECT 17.160 11.360 17.480 11.680 ;
        RECT 18.260 11.360 18.580 11.680 ;
        RECT 15.510 10.630 15.830 10.950 ;
        RECT 16.610 10.630 16.930 10.950 ;
        RECT 17.700 10.630 18.020 10.950 ;
        RECT 15.500 9.290 15.820 9.610 ;
        RECT 16.610 9.280 16.930 9.600 ;
        RECT 17.700 9.260 18.020 9.580 ;
        RECT 16.060 8.590 16.380 8.910 ;
        RECT 17.160 8.580 17.480 8.900 ;
        RECT 18.250 8.580 18.570 8.900 ;
        RECT 15.070 6.930 15.360 7.280 ;
        RECT 15.080 1.640 15.340 6.930 ;
        RECT 18.860 6.290 19.180 6.610 ;
        RECT 21.020 6.570 21.260 21.230 ;
        RECT 21.470 20.560 21.690 42.160 ;
        RECT 21.870 23.170 22.090 46.050 ;
        RECT 22.490 46.830 22.740 47.620 ;
        RECT 22.490 46.510 22.780 46.830 ;
        RECT 22.490 45.910 22.740 46.510 ;
        RECT 22.490 45.590 22.780 45.910 ;
        RECT 22.490 44.990 22.740 45.590 ;
        RECT 22.490 44.670 22.750 44.990 ;
        RECT 22.490 24.320 22.740 44.670 ;
        RECT 23.110 43.900 23.370 48.440 ;
        RECT 38.880 46.740 39.270 47.110 ;
        RECT 38.300 45.250 38.690 45.640 ;
        RECT 23.110 43.580 23.390 43.900 ;
        RECT 37.660 43.660 38.050 44.040 ;
        RECT 37.690 43.650 38.030 43.660 ;
        RECT 23.110 42.940 23.370 43.580 ;
        RECT 37.050 43.460 37.390 43.470 ;
        RECT 37.040 43.070 37.400 43.460 ;
        RECT 23.110 42.620 23.400 42.940 ;
        RECT 23.110 41.980 23.370 42.620 ;
        RECT 23.110 41.660 23.390 41.980 ;
        RECT 22.490 24.300 22.750 24.320 ;
        RECT 22.480 24.020 22.760 24.300 ;
        RECT 22.490 24.000 22.750 24.020 ;
        RECT 21.830 22.850 22.150 23.170 ;
        RECT 21.430 20.240 21.710 20.560 ;
        RECT 21.470 7.270 21.690 20.240 ;
        RECT 21.870 15.030 22.090 22.850 ;
        RECT 21.870 14.550 22.160 15.030 ;
        RECT 21.870 12.590 22.090 14.550 ;
        RECT 21.850 12.170 22.110 12.590 ;
        RECT 21.870 7.550 22.090 12.170 ;
        RECT 22.490 8.930 22.740 24.000 ;
        RECT 23.110 19.990 23.370 41.660 ;
        RECT 36.430 41.510 36.790 41.900 ;
        RECT 35.780 39.970 36.190 40.370 ;
        RECT 35.250 38.410 35.610 38.800 ;
        RECT 34.670 33.350 35.000 33.370 ;
        RECT 34.610 32.930 35.000 33.350 ;
        RECT 34.040 31.740 34.370 31.760 ;
        RECT 33.990 31.350 34.380 31.740 ;
        RECT 33.420 30.190 33.750 30.200 ;
        RECT 33.390 29.800 33.750 30.190 ;
        RECT 32.770 28.320 33.160 28.720 ;
        RECT 32.100 23.150 32.530 23.550 ;
        RECT 31.440 21.580 31.850 21.980 ;
        RECT 23.100 19.670 23.410 19.990 ;
        RECT 30.830 19.940 31.220 20.340 ;
        RECT 22.450 8.530 22.750 8.930 ;
        RECT 21.870 7.410 22.110 7.550 ;
        RECT 21.430 6.920 21.740 7.270 ;
        RECT 21.880 6.780 22.110 7.410 ;
        RECT 15.550 5.850 15.870 6.170 ;
        RECT 16.650 5.860 16.970 6.180 ;
        RECT 17.740 5.860 18.060 6.180 ;
        RECT 18.870 5.820 19.190 6.140 ;
        RECT 20.230 6.010 21.260 6.570 ;
        RECT 21.870 6.750 22.110 6.780 ;
        RECT 20.230 5.900 21.020 6.010 ;
        RECT 16.100 5.180 16.420 5.500 ;
        RECT 17.200 5.180 17.520 5.500 ;
        RECT 18.300 5.180 18.620 5.500 ;
        RECT 21.870 5.360 22.090 6.750 ;
        RECT 16.100 3.810 16.420 4.130 ;
        RECT 17.200 3.810 17.520 4.130 ;
        RECT 18.300 3.810 18.620 4.130 ;
        RECT 15.550 3.080 15.870 3.400 ;
        RECT 16.650 3.080 16.970 3.400 ;
        RECT 17.740 3.080 18.060 3.400 ;
        RECT 15.540 1.740 15.860 2.060 ;
        RECT 16.650 1.730 16.970 2.050 ;
        RECT 17.740 1.710 18.060 2.030 ;
        RECT 20.340 1.680 22.760 5.360 ;
        RECT 15.030 0.830 15.340 1.640 ;
        RECT 23.110 1.390 23.370 19.670 ;
        RECT 30.140 18.500 30.550 18.890 ;
        RECT 25.930 13.350 26.860 15.000 ;
        RECT 26.020 12.870 26.760 13.350 ;
        RECT 16.100 1.040 16.420 1.360 ;
        RECT 17.200 1.030 17.520 1.350 ;
        RECT 18.290 1.030 18.610 1.350 ;
        RECT 23.020 0.980 23.370 1.390 ;
        RECT 15.080 0.630 15.340 0.830 ;
        RECT 4.090 0.010 4.650 0.530 ;
        RECT 30.200 -4.840 30.530 18.500 ;
        RECT 30.150 -4.850 30.580 -4.840 ;
        RECT 30.120 -5.310 30.610 -4.850 ;
        RECT 30.150 -5.330 30.580 -5.310 ;
        RECT 30.850 -5.630 31.180 19.940 ;
        RECT 30.760 -6.120 31.250 -5.630 ;
        RECT 31.500 -6.340 31.830 21.580 ;
        RECT 31.470 -6.800 31.870 -6.340 ;
        RECT 31.260 -7.290 31.840 -7.180 ;
        RECT 32.170 -7.290 32.500 23.150 ;
        RECT 32.810 -2.710 33.140 28.320 ;
        RECT 32.810 -7.170 33.130 -2.710 ;
        RECT 33.420 -6.560 33.750 29.800 ;
        RECT 34.040 -6.310 34.370 31.350 ;
        RECT 34.670 -5.280 35.000 32.930 ;
        RECT 35.270 -4.980 35.600 38.410 ;
        RECT 35.850 -4.410 36.180 39.970 ;
        RECT 36.460 -3.380 36.790 41.510 ;
        RECT 37.050 -2.770 37.380 43.070 ;
        RECT 37.690 -2.100 38.020 43.650 ;
        RECT 38.310 -1.450 38.640 45.250 ;
        RECT 38.910 -0.820 39.240 46.740 ;
        RECT 39.540 -0.210 39.870 48.460 ;
        RECT 40.930 47.380 41.340 47.710 ;
        RECT 40.930 45.630 41.340 45.960 ;
        RECT 40.930 43.880 41.340 44.210 ;
        RECT 40.930 43.080 41.340 43.410 ;
        RECT 40.930 41.330 41.340 41.660 ;
        RECT 40.930 39.580 41.340 39.910 ;
        RECT 40.930 37.830 41.340 38.160 ;
        RECT 41.670 37.550 41.910 49.630 ;
        RECT 44.510 49.560 44.920 50.700 ;
        RECT 46.830 50.270 47.140 50.280 ;
        RECT 46.830 50.000 47.150 50.270 ;
        RECT 47.870 50.040 48.190 50.340 ;
        RECT 46.850 49.990 47.140 50.000 ;
        RECT 43.090 48.240 43.440 48.530 ;
        RECT 43.090 48.220 43.290 48.240 ;
        RECT 43.090 46.490 43.440 46.780 ;
        RECT 43.090 46.470 43.290 46.490 ;
        RECT 43.090 44.740 43.440 45.030 ;
        RECT 43.090 44.720 43.290 44.740 ;
        RECT 43.090 42.550 43.290 42.570 ;
        RECT 43.090 42.260 43.440 42.550 ;
        RECT 43.090 40.800 43.290 40.820 ;
        RECT 43.090 40.510 43.440 40.800 ;
        RECT 43.090 39.050 43.290 39.070 ;
        RECT 43.090 38.760 43.440 39.050 ;
        RECT 44.610 37.620 44.920 49.560 ;
        RECT 45.170 49.240 45.450 49.570 ;
        RECT 46.830 48.520 47.140 48.530 ;
        RECT 46.830 48.250 47.150 48.520 ;
        RECT 47.870 48.290 48.190 48.590 ;
        RECT 46.850 48.240 47.140 48.250 ;
        RECT 45.170 47.490 45.450 47.820 ;
        RECT 46.830 46.770 47.140 46.780 ;
        RECT 46.830 46.500 47.150 46.770 ;
        RECT 47.870 46.540 48.190 46.840 ;
        RECT 46.850 46.490 47.140 46.500 ;
        RECT 45.170 45.740 45.450 46.070 ;
        RECT 46.830 45.020 47.140 45.030 ;
        RECT 46.830 44.750 47.150 45.020 ;
        RECT 47.870 44.790 48.190 45.090 ;
        RECT 46.850 44.740 47.140 44.750 ;
        RECT 45.170 43.990 45.450 44.320 ;
        RECT 45.170 42.970 45.450 43.300 ;
        RECT 46.850 42.540 47.140 42.550 ;
        RECT 46.830 42.270 47.150 42.540 ;
        RECT 46.830 42.260 47.140 42.270 ;
        RECT 47.870 42.200 48.190 42.500 ;
        RECT 45.170 41.220 45.450 41.550 ;
        RECT 46.850 40.790 47.140 40.800 ;
        RECT 46.830 40.520 47.150 40.790 ;
        RECT 46.830 40.510 47.140 40.520 ;
        RECT 47.870 40.450 48.190 40.750 ;
        RECT 45.170 39.470 45.450 39.800 ;
        RECT 46.850 39.040 47.140 39.050 ;
        RECT 46.830 38.770 47.150 39.040 ;
        RECT 46.830 38.760 47.140 38.770 ;
        RECT 47.870 38.700 48.190 39.000 ;
        RECT 45.170 37.720 45.450 38.050 ;
        RECT 41.570 36.590 41.910 37.550 ;
        RECT 43.090 37.300 43.290 37.320 ;
        RECT 43.090 37.010 43.440 37.300 ;
        RECT 44.510 36.590 44.920 37.620 ;
        RECT 46.850 37.290 47.140 37.300 ;
        RECT 46.830 37.020 47.150 37.290 ;
        RECT 46.830 37.010 47.140 37.020 ;
        RECT 47.870 36.950 48.190 37.250 ;
        RECT 41.570 33.460 41.810 36.590 ;
        RECT 44.510 33.460 44.820 36.590 ;
        RECT 40.930 32.950 41.340 33.280 ;
        RECT 41.570 33.180 41.910 33.460 ;
        RECT 40.930 31.200 41.340 31.530 ;
        RECT 40.930 29.450 41.340 29.780 ;
        RECT 40.930 27.700 41.340 28.030 ;
        RECT 41.670 27.420 41.910 33.180 ;
        RECT 44.510 33.110 44.920 33.460 ;
        RECT 43.090 32.420 43.290 32.440 ;
        RECT 43.090 32.130 43.440 32.420 ;
        RECT 43.090 30.670 43.290 30.690 ;
        RECT 43.090 30.380 43.440 30.670 ;
        RECT 43.090 28.920 43.290 28.940 ;
        RECT 43.090 28.630 43.440 28.920 ;
        RECT 44.610 27.490 44.920 33.110 ;
        RECT 45.170 32.840 45.450 33.170 ;
        RECT 46.850 32.410 47.140 32.420 ;
        RECT 46.830 32.140 47.150 32.410 ;
        RECT 46.830 32.130 47.140 32.140 ;
        RECT 47.870 32.070 48.190 32.370 ;
        RECT 45.170 31.090 45.450 31.420 ;
        RECT 46.850 30.660 47.140 30.670 ;
        RECT 46.830 30.390 47.150 30.660 ;
        RECT 46.830 30.380 47.140 30.390 ;
        RECT 47.870 30.320 48.190 30.620 ;
        RECT 45.170 29.340 45.450 29.670 ;
        RECT 46.850 28.910 47.140 28.920 ;
        RECT 46.830 28.640 47.150 28.910 ;
        RECT 46.830 28.630 47.140 28.640 ;
        RECT 47.870 28.570 48.190 28.870 ;
        RECT 45.170 27.590 45.450 27.920 ;
        RECT 40.890 23.890 41.300 24.220 ;
        RECT 41.570 23.650 41.910 27.420 ;
        RECT 43.090 27.170 43.290 27.190 ;
        RECT 43.090 26.880 43.440 27.170 ;
        RECT 44.510 23.650 44.920 27.490 ;
        RECT 46.850 27.160 47.140 27.170 ;
        RECT 46.830 26.890 47.150 27.160 ;
        RECT 46.830 26.880 47.140 26.890 ;
        RECT 47.870 26.820 48.190 27.120 ;
        RECT 48.940 24.400 49.230 57.180 ;
        RECT 50.130 56.190 50.630 56.630 ;
        RECT 50.400 43.460 50.590 56.190 ;
        RECT 50.120 42.970 50.590 43.460 ;
        RECT 50.980 43.320 51.350 43.340 ;
        RECT 50.930 43.060 51.350 43.320 ;
        RECT 50.980 43.050 51.350 43.060 ;
        RECT 49.940 42.530 50.260 42.810 ;
        RECT 50.400 42.710 50.590 42.970 ;
        RECT 50.400 42.420 50.630 42.710 ;
        RECT 50.400 41.650 50.590 42.420 ;
        RECT 49.940 41.260 50.260 41.540 ;
        RECT 50.400 41.360 50.630 41.650 ;
        RECT 50.400 41.100 50.590 41.360 ;
        RECT 50.120 40.610 50.590 41.100 ;
        RECT 50.980 41.010 51.350 41.020 ;
        RECT 50.930 40.750 51.350 41.010 ;
        RECT 50.980 40.730 51.350 40.750 ;
        RECT 50.400 40.260 50.590 40.610 ;
        RECT 50.120 39.770 50.590 40.260 ;
        RECT 50.980 40.120 51.350 40.140 ;
        RECT 50.930 39.860 51.350 40.120 ;
        RECT 50.980 39.850 51.350 39.860 ;
        RECT 49.940 39.330 50.260 39.610 ;
        RECT 50.400 39.510 50.590 39.770 ;
        RECT 50.400 39.220 50.630 39.510 ;
        RECT 50.400 38.450 50.590 39.220 ;
        RECT 49.940 38.060 50.260 38.340 ;
        RECT 50.400 38.160 50.630 38.450 ;
        RECT 50.400 37.900 50.590 38.160 ;
        RECT 50.120 37.410 50.590 37.900 ;
        RECT 50.980 37.810 51.350 37.820 ;
        RECT 50.930 37.550 51.350 37.810 ;
        RECT 50.980 37.530 51.350 37.550 ;
        RECT 50.400 33.640 50.590 37.410 ;
        RECT 51.710 33.740 51.940 43.680 ;
        RECT 54.680 43.460 54.930 57.180 ;
        RECT 64.560 56.160 65.000 56.660 ;
        RECT 58.760 52.410 59.100 52.700 ;
        RECT 58.810 52.380 59.070 52.410 ;
        RECT 56.930 48.850 57.190 49.170 ;
        RECT 56.960 45.350 57.150 48.850 ;
        RECT 58.830 46.440 59.040 52.380 ;
        RECT 62.400 51.780 62.660 51.790 ;
        RECT 62.380 51.480 62.680 51.780 ;
        RECT 62.400 51.470 62.660 51.480 ;
        RECT 59.230 50.450 59.570 50.770 ;
        RECT 58.360 45.990 58.670 46.430 ;
        RECT 58.820 46.150 59.050 46.440 ;
        RECT 56.930 45.320 57.150 45.350 ;
        RECT 56.920 45.050 57.170 45.320 ;
        RECT 56.920 45.040 57.160 45.050 ;
        RECT 56.930 44.800 57.160 45.040 ;
        RECT 53.440 43.300 53.780 43.350 ;
        RECT 53.440 43.280 54.000 43.300 ;
        RECT 53.320 43.110 54.000 43.280 ;
        RECT 53.440 43.070 54.000 43.110 ;
        RECT 53.440 43.030 53.780 43.070 ;
        RECT 54.680 42.390 55.320 43.460 ;
        RECT 56.960 42.770 57.120 44.800 ;
        RECT 57.960 44.460 58.280 44.780 ;
        RECT 58.830 44.450 59.040 46.150 ;
        RECT 59.300 45.880 59.490 50.450 ;
        RECT 59.670 48.360 59.960 48.680 ;
        RECT 59.290 45.590 59.520 45.880 ;
        RECT 57.310 43.950 57.550 44.370 ;
        RECT 58.820 44.160 59.050 44.450 ;
        RECT 58.830 44.020 59.040 44.160 ;
        RECT 57.280 43.630 57.550 43.950 ;
        RECT 57.310 43.200 57.550 43.630 ;
        RECT 59.300 43.560 59.490 45.590 ;
        RECT 59.710 44.090 59.920 48.360 ;
        RECT 60.710 47.880 61.050 48.200 ;
        RECT 59.680 43.580 59.920 44.090 ;
        RECT 58.850 43.380 59.040 43.510 ;
        RECT 58.830 43.090 59.060 43.380 ;
        RECT 59.290 43.270 59.520 43.560 ;
        RECT 57.950 42.770 58.270 43.090 ;
        RECT 56.930 42.530 57.160 42.770 ;
        RECT 56.920 42.520 57.160 42.530 ;
        RECT 54.680 41.680 54.930 42.390 ;
        RECT 56.920 42.250 57.170 42.520 ;
        RECT 56.930 42.220 57.150 42.250 ;
        RECT 53.440 41.000 53.780 41.040 ;
        RECT 53.440 40.960 54.000 41.000 ;
        RECT 53.320 40.790 54.000 40.960 ;
        RECT 53.440 40.770 54.000 40.790 ;
        RECT 53.440 40.720 53.780 40.770 ;
        RECT 54.680 40.610 55.320 41.680 ;
        RECT 56.960 40.780 57.150 42.220 ;
        RECT 58.360 41.140 58.670 41.580 ;
        RECT 58.850 41.470 59.040 43.090 ;
        RECT 59.300 41.980 59.490 43.270 ;
        RECT 59.280 41.690 59.510 41.980 ;
        RECT 58.850 41.260 59.080 41.470 ;
        RECT 58.840 41.180 59.080 41.260 ;
        RECT 56.960 40.760 57.160 40.780 ;
        RECT 58.840 40.760 59.070 41.180 ;
        RECT 59.300 40.760 59.490 41.690 ;
        RECT 59.710 40.760 59.920 43.580 ;
        RECT 60.790 42.280 60.970 47.880 ;
        RECT 61.510 44.810 61.770 45.600 ;
        RECT 60.730 41.940 61.020 42.280 ;
        RECT 60.790 40.760 60.970 41.940 ;
        RECT 61.510 41.870 61.770 42.660 ;
        RECT 62.430 41.240 62.630 51.470 ;
        RECT 62.410 41.110 62.630 41.240 ;
        RECT 64.660 41.110 64.890 56.160 ;
        RECT 65.560 52.390 65.840 52.710 ;
        RECT 65.120 51.480 65.400 51.800 ;
        RECT 62.360 40.780 62.690 41.110 ;
        RECT 64.610 40.810 64.930 41.110 ;
        RECT 54.680 40.260 54.930 40.610 ;
        RECT 53.440 40.100 53.780 40.150 ;
        RECT 53.440 40.080 54.000 40.100 ;
        RECT 53.320 39.910 54.000 40.080 ;
        RECT 53.440 39.870 54.000 39.910 ;
        RECT 53.440 39.830 53.780 39.870 ;
        RECT 54.680 39.190 55.320 40.260 ;
        RECT 56.970 39.320 57.160 40.760 ;
        RECT 58.370 39.960 58.680 40.400 ;
        RECT 63.450 39.570 63.680 40.780 ;
        RECT 64.660 40.760 64.900 40.810 ;
        RECT 64.670 39.810 64.900 40.760 ;
        RECT 65.150 39.940 65.370 51.480 ;
        RECT 65.140 39.870 65.370 39.940 ;
        RECT 56.940 39.290 57.160 39.320 ;
        RECT 54.680 38.480 54.930 39.190 ;
        RECT 56.930 39.020 57.180 39.290 ;
        RECT 56.930 39.010 57.170 39.020 ;
        RECT 56.940 38.770 57.170 39.010 ;
        RECT 58.210 39.000 58.530 39.320 ;
        RECT 63.420 38.780 63.680 39.570 ;
        RECT 64.660 39.560 64.900 39.810 ;
        RECT 53.440 37.800 53.780 37.840 ;
        RECT 53.440 37.760 54.000 37.800 ;
        RECT 53.320 37.590 54.000 37.760 ;
        RECT 53.440 37.570 54.000 37.590 ;
        RECT 53.440 37.520 53.780 37.570 ;
        RECT 54.680 37.410 55.320 38.480 ;
        RECT 54.680 33.750 54.930 37.410 ;
        RECT 56.970 36.740 57.130 38.770 ;
        RECT 57.320 38.210 57.560 38.340 ;
        RECT 57.300 37.890 57.560 38.210 ;
        RECT 57.300 37.290 57.560 37.610 ;
        RECT 57.320 37.170 57.560 37.290 ;
        RECT 56.940 36.500 57.170 36.740 ;
        RECT 63.450 36.630 63.680 38.780 ;
        RECT 56.930 36.490 57.170 36.500 ;
        RECT 56.930 36.220 57.180 36.490 ;
        RECT 58.210 36.240 58.530 36.560 ;
        RECT 56.940 36.190 57.160 36.220 ;
        RECT 56.970 34.320 57.160 36.190 ;
        RECT 63.420 35.840 63.680 36.630 ;
        RECT 58.370 35.110 58.680 35.550 ;
        RECT 58.970 34.480 59.360 34.500 ;
        RECT 58.960 34.390 59.360 34.480 ;
        RECT 58.810 34.380 59.360 34.390 ;
        RECT 56.970 34.130 58.570 34.320 ;
        RECT 50.380 33.140 50.590 33.640 ;
        RECT 51.690 33.330 51.940 33.740 ;
        RECT 54.660 33.330 54.930 33.750 ;
        RECT 50.380 32.990 50.570 33.140 ;
        RECT 50.100 32.500 50.570 32.990 ;
        RECT 50.960 32.850 51.330 32.870 ;
        RECT 50.910 32.590 51.330 32.850 ;
        RECT 50.960 32.580 51.330 32.590 ;
        RECT 49.920 32.060 50.240 32.340 ;
        RECT 50.380 32.240 50.570 32.500 ;
        RECT 50.380 31.950 50.610 32.240 ;
        RECT 50.380 31.180 50.570 31.950 ;
        RECT 49.920 30.790 50.240 31.070 ;
        RECT 50.380 30.890 50.610 31.180 ;
        RECT 50.380 30.630 50.570 30.890 ;
        RECT 50.100 30.140 50.570 30.630 ;
        RECT 50.960 30.540 51.330 30.550 ;
        RECT 50.910 30.280 51.330 30.540 ;
        RECT 50.960 30.260 51.330 30.280 ;
        RECT 50.380 29.790 50.570 30.140 ;
        RECT 50.100 29.300 50.570 29.790 ;
        RECT 50.960 29.650 51.330 29.670 ;
        RECT 50.910 29.390 51.330 29.650 ;
        RECT 50.960 29.380 51.330 29.390 ;
        RECT 49.920 28.860 50.240 29.140 ;
        RECT 50.380 29.040 50.570 29.300 ;
        RECT 50.380 28.750 50.610 29.040 ;
        RECT 50.380 27.980 50.570 28.750 ;
        RECT 49.920 27.590 50.240 27.870 ;
        RECT 50.380 27.690 50.610 27.980 ;
        RECT 50.380 27.470 50.570 27.690 ;
        RECT 51.690 27.510 51.920 33.330 ;
        RECT 54.660 32.990 54.910 33.330 ;
        RECT 53.420 32.830 53.760 32.880 ;
        RECT 53.420 32.810 53.980 32.830 ;
        RECT 53.300 32.640 53.980 32.810 ;
        RECT 53.420 32.600 53.980 32.640 ;
        RECT 53.420 32.560 53.760 32.600 ;
        RECT 54.660 31.920 55.300 32.990 ;
        RECT 58.380 32.210 58.570 34.130 ;
        RECT 58.780 34.140 59.360 34.380 ;
        RECT 58.780 34.120 59.350 34.140 ;
        RECT 58.780 34.110 58.970 34.120 ;
        RECT 58.780 33.270 58.950 34.110 ;
        RECT 63.450 34.050 63.680 35.840 ;
        RECT 64.670 37.670 64.900 39.560 ;
        RECT 65.130 39.270 65.330 39.870 ;
        RECT 65.580 39.730 65.810 52.390 ;
        RECT 66.950 46.660 67.370 58.770 ;
        RECT 67.980 46.660 68.400 58.770 ;
        RECT 70.360 56.120 70.800 56.620 ;
        RECT 70.460 49.140 70.690 56.120 ;
        RECT 74.880 50.870 76.160 62.840 ;
        RECT 78.640 57.650 78.920 57.770 ;
        RECT 78.640 57.150 78.970 57.650 ;
        RECT 74.880 50.790 76.180 50.870 ;
        RECT 74.870 50.490 76.180 50.790 ;
        RECT 71.650 49.840 71.950 50.160 ;
        RECT 70.330 49.130 70.690 49.140 ;
        RECT 70.300 48.240 70.690 49.130 ;
        RECT 66.950 46.520 68.400 46.660 ;
        RECT 66.950 40.780 67.370 46.520 ;
        RECT 67.980 40.780 68.400 46.520 ;
        RECT 70.460 41.110 70.690 48.240 ;
        RECT 71.680 45.600 71.910 49.840 ;
        RECT 77.960 49.290 78.390 49.630 ;
        RECT 76.680 45.990 76.990 46.430 ;
        RECT 71.680 44.810 71.940 45.600 ;
        RECT 78.200 45.350 78.390 49.290 ;
        RECT 78.640 46.790 78.920 57.150 ;
        RECT 80.340 52.390 80.600 52.710 ;
        RECT 79.450 51.520 79.710 51.840 ;
        RECT 79.480 47.800 79.670 51.520 ;
        RECT 80.360 47.800 80.580 52.390 ;
        RECT 82.330 49.170 82.670 65.390 ;
        RECT 102.730 62.870 105.920 63.990 ;
        RECT 86.830 61.930 87.200 61.940 ;
        RECT 86.780 61.480 87.280 61.930 ;
        RECT 82.980 53.070 83.300 53.440 ;
        RECT 82.280 49.090 82.670 49.170 ;
        RECT 82.270 48.320 82.670 49.090 ;
        RECT 82.280 48.250 82.670 48.320 ;
        RECT 79.310 47.110 79.990 47.800 ;
        RECT 80.350 47.110 81.030 47.800 ;
        RECT 78.640 46.490 78.980 46.790 ;
        RECT 78.640 46.160 78.920 46.490 ;
        RECT 80.390 46.470 80.710 46.790 ;
        RECT 81.370 46.220 81.690 46.540 ;
        RECT 78.530 45.560 78.920 46.160 ;
        RECT 80.540 45.640 80.860 45.960 ;
        RECT 81.320 45.570 81.640 45.890 ;
        RECT 76.830 45.030 77.150 45.350 ;
        RECT 78.200 45.320 78.420 45.350 ;
        RECT 78.180 45.050 78.430 45.320 ;
        RECT 78.190 45.040 78.430 45.050 ;
        RECT 71.680 42.660 71.910 44.810 ;
        RECT 78.190 44.800 78.420 45.040 ;
        RECT 77.800 44.240 78.040 44.370 ;
        RECT 77.800 43.920 78.060 44.240 ;
        RECT 77.800 43.320 78.060 43.640 ;
        RECT 77.800 43.200 78.040 43.320 ;
        RECT 78.230 42.770 78.390 44.800 ;
        RECT 78.640 43.960 78.920 45.560 ;
        RECT 79.430 45.110 79.750 45.430 ;
        RECT 80.650 44.950 80.860 45.060 ;
        RECT 80.630 44.630 80.890 44.950 ;
        RECT 81.320 44.720 81.640 45.040 ;
        RECT 78.640 43.640 79.000 43.960 ;
        RECT 80.160 43.830 80.480 44.150 ;
        RECT 71.680 41.870 71.940 42.660 ;
        RECT 76.830 42.270 77.150 42.590 ;
        RECT 78.190 42.530 78.420 42.770 ;
        RECT 78.190 42.520 78.430 42.530 ;
        RECT 78.180 42.250 78.430 42.520 ;
        RECT 78.200 42.220 78.420 42.250 ;
        RECT 70.410 40.810 70.730 41.110 ;
        RECT 66.950 40.760 68.400 40.780 ;
        RECT 65.470 39.420 65.810 39.730 ;
        RECT 66.960 40.620 68.400 40.760 ;
        RECT 65.470 39.410 65.790 39.420 ;
        RECT 65.140 39.240 65.370 39.270 ;
        RECT 64.670 37.370 65.000 37.670 ;
        RECT 64.670 37.200 64.920 37.370 ;
        RECT 64.670 34.080 64.900 37.200 ;
        RECT 65.150 36.040 65.370 39.240 ;
        RECT 65.150 35.730 65.820 36.040 ;
        RECT 65.500 35.720 65.820 35.730 ;
        RECT 66.960 34.740 67.380 40.620 ;
        RECT 62.930 33.980 63.680 34.050 ;
        RECT 62.900 33.820 63.680 33.980 ;
        RECT 64.650 34.020 64.900 34.080 ;
        RECT 67.980 34.150 68.400 40.620 ;
        RECT 70.460 37.620 70.690 40.810 ;
        RECT 71.680 39.570 71.910 41.870 ;
        RECT 76.680 41.140 76.990 41.580 ;
        RECT 76.680 39.960 76.990 40.400 ;
        RECT 71.680 38.780 71.940 39.570 ;
        RECT 78.200 39.320 78.390 42.220 ;
        RECT 78.640 42.010 78.920 43.640 ;
        RECT 80.650 43.340 80.860 44.630 ;
        RECT 81.370 44.070 81.690 44.390 ;
        RECT 80.630 43.050 80.860 43.340 ;
        RECT 81.370 43.220 81.690 43.540 ;
        RECT 81.320 42.570 81.640 42.890 ;
        RECT 78.530 41.410 78.920 42.010 ;
        RECT 81.320 41.720 81.640 42.040 ;
        RECT 78.640 40.730 78.920 41.410 ;
        RECT 80.800 40.960 81.120 41.260 ;
        RECT 81.370 41.070 81.690 41.390 ;
        RECT 82.330 40.960 82.670 48.250 ;
        RECT 83.000 47.690 83.270 53.070 ;
        RECT 83.000 47.190 83.680 47.690 ;
        RECT 83.000 46.810 83.270 47.190 ;
        RECT 82.990 46.660 83.270 46.810 ;
        RECT 80.800 40.930 81.230 40.960 ;
        RECT 81.830 40.930 82.670 40.960 ;
        RECT 80.800 40.900 82.670 40.930 ;
        RECT 80.950 40.850 82.670 40.900 ;
        RECT 80.980 40.820 82.670 40.850 ;
        RECT 81.010 40.800 82.670 40.820 ;
        RECT 81.080 40.790 82.040 40.800 ;
        RECT 78.640 40.430 78.960 40.730 ;
        RECT 80.390 40.440 80.710 40.760 ;
        RECT 78.640 40.130 78.920 40.430 ;
        RECT 81.370 40.190 81.690 40.510 ;
        RECT 78.530 39.530 78.920 40.130 ;
        RECT 80.540 39.610 80.860 39.930 ;
        RECT 81.320 39.540 81.640 39.860 ;
        RECT 76.830 39.000 77.150 39.320 ;
        RECT 78.200 39.290 78.420 39.320 ;
        RECT 78.180 39.020 78.430 39.290 ;
        RECT 78.190 39.010 78.430 39.020 ;
        RECT 70.380 37.300 70.700 37.620 ;
        RECT 70.460 35.090 70.690 37.300 ;
        RECT 71.680 36.630 71.910 38.780 ;
        RECT 78.190 38.770 78.420 39.010 ;
        RECT 77.800 38.210 78.040 38.340 ;
        RECT 77.800 37.890 78.060 38.210 ;
        RECT 77.800 37.290 78.060 37.610 ;
        RECT 77.800 37.170 78.040 37.290 ;
        RECT 78.230 36.740 78.390 38.770 ;
        RECT 78.640 37.930 78.920 39.530 ;
        RECT 79.430 39.080 79.750 39.400 ;
        RECT 80.650 38.920 80.860 39.030 ;
        RECT 80.630 38.600 80.890 38.920 ;
        RECT 81.320 38.690 81.640 39.010 ;
        RECT 78.640 37.610 79.000 37.930 ;
        RECT 80.160 37.800 80.480 38.120 ;
        RECT 71.680 35.840 71.940 36.630 ;
        RECT 76.830 36.240 77.150 36.560 ;
        RECT 78.190 36.500 78.420 36.740 ;
        RECT 78.190 36.490 78.430 36.500 ;
        RECT 78.180 36.220 78.430 36.490 ;
        RECT 78.200 36.190 78.420 36.220 ;
        RECT 70.380 34.790 70.700 35.090 ;
        RECT 62.900 33.370 63.310 33.820 ;
        RECT 58.780 32.520 58.940 33.270 ;
        RECT 58.740 32.500 58.940 32.520 ;
        RECT 59.760 32.510 60.080 32.830 ;
        RECT 58.730 32.260 58.960 32.500 ;
        RECT 58.730 32.210 58.940 32.260 ;
        RECT 58.380 32.090 58.550 32.210 ;
        RECT 54.660 31.210 54.910 31.920 ;
        RECT 53.420 30.530 53.760 30.570 ;
        RECT 53.420 30.490 53.980 30.530 ;
        RECT 53.300 30.320 53.980 30.490 ;
        RECT 53.420 30.300 53.980 30.320 ;
        RECT 53.420 30.250 53.760 30.300 ;
        RECT 54.660 30.140 55.300 31.210 ;
        RECT 58.380 31.160 58.540 32.090 ;
        RECT 58.380 31.040 58.550 31.160 ;
        RECT 58.780 31.040 58.940 32.210 ;
        RECT 59.760 31.960 60.080 32.280 ;
        RECT 60.720 31.870 60.960 33.260 ;
        RECT 54.660 29.790 54.910 30.140 ;
        RECT 58.380 30.120 58.570 31.040 ;
        RECT 58.730 30.990 58.940 31.040 ;
        RECT 58.730 30.750 58.960 30.990 ;
        RECT 59.760 30.970 60.080 31.290 ;
        RECT 60.710 31.210 60.980 31.870 ;
        RECT 58.740 30.730 58.940 30.750 ;
        RECT 58.350 30.100 58.590 30.120 ;
        RECT 58.780 30.100 58.940 30.730 ;
        RECT 59.760 30.420 60.080 30.740 ;
        RECT 58.350 29.910 58.940 30.100 ;
        RECT 58.350 29.890 58.590 29.910 ;
        RECT 53.420 29.630 53.760 29.680 ;
        RECT 53.420 29.610 53.980 29.630 ;
        RECT 53.300 29.440 53.980 29.610 ;
        RECT 53.420 29.400 53.980 29.440 ;
        RECT 53.420 29.360 53.760 29.400 ;
        RECT 54.660 28.720 55.300 29.790 ;
        RECT 58.380 28.970 58.570 29.890 ;
        RECT 58.780 29.280 58.940 29.910 ;
        RECT 58.740 29.260 58.940 29.280 ;
        RECT 59.760 29.270 60.080 29.590 ;
        RECT 58.730 29.020 58.960 29.260 ;
        RECT 58.730 28.970 58.940 29.020 ;
        RECT 58.380 28.850 58.550 28.970 ;
        RECT 54.660 28.010 54.910 28.720 ;
        RECT 50.380 27.430 50.590 27.470 ;
        RECT 50.100 26.940 50.590 27.430 ;
        RECT 50.960 27.340 51.330 27.350 ;
        RECT 50.910 27.080 51.330 27.340 ;
        RECT 50.960 27.060 51.330 27.080 ;
        RECT 50.380 26.720 50.590 26.940 ;
        RECT 51.690 26.720 51.940 27.510 ;
        RECT 53.420 27.330 53.760 27.370 ;
        RECT 53.420 27.290 53.980 27.330 ;
        RECT 53.300 27.120 53.980 27.290 ;
        RECT 53.420 27.100 53.980 27.120 ;
        RECT 53.420 27.050 53.760 27.100 ;
        RECT 54.660 26.940 55.300 28.010 ;
        RECT 58.380 27.930 58.540 28.850 ;
        RECT 58.380 27.810 58.550 27.930 ;
        RECT 58.780 27.810 58.940 28.970 ;
        RECT 59.760 28.720 60.080 29.040 ;
        RECT 60.720 28.620 60.960 31.210 ;
        RECT 62.900 31.110 63.280 33.370 ;
        RECT 64.650 31.850 64.890 34.020 ;
        RECT 67.980 33.970 68.410 34.150 ;
        RECT 67.980 33.580 68.420 33.970 ;
        RECT 70.460 33.760 70.690 34.790 ;
        RECT 68.010 33.370 68.420 33.580 ;
        RECT 66.930 32.890 67.330 33.260 ;
        RECT 68.010 32.890 68.410 33.370 ;
        RECT 66.930 32.670 68.410 32.890 ;
        RECT 64.640 31.190 64.900 31.850 ;
        RECT 62.900 29.250 63.290 31.110 ;
        RECT 60.710 28.300 60.970 28.620 ;
        RECT 54.660 26.720 54.930 26.940 ;
        RECT 58.380 26.820 58.570 27.810 ;
        RECT 58.730 27.760 58.940 27.810 ;
        RECT 58.730 27.520 58.960 27.760 ;
        RECT 59.760 27.740 60.080 28.060 ;
        RECT 60.720 27.620 60.960 28.300 ;
        RECT 62.900 27.760 63.280 29.250 ;
        RECT 64.650 28.580 64.890 31.190 ;
        RECT 64.640 28.260 64.900 28.580 ;
        RECT 58.740 27.500 58.940 27.520 ;
        RECT 58.780 26.770 58.940 27.500 ;
        RECT 59.760 27.190 60.080 27.510 ;
        RECT 60.720 26.760 60.990 27.620 ;
        RECT 62.900 26.760 63.310 27.760 ;
        RECT 64.650 27.620 64.890 28.260 ;
        RECT 66.930 27.780 67.330 32.670 ;
        RECT 64.650 26.760 64.920 27.620 ;
        RECT 66.930 26.760 67.360 27.780 ;
        RECT 68.010 26.760 68.410 32.670 ;
        RECT 70.450 31.850 70.690 33.760 ;
        RECT 71.680 34.070 71.910 35.840 ;
        RECT 76.680 35.110 76.990 35.550 ;
        RECT 71.680 33.690 72.440 34.070 ;
        RECT 78.200 33.940 78.390 36.190 ;
        RECT 78.640 35.980 78.920 37.610 ;
        RECT 80.650 37.310 80.860 38.600 ;
        RECT 81.370 38.040 81.690 38.360 ;
        RECT 80.630 37.020 80.860 37.310 ;
        RECT 81.370 37.190 81.690 37.510 ;
        RECT 81.320 36.540 81.640 36.860 ;
        RECT 78.530 35.380 78.920 35.980 ;
        RECT 81.320 35.690 81.640 36.010 ;
        RECT 70.440 31.190 70.700 31.850 ;
        RECT 70.450 28.580 70.690 31.190 ;
        RECT 72.060 31.110 72.440 33.690 ;
        RECT 76.370 33.570 76.650 33.890 ;
        RECT 76.800 33.750 78.390 33.940 ;
        RECT 74.380 31.870 74.620 33.260 ;
        RECT 75.260 32.510 75.580 32.830 ;
        RECT 76.400 32.520 76.560 33.570 ;
        RECT 76.800 33.420 76.990 33.750 ;
        RECT 78.640 33.560 78.920 35.380 ;
        RECT 80.820 34.930 81.150 35.220 ;
        RECT 81.370 35.040 81.690 35.360 ;
        RECT 82.330 34.930 82.670 40.800 ;
        RECT 83.000 45.230 83.270 46.660 ;
        RECT 83.620 46.240 83.940 46.560 ;
        RECT 83.000 44.940 83.280 45.230 ;
        RECT 83.000 42.640 83.270 44.940 ;
        RECT 83.670 44.020 83.990 44.340 ;
        RECT 83.660 43.300 83.980 43.620 ;
        RECT 83.000 42.350 83.280 42.640 ;
        RECT 83.000 40.780 83.270 42.350 ;
        RECT 83.580 41.050 83.900 41.370 ;
        RECT 82.990 40.630 83.270 40.780 ;
        RECT 80.810 34.900 81.230 34.930 ;
        RECT 81.830 34.900 82.670 34.930 ;
        RECT 80.810 34.790 82.670 34.900 ;
        RECT 81.090 34.760 81.990 34.790 ;
        RECT 82.330 34.730 82.670 34.790 ;
        RECT 83.000 39.200 83.270 40.630 ;
        RECT 83.620 40.210 83.940 40.530 ;
        RECT 83.000 38.910 83.280 39.200 ;
        RECT 83.000 36.610 83.270 38.910 ;
        RECT 83.670 37.990 83.990 38.310 ;
        RECT 83.660 37.270 83.980 37.590 ;
        RECT 83.000 36.320 83.280 36.610 ;
        RECT 83.000 34.730 83.270 36.320 ;
        RECT 83.580 35.020 83.900 35.340 ;
        RECT 86.830 34.570 87.200 61.480 ;
        RECT 87.620 58.030 88.080 58.460 ;
        RECT 86.800 34.110 87.250 34.570 ;
        RECT 86.830 34.070 87.200 34.110 ;
        RECT 87.640 33.980 88.010 58.030 ;
        RECT 88.390 53.320 88.840 53.750 ;
        RECT 77.250 33.550 78.920 33.560 ;
        RECT 76.770 33.310 76.990 33.420 ;
        RECT 76.400 32.500 76.600 32.520 ;
        RECT 75.260 31.960 75.580 32.280 ;
        RECT 76.380 32.260 76.610 32.500 ;
        RECT 76.400 32.210 76.610 32.260 ;
        RECT 76.770 32.210 76.960 33.310 ;
        RECT 77.210 33.280 78.920 33.550 ;
        RECT 87.610 33.520 88.050 33.980 ;
        RECT 87.640 33.470 88.010 33.520 ;
        RECT 77.210 33.140 77.370 33.280 ;
        RECT 77.210 32.860 77.540 33.140 ;
        RECT 77.210 32.550 77.370 32.860 ;
        RECT 74.360 31.210 74.630 31.870 ;
        RECT 72.050 29.250 72.440 31.110 ;
        RECT 70.440 28.260 70.700 28.580 ;
        RECT 70.450 27.620 70.690 28.260 ;
        RECT 70.450 26.760 70.720 27.620 ;
        RECT 72.060 26.760 72.440 29.250 ;
        RECT 74.380 28.620 74.620 31.210 ;
        RECT 75.260 30.970 75.580 31.290 ;
        RECT 76.400 31.040 76.560 32.210 ;
        RECT 76.790 32.090 76.960 32.210 ;
        RECT 76.800 31.160 76.960 32.090 ;
        RECT 77.100 32.000 77.370 32.550 ;
        RECT 77.100 31.950 77.380 32.000 ;
        RECT 77.210 31.860 77.380 31.950 ;
        RECT 77.210 31.390 77.370 31.860 ;
        RECT 88.410 31.630 88.780 53.320 ;
        RECT 94.960 52.270 95.540 52.830 ;
        RECT 91.750 50.700 92.310 51.350 ;
        RECT 92.700 51.190 93.260 51.770 ;
        RECT 93.780 51.650 94.340 52.240 ;
        RECT 89.280 48.240 89.710 48.680 ;
        RECT 88.380 31.620 88.780 31.630 ;
        RECT 77.210 31.300 77.380 31.390 ;
        RECT 76.790 31.040 76.960 31.160 ;
        RECT 76.400 30.990 76.610 31.040 ;
        RECT 76.380 30.750 76.610 30.990 ;
        RECT 75.260 30.420 75.580 30.740 ;
        RECT 76.400 30.730 76.600 30.750 ;
        RECT 76.400 30.100 76.560 30.730 ;
        RECT 76.770 30.120 76.960 31.040 ;
        RECT 77.100 31.250 77.380 31.300 ;
        RECT 77.100 30.700 77.370 31.250 ;
        RECT 88.370 31.200 88.790 31.620 ;
        RECT 88.410 31.190 88.780 31.200 ;
        RECT 76.750 30.100 76.990 30.120 ;
        RECT 76.400 29.910 76.990 30.100 ;
        RECT 75.260 29.270 75.580 29.590 ;
        RECT 76.400 29.280 76.560 29.910 ;
        RECT 76.750 29.890 76.990 29.910 ;
        RECT 76.400 29.260 76.600 29.280 ;
        RECT 75.260 28.720 75.580 29.040 ;
        RECT 76.380 29.020 76.610 29.260 ;
        RECT 76.400 28.970 76.610 29.020 ;
        RECT 76.770 28.970 76.960 29.890 ;
        RECT 77.210 29.310 77.370 30.700 ;
        RECT 74.370 28.300 74.630 28.620 ;
        RECT 74.380 26.760 74.620 28.300 ;
        RECT 75.260 27.740 75.580 28.060 ;
        RECT 76.400 27.810 76.560 28.970 ;
        RECT 76.790 28.850 76.960 28.970 ;
        RECT 76.800 27.930 76.960 28.850 ;
        RECT 77.100 28.760 77.370 29.310 ;
        RECT 77.100 28.710 77.380 28.760 ;
        RECT 77.210 28.620 77.380 28.710 ;
        RECT 77.210 28.160 77.370 28.620 ;
        RECT 77.210 28.070 77.380 28.160 ;
        RECT 76.790 27.810 76.960 27.930 ;
        RECT 76.400 27.760 76.610 27.810 ;
        RECT 76.380 27.520 76.610 27.760 ;
        RECT 75.260 27.190 75.580 27.510 ;
        RECT 76.400 27.500 76.600 27.520 ;
        RECT 76.400 26.770 76.560 27.500 ;
        RECT 76.770 26.820 76.960 27.810 ;
        RECT 77.100 28.020 77.380 28.070 ;
        RECT 77.100 27.470 77.370 28.020 ;
        RECT 77.210 26.770 77.370 27.470 ;
        RECT 45.130 23.780 45.410 24.110 ;
        RECT 41.630 23.410 41.910 23.650 ;
        RECT 40.890 22.140 41.300 22.470 ;
        RECT 40.890 20.390 41.300 20.720 ;
        RECT 40.890 18.640 41.300 18.970 ;
        RECT 41.630 17.650 41.870 23.410 ;
        RECT 44.570 23.380 44.920 23.650 ;
        RECT 48.900 23.650 49.230 24.400 ;
        RECT 50.400 23.940 50.590 26.720 ;
        RECT 51.710 26.430 51.940 26.720 ;
        RECT 51.620 25.950 51.950 26.430 ;
        RECT 51.710 23.940 51.940 25.950 ;
        RECT 54.680 23.940 54.930 26.720 ;
        RECT 50.400 23.720 50.600 23.940 ;
        RECT 43.050 23.360 43.250 23.380 ;
        RECT 43.050 23.070 43.400 23.360 ;
        RECT 43.050 21.610 43.250 21.630 ;
        RECT 43.050 21.320 43.400 21.610 ;
        RECT 43.050 19.860 43.250 19.880 ;
        RECT 43.050 19.570 43.400 19.860 ;
        RECT 43.050 18.110 43.250 18.130 ;
        RECT 43.050 17.820 43.400 18.110 ;
        RECT 44.570 17.720 44.880 23.380 ;
        RECT 46.810 23.350 47.100 23.360 ;
        RECT 46.790 23.080 47.110 23.350 ;
        RECT 46.790 23.070 47.100 23.080 ;
        RECT 47.830 23.010 48.150 23.310 ;
        RECT 45.130 22.030 45.410 22.360 ;
        RECT 46.810 21.600 47.100 21.610 ;
        RECT 46.790 21.330 47.110 21.600 ;
        RECT 46.790 21.320 47.100 21.330 ;
        RECT 47.830 21.260 48.150 21.560 ;
        RECT 45.130 20.280 45.410 20.610 ;
        RECT 46.810 19.850 47.100 19.860 ;
        RECT 46.790 19.580 47.110 19.850 ;
        RECT 46.790 19.570 47.100 19.580 ;
        RECT 47.830 19.510 48.150 19.810 ;
        RECT 45.130 18.530 45.410 18.860 ;
        RECT 46.810 18.100 47.100 18.110 ;
        RECT 46.790 17.830 47.110 18.100 ;
        RECT 46.790 17.820 47.100 17.830 ;
        RECT 47.830 17.760 48.150 18.060 ;
        RECT 41.570 17.400 41.870 17.650 ;
        RECT 44.510 17.400 44.880 17.720 ;
        RECT 48.900 17.700 49.190 23.650 ;
        RECT 50.130 23.230 50.600 23.720 ;
        RECT 50.990 23.580 51.360 23.600 ;
        RECT 50.940 23.320 51.360 23.580 ;
        RECT 51.710 23.340 51.950 23.940 ;
        RECT 54.680 23.720 54.940 23.940 ;
        RECT 60.750 23.930 60.990 26.760 ;
        RECT 53.450 23.560 53.790 23.610 ;
        RECT 53.450 23.540 54.010 23.560 ;
        RECT 54.680 23.550 55.330 23.720 ;
        RECT 53.330 23.370 54.010 23.540 ;
        RECT 50.990 23.310 51.360 23.320 ;
        RECT 49.950 22.790 50.270 23.070 ;
        RECT 50.410 22.970 50.600 23.230 ;
        RECT 50.410 22.680 50.640 22.970 ;
        RECT 50.410 21.910 50.600 22.680 ;
        RECT 49.950 21.520 50.270 21.800 ;
        RECT 50.410 21.620 50.640 21.910 ;
        RECT 50.410 21.360 50.600 21.620 ;
        RECT 50.130 20.870 50.600 21.360 ;
        RECT 50.990 21.270 51.360 21.280 ;
        RECT 50.940 21.010 51.360 21.270 ;
        RECT 50.990 20.990 51.360 21.010 ;
        RECT 50.410 20.520 50.600 20.870 ;
        RECT 50.130 20.030 50.600 20.520 ;
        RECT 50.990 20.380 51.360 20.400 ;
        RECT 50.940 20.120 51.360 20.380 ;
        RECT 50.990 20.110 51.360 20.120 ;
        RECT 49.950 19.590 50.270 19.870 ;
        RECT 50.410 19.770 50.600 20.030 ;
        RECT 50.410 19.480 50.640 19.770 ;
        RECT 50.410 18.710 50.600 19.480 ;
        RECT 49.950 18.320 50.270 18.600 ;
        RECT 50.410 18.420 50.640 18.710 ;
        RECT 50.410 18.160 50.600 18.420 ;
        RECT 48.900 17.400 49.230 17.700 ;
        RECT 50.130 17.670 50.600 18.160 ;
        RECT 50.990 18.070 51.360 18.080 ;
        RECT 50.940 17.810 51.360 18.070 ;
        RECT 50.990 17.790 51.360 17.810 ;
        RECT 50.400 17.450 50.600 17.670 ;
        RECT 51.720 17.450 51.950 23.340 ;
        RECT 53.450 23.330 54.010 23.370 ;
        RECT 53.450 23.290 53.790 23.330 ;
        RECT 54.690 22.650 55.330 23.550 ;
        RECT 58.410 22.880 58.600 23.870 ;
        RECT 58.810 23.190 58.970 23.920 ;
        RECT 60.750 23.900 61.120 23.930 ;
        RECT 60.730 23.650 61.120 23.900 ;
        RECT 58.770 23.170 58.970 23.190 ;
        RECT 59.790 23.180 60.110 23.500 ;
        RECT 58.760 22.930 58.990 23.170 ;
        RECT 60.430 23.080 60.690 23.400 ;
        RECT 58.760 22.880 58.970 22.930 ;
        RECT 58.410 22.760 58.580 22.880 ;
        RECT 54.690 21.940 54.940 22.650 ;
        RECT 56.030 22.220 56.350 22.560 ;
        RECT 53.450 21.260 53.790 21.300 ;
        RECT 53.450 21.220 54.010 21.260 ;
        RECT 53.330 21.050 54.010 21.220 ;
        RECT 53.450 21.030 54.010 21.050 ;
        RECT 53.450 20.980 53.790 21.030 ;
        RECT 54.690 20.870 55.330 21.940 ;
        RECT 54.690 20.520 54.940 20.870 ;
        RECT 53.450 20.360 53.790 20.410 ;
        RECT 53.450 20.340 54.010 20.360 ;
        RECT 53.330 20.170 54.010 20.340 ;
        RECT 53.450 20.130 54.010 20.170 ;
        RECT 53.450 20.090 53.790 20.130 ;
        RECT 54.690 19.450 55.330 20.520 ;
        RECT 54.690 18.740 54.940 19.450 ;
        RECT 53.450 18.060 53.790 18.100 ;
        RECT 53.450 18.020 54.010 18.060 ;
        RECT 53.330 17.850 54.010 18.020 ;
        RECT 53.450 17.830 54.010 17.850 ;
        RECT 53.450 17.780 53.790 17.830 ;
        RECT 54.690 17.770 55.330 18.740 ;
        RECT 54.680 17.670 55.330 17.770 ;
        RECT 54.680 17.450 54.940 17.670 ;
        RECT 56.110 17.460 56.320 22.220 ;
        RECT 58.410 21.850 58.570 22.760 ;
        RECT 57.140 21.730 57.400 21.850 ;
        RECT 57.130 21.530 57.400 21.730 ;
        RECT 58.410 21.730 58.580 21.850 ;
        RECT 58.810 21.730 58.970 22.880 ;
        RECT 59.790 22.630 60.110 22.950 ;
        RECT 60.430 22.350 60.640 23.080 ;
        RECT 60.410 22.030 60.670 22.350 ;
        RECT 57.130 20.840 57.340 21.530 ;
        RECT 57.120 20.780 57.380 20.840 ;
        RECT 58.410 20.810 58.600 21.730 ;
        RECT 58.760 21.680 58.970 21.730 ;
        RECT 58.760 21.440 58.990 21.680 ;
        RECT 59.790 21.660 60.110 21.980 ;
        RECT 58.770 21.420 58.970 21.440 ;
        RECT 58.380 20.780 58.620 20.810 ;
        RECT 58.810 20.780 58.970 21.420 ;
        RECT 59.790 21.110 60.110 21.430 ;
        RECT 57.120 20.530 57.760 20.780 ;
        RECT 58.380 20.610 58.970 20.780 ;
        RECT 58.380 20.580 58.620 20.610 ;
        RECT 57.120 20.520 57.380 20.530 ;
        RECT 56.650 19.430 56.990 19.770 ;
        RECT 56.690 19.410 56.910 19.430 ;
        RECT 41.570 5.020 41.810 17.400 ;
        RECT 44.510 16.570 44.820 17.400 ;
        RECT 48.940 17.080 49.230 17.400 ;
        RECT 49.440 17.100 49.780 17.420 ;
        RECT 48.910 16.730 49.260 17.080 ;
        RECT 44.470 16.240 44.840 16.570 ;
        RECT 48.940 16.270 49.230 16.730 ;
        RECT 49.440 16.490 49.690 17.100 ;
        RECT 50.400 16.510 50.590 17.450 ;
        RECT 54.680 17.040 54.930 17.450 ;
        RECT 56.080 17.140 56.360 17.460 ;
        RECT 56.690 17.130 56.890 19.410 ;
        RECT 57.040 18.480 57.360 18.800 ;
        RECT 57.150 17.840 57.340 17.950 ;
        RECT 57.090 17.520 57.410 17.840 ;
        RECT 54.650 16.750 54.990 17.040 ;
        RECT 56.650 16.810 56.930 17.130 ;
        RECT 57.110 17.120 57.390 17.520 ;
        RECT 44.510 15.030 44.820 16.240 ;
        RECT 48.370 15.990 49.230 16.270 ;
        RECT 48.290 15.980 49.230 15.990 ;
        RECT 49.390 16.380 49.690 16.490 ;
        RECT 48.290 15.510 48.750 15.980 ;
        RECT 44.460 14.550 44.880 15.030 ;
        RECT 49.390 14.870 49.580 16.380 ;
        RECT 50.340 16.190 50.660 16.510 ;
        RECT 57.580 15.900 57.760 20.530 ;
        RECT 58.410 19.640 58.600 20.580 ;
        RECT 58.810 19.950 58.970 20.610 ;
        RECT 58.770 19.930 58.970 19.950 ;
        RECT 59.790 19.940 60.110 20.260 ;
        RECT 60.410 20.150 60.670 20.470 ;
        RECT 58.760 19.690 58.990 19.930 ;
        RECT 58.760 19.640 58.970 19.690 ;
        RECT 58.410 19.520 58.580 19.640 ;
        RECT 58.410 18.600 58.570 19.520 ;
        RECT 58.410 18.480 58.580 18.600 ;
        RECT 58.810 18.480 58.970 19.640 ;
        RECT 59.790 19.390 60.110 19.710 ;
        RECT 60.410 19.290 60.570 20.150 ;
        RECT 60.280 18.970 60.570 19.290 ;
        RECT 60.870 19.220 61.120 23.650 ;
        RECT 62.930 21.740 63.310 26.760 ;
        RECT 64.680 23.930 64.920 26.760 ;
        RECT 64.680 23.610 65.150 23.930 ;
        RECT 62.930 19.880 63.320 21.740 ;
        RECT 60.850 19.190 61.130 19.220 ;
        RECT 60.840 18.910 61.140 19.190 ;
        RECT 60.850 18.890 61.130 18.910 ;
        RECT 58.410 17.490 58.600 18.480 ;
        RECT 58.760 18.430 58.970 18.480 ;
        RECT 58.760 18.190 58.990 18.430 ;
        RECT 59.790 18.410 60.110 18.730 ;
        RECT 58.770 18.170 58.970 18.190 ;
        RECT 58.810 17.440 58.970 18.170 ;
        RECT 59.790 17.860 60.110 18.180 ;
        RECT 58.900 17.060 59.160 17.090 ;
        RECT 58.880 16.760 59.180 17.060 ;
        RECT 58.900 16.750 59.160 16.760 ;
        RECT 49.750 15.520 50.070 15.840 ;
        RECT 50.840 15.520 51.160 15.840 ;
        RECT 51.940 15.510 52.260 15.830 ;
        RECT 54.780 15.510 55.100 15.830 ;
        RECT 55.880 15.520 56.200 15.840 ;
        RECT 56.970 15.520 57.290 15.840 ;
        RECT 57.580 15.600 58.060 15.900 ;
        RECT 58.910 15.830 59.130 16.750 ;
        RECT 60.870 16.620 61.120 18.890 ;
        RECT 62.930 17.430 63.310 19.880 ;
        RECT 64.880 19.190 65.150 23.610 ;
        RECT 64.860 18.880 65.170 19.190 ;
        RECT 64.880 16.640 65.150 18.880 ;
        RECT 66.960 17.430 67.360 26.760 ;
        RECT 70.480 25.110 70.720 26.760 ;
        RECT 89.290 26.450 89.660 48.240 ;
        RECT 89.250 25.940 89.740 26.450 ;
        RECT 89.290 25.910 89.660 25.940 ;
        RECT 70.480 24.870 71.060 25.110 ;
        RECT 68.480 22.880 68.800 23.200 ;
        RECT 68.630 22.200 68.950 22.520 ;
        RECT 68.630 21.310 68.950 21.630 ;
        RECT 68.480 20.630 68.800 20.950 ;
        RECT 68.480 20.110 68.800 20.430 ;
        RECT 68.630 19.430 68.950 19.750 ;
        RECT 68.630 18.540 68.950 18.860 ;
        RECT 68.480 17.860 68.800 18.180 ;
        RECT 69.560 17.610 69.790 23.660 ;
        RECT 70.820 23.530 71.060 24.870 ;
        RECT 70.820 19.310 71.050 23.530 ;
        RECT 75.940 22.470 76.200 22.530 ;
        RECT 75.930 22.210 76.200 22.470 ;
        RECT 75.420 21.280 75.680 21.600 ;
        RECT 74.950 19.440 75.210 19.760 ;
        RECT 70.780 19.300 71.060 19.310 ;
        RECT 70.780 18.980 71.080 19.300 ;
        RECT 67.700 17.070 68.130 17.470 ;
        RECT 60.860 16.360 61.180 16.620 ;
        RECT 64.880 16.330 65.230 16.640 ;
        RECT 57.660 15.490 58.060 15.600 ;
        RECT 58.850 15.430 59.190 15.830 ;
        RECT 59.560 15.550 59.880 15.870 ;
        RECT 60.650 15.550 60.970 15.870 ;
        RECT 61.750 15.540 62.070 15.860 ;
        RECT 64.590 15.540 64.910 15.860 ;
        RECT 65.690 15.550 66.010 15.870 ;
        RECT 66.780 15.550 67.100 15.870 ;
        RECT 58.910 15.350 59.130 15.430 ;
        RECT 67.740 15.280 68.090 17.070 ;
        RECT 69.560 16.510 69.780 17.610 ;
        RECT 70.820 17.110 71.050 18.980 ;
        RECT 74.450 18.510 74.710 18.830 ;
        RECT 70.820 16.880 74.030 17.110 ;
        RECT 70.820 16.870 71.050 16.880 ;
        RECT 69.270 16.270 69.780 16.510 ;
        RECT 48.950 14.550 49.580 14.870 ;
        RECT 50.300 14.840 50.620 15.160 ;
        RECT 51.390 14.820 51.710 15.140 ;
        RECT 55.330 14.820 55.650 15.140 ;
        RECT 56.420 14.840 56.740 15.160 ;
        RECT 60.110 14.870 60.430 15.190 ;
        RECT 61.200 14.850 61.520 15.170 ;
        RECT 65.140 14.850 65.460 15.170 ;
        RECT 66.230 14.870 66.550 15.190 ;
        RECT 69.270 15.020 69.500 16.270 ;
        RECT 73.800 15.910 74.030 16.880 ;
        RECT 70.330 15.530 70.650 15.850 ;
        RECT 71.430 15.540 71.750 15.860 ;
        RECT 72.520 15.540 72.840 15.860 ;
        RECT 73.750 15.510 74.060 15.910 ;
        RECT 69.160 14.580 69.620 15.020 ;
        RECT 69.770 14.830 70.090 15.150 ;
        RECT 70.880 14.840 71.200 15.160 ;
        RECT 71.970 14.860 72.290 15.180 ;
        RECT 48.950 14.450 49.390 14.550 ;
        RECT 50.300 13.470 50.620 13.790 ;
        RECT 51.390 13.470 51.710 13.790 ;
        RECT 55.330 13.470 55.650 13.790 ;
        RECT 56.420 13.470 56.740 13.790 ;
        RECT 60.110 13.500 60.430 13.820 ;
        RECT 61.200 13.500 61.520 13.820 ;
        RECT 65.140 13.500 65.460 13.820 ;
        RECT 66.230 13.500 66.550 13.820 ;
        RECT 69.780 13.490 70.100 13.810 ;
        RECT 70.880 13.490 71.200 13.810 ;
        RECT 71.970 13.490 72.290 13.810 ;
        RECT 49.740 12.740 50.060 13.060 ;
        RECT 50.840 12.740 51.160 13.060 ;
        RECT 51.940 12.740 52.260 13.060 ;
        RECT 54.780 12.740 55.100 13.060 ;
        RECT 55.880 12.740 56.200 13.060 ;
        RECT 56.980 12.740 57.300 13.060 ;
        RECT 59.550 12.770 59.870 13.090 ;
        RECT 60.650 12.770 60.970 13.090 ;
        RECT 61.750 12.770 62.070 13.090 ;
        RECT 64.590 12.770 64.910 13.090 ;
        RECT 65.690 12.770 66.010 13.090 ;
        RECT 66.790 12.770 67.110 13.090 ;
        RECT 70.330 12.760 70.650 13.080 ;
        RECT 71.430 12.760 71.750 13.080 ;
        RECT 72.530 12.760 72.850 13.080 ;
        RECT 73.260 12.730 73.530 12.760 ;
        RECT 73.250 12.200 73.530 12.730 ;
        RECT 73.800 12.340 74.030 15.510 ;
        RECT 73.670 12.200 74.030 12.340 ;
        RECT 73.250 11.900 74.030 12.200 ;
        RECT 73.240 11.890 74.030 11.900 ;
        RECT 73.240 11.880 74.010 11.890 ;
        RECT 49.740 11.370 50.060 11.690 ;
        RECT 50.840 11.370 51.160 11.690 ;
        RECT 51.940 11.370 52.260 11.690 ;
        RECT 54.780 11.370 55.100 11.690 ;
        RECT 55.880 11.370 56.200 11.690 ;
        RECT 56.980 11.370 57.300 11.690 ;
        RECT 59.550 11.400 59.870 11.720 ;
        RECT 60.650 11.400 60.970 11.720 ;
        RECT 61.750 11.400 62.070 11.720 ;
        RECT 64.590 11.400 64.910 11.720 ;
        RECT 65.690 11.400 66.010 11.720 ;
        RECT 66.790 11.400 67.110 11.720 ;
        RECT 70.330 11.390 70.650 11.710 ;
        RECT 71.430 11.390 71.750 11.710 ;
        RECT 72.530 11.390 72.850 11.710 ;
        RECT 73.240 11.450 73.530 11.880 ;
        RECT 49.170 11.020 49.490 11.050 ;
        RECT 57.550 11.040 57.870 11.050 ;
        RECT 49.160 10.730 49.490 11.020 ;
        RECT 49.160 10.580 49.480 10.730 ;
        RECT 50.300 10.690 50.620 11.010 ;
        RECT 51.390 10.690 51.710 11.010 ;
        RECT 55.330 10.690 55.650 11.010 ;
        RECT 56.420 10.690 56.740 11.010 ;
        RECT 49.160 10.260 49.500 10.580 ;
        RECT 49.160 9.270 49.480 10.260 ;
        RECT 49.040 8.670 49.580 9.270 ;
        RECT 57.530 8.250 57.870 11.040 ;
        RECT 58.980 11.030 59.300 11.080 ;
        RECT 58.960 10.610 59.300 11.030 ;
        RECT 60.110 10.720 60.430 11.040 ;
        RECT 61.200 10.720 61.520 11.040 ;
        RECT 65.140 10.720 65.460 11.040 ;
        RECT 66.230 10.720 66.550 11.040 ;
        RECT 67.360 10.760 67.680 11.080 ;
        RECT 67.380 10.610 67.650 10.760 ;
        RECT 69.780 10.720 70.100 11.040 ;
        RECT 70.880 10.710 71.200 11.030 ;
        RECT 71.970 10.710 72.290 11.030 ;
        RECT 73.100 10.750 73.420 11.070 ;
        RECT 74.450 10.670 74.700 18.510 ;
        RECT 74.950 11.570 75.200 19.440 ;
        RECT 75.430 12.480 75.680 21.280 ;
        RECT 75.930 13.370 76.180 22.210 ;
        RECT 91.770 14.870 92.270 50.700 ;
        RECT 92.700 20.150 93.200 51.190 ;
        RECT 93.830 25.380 94.330 51.650 ;
        RECT 94.960 30.550 95.460 52.270 ;
        RECT 103.820 50.670 105.100 62.870 ;
        RECT 103.810 49.330 105.100 50.670 ;
        RECT 103.820 48.840 105.100 49.330 ;
        RECT 108.180 47.660 108.380 47.690 ;
        RECT 108.090 47.160 108.400 47.660 ;
        RECT 104.270 45.890 104.620 46.370 ;
        RECT 100.280 42.690 100.750 43.180 ;
        RECT 94.910 29.990 95.460 30.550 ;
        RECT 93.820 24.820 94.340 25.380 ;
        RECT 92.690 19.630 93.210 20.150 ;
        RECT 91.610 14.300 92.270 14.870 ;
        RECT 75.880 12.790 76.250 13.370 ;
        RECT 75.350 11.900 75.720 12.480 ;
        RECT 74.860 10.990 75.230 11.570 ;
        RECT 58.960 10.290 59.310 10.610 ;
        RECT 67.350 10.290 67.670 10.610 ;
        RECT 73.090 10.450 73.410 10.600 ;
        RECT 57.470 7.730 57.930 8.250 ;
        RECT 58.960 7.360 59.300 10.290 ;
        RECT 58.870 6.840 59.390 7.360 ;
        RECT 67.380 6.480 67.650 10.290 ;
        RECT 73.090 10.280 73.450 10.450 ;
        RECT 67.270 5.920 67.760 6.480 ;
        RECT 41.170 3.700 41.820 5.020 ;
        RECT 73.120 0.460 73.450 10.280 ;
        RECT 74.390 10.100 74.740 10.670 ;
        RECT 91.770 5.990 92.270 14.300 ;
        RECT 92.700 6.900 93.200 19.630 ;
        RECT 93.830 7.770 94.330 24.820 ;
        RECT 94.960 9.280 95.460 29.990 ;
        RECT 97.850 16.840 98.430 17.400 ;
        RECT 97.880 16.830 98.390 16.840 ;
        RECT 94.960 8.720 95.520 9.280 ;
        RECT 94.960 8.590 95.460 8.720 ;
        RECT 97.880 4.960 98.380 16.830 ;
        RECT 97.250 3.680 98.380 4.960 ;
        RECT 73.060 0.070 73.490 0.460 ;
        RECT 39.520 -0.590 39.890 -0.210 ;
        RECT 100.330 -0.660 100.730 42.690 ;
        RECT 101.250 42.080 101.670 42.440 ;
        RECT 38.870 -1.210 39.260 -0.820 ;
        RECT 100.320 -1.120 100.790 -0.660 ;
        RECT 38.270 -1.840 38.650 -1.450 ;
        RECT 101.260 -1.460 101.650 42.080 ;
        RECT 102.170 39.690 102.620 40.120 ;
        RECT 101.230 -1.930 101.690 -1.460 ;
        RECT 37.680 -2.470 38.030 -2.100 ;
        RECT 102.190 -2.280 102.580 39.690 ;
        RECT 103.030 39.430 103.410 39.440 ;
        RECT 103.010 39.130 103.430 39.430 ;
        RECT 102.170 -2.740 102.640 -2.280 ;
        RECT 37.040 -3.150 37.400 -2.770 ;
        RECT 103.030 -3.080 103.410 39.130 ;
        RECT 104.370 15.900 104.600 45.890 ;
        RECT 108.180 43.320 108.380 47.160 ;
        RECT 109.080 43.760 109.400 44.080 ;
        RECT 110.080 43.640 110.310 43.930 ;
        RECT 110.650 43.760 110.970 44.080 ;
        RECT 111.210 43.650 111.440 43.940 ;
        RECT 107.670 43.100 107.900 43.290 ;
        RECT 107.670 43.000 108.020 43.100 ;
        RECT 108.170 43.030 108.400 43.320 ;
        RECT 110.100 43.170 110.290 43.640 ;
        RECT 107.680 42.780 108.020 43.000 ;
        RECT 107.680 42.270 108.020 42.490 ;
        RECT 107.670 42.170 108.020 42.270 ;
        RECT 108.180 42.240 108.380 43.030 ;
        RECT 110.030 42.850 110.290 43.170 ;
        RECT 111.210 43.160 111.400 43.650 ;
        RECT 111.690 43.320 111.880 64.190 ;
        RECT 115.030 55.340 115.850 55.430 ;
        RECT 114.970 54.650 115.850 55.340 ;
        RECT 111.030 42.910 111.400 43.160 ;
        RECT 111.670 43.030 111.900 43.320 ;
        RECT 111.030 42.840 111.300 42.910 ;
        RECT 107.670 41.980 107.900 42.170 ;
        RECT 108.170 41.950 108.400 42.240 ;
        RECT 110.030 42.100 110.290 42.420 ;
        RECT 111.030 42.360 111.300 42.430 ;
        RECT 111.030 42.110 111.400 42.360 ;
        RECT 111.690 42.240 111.880 43.030 ;
        RECT 108.180 40.120 108.380 41.950 ;
        RECT 110.100 41.630 110.290 42.100 ;
        RECT 109.080 41.190 109.400 41.510 ;
        RECT 110.080 41.340 110.310 41.630 ;
        RECT 111.210 41.620 111.400 42.110 ;
        RECT 111.670 41.950 111.900 42.240 ;
        RECT 110.650 41.190 110.970 41.510 ;
        RECT 111.210 41.330 111.440 41.620 ;
        RECT 109.080 40.560 109.400 40.880 ;
        RECT 110.080 40.440 110.310 40.730 ;
        RECT 110.650 40.560 110.970 40.880 ;
        RECT 111.210 40.450 111.440 40.740 ;
        RECT 107.670 39.900 107.900 40.090 ;
        RECT 107.670 39.800 108.020 39.900 ;
        RECT 108.170 39.830 108.400 40.120 ;
        RECT 110.100 39.970 110.290 40.440 ;
        RECT 107.680 39.580 108.020 39.800 ;
        RECT 107.680 39.070 108.020 39.290 ;
        RECT 107.670 38.970 108.020 39.070 ;
        RECT 108.180 39.040 108.380 39.830 ;
        RECT 110.030 39.650 110.290 39.970 ;
        RECT 111.210 39.960 111.400 40.450 ;
        RECT 111.690 40.120 111.880 41.950 ;
        RECT 111.030 39.710 111.400 39.960 ;
        RECT 111.670 39.830 111.900 40.120 ;
        RECT 111.030 39.640 111.300 39.710 ;
        RECT 107.670 38.780 107.900 38.970 ;
        RECT 108.170 38.750 108.400 39.040 ;
        RECT 110.030 38.900 110.290 39.220 ;
        RECT 111.030 39.160 111.300 39.230 ;
        RECT 111.030 38.910 111.400 39.160 ;
        RECT 111.690 39.040 111.880 39.830 ;
        RECT 108.180 37.830 108.380 38.750 ;
        RECT 110.100 38.430 110.290 38.900 ;
        RECT 109.080 37.990 109.400 38.310 ;
        RECT 110.080 38.140 110.310 38.430 ;
        RECT 111.210 38.420 111.400 38.910 ;
        RECT 111.670 38.750 111.900 39.040 ;
        RECT 110.650 37.990 110.970 38.310 ;
        RECT 111.210 38.130 111.440 38.420 ;
        RECT 111.690 37.830 111.880 38.750 ;
        RECT 114.970 35.650 115.680 54.650 ;
        RECT 114.840 34.860 115.680 35.650 ;
        RECT 110.560 16.820 111.280 17.390 ;
        RECT 104.370 15.670 104.610 15.900 ;
        RECT 104.370 8.020 104.600 15.670 ;
        RECT 110.620 9.810 111.130 16.820 ;
        RECT 110.480 9.760 111.130 9.810 ;
        RECT 110.470 9.580 111.130 9.760 ;
        RECT 110.440 9.570 111.130 9.580 ;
        RECT 110.440 9.200 111.040 9.570 ;
        RECT 104.360 7.790 104.650 8.020 ;
        RECT 104.370 6.410 104.600 7.790 ;
        RECT 110.440 7.330 111.020 9.200 ;
        RECT 109.870 7.010 111.020 7.330 ;
        RECT 110.090 6.660 111.020 7.010 ;
        RECT 104.360 6.180 104.650 6.410 ;
        RECT 109.870 6.340 111.020 6.660 ;
        RECT 104.370 4.810 104.600 6.180 ;
        RECT 110.440 5.560 111.020 6.340 ;
        RECT 110.030 5.370 110.350 5.420 ;
        RECT 109.800 5.140 110.350 5.370 ;
        RECT 110.030 5.100 110.350 5.140 ;
        RECT 110.490 4.960 111.020 5.560 ;
        RECT 110.450 4.950 111.020 4.960 ;
        RECT 104.360 4.580 104.650 4.810 ;
        RECT 104.370 3.190 104.600 4.580 ;
        RECT 110.440 3.950 111.020 4.950 ;
        RECT 110.030 3.760 110.350 3.810 ;
        RECT 106.080 3.670 108.090 3.700 ;
        RECT 105.590 3.500 108.090 3.670 ;
        RECT 109.800 3.530 110.350 3.760 ;
        RECT 105.590 3.450 106.100 3.500 ;
        RECT 105.590 3.440 105.880 3.450 ;
        RECT 104.360 2.960 104.650 3.190 ;
        RECT 104.370 1.590 104.600 2.960 ;
        RECT 105.090 1.980 105.410 2.060 ;
        RECT 106.670 1.980 107.180 2.030 ;
        RECT 105.090 1.800 107.180 1.980 ;
        RECT 104.360 1.360 104.650 1.590 ;
        RECT 104.370 -0.030 104.600 1.360 ;
        RECT 107.920 0.450 108.090 3.500 ;
        RECT 110.030 3.490 110.350 3.530 ;
        RECT 110.490 3.350 111.020 3.950 ;
        RECT 110.440 2.340 111.020 3.350 ;
        RECT 110.020 2.150 110.340 2.200 ;
        RECT 109.790 1.920 110.340 2.150 ;
        RECT 110.020 1.880 110.340 1.920 ;
        RECT 110.480 1.740 111.020 2.340 ;
        RECT 110.440 0.720 111.020 1.740 ;
        RECT 110.030 0.530 110.350 0.580 ;
        RECT 107.500 0.250 108.090 0.450 ;
        RECT 109.800 0.300 110.350 0.530 ;
        RECT 110.030 0.260 110.350 0.300 ;
        RECT 107.500 0.230 108.010 0.250 ;
        RECT 107.500 0.220 107.790 0.230 ;
        RECT 110.490 0.120 111.020 0.720 ;
        RECT 104.360 -0.260 104.650 -0.030 ;
        RECT 104.370 -1.630 104.600 -0.260 ;
        RECT 110.440 -0.890 111.020 0.120 ;
        RECT 110.020 -1.080 110.340 -1.030 ;
        RECT 109.790 -1.310 110.340 -1.080 ;
        RECT 110.020 -1.350 110.340 -1.310 ;
        RECT 110.480 -1.490 111.020 -0.890 ;
        RECT 104.360 -1.860 104.650 -1.630 ;
        RECT 36.450 -3.390 36.790 -3.380 ;
        RECT 36.430 -3.760 36.810 -3.390 ;
        RECT 103.000 -3.540 103.440 -3.080 ;
        RECT 104.370 -3.250 104.600 -1.860 ;
        RECT 109.610 -3.000 109.930 -2.680 ;
        RECT 109.660 -3.230 109.890 -3.000 ;
        RECT 104.360 -3.480 104.650 -3.250 ;
        RECT 110.440 -3.360 111.020 -1.490 ;
        RECT 36.450 -3.770 36.780 -3.760 ;
        RECT 110.020 -4.280 110.340 -4.230 ;
        RECT 109.790 -4.510 110.340 -4.280 ;
        RECT 110.020 -4.550 110.340 -4.510 ;
        RECT 34.670 -5.610 35.020 -5.280 ;
        RECT 110.480 -5.570 111.020 -3.360 ;
        RECT 34.690 -5.670 35.020 -5.610 ;
        RECT 106.780 -5.990 107.100 -5.940 ;
        RECT 107.720 -5.990 108.040 -5.940 ;
        RECT 106.550 -6.220 107.100 -5.990 ;
        RECT 107.490 -6.220 108.040 -5.990 ;
        RECT 108.670 -6.010 108.990 -5.960 ;
        RECT 109.980 -5.990 110.300 -5.940 ;
        RECT 106.780 -6.260 107.100 -6.220 ;
        RECT 107.720 -6.260 108.040 -6.220 ;
        RECT 108.440 -6.240 108.990 -6.010 ;
        RECT 109.750 -6.220 110.300 -5.990 ;
        RECT 108.670 -6.280 108.990 -6.240 ;
        RECT 109.980 -6.260 110.300 -6.220 ;
        RECT 33.400 -6.890 33.750 -6.560 ;
        RECT 33.400 -6.960 33.730 -6.890 ;
        RECT 31.260 -7.620 32.500 -7.290 ;
        RECT 32.790 -7.590 33.230 -7.170 ;
        RECT 31.260 -7.730 31.840 -7.620 ;
      LAYER via ;
        RECT 4.210 62.150 4.600 62.540 ;
        RECT 6.630 61.230 6.890 61.490 ;
        RECT 9.490 61.280 9.750 61.540 ;
        RECT 6.620 60.200 6.880 60.460 ;
        RECT 7.340 60.170 7.600 60.430 ;
        RECT 8.030 60.210 8.290 60.470 ;
        RECT 6.620 59.750 6.880 60.010 ;
        RECT 8.030 59.770 8.290 60.030 ;
        RECT 6.620 59.330 6.880 59.590 ;
        RECT 7.340 59.330 7.600 59.590 ;
        RECT 8.050 59.350 8.310 59.610 ;
        RECT 4.290 58.700 4.680 59.090 ;
        RECT 6.620 57.980 6.880 58.240 ;
        RECT 5.670 57.530 5.930 57.790 ;
        RECT 9.180 59.740 9.440 60.000 ;
        RECT 22.730 59.430 22.990 59.690 ;
        RECT 24.090 59.510 24.350 59.770 ;
        RECT 24.780 59.500 25.040 59.760 ;
        RECT 8.760 57.730 9.020 57.990 ;
        RECT 7.320 56.530 7.580 56.790 ;
        RECT 8.750 56.550 9.010 56.810 ;
        RECT 6.530 55.950 6.790 56.210 ;
        RECT 7.460 55.950 7.720 56.210 ;
        RECT 8.160 55.950 8.420 56.210 ;
        RECT 8.900 55.950 9.160 56.210 ;
        RECT 9.610 55.940 9.870 56.200 ;
        RECT 5.590 54.830 6.010 55.250 ;
        RECT 22.010 55.770 22.270 56.030 ;
        RECT 11.540 53.430 11.830 54.010 ;
        RECT 24.830 52.370 25.090 52.630 ;
        RECT 19.910 46.630 20.170 46.890 ;
        RECT 21.000 46.640 21.260 46.900 ;
        RECT 18.750 46.120 19.010 46.380 ;
        RECT 19.480 46.130 19.740 46.390 ;
        RECT 19.920 45.640 20.180 45.900 ;
        RECT 21.010 45.650 21.270 45.910 ;
        RECT 18.720 45.200 18.980 45.460 ;
        RECT 19.460 45.210 19.720 45.470 ;
        RECT 19.920 44.650 20.180 44.910 ;
        RECT 21.010 44.660 21.270 44.920 ;
        RECT 18.730 44.280 18.990 44.540 ;
        RECT 18.080 43.260 18.340 43.520 ;
        RECT 18.040 42.300 18.300 42.560 ;
        RECT 18.080 41.340 18.340 41.600 ;
        RECT 19.440 44.220 19.700 44.480 ;
        RECT 19.730 43.720 19.990 43.980 ;
        RECT 21.030 43.620 21.290 43.880 ;
        RECT 19.700 43.260 19.960 43.520 ;
        RECT 19.730 42.730 19.990 42.990 ;
        RECT 21.030 42.630 21.290 42.890 ;
        RECT 19.700 42.270 19.960 42.530 ;
        RECT 31.870 55.790 32.130 56.050 ;
        RECT 30.620 51.940 30.930 52.250 ;
        RECT 47.200 59.580 47.620 60.000 ;
        RECT 43.350 58.820 43.770 59.240 ;
        RECT 66.970 58.820 68.320 59.240 ;
        RECT 48.870 57.210 49.310 57.650 ;
        RECT 54.590 57.210 55.030 57.650 ;
        RECT 44.450 56.190 44.890 56.630 ;
        RECT 41.690 53.170 41.950 53.430 ;
        RECT 34.620 52.480 34.880 52.740 ;
        RECT 33.450 51.490 33.720 51.750 ;
        RECT 22.120 50.710 22.470 51.060 ;
        RECT 27.370 51.020 27.630 51.280 ;
        RECT 43.140 50.000 43.400 50.260 ;
        RECT 41.040 49.160 41.300 49.420 ;
        RECT 23.140 48.470 23.400 48.860 ;
        RECT 39.540 48.480 39.870 48.740 ;
        RECT 22.500 47.650 22.760 48.050 ;
        RECT 19.730 41.740 19.990 42.000 ;
        RECT 21.030 41.640 21.290 41.900 ;
        RECT 19.700 41.280 19.960 41.540 ;
        RECT 18.040 26.060 18.300 26.530 ;
        RECT 18.680 26.060 18.940 26.530 ;
        RECT 16.680 25.030 16.940 25.290 ;
        RECT 16.160 24.630 16.420 24.890 ;
        RECT 6.880 23.380 7.540 24.040 ;
        RECT 18.760 25.010 19.020 25.270 ;
        RECT 20.520 25.020 20.790 25.290 ;
        RECT 18.100 24.650 18.360 24.910 ;
        RECT 18.850 24.050 19.110 24.310 ;
        RECT 19.500 24.050 19.760 24.310 ;
        RECT 17.630 23.610 17.890 23.870 ;
        RECT 18.330 23.610 18.590 23.870 ;
        RECT 20.010 22.880 20.270 23.140 ;
        RECT 17.180 22.260 17.440 22.520 ;
        RECT 16.180 20.720 16.440 20.980 ;
        RECT 12.090 18.860 12.460 19.230 ;
        RECT 6.920 17.520 7.580 18.180 ;
        RECT 19.930 21.750 20.190 22.010 ;
        RECT 21.020 24.630 21.280 24.890 ;
        RECT 19.940 21.210 20.200 21.470 ;
        RECT 17.180 20.710 17.440 20.970 ;
        RECT 19.990 20.260 20.250 20.520 ;
        RECT 17.660 19.730 17.920 19.990 ;
        RECT 18.350 19.720 18.610 19.980 ;
        RECT 18.830 18.950 19.090 19.210 ;
        RECT 19.540 18.890 19.800 19.150 ;
        RECT 18.850 13.870 19.110 14.130 ;
        RECT 15.540 13.430 15.800 13.690 ;
        RECT 16.640 13.440 16.900 13.700 ;
        RECT 17.730 13.440 17.990 13.700 ;
        RECT 18.860 13.400 19.120 13.660 ;
        RECT 12.080 12.620 12.450 12.990 ;
        RECT 16.090 12.760 16.350 13.020 ;
        RECT 17.190 12.760 17.450 13.020 ;
        RECT 18.290 12.760 18.550 13.020 ;
        RECT 19.620 12.200 19.880 12.560 ;
        RECT 16.090 11.390 16.350 11.650 ;
        RECT 17.190 11.390 17.450 11.650 ;
        RECT 18.290 11.390 18.550 11.650 ;
        RECT 15.540 10.660 15.800 10.920 ;
        RECT 16.640 10.660 16.900 10.920 ;
        RECT 17.730 10.660 17.990 10.920 ;
        RECT 15.530 9.320 15.790 9.580 ;
        RECT 16.640 9.310 16.900 9.570 ;
        RECT 17.730 9.290 17.990 9.550 ;
        RECT 16.090 8.620 16.350 8.880 ;
        RECT 17.190 8.610 17.450 8.870 ;
        RECT 18.280 8.610 18.540 8.870 ;
        RECT 15.070 6.960 15.360 7.250 ;
        RECT 18.890 6.320 19.150 6.580 ;
        RECT 22.520 46.540 22.780 46.800 ;
        RECT 22.520 45.620 22.780 45.880 ;
        RECT 22.490 44.700 22.750 44.960 ;
        RECT 38.910 46.760 39.240 47.090 ;
        RECT 38.340 45.280 38.670 45.610 ;
        RECT 23.130 43.610 23.390 43.870 ;
        RECT 37.700 43.680 38.030 44.010 ;
        RECT 37.060 43.110 37.390 43.440 ;
        RECT 23.140 42.650 23.400 42.910 ;
        RECT 23.130 41.690 23.390 41.950 ;
        RECT 22.490 24.030 22.750 24.290 ;
        RECT 21.870 22.880 22.130 23.140 ;
        RECT 21.450 20.270 21.710 20.530 ;
        RECT 21.890 14.580 22.150 15.000 ;
        RECT 21.850 12.200 22.110 12.560 ;
        RECT 36.450 41.540 36.780 41.870 ;
        RECT 35.820 40.010 36.150 40.340 ;
        RECT 35.260 38.440 35.590 38.770 ;
        RECT 34.640 32.970 34.970 33.300 ;
        RECT 34.010 31.380 34.340 31.710 ;
        RECT 33.390 29.830 33.720 30.160 ;
        RECT 32.790 28.350 33.120 28.680 ;
        RECT 32.150 23.180 32.480 23.510 ;
        RECT 31.480 21.610 31.810 21.940 ;
        RECT 23.130 19.700 23.390 19.960 ;
        RECT 30.860 19.970 31.190 20.300 ;
        RECT 22.470 8.570 22.730 8.900 ;
        RECT 21.440 6.950 21.730 7.240 ;
        RECT 15.580 5.880 15.840 6.140 ;
        RECT 16.680 5.890 16.940 6.150 ;
        RECT 17.770 5.890 18.030 6.150 ;
        RECT 18.900 5.850 19.160 6.110 ;
        RECT 20.280 5.940 20.880 6.540 ;
        RECT 16.130 5.210 16.390 5.470 ;
        RECT 17.230 5.210 17.490 5.470 ;
        RECT 18.330 5.210 18.590 5.470 ;
        RECT 16.130 3.840 16.390 4.100 ;
        RECT 17.230 3.840 17.490 4.100 ;
        RECT 18.330 3.840 18.590 4.100 ;
        RECT 15.580 3.110 15.840 3.370 ;
        RECT 16.680 3.110 16.940 3.370 ;
        RECT 17.770 3.110 18.030 3.370 ;
        RECT 15.570 1.770 15.830 2.030 ;
        RECT 16.680 1.760 16.940 2.020 ;
        RECT 17.770 1.740 18.030 2.000 ;
        RECT 30.180 18.530 30.510 18.860 ;
        RECT 26.140 14.170 26.720 14.880 ;
        RECT 16.130 1.070 16.390 1.330 ;
        RECT 17.230 1.060 17.490 1.320 ;
        RECT 18.320 1.060 18.580 1.320 ;
        RECT 23.060 1.010 23.320 1.350 ;
        RECT 4.150 0.070 4.540 0.460 ;
        RECT 30.150 -5.300 30.580 -4.870 ;
        RECT 30.800 -6.090 31.230 -5.660 ;
        RECT 31.470 -6.770 31.870 -6.370 ;
        RECT 31.300 -7.710 31.810 -7.200 ;
        RECT 41.040 47.410 41.300 47.670 ;
        RECT 41.040 45.660 41.300 45.920 ;
        RECT 41.040 43.910 41.300 44.170 ;
        RECT 41.040 43.120 41.300 43.380 ;
        RECT 41.040 41.370 41.300 41.630 ;
        RECT 41.040 39.620 41.300 39.880 ;
        RECT 41.040 37.870 41.300 38.130 ;
        RECT 46.860 50.010 47.120 50.270 ;
        RECT 47.900 50.050 48.160 50.310 ;
        RECT 43.140 48.250 43.400 48.510 ;
        RECT 43.140 46.500 43.400 46.760 ;
        RECT 43.140 44.750 43.400 45.010 ;
        RECT 43.140 42.280 43.400 42.540 ;
        RECT 43.140 40.530 43.400 40.790 ;
        RECT 43.140 38.780 43.400 39.040 ;
        RECT 45.180 49.280 45.440 49.540 ;
        RECT 46.860 48.260 47.120 48.520 ;
        RECT 47.900 48.300 48.160 48.560 ;
        RECT 45.180 47.530 45.440 47.790 ;
        RECT 46.860 46.510 47.120 46.770 ;
        RECT 47.900 46.550 48.160 46.810 ;
        RECT 45.180 45.780 45.440 46.040 ;
        RECT 46.860 44.760 47.120 45.020 ;
        RECT 47.900 44.800 48.160 45.060 ;
        RECT 45.180 44.030 45.440 44.290 ;
        RECT 45.180 43.000 45.440 43.260 ;
        RECT 46.860 42.270 47.120 42.530 ;
        RECT 47.900 42.230 48.160 42.490 ;
        RECT 45.180 41.250 45.440 41.510 ;
        RECT 46.860 40.520 47.120 40.780 ;
        RECT 47.900 40.480 48.160 40.740 ;
        RECT 45.180 39.500 45.440 39.760 ;
        RECT 46.860 38.770 47.120 39.030 ;
        RECT 47.900 38.730 48.160 38.990 ;
        RECT 45.180 37.750 45.440 38.010 ;
        RECT 43.140 37.030 43.400 37.290 ;
        RECT 46.860 37.020 47.120 37.280 ;
        RECT 47.900 36.980 48.160 37.240 ;
        RECT 41.040 32.990 41.300 33.250 ;
        RECT 41.040 31.240 41.300 31.500 ;
        RECT 41.040 29.490 41.300 29.750 ;
        RECT 41.040 27.740 41.300 28.000 ;
        RECT 43.140 32.150 43.400 32.410 ;
        RECT 43.140 30.400 43.400 30.660 ;
        RECT 43.140 28.650 43.400 28.910 ;
        RECT 45.180 32.870 45.440 33.130 ;
        RECT 46.860 32.140 47.120 32.400 ;
        RECT 47.900 32.100 48.160 32.360 ;
        RECT 45.180 31.120 45.440 31.380 ;
        RECT 46.860 30.390 47.120 30.650 ;
        RECT 47.900 30.350 48.160 30.610 ;
        RECT 45.180 29.370 45.440 29.630 ;
        RECT 46.860 28.640 47.120 28.900 ;
        RECT 47.900 28.600 48.160 28.860 ;
        RECT 45.180 27.620 45.440 27.880 ;
        RECT 41.000 23.930 41.260 24.190 ;
        RECT 43.140 26.900 43.400 27.160 ;
        RECT 46.860 26.890 47.120 27.150 ;
        RECT 47.900 26.850 48.160 27.110 ;
        RECT 50.160 56.190 50.600 56.630 ;
        RECT 51.060 43.060 51.320 43.320 ;
        RECT 49.970 42.540 50.230 42.800 ;
        RECT 49.970 41.270 50.230 41.530 ;
        RECT 51.060 40.750 51.320 41.010 ;
        RECT 51.060 39.860 51.320 40.120 ;
        RECT 49.970 39.340 50.230 39.600 ;
        RECT 49.970 38.070 50.230 38.330 ;
        RECT 51.060 37.550 51.320 37.810 ;
        RECT 64.560 56.190 65.000 56.630 ;
        RECT 58.810 52.410 59.070 52.670 ;
        RECT 56.930 48.880 57.190 49.140 ;
        RECT 62.400 51.500 62.660 51.760 ;
        RECT 59.270 50.480 59.530 50.740 ;
        RECT 58.380 46.020 58.640 46.280 ;
        RECT 53.470 43.060 53.730 43.320 ;
        RECT 57.990 44.490 58.250 44.750 ;
        RECT 59.690 48.390 59.950 48.650 ;
        RECT 57.280 43.660 57.540 43.920 ;
        RECT 60.750 47.910 61.010 48.170 ;
        RECT 57.980 42.800 58.240 43.060 ;
        RECT 53.470 40.750 53.730 41.010 ;
        RECT 58.380 41.290 58.640 41.550 ;
        RECT 65.570 52.420 65.830 52.680 ;
        RECT 65.130 51.510 65.390 51.770 ;
        RECT 62.390 40.810 62.660 41.080 ;
        RECT 64.640 40.830 64.900 41.090 ;
        RECT 53.470 39.860 53.730 40.120 ;
        RECT 58.390 39.990 58.650 40.250 ;
        RECT 58.240 39.030 58.500 39.290 ;
        RECT 53.470 37.550 53.730 37.810 ;
        RECT 57.300 37.920 57.560 38.180 ;
        RECT 57.300 37.320 57.560 37.580 ;
        RECT 58.240 36.270 58.500 36.530 ;
        RECT 58.390 35.260 58.650 35.520 ;
        RECT 51.040 32.590 51.300 32.850 ;
        RECT 49.950 32.070 50.210 32.330 ;
        RECT 49.950 30.800 50.210 31.060 ;
        RECT 51.040 30.280 51.300 30.540 ;
        RECT 51.040 29.390 51.300 29.650 ;
        RECT 49.950 28.870 50.210 29.130 ;
        RECT 49.950 27.600 50.210 27.860 ;
        RECT 53.450 32.590 53.710 32.850 ;
        RECT 59.030 34.170 59.310 34.450 ;
        RECT 70.360 56.150 70.800 56.590 ;
        RECT 78.690 57.180 78.970 57.620 ;
        RECT 74.910 50.520 76.130 50.780 ;
        RECT 71.670 49.870 71.930 50.130 ;
        RECT 78.000 49.330 78.260 49.590 ;
        RECT 76.710 46.020 76.970 46.280 ;
        RECT 80.340 52.420 80.600 52.680 ;
        RECT 79.450 51.550 79.710 51.810 ;
        RECT 86.860 61.520 87.230 61.890 ;
        RECT 83.010 53.130 83.270 53.400 ;
        RECT 79.450 47.340 79.710 47.600 ;
        RECT 80.470 47.350 80.730 47.610 ;
        RECT 78.690 46.510 78.950 46.770 ;
        RECT 80.420 46.500 80.680 46.760 ;
        RECT 81.400 46.250 81.660 46.510 ;
        RECT 80.570 45.670 80.830 45.930 ;
        RECT 81.350 45.600 81.610 45.860 ;
        RECT 76.860 45.060 77.120 45.320 ;
        RECT 77.800 43.950 78.060 44.210 ;
        RECT 77.800 43.350 78.060 43.610 ;
        RECT 79.460 45.140 79.720 45.400 ;
        RECT 80.630 44.660 80.890 44.920 ;
        RECT 81.350 44.750 81.610 45.010 ;
        RECT 78.740 43.670 79.000 43.930 ;
        RECT 80.190 43.860 80.450 44.120 ;
        RECT 76.860 42.300 77.120 42.560 ;
        RECT 70.440 40.830 70.700 41.090 ;
        RECT 65.500 39.440 65.760 39.700 ;
        RECT 64.710 37.390 64.970 37.650 ;
        RECT 65.530 35.750 65.790 36.010 ;
        RECT 76.710 41.290 76.970 41.550 ;
        RECT 76.710 39.990 76.970 40.250 ;
        RECT 81.400 44.100 81.660 44.360 ;
        RECT 81.400 43.250 81.660 43.510 ;
        RECT 81.350 42.600 81.610 42.860 ;
        RECT 81.350 41.750 81.610 42.010 ;
        RECT 80.830 40.980 81.090 41.240 ;
        RECT 81.400 41.100 81.660 41.360 ;
        RECT 83.220 47.230 83.650 47.660 ;
        RECT 78.670 40.450 78.930 40.710 ;
        RECT 80.420 40.470 80.680 40.730 ;
        RECT 81.400 40.220 81.660 40.480 ;
        RECT 80.570 39.640 80.830 39.900 ;
        RECT 81.350 39.570 81.610 39.830 ;
        RECT 76.860 39.030 77.120 39.290 ;
        RECT 70.410 37.330 70.670 37.590 ;
        RECT 77.800 37.920 78.060 38.180 ;
        RECT 77.800 37.320 78.060 37.580 ;
        RECT 79.460 39.110 79.720 39.370 ;
        RECT 80.630 38.630 80.890 38.890 ;
        RECT 81.350 38.720 81.610 38.980 ;
        RECT 78.740 37.640 79.000 37.900 ;
        RECT 80.190 37.830 80.450 38.090 ;
        RECT 76.860 36.270 77.120 36.530 ;
        RECT 70.410 34.810 70.670 35.070 ;
        RECT 59.790 32.540 60.050 32.800 ;
        RECT 53.450 30.280 53.710 30.540 ;
        RECT 59.790 31.990 60.050 32.250 ;
        RECT 59.790 31.000 60.050 31.260 ;
        RECT 59.790 30.450 60.050 30.710 ;
        RECT 53.450 29.390 53.710 29.650 ;
        RECT 59.790 29.300 60.050 29.560 ;
        RECT 51.040 27.080 51.300 27.340 ;
        RECT 53.450 27.080 53.710 27.340 ;
        RECT 59.790 28.750 60.050 29.010 ;
        RECT 60.710 28.330 60.970 28.590 ;
        RECT 59.790 27.770 60.050 28.030 ;
        RECT 64.640 28.290 64.900 28.550 ;
        RECT 59.790 27.220 60.050 27.480 ;
        RECT 76.710 35.260 76.970 35.520 ;
        RECT 81.400 38.070 81.660 38.330 ;
        RECT 81.400 37.220 81.660 37.480 ;
        RECT 81.350 36.570 81.610 36.830 ;
        RECT 81.350 35.720 81.610 35.980 ;
        RECT 76.380 33.600 76.640 33.860 ;
        RECT 75.290 32.540 75.550 32.800 ;
        RECT 80.850 34.940 81.120 35.200 ;
        RECT 81.400 35.070 81.660 35.330 ;
        RECT 83.650 46.270 83.910 46.530 ;
        RECT 83.700 44.050 83.960 44.310 ;
        RECT 83.690 43.330 83.950 43.590 ;
        RECT 83.610 41.080 83.870 41.340 ;
        RECT 83.650 40.240 83.910 40.500 ;
        RECT 83.700 38.020 83.960 38.280 ;
        RECT 83.690 37.300 83.950 37.560 ;
        RECT 83.610 35.050 83.870 35.310 ;
        RECT 87.680 58.060 88.050 58.430 ;
        RECT 86.870 34.150 87.240 34.520 ;
        RECT 88.450 53.350 88.820 53.720 ;
        RECT 75.290 31.990 75.550 32.250 ;
        RECT 87.640 33.560 88.010 33.930 ;
        RECT 77.250 32.870 77.510 33.130 ;
        RECT 70.440 28.290 70.700 28.550 ;
        RECT 75.290 31.000 75.550 31.260 ;
        RECT 95.000 52.300 95.500 52.800 ;
        RECT 91.780 50.740 92.280 51.240 ;
        RECT 92.730 51.230 93.230 51.730 ;
        RECT 93.810 51.700 94.310 52.200 ;
        RECT 89.330 48.280 89.700 48.650 ;
        RECT 75.290 30.450 75.550 30.710 ;
        RECT 88.380 31.230 88.750 31.600 ;
        RECT 75.290 29.300 75.550 29.560 ;
        RECT 75.290 28.750 75.550 29.010 ;
        RECT 74.370 28.330 74.630 28.590 ;
        RECT 75.290 27.770 75.550 28.030 ;
        RECT 75.290 27.220 75.550 27.480 ;
        RECT 45.140 23.810 45.400 24.070 ;
        RECT 41.000 22.180 41.260 22.440 ;
        RECT 41.000 20.430 41.260 20.690 ;
        RECT 41.000 18.680 41.260 18.940 ;
        RECT 51.660 25.980 51.920 26.390 ;
        RECT 43.100 23.090 43.360 23.350 ;
        RECT 43.100 21.340 43.360 21.600 ;
        RECT 43.100 19.590 43.360 19.850 ;
        RECT 43.100 17.840 43.360 18.100 ;
        RECT 46.820 23.080 47.080 23.340 ;
        RECT 47.860 23.040 48.120 23.300 ;
        RECT 45.140 22.060 45.400 22.320 ;
        RECT 46.820 21.330 47.080 21.590 ;
        RECT 47.860 21.290 48.120 21.550 ;
        RECT 45.140 20.310 45.400 20.570 ;
        RECT 46.820 19.580 47.080 19.840 ;
        RECT 47.860 19.540 48.120 19.800 ;
        RECT 45.140 18.560 45.400 18.820 ;
        RECT 46.820 17.830 47.080 18.090 ;
        RECT 47.860 17.790 48.120 18.050 ;
        RECT 51.070 23.320 51.330 23.580 ;
        RECT 49.980 22.800 50.240 23.060 ;
        RECT 49.980 21.530 50.240 21.790 ;
        RECT 51.070 21.010 51.330 21.270 ;
        RECT 51.070 20.120 51.330 20.380 ;
        RECT 49.980 19.600 50.240 19.860 ;
        RECT 49.980 18.330 50.240 18.590 ;
        RECT 51.070 17.810 51.330 18.070 ;
        RECT 53.480 23.320 53.740 23.580 ;
        RECT 59.820 23.210 60.080 23.470 ;
        RECT 60.430 23.110 60.690 23.370 ;
        RECT 56.060 22.260 56.320 22.520 ;
        RECT 53.480 21.010 53.740 21.270 ;
        RECT 53.480 20.120 53.740 20.380 ;
        RECT 53.480 17.810 53.740 18.070 ;
        RECT 57.140 21.560 57.400 21.820 ;
        RECT 59.820 22.660 60.080 22.920 ;
        RECT 60.410 22.060 60.670 22.320 ;
        RECT 59.820 21.690 60.080 21.950 ;
        RECT 57.120 20.550 57.380 20.810 ;
        RECT 59.820 21.140 60.080 21.400 ;
        RECT 56.690 19.480 56.950 19.740 ;
        RECT 49.480 17.130 49.740 17.390 ;
        RECT 48.940 16.760 49.230 17.050 ;
        RECT 44.500 16.250 44.810 16.560 ;
        RECT 56.090 17.170 56.350 17.430 ;
        RECT 57.070 18.510 57.330 18.770 ;
        RECT 57.120 17.550 57.380 17.810 ;
        RECT 57.120 17.160 57.380 17.420 ;
        RECT 54.690 16.760 54.950 17.020 ;
        RECT 56.660 16.840 56.920 17.100 ;
        RECT 48.310 15.540 48.730 15.960 ;
        RECT 44.460 14.580 44.880 15.000 ;
        RECT 50.370 16.220 50.630 16.480 ;
        RECT 59.820 19.970 60.080 20.230 ;
        RECT 60.410 20.180 60.670 20.440 ;
        RECT 59.820 19.420 60.080 19.680 ;
        RECT 60.280 19.000 60.540 19.260 ;
        RECT 60.860 18.920 61.120 19.180 ;
        RECT 59.820 18.440 60.080 18.700 ;
        RECT 59.820 17.890 60.080 18.150 ;
        RECT 58.900 16.780 59.160 17.040 ;
        RECT 49.780 15.550 50.040 15.810 ;
        RECT 50.870 15.550 51.130 15.810 ;
        RECT 51.970 15.540 52.230 15.800 ;
        RECT 54.810 15.540 55.070 15.800 ;
        RECT 55.910 15.550 56.170 15.810 ;
        RECT 57.000 15.550 57.260 15.810 ;
        RECT 57.700 15.530 58.030 15.860 ;
        RECT 64.880 18.900 65.150 19.160 ;
        RECT 89.310 25.980 89.680 26.390 ;
        RECT 68.510 22.910 68.770 23.170 ;
        RECT 68.660 22.230 68.920 22.490 ;
        RECT 68.660 21.340 68.920 21.600 ;
        RECT 68.510 20.660 68.770 20.920 ;
        RECT 68.510 20.140 68.770 20.400 ;
        RECT 68.660 19.460 68.920 19.720 ;
        RECT 68.660 18.570 68.920 18.830 ;
        RECT 68.510 17.890 68.770 18.150 ;
        RECT 75.940 22.240 76.200 22.500 ;
        RECT 75.420 21.310 75.680 21.570 ;
        RECT 74.950 19.470 75.210 19.730 ;
        RECT 70.790 19.010 71.060 19.280 ;
        RECT 67.740 17.090 68.090 17.440 ;
        RECT 60.890 16.360 61.150 16.620 ;
        RECT 64.930 16.330 65.200 16.600 ;
        RECT 58.850 15.460 59.190 15.800 ;
        RECT 59.590 15.580 59.850 15.840 ;
        RECT 60.680 15.580 60.940 15.840 ;
        RECT 61.780 15.570 62.040 15.830 ;
        RECT 64.620 15.570 64.880 15.830 ;
        RECT 65.720 15.580 65.980 15.840 ;
        RECT 66.810 15.580 67.070 15.840 ;
        RECT 74.450 18.540 74.710 18.800 ;
        RECT 67.780 15.320 68.040 15.640 ;
        RECT 50.330 14.870 50.590 15.130 ;
        RECT 51.420 14.850 51.680 15.110 ;
        RECT 55.360 14.850 55.620 15.110 ;
        RECT 56.450 14.870 56.710 15.130 ;
        RECT 60.140 14.900 60.400 15.160 ;
        RECT 61.230 14.880 61.490 15.140 ;
        RECT 65.170 14.880 65.430 15.140 ;
        RECT 66.260 14.900 66.520 15.160 ;
        RECT 70.360 15.560 70.620 15.820 ;
        RECT 71.460 15.570 71.720 15.830 ;
        RECT 72.550 15.570 72.810 15.830 ;
        RECT 73.770 15.540 74.030 15.880 ;
        RECT 48.990 14.490 49.310 14.810 ;
        RECT 69.200 14.610 69.580 14.990 ;
        RECT 69.800 14.860 70.060 15.120 ;
        RECT 70.910 14.870 71.170 15.130 ;
        RECT 72.000 14.890 72.260 15.150 ;
        RECT 50.330 13.500 50.590 13.760 ;
        RECT 51.420 13.500 51.680 13.760 ;
        RECT 55.360 13.500 55.620 13.760 ;
        RECT 56.450 13.500 56.710 13.760 ;
        RECT 60.140 13.530 60.400 13.790 ;
        RECT 61.230 13.530 61.490 13.790 ;
        RECT 65.170 13.530 65.430 13.790 ;
        RECT 66.260 13.530 66.520 13.790 ;
        RECT 69.810 13.520 70.070 13.780 ;
        RECT 70.910 13.520 71.170 13.780 ;
        RECT 72.000 13.520 72.260 13.780 ;
        RECT 49.770 12.770 50.030 13.030 ;
        RECT 50.870 12.770 51.130 13.030 ;
        RECT 51.970 12.770 52.230 13.030 ;
        RECT 54.810 12.770 55.070 13.030 ;
        RECT 55.910 12.770 56.170 13.030 ;
        RECT 57.010 12.770 57.270 13.030 ;
        RECT 59.580 12.800 59.840 13.060 ;
        RECT 60.680 12.800 60.940 13.060 ;
        RECT 61.780 12.800 62.040 13.060 ;
        RECT 64.620 12.800 64.880 13.060 ;
        RECT 65.720 12.800 65.980 13.060 ;
        RECT 66.820 12.800 67.080 13.060 ;
        RECT 70.360 12.790 70.620 13.050 ;
        RECT 71.460 12.790 71.720 13.050 ;
        RECT 72.560 12.790 72.820 13.050 ;
        RECT 49.770 11.400 50.030 11.660 ;
        RECT 50.870 11.400 51.130 11.660 ;
        RECT 51.970 11.400 52.230 11.660 ;
        RECT 54.810 11.400 55.070 11.660 ;
        RECT 55.910 11.400 56.170 11.660 ;
        RECT 57.010 11.400 57.270 11.660 ;
        RECT 59.580 11.430 59.840 11.690 ;
        RECT 60.680 11.430 60.940 11.690 ;
        RECT 61.780 11.430 62.040 11.690 ;
        RECT 64.620 11.430 64.880 11.690 ;
        RECT 65.720 11.430 65.980 11.690 ;
        RECT 66.820 11.430 67.080 11.690 ;
        RECT 70.360 11.420 70.620 11.680 ;
        RECT 71.460 11.420 71.720 11.680 ;
        RECT 72.560 11.420 72.820 11.680 ;
        RECT 49.200 10.760 49.460 11.020 ;
        RECT 50.330 10.720 50.590 10.980 ;
        RECT 51.420 10.720 51.680 10.980 ;
        RECT 55.360 10.720 55.620 10.980 ;
        RECT 56.450 10.720 56.710 10.980 ;
        RECT 57.580 10.760 57.840 11.020 ;
        RECT 49.210 10.290 49.470 10.550 ;
        RECT 57.570 10.290 57.830 10.550 ;
        RECT 49.090 8.710 49.550 9.170 ;
        RECT 59.010 10.790 59.270 11.050 ;
        RECT 60.140 10.750 60.400 11.010 ;
        RECT 61.230 10.750 61.490 11.010 ;
        RECT 65.170 10.750 65.430 11.010 ;
        RECT 66.260 10.750 66.520 11.010 ;
        RECT 67.390 10.790 67.650 11.050 ;
        RECT 69.810 10.750 70.070 11.010 ;
        RECT 70.910 10.740 71.170 11.000 ;
        RECT 72.000 10.740 72.260 11.000 ;
        RECT 73.130 10.780 73.390 11.040 ;
        RECT 103.810 49.360 105.090 50.640 ;
        RECT 108.130 47.200 108.390 47.630 ;
        RECT 104.300 45.920 104.560 46.340 ;
        RECT 100.300 42.720 100.700 43.120 ;
        RECT 94.910 30.020 95.410 30.520 ;
        RECT 93.830 24.830 94.330 25.300 ;
        RECT 92.700 19.640 93.200 20.140 ;
        RECT 91.650 14.340 92.150 14.840 ;
        RECT 75.920 12.830 76.180 13.330 ;
        RECT 75.380 11.930 75.640 12.430 ;
        RECT 74.910 11.030 75.170 11.530 ;
        RECT 59.020 10.320 59.280 10.580 ;
        RECT 67.380 10.320 67.640 10.580 ;
        RECT 73.120 10.310 73.380 10.570 ;
        RECT 57.470 7.760 57.930 8.220 ;
        RECT 58.900 6.870 59.360 7.330 ;
        RECT 67.290 5.960 67.750 6.420 ;
        RECT 41.220 3.730 41.480 4.850 ;
        RECT 74.430 10.130 74.690 10.630 ;
        RECT 97.890 16.860 98.390 17.360 ;
        RECT 95.020 8.750 95.520 9.250 ;
        RECT 93.830 7.800 94.330 8.260 ;
        RECT 92.700 6.930 93.200 7.390 ;
        RECT 91.770 6.020 92.270 6.480 ;
        RECT 97.310 3.730 98.250 4.850 ;
        RECT 73.100 0.100 73.430 0.430 ;
        RECT 39.540 -0.560 39.870 -0.230 ;
        RECT 101.280 42.080 101.640 42.440 ;
        RECT 38.920 -1.180 39.250 -0.850 ;
        RECT 100.360 -1.090 100.760 -0.690 ;
        RECT 102.200 39.710 102.590 40.100 ;
        RECT 38.290 -1.810 38.620 -1.480 ;
        RECT 101.270 -1.890 101.660 -1.500 ;
        RECT 37.690 -2.440 38.020 -2.110 ;
        RECT 103.030 39.150 103.410 39.410 ;
        RECT 102.200 -2.710 102.590 -2.320 ;
        RECT 37.050 -3.120 37.380 -2.790 ;
        RECT 109.110 43.790 109.370 44.050 ;
        RECT 110.680 43.790 110.940 44.050 ;
        RECT 107.760 42.810 108.020 43.070 ;
        RECT 115.080 54.690 115.790 55.400 ;
        RECT 107.760 42.200 108.020 42.460 ;
        RECT 110.030 42.880 110.290 43.140 ;
        RECT 111.040 42.870 111.300 43.130 ;
        RECT 110.030 42.130 110.290 42.390 ;
        RECT 111.040 42.140 111.300 42.400 ;
        RECT 109.110 41.220 109.370 41.480 ;
        RECT 110.680 41.220 110.940 41.480 ;
        RECT 109.110 40.590 109.370 40.850 ;
        RECT 110.680 40.590 110.940 40.850 ;
        RECT 107.760 39.610 108.020 39.870 ;
        RECT 107.760 39.000 108.020 39.260 ;
        RECT 110.030 39.680 110.290 39.940 ;
        RECT 111.040 39.670 111.300 39.930 ;
        RECT 110.030 38.930 110.290 39.190 ;
        RECT 111.040 38.940 111.300 39.200 ;
        RECT 109.110 38.020 109.370 38.280 ;
        RECT 110.680 38.020 110.940 38.280 ;
        RECT 114.890 34.900 115.600 35.610 ;
        RECT 110.690 16.850 111.200 17.360 ;
        RECT 109.900 7.040 110.160 7.300 ;
        RECT 109.900 6.370 110.160 6.630 ;
        RECT 110.060 5.130 110.320 5.390 ;
        RECT 105.120 1.800 105.380 2.060 ;
        RECT 110.060 3.520 110.320 3.780 ;
        RECT 110.050 1.910 110.310 2.170 ;
        RECT 110.060 0.290 110.320 0.550 ;
        RECT 110.050 -1.320 110.310 -1.060 ;
        RECT 36.450 -3.740 36.780 -3.410 ;
        RECT 103.020 -3.500 103.400 -3.120 ;
        RECT 109.640 -2.970 109.900 -2.710 ;
        RECT 35.850 -4.380 36.180 -4.050 ;
        RECT 110.050 -4.520 110.310 -4.260 ;
        RECT 35.270 -4.950 35.600 -4.620 ;
        RECT 34.690 -5.640 35.020 -5.310 ;
        RECT 34.040 -6.280 34.370 -5.950 ;
        RECT 106.810 -6.230 107.070 -5.970 ;
        RECT 107.750 -6.230 108.010 -5.970 ;
        RECT 108.700 -6.250 108.960 -5.990 ;
        RECT 110.010 -6.230 110.270 -5.970 ;
        RECT 33.400 -6.930 33.730 -6.590 ;
        RECT 32.820 -7.570 33.190 -7.200 ;
      LAYER met2 ;
        RECT 9.460 61.490 9.780 61.540 ;
        RECT 6.600 61.250 9.780 61.490 ;
        RECT 6.600 61.230 6.920 61.250 ;
        RECT 34.590 52.740 34.900 52.760 ;
        RECT 24.800 52.660 25.120 52.670 ;
        RECT 34.590 52.660 34.910 52.740 ;
        RECT 58.770 52.670 59.090 52.690 ;
        RECT 58.770 52.660 59.100 52.670 ;
        RECT 65.540 52.660 65.860 52.690 ;
        RECT 80.310 52.660 80.630 52.680 ;
        RECT 94.970 52.660 95.530 52.800 ;
        RECT 24.800 52.430 95.530 52.660 ;
        RECT 24.800 52.350 25.120 52.430 ;
        RECT 34.590 52.420 34.900 52.430 ;
        RECT 58.770 52.410 59.100 52.430 ;
        RECT 65.540 52.410 65.860 52.430 ;
        RECT 80.310 52.420 80.630 52.430 ;
        RECT 94.970 52.290 95.530 52.430 ;
        RECT 62.390 51.760 62.670 51.770 ;
        RECT 33.420 51.750 33.730 51.760 ;
        RECT 62.370 51.750 62.690 51.760 ;
        RECT 65.100 51.750 65.420 51.780 ;
        RECT 79.420 51.750 79.740 51.810 ;
        RECT 92.710 51.750 93.250 51.760 ;
        RECT 33.420 51.520 93.250 51.750 ;
        RECT 33.420 51.490 33.750 51.520 ;
        RECT 62.370 51.500 62.690 51.520 ;
        RECT 65.100 51.500 65.420 51.520 ;
        RECT 62.390 51.490 62.670 51.500 ;
        RECT 33.420 51.470 33.730 51.490 ;
        RECT 92.710 51.200 93.250 51.520 ;
        RECT 43.140 49.490 43.400 50.290 ;
        RECT 45.140 49.490 45.480 49.550 ;
        RECT 43.040 49.270 45.480 49.490 ;
        RECT 59.660 48.650 59.970 48.660 ;
        RECT 59.660 48.620 59.980 48.650 ;
        RECT 43.140 47.740 43.400 48.540 ;
        RECT 52.410 48.420 59.980 48.620 ;
        RECT 45.140 47.740 45.480 47.800 ;
        RECT 43.040 47.520 45.480 47.740 ;
        RECT 43.140 45.990 43.400 46.790 ;
        RECT 46.840 46.770 47.160 46.780 ;
        RECT 46.830 46.760 47.160 46.770 ;
        RECT 47.870 46.760 48.190 46.810 ;
        RECT 52.410 46.760 52.610 48.420 ;
        RECT 59.660 48.390 59.980 48.420 ;
        RECT 59.660 48.380 59.970 48.390 ;
        RECT 60.720 48.140 61.040 48.180 ;
        RECT 46.830 46.560 52.610 46.760 ;
        RECT 52.960 47.940 61.120 48.140 ;
        RECT 46.830 46.510 47.160 46.560 ;
        RECT 47.870 46.550 48.190 46.560 ;
        RECT 46.840 46.490 47.160 46.510 ;
        RECT 45.140 45.990 45.480 46.050 ;
        RECT 43.040 45.770 45.480 45.990 ;
        RECT 43.140 44.240 43.400 45.040 ;
        RECT 46.840 45.020 47.160 45.030 ;
        RECT 46.830 45.010 47.160 45.020 ;
        RECT 47.870 45.010 48.190 45.060 ;
        RECT 52.960 45.010 53.160 47.940 ;
        RECT 60.720 47.900 61.040 47.940 ;
        RECT 79.360 47.340 79.940 47.780 ;
        RECT 79.360 47.150 80.000 47.340 ;
        RECT 79.760 46.790 80.000 47.150 ;
        RECT 80.380 47.140 80.960 47.770 ;
        RECT 80.400 46.790 80.710 46.800 ;
        RECT 79.760 46.540 80.710 46.790 ;
        RECT 80.400 46.470 80.710 46.540 ;
        RECT 81.370 46.470 81.680 46.550 ;
        RECT 83.620 46.470 83.930 46.570 ;
        RECT 58.600 46.320 58.920 46.330 ;
        RECT 46.830 44.810 53.160 45.010 ;
        RECT 56.110 46.310 56.400 46.320 ;
        RECT 58.360 46.310 58.920 46.320 ;
        RECT 76.680 46.310 76.990 46.320 ;
        RECT 56.110 46.130 79.160 46.310 ;
        RECT 81.370 46.240 83.930 46.470 ;
        RECT 81.370 46.220 81.680 46.240 ;
        RECT 46.830 44.760 47.160 44.810 ;
        RECT 47.870 44.800 48.190 44.810 ;
        RECT 46.840 44.740 47.160 44.760 ;
        RECT 45.140 44.240 45.480 44.300 ;
        RECT 43.040 44.020 45.480 44.240 ;
        RECT 51.030 43.300 51.350 43.350 ;
        RECT 53.440 43.300 53.760 43.320 ;
        RECT 56.110 43.300 56.290 46.130 ;
        RECT 58.360 45.990 58.670 46.130 ;
        RECT 76.680 45.990 76.990 46.130 ;
        RECT 80.550 45.930 80.860 45.970 ;
        RECT 80.370 45.820 81.090 45.930 ;
        RECT 81.320 45.820 81.630 45.900 ;
        RECT 80.370 45.680 81.630 45.820 ;
        RECT 80.550 45.640 81.630 45.680 ;
        RECT 80.820 45.610 81.630 45.640 ;
        RECT 80.820 45.570 81.090 45.610 ;
        RECT 81.320 45.570 81.630 45.610 ;
        RECT 76.830 45.290 77.140 45.360 ;
        RECT 79.430 45.290 79.740 45.430 ;
        RECT 76.830 45.100 79.740 45.290 ;
        RECT 76.830 45.070 79.430 45.100 ;
        RECT 76.830 45.030 77.140 45.070 ;
        RECT 80.890 45.000 81.090 45.010 ;
        RECT 81.320 45.000 81.630 45.040 ;
        RECT 80.890 44.920 81.630 45.000 ;
        RECT 80.600 44.900 81.630 44.920 ;
        RECT 80.550 44.790 81.630 44.900 ;
        RECT 57.970 44.770 58.280 44.790 ;
        RECT 67.700 44.770 75.690 44.780 ;
        RECT 57.970 44.580 75.690 44.770 ;
        RECT 80.550 44.660 81.110 44.790 ;
        RECT 81.320 44.710 81.630 44.790 ;
        RECT 80.550 44.650 81.020 44.660 ;
        RECT 57.970 44.460 58.280 44.580 ;
        RECT 57.250 43.890 57.570 43.920 ;
        RECT 74.290 43.900 74.510 43.910 ;
        RECT 67.710 43.890 74.540 43.900 ;
        RECT 57.250 43.660 74.540 43.890 ;
        RECT 75.470 43.860 75.690 44.580 ;
        RECT 81.370 44.330 81.680 44.390 ;
        RECT 83.670 44.330 83.980 44.350 ;
        RECT 80.460 44.150 81.060 44.270 ;
        RECT 80.160 44.110 81.060 44.150 ;
        RECT 79.840 43.870 81.060 44.110 ;
        RECT 81.370 44.100 89.290 44.330 ;
        RECT 89.660 44.100 98.810 44.330 ;
        RECT 81.370 44.060 81.680 44.100 ;
        RECT 83.670 44.020 83.980 44.100 ;
        RECT 67.710 43.650 74.540 43.660 ;
        RECT 43.040 43.050 45.480 43.270 ;
        RECT 43.140 42.250 43.400 43.050 ;
        RECT 45.140 42.990 45.480 43.050 ;
        RECT 51.030 43.130 56.290 43.300 ;
        RECT 51.030 43.110 53.760 43.130 ;
        RECT 51.030 43.030 51.350 43.110 ;
        RECT 53.440 43.060 53.760 43.110 ;
        RECT 57.960 42.910 58.270 43.100 ;
        RECT 67.710 42.910 71.220 42.920 ;
        RECT 46.840 42.530 47.160 42.550 ;
        RECT 46.830 42.480 47.160 42.530 ;
        RECT 49.680 42.520 50.270 42.820 ;
        RECT 57.960 42.770 71.220 42.910 ;
        RECT 57.990 42.730 71.220 42.770 ;
        RECT 57.990 42.720 67.710 42.730 ;
        RECT 49.680 42.500 50.030 42.520 ;
        RECT 47.870 42.480 48.190 42.490 ;
        RECT 49.680 42.480 49.880 42.500 ;
        RECT 46.830 42.280 49.880 42.480 ;
        RECT 46.830 42.270 47.160 42.280 ;
        RECT 46.840 42.260 47.160 42.270 ;
        RECT 47.870 42.230 48.190 42.280 ;
        RECT 70.990 42.130 71.220 42.730 ;
        RECT 74.250 42.480 74.540 43.650 ;
        RECT 75.440 43.820 75.690 43.860 ;
        RECT 80.160 43.820 81.060 43.870 ;
        RECT 75.440 43.180 75.700 43.820 ;
        RECT 80.460 43.710 81.060 43.820 ;
        RECT 98.520 44.000 98.810 44.100 ;
        RECT 108.310 44.080 109.430 44.090 ;
        RECT 106.500 44.000 110.960 44.080 ;
        RECT 98.520 43.880 110.960 44.000 ;
        RECT 98.520 43.800 106.850 43.880 ;
        RECT 108.310 43.870 109.430 43.880 ;
        RECT 98.520 43.790 98.810 43.800 ;
        RECT 109.080 43.750 109.390 43.870 ;
        RECT 110.650 43.750 110.960 43.880 ;
        RECT 81.370 43.500 81.680 43.550 ;
        RECT 83.660 43.500 83.970 43.630 ;
        RECT 81.370 43.280 89.290 43.500 ;
        RECT 89.660 43.280 97.870 43.500 ;
        RECT 81.370 43.220 81.680 43.280 ;
        RECT 75.440 42.970 79.570 43.180 ;
        RECT 79.360 42.830 79.570 42.970 ;
        RECT 81.320 42.830 81.630 42.900 ;
        RECT 79.360 42.620 81.630 42.830 ;
        RECT 81.020 42.610 81.630 42.620 ;
        RECT 76.830 42.530 77.140 42.600 ;
        RECT 81.320 42.570 81.630 42.610 ;
        RECT 76.830 42.480 79.160 42.530 ;
        RECT 74.250 42.320 79.160 42.480 ;
        RECT 74.250 42.260 77.140 42.320 ;
        RECT 74.250 42.250 74.540 42.260 ;
        RECT 70.990 41.980 71.210 42.130 ;
        RECT 81.320 42.030 81.630 42.040 ;
        RECT 75.360 41.980 81.630 42.030 ;
        RECT 70.990 41.820 81.630 41.980 ;
        RECT 70.990 41.760 75.750 41.820 ;
        RECT 81.020 41.790 81.630 41.820 ;
        RECT 81.320 41.710 81.630 41.790 ;
        RECT 43.040 41.300 45.480 41.520 ;
        RECT 49.930 41.480 50.270 41.550 ;
        RECT 43.140 40.500 43.400 41.300 ;
        RECT 45.140 41.240 45.480 41.300 ;
        RECT 49.630 41.250 50.270 41.480 ;
        RECT 58.360 41.440 58.670 41.580 ;
        RECT 56.190 41.430 58.670 41.440 ;
        RECT 76.680 41.440 76.990 41.580 ;
        RECT 76.680 41.430 79.160 41.440 ;
        RECT 55.670 41.280 79.160 41.430 ;
        RECT 97.650 41.400 97.870 43.280 ;
        RECT 109.080 41.400 109.390 41.520 ;
        RECT 97.650 41.390 99.250 41.400 ;
        RECT 108.310 41.390 109.430 41.400 ;
        RECT 110.650 41.390 110.960 41.520 ;
        RECT 55.670 41.260 58.670 41.280 ;
        RECT 55.670 41.250 56.400 41.260 ;
        RECT 58.360 41.250 58.670 41.260 ;
        RECT 76.680 41.260 79.160 41.280 ;
        RECT 81.370 41.340 81.680 41.390 ;
        RECT 83.580 41.340 83.890 41.380 ;
        RECT 76.680 41.250 76.990 41.260 ;
        RECT 46.840 40.780 47.160 40.800 ;
        RECT 46.830 40.730 47.160 40.780 ;
        RECT 47.870 40.730 48.190 40.740 ;
        RECT 49.630 40.730 49.830 41.250 ;
        RECT 55.670 41.040 55.850 41.250 ;
        RECT 81.370 41.110 84.080 41.340 ;
        RECT 97.650 41.190 110.960 41.390 ;
        RECT 97.650 41.180 99.250 41.190 ;
        RECT 108.310 41.180 109.430 41.190 ;
        RECT 62.370 41.090 62.680 41.100 ;
        RECT 46.830 40.530 49.830 40.730 ;
        RECT 51.030 40.960 51.350 41.040 ;
        RECT 53.510 41.010 55.850 41.040 ;
        RECT 62.360 41.030 62.690 41.090 ;
        RECT 81.370 41.060 81.680 41.110 ;
        RECT 83.580 41.050 83.890 41.110 ;
        RECT 53.440 40.960 55.850 41.010 ;
        RECT 62.010 40.980 62.690 41.030 ;
        RECT 51.030 40.880 55.850 40.960 ;
        RECT 51.030 40.770 53.760 40.880 ;
        RECT 54.240 40.870 55.850 40.880 ;
        RECT 54.940 40.860 55.850 40.870 ;
        RECT 51.030 40.720 51.350 40.770 ;
        RECT 53.440 40.750 53.760 40.770 ;
        RECT 58.780 40.810 62.690 40.980 ;
        RECT 84.840 40.820 89.290 40.980 ;
        RECT 58.780 40.760 62.680 40.810 ;
        RECT 84.810 40.780 89.290 40.820 ;
        RECT 89.660 40.880 106.850 40.980 ;
        RECT 108.310 40.880 109.430 40.890 ;
        RECT 89.660 40.780 110.960 40.880 ;
        RECT 79.400 40.760 79.960 40.780 ;
        RECT 80.400 40.760 80.710 40.770 ;
        RECT 46.830 40.520 47.160 40.530 ;
        RECT 46.840 40.510 47.160 40.520 ;
        RECT 47.870 40.480 48.190 40.530 ;
        RECT 79.400 40.510 80.710 40.760 ;
        RECT 58.370 40.280 58.680 40.290 ;
        RECT 76.680 40.280 76.990 40.290 ;
        RECT 51.030 40.100 51.350 40.150 ;
        RECT 53.440 40.100 53.760 40.120 ;
        RECT 51.030 40.080 53.760 40.100 ;
        RECT 55.770 40.100 79.160 40.280 ;
        RECT 79.400 40.240 79.960 40.510 ;
        RECT 80.400 40.440 80.710 40.510 ;
        RECT 81.370 40.440 81.680 40.520 ;
        RECT 83.620 40.440 83.930 40.540 ;
        RECT 81.370 40.210 83.930 40.440 ;
        RECT 81.370 40.190 81.680 40.210 ;
        RECT 55.770 40.080 55.950 40.100 ;
        RECT 51.030 39.920 55.950 40.080 ;
        RECT 58.370 39.960 58.680 40.100 ;
        RECT 76.680 39.960 76.990 40.100 ;
        RECT 51.030 39.910 53.760 39.920 ;
        RECT 51.030 39.830 51.350 39.910 ;
        RECT 53.440 39.860 53.760 39.910 ;
        RECT 80.550 39.900 80.860 39.940 ;
        RECT 80.370 39.790 81.090 39.900 ;
        RECT 81.320 39.790 81.630 39.870 ;
        RECT 43.040 39.550 45.480 39.770 ;
        RECT 65.480 39.700 65.790 39.740 ;
        RECT 65.100 39.680 65.940 39.700 ;
        RECT 49.790 39.610 50.270 39.620 ;
        RECT 43.140 38.750 43.400 39.550 ;
        RECT 45.140 39.490 45.480 39.550 ;
        RECT 49.660 39.320 50.270 39.610 ;
        RECT 65.100 39.500 67.730 39.680 ;
        RECT 80.370 39.650 81.630 39.790 ;
        RECT 80.550 39.610 81.630 39.650 ;
        RECT 80.820 39.580 81.630 39.610 ;
        RECT 80.820 39.540 81.090 39.580 ;
        RECT 81.320 39.540 81.630 39.580 ;
        RECT 65.480 39.410 65.790 39.500 ;
        RECT 49.660 39.170 49.980 39.320 ;
        RECT 58.220 39.260 58.530 39.330 ;
        RECT 56.200 39.250 58.530 39.260 ;
        RECT 76.830 39.260 77.140 39.330 ;
        RECT 79.430 39.260 79.740 39.400 ;
        RECT 46.840 39.030 47.160 39.050 ;
        RECT 46.830 38.980 47.160 39.030 ;
        RECT 47.870 38.980 48.190 38.990 ;
        RECT 49.660 38.980 49.860 39.170 ;
        RECT 56.200 39.040 75.690 39.250 ;
        RECT 57.510 39.030 75.690 39.040 ;
        RECT 58.220 39.000 58.530 39.030 ;
        RECT 46.830 38.780 49.860 38.980 ;
        RECT 46.830 38.770 47.160 38.780 ;
        RECT 46.840 38.760 47.160 38.770 ;
        RECT 47.870 38.730 48.190 38.780 ;
        RECT 49.930 38.280 50.270 38.350 ;
        RECT 49.790 38.230 50.270 38.280 ;
        RECT 49.590 38.050 50.270 38.230 ;
        RECT 57.270 38.060 74.510 38.280 ;
        RECT 43.040 37.800 45.480 38.020 ;
        RECT 43.140 37.000 43.400 37.800 ;
        RECT 45.140 37.740 45.480 37.800 ;
        RECT 46.840 37.280 47.160 37.300 ;
        RECT 46.830 37.230 47.160 37.280 ;
        RECT 47.870 37.230 48.190 37.240 ;
        RECT 49.590 37.230 49.770 38.050 ;
        RECT 57.270 37.920 57.590 38.060 ;
        RECT 51.030 37.760 51.350 37.840 ;
        RECT 53.440 37.780 53.760 37.810 ;
        RECT 53.440 37.760 56.050 37.780 ;
        RECT 51.030 37.600 56.050 37.760 ;
        RECT 51.030 37.570 53.760 37.600 ;
        RECT 51.030 37.520 51.350 37.570 ;
        RECT 53.440 37.550 53.760 37.570 ;
        RECT 46.830 37.030 49.780 37.230 ;
        RECT 46.830 37.020 47.160 37.030 ;
        RECT 46.840 37.010 47.160 37.020 ;
        RECT 47.870 36.980 48.190 37.030 ;
        RECT 55.870 35.410 56.050 37.600 ;
        RECT 57.290 37.580 57.550 37.920 ;
        RECT 57.270 37.320 57.590 37.580 ;
        RECT 58.220 36.500 58.530 36.570 ;
        RECT 56.200 36.290 71.210 36.500 ;
        RECT 57.510 36.280 71.210 36.290 ;
        RECT 58.220 36.240 58.530 36.280 ;
        RECT 65.510 35.990 65.820 36.050 ;
        RECT 65.050 35.980 65.820 35.990 ;
        RECT 65.050 35.970 65.940 35.980 ;
        RECT 65.050 35.760 67.730 35.970 ;
        RECT 70.990 35.950 71.210 36.280 ;
        RECT 74.290 36.450 74.510 38.060 ;
        RECT 75.470 37.830 75.690 39.030 ;
        RECT 76.830 39.070 79.740 39.260 ;
        RECT 76.830 39.040 79.430 39.070 ;
        RECT 76.830 39.000 77.140 39.040 ;
        RECT 80.890 38.970 81.090 38.980 ;
        RECT 81.320 38.970 81.630 39.010 ;
        RECT 80.890 38.890 81.630 38.970 ;
        RECT 80.600 38.870 81.630 38.890 ;
        RECT 80.550 38.760 81.630 38.870 ;
        RECT 80.550 38.630 81.110 38.760 ;
        RECT 81.320 38.680 81.630 38.760 ;
        RECT 80.550 38.620 81.020 38.630 ;
        RECT 81.370 38.300 81.680 38.360 ;
        RECT 83.670 38.300 83.980 38.320 ;
        RECT 84.810 38.300 85.040 40.780 ;
        RECT 106.550 40.680 110.960 40.780 ;
        RECT 108.310 40.670 109.430 40.680 ;
        RECT 109.080 40.550 109.390 40.670 ;
        RECT 110.650 40.550 110.960 40.680 ;
        RECT 80.440 38.120 81.060 38.220 ;
        RECT 80.160 38.080 81.060 38.120 ;
        RECT 79.840 37.840 81.060 38.080 ;
        RECT 81.370 38.070 85.040 38.300 ;
        RECT 85.650 38.170 89.290 38.370 ;
        RECT 89.660 38.190 106.850 38.370 ;
        RECT 109.080 38.200 109.390 38.320 ;
        RECT 108.310 38.190 109.430 38.200 ;
        RECT 110.650 38.190 110.960 38.320 ;
        RECT 89.660 38.170 110.960 38.190 ;
        RECT 81.370 38.030 81.680 38.070 ;
        RECT 83.670 37.990 83.980 38.070 ;
        RECT 75.440 37.790 75.690 37.830 ;
        RECT 80.160 37.790 81.060 37.840 ;
        RECT 75.440 37.150 75.700 37.790 ;
        RECT 80.440 37.690 81.060 37.790 ;
        RECT 81.370 37.470 81.680 37.520 ;
        RECT 83.660 37.470 83.970 37.600 ;
        RECT 85.650 37.470 85.850 38.170 ;
        RECT 106.590 37.990 110.960 38.170 ;
        RECT 108.310 37.980 109.430 37.990 ;
        RECT 81.370 37.320 85.850 37.470 ;
        RECT 81.370 37.250 85.820 37.320 ;
        RECT 81.370 37.190 81.680 37.250 ;
        RECT 75.440 36.940 79.570 37.150 ;
        RECT 79.360 36.800 79.570 36.940 ;
        RECT 81.320 36.800 81.630 36.870 ;
        RECT 79.360 36.590 81.630 36.800 ;
        RECT 81.020 36.580 81.630 36.590 ;
        RECT 76.830 36.500 77.140 36.570 ;
        RECT 81.320 36.540 81.630 36.580 ;
        RECT 76.830 36.450 79.160 36.500 ;
        RECT 74.290 36.290 79.160 36.450 ;
        RECT 74.290 36.230 77.140 36.290 ;
        RECT 81.320 36.000 81.630 36.010 ;
        RECT 75.360 35.950 81.630 36.000 ;
        RECT 70.990 35.790 81.630 35.950 ;
        RECT 65.050 35.740 65.940 35.760 ;
        RECT 65.510 35.720 65.820 35.740 ;
        RECT 70.990 35.730 75.750 35.790 ;
        RECT 81.020 35.760 81.630 35.790 ;
        RECT 81.320 35.680 81.630 35.760 ;
        RECT 58.370 35.410 58.680 35.550 ;
        RECT 55.870 35.400 58.680 35.410 ;
        RECT 76.680 35.410 76.990 35.550 ;
        RECT 76.680 35.400 79.160 35.410 ;
        RECT 55.870 35.250 79.160 35.400 ;
        RECT 55.870 35.230 58.680 35.250 ;
        RECT 58.370 35.220 58.680 35.230 ;
        RECT 76.680 35.230 79.160 35.250 ;
        RECT 81.370 35.310 81.680 35.360 ;
        RECT 83.580 35.310 83.890 35.350 ;
        RECT 76.680 35.220 76.990 35.230 ;
        RECT 81.370 35.080 84.080 35.310 ;
        RECT 81.370 35.030 81.680 35.080 ;
        RECT 83.580 35.020 83.890 35.080 ;
        RECT 43.040 32.920 45.480 33.140 ;
        RECT 43.140 32.120 43.400 32.920 ;
        RECT 45.140 32.860 45.480 32.920 ;
        RECT 51.010 32.830 51.330 32.880 ;
        RECT 53.420 32.830 53.740 32.850 ;
        RECT 51.010 32.810 55.490 32.830 ;
        RECT 55.790 32.810 55.970 32.820 ;
        RECT 51.010 32.700 55.970 32.810 ;
        RECT 59.770 32.700 60.080 32.840 ;
        RECT 75.260 32.700 75.570 32.840 ;
        RECT 51.010 32.660 77.730 32.700 ;
        RECT 51.010 32.640 53.740 32.660 ;
        RECT 51.010 32.560 51.330 32.640 ;
        RECT 53.420 32.590 53.740 32.640 ;
        RECT 55.450 32.630 77.730 32.660 ;
        RECT 55.790 32.520 77.730 32.630 ;
        RECT 59.770 32.510 60.080 32.520 ;
        RECT 75.260 32.510 75.570 32.520 ;
        RECT 46.840 32.400 47.160 32.420 ;
        RECT 46.830 32.350 47.160 32.400 ;
        RECT 47.870 32.350 48.190 32.360 ;
        RECT 46.830 32.150 50.250 32.350 ;
        RECT 77.580 32.320 78.140 32.500 ;
        RECT 59.770 32.270 60.080 32.290 ;
        RECT 75.260 32.270 75.570 32.290 ;
        RECT 46.830 32.140 47.160 32.150 ;
        RECT 46.840 32.130 47.160 32.140 ;
        RECT 47.870 32.100 48.190 32.150 ;
        RECT 49.770 32.120 50.250 32.150 ;
        RECT 49.910 32.050 50.250 32.120 ;
        RECT 57.610 32.260 60.170 32.270 ;
        RECT 75.170 32.260 77.730 32.270 ;
        RECT 57.610 32.090 77.730 32.260 ;
        RECT 59.770 32.080 75.570 32.090 ;
        RECT 59.770 31.960 60.080 32.080 ;
        RECT 75.260 31.960 75.570 32.080 ;
        RECT 43.040 31.170 45.480 31.390 ;
        RECT 43.140 30.370 43.400 31.170 ;
        RECT 45.140 31.110 45.480 31.170 ;
        RECT 49.910 31.010 50.250 31.080 ;
        RECT 49.770 30.960 50.250 31.010 ;
        RECT 49.570 30.950 50.250 30.960 ;
        RECT 49.550 30.780 50.250 30.950 ;
        RECT 46.840 30.650 47.160 30.670 ;
        RECT 46.830 30.600 47.160 30.650 ;
        RECT 47.870 30.600 48.190 30.610 ;
        RECT 49.550 30.600 49.750 30.780 ;
        RECT 59.770 30.730 60.080 30.740 ;
        RECT 75.260 30.730 75.570 30.740 ;
        RECT 46.830 30.400 49.750 30.600 ;
        RECT 55.530 30.570 77.730 30.730 ;
        RECT 51.010 30.490 51.330 30.570 ;
        RECT 53.490 30.550 77.730 30.570 ;
        RECT 53.490 30.540 55.710 30.550 ;
        RECT 53.420 30.490 55.710 30.540 ;
        RECT 51.010 30.410 55.710 30.490 ;
        RECT 59.770 30.410 60.080 30.550 ;
        RECT 75.260 30.410 75.570 30.550 ;
        RECT 94.880 30.500 95.480 30.560 ;
        RECT 117.600 30.500 118.500 31.530 ;
        RECT 46.830 30.390 47.160 30.400 ;
        RECT 46.840 30.380 47.160 30.390 ;
        RECT 47.870 30.350 48.190 30.400 ;
        RECT 51.010 30.300 53.740 30.410 ;
        RECT 54.220 30.400 55.710 30.410 ;
        RECT 54.920 30.390 55.710 30.400 ;
        RECT 51.010 30.250 51.330 30.300 ;
        RECT 53.420 30.280 53.740 30.300 ;
        RECT 94.880 30.030 118.500 30.500 ;
        RECT 94.880 29.980 95.480 30.030 ;
        RECT 43.040 29.420 45.480 29.640 ;
        RECT 43.140 28.620 43.400 29.420 ;
        RECT 45.140 29.360 45.480 29.420 ;
        RECT 51.010 29.630 51.330 29.680 ;
        RECT 53.420 29.630 53.740 29.650 ;
        RECT 51.010 29.610 53.740 29.630 ;
        RECT 51.010 29.600 55.730 29.610 ;
        RECT 51.010 29.460 55.740 29.600 ;
        RECT 59.770 29.460 60.080 29.600 ;
        RECT 75.260 29.460 75.570 29.600 ;
        RECT 51.010 29.450 77.730 29.460 ;
        RECT 51.010 29.440 53.740 29.450 ;
        RECT 51.010 29.360 51.330 29.440 ;
        RECT 53.420 29.390 53.740 29.440 ;
        RECT 55.560 29.280 77.730 29.450 ;
        RECT 117.600 29.440 118.500 30.030 ;
        RECT 59.770 29.270 60.080 29.280 ;
        RECT 75.260 29.270 75.570 29.280 ;
        RECT 49.770 29.130 50.250 29.150 ;
        RECT 46.840 28.900 47.160 28.920 ;
        RECT 46.830 28.850 47.160 28.900 ;
        RECT 47.870 28.850 48.190 28.860 ;
        RECT 49.500 28.850 50.250 29.130 ;
        RECT 59.770 29.030 60.080 29.050 ;
        RECT 75.260 29.030 75.570 29.050 ;
        RECT 57.610 28.850 77.730 29.030 ;
        RECT 46.830 28.800 49.990 28.850 ;
        RECT 46.830 28.650 49.850 28.800 ;
        RECT 59.770 28.720 60.080 28.850 ;
        RECT 75.260 28.720 75.570 28.850 ;
        RECT 46.830 28.640 47.160 28.650 ;
        RECT 46.840 28.630 47.160 28.640 ;
        RECT 47.870 28.600 48.190 28.650 ;
        RECT 59.770 27.930 60.080 28.060 ;
        RECT 75.260 27.930 75.570 28.060 ;
        RECT 43.040 27.670 45.480 27.890 ;
        RECT 49.910 27.810 50.250 27.880 ;
        RECT 43.140 26.870 43.400 27.670 ;
        RECT 45.140 27.610 45.480 27.670 ;
        RECT 49.540 27.580 50.250 27.810 ;
        RECT 57.610 27.750 77.730 27.930 ;
        RECT 59.770 27.730 60.080 27.750 ;
        RECT 75.260 27.730 75.570 27.750 ;
        RECT 46.840 27.150 47.160 27.170 ;
        RECT 46.830 27.100 47.160 27.150 ;
        RECT 47.870 27.100 48.190 27.110 ;
        RECT 49.540 27.100 49.740 27.580 ;
        RECT 59.770 27.500 60.080 27.510 ;
        RECT 75.260 27.500 75.570 27.510 ;
        RECT 46.830 26.900 49.740 27.100 ;
        RECT 51.010 27.290 51.330 27.370 ;
        RECT 53.420 27.310 53.740 27.340 ;
        RECT 55.530 27.330 77.730 27.500 ;
        RECT 55.530 27.320 60.080 27.330 ;
        RECT 55.540 27.310 55.720 27.320 ;
        RECT 53.420 27.290 55.720 27.310 ;
        RECT 51.010 27.130 55.720 27.290 ;
        RECT 59.770 27.180 60.080 27.320 ;
        RECT 75.260 27.320 77.730 27.330 ;
        RECT 75.260 27.180 75.570 27.320 ;
        RECT 51.010 27.100 53.740 27.130 ;
        RECT 51.010 27.050 51.330 27.100 ;
        RECT 53.420 27.080 53.740 27.100 ;
        RECT 46.830 26.890 47.160 26.900 ;
        RECT 46.840 26.880 47.160 26.890 ;
        RECT 47.870 26.850 48.190 26.900 ;
        RECT 43.000 23.860 45.440 24.080 ;
        RECT 43.100 23.060 43.360 23.860 ;
        RECT 45.100 23.800 45.440 23.860 ;
        RECT 51.040 23.560 51.360 23.610 ;
        RECT 53.450 23.560 53.770 23.580 ;
        RECT 51.040 23.550 55.520 23.560 ;
        RECT 51.040 23.390 55.650 23.550 ;
        RECT 51.040 23.370 53.770 23.390 ;
        RECT 55.340 23.370 55.650 23.390 ;
        RECT 59.800 23.370 60.110 23.510 ;
        RECT 46.800 23.340 47.120 23.360 ;
        RECT 46.790 23.290 47.120 23.340 ;
        RECT 47.830 23.290 48.150 23.300 ;
        RECT 51.040 23.290 51.360 23.370 ;
        RECT 53.450 23.320 53.770 23.370 ;
        RECT 46.790 23.090 49.870 23.290 ;
        RECT 55.470 23.190 60.110 23.370 ;
        RECT 59.800 23.180 60.110 23.190 ;
        RECT 60.400 23.350 60.720 23.370 ;
        RECT 60.400 23.160 68.320 23.350 ;
        RECT 68.480 23.160 68.790 23.200 ;
        RECT 60.400 23.140 68.790 23.160 ;
        RECT 60.400 23.110 60.720 23.140 ;
        RECT 46.790 23.080 47.120 23.090 ;
        RECT 46.800 23.070 47.120 23.080 ;
        RECT 47.830 23.040 48.150 23.090 ;
        RECT 49.670 23.080 49.870 23.090 ;
        RECT 49.670 22.850 50.280 23.080 ;
        RECT 68.110 22.950 68.790 23.140 ;
        RECT 68.480 22.870 68.790 22.950 ;
        RECT 49.940 22.780 50.280 22.850 ;
        RECT 57.130 22.710 57.280 22.730 ;
        RECT 56.110 22.560 57.280 22.710 ;
        RECT 43.000 22.110 45.440 22.330 ;
        RECT 56.050 22.230 56.330 22.560 ;
        RECT 57.130 22.310 57.280 22.560 ;
        RECT 60.380 22.310 60.700 22.320 ;
        RECT 57.130 22.160 60.700 22.310 ;
        RECT 43.100 21.310 43.360 22.110 ;
        RECT 45.100 22.050 45.440 22.110 ;
        RECT 60.260 22.060 60.700 22.160 ;
        RECT 49.940 21.740 50.280 21.810 ;
        RECT 49.800 21.700 50.280 21.740 ;
        RECT 46.800 21.590 47.120 21.610 ;
        RECT 46.790 21.540 47.120 21.590 ;
        RECT 47.830 21.540 48.150 21.550 ;
        RECT 49.660 21.540 50.280 21.700 ;
        RECT 57.110 21.560 57.430 21.830 ;
        RECT 46.790 21.510 50.280 21.540 ;
        RECT 46.790 21.340 49.980 21.510 ;
        RECT 59.800 21.420 60.110 21.430 ;
        RECT 46.790 21.330 47.120 21.340 ;
        RECT 46.800 21.320 47.120 21.330 ;
        RECT 47.830 21.290 48.150 21.340 ;
        RECT 55.450 21.300 60.110 21.420 ;
        RECT 51.040 21.220 51.360 21.300 ;
        RECT 53.520 21.270 60.110 21.300 ;
        RECT 53.450 21.260 60.110 21.270 ;
        RECT 53.450 21.240 60.200 21.260 ;
        RECT 53.450 21.220 55.630 21.240 ;
        RECT 51.040 21.140 55.630 21.220 ;
        RECT 51.040 21.030 53.770 21.140 ;
        RECT 54.250 21.130 55.630 21.140 ;
        RECT 54.950 21.120 55.630 21.130 ;
        RECT 51.040 20.980 51.360 21.030 ;
        RECT 53.450 21.010 53.770 21.030 ;
        RECT 55.310 21.090 55.630 21.120 ;
        RECT 59.800 21.120 60.200 21.240 ;
        RECT 59.800 21.100 60.110 21.120 ;
        RECT 55.310 21.010 55.490 21.090 ;
        RECT 60.340 21.080 60.570 21.090 ;
        RECT 60.340 21.050 67.910 21.080 ;
        RECT 60.340 20.880 67.970 21.050 ;
        RECT 68.480 20.880 68.790 20.960 ;
        RECT 57.090 20.780 57.410 20.810 ;
        RECT 60.340 20.780 60.580 20.880 ;
        RECT 57.090 20.600 60.580 20.780 ;
        RECT 67.780 20.680 68.790 20.880 ;
        RECT 68.380 20.670 68.790 20.680 ;
        RECT 68.480 20.630 68.790 20.670 ;
        RECT 57.090 20.580 60.500 20.600 ;
        RECT 43.000 20.360 45.440 20.580 ;
        RECT 57.090 20.550 57.410 20.580 ;
        RECT 43.100 19.560 43.360 20.360 ;
        RECT 45.100 20.300 45.440 20.360 ;
        RECT 51.040 20.360 51.360 20.410 ;
        RECT 60.380 20.400 60.700 20.440 ;
        RECT 60.380 20.380 67.930 20.400 ;
        RECT 68.480 20.390 68.790 20.430 ;
        RECT 68.380 20.380 68.790 20.390 ;
        RECT 53.450 20.360 53.770 20.380 ;
        RECT 51.040 20.340 53.770 20.360 ;
        RECT 51.040 20.180 55.560 20.340 ;
        RECT 51.040 20.170 53.770 20.180 ;
        RECT 51.040 20.090 51.360 20.170 ;
        RECT 53.450 20.120 53.770 20.170 ;
        RECT 55.380 20.130 55.560 20.180 ;
        RECT 59.800 20.140 60.110 20.270 ;
        RECT 60.380 20.180 68.790 20.380 ;
        RECT 60.480 20.170 60.800 20.180 ;
        RECT 59.800 20.130 60.230 20.140 ;
        RECT 55.380 19.970 60.230 20.130 ;
        RECT 68.480 20.100 68.790 20.180 ;
        RECT 92.670 20.140 93.220 20.150 ;
        RECT 92.670 20.120 93.230 20.140 ;
        RECT 117.600 20.120 118.500 21.270 ;
        RECT 55.380 19.950 60.110 19.970 ;
        RECT 59.800 19.940 60.110 19.950 ;
        RECT 46.800 19.840 47.120 19.860 ;
        RECT 46.790 19.790 47.120 19.840 ;
        RECT 47.830 19.790 48.150 19.800 ;
        RECT 49.800 19.790 50.280 19.880 ;
        RECT 46.790 19.590 50.280 19.790 ;
        RECT 46.790 19.580 47.120 19.590 ;
        RECT 46.800 19.570 47.120 19.580 ;
        RECT 47.830 19.540 48.150 19.590 ;
        RECT 49.740 19.580 50.280 19.590 ;
        RECT 56.660 19.720 56.980 19.760 ;
        RECT 49.740 19.500 50.030 19.580 ;
        RECT 56.660 19.440 57.270 19.720 ;
        RECT 59.800 19.700 60.110 19.720 ;
        RECT 57.640 19.530 66.940 19.700 ;
        RECT 92.670 19.650 118.500 20.120 ;
        RECT 92.670 19.640 93.230 19.650 ;
        RECT 92.670 19.620 93.220 19.640 ;
        RECT 57.640 19.520 60.200 19.530 ;
        RECT 57.070 19.220 57.270 19.440 ;
        RECT 59.800 19.390 60.110 19.520 ;
        RECT 60.250 19.220 60.570 19.260 ;
        RECT 57.070 19.020 60.620 19.220 ;
        RECT 117.600 19.180 118.500 19.650 ;
        RECT 60.250 19.000 60.570 19.020 ;
        RECT 43.000 18.610 45.440 18.830 ;
        RECT 49.720 18.620 50.020 18.660 ;
        RECT 43.100 17.810 43.360 18.610 ;
        RECT 45.100 18.550 45.440 18.610 ;
        RECT 49.710 18.610 50.020 18.620 ;
        RECT 49.710 18.310 50.280 18.610 ;
        RECT 57.040 18.480 57.350 18.810 ;
        RECT 46.800 18.090 47.120 18.110 ;
        RECT 46.790 18.040 47.120 18.090 ;
        RECT 47.830 18.040 48.150 18.050 ;
        RECT 49.710 18.040 49.910 18.310 ;
        RECT 59.800 18.170 60.110 18.180 ;
        RECT 46.790 17.840 49.910 18.040 ;
        RECT 51.040 18.020 51.360 18.100 ;
        RECT 53.450 18.040 53.770 18.070 ;
        RECT 55.620 18.040 60.110 18.170 ;
        RECT 68.480 18.130 68.790 18.190 ;
        RECT 67.930 18.120 68.790 18.130 ;
        RECT 53.450 18.020 60.110 18.040 ;
        RECT 51.040 17.990 60.110 18.020 ;
        RECT 51.040 17.860 55.800 17.990 ;
        RECT 46.790 17.830 47.120 17.840 ;
        RECT 46.800 17.820 47.120 17.830 ;
        RECT 47.830 17.790 48.150 17.840 ;
        RECT 51.040 17.830 53.770 17.860 ;
        RECT 59.800 17.850 60.110 17.990 ;
        RECT 60.350 17.900 68.790 18.120 ;
        RECT 60.350 17.890 67.940 17.900 ;
        RECT 60.350 17.880 61.120 17.890 ;
        RECT 51.040 17.780 51.360 17.830 ;
        RECT 53.450 17.810 53.770 17.830 ;
        RECT 57.090 17.840 57.400 17.850 ;
        RECT 57.090 17.710 57.450 17.840 ;
        RECT 60.350 17.710 60.590 17.880 ;
        RECT 68.480 17.860 68.790 17.900 ;
        RECT 57.090 17.470 60.590 17.710 ;
        RECT 49.450 17.340 49.770 17.390 ;
        RECT 56.060 17.340 56.380 17.440 ;
        RECT 49.450 17.180 56.380 17.340 ;
        RECT 49.450 17.130 49.770 17.180 ;
        RECT 56.060 17.160 56.380 17.180 ;
        RECT 57.090 17.340 57.410 17.470 ;
        RECT 67.710 17.340 68.120 17.450 ;
        RECT 57.090 17.180 68.120 17.340 ;
        RECT 57.090 17.150 57.410 17.180 ;
        RECT 56.650 17.100 56.930 17.110 ;
        RECT 56.630 17.010 56.950 17.100 ;
        RECT 67.710 17.080 68.120 17.180 ;
        RECT 58.870 17.010 59.190 17.040 ;
        RECT 56.600 16.850 59.190 17.010 ;
        RECT 56.630 16.840 56.950 16.850 ;
        RECT 56.650 16.830 56.930 16.840 ;
        RECT 58.870 16.780 59.190 16.850 ;
        RECT 58.890 16.770 59.170 16.780 ;
        RECT 57.670 15.860 58.050 15.890 ;
        RECT 59.020 15.880 62.080 15.890 ;
        RECT 49.210 15.850 52.270 15.860 ;
        RECT 49.120 15.520 52.270 15.850 ;
        RECT 54.770 15.520 58.050 15.860 ;
        RECT 58.930 15.800 62.080 15.880 ;
        RECT 49.120 14.840 49.440 15.520 ;
        RECT 51.940 15.510 52.250 15.520 ;
        RECT 54.790 15.510 55.100 15.520 ;
        RECT 48.970 14.460 49.440 14.840 ;
        RECT 49.120 13.070 49.440 14.460 ;
        RECT 57.600 15.500 58.050 15.520 ;
        RECT 58.820 15.550 62.080 15.800 ;
        RECT 64.580 15.880 67.640 15.890 ;
        RECT 64.580 15.660 67.730 15.880 ;
        RECT 64.580 15.550 68.070 15.660 ;
        RECT 57.600 13.070 57.920 15.500 ;
        RECT 58.820 15.460 59.250 15.550 ;
        RECT 61.750 15.540 62.060 15.550 ;
        RECT 64.600 15.540 64.910 15.550 ;
        RECT 49.120 12.740 52.280 13.070 ;
        RECT 54.760 12.740 57.920 13.070 ;
        RECT 49.120 11.700 49.440 12.740 ;
        RECT 57.600 11.700 57.920 12.740 ;
        RECT 49.120 11.380 52.280 11.700 ;
        RECT 54.760 11.380 57.920 11.700 ;
        RECT 58.930 13.100 59.250 15.460 ;
        RECT 67.410 15.300 68.070 15.550 ;
        RECT 67.410 13.100 67.730 15.300 ;
        RECT 70.890 15.160 71.200 15.170 ;
        RECT 71.980 15.160 72.290 15.190 ;
        RECT 69.340 15.010 72.290 15.160 ;
        RECT 69.160 14.860 72.290 15.010 ;
        RECT 69.160 14.820 70.090 14.860 ;
        RECT 70.890 14.840 71.200 14.860 ;
        RECT 69.160 14.690 69.720 14.820 ;
        RECT 69.160 14.580 69.690 14.690 ;
        RECT 58.930 12.770 62.090 13.100 ;
        RECT 64.570 12.770 67.730 13.100 ;
        RECT 58.930 11.730 59.250 12.770 ;
        RECT 67.410 11.730 67.730 12.770 ;
        RECT 58.930 11.410 62.090 11.730 ;
        RECT 64.570 11.410 67.730 11.730 ;
        RECT 69.340 13.820 69.690 14.580 ;
        RECT 69.340 13.490 72.290 13.820 ;
        RECT 59.550 11.400 59.860 11.410 ;
        RECT 60.650 11.400 60.960 11.410 ;
        RECT 61.750 11.400 62.060 11.410 ;
        RECT 64.600 11.400 64.910 11.410 ;
        RECT 65.700 11.400 66.010 11.410 ;
        RECT 66.800 11.400 67.110 11.410 ;
        RECT 49.740 11.370 50.050 11.380 ;
        RECT 50.840 11.370 51.150 11.380 ;
        RECT 51.940 11.370 52.250 11.380 ;
        RECT 54.790 11.370 55.100 11.380 ;
        RECT 55.890 11.370 56.200 11.380 ;
        RECT 56.990 11.370 57.300 11.380 ;
        RECT 48.880 10.590 49.480 11.080 ;
        RECT 58.690 10.620 59.290 11.110 ;
        RECT 69.340 11.050 69.690 13.490 ;
        RECT 69.340 11.040 72.280 11.050 ;
        RECT 69.340 10.730 72.290 11.040 ;
        RECT 69.570 10.720 72.290 10.730 ;
        RECT 70.890 10.710 71.200 10.720 ;
        RECT 71.980 10.710 72.290 10.720 ;
        RECT 48.880 10.260 49.490 10.590 ;
        RECT 58.690 10.290 59.300 10.620 ;
        RECT 49.060 9.230 49.560 9.240 ;
        RECT 94.990 9.230 95.550 9.250 ;
        RECT 49.060 8.770 95.550 9.230 ;
        RECT 49.060 8.710 49.580 8.770 ;
        RECT 94.990 8.750 95.550 8.770 ;
        RECT 49.060 8.690 49.560 8.710 ;
        RECT 58.810 7.340 93.360 7.410 ;
        RECT 58.800 6.950 93.360 7.340 ;
        RECT 58.800 6.820 59.450 6.950 ;
        RECT 92.670 6.930 93.230 6.950 ;
        RECT 2.770 -2.960 4.040 -1.080 ;
        RECT 2.840 -7.710 4.110 -5.830 ;
        RECT 106.780 -6.260 107.100 -5.940 ;
        RECT 107.720 -6.260 108.040 -5.940 ;
      LAYER via2 ;
        RECT 79.480 47.310 79.800 47.630 ;
        RECT 80.510 47.300 80.830 47.620 ;
        RECT 80.590 43.820 80.930 44.160 ;
        RECT 79.520 40.340 79.850 40.690 ;
        RECT 80.610 37.770 80.950 38.130 ;
  END
END sky130_hilas_TopLevelTextStructure

MACRO sky130_hilas_capacitorArray01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_capacitorArray01 ;
  ORIGIN 13.040 0.790 ;
  SIZE 36.700 BY 6.500 ;
  PIN CAPTERM2
    USE ANALOG ;
    PORT
      LAYER met3 ;
        RECT 22.190 1.630 23.340 3.270 ;
        RECT 22.640 1.620 23.340 1.630 ;
    END
  END CAPTERM2
  PIN CAPTERM1
    USE ANALOG ;
    ANTENNAGATEAREA 0.720000 ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met3 ;
        RECT -1.790 5.170 -1.410 5.460 ;
        RECT -1.870 3.920 -1.330 5.170 ;
    END
  END CAPTERM1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -5.520 5.480 -2.960 5.710 ;
        RECT -5.520 -0.560 22.380 5.480 ;
        RECT -5.520 -0.790 -2.960 -0.560 ;
        RECT -1.040 -0.570 22.380 -0.560 ;
      LAYER met1 ;
        RECT -3.480 5.000 -3.320 5.700 ;
        RECT -3.590 4.450 -3.320 5.000 ;
        RECT -3.590 4.400 -3.310 4.450 ;
        RECT -3.480 4.310 -3.310 4.400 ;
        RECT -3.480 3.840 -3.320 4.310 ;
        RECT -3.480 3.750 -3.310 3.840 ;
        RECT -3.590 3.700 -3.310 3.750 ;
        RECT -3.590 3.150 -3.320 3.700 ;
        RECT -3.480 1.760 -3.320 3.150 ;
        RECT -3.590 1.210 -3.320 1.760 ;
        RECT -3.590 1.160 -3.310 1.210 ;
        RECT -3.480 1.070 -3.310 1.160 ;
        RECT -3.480 0.610 -3.320 1.070 ;
        RECT -3.480 0.520 -3.310 0.610 ;
        RECT -3.590 0.470 -3.310 0.520 ;
        RECT -3.590 -0.080 -3.320 0.470 ;
        RECT -3.480 -0.780 -3.320 -0.080 ;
    END
  END VINJ
  PIN GATESELECT
    ANTENNAGATEAREA 0.720000 ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met2 ;
        RECT -2.300 5.450 -1.790 5.480 ;
        RECT -4.370 5.360 -4.050 5.430 ;
        RECT -2.300 5.360 -1.370 5.450 ;
        RECT -4.370 5.170 -1.370 5.360 ;
        RECT -1.870 5.150 -1.370 5.170 ;
      LAYER via2 ;
        RECT -1.740 5.150 -1.460 5.430 ;
    END
  END GATESELECT
  PIN VTUN
    ANTENNADIFFAREA 2.237600 ;
    PORT
      LAYER nwell ;
        RECT -13.030 3.120 -11.300 5.700 ;
        RECT -13.040 2.940 -11.300 3.120 ;
        RECT -13.030 -0.790 -11.300 2.940 ;
      LAYER met1 ;
        RECT -12.680 -0.790 -12.280 5.710 ;
    END
  END VTUN
  PIN GATE
    USE ANALOG ;
    ANTENNADIFFAREA 3.253900 ;
    PORT
      LAYER nwell ;
        RECT -9.280 -0.790 -7.050 5.700 ;
      LAYER met1 ;
        RECT -8.630 3.560 -8.250 5.710 ;
        RECT -8.640 1.700 -8.250 3.560 ;
        RECT -8.630 -0.420 -8.250 1.700 ;
        RECT -8.640 -0.570 -8.250 -0.420 ;
        RECT -8.630 -0.790 -8.250 -0.570 ;
    END
  END GATE
  PIN DRAIN2
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT -5.430 3.180 -5.120 3.190 ;
        RECT -13.030 3.120 -2.960 3.180 ;
        RECT 22.650 3.120 23.660 3.130 ;
        RECT -13.040 3.000 23.660 3.120 ;
        RECT -13.040 2.940 -12.920 3.000 ;
        RECT -5.430 2.860 -5.120 3.000 ;
        RECT -4.100 2.940 23.660 3.000 ;
    END
  END DRAIN2
  PIN DRAIN1
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT -5.430 5.150 -5.120 5.290 ;
        RECT -13.030 4.980 -2.960 5.150 ;
        RECT -13.030 4.970 23.660 4.980 ;
        RECT -13.030 4.800 -12.920 4.970 ;
        RECT -5.430 4.960 -5.120 4.970 ;
        RECT -4.060 4.800 23.660 4.970 ;
    END
  END DRAIN1
  PIN DRAIN4
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT -13.020 -0.050 -12.920 0.120 ;
        RECT -5.430 -0.050 -5.120 -0.040 ;
        RECT -4.230 -0.050 23.660 0.120 ;
        RECT -13.030 -0.220 -2.960 -0.050 ;
        RECT -5.430 -0.230 -2.960 -0.220 ;
        RECT -5.430 -0.370 -5.120 -0.230 ;
    END
  END DRAIN4
  PIN DRAIN3
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT -13.020 1.910 -12.920 1.960 ;
        RECT -5.430 1.910 -5.120 2.050 ;
        RECT -4.270 1.910 23.660 1.960 ;
        RECT -13.030 1.790 23.660 1.910 ;
        RECT -13.030 1.730 -2.960 1.790 ;
        RECT -5.430 1.720 -5.120 1.730 ;
    END
  END DRAIN3
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT -10.280 0.990 -9.960 1.000 ;
        RECT -6.350 0.990 -6.030 1.050 ;
        RECT -10.280 0.810 -6.030 0.990 ;
        RECT -10.280 0.740 -9.960 0.810 ;
        RECT -6.350 0.760 -6.030 0.810 ;
    END
    PORT
      LAYER met1 ;
        RECT -6.310 4.320 -6.070 5.710 ;
        RECT -6.330 3.660 -6.060 4.320 ;
        RECT -6.310 1.070 -6.070 3.660 ;
        RECT -6.320 0.750 -6.060 1.070 ;
        RECT -6.310 -0.790 -6.070 0.750 ;
      LAYER via ;
        RECT -6.320 0.780 -6.060 1.040 ;
    END
    PORT
      LAYER met1 ;
        RECT -10.240 4.300 -10.000 5.710 ;
        RECT -10.250 3.640 -9.990 4.300 ;
        RECT -10.240 1.030 -10.000 3.640 ;
        RECT -10.250 0.710 -9.990 1.030 ;
        RECT -10.240 -0.790 -10.000 0.710 ;
      LAYER via ;
        RECT -10.250 0.740 -9.990 1.000 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT -5.420 5.240 -5.100 5.250 ;
        RECT -5.420 5.070 -4.840 5.240 ;
        RECT -5.420 5.020 -5.090 5.070 ;
        RECT -5.420 4.990 -5.100 5.020 ;
        RECT -3.560 4.970 -3.360 5.320 ;
        RECT -5.420 4.660 -5.100 4.700 ;
        RECT -5.420 4.620 -5.090 4.660 ;
        RECT -5.420 4.450 -4.840 4.620 ;
        RECT -5.420 4.440 -5.100 4.450 ;
        RECT -4.290 4.350 -4.090 4.950 ;
        RECT -3.560 4.940 -3.350 4.970 ;
        RECT -3.570 4.350 -3.350 4.940 ;
        RECT -10.210 3.730 -10.040 4.260 ;
        RECT -6.270 3.720 -6.100 4.250 ;
        RECT -5.420 3.700 -5.100 3.710 ;
        RECT -5.420 3.530 -4.840 3.700 ;
        RECT -5.420 3.490 -5.090 3.530 ;
        RECT -5.420 3.450 -5.100 3.490 ;
        RECT -4.290 3.200 -4.090 3.800 ;
        RECT -3.570 3.210 -3.350 3.800 ;
        RECT -3.560 3.180 -3.350 3.210 ;
        RECT -5.420 3.130 -5.100 3.160 ;
        RECT -5.420 3.080 -5.090 3.130 ;
        RECT -12.610 2.230 -12.060 2.660 ;
        RECT -10.200 2.020 -10.030 3.030 ;
        RECT -5.420 2.910 -4.840 3.080 ;
        RECT -5.420 2.900 -5.100 2.910 ;
        RECT -8.580 2.160 -8.030 2.590 ;
        RECT -6.270 1.880 -6.100 2.890 ;
        RECT -3.560 2.830 -3.360 3.180 ;
        RECT -4.170 2.370 -3.730 2.540 ;
        RECT -5.420 2.000 -5.100 2.010 ;
        RECT -5.420 1.830 -4.840 2.000 ;
        RECT -5.420 1.780 -5.090 1.830 ;
        RECT -5.420 1.750 -5.100 1.780 ;
        RECT -3.560 1.730 -3.360 2.080 ;
        RECT -5.420 1.420 -5.100 1.460 ;
        RECT -5.420 1.380 -5.090 1.420 ;
        RECT -5.420 1.210 -4.840 1.380 ;
        RECT -5.420 1.200 -5.100 1.210 ;
        RECT -4.290 1.110 -4.090 1.710 ;
        RECT -3.560 1.700 -3.350 1.730 ;
        RECT -3.570 1.110 -3.350 1.700 ;
        RECT -5.420 0.470 -5.100 0.480 ;
        RECT -5.420 0.300 -4.840 0.470 ;
        RECT -5.420 0.260 -5.090 0.300 ;
        RECT -5.420 0.220 -5.100 0.260 ;
        RECT -4.290 -0.030 -4.090 0.570 ;
        RECT -3.570 -0.020 -3.350 0.570 ;
        RECT -3.560 -0.050 -3.350 -0.020 ;
        RECT -5.420 -0.100 -5.100 -0.070 ;
        RECT -5.420 -0.150 -5.090 -0.100 ;
        RECT -5.420 -0.320 -4.840 -0.150 ;
        RECT -5.420 -0.330 -5.100 -0.320 ;
        RECT -3.560 -0.400 -3.360 -0.050 ;
      LAYER mcon ;
        RECT -5.360 5.030 -5.190 5.200 ;
        RECT -4.280 4.740 -4.110 4.910 ;
        RECT -5.360 4.480 -5.190 4.650 ;
        RECT -3.550 4.770 -3.380 4.940 ;
        RECT -10.210 4.090 -10.040 4.260 ;
        RECT -6.270 4.080 -6.100 4.250 ;
        RECT -5.360 3.500 -5.190 3.670 ;
        RECT -4.280 3.240 -4.110 3.410 ;
        RECT -3.550 3.210 -3.380 3.380 ;
        RECT -5.360 2.950 -5.190 3.120 ;
        RECT -12.610 2.310 -12.340 2.580 ;
        RECT -10.200 2.630 -10.030 2.800 ;
        RECT -10.200 2.270 -10.030 2.440 ;
        RECT -8.580 2.240 -8.310 2.510 ;
        RECT -6.270 2.490 -6.100 2.660 ;
        RECT -3.910 2.370 -3.730 2.540 ;
        RECT -6.270 2.130 -6.100 2.300 ;
        RECT -5.360 1.790 -5.190 1.960 ;
        RECT -4.280 1.500 -4.110 1.670 ;
        RECT -5.360 1.240 -5.190 1.410 ;
        RECT -3.550 1.530 -3.380 1.700 ;
        RECT -5.360 0.270 -5.190 0.440 ;
        RECT -4.280 0.010 -4.110 0.180 ;
        RECT -3.550 -0.020 -3.380 0.150 ;
        RECT -5.360 -0.280 -5.190 -0.110 ;
      LAYER met1 ;
        RECT -4.290 5.460 -4.130 5.700 ;
        RECT -5.430 4.960 -5.110 5.280 ;
        RECT -4.340 5.140 -4.080 5.460 ;
        RECT -4.290 4.970 -4.130 5.140 ;
        RECT -4.290 4.950 -4.090 4.970 ;
        RECT -5.430 4.410 -5.110 4.730 ;
        RECT -4.310 4.710 -4.080 4.950 ;
        RECT -4.290 4.660 -4.080 4.710 ;
        RECT -3.920 4.660 -3.730 5.650 ;
        RECT -5.430 3.420 -5.110 3.740 ;
        RECT -4.290 3.490 -4.130 4.660 ;
        RECT -3.900 4.540 -3.730 4.660 ;
        RECT -3.890 3.610 -3.730 4.540 ;
        RECT -3.900 3.490 -3.730 3.610 ;
        RECT -4.290 3.440 -4.080 3.490 ;
        RECT -4.310 3.200 -4.080 3.440 ;
        RECT -5.430 2.870 -5.110 3.190 ;
        RECT -4.290 3.180 -4.090 3.200 ;
        RECT -4.290 2.550 -4.130 3.180 ;
        RECT -3.920 2.570 -3.730 3.490 ;
        RECT -3.940 2.550 -3.700 2.570 ;
        RECT -4.290 2.360 -3.700 2.550 ;
        RECT -5.430 1.720 -5.110 2.040 ;
        RECT -4.290 1.730 -4.130 2.360 ;
        RECT -3.940 2.340 -3.700 2.360 ;
        RECT -4.290 1.710 -4.090 1.730 ;
        RECT -5.430 1.170 -5.110 1.490 ;
        RECT -4.310 1.470 -4.080 1.710 ;
        RECT -4.290 1.420 -4.080 1.470 ;
        RECT -3.920 1.420 -3.730 2.340 ;
        RECT -5.430 0.190 -5.110 0.510 ;
        RECT -4.290 0.260 -4.130 1.420 ;
        RECT -3.900 1.300 -3.730 1.420 ;
        RECT -3.890 0.380 -3.730 1.300 ;
        RECT -3.900 0.260 -3.730 0.380 ;
        RECT -4.290 0.210 -4.080 0.260 ;
        RECT -4.310 -0.030 -4.080 0.210 ;
        RECT -5.430 -0.360 -5.110 -0.040 ;
        RECT -4.290 -0.050 -4.090 -0.030 ;
        RECT -4.290 -0.780 -4.130 -0.050 ;
        RECT -3.920 -0.730 -3.730 0.260 ;
      LAYER via ;
        RECT -5.400 4.990 -5.140 5.250 ;
        RECT -4.340 5.170 -4.080 5.430 ;
        RECT -5.400 4.440 -5.140 4.700 ;
        RECT -5.400 3.450 -5.140 3.710 ;
        RECT -5.400 2.900 -5.140 3.160 ;
        RECT -5.400 1.750 -5.140 2.010 ;
        RECT -5.400 1.200 -5.140 1.460 ;
        RECT -5.400 0.220 -5.140 0.480 ;
        RECT -5.400 -0.330 -5.140 -0.070 ;
      LAYER met2 ;
        RECT -5.430 4.720 -5.120 4.740 ;
        RECT -5.520 4.710 -2.960 4.720 ;
        RECT -13.030 4.550 -2.960 4.710 ;
        RECT -13.030 4.540 23.660 4.550 ;
        RECT -13.030 4.530 -5.120 4.540 ;
        RECT -5.430 4.410 -5.120 4.530 ;
        RECT -4.120 4.370 23.660 4.540 ;
        RECT -5.430 3.610 -5.120 3.740 ;
        RECT -3.160 3.610 -2.790 3.720 ;
        RECT -13.030 3.550 -2.790 3.610 ;
        RECT -13.030 3.430 23.660 3.550 ;
        RECT -5.430 3.410 -5.120 3.430 ;
        RECT -4.060 3.370 23.660 3.430 ;
        RECT -3.160 3.320 -2.790 3.370 ;
        RECT 22.970 2.220 23.660 2.630 ;
        RECT -3.200 1.540 -2.830 1.630 ;
        RECT -5.430 1.480 -5.120 1.500 ;
        RECT -4.170 1.480 23.660 1.540 ;
        RECT -13.030 1.370 23.660 1.480 ;
        RECT -13.030 1.300 -2.830 1.370 ;
        RECT -5.430 1.170 -5.120 1.300 ;
        RECT -3.200 1.230 -2.830 1.300 ;
        RECT -2.110 0.560 -1.740 0.760 ;
        RECT -5.430 0.380 -5.120 0.510 ;
        RECT -4.190 0.390 23.660 0.560 ;
        RECT -13.030 0.200 -2.960 0.380 ;
        RECT -2.110 0.360 -1.740 0.390 ;
        RECT -5.430 0.180 -5.120 0.200 ;
      LAYER via2 ;
        RECT -3.110 3.380 -2.830 3.660 ;
        RECT 23.040 2.280 23.330 2.560 ;
        RECT -3.150 1.290 -2.870 1.570 ;
        RECT -2.060 0.420 -1.780 0.700 ;
      LAYER met3 ;
        RECT -3.380 3.120 -2.590 3.870 ;
        RECT -3.420 1.730 -2.630 1.780 ;
        RECT -3.420 1.430 -2.490 1.730 ;
        RECT -3.420 1.030 -2.630 1.430 ;
        RECT -2.330 0.520 -1.540 0.910 ;
        RECT -2.330 0.220 -1.400 0.520 ;
        RECT -2.330 0.160 -1.540 0.220 ;
      LAYER via3 ;
        RECT -3.190 3.270 -2.760 3.750 ;
        RECT -3.230 1.180 -2.800 1.660 ;
        RECT -2.140 0.310 -1.710 0.790 ;
      LAYER met4 ;
        RECT -0.250 4.810 3.850 5.110 ;
        RECT -1.940 4.200 0.760 4.310 ;
        RECT -1.940 3.900 0.970 4.200 ;
        RECT -3.290 3.480 -2.630 3.840 ;
        RECT 0.460 3.560 0.970 3.900 ;
        RECT 3.470 3.610 3.850 4.810 ;
        RECT 6.310 3.640 9.590 3.940 ;
        RECT -3.290 3.180 -1.270 3.480 ;
        RECT -1.570 2.620 -1.270 3.180 ;
        RECT 6.310 2.620 6.610 3.640 ;
        RECT 9.290 2.620 9.590 3.640 ;
        RECT -1.570 2.320 9.590 2.620 ;
        RECT 11.990 3.620 20.880 3.920 ;
        RECT -3.330 1.730 -2.670 1.750 ;
        RECT 0.670 1.730 3.860 1.760 ;
        RECT 6.310 1.730 6.610 1.760 ;
        RECT -3.330 1.430 9.530 1.730 ;
        RECT -3.330 1.090 -2.670 1.430 ;
        RECT 0.670 1.060 0.970 1.430 ;
        RECT 3.560 1.090 3.860 1.430 ;
        RECT 6.310 1.090 6.610 1.430 ;
        RECT 3.560 1.060 6.610 1.090 ;
        RECT 9.230 1.060 9.530 1.430 ;
        RECT -2.240 0.520 -1.580 0.880 ;
        RECT 0.670 0.760 9.530 1.060 ;
        RECT 11.990 1.100 12.290 3.620 ;
        RECT 14.820 3.590 17.930 3.620 ;
        RECT 14.820 1.100 15.120 3.590 ;
        RECT 17.630 1.100 17.930 3.590 ;
        RECT 20.580 1.100 20.880 3.620 ;
        RECT 11.990 0.800 20.940 1.100 ;
        RECT 17.630 0.790 20.940 0.800 ;
        RECT -2.240 0.220 -1.190 0.520 ;
        RECT -1.490 -0.020 -1.190 0.220 ;
        RECT 20.640 -0.020 20.940 0.790 ;
        RECT -1.490 -0.320 20.940 -0.020 ;
  END
END sky130_hilas_capacitorArray01

MACRO sky130_hilas_TA2Cell_1FG
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TA2Cell_1FG ;
  ORIGIN 26.160 -1.350 ;
  SIZE 28.090 BY 6.150 ;
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -16.850 2.660 -16.540 2.720 ;
        RECT -17.310 2.650 -16.540 2.660 ;
        RECT -17.310 2.640 -16.420 2.650 ;
        RECT -17.310 2.430 -14.630 2.640 ;
        RECT -17.310 2.410 -16.420 2.430 ;
        RECT -16.850 2.390 -16.540 2.410 ;
    END
  END VIN12
  PIN VIN11
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -16.880 6.370 -16.570 6.410 ;
        RECT -17.260 6.350 -16.420 6.370 ;
        RECT -17.260 6.170 -14.630 6.350 ;
        RECT -16.880 6.080 -16.570 6.170 ;
    END
  END VIN11
  PIN VIN21
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -2.200 4.750 -1.890 4.790 ;
        RECT -2.520 4.740 -1.860 4.750 ;
        RECT -2.520 4.510 -1.420 4.740 ;
        RECT -2.200 4.460 -1.890 4.510 ;
    END
  END VIN21
  PIN VIN22
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -1.960 7.430 -1.650 7.440 ;
        RECT -2.530 7.420 -1.650 7.430 ;
        RECT -2.600 7.180 -1.650 7.420 ;
        RECT -1.960 7.110 -1.650 7.180 ;
    END
  END VIN22
  PIN VPWR
    USE ANALOG ;
    ANTENNADIFFAREA 1.373600 ;
    PORT
      LAYER nwell ;
        RECT 0.650 1.400 1.930 7.450 ;
      LAYER met1 ;
        RECT 0.630 7.300 0.910 7.450 ;
        RECT 0.640 5.870 0.910 7.300 ;
        RECT 0.640 5.580 0.920 5.870 ;
        RECT 0.640 3.280 0.910 5.580 ;
        RECT 0.640 2.990 0.920 3.280 ;
        RECT 0.640 1.400 0.910 2.990 ;
    END
  END VPWR
  PIN VGND
    USE ANALOG ;
    ANTENNADIFFAREA 5.718600 ;
    PORT
      LAYER met2 ;
        RECT -17.680 4.290 -17.360 4.340 ;
        RECT -17.680 4.040 -11.660 4.290 ;
        RECT -11.980 3.970 -11.660 4.040 ;
        RECT -11.980 1.750 -11.660 1.760 ;
        RECT -1.540 1.750 -1.210 1.890 ;
        RECT -11.980 1.590 -1.210 1.750 ;
        RECT -11.980 1.580 -11.290 1.590 ;
        RECT -11.980 1.460 -11.660 1.580 ;
    END
    PORT
      LAYER met1 ;
        RECT -1.540 1.600 -1.210 1.890 ;
        RECT -0.030 1.600 0.310 7.450 ;
        RECT -1.550 1.570 -1.130 1.600 ;
        RECT -0.530 1.570 0.310 1.600 ;
        RECT -1.550 1.460 0.310 1.570 ;
        RECT -1.270 1.430 -0.370 1.460 ;
        RECT -0.030 1.400 0.310 1.460 ;
      LAYER via ;
        RECT -1.510 1.610 -1.240 1.870 ;
    END
    PORT
      LAYER met1 ;
        RECT -17.690 6.480 -17.460 7.450 ;
        RECT -17.700 6.230 -17.460 6.480 ;
        RECT -17.690 4.340 -17.460 6.230 ;
        RECT -17.690 4.040 -17.360 4.340 ;
        RECT -17.690 3.870 -17.440 4.040 ;
        RECT -17.690 1.400 -17.460 3.870 ;
      LAYER via ;
        RECT -17.650 4.060 -17.390 4.320 ;
    END
    PORT
      LAYER met1 ;
        RECT -11.900 4.290 -11.670 7.450 ;
        RECT -11.980 3.970 -11.660 4.290 ;
        RECT -11.900 1.760 -11.670 3.970 ;
        RECT -11.980 1.460 -11.660 1.760 ;
        RECT -11.900 1.400 -11.670 1.460 ;
      LAYER via ;
        RECT -11.950 4.000 -11.690 4.260 ;
        RECT -11.950 1.480 -11.690 1.740 ;
    END
  END VGND
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -26.160 1.350 -22.850 7.500 ;
        RECT -6.510 7.450 -3.200 7.500 ;
        RECT -6.510 7.440 -1.730 7.450 ;
        RECT -6.510 1.400 -1.350 7.440 ;
        RECT -6.510 1.350 -3.200 1.400 ;
      LAYER met2 ;
        RECT -25.920 7.280 -25.600 7.400 ;
        RECT -3.720 7.280 -3.400 7.400 ;
        RECT -25.920 7.100 -3.400 7.280 ;
        RECT -4.590 4.590 -4.270 4.850 ;
        RECT -4.550 4.570 -3.370 4.590 ;
        RECT -4.550 4.310 -3.330 4.570 ;
        RECT -4.550 4.250 -3.370 4.310 ;
        RECT -4.590 4.240 -3.370 4.250 ;
        RECT -4.590 3.990 -4.270 4.240 ;
    END
    PORT
      LAYER met1 ;
        RECT -3.720 7.400 -3.440 7.450 ;
        RECT -3.720 7.100 -3.400 7.400 ;
        RECT -3.720 6.800 -3.440 7.100 ;
        RECT -3.830 6.200 -3.440 6.800 ;
        RECT -3.720 4.600 -3.440 6.200 ;
        RECT -3.720 4.280 -3.360 4.600 ;
        RECT -3.720 2.650 -3.440 4.280 ;
        RECT -3.830 2.050 -3.440 2.650 ;
        RECT -3.720 1.400 -3.440 2.050 ;
      LAYER via ;
        RECT -3.690 7.120 -3.430 7.380 ;
        RECT -3.620 4.310 -3.360 4.570 ;
    END
    PORT
      LAYER met1 ;
        RECT -25.920 7.400 -25.640 7.450 ;
        RECT -25.920 7.120 -25.600 7.400 ;
        RECT -25.920 6.800 -25.640 7.120 ;
        RECT -25.920 6.200 -25.530 6.800 ;
        RECT -25.920 2.650 -25.640 6.200 ;
        RECT -25.920 2.050 -25.530 2.650 ;
        RECT -25.920 1.400 -25.640 2.050 ;
      LAYER via ;
        RECT -25.890 7.130 -25.630 7.390 ;
    END
  END VINJ
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.308800 ;
    PORT
      LAYER met2 ;
        RECT -0.990 4.970 -0.680 5.030 ;
        RECT 1.310 4.970 1.620 4.990 ;
        RECT -0.990 4.740 1.930 4.970 ;
        RECT -0.990 4.700 -0.680 4.740 ;
        RECT 1.310 4.660 1.620 4.740 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.308800 ;
    PORT
      LAYER met2 ;
        RECT -0.990 4.140 -0.680 4.190 ;
        RECT 1.300 4.140 1.610 4.270 ;
        RECT -0.990 3.920 1.930 4.140 ;
        RECT -0.990 3.860 -0.680 3.920 ;
    END
  END OUTPUT2
  PIN DRAIN1
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER met2 ;
        RECT -23.990 6.950 -23.680 6.960 ;
        RECT -5.680 6.950 -5.370 6.960 ;
        RECT -26.160 6.770 -3.200 6.950 ;
        RECT -23.990 6.630 -23.680 6.770 ;
        RECT -5.680 6.630 -5.370 6.770 ;
    END
  END DRAIN1
  PIN DRAIN2
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER met2 ;
        RECT -23.990 2.080 -23.680 2.220 ;
        RECT -26.160 2.070 -23.680 2.080 ;
        RECT -5.680 2.080 -5.370 2.220 ;
        RECT -5.680 2.070 -3.200 2.080 ;
        RECT -26.160 1.920 -3.200 2.070 ;
        RECT -26.160 1.900 -23.680 1.920 ;
        RECT -23.990 1.890 -23.680 1.900 ;
        RECT -5.680 1.900 -3.200 1.920 ;
        RECT -5.680 1.890 -5.370 1.900 ;
    END
  END DRAIN2
  PIN COLSEL2
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT -25.390 5.990 -25.200 7.450 ;
        RECT -25.420 5.960 -25.200 5.990 ;
        RECT -25.430 5.690 -25.180 5.960 ;
        RECT -25.430 5.680 -25.190 5.690 ;
        RECT -25.420 5.440 -25.190 5.680 ;
        RECT -25.390 3.410 -25.230 5.440 ;
        RECT -25.420 3.170 -25.190 3.410 ;
        RECT -25.430 3.160 -25.190 3.170 ;
        RECT -25.430 2.890 -25.180 3.160 ;
        RECT -25.420 2.860 -25.200 2.890 ;
        RECT -25.390 1.400 -25.200 2.860 ;
    END
  END COLSEL2
  PIN GATE2
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT -21.120 5.060 -18.400 6.710 ;
        RECT -21.110 5.020 -18.400 5.060 ;
        RECT -21.110 3.690 -18.400 3.730 ;
        RECT -21.120 2.040 -18.400 3.690 ;
      LAYER met1 ;
        RECT -18.910 6.240 -18.680 7.450 ;
        RECT -18.940 5.450 -18.680 6.240 ;
        RECT -18.910 3.300 -18.680 5.450 ;
        RECT -18.940 2.510 -18.680 3.300 ;
        RECT -18.910 1.400 -18.680 2.510 ;
    END
  END GATE2
  PIN GATE1
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT -10.960 5.060 -8.240 6.710 ;
        RECT -10.960 5.020 -8.250 5.060 ;
        RECT -10.960 3.690 -8.250 3.730 ;
        RECT -10.960 2.040 -8.240 3.690 ;
      LAYER met1 ;
        RECT -10.680 6.240 -10.450 7.450 ;
        RECT -10.680 5.450 -10.420 6.240 ;
        RECT -10.680 3.300 -10.450 5.450 ;
        RECT -10.680 2.510 -10.420 3.300 ;
        RECT -10.680 1.400 -10.450 2.510 ;
    END
  END GATE1
  PIN COLSEL1
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT -4.160 5.990 -3.970 7.450 ;
        RECT -4.160 5.960 -3.940 5.990 ;
        RECT -4.180 5.690 -3.930 5.960 ;
        RECT -4.170 5.680 -3.930 5.690 ;
        RECT -4.170 5.440 -3.940 5.680 ;
        RECT -4.130 3.410 -3.970 5.440 ;
        RECT -4.170 3.170 -3.940 3.410 ;
        RECT -4.170 3.160 -3.930 3.170 ;
        RECT -4.180 2.890 -3.930 3.160 ;
        RECT -4.160 2.860 -3.940 2.890 ;
        RECT -4.160 1.400 -3.970 2.860 ;
    END
  END COLSEL1
  PIN VTUN
    ANTENNADIFFAREA 5.032200 ;
    PORT
      LAYER nwell ;
        RECT -16.370 6.700 -12.990 7.450 ;
        RECT -16.380 3.130 -12.980 6.700 ;
        RECT -16.370 1.410 -12.990 3.130 ;
      LAYER met1 ;
        RECT -15.400 7.290 -13.960 7.450 ;
        RECT -15.400 1.410 -14.980 7.290 ;
        RECT -14.380 1.400 -13.960 7.290 ;
    END
  END VTUN
  OBS
      LAYER li1 ;
        RECT -2.220 7.400 -2.050 7.450 ;
        RECT -25.760 6.770 -25.560 7.120 ;
        RECT -24.280 6.870 -23.750 7.040 ;
        RECT -25.770 6.740 -25.560 6.770 ;
        RECT -25.770 6.160 -25.550 6.740 ;
        RECT -25.770 6.150 -25.560 6.160 ;
        RECT -25.390 5.980 -25.200 5.990 ;
        RECT -25.400 5.690 -25.200 5.980 ;
        RECT -25.480 5.360 -25.190 5.690 ;
        RECT -25.000 4.880 -24.830 6.490 ;
        RECT -25.010 4.690 -24.830 4.880 ;
        RECT -24.170 5.960 -24.000 6.480 ;
        RECT -21.560 6.440 -16.500 7.270 ;
        RECT -2.220 7.140 -1.660 7.400 ;
        RECT -0.750 7.150 -0.550 7.190 ;
        RECT -2.220 7.120 -2.050 7.140 ;
        RECT -5.610 6.870 -5.080 7.040 ;
        RECT -3.800 6.770 -3.600 7.120 ;
        RECT -3.800 6.740 -3.590 6.770 ;
        RECT -17.050 6.360 -16.570 6.440 ;
        RECT -24.170 5.700 -23.840 5.960 ;
        RECT -24.170 4.790 -24.000 5.700 ;
        RECT -18.930 5.500 -18.700 6.190 ;
        RECT -17.050 6.110 -16.580 6.360 ;
        RECT -15.620 5.310 -15.070 5.740 ;
        RECT -14.290 5.310 -13.740 5.740 ;
        RECT -10.660 5.500 -10.430 6.190 ;
        RECT -5.360 5.960 -5.190 6.480 ;
        RECT -5.520 5.700 -5.190 5.960 ;
        RECT -17.860 4.470 -17.470 4.880 ;
        RECT -21.220 4.290 -17.470 4.470 ;
        RECT -25.010 3.970 -24.830 4.160 ;
        RECT -25.480 3.160 -25.190 3.490 ;
        RECT -25.400 2.870 -25.200 3.160 ;
        RECT -25.390 2.860 -25.200 2.870 ;
        RECT -25.770 2.690 -25.560 2.700 ;
        RECT -25.770 2.110 -25.550 2.690 ;
        RECT -25.000 2.360 -24.830 3.970 ;
        RECT -24.170 3.200 -24.000 4.060 ;
        RECT -17.860 3.870 -17.470 4.290 ;
        RECT -11.920 4.470 -11.500 4.880 ;
        RECT -5.360 4.790 -5.190 5.700 ;
        RECT -4.530 4.880 -4.360 6.490 ;
        RECT -3.810 6.160 -3.590 6.740 ;
        RECT -3.800 6.150 -3.590 6.160 ;
        RECT -2.800 6.040 -2.620 6.970 ;
        RECT -0.980 6.890 -0.550 7.150 ;
        RECT -2.070 6.710 -1.740 6.880 ;
        RECT -0.750 6.860 -0.550 6.890 ;
        RECT -1.990 6.570 -1.740 6.710 ;
        RECT -1.990 6.310 -1.510 6.570 ;
        RECT -1.160 6.500 -0.990 6.540 ;
        RECT -0.750 6.500 -0.550 6.530 ;
        RECT -2.920 6.010 -2.600 6.040 ;
        RECT -4.160 5.980 -3.970 5.990 ;
        RECT -4.160 5.690 -3.960 5.980 ;
        RECT -2.920 5.820 -2.590 6.010 ;
        RECT -2.920 5.780 -2.600 5.820 ;
        RECT -4.170 5.360 -3.880 5.690 ;
        RECT -4.530 4.690 -4.350 4.880 ;
        RECT -11.920 4.290 -8.140 4.470 ;
        RECT -15.620 3.580 -15.070 4.010 ;
        RECT -14.290 3.580 -13.740 4.010 ;
        RECT -11.920 3.870 -11.500 4.290 ;
        RECT -24.170 2.940 -23.840 3.200 ;
        RECT -24.170 2.370 -24.000 2.940 ;
        RECT -18.930 2.560 -18.700 3.290 ;
        RECT -16.890 2.430 -16.550 2.680 ;
        RECT -10.660 2.560 -10.430 3.290 ;
        RECT -5.360 3.200 -5.190 4.060 ;
        RECT -5.520 2.940 -5.190 3.200 ;
        RECT -16.890 2.350 -16.540 2.430 ;
        RECT -5.360 2.370 -5.190 2.940 ;
        RECT -4.530 3.970 -4.350 4.160 ;
        RECT -4.530 2.360 -4.360 3.970 ;
        RECT -4.170 3.160 -3.880 3.490 ;
        RECT -4.160 2.870 -3.960 3.160 ;
        RECT -4.160 2.860 -3.970 2.870 ;
        RECT -3.800 2.690 -3.590 2.700 ;
        RECT -25.770 2.080 -25.560 2.110 ;
        RECT -25.760 1.730 -25.560 2.080 ;
        RECT -24.280 1.810 -23.750 1.980 ;
        RECT -21.590 1.500 -16.540 2.350 ;
        RECT -3.810 2.110 -3.590 2.690 ;
        RECT -3.800 2.080 -3.590 2.110 ;
        RECT -5.610 1.810 -5.080 1.980 ;
        RECT -3.800 1.730 -3.600 2.080 ;
        RECT -2.800 1.870 -2.620 5.780 ;
        RECT -1.990 4.930 -1.820 6.310 ;
        RECT -1.160 6.240 -0.550 6.500 ;
        RECT -1.160 6.210 -0.990 6.240 ;
        RECT -0.750 6.200 -0.550 6.240 ;
        RECT -0.160 6.200 0.390 7.190 ;
        RECT 1.210 7.040 1.840 7.210 ;
        RECT 1.210 6.940 1.600 7.040 ;
        RECT 1.210 6.910 1.590 6.940 ;
        RECT 1.210 6.760 1.570 6.910 ;
        RECT 0.860 6.590 1.570 6.760 ;
        RECT 0.860 5.840 1.560 6.150 ;
        RECT -1.160 5.650 -0.990 5.680 ;
        RECT -0.750 5.650 -0.550 5.690 ;
        RECT -1.160 5.390 -0.550 5.650 ;
        RECT -1.160 5.350 -0.990 5.390 ;
        RECT -0.750 5.360 -0.550 5.390 ;
        RECT -0.750 5.000 -0.550 5.030 ;
        RECT -2.190 4.730 -1.870 4.760 ;
        RECT -0.980 4.740 -0.550 5.000 ;
        RECT -2.190 4.540 -1.860 4.730 ;
        RECT -0.750 4.700 -0.550 4.740 ;
        RECT -0.160 4.700 0.390 5.690 ;
        RECT 0.710 5.610 1.560 5.840 ;
        RECT 0.860 5.270 1.560 5.610 ;
        RECT 1.320 4.910 1.640 4.950 ;
        RECT 1.320 4.850 1.650 4.910 ;
        RECT 0.850 4.720 1.650 4.850 ;
        RECT 0.850 4.690 1.640 4.720 ;
        RECT 0.850 4.670 1.550 4.690 ;
        RECT -2.190 4.500 -1.870 4.540 ;
        RECT -2.190 4.420 -2.020 4.500 ;
        RECT -2.240 4.250 -2.020 4.420 ;
        RECT -2.240 4.090 -2.070 4.250 ;
        RECT 1.310 4.190 1.630 4.230 ;
        RECT -0.750 4.150 -0.550 4.190 ;
        RECT -1.710 3.830 -1.520 3.950 ;
        RECT -0.980 3.890 -0.550 4.150 ;
        RECT -0.750 3.860 -0.550 3.890 ;
        RECT -2.070 3.720 -1.520 3.830 ;
        RECT -2.070 3.660 -1.530 3.720 ;
        RECT -1.990 1.880 -1.820 3.660 ;
        RECT -1.160 3.500 -0.990 3.540 ;
        RECT -0.750 3.500 -0.550 3.530 ;
        RECT -1.160 3.240 -0.550 3.500 ;
        RECT -1.160 3.210 -0.990 3.240 ;
        RECT -0.750 3.200 -0.550 3.240 ;
        RECT -0.160 3.200 0.390 4.190 ;
        RECT 0.850 4.010 1.640 4.190 ;
        RECT 1.310 4.000 1.640 4.010 ;
        RECT 1.310 3.970 1.630 4.000 ;
        RECT 0.860 3.250 1.560 3.590 ;
        RECT 0.710 3.020 1.560 3.250 ;
        RECT 0.860 2.710 1.560 3.020 ;
        RECT -1.160 2.650 -0.990 2.680 ;
        RECT -0.750 2.650 -0.550 2.690 ;
        RECT -1.160 2.390 -0.550 2.650 ;
        RECT -1.160 2.350 -0.990 2.390 ;
        RECT -0.750 2.360 -0.550 2.390 ;
        RECT -0.750 2.000 -0.550 2.030 ;
        RECT -0.980 1.740 -0.550 2.000 ;
        RECT -0.750 1.700 -0.550 1.740 ;
        RECT -0.160 1.700 0.390 2.690 ;
        RECT 0.860 2.100 1.570 2.270 ;
        RECT 1.210 1.820 1.570 2.100 ;
        RECT 1.210 1.650 1.840 1.820 ;
      LAYER mcon ;
        RECT -23.930 6.870 -23.750 7.040 ;
        RECT -25.740 6.570 -25.570 6.740 ;
        RECT -25.390 5.730 -25.210 5.920 ;
        RECT -1.890 7.180 -1.720 7.350 ;
        RECT -3.790 6.570 -3.620 6.740 ;
        RECT -18.900 5.990 -18.730 6.160 ;
        RECT -16.810 6.150 -16.640 6.320 ;
        RECT -24.070 5.740 -23.900 5.910 ;
        RECT -10.630 5.990 -10.460 6.160 ;
        RECT -18.900 5.540 -18.730 5.710 ;
        RECT -15.340 5.390 -15.070 5.660 ;
        RECT -14.290 5.390 -14.020 5.660 ;
        RECT -10.630 5.540 -10.460 5.710 ;
        RECT -5.460 5.740 -5.290 5.910 ;
        RECT -17.660 4.640 -17.490 4.810 ;
        RECT -17.660 4.280 -17.490 4.450 ;
        RECT -25.390 2.930 -25.210 3.120 ;
        RECT -17.650 3.920 -17.480 4.090 ;
        RECT -11.870 4.640 -11.700 4.810 ;
        RECT -0.920 6.930 -0.750 7.100 ;
        RECT 0.060 6.610 0.230 6.780 ;
        RECT 1.330 6.950 1.500 7.120 ;
        RECT -1.740 6.350 -1.570 6.520 ;
        RECT -4.150 5.730 -3.970 5.920 ;
        RECT -2.860 5.830 -2.690 6.000 ;
        RECT -11.870 4.280 -11.700 4.450 ;
        RECT -15.340 3.660 -15.070 3.930 ;
        RECT -14.290 3.660 -14.020 3.930 ;
        RECT -11.870 3.920 -11.700 4.090 ;
        RECT -24.070 2.980 -23.900 3.150 ;
        RECT -18.900 3.040 -18.730 3.210 ;
        RECT -18.900 2.590 -18.730 2.760 ;
        RECT -10.630 3.040 -10.460 3.210 ;
        RECT -5.460 2.980 -5.290 3.150 ;
        RECT -16.780 2.460 -16.610 2.630 ;
        RECT -10.630 2.590 -10.460 2.760 ;
        RECT -4.150 2.930 -3.970 3.120 ;
        RECT -25.740 2.110 -25.570 2.280 ;
        RECT -23.930 1.810 -23.750 1.980 ;
        RECT -3.790 2.110 -3.620 2.280 ;
        RECT -0.970 6.280 -0.800 6.450 ;
        RECT -0.970 5.440 -0.800 5.610 ;
        RECT 0.720 5.640 0.890 5.810 ;
        RECT 0.060 5.110 0.230 5.280 ;
        RECT -0.920 4.790 -0.750 4.960 ;
        RECT -2.130 4.550 -1.960 4.720 ;
        RECT 1.380 4.730 1.550 4.900 ;
        RECT -1.700 3.750 -1.530 3.920 ;
        RECT -0.920 3.930 -0.750 4.100 ;
        RECT 1.370 4.010 1.540 4.180 ;
        RECT 0.060 3.610 0.230 3.780 ;
        RECT -0.970 3.280 -0.800 3.450 ;
        RECT 0.720 3.050 0.890 3.220 ;
        RECT -0.970 2.440 -0.800 2.610 ;
        RECT 0.060 2.110 0.230 2.280 ;
        RECT -0.920 1.790 -0.750 1.960 ;
        RECT 1.290 1.760 1.460 1.930 ;
      LAYER met1 ;
        RECT -1.970 7.110 -1.650 7.430 ;
        RECT -23.990 6.630 -23.680 7.070 ;
        RECT -5.680 6.630 -5.370 7.070 ;
        RECT -0.990 6.860 -0.670 7.180 ;
        RECT 1.260 6.880 1.580 7.200 ;
        RECT -16.890 6.080 -16.570 6.400 ;
        RECT -1.820 6.280 -1.500 6.600 ;
        RECT -1.040 6.210 -0.720 6.530 ;
        RECT -24.150 5.670 -23.830 5.990 ;
        RECT -5.530 5.670 -5.210 5.990 ;
        RECT -2.930 5.750 -2.610 6.070 ;
        RECT -1.710 5.590 -1.500 5.700 ;
        RECT -1.730 5.270 -1.470 5.590 ;
        RECT -1.040 5.360 -0.720 5.680 ;
        RECT -25.040 4.880 -24.800 5.010 ;
        RECT -25.060 4.560 -24.800 4.880 ;
        RECT -4.560 4.880 -4.320 5.010 ;
        RECT -4.560 4.560 -4.300 4.880 ;
        RECT -2.200 4.470 -1.880 4.790 ;
        RECT -25.060 3.960 -24.800 4.280 ;
        RECT -25.040 3.840 -24.800 3.960 ;
        RECT -4.560 3.960 -4.300 4.280 ;
        RECT -1.710 3.980 -1.500 5.270 ;
        RECT -0.990 4.710 -0.670 5.030 ;
        RECT 1.310 4.660 1.630 4.980 ;
        RECT -4.560 3.840 -4.320 3.960 ;
        RECT -1.730 3.690 -1.500 3.980 ;
        RECT -0.990 3.860 -0.670 4.180 ;
        RECT 1.300 3.940 1.620 4.260 ;
        RECT -24.150 2.910 -23.830 3.230 ;
        RECT -5.530 2.910 -5.210 3.230 ;
        RECT -1.040 3.210 -0.720 3.530 ;
        RECT -16.860 2.390 -16.540 2.710 ;
        RECT -1.040 2.360 -0.720 2.680 ;
        RECT -23.990 1.780 -23.680 2.220 ;
        RECT -5.680 1.780 -5.370 2.220 ;
        RECT -0.990 1.710 -0.670 2.030 ;
        RECT 1.220 1.690 1.540 2.010 ;
      LAYER via ;
        RECT -1.940 7.140 -1.680 7.400 ;
        RECT -23.970 6.660 -23.710 6.920 ;
        RECT -5.650 6.660 -5.390 6.920 ;
        RECT -0.960 6.890 -0.700 7.150 ;
        RECT 1.290 6.910 1.550 7.170 ;
        RECT -16.860 6.110 -16.600 6.370 ;
        RECT -1.790 6.310 -1.530 6.570 ;
        RECT -1.010 6.240 -0.750 6.500 ;
        RECT -24.120 5.700 -23.860 5.960 ;
        RECT -5.500 5.700 -5.240 5.960 ;
        RECT -2.900 5.780 -2.640 6.040 ;
        RECT -1.730 5.300 -1.470 5.560 ;
        RECT -1.010 5.390 -0.750 5.650 ;
        RECT -25.060 4.590 -24.800 4.850 ;
        RECT -4.560 4.590 -4.300 4.850 ;
        RECT -2.170 4.500 -1.910 4.760 ;
        RECT -25.060 3.990 -24.800 4.250 ;
        RECT -4.560 3.990 -4.300 4.250 ;
        RECT -0.960 4.740 -0.700 5.000 ;
        RECT 1.340 4.690 1.600 4.950 ;
        RECT -0.960 3.890 -0.700 4.150 ;
        RECT 1.330 3.970 1.590 4.230 ;
        RECT -1.010 3.240 -0.750 3.500 ;
        RECT -24.120 2.940 -23.860 3.200 ;
        RECT -5.500 2.940 -5.240 3.200 ;
        RECT -16.830 2.420 -16.570 2.680 ;
        RECT -1.010 2.390 -0.750 2.650 ;
        RECT -23.970 1.930 -23.710 2.190 ;
        RECT -5.650 1.930 -5.390 2.190 ;
        RECT -0.960 1.740 -0.700 2.000 ;
        RECT 1.250 1.720 1.510 1.980 ;
      LAYER met2 ;
        RECT -0.990 7.110 -0.680 7.190 ;
        RECT 1.260 7.110 1.570 7.210 ;
        RECT -0.990 6.880 1.570 7.110 ;
        RECT -0.990 6.860 -0.680 6.880 ;
        RECT -1.810 6.570 -1.500 6.610 ;
        RECT -1.990 6.460 -1.270 6.570 ;
        RECT -1.040 6.460 -0.730 6.540 ;
        RECT -1.990 6.320 -0.730 6.460 ;
        RECT -1.810 6.280 -0.730 6.320 ;
        RECT -1.540 6.250 -0.730 6.280 ;
        RECT -1.540 6.210 -1.270 6.250 ;
        RECT -1.040 6.210 -0.730 6.250 ;
        RECT -24.140 5.930 -23.830 6.000 ;
        RECT -26.160 5.920 -23.830 5.930 ;
        RECT -5.530 5.930 -5.220 6.000 ;
        RECT -2.930 5.930 -2.620 6.070 ;
        RECT -26.160 5.710 -6.670 5.920 ;
        RECT -24.850 5.700 -6.670 5.710 ;
        RECT -24.140 5.670 -23.830 5.700 ;
        RECT -25.090 4.730 -7.850 4.950 ;
        RECT -25.090 4.590 -24.770 4.730 ;
        RECT -25.070 4.250 -24.810 4.590 ;
        RECT -25.090 3.990 -24.770 4.250 ;
        RECT -24.140 3.170 -23.830 3.240 ;
        RECT -26.160 2.960 -11.150 3.170 ;
        RECT -24.850 2.950 -11.150 2.960 ;
        RECT -24.140 2.910 -23.830 2.950 ;
        RECT -11.370 2.620 -11.150 2.950 ;
        RECT -8.070 3.120 -7.850 4.730 ;
        RECT -6.890 4.500 -6.670 5.700 ;
        RECT -5.530 5.740 -2.620 5.930 ;
        RECT -5.530 5.710 -2.930 5.740 ;
        RECT -5.530 5.670 -5.220 5.710 ;
        RECT -1.470 5.640 -1.270 5.650 ;
        RECT -1.040 5.640 -0.730 5.680 ;
        RECT -1.470 5.560 -0.730 5.640 ;
        RECT -1.760 5.540 -0.730 5.560 ;
        RECT -1.810 5.430 -0.730 5.540 ;
        RECT -1.810 5.300 -1.250 5.430 ;
        RECT -1.040 5.350 -0.730 5.430 ;
        RECT -1.810 5.290 -1.340 5.300 ;
        RECT -6.920 4.460 -6.670 4.500 ;
        RECT -6.920 3.820 -6.660 4.460 ;
        RECT -6.920 3.610 -2.790 3.820 ;
        RECT -3.000 3.470 -2.790 3.610 ;
        RECT -1.040 3.470 -0.730 3.540 ;
        RECT -3.000 3.260 -0.730 3.470 ;
        RECT -1.340 3.250 -0.730 3.260 ;
        RECT -5.530 3.170 -5.220 3.240 ;
        RECT -1.040 3.210 -0.730 3.250 ;
        RECT -5.530 3.120 -3.200 3.170 ;
        RECT -8.070 2.960 -3.200 3.120 ;
        RECT -8.070 2.900 -5.220 2.960 ;
        RECT -1.040 2.670 -0.730 2.680 ;
        RECT -7.000 2.620 -0.730 2.670 ;
        RECT -11.370 2.460 -0.730 2.620 ;
        RECT -11.370 2.400 -6.610 2.460 ;
        RECT -1.340 2.430 -0.730 2.460 ;
        RECT -1.040 2.350 -0.730 2.430 ;
        RECT -0.990 1.980 -0.680 2.030 ;
        RECT 1.220 1.980 1.530 2.020 ;
        RECT -0.990 1.750 1.720 1.980 ;
        RECT -0.990 1.700 -0.680 1.750 ;
        RECT 1.220 1.690 1.530 1.750 ;
  END
END sky130_hilas_TA2Cell_1FG

MACRO sky130_hilas_FGBiasWeakGate2x1cell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_FGBiasWeakGate2x1cell ;
  ORIGIN 3.960 3.870 ;
  SIZE 11.530 BY 6.150 ;
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 5.090 1.730 5.400 1.740 ;
        RECT -3.960 1.550 7.570 1.730 ;
        RECT 5.090 1.410 5.400 1.550 ;
    END
  END DRAIN1
  PIN VIN11
    PORT
      LAYER met2 ;
        RECT -2.020 1.140 -1.710 1.190 ;
        RECT -2.170 1.130 -1.710 1.140 ;
        RECT -3.960 0.950 -1.710 1.130 ;
        RECT -2.020 0.860 -1.710 0.950 ;
    END
  END VIN11
  PIN ROW1
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 5.240 0.710 5.550 0.780 ;
        RECT 5.240 0.700 7.570 0.710 ;
        RECT -3.960 0.490 7.570 0.700 ;
        RECT -3.960 0.480 6.260 0.490 ;
        RECT 5.240 0.450 5.550 0.480 ;
    END
  END ROW1
  PIN ROW2
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 5.240 -2.050 5.550 -1.980 ;
        RECT -3.960 -2.260 7.570 -2.050 ;
        RECT -3.960 -2.270 6.260 -2.260 ;
        RECT 5.240 -2.310 5.550 -2.270 ;
    END
  END ROW2
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 4.260 -3.870 7.570 2.280 ;
      LAYER met1 ;
        RECT 7.050 1.580 7.330 2.230 ;
        RECT 6.940 0.980 7.330 1.580 ;
        RECT 7.050 -2.570 7.330 0.980 ;
        RECT 6.940 -3.170 7.330 -2.570 ;
        RECT 7.050 -3.820 7.330 -3.170 ;
    END
  END VINJ
  PIN COLSEL1
    USE ANALOG ;
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT 6.610 0.770 6.800 2.230 ;
        RECT 6.610 0.740 6.830 0.770 ;
        RECT 6.590 0.470 6.840 0.740 ;
        RECT 6.600 0.460 6.840 0.470 ;
        RECT 6.600 0.220 6.830 0.460 ;
        RECT 6.640 -1.810 6.800 0.220 ;
        RECT 6.600 -2.050 6.830 -1.810 ;
        RECT 6.600 -2.060 6.840 -2.050 ;
        RECT 6.590 -2.330 6.840 -2.060 ;
        RECT 6.610 -2.360 6.830 -2.330 ;
        RECT 6.610 -3.820 6.800 -2.360 ;
    END
  END COLSEL1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT -1.130 1.260 -0.900 2.230 ;
        RECT -1.130 1.010 -0.890 1.260 ;
        RECT -1.130 -3.820 -0.900 1.010 ;
    END
  END VGND
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT -0.190 -0.160 2.530 1.490 ;
        RECT -0.190 -0.200 2.520 -0.160 ;
        RECT -0.190 -1.530 2.520 -1.490 ;
        RECT -0.190 -3.180 2.530 -1.530 ;
      LAYER met1 ;
        RECT 0.090 1.020 0.320 2.230 ;
        RECT 0.090 0.230 0.350 1.020 ;
        RECT 0.090 -1.920 0.320 0.230 ;
        RECT 0.090 -2.710 0.350 -1.920 ;
        RECT 0.090 -3.820 0.320 -2.710 ;
    END
  END GATE1
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 2.516100 ;
    PORT
      LAYER nwell ;
        RECT -3.950 1.480 -2.220 2.230 ;
        RECT -3.950 0.330 -2.210 1.480 ;
        RECT -3.940 -1.910 -2.210 0.330 ;
        RECT -3.950 -2.090 -2.210 -1.910 ;
        RECT -3.950 -3.810 -2.220 -2.090 ;
      LAYER met1 ;
        RECT -3.610 -3.810 -3.190 2.230 ;
    END
  END VTUN
  PIN DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 5.090 -3.140 5.400 -3.000 ;
        RECT 5.090 -3.150 7.570 -3.140 ;
        RECT -3.960 -3.300 7.570 -3.150 ;
        RECT 5.090 -3.320 7.570 -3.300 ;
        RECT 5.090 -3.330 5.400 -3.320 ;
    END
  END DRAIN2
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -2.050 -2.580 -1.740 -2.500 ;
        RECT -3.960 -2.790 -1.740 -2.580 ;
        RECT -2.050 -2.830 -1.740 -2.790 ;
    END
  END VIN12
  PIN COMMONSOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 1.030400 ;
    PORT
      LAYER met2 ;
        RECT -3.960 -0.490 6.500 -0.270 ;
        RECT 6.180 -0.630 6.500 -0.490 ;
        RECT 6.220 -0.970 6.480 -0.630 ;
        RECT 6.180 -1.230 6.500 -0.970 ;
    END
  END COMMONSOURCE
  OBS
      LAYER li1 ;
        RECT -2.090 1.220 2.970 2.050 ;
        RECT 5.160 1.650 5.690 1.820 ;
        RECT 6.970 1.550 7.170 1.900 ;
        RECT 6.970 1.520 7.180 1.550 ;
        RECT -2.020 1.140 -1.540 1.220 ;
        RECT -2.010 0.890 -1.540 1.140 ;
        RECT -3.520 0.090 -2.970 0.520 ;
        RECT 0.110 0.280 0.340 0.970 ;
        RECT 5.410 0.740 5.580 1.260 ;
        RECT 5.250 0.480 5.580 0.740 ;
        RECT -0.920 -0.740 -0.730 -0.340 ;
        RECT 5.410 -0.430 5.580 0.480 ;
        RECT 6.240 -0.340 6.410 1.270 ;
        RECT 6.960 0.940 7.180 1.520 ;
        RECT 6.970 0.930 7.180 0.940 ;
        RECT 6.610 0.760 6.800 0.770 ;
        RECT 6.610 0.470 6.810 0.760 ;
        RECT 6.600 0.140 6.890 0.470 ;
        RECT 6.240 -0.530 6.420 -0.340 ;
        RECT -1.110 -0.750 -0.730 -0.740 ;
        RECT -1.110 -0.930 2.630 -0.750 ;
        RECT -1.110 -0.970 -0.730 -0.930 ;
        RECT -3.520 -1.640 -2.970 -1.210 ;
        RECT -0.920 -1.350 -0.730 -0.970 ;
        RECT -2.040 -2.790 -1.700 -2.540 ;
        RECT 0.110 -2.660 0.340 -1.930 ;
        RECT 5.410 -2.020 5.580 -1.160 ;
        RECT 5.250 -2.280 5.580 -2.020 ;
        RECT -2.050 -2.870 -1.700 -2.790 ;
        RECT 5.410 -2.850 5.580 -2.280 ;
        RECT 6.240 -1.250 6.420 -1.060 ;
        RECT 6.240 -2.860 6.410 -1.250 ;
        RECT 6.600 -2.060 6.890 -1.730 ;
        RECT 6.610 -2.350 6.810 -2.060 ;
        RECT 6.610 -2.360 6.800 -2.350 ;
        RECT 6.970 -2.530 7.180 -2.520 ;
        RECT -2.050 -3.720 3.000 -2.870 ;
        RECT 6.960 -3.110 7.180 -2.530 ;
        RECT 6.970 -3.140 7.180 -3.110 ;
        RECT 5.160 -3.410 5.690 -3.240 ;
        RECT 6.970 -3.490 7.170 -3.140 ;
      LAYER mcon ;
        RECT 6.980 1.350 7.150 1.520 ;
        RECT -1.950 0.930 -1.780 1.100 ;
        RECT 0.140 0.770 0.310 0.940 ;
        RECT -3.520 0.170 -3.250 0.440 ;
        RECT 0.140 0.320 0.310 0.490 ;
        RECT 5.310 0.520 5.480 0.690 ;
        RECT 6.620 0.510 6.800 0.700 ;
        RECT -1.100 -0.940 -0.930 -0.770 ;
        RECT -3.520 -1.560 -3.250 -1.290 ;
        RECT 0.140 -2.180 0.310 -2.010 ;
        RECT 5.310 -2.240 5.480 -2.070 ;
        RECT -1.980 -2.760 -1.810 -2.590 ;
        RECT 0.140 -2.630 0.310 -2.460 ;
        RECT 6.620 -2.290 6.800 -2.100 ;
        RECT 6.980 -3.110 7.150 -2.940 ;
      LAYER met1 ;
        RECT 5.090 1.410 5.400 1.850 ;
        RECT -2.020 0.860 -1.700 1.180 ;
        RECT 5.240 0.450 5.560 0.770 ;
        RECT 6.210 -0.340 6.450 -0.210 ;
        RECT 6.210 -0.660 6.470 -0.340 ;
        RECT 6.210 -1.260 6.470 -0.940 ;
        RECT 6.210 -1.380 6.450 -1.260 ;
        RECT 5.240 -2.310 5.560 -1.990 ;
        RECT -2.050 -2.830 -1.730 -2.510 ;
        RECT 5.090 -3.440 5.400 -3.000 ;
      LAYER via ;
        RECT 5.120 1.440 5.380 1.700 ;
        RECT -1.990 0.890 -1.730 1.150 ;
        RECT 5.270 0.480 5.530 0.740 ;
        RECT 6.210 -0.630 6.470 -0.370 ;
        RECT 6.210 -1.230 6.470 -0.970 ;
        RECT 5.270 -2.280 5.530 -2.020 ;
        RECT -2.020 -2.800 -1.760 -2.540 ;
        RECT 5.120 -3.290 5.380 -3.030 ;
  END
END sky130_hilas_FGBiasWeakGate2x1cell

MACRO sky130_hilas_swc4x1cellOverlap
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc4x1cellOverlap ;
  ORIGIN 2.640 4.130 ;
  SIZE 10.080 BY 6.710 ;
  OBS
      LAYER nwell ;
        RECT 2.230 2.290 4.950 2.520 ;
        RECT -2.630 -3.820 -0.900 2.230 ;
        RECT 2.230 -0.570 7.440 2.290 ;
        RECT 2.220 -3.870 7.440 -0.570 ;
        RECT 2.220 -4.070 4.940 -3.870 ;
      LAYER li1 ;
        RECT 2.630 0.950 4.580 2.120 ;
        RECT 4.980 1.820 5.300 1.830 ;
        RECT 4.980 1.650 5.560 1.820 ;
        RECT 4.980 1.600 5.310 1.650 ;
        RECT 4.980 1.570 5.300 1.600 ;
        RECT 6.840 1.550 7.040 1.900 ;
        RECT 4.980 1.240 5.300 1.280 ;
        RECT 4.980 1.200 5.310 1.240 ;
        RECT 4.980 1.030 5.560 1.200 ;
        RECT 4.980 1.020 5.300 1.030 ;
        RECT 6.110 0.930 6.310 1.530 ;
        RECT 6.840 1.520 7.050 1.550 ;
        RECT 6.830 0.930 7.050 1.520 ;
        RECT 2.630 -0.580 4.580 0.590 ;
        RECT 4.980 0.390 5.300 0.400 ;
        RECT 4.980 0.220 5.560 0.390 ;
        RECT 4.980 0.180 5.310 0.220 ;
        RECT 4.980 0.140 5.300 0.180 ;
        RECT 6.110 -0.110 6.310 0.490 ;
        RECT 6.830 -0.100 7.050 0.490 ;
        RECT 6.840 -0.130 7.050 -0.100 ;
        RECT 4.980 -0.180 5.300 -0.150 ;
        RECT 4.980 -0.230 5.310 -0.180 ;
        RECT 4.980 -0.400 5.560 -0.230 ;
        RECT 4.980 -0.410 5.300 -0.400 ;
        RECT 6.840 -0.480 7.040 -0.130 ;
        RECT -2.210 -1.020 -1.660 -0.590 ;
        RECT 6.230 -0.880 6.670 -0.710 ;
        RECT 2.620 -2.140 4.570 -0.970 ;
        RECT 4.980 -1.190 5.300 -1.180 ;
        RECT 4.980 -1.360 5.560 -1.190 ;
        RECT 4.980 -1.410 5.310 -1.360 ;
        RECT 4.980 -1.440 5.300 -1.410 ;
        RECT 6.840 -1.460 7.040 -1.110 ;
        RECT 4.980 -1.770 5.300 -1.730 ;
        RECT 4.980 -1.810 5.310 -1.770 ;
        RECT 4.980 -1.980 5.560 -1.810 ;
        RECT 4.980 -1.990 5.300 -1.980 ;
        RECT 6.110 -2.080 6.310 -1.480 ;
        RECT 6.840 -1.490 7.050 -1.460 ;
        RECT 6.830 -2.080 7.050 -1.490 ;
        RECT 2.620 -3.680 4.570 -2.510 ;
        RECT 4.980 -2.610 5.300 -2.600 ;
        RECT 4.980 -2.780 5.560 -2.610 ;
        RECT 4.980 -2.820 5.310 -2.780 ;
        RECT 4.980 -2.860 5.300 -2.820 ;
        RECT 6.110 -3.110 6.310 -2.510 ;
        RECT 6.830 -3.100 7.050 -2.510 ;
        RECT 6.840 -3.130 7.050 -3.100 ;
        RECT 4.980 -3.180 5.300 -3.150 ;
        RECT 4.980 -3.230 5.310 -3.180 ;
        RECT 4.980 -3.400 5.560 -3.230 ;
        RECT 4.980 -3.410 5.300 -3.400 ;
        RECT 6.840 -3.480 7.040 -3.130 ;
      LAYER mcon ;
        RECT 3.110 1.780 3.280 1.950 ;
        RECT 3.110 1.440 3.280 1.610 ;
        RECT 5.040 1.610 5.210 1.780 ;
        RECT 6.120 1.320 6.290 1.490 ;
        RECT 3.110 1.100 3.280 1.270 ;
        RECT 5.040 1.060 5.210 1.230 ;
        RECT 6.850 1.350 7.020 1.520 ;
        RECT 3.110 0.250 3.280 0.420 ;
        RECT 5.040 0.190 5.210 0.360 ;
        RECT 3.110 -0.090 3.280 0.080 ;
        RECT 6.120 -0.070 6.290 0.100 ;
        RECT 6.850 -0.100 7.020 0.070 ;
        RECT 3.110 -0.430 3.280 -0.260 ;
        RECT 5.040 -0.360 5.210 -0.190 ;
        RECT -2.210 -0.940 -1.940 -0.670 ;
        RECT 6.490 -0.880 6.670 -0.710 ;
        RECT 3.100 -1.310 3.270 -1.140 ;
        RECT 5.040 -1.400 5.210 -1.230 ;
        RECT 3.100 -1.650 3.270 -1.480 ;
        RECT 6.120 -1.690 6.290 -1.520 ;
        RECT 3.100 -1.990 3.270 -1.820 ;
        RECT 5.040 -1.950 5.210 -1.780 ;
        RECT 6.850 -1.660 7.020 -1.490 ;
        RECT 3.100 -2.850 3.270 -2.680 ;
        RECT 5.040 -2.810 5.210 -2.640 ;
        RECT 3.100 -3.190 3.270 -3.020 ;
        RECT 6.120 -3.070 6.290 -2.900 ;
        RECT 6.850 -3.100 7.020 -2.930 ;
        RECT 3.100 -3.530 3.270 -3.360 ;
        RECT 5.040 -3.360 5.210 -3.190 ;
      LAYER met1 ;
        RECT -2.280 -3.820 -1.880 2.170 ;
        RECT 3.070 1.530 3.330 2.010 ;
        RECT 4.970 1.540 5.290 1.860 ;
        RECT 6.110 1.550 6.270 2.280 ;
        RECT 6.110 1.530 6.310 1.550 ;
        RECT 3.060 1.010 3.330 1.530 ;
        RECT 3.060 0.560 3.320 1.010 ;
        RECT 4.970 0.990 5.290 1.310 ;
        RECT 6.090 1.290 6.320 1.530 ;
        RECT 6.110 1.240 6.320 1.290 ;
        RECT 6.480 1.240 6.670 2.230 ;
        RECT 6.920 1.580 7.080 2.280 ;
        RECT 3.070 0.000 3.330 0.480 ;
        RECT 4.970 0.110 5.290 0.430 ;
        RECT 6.110 0.180 6.270 1.240 ;
        RECT 6.500 1.120 6.670 1.240 ;
        RECT 6.510 0.300 6.670 1.120 ;
        RECT 6.810 1.030 7.080 1.580 ;
        RECT 6.810 0.980 7.090 1.030 ;
        RECT 6.920 0.890 7.090 0.980 ;
        RECT 6.920 0.530 7.080 0.890 ;
        RECT 6.920 0.440 7.090 0.530 ;
        RECT 6.500 0.180 6.670 0.300 ;
        RECT 6.110 0.130 6.320 0.180 ;
        RECT 3.060 -0.520 3.330 0.000 ;
        RECT 6.090 -0.110 6.320 0.130 ;
        RECT 4.970 -0.440 5.290 -0.120 ;
        RECT 6.110 -0.130 6.310 -0.110 ;
        RECT 3.060 -0.970 3.320 -0.520 ;
        RECT 3.060 -1.560 3.320 -1.080 ;
        RECT 4.970 -1.470 5.290 -1.150 ;
        RECT 6.110 -1.460 6.270 -0.130 ;
        RECT 6.480 -0.680 6.670 0.180 ;
        RECT 6.810 0.390 7.090 0.440 ;
        RECT 6.810 -0.160 7.080 0.390 ;
        RECT 6.460 -0.910 6.700 -0.680 ;
        RECT 6.110 -1.480 6.310 -1.460 ;
        RECT 3.050 -2.080 3.320 -1.560 ;
        RECT 4.970 -2.020 5.290 -1.700 ;
        RECT 6.090 -1.720 6.320 -1.480 ;
        RECT 6.110 -1.770 6.320 -1.720 ;
        RECT 6.480 -1.770 6.670 -0.910 ;
        RECT 6.920 -1.430 7.080 -0.160 ;
        RECT 3.050 -2.530 3.310 -2.080 ;
        RECT 3.060 -3.100 3.320 -2.620 ;
        RECT 4.970 -2.890 5.290 -2.570 ;
        RECT 6.110 -2.820 6.270 -1.770 ;
        RECT 6.500 -1.890 6.670 -1.770 ;
        RECT 6.510 -2.700 6.670 -1.890 ;
        RECT 6.810 -1.980 7.080 -1.430 ;
        RECT 6.810 -2.030 7.090 -1.980 ;
        RECT 6.920 -2.120 7.090 -2.030 ;
        RECT 6.920 -2.470 7.080 -2.120 ;
        RECT 6.920 -2.560 7.090 -2.470 ;
        RECT 6.500 -2.820 6.670 -2.700 ;
        RECT 6.110 -2.870 6.320 -2.820 ;
        RECT 3.050 -3.620 3.320 -3.100 ;
        RECT 6.090 -3.110 6.320 -2.870 ;
        RECT 4.970 -3.440 5.290 -3.120 ;
        RECT 6.110 -3.130 6.310 -3.110 ;
        RECT 3.050 -4.070 3.310 -3.620 ;
        RECT 6.110 -3.860 6.270 -3.130 ;
        RECT 6.480 -3.810 6.670 -2.820 ;
        RECT 6.810 -2.610 7.090 -2.560 ;
        RECT 6.810 -3.160 7.080 -2.610 ;
        RECT 6.920 -3.860 7.080 -3.160 ;
      LAYER via ;
        RECT 5.000 1.570 5.260 1.830 ;
        RECT 5.000 1.020 5.260 1.280 ;
        RECT 5.000 0.140 5.260 0.400 ;
        RECT 5.000 -0.410 5.260 -0.150 ;
        RECT 5.000 -1.440 5.260 -1.180 ;
        RECT 5.000 -1.990 5.260 -1.730 ;
        RECT 5.000 -2.860 5.260 -2.600 ;
        RECT 5.000 -3.410 5.260 -3.150 ;
      LAYER met2 ;
        RECT 4.970 1.730 5.280 1.870 ;
        RECT -2.640 1.550 7.440 1.730 ;
        RECT 4.970 1.540 5.280 1.550 ;
        RECT 4.970 1.300 5.280 1.320 ;
        RECT -2.640 1.120 7.440 1.300 ;
        RECT 4.970 0.990 5.280 1.120 ;
        RECT 4.970 0.300 5.280 0.430 ;
        RECT -2.640 0.120 7.440 0.300 ;
        RECT 4.970 0.100 5.280 0.120 ;
        RECT 4.970 -0.130 5.280 -0.120 ;
        RECT -2.640 -0.200 4.960 -0.130 ;
        RECT 4.970 -0.200 7.440 -0.130 ;
        RECT -2.640 -0.310 7.440 -0.200 ;
        RECT 4.970 -0.450 5.280 -0.310 ;
        RECT 4.970 -1.280 5.280 -1.140 ;
        RECT 4.970 -1.290 7.440 -1.280 ;
        RECT -2.620 -1.460 7.440 -1.290 ;
        RECT 4.970 -1.470 5.280 -1.460 ;
        RECT 4.970 -1.710 5.280 -1.690 ;
        RECT -2.620 -1.880 7.440 -1.710 ;
        RECT 4.880 -1.890 7.440 -1.880 ;
        RECT 4.970 -2.020 5.280 -1.890 ;
        RECT 4.970 -2.690 5.280 -2.570 ;
        RECT -2.620 -2.700 5.280 -2.690 ;
        RECT -2.620 -2.860 7.440 -2.700 ;
        RECT -1.840 -2.950 -0.300 -2.860 ;
        RECT 4.880 -2.880 7.440 -2.860 ;
        RECT 4.970 -2.900 5.280 -2.880 ;
        RECT 4.970 -3.130 5.280 -3.120 ;
        RECT -2.620 -3.300 7.440 -3.130 ;
        RECT 4.970 -3.310 7.440 -3.300 ;
        RECT 4.970 -3.450 5.280 -3.310 ;
  END
END sky130_hilas_swc4x1cellOverlap

MACRO sky130_hilas_nFETLarge
  CLASS BLOCK ;
  FOREIGN sky130_hilas_nFETLarge ;
  ORIGIN -0.640 -4.200 ;
  SIZE 4.370 BY 5.830 ;
  PIN GATE
    USE ANALOG ;
    ANTENNAGATEAREA 6.396000 ;
    PORT
      LAYER met2 ;
        RECT 0.640 4.530 1.240 5.020 ;
        RECT 0.640 4.200 1.250 4.530 ;
    END
  END GATE
  PIN SOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 4.231200 ;
    PORT
      LAYER met2 ;
        RECT 0.970 9.790 4.030 9.800 ;
        RECT 0.880 9.460 4.030 9.790 ;
        RECT 0.880 7.010 1.200 9.460 ;
        RECT 3.700 9.450 4.010 9.460 ;
        RECT 0.880 6.680 4.040 7.010 ;
        RECT 0.880 5.640 1.200 6.680 ;
        RECT 0.880 5.320 4.040 5.640 ;
        RECT 1.500 5.310 1.810 5.320 ;
        RECT 2.600 5.310 2.910 5.320 ;
        RECT 3.700 5.310 4.010 5.320 ;
    END
  END SOURCE
  PIN DRAIN
    USE ANALOG ;
    ANTENNADIFFAREA 4.231200 ;
    PORT
      LAYER met2 ;
        RECT 2.060 9.080 2.370 9.110 ;
        RECT 3.150 9.080 3.460 9.090 ;
        RECT 2.060 8.780 5.010 9.080 ;
        RECT 3.150 8.760 3.460 8.780 ;
        RECT 4.260 8.740 5.010 8.780 ;
        RECT 4.630 8.610 5.010 8.740 ;
        RECT 4.660 7.740 5.010 8.610 ;
        RECT 2.060 7.410 5.010 7.740 ;
        RECT 4.660 4.970 5.010 7.410 ;
        RECT 2.070 4.960 5.010 4.970 ;
        RECT 2.060 4.650 5.010 4.960 ;
        RECT 2.060 4.640 4.780 4.650 ;
        RECT 2.060 4.630 2.370 4.640 ;
        RECT 3.150 4.630 3.460 4.640 ;
    END
  END DRAIN
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.820 6.650 1.090 6.680 ;
        RECT 0.820 6.120 1.100 6.650 ;
        RECT 0.640 5.820 1.100 6.120 ;
        RECT 0.640 5.800 1.110 5.820 ;
        RECT 0.820 5.370 1.110 5.800 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.590 9.750 1.760 9.780 ;
        RECT 1.520 9.710 1.840 9.750 ;
        RECT 1.520 9.520 1.850 9.710 ;
        RECT 1.520 9.490 1.840 9.520 ;
        RECT 1.590 6.970 1.760 9.490 ;
        RECT 2.140 9.070 2.310 9.780 ;
        RECT 2.690 9.750 2.860 9.780 ;
        RECT 2.610 9.710 2.930 9.750 ;
        RECT 2.610 9.520 2.940 9.710 ;
        RECT 2.610 9.490 2.930 9.520 ;
        RECT 2.070 9.030 2.390 9.070 ;
        RECT 2.070 8.840 2.400 9.030 ;
        RECT 2.070 8.810 2.390 8.840 ;
        RECT 2.140 7.700 2.310 8.810 ;
        RECT 2.070 7.660 2.390 7.700 ;
        RECT 2.070 7.470 2.400 7.660 ;
        RECT 2.070 7.440 2.390 7.470 ;
        RECT 1.510 6.930 1.830 6.970 ;
        RECT 1.510 6.740 1.840 6.930 ;
        RECT 1.510 6.710 1.830 6.740 ;
        RECT 0.880 5.400 1.050 6.620 ;
        RECT 1.590 5.600 1.760 6.710 ;
        RECT 1.510 5.560 1.830 5.600 ;
        RECT 1.510 5.370 1.840 5.560 ;
        RECT 1.510 5.340 1.830 5.370 ;
        RECT 0.830 4.950 1.340 5.210 ;
        RECT 0.830 4.880 1.350 4.950 ;
        RECT 0.840 4.200 1.350 4.880 ;
        RECT 1.590 4.600 1.760 5.340 ;
        RECT 2.140 4.920 2.310 7.440 ;
        RECT 2.690 6.970 2.860 9.490 ;
        RECT 3.240 9.050 3.410 9.780 ;
        RECT 3.790 9.740 3.960 9.780 ;
        RECT 3.710 9.700 4.030 9.740 ;
        RECT 3.710 9.510 4.040 9.700 ;
        RECT 3.710 9.480 4.030 9.510 ;
        RECT 3.160 9.010 3.480 9.050 ;
        RECT 3.160 8.820 3.490 9.010 ;
        RECT 3.160 8.790 3.480 8.820 ;
        RECT 3.240 7.700 3.410 8.790 ;
        RECT 3.160 7.660 3.480 7.700 ;
        RECT 3.160 7.470 3.490 7.660 ;
        RECT 3.160 7.440 3.480 7.470 ;
        RECT 2.610 6.930 2.930 6.970 ;
        RECT 2.610 6.740 2.940 6.930 ;
        RECT 2.610 6.710 2.930 6.740 ;
        RECT 2.690 5.600 2.860 6.710 ;
        RECT 2.610 5.560 2.930 5.600 ;
        RECT 2.610 5.370 2.940 5.560 ;
        RECT 2.610 5.340 2.930 5.370 ;
        RECT 2.070 4.880 2.390 4.920 ;
        RECT 2.070 4.690 2.400 4.880 ;
        RECT 2.070 4.660 2.390 4.690 ;
        RECT 2.140 4.600 2.310 4.660 ;
        RECT 2.690 4.600 2.860 5.340 ;
        RECT 3.240 4.920 3.410 7.440 ;
        RECT 3.790 6.970 3.960 9.480 ;
        RECT 4.340 9.040 4.510 9.780 ;
        RECT 4.270 9.000 4.590 9.040 ;
        RECT 4.270 8.810 4.600 9.000 ;
        RECT 4.270 8.780 4.590 8.810 ;
        RECT 4.340 7.700 4.510 8.780 ;
        RECT 4.260 7.660 4.580 7.700 ;
        RECT 4.260 7.470 4.590 7.660 ;
        RECT 4.260 7.440 4.580 7.470 ;
        RECT 3.710 6.930 4.030 6.970 ;
        RECT 3.710 6.740 4.040 6.930 ;
        RECT 3.710 6.710 4.030 6.740 ;
        RECT 3.790 5.600 3.960 6.710 ;
        RECT 3.710 5.560 4.030 5.600 ;
        RECT 3.710 5.370 4.040 5.560 ;
        RECT 3.710 5.340 4.030 5.370 ;
        RECT 3.160 4.880 3.480 4.920 ;
        RECT 3.160 4.690 3.490 4.880 ;
        RECT 3.160 4.660 3.480 4.690 ;
        RECT 3.240 4.600 3.410 4.660 ;
        RECT 3.790 4.600 3.960 5.340 ;
        RECT 4.340 4.930 4.510 7.440 ;
        RECT 4.260 4.890 4.580 4.930 ;
        RECT 4.260 4.700 4.590 4.890 ;
        RECT 4.260 4.670 4.580 4.700 ;
        RECT 4.340 4.600 4.510 4.670 ;
      LAYER mcon ;
        RECT 1.580 9.530 1.750 9.700 ;
        RECT 2.670 9.530 2.840 9.700 ;
        RECT 2.130 8.850 2.300 9.020 ;
        RECT 2.130 7.480 2.300 7.650 ;
        RECT 1.570 6.750 1.740 6.920 ;
        RECT 0.880 6.450 1.050 6.620 ;
        RECT 0.880 6.090 1.050 6.260 ;
        RECT 1.570 5.380 1.740 5.550 ;
        RECT 1.000 4.740 1.170 4.910 ;
        RECT 3.770 9.520 3.940 9.690 ;
        RECT 3.220 8.830 3.390 9.000 ;
        RECT 3.220 7.480 3.390 7.650 ;
        RECT 2.670 6.750 2.840 6.920 ;
        RECT 2.670 5.380 2.840 5.550 ;
        RECT 2.130 4.700 2.300 4.870 ;
        RECT 4.330 8.820 4.500 8.990 ;
        RECT 4.320 7.480 4.490 7.650 ;
        RECT 3.770 6.750 3.940 6.920 ;
        RECT 3.770 5.380 3.940 5.550 ;
        RECT 3.220 4.700 3.390 4.870 ;
        RECT 4.320 4.710 4.490 4.880 ;
        RECT 1.010 4.270 1.180 4.440 ;
      LAYER met1 ;
        RECT 1.510 9.460 1.830 9.780 ;
        RECT 2.600 9.460 2.920 9.780 ;
        RECT 3.700 9.450 4.020 9.770 ;
        RECT 2.060 8.780 2.380 9.100 ;
        RECT 3.150 8.760 3.470 9.080 ;
        RECT 4.260 8.750 4.580 9.070 ;
        RECT 2.060 7.410 2.380 7.730 ;
        RECT 3.150 7.410 3.470 7.730 ;
        RECT 4.250 7.410 4.570 7.730 ;
        RECT 1.500 6.680 1.820 7.000 ;
        RECT 2.600 6.680 2.920 7.000 ;
        RECT 3.700 6.680 4.020 7.000 ;
        RECT 1.500 5.310 1.820 5.630 ;
        RECT 2.600 5.310 2.920 5.630 ;
        RECT 3.700 5.310 4.020 5.630 ;
        RECT 0.930 4.670 1.250 4.990 ;
        RECT 2.060 4.630 2.380 4.950 ;
        RECT 3.150 4.630 3.470 4.950 ;
        RECT 4.250 4.640 4.570 4.960 ;
        RECT 0.940 4.200 1.260 4.520 ;
      LAYER via ;
        RECT 1.540 9.490 1.800 9.750 ;
        RECT 2.630 9.490 2.890 9.750 ;
        RECT 3.730 9.480 3.990 9.740 ;
        RECT 2.090 8.810 2.350 9.070 ;
        RECT 3.180 8.790 3.440 9.050 ;
        RECT 4.290 8.780 4.550 9.040 ;
        RECT 2.090 7.440 2.350 7.700 ;
        RECT 3.180 7.440 3.440 7.700 ;
        RECT 4.280 7.440 4.540 7.700 ;
        RECT 1.530 6.710 1.790 6.970 ;
        RECT 2.630 6.710 2.890 6.970 ;
        RECT 3.730 6.710 3.990 6.970 ;
        RECT 1.530 5.340 1.790 5.600 ;
        RECT 2.630 5.340 2.890 5.600 ;
        RECT 3.730 5.340 3.990 5.600 ;
        RECT 0.960 4.700 1.220 4.960 ;
        RECT 2.090 4.660 2.350 4.920 ;
        RECT 3.180 4.660 3.440 4.920 ;
        RECT 4.280 4.670 4.540 4.930 ;
        RECT 0.970 4.230 1.230 4.490 ;
  END
END sky130_hilas_nFETLarge

MACRO sky130_hilas_pFETLarge
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pFETLarge ;
  ORIGIN -0.640 -4.190 ;
  SIZE 4.640 BY 5.990 ;
  PIN GATE
    ANTENNAGATEAREA 6.526000 ;
    PORT
      LAYER met2 ;
        RECT 0.640 4.530 1.240 5.020 ;
        RECT 0.640 4.200 1.250 4.530 ;
    END
  END GATE
  PIN SOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 4.367400 ;
    PORT
      LAYER met2 ;
        RECT 0.970 9.790 4.030 9.800 ;
        RECT 0.880 9.460 4.030 9.790 ;
        RECT 0.880 7.010 1.200 9.460 ;
        RECT 3.700 9.450 4.010 9.460 ;
        RECT 0.880 6.680 4.040 7.010 ;
        RECT 0.880 5.640 1.200 6.680 ;
        RECT 0.880 5.320 4.040 5.640 ;
        RECT 1.500 5.310 1.810 5.320 ;
        RECT 2.600 5.310 2.910 5.320 ;
        RECT 3.700 5.310 4.010 5.320 ;
    END
  END SOURCE
  PIN DRAIN
    USE ANALOG ;
    ANTENNADIFFAREA 4.317200 ;
    PORT
      LAYER met2 ;
        RECT 2.060 9.080 2.370 9.110 ;
        RECT 3.150 9.080 3.460 9.090 ;
        RECT 2.060 8.780 5.010 9.080 ;
        RECT 3.150 8.760 3.460 8.780 ;
        RECT 4.260 8.740 5.010 8.780 ;
        RECT 4.630 8.610 5.010 8.740 ;
        RECT 4.660 7.740 5.010 8.610 ;
        RECT 2.060 7.410 5.010 7.740 ;
        RECT 4.660 4.970 5.010 7.410 ;
        RECT 2.070 4.960 5.010 4.970 ;
        RECT 2.060 4.650 5.010 4.960 ;
        RECT 2.060 4.640 4.780 4.650 ;
        RECT 2.060 4.630 2.370 4.640 ;
        RECT 3.150 4.630 3.460 4.640 ;
    END
  END DRAIN
  PIN WELL
    USE ANALOG ;
    ANTENNADIFFAREA 0.213200 ;
    PORT
      LAYER nwell ;
        RECT 1.360 4.370 5.280 10.070 ;
      LAYER met1 ;
        RECT 4.780 9.980 5.040 10.180 ;
        RECT 4.780 9.170 5.090 9.980 ;
        RECT 4.780 4.190 5.040 9.170 ;
    END
  END WELL
  OBS
      LAYER li1 ;
        RECT 1.600 9.750 1.770 9.840 ;
        RECT 1.520 9.710 1.840 9.750 ;
        RECT 1.520 9.520 1.850 9.710 ;
        RECT 1.520 9.490 1.840 9.520 ;
        RECT 1.600 6.970 1.770 9.490 ;
        RECT 2.150 9.070 2.320 9.840 ;
        RECT 2.700 9.750 2.870 9.840 ;
        RECT 2.610 9.710 2.930 9.750 ;
        RECT 2.610 9.520 2.940 9.710 ;
        RECT 2.610 9.490 2.930 9.520 ;
        RECT 2.070 9.030 2.390 9.070 ;
        RECT 2.070 8.840 2.400 9.030 ;
        RECT 2.070 8.810 2.390 8.840 ;
        RECT 2.150 7.700 2.320 8.810 ;
        RECT 2.070 7.660 2.390 7.700 ;
        RECT 2.070 7.470 2.400 7.660 ;
        RECT 2.070 7.440 2.390 7.470 ;
        RECT 1.510 6.930 1.830 6.970 ;
        RECT 1.510 6.740 1.840 6.930 ;
        RECT 1.510 6.710 1.830 6.740 ;
        RECT 1.600 5.600 1.770 6.710 ;
        RECT 1.510 5.560 1.830 5.600 ;
        RECT 1.510 5.370 1.840 5.560 ;
        RECT 1.510 5.340 1.830 5.370 ;
        RECT 0.830 5.130 1.340 5.210 ;
        RECT 0.830 4.880 1.350 5.130 ;
        RECT 0.840 4.200 1.350 4.880 ;
        RECT 1.600 4.520 1.770 5.340 ;
        RECT 2.150 4.920 2.320 7.440 ;
        RECT 2.700 6.970 2.870 9.490 ;
        RECT 3.250 9.050 3.420 9.840 ;
        RECT 3.800 9.740 3.970 9.840 ;
        RECT 3.710 9.700 4.030 9.740 ;
        RECT 3.710 9.510 4.040 9.700 ;
        RECT 3.710 9.480 4.030 9.510 ;
        RECT 3.160 9.010 3.480 9.050 ;
        RECT 3.160 8.820 3.490 9.010 ;
        RECT 3.160 8.790 3.480 8.820 ;
        RECT 3.250 7.700 3.420 8.790 ;
        RECT 3.160 7.660 3.480 7.700 ;
        RECT 3.160 7.470 3.490 7.660 ;
        RECT 3.160 7.440 3.480 7.470 ;
        RECT 2.610 6.930 2.930 6.970 ;
        RECT 2.610 6.740 2.940 6.930 ;
        RECT 2.610 6.710 2.930 6.740 ;
        RECT 2.700 5.600 2.870 6.710 ;
        RECT 2.610 5.560 2.930 5.600 ;
        RECT 2.610 5.370 2.940 5.560 ;
        RECT 2.610 5.340 2.930 5.370 ;
        RECT 2.070 4.880 2.390 4.920 ;
        RECT 2.070 4.690 2.400 4.880 ;
        RECT 2.070 4.660 2.390 4.690 ;
        RECT 2.150 4.510 2.320 4.660 ;
        RECT 2.700 4.510 2.870 5.340 ;
        RECT 3.250 4.920 3.420 7.440 ;
        RECT 3.800 6.970 3.970 9.480 ;
        RECT 4.350 9.040 4.520 9.840 ;
        RECT 4.890 9.110 5.060 9.870 ;
        RECT 4.270 9.000 4.590 9.040 ;
        RECT 4.270 8.810 4.600 9.000 ;
        RECT 4.270 8.780 4.590 8.810 ;
        RECT 4.350 7.700 4.520 8.780 ;
        RECT 4.260 7.660 4.580 7.700 ;
        RECT 4.260 7.470 4.590 7.660 ;
        RECT 4.260 7.440 4.580 7.470 ;
        RECT 3.710 6.930 4.030 6.970 ;
        RECT 3.710 6.740 4.040 6.930 ;
        RECT 3.710 6.710 4.030 6.740 ;
        RECT 3.800 5.600 3.970 6.710 ;
        RECT 3.710 5.560 4.030 5.600 ;
        RECT 3.710 5.370 4.040 5.560 ;
        RECT 3.710 5.340 4.030 5.370 ;
        RECT 3.160 4.880 3.480 4.920 ;
        RECT 3.160 4.690 3.490 4.880 ;
        RECT 3.160 4.660 3.480 4.690 ;
        RECT 3.250 4.510 3.420 4.660 ;
        RECT 3.800 4.510 3.970 5.340 ;
        RECT 4.350 4.930 4.520 7.440 ;
        RECT 4.260 4.890 4.580 4.930 ;
        RECT 4.260 4.700 4.590 4.890 ;
        RECT 4.260 4.670 4.580 4.700 ;
        RECT 4.350 4.510 4.520 4.670 ;
      LAYER mcon ;
        RECT 1.580 9.530 1.750 9.700 ;
        RECT 2.670 9.530 2.840 9.700 ;
        RECT 2.130 8.850 2.300 9.020 ;
        RECT 2.130 7.480 2.300 7.650 ;
        RECT 1.570 6.750 1.740 6.920 ;
        RECT 1.570 5.380 1.740 5.550 ;
        RECT 1.000 4.740 1.170 4.910 ;
        RECT 3.770 9.520 3.940 9.690 ;
        RECT 3.220 8.830 3.390 9.000 ;
        RECT 3.220 7.480 3.390 7.650 ;
        RECT 2.670 6.750 2.840 6.920 ;
        RECT 2.670 5.380 2.840 5.550 ;
        RECT 2.130 4.700 2.300 4.870 ;
        RECT 4.890 9.700 5.060 9.870 ;
        RECT 4.890 9.340 5.060 9.510 ;
        RECT 4.330 8.820 4.500 8.990 ;
        RECT 4.320 7.480 4.490 7.650 ;
        RECT 3.770 6.750 3.940 6.920 ;
        RECT 3.770 5.380 3.940 5.550 ;
        RECT 3.220 4.700 3.390 4.870 ;
        RECT 4.320 4.710 4.490 4.880 ;
        RECT 1.010 4.270 1.180 4.440 ;
      LAYER met1 ;
        RECT 1.510 9.460 1.830 9.780 ;
        RECT 2.600 9.460 2.920 9.780 ;
        RECT 3.700 9.450 4.020 9.770 ;
        RECT 2.060 8.780 2.380 9.100 ;
        RECT 3.150 8.760 3.470 9.080 ;
        RECT 4.260 8.750 4.580 9.070 ;
        RECT 2.060 7.410 2.380 7.730 ;
        RECT 3.150 7.410 3.470 7.730 ;
        RECT 4.250 7.410 4.570 7.730 ;
        RECT 1.500 6.680 1.820 7.000 ;
        RECT 2.600 6.680 2.920 7.000 ;
        RECT 3.700 6.680 4.020 7.000 ;
        RECT 1.500 5.310 1.820 5.630 ;
        RECT 2.600 5.310 2.920 5.630 ;
        RECT 3.700 5.310 4.020 5.630 ;
        RECT 0.930 4.670 1.250 4.990 ;
        RECT 2.060 4.630 2.380 4.950 ;
        RECT 3.150 4.630 3.470 4.950 ;
        RECT 4.250 4.640 4.570 4.960 ;
        RECT 0.940 4.200 1.260 4.520 ;
      LAYER via ;
        RECT 1.540 9.490 1.800 9.750 ;
        RECT 2.630 9.490 2.890 9.750 ;
        RECT 3.730 9.480 3.990 9.740 ;
        RECT 2.090 8.810 2.350 9.070 ;
        RECT 3.180 8.790 3.440 9.050 ;
        RECT 4.290 8.780 4.550 9.040 ;
        RECT 2.090 7.440 2.350 7.700 ;
        RECT 3.180 7.440 3.440 7.700 ;
        RECT 4.280 7.440 4.540 7.700 ;
        RECT 1.530 6.710 1.790 6.970 ;
        RECT 2.630 6.710 2.890 6.970 ;
        RECT 3.730 6.710 3.990 6.970 ;
        RECT 1.530 5.340 1.790 5.600 ;
        RECT 2.630 5.340 2.890 5.600 ;
        RECT 3.730 5.340 3.990 5.600 ;
        RECT 0.960 4.700 1.220 4.960 ;
        RECT 2.090 4.660 2.350 4.920 ;
        RECT 3.180 4.660 3.440 4.920 ;
        RECT 4.280 4.670 4.540 4.930 ;
        RECT 0.970 4.230 1.230 4.490 ;
  END
END sky130_hilas_pFETLarge

MACRO sky130_hilas_polyresistorGND
  CLASS BLOCK ;
  FOREIGN sky130_hilas_polyresistorGND ;
  ORIGIN 27.490 0.570 ;
  SIZE 55.470 BY 10.890 ;
  PIN INPUT
    PORT
      LAYER met1 ;
        RECT -6.430 9.680 -4.020 10.320 ;
        RECT -6.410 8.330 -6.000 9.680 ;
    END
  END INPUT
  PIN OUTPUT
    ANTENNADIFFAREA 16.452000 ;
    PORT
      LAYER met2 ;
        RECT -27.490 6.810 27.980 8.200 ;
    END
  END OUTPUT
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.320 9.020 0.730 9.790 ;
        RECT 0.050 8.750 0.730 9.020 ;
        RECT 0.050 8.320 1.740 8.750 ;
        RECT -27.160 8.140 -2.790 8.160 ;
        RECT -27.220 7.750 -2.790 8.140 ;
        RECT -27.220 -0.500 -26.810 7.750 ;
        RECT -0.620 0.250 1.740 8.320 ;
        RECT 6.010 8.150 27.370 8.160 ;
        RECT 5.950 7.760 27.370 8.150 ;
        RECT 5.950 7.750 27.210 7.760 ;
        RECT -0.740 -0.570 1.740 0.250 ;
      LAYER via ;
        RECT -26.670 7.840 -2.870 8.100 ;
        RECT 6.010 7.840 26.870 8.100 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT -6.350 8.550 -6.130 9.670 ;
        RECT -6.400 8.360 -6.070 8.550 ;
        RECT 0.390 8.360 0.630 9.710 ;
        RECT -27.110 7.890 27.630 8.160 ;
        RECT -27.110 7.760 -2.770 7.890 ;
        RECT 5.920 7.760 27.630 7.890 ;
        RECT -27.110 0.160 -26.940 7.760 ;
        RECT 27.460 0.680 27.630 7.760 ;
        RECT -0.670 -0.180 1.690 -0.010 ;
      LAYER mcon ;
        RECT -6.320 9.470 -6.150 9.640 ;
        RECT -6.320 9.110 -6.150 9.280 ;
        RECT -6.320 8.750 -6.150 8.920 ;
        RECT -6.320 8.390 -6.150 8.560 ;
        RECT 0.430 9.300 0.600 9.470 ;
        RECT 0.430 8.940 0.600 9.110 ;
        RECT 0.430 8.580 0.600 8.750 ;
        RECT -26.770 7.780 -2.870 7.950 ;
        RECT 6.010 7.780 27.180 7.950 ;
        RECT -0.300 -0.180 -0.130 -0.010 ;
        RECT 0.070 -0.180 0.240 -0.010 ;
        RECT 0.430 -0.180 0.600 -0.010 ;
        RECT 0.790 -0.180 0.960 -0.010 ;
        RECT 1.150 -0.180 1.330 -0.010 ;
        RECT 1.520 -0.180 1.690 -0.010 ;
      LAYER met2 ;
        RECT -27.490 0.510 27.980 1.910 ;
  END
END sky130_hilas_polyresistorGND

MACRO sky130_hilas_LevelShift4InputUp
  CLASS BLOCK ;
  FOREIGN sky130_hilas_LevelShift4InputUp ;
  ORIGIN 0.300 1.060 ;
  SIZE 8.700 BY 7.000 ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 6.070 -1.060 7.840 5.940 ;
      LAYER met1 ;
        RECT 7.360 -1.060 7.600 5.940 ;
    END
  END VPWR
  PIN VINJ
    ANTENNADIFFAREA 1.900800 ;
    PORT
      LAYER nwell ;
        RECT -0.300 -1.060 2.200 5.940 ;
      LAYER met1 ;
        RECT 0.040 -1.060 0.330 5.940 ;
    END
  END VINJ
  PIN OUTPUT4
    ANTENNAGATEAREA 0.180000 ;
    ANTENNADIFFAREA 0.223200 ;
    PORT
      LAYER met2 ;
        RECT 1.080 0.250 1.400 0.300 ;
        RECT 2.110 0.260 2.430 0.270 ;
        RECT 2.110 0.250 2.440 0.260 ;
        RECT -0.230 0.050 2.440 0.250 ;
        RECT 1.080 0.040 1.400 0.050 ;
        RECT 2.110 0.000 2.440 0.050 ;
        RECT 2.110 -0.020 2.430 0.000 ;
    END
  END OUTPUT4
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 4.350 -1.060 4.660 5.940 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.980 5.430 1.430 5.580 ;
        RECT 0.040 5.250 0.370 5.420 ;
        RECT 0.830 5.260 1.430 5.430 ;
        RECT 0.110 4.790 0.290 5.250 ;
        RECT 1.630 4.820 1.800 5.580 ;
        RECT 2.130 5.490 2.420 5.510 ;
        RECT 2.130 5.450 2.590 5.490 ;
        RECT 2.130 5.430 3.570 5.450 ;
        RECT 2.130 5.270 3.610 5.430 ;
        RECT 2.420 5.260 3.610 5.270 ;
        RECT 4.060 5.400 4.520 5.430 ;
        RECT 5.830 5.400 6.180 5.500 ;
        RECT 4.060 5.260 5.170 5.400 ;
        RECT 4.350 5.230 5.170 5.260 ;
        RECT 5.410 5.230 6.580 5.400 ;
        RECT 6.830 5.230 7.590 5.400 ;
        RECT 4.350 5.090 4.610 5.230 ;
        RECT 3.430 4.920 4.610 5.090 ;
        RECT 7.360 5.220 7.590 5.230 ;
        RECT 1.630 4.810 2.010 4.820 ;
        RECT 0.110 4.620 1.070 4.790 ;
        RECT 1.540 4.750 2.010 4.810 ;
        RECT 1.540 4.640 2.880 4.750 ;
        RECT 1.620 4.580 2.880 4.640 ;
        RECT 1.620 4.530 2.010 4.580 ;
        RECT 3.430 4.480 3.610 4.920 ;
        RECT 4.350 4.780 4.610 4.920 ;
        RECT 5.820 4.780 6.150 5.040 ;
        RECT 7.360 4.780 7.630 5.220 ;
        RECT 3.850 4.420 4.060 4.750 ;
        RECT 4.350 4.610 4.680 4.780 ;
        RECT 4.920 4.610 7.080 4.780 ;
        RECT 4.350 4.560 4.520 4.610 ;
        RECT 7.330 4.600 7.660 4.780 ;
        RECT 8.010 4.640 8.180 4.700 ;
        RECT 7.990 4.420 8.210 4.640 ;
        RECT 8.010 4.370 8.180 4.420 ;
        RECT 0.980 3.680 1.430 3.830 ;
        RECT 0.040 3.500 0.370 3.670 ;
        RECT 0.830 3.510 1.430 3.680 ;
        RECT 0.110 3.040 0.290 3.500 ;
        RECT 1.630 3.070 1.800 3.830 ;
        RECT 2.130 3.740 2.420 3.760 ;
        RECT 2.130 3.700 2.590 3.740 ;
        RECT 2.130 3.680 3.570 3.700 ;
        RECT 2.130 3.520 3.610 3.680 ;
        RECT 2.420 3.510 3.610 3.520 ;
        RECT 4.060 3.650 4.520 3.680 ;
        RECT 5.830 3.650 6.180 3.750 ;
        RECT 4.060 3.510 5.170 3.650 ;
        RECT 4.350 3.480 5.170 3.510 ;
        RECT 5.410 3.480 6.580 3.650 ;
        RECT 6.830 3.480 7.590 3.650 ;
        RECT 4.350 3.340 4.610 3.480 ;
        RECT 3.430 3.170 4.610 3.340 ;
        RECT 7.360 3.470 7.590 3.480 ;
        RECT 1.630 3.060 2.010 3.070 ;
        RECT 0.110 2.870 1.070 3.040 ;
        RECT 1.540 3.000 2.010 3.060 ;
        RECT 1.540 2.890 2.880 3.000 ;
        RECT 1.620 2.830 2.880 2.890 ;
        RECT 1.620 2.780 2.010 2.830 ;
        RECT 3.430 2.730 3.610 3.170 ;
        RECT 4.350 3.030 4.610 3.170 ;
        RECT 5.820 3.030 6.150 3.290 ;
        RECT 7.360 3.030 7.630 3.470 ;
        RECT 3.850 2.670 4.060 3.000 ;
        RECT 4.350 2.860 4.680 3.030 ;
        RECT 4.920 2.860 7.080 3.030 ;
        RECT 4.350 2.810 4.520 2.860 ;
        RECT 7.330 2.850 7.660 3.030 ;
        RECT 8.010 2.890 8.180 2.950 ;
        RECT 7.990 2.670 8.210 2.890 ;
        RECT 8.010 2.620 8.180 2.670 ;
        RECT 0.980 1.930 1.430 2.080 ;
        RECT 0.040 1.750 0.370 1.920 ;
        RECT 0.830 1.760 1.430 1.930 ;
        RECT 0.110 1.290 0.290 1.750 ;
        RECT 1.630 1.320 1.800 2.080 ;
        RECT 2.130 1.990 2.420 2.010 ;
        RECT 2.130 1.950 2.590 1.990 ;
        RECT 2.130 1.930 3.570 1.950 ;
        RECT 2.130 1.770 3.610 1.930 ;
        RECT 2.420 1.760 3.610 1.770 ;
        RECT 4.060 1.900 4.520 1.930 ;
        RECT 5.830 1.900 6.180 2.000 ;
        RECT 4.060 1.760 5.170 1.900 ;
        RECT 4.350 1.730 5.170 1.760 ;
        RECT 5.410 1.730 6.580 1.900 ;
        RECT 6.830 1.730 7.590 1.900 ;
        RECT 4.350 1.590 4.610 1.730 ;
        RECT 3.430 1.420 4.610 1.590 ;
        RECT 7.360 1.720 7.590 1.730 ;
        RECT 1.630 1.310 2.010 1.320 ;
        RECT 0.110 1.120 1.070 1.290 ;
        RECT 1.540 1.250 2.010 1.310 ;
        RECT 1.540 1.140 2.880 1.250 ;
        RECT 1.620 1.080 2.880 1.140 ;
        RECT 1.620 1.030 2.010 1.080 ;
        RECT 3.430 0.980 3.610 1.420 ;
        RECT 4.350 1.280 4.610 1.420 ;
        RECT 5.820 1.280 6.150 1.540 ;
        RECT 7.360 1.280 7.630 1.720 ;
        RECT 3.850 0.920 4.060 1.250 ;
        RECT 4.350 1.110 4.680 1.280 ;
        RECT 4.920 1.110 7.080 1.280 ;
        RECT 4.350 1.060 4.520 1.110 ;
        RECT 7.330 1.100 7.660 1.280 ;
        RECT 8.010 1.140 8.180 1.200 ;
        RECT 7.990 0.920 8.210 1.140 ;
        RECT 8.010 0.870 8.180 0.920 ;
        RECT 0.980 0.180 1.430 0.330 ;
        RECT 0.040 0.000 0.370 0.170 ;
        RECT 0.830 0.010 1.430 0.180 ;
        RECT 0.110 -0.460 0.290 0.000 ;
        RECT 1.630 -0.430 1.800 0.330 ;
        RECT 2.130 0.240 2.420 0.260 ;
        RECT 2.130 0.200 2.590 0.240 ;
        RECT 2.130 0.180 3.570 0.200 ;
        RECT 2.130 0.020 3.610 0.180 ;
        RECT 2.420 0.010 3.610 0.020 ;
        RECT 4.060 0.150 4.520 0.180 ;
        RECT 5.830 0.150 6.180 0.250 ;
        RECT 4.060 0.010 5.170 0.150 ;
        RECT 4.350 -0.020 5.170 0.010 ;
        RECT 5.410 -0.020 6.580 0.150 ;
        RECT 6.830 -0.020 7.590 0.150 ;
        RECT 4.350 -0.160 4.610 -0.020 ;
        RECT 3.430 -0.330 4.610 -0.160 ;
        RECT 7.360 -0.030 7.590 -0.020 ;
        RECT 1.630 -0.440 2.010 -0.430 ;
        RECT 0.110 -0.630 1.070 -0.460 ;
        RECT 1.540 -0.500 2.010 -0.440 ;
        RECT 1.540 -0.610 2.880 -0.500 ;
        RECT 1.620 -0.670 2.880 -0.610 ;
        RECT 1.620 -0.720 2.010 -0.670 ;
        RECT 3.430 -0.770 3.610 -0.330 ;
        RECT 4.350 -0.470 4.610 -0.330 ;
        RECT 5.820 -0.470 6.150 -0.210 ;
        RECT 7.360 -0.470 7.630 -0.030 ;
        RECT 3.850 -0.830 4.060 -0.500 ;
        RECT 4.350 -0.640 4.680 -0.470 ;
        RECT 4.920 -0.640 7.080 -0.470 ;
        RECT 4.350 -0.690 4.520 -0.640 ;
        RECT 7.330 -0.650 7.660 -0.470 ;
        RECT 8.010 -0.610 8.180 -0.550 ;
        RECT 7.990 -0.830 8.210 -0.610 ;
        RECT 8.010 -0.880 8.180 -0.830 ;
      LAYER mcon ;
        RECT 1.150 5.330 1.320 5.500 ;
        RECT 0.110 4.990 0.280 5.160 ;
        RECT 2.190 5.290 2.360 5.460 ;
        RECT 5.890 5.270 6.100 5.480 ;
        RECT 0.110 4.630 0.280 4.800 ;
        RECT 7.400 4.900 7.570 5.070 ;
        RECT 1.150 3.580 1.320 3.750 ;
        RECT 0.110 3.240 0.280 3.410 ;
        RECT 2.190 3.540 2.360 3.710 ;
        RECT 5.890 3.520 6.100 3.730 ;
        RECT 0.110 2.880 0.280 3.050 ;
        RECT 7.400 3.150 7.570 3.320 ;
        RECT 1.150 1.830 1.320 2.000 ;
        RECT 0.110 1.490 0.280 1.660 ;
        RECT 2.190 1.790 2.360 1.960 ;
        RECT 5.890 1.770 6.100 1.980 ;
        RECT 0.110 1.130 0.280 1.300 ;
        RECT 7.400 1.400 7.570 1.570 ;
        RECT 1.150 0.080 1.320 0.250 ;
        RECT 0.110 -0.260 0.280 -0.090 ;
        RECT 2.190 0.040 2.360 0.210 ;
        RECT 5.890 0.020 6.100 0.230 ;
        RECT 0.110 -0.620 0.280 -0.450 ;
        RECT 7.400 -0.350 7.570 -0.180 ;
      LAYER met1 ;
        RECT 1.080 5.280 1.400 5.580 ;
        RECT 2.130 5.510 2.440 5.520 ;
        RECT 2.120 5.240 2.440 5.510 ;
        RECT 2.130 5.230 2.420 5.240 ;
        RECT 5.830 5.230 6.180 5.520 ;
        RECT 5.980 5.210 6.180 5.230 ;
        RECT 3.820 4.480 4.100 4.810 ;
        RECT 7.930 4.370 8.340 4.700 ;
        RECT 1.080 3.530 1.400 3.830 ;
        RECT 2.130 3.760 2.440 3.770 ;
        RECT 2.120 3.490 2.440 3.760 ;
        RECT 2.130 3.480 2.420 3.490 ;
        RECT 5.830 3.480 6.180 3.770 ;
        RECT 5.980 3.460 6.180 3.480 ;
        RECT 3.820 2.730 4.100 3.060 ;
        RECT 7.930 2.620 8.340 2.950 ;
        RECT 1.080 1.780 1.400 2.080 ;
        RECT 2.130 2.010 2.440 2.020 ;
        RECT 2.120 1.740 2.440 2.010 ;
        RECT 2.130 1.730 2.420 1.740 ;
        RECT 5.830 1.730 6.180 2.020 ;
        RECT 5.980 1.710 6.180 1.730 ;
        RECT 3.820 0.980 4.100 1.310 ;
        RECT 7.930 0.870 8.340 1.200 ;
        RECT 1.080 0.030 1.400 0.330 ;
        RECT 2.130 0.260 2.440 0.270 ;
        RECT 2.120 -0.010 2.440 0.260 ;
        RECT 2.130 -0.020 2.420 -0.010 ;
        RECT 5.830 -0.020 6.180 0.270 ;
        RECT 5.980 -0.040 6.180 -0.020 ;
        RECT 3.820 -0.770 4.100 -0.440 ;
        RECT 7.930 -0.880 8.340 -0.550 ;
      LAYER via ;
        RECT 1.110 5.290 1.370 5.550 ;
        RECT 2.150 5.250 2.410 5.510 ;
        RECT 5.870 5.240 6.130 5.500 ;
        RECT 3.830 4.520 4.090 4.780 ;
        RECT 7.970 4.400 8.230 4.660 ;
        RECT 1.110 3.540 1.370 3.800 ;
        RECT 2.150 3.500 2.410 3.760 ;
        RECT 5.870 3.490 6.130 3.750 ;
        RECT 3.830 2.770 4.090 3.030 ;
        RECT 7.970 2.650 8.230 2.910 ;
        RECT 1.110 1.790 1.370 2.050 ;
        RECT 2.150 1.750 2.410 2.010 ;
        RECT 5.870 1.740 6.130 2.000 ;
        RECT 3.830 1.020 4.090 1.280 ;
        RECT 7.970 0.900 8.230 1.160 ;
        RECT 1.110 0.040 1.370 0.300 ;
        RECT 2.150 0.000 2.410 0.260 ;
        RECT 5.870 -0.010 6.130 0.250 ;
        RECT 3.830 -0.730 4.090 -0.470 ;
        RECT 7.970 -0.850 8.230 -0.590 ;
      LAYER met2 ;
        RECT 1.080 5.500 1.400 5.550 ;
        RECT 2.110 5.510 2.430 5.520 ;
        RECT 2.110 5.500 2.440 5.510 ;
        RECT -0.230 5.300 2.440 5.500 ;
        RECT 1.080 5.290 1.400 5.300 ;
        RECT 2.110 5.250 2.440 5.300 ;
        RECT 2.110 5.230 2.430 5.250 ;
        RECT 3.790 4.730 4.130 4.790 ;
        RECT 5.870 4.730 6.130 5.530 ;
        RECT 3.790 4.510 6.230 4.730 ;
        RECT 7.940 4.370 8.400 4.690 ;
        RECT 1.080 3.750 1.400 3.800 ;
        RECT 2.110 3.760 2.430 3.770 ;
        RECT 2.110 3.750 2.440 3.760 ;
        RECT -0.230 3.550 2.440 3.750 ;
        RECT 1.080 3.540 1.400 3.550 ;
        RECT 2.110 3.500 2.440 3.550 ;
        RECT 2.110 3.480 2.430 3.500 ;
        RECT 3.790 2.980 4.130 3.040 ;
        RECT 5.870 2.980 6.130 3.780 ;
        RECT 3.790 2.760 6.230 2.980 ;
        RECT 7.940 2.620 8.400 2.940 ;
        RECT 1.080 2.000 1.400 2.050 ;
        RECT 2.110 2.010 2.430 2.020 ;
        RECT 2.110 2.000 2.440 2.010 ;
        RECT -0.230 1.800 2.440 2.000 ;
        RECT 1.080 1.790 1.400 1.800 ;
        RECT 2.110 1.750 2.440 1.800 ;
        RECT 2.110 1.730 2.430 1.750 ;
        RECT 3.790 1.230 4.130 1.290 ;
        RECT 5.870 1.230 6.130 2.030 ;
        RECT 3.790 1.010 6.230 1.230 ;
        RECT 7.940 0.870 8.400 1.190 ;
        RECT 3.790 -0.520 4.130 -0.460 ;
        RECT 5.870 -0.520 6.130 0.280 ;
        RECT 3.790 -0.740 6.230 -0.520 ;
        RECT 7.940 -0.880 8.400 -0.560 ;
  END
END sky130_hilas_LevelShift4InputUp

MACRO sky130_hilas_swc4x2cell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc4x2cell ;
  ORIGIN 10.040 0.260 ;
  SIZE 20.120 BY 6.500 ;
  PIN GATE2
    USE ANALOG ;
    ANTENNADIFFAREA 3.253900 ;
    PORT
      LAYER nwell ;
        RECT 3.760 -0.260 5.990 6.230 ;
      LAYER met1 ;
        RECT 4.410 4.090 4.790 6.240 ;
        RECT 4.400 2.230 4.790 4.090 ;
        RECT 4.410 -0.260 4.790 2.230 ;
    END
  END GATE2
  PIN VTUN
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -1.700 -0.260 1.740 6.230 ;
      LAYER met1 ;
        RECT -0.720 5.870 -0.320 6.240 ;
        RECT 0.360 5.870 0.760 6.240 ;
        RECT -0.720 5.650 0.760 5.870 ;
        RECT -0.720 -0.260 -0.320 5.650 ;
        RECT 0.360 -0.260 0.760 5.650 ;
    END
  END VTUN
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 3.253900 ;
    PORT
      LAYER nwell ;
        RECT -5.950 -0.260 -3.720 6.230 ;
      LAYER met1 ;
        RECT -4.750 4.090 -4.370 6.240 ;
        RECT -4.750 2.230 -4.360 4.090 ;
        RECT -4.750 -0.260 -4.370 2.230 ;
    END
  END GATE1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -10.040 -0.260 -7.480 6.240 ;
        RECT 7.520 -0.260 10.080 6.240 ;
      LAYER met2 ;
        RECT -9.840 5.960 9.900 6.140 ;
        RECT -9.840 5.820 -9.420 5.960 ;
        RECT 9.560 5.830 9.900 5.960 ;
    END
  END VINJ
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 9.560 6.120 9.720 6.230 ;
        RECT 9.560 5.840 9.890 6.120 ;
        RECT 9.560 5.530 9.720 5.840 ;
        RECT 9.450 4.980 9.720 5.530 ;
        RECT 9.450 4.930 9.730 4.980 ;
        RECT 9.560 4.840 9.730 4.930 ;
        RECT 9.560 4.370 9.720 4.840 ;
        RECT 9.560 4.280 9.730 4.370 ;
        RECT 9.450 4.230 9.730 4.280 ;
        RECT 9.450 3.680 9.720 4.230 ;
        RECT 9.560 2.290 9.720 3.680 ;
        RECT 9.450 1.740 9.720 2.290 ;
        RECT 9.450 1.690 9.730 1.740 ;
        RECT 9.560 1.600 9.730 1.690 ;
        RECT 9.560 1.140 9.720 1.600 ;
        RECT 9.560 1.050 9.730 1.140 ;
        RECT 9.450 1.000 9.730 1.050 ;
        RECT 9.450 0.450 9.720 1.000 ;
        RECT 9.560 -0.250 9.720 0.450 ;
      LAYER via ;
        RECT 9.600 5.850 9.860 6.110 ;
    END
    PORT
      LAYER met1 ;
        RECT -9.680 6.110 -9.520 6.230 ;
        RECT -9.830 5.970 -9.520 6.110 ;
        RECT -9.840 5.820 -9.520 5.970 ;
        RECT -9.680 5.530 -9.520 5.820 ;
        RECT -9.680 4.980 -9.410 5.530 ;
        RECT -9.690 4.930 -9.410 4.980 ;
        RECT -9.690 4.840 -9.520 4.930 ;
        RECT -9.680 4.370 -9.520 4.840 ;
        RECT -9.690 4.280 -9.520 4.370 ;
        RECT -9.690 4.230 -9.410 4.280 ;
        RECT -9.680 3.680 -9.410 4.230 ;
        RECT -9.680 2.290 -9.520 3.680 ;
        RECT -9.680 1.740 -9.410 2.290 ;
        RECT -9.690 1.690 -9.410 1.740 ;
        RECT -9.690 1.600 -9.520 1.690 ;
        RECT -9.680 1.140 -9.520 1.600 ;
        RECT -9.690 1.050 -9.520 1.140 ;
        RECT -9.690 1.000 -9.410 1.050 ;
        RECT -9.680 0.450 -9.410 1.000 ;
        RECT -9.680 -0.250 -9.520 0.450 ;
      LAYER via ;
        RECT -9.800 5.840 -9.540 6.100 ;
    END
  END VINJ
  PIN GATESELECT1
    USE ANALOG ;
    ANTENNAGATEAREA 0.720000 ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met1 ;
        RECT -9.270 5.190 -9.080 6.180 ;
        RECT -8.870 5.500 -8.710 6.230 ;
        RECT -8.910 5.480 -8.710 5.500 ;
        RECT -8.920 5.240 -8.690 5.480 ;
        RECT -8.920 5.190 -8.710 5.240 ;
        RECT -9.270 5.070 -9.100 5.190 ;
        RECT -9.270 4.140 -9.110 5.070 ;
        RECT -9.270 4.020 -9.100 4.140 ;
        RECT -8.870 4.020 -8.710 5.190 ;
        RECT -9.270 3.100 -9.080 4.020 ;
        RECT -8.920 3.970 -8.710 4.020 ;
        RECT -8.920 3.730 -8.690 3.970 ;
        RECT -8.910 3.710 -8.710 3.730 ;
        RECT -9.300 3.080 -9.060 3.100 ;
        RECT -8.870 3.080 -8.710 3.710 ;
        RECT -9.300 2.890 -8.710 3.080 ;
        RECT -9.300 2.870 -9.060 2.890 ;
        RECT -9.270 1.950 -9.080 2.870 ;
        RECT -8.870 2.260 -8.710 2.890 ;
        RECT -8.910 2.240 -8.710 2.260 ;
        RECT -8.920 2.000 -8.690 2.240 ;
        RECT -8.920 1.950 -8.710 2.000 ;
        RECT -9.270 1.830 -9.100 1.950 ;
        RECT -9.270 0.910 -9.110 1.830 ;
        RECT -9.270 0.790 -9.100 0.910 ;
        RECT -8.870 0.790 -8.710 1.950 ;
        RECT -9.270 -0.200 -9.080 0.790 ;
        RECT -8.920 0.740 -8.710 0.790 ;
        RECT -8.920 0.500 -8.690 0.740 ;
        RECT -8.910 0.480 -8.710 0.500 ;
        RECT -8.870 -0.250 -8.710 0.480 ;
    END
  END GATESELECT1
  PIN GATESELECT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.720000 ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met1 ;
        RECT 8.750 5.500 8.910 6.230 ;
        RECT 8.750 5.480 8.950 5.500 ;
        RECT 8.730 5.240 8.960 5.480 ;
        RECT 8.750 5.190 8.960 5.240 ;
        RECT 9.120 5.190 9.310 6.180 ;
        RECT 8.750 4.020 8.910 5.190 ;
        RECT 9.140 5.070 9.310 5.190 ;
        RECT 9.150 4.140 9.310 5.070 ;
        RECT 9.140 4.020 9.310 4.140 ;
        RECT 8.750 3.970 8.960 4.020 ;
        RECT 8.730 3.730 8.960 3.970 ;
        RECT 8.750 3.710 8.950 3.730 ;
        RECT 8.750 3.080 8.910 3.710 ;
        RECT 9.120 3.100 9.310 4.020 ;
        RECT 9.100 3.080 9.340 3.100 ;
        RECT 8.750 2.890 9.340 3.080 ;
        RECT 8.750 2.260 8.910 2.890 ;
        RECT 9.100 2.870 9.340 2.890 ;
        RECT 8.750 2.240 8.950 2.260 ;
        RECT 8.730 2.000 8.960 2.240 ;
        RECT 8.750 1.950 8.960 2.000 ;
        RECT 9.120 1.950 9.310 2.870 ;
        RECT 8.750 0.790 8.910 1.950 ;
        RECT 9.140 1.830 9.310 1.950 ;
        RECT 9.150 0.910 9.310 1.830 ;
        RECT 9.140 0.790 9.310 0.910 ;
        RECT 8.750 0.740 8.960 0.790 ;
        RECT 8.730 0.500 8.960 0.740 ;
        RECT 8.750 0.480 8.950 0.500 ;
        RECT 8.750 -0.250 8.910 0.480 ;
        RECT 9.120 -0.200 9.310 0.790 ;
    END
  END GATESELECT2
  PIN ROW1
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT -7.880 5.250 -7.570 5.270 ;
        RECT 7.610 5.250 7.920 5.270 ;
        RECT -10.040 5.240 -7.480 5.250 ;
        RECT 7.520 5.240 10.080 5.250 ;
        RECT -10.040 5.070 10.080 5.240 ;
        RECT -7.880 5.060 7.920 5.070 ;
        RECT -7.880 4.940 -7.570 5.060 ;
        RECT 7.610 4.940 7.920 5.060 ;
    END
  END ROW1
  PIN ROW2
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT -7.880 4.140 -7.570 4.270 ;
        RECT 7.610 4.140 7.920 4.270 ;
        RECT -10.040 3.960 10.080 4.140 ;
        RECT -7.880 3.940 -7.570 3.960 ;
        RECT 7.610 3.940 7.920 3.960 ;
    END
  END ROW2
  PIN DRAIN1
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT -7.880 5.680 -7.570 5.820 ;
        RECT 7.610 5.680 7.920 5.820 ;
        RECT -10.040 5.500 10.080 5.680 ;
        RECT -7.880 5.490 -7.570 5.500 ;
        RECT 7.610 5.490 7.920 5.500 ;
    END
  END DRAIN1
  PIN DRAIN2
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT -7.880 3.710 -7.570 3.720 ;
        RECT 7.610 3.710 7.920 3.720 ;
        RECT -10.040 3.530 10.080 3.710 ;
        RECT -7.880 3.390 -7.570 3.530 ;
        RECT 7.610 3.390 7.920 3.530 ;
    END
  END DRAIN2
  PIN DRAIN3
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT -7.880 2.440 -7.570 2.580 ;
        RECT 7.610 2.440 7.920 2.580 ;
        RECT -10.040 2.260 10.080 2.440 ;
        RECT -7.880 2.250 -7.570 2.260 ;
        RECT 7.610 2.250 7.920 2.260 ;
    END
  END DRAIN3
  PIN ROW3
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT -7.880 2.010 -7.570 2.030 ;
        RECT 7.610 2.010 7.920 2.030 ;
        RECT -10.040 1.830 10.080 2.010 ;
        RECT -7.880 1.700 -7.570 1.830 ;
        RECT 7.610 1.700 7.920 1.830 ;
    END
  END ROW3
  PIN ROW4
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT -7.880 0.910 -7.570 1.040 ;
        RECT 7.610 0.910 7.920 1.040 ;
        RECT -10.040 0.730 10.080 0.910 ;
        RECT -7.880 0.710 -7.570 0.730 ;
        RECT 7.610 0.710 7.920 0.730 ;
    END
  END ROW4
  PIN DRAIN4
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT -7.880 0.480 -7.570 0.490 ;
        RECT 7.610 0.480 7.920 0.490 ;
        RECT -10.040 0.310 10.080 0.480 ;
        RECT -10.040 0.300 -7.570 0.310 ;
        RECT -7.880 0.160 -7.570 0.300 ;
        RECT 7.610 0.300 10.080 0.310 ;
        RECT 7.610 0.160 7.920 0.300 ;
    END
  END DRAIN4
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT -6.970 1.520 -6.650 1.580 ;
        RECT -3.040 1.520 -2.720 1.530 ;
        RECT 2.760 1.520 3.080 1.530 ;
        RECT 6.690 1.520 7.010 1.580 ;
        RECT -6.970 1.340 7.010 1.520 ;
        RECT -6.970 1.290 -6.650 1.340 ;
        RECT -3.040 1.270 -2.720 1.340 ;
        RECT 2.760 1.270 3.080 1.340 ;
        RECT 6.690 1.290 7.010 1.340 ;
    END
    PORT
      LAYER met1 ;
        RECT -6.930 4.850 -6.690 6.240 ;
        RECT -6.940 4.190 -6.670 4.850 ;
        RECT -6.930 1.600 -6.690 4.190 ;
        RECT -6.940 1.280 -6.680 1.600 ;
        RECT -6.930 -0.260 -6.690 1.280 ;
      LAYER via ;
        RECT -6.940 1.310 -6.680 1.570 ;
    END
    PORT
      LAYER met1 ;
        RECT -3.000 4.830 -2.760 6.240 ;
        RECT -3.010 4.170 -2.750 4.830 ;
        RECT -3.000 1.560 -2.760 4.170 ;
        RECT -3.010 1.240 -2.750 1.560 ;
        RECT -3.000 -0.260 -2.760 1.240 ;
      LAYER via ;
        RECT -3.010 1.270 -2.750 1.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.800 4.830 3.040 6.240 ;
        RECT 2.790 4.170 3.050 4.830 ;
        RECT 2.800 1.560 3.040 4.170 ;
        RECT 2.790 1.240 3.050 1.560 ;
        RECT 2.800 -0.260 3.040 1.240 ;
      LAYER via ;
        RECT 2.790 1.270 3.050 1.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.730 4.850 6.970 6.240 ;
        RECT 6.710 4.190 6.980 4.850 ;
        RECT 6.730 1.600 6.970 4.190 ;
        RECT 6.720 1.280 6.980 1.600 ;
        RECT 6.730 -0.260 6.970 1.280 ;
      LAYER via ;
        RECT 6.720 1.310 6.980 1.570 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT -9.640 5.500 -9.440 5.850 ;
        RECT -7.900 5.770 -7.580 5.780 ;
        RECT -8.160 5.600 -7.580 5.770 ;
        RECT -7.910 5.550 -7.580 5.600 ;
        RECT -7.900 5.520 -7.580 5.550 ;
        RECT 7.620 5.770 7.940 5.780 ;
        RECT 7.620 5.600 8.200 5.770 ;
        RECT 7.620 5.550 7.950 5.600 ;
        RECT 7.620 5.520 7.940 5.550 ;
        RECT -9.650 5.470 -9.440 5.500 ;
        RECT 9.480 5.500 9.680 5.850 ;
        RECT -9.650 4.880 -9.430 5.470 ;
        RECT -8.910 4.880 -8.710 5.480 ;
        RECT -7.900 5.190 -7.580 5.230 ;
        RECT -7.910 5.150 -7.580 5.190 ;
        RECT -8.160 4.980 -7.580 5.150 ;
        RECT -7.900 4.970 -7.580 4.980 ;
        RECT 7.620 5.190 7.940 5.230 ;
        RECT 7.620 5.150 7.950 5.190 ;
        RECT 7.620 4.980 8.200 5.150 ;
        RECT 7.620 4.970 7.940 4.980 ;
        RECT 8.750 4.880 8.950 5.480 ;
        RECT 9.480 5.470 9.690 5.500 ;
        RECT 9.470 4.880 9.690 5.470 ;
        RECT -9.650 3.740 -9.430 4.330 ;
        RECT -9.650 3.710 -9.440 3.740 ;
        RECT -8.910 3.730 -8.710 4.330 ;
        RECT -6.900 4.250 -6.730 4.780 ;
        RECT -2.960 4.260 -2.790 4.790 ;
        RECT 2.830 4.260 3.000 4.790 ;
        RECT 6.770 4.250 6.940 4.780 ;
        RECT -7.900 4.230 -7.580 4.240 ;
        RECT -8.160 4.060 -7.580 4.230 ;
        RECT -7.910 4.020 -7.580 4.060 ;
        RECT -7.900 3.980 -7.580 4.020 ;
        RECT 7.620 4.230 7.940 4.240 ;
        RECT 7.620 4.060 8.200 4.230 ;
        RECT 7.620 4.020 7.950 4.060 ;
        RECT 7.620 3.980 7.940 4.020 ;
        RECT 8.750 3.730 8.950 4.330 ;
        RECT 9.470 3.740 9.690 4.330 ;
        RECT -9.640 3.360 -9.440 3.710 ;
        RECT 9.480 3.710 9.690 3.740 ;
        RECT -7.900 3.660 -7.580 3.690 ;
        RECT -7.910 3.610 -7.580 3.660 ;
        RECT -8.160 3.440 -7.580 3.610 ;
        RECT 7.620 3.660 7.940 3.690 ;
        RECT 7.620 3.610 7.950 3.660 ;
        RECT -7.900 3.430 -7.580 3.440 ;
        RECT -9.270 2.900 -8.830 3.070 ;
        RECT -9.640 2.260 -9.440 2.610 ;
        RECT -7.900 2.530 -7.580 2.540 ;
        RECT -8.160 2.360 -7.580 2.530 ;
        RECT -6.900 2.410 -6.730 3.420 ;
        RECT -4.970 2.690 -4.420 3.120 ;
        RECT -2.970 2.550 -2.800 3.560 ;
        RECT -0.940 2.760 -0.390 3.190 ;
        RECT 0.430 2.760 0.980 3.190 ;
        RECT 2.840 2.550 3.010 3.560 ;
        RECT 7.620 3.440 8.200 3.610 ;
        RECT 7.620 3.430 7.940 3.440 ;
        RECT 4.460 2.690 5.010 3.120 ;
        RECT 6.770 2.410 6.940 3.420 ;
        RECT 9.480 3.360 9.680 3.710 ;
        RECT 8.870 2.900 9.310 3.070 ;
        RECT 7.620 2.530 7.940 2.540 ;
        RECT -7.910 2.310 -7.580 2.360 ;
        RECT -7.900 2.280 -7.580 2.310 ;
        RECT 7.620 2.360 8.200 2.530 ;
        RECT 7.620 2.310 7.950 2.360 ;
        RECT 7.620 2.280 7.940 2.310 ;
        RECT -9.650 2.230 -9.440 2.260 ;
        RECT 9.480 2.260 9.680 2.610 ;
        RECT -9.650 1.640 -9.430 2.230 ;
        RECT -8.910 1.640 -8.710 2.240 ;
        RECT -7.900 1.950 -7.580 1.990 ;
        RECT -7.910 1.910 -7.580 1.950 ;
        RECT -8.160 1.740 -7.580 1.910 ;
        RECT -7.900 1.730 -7.580 1.740 ;
        RECT 7.620 1.950 7.940 1.990 ;
        RECT 7.620 1.910 7.950 1.950 ;
        RECT 7.620 1.740 8.200 1.910 ;
        RECT 7.620 1.730 7.940 1.740 ;
        RECT 8.750 1.640 8.950 2.240 ;
        RECT 9.480 2.230 9.690 2.260 ;
        RECT 9.470 1.640 9.690 2.230 ;
        RECT -9.650 0.510 -9.430 1.100 ;
        RECT -9.650 0.480 -9.440 0.510 ;
        RECT -8.910 0.500 -8.710 1.100 ;
        RECT -7.900 1.000 -7.580 1.010 ;
        RECT -8.160 0.830 -7.580 1.000 ;
        RECT -7.910 0.790 -7.580 0.830 ;
        RECT -7.900 0.750 -7.580 0.790 ;
        RECT 7.620 1.000 7.940 1.010 ;
        RECT 7.620 0.830 8.200 1.000 ;
        RECT 7.620 0.790 7.950 0.830 ;
        RECT 7.620 0.750 7.940 0.790 ;
        RECT 8.750 0.500 8.950 1.100 ;
        RECT 9.470 0.510 9.690 1.100 ;
        RECT -9.640 0.130 -9.440 0.480 ;
        RECT 9.480 0.480 9.690 0.510 ;
        RECT -7.900 0.430 -7.580 0.460 ;
        RECT -7.910 0.380 -7.580 0.430 ;
        RECT -8.160 0.210 -7.580 0.380 ;
        RECT -7.900 0.200 -7.580 0.210 ;
        RECT 7.620 0.430 7.940 0.460 ;
        RECT 7.620 0.380 7.950 0.430 ;
        RECT 7.620 0.210 8.200 0.380 ;
        RECT 7.620 0.200 7.940 0.210 ;
        RECT 9.480 0.130 9.680 0.480 ;
      LAYER mcon ;
        RECT -7.810 5.560 -7.640 5.730 ;
        RECT 7.680 5.560 7.850 5.730 ;
        RECT -9.620 5.300 -9.450 5.470 ;
        RECT -8.890 5.270 -8.720 5.440 ;
        RECT 8.760 5.270 8.930 5.440 ;
        RECT -7.810 5.010 -7.640 5.180 ;
        RECT 7.680 5.010 7.850 5.180 ;
        RECT 9.490 5.300 9.660 5.470 ;
        RECT -6.900 4.610 -6.730 4.780 ;
        RECT -9.620 3.740 -9.450 3.910 ;
        RECT -2.960 4.620 -2.790 4.790 ;
        RECT 2.830 4.620 3.000 4.790 ;
        RECT 6.770 4.610 6.940 4.780 ;
        RECT -7.810 4.030 -7.640 4.200 ;
        RECT 7.680 4.030 7.850 4.200 ;
        RECT -8.890 3.770 -8.720 3.940 ;
        RECT 8.760 3.770 8.930 3.940 ;
        RECT 9.490 3.740 9.660 3.910 ;
        RECT -7.810 3.480 -7.640 3.650 ;
        RECT -6.900 3.020 -6.730 3.190 ;
        RECT -2.970 3.160 -2.800 3.330 ;
        RECT 7.680 3.480 7.850 3.650 ;
        RECT -6.900 2.660 -6.730 2.830 ;
        RECT -4.690 2.770 -4.420 3.040 ;
        RECT -2.970 2.800 -2.800 2.970 ;
        RECT -7.810 2.320 -7.640 2.490 ;
        RECT -0.660 2.840 -0.390 3.110 ;
        RECT 0.430 2.840 0.700 3.110 ;
        RECT 2.840 3.160 3.010 3.330 ;
        RECT 2.840 2.800 3.010 2.970 ;
        RECT 4.460 2.770 4.730 3.040 ;
        RECT 6.770 3.020 6.940 3.190 ;
        RECT 9.130 2.900 9.310 3.070 ;
        RECT 6.770 2.660 6.940 2.830 ;
        RECT 7.680 2.320 7.850 2.490 ;
        RECT -9.620 2.060 -9.450 2.230 ;
        RECT -8.890 2.030 -8.720 2.200 ;
        RECT 8.760 2.030 8.930 2.200 ;
        RECT -7.810 1.770 -7.640 1.940 ;
        RECT 7.680 1.770 7.850 1.940 ;
        RECT 9.490 2.060 9.660 2.230 ;
        RECT -9.620 0.510 -9.450 0.680 ;
        RECT -7.810 0.800 -7.640 0.970 ;
        RECT 7.680 0.800 7.850 0.970 ;
        RECT -8.890 0.540 -8.720 0.710 ;
        RECT 8.760 0.540 8.930 0.710 ;
        RECT 9.490 0.510 9.660 0.680 ;
        RECT -7.810 0.250 -7.640 0.420 ;
        RECT 7.680 0.250 7.850 0.420 ;
      LAYER met1 ;
        RECT -7.890 5.490 -7.570 5.810 ;
        RECT 7.610 5.490 7.930 5.810 ;
        RECT -7.890 4.940 -7.570 5.260 ;
        RECT 7.610 4.940 7.930 5.260 ;
        RECT -7.890 3.950 -7.570 4.270 ;
        RECT 7.610 3.950 7.930 4.270 ;
        RECT -7.890 3.400 -7.570 3.720 ;
        RECT 7.610 3.400 7.930 3.720 ;
        RECT -7.890 2.250 -7.570 2.570 ;
        RECT 7.610 2.250 7.930 2.570 ;
        RECT -7.890 1.700 -7.570 2.020 ;
        RECT 7.610 1.700 7.930 2.020 ;
        RECT -7.890 0.720 -7.570 1.040 ;
        RECT 7.610 0.720 7.930 1.040 ;
        RECT -7.890 0.170 -7.570 0.490 ;
        RECT 7.610 0.170 7.930 0.490 ;
      LAYER via ;
        RECT -7.860 5.520 -7.600 5.780 ;
        RECT 7.640 5.520 7.900 5.780 ;
        RECT -7.860 4.970 -7.600 5.230 ;
        RECT 7.640 4.970 7.900 5.230 ;
        RECT -7.860 3.980 -7.600 4.240 ;
        RECT 7.640 3.980 7.900 4.240 ;
        RECT -7.860 3.430 -7.600 3.690 ;
        RECT 7.640 3.430 7.900 3.690 ;
        RECT -7.860 2.280 -7.600 2.540 ;
        RECT 7.640 2.280 7.900 2.540 ;
        RECT -7.860 1.730 -7.600 1.990 ;
        RECT 7.640 1.730 7.900 1.990 ;
        RECT -7.860 0.750 -7.600 1.010 ;
        RECT 7.640 0.750 7.900 1.010 ;
        RECT -7.860 0.200 -7.600 0.460 ;
        RECT 7.640 0.200 7.900 0.460 ;
  END
END sky130_hilas_swc4x2cell

MACRO sky130_hilas_Trans4small
  CLASS BLOCK ;
  FOREIGN sky130_hilas_Trans4small ;
  ORIGIN -1.910 1.500 ;
  SIZE 2.800 BY 6.050 ;
  PIN NFET_SOURCE1
    USE ANALOG ;
    ANTENNADIFFAREA 0.130200 ;
    PORT
      LAYER met2 ;
        RECT 2.500 4.250 2.810 4.340 ;
        RECT 1.910 4.080 2.810 4.250 ;
        RECT 1.910 3.980 2.050 4.080 ;
        RECT 2.500 4.010 2.810 4.080 ;
    END
  END NFET_SOURCE1
  PIN NFET_GATE1
    USE ANALOG ;
    ANTENNAGATEAREA 0.113400 ;
    PORT
      LAYER met2 ;
        RECT 2.070 3.740 2.380 3.840 ;
        RECT 1.910 3.570 2.380 3.740 ;
        RECT 2.070 3.510 2.380 3.570 ;
    END
  END NFET_GATE1
  PIN NFET_SOURCE2
    USE ANALOG ;
    ANTENNADIFFAREA 0.130200 ;
    PORT
      LAYER met2 ;
        RECT 2.510 3.260 2.820 3.350 ;
        RECT 1.980 3.230 2.820 3.260 ;
        RECT 1.910 3.090 2.820 3.230 ;
        RECT 1.910 3.060 2.050 3.090 ;
        RECT 2.510 3.020 2.820 3.090 ;
    END
  END NFET_SOURCE2
  PIN NFET_GATE2
    USE ANALOG ;
    ANTENNAGATEAREA 0.113400 ;
    PORT
      LAYER met2 ;
        RECT 2.050 2.820 2.360 2.920 ;
        RECT 1.910 2.650 2.360 2.820 ;
        RECT 2.050 2.590 2.360 2.650 ;
    END
  END NFET_GATE2
  PIN NFET_SOURCE3
    USE ANALOG ;
    ANTENNADIFFAREA 0.130200 ;
    PORT
      LAYER met2 ;
        RECT 1.910 2.280 2.050 2.310 ;
        RECT 1.910 2.270 2.120 2.280 ;
        RECT 2.510 2.270 2.820 2.360 ;
        RECT 1.910 2.140 2.820 2.270 ;
        RECT 1.980 2.100 2.820 2.140 ;
        RECT 2.510 2.030 2.820 2.100 ;
    END
  END NFET_SOURCE3
  PIN NFET_GATE3
    USE ANALOG ;
    ANTENNAGATEAREA 0.113400 ;
    PORT
      LAYER met2 ;
        RECT 2.030 1.900 2.340 1.930 ;
        RECT 1.910 1.730 2.340 1.900 ;
        RECT 2.030 1.600 2.340 1.730 ;
    END
  END NFET_GATE3
  PIN PFET_SOURCE1
    USE ANALOG ;
    ANTENNADIFFAREA 0.117600 ;
    PORT
      LAYER met2 ;
        RECT 2.320 1.320 2.630 1.430 ;
        RECT 1.980 1.310 2.630 1.320 ;
        RECT 1.910 1.130 2.630 1.310 ;
        RECT 1.910 1.120 2.050 1.130 ;
        RECT 2.320 1.100 2.630 1.130 ;
    END
  END PFET_SOURCE1
  PIN PFET_GATE1
    USE ANALOG ;
    ANTENNAGATEAREA 0.163800 ;
    PORT
      LAYER met2 ;
        RECT 2.290 0.900 2.610 0.960 ;
        RECT 1.980 0.890 2.610 0.900 ;
        RECT 1.910 0.710 2.610 0.890 ;
        RECT 1.910 0.700 2.050 0.710 ;
        RECT 2.290 0.640 2.610 0.710 ;
    END
  END PFET_GATE1
  PIN PFET_SOURCE2
    USE ANALOG ;
    ANTENNADIFFAREA 0.117600 ;
    PORT
      LAYER met2 ;
        RECT 1.910 0.330 2.050 0.350 ;
        RECT 2.320 0.330 2.630 0.440 ;
        RECT 1.910 0.160 2.630 0.330 ;
        RECT 1.980 0.140 2.630 0.160 ;
        RECT 2.320 0.110 2.630 0.140 ;
    END
  END PFET_SOURCE2
  PIN PFET_GATE2
    USE ANALOG ;
    ANTENNAGATEAREA 0.163800 ;
    PORT
      LAYER met2 ;
        RECT 1.910 -0.090 2.050 -0.070 ;
        RECT 2.290 -0.090 2.610 -0.030 ;
        RECT 1.910 -0.260 2.610 -0.090 ;
        RECT 1.980 -0.280 2.610 -0.260 ;
        RECT 2.290 -0.350 2.610 -0.280 ;
    END
  END PFET_GATE2
  PIN PFET_SOURCE3
    USE ANALOG ;
    ANTENNADIFFAREA 0.117600 ;
    PORT
      LAYER met2 ;
        RECT 1.910 -0.660 2.050 -0.610 ;
        RECT 2.320 -0.660 2.630 -0.550 ;
        RECT 1.910 -0.800 2.630 -0.660 ;
        RECT 1.980 -0.850 2.630 -0.800 ;
        RECT 2.320 -0.880 2.630 -0.850 ;
    END
  END PFET_SOURCE3
  PIN PFET_GATE3
    USE ANALOG ;
    ANTENNAGATEAREA 0.163800 ;
    PORT
      LAYER met2 ;
        RECT 1.910 -1.050 2.050 -1.030 ;
        RECT 1.910 -1.080 2.060 -1.050 ;
        RECT 2.290 -1.080 2.610 -1.020 ;
        RECT 1.910 -1.220 2.610 -1.080 ;
        RECT 1.980 -1.270 2.610 -1.220 ;
        RECT 2.290 -1.340 2.610 -1.270 ;
    END
  END PFET_GATE3
  PIN WELL
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 1.980 1.590 4.010 1.600 ;
        RECT 1.980 -1.500 4.550 1.590 ;
      LAYER met1 ;
        RECT 4.090 -0.200 4.310 4.380 ;
        RECT 4.040 -0.430 4.330 -0.200 ;
        RECT 4.090 -1.500 4.310 -0.430 ;
    END
  END WELL
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 4.490 3.750 4.710 4.380 ;
        RECT 4.480 3.460 4.710 3.750 ;
        RECT 4.490 -1.500 4.710 3.460 ;
    END
  END VGND
  PIN PFET_DRAIN3
    USE ANALOG ;
    ANTENNADIFFAREA 0.113400 ;
    PORT
      LAYER met2 ;
        RECT 3.620 -0.670 3.930 -0.650 ;
        RECT 3.620 -0.870 4.710 -0.670 ;
        RECT 3.620 -0.980 3.930 -0.870 ;
    END
  END PFET_DRAIN3
  PIN PFET_DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.113400 ;
    PORT
      LAYER met2 ;
        RECT 3.620 0.290 3.930 0.340 ;
        RECT 3.620 0.090 4.710 0.290 ;
        RECT 3.620 0.010 3.930 0.090 ;
    END
  END PFET_DRAIN2
  PIN PFET_DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.113400 ;
    PORT
      LAYER met2 ;
        RECT 3.620 1.250 3.930 1.330 ;
        RECT 3.620 1.050 4.710 1.250 ;
        RECT 3.620 1.000 3.930 1.050 ;
    END
  END PFET_DRAIN1
  PIN NFET_DRAIN3
    USE ANALOG ;
    ANTENNADIFFAREA 0.130200 ;
    PORT
      LAYER met2 ;
        RECT 3.600 2.320 3.910 2.370 ;
        RECT 3.600 2.150 4.710 2.320 ;
        RECT 3.600 2.110 4.060 2.150 ;
        RECT 3.600 2.040 3.910 2.110 ;
    END
  END NFET_DRAIN3
  PIN NFET_DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.130200 ;
    PORT
      LAYER met2 ;
        RECT 3.600 3.270 3.910 3.360 ;
        RECT 3.600 3.240 4.060 3.270 ;
        RECT 3.600 3.070 4.710 3.240 ;
        RECT 3.600 3.030 3.910 3.070 ;
    END
  END NFET_DRAIN2
  PIN NFET_DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.130200 ;
    PORT
      LAYER met2 ;
        RECT 3.590 4.260 3.900 4.350 ;
        RECT 3.590 4.160 4.050 4.260 ;
        RECT 3.590 4.020 4.710 4.160 ;
        RECT 3.890 3.990 4.710 4.020 ;
    END
  END NFET_DRAIN1
  OBS
      LAYER li1 ;
        RECT 2.820 4.300 3.020 4.340 ;
        RECT 2.510 4.040 3.020 4.300 ;
        RECT 2.820 4.010 3.020 4.040 ;
        RECT 3.410 4.310 3.610 4.340 ;
        RECT 3.410 4.270 3.920 4.310 ;
        RECT 3.410 4.080 3.930 4.270 ;
        RECT 3.410 4.050 3.920 4.080 ;
        RECT 3.410 4.010 3.610 4.050 ;
        RECT 2.240 3.800 2.600 3.870 ;
        RECT 2.080 3.700 2.600 3.800 ;
        RECT 4.110 3.760 4.280 3.810 ;
        RECT 4.100 3.730 4.280 3.760 ;
        RECT 4.100 3.720 4.530 3.730 ;
        RECT 2.080 3.620 2.450 3.700 ;
        RECT 2.080 3.570 2.410 3.620 ;
        RECT 2.080 3.540 2.400 3.570 ;
        RECT 4.100 3.490 4.690 3.720 ;
        RECT 4.100 3.480 4.530 3.490 ;
        RECT 4.100 3.450 4.290 3.480 ;
        RECT 4.110 3.420 4.290 3.450 ;
        RECT 2.830 3.310 3.030 3.350 ;
        RECT 2.520 3.050 3.030 3.310 ;
        RECT 2.830 3.020 3.030 3.050 ;
        RECT 3.420 3.320 3.620 3.350 ;
        RECT 3.420 3.280 3.930 3.320 ;
        RECT 3.420 3.090 3.940 3.280 ;
        RECT 3.420 3.060 3.930 3.090 ;
        RECT 3.420 3.020 3.620 3.060 ;
        RECT 2.060 2.710 2.610 2.880 ;
        RECT 2.060 2.650 2.390 2.710 ;
        RECT 2.060 2.620 2.380 2.650 ;
        RECT 2.830 2.320 3.030 2.360 ;
        RECT 2.520 2.060 3.030 2.320 ;
        RECT 2.830 2.030 3.030 2.060 ;
        RECT 3.420 2.330 3.620 2.360 ;
        RECT 3.420 2.290 3.930 2.330 ;
        RECT 3.420 2.100 3.940 2.290 ;
        RECT 3.420 2.070 3.930 2.100 ;
        RECT 3.420 2.030 3.620 2.070 ;
        RECT 2.040 1.720 2.610 1.890 ;
        RECT 2.040 1.660 2.370 1.720 ;
        RECT 2.040 1.630 2.360 1.660 ;
        RECT 2.330 1.350 2.650 1.390 ;
        RECT 2.330 1.330 2.660 1.350 ;
        RECT 2.330 1.130 2.950 1.330 ;
        RECT 2.780 1.000 2.950 1.130 ;
        RECT 3.460 1.290 3.630 1.330 ;
        RECT 3.460 1.250 3.950 1.290 ;
        RECT 3.460 1.060 3.960 1.250 ;
        RECT 3.460 1.030 3.950 1.060 ;
        RECT 3.460 1.000 3.630 1.030 ;
        RECT 2.140 0.890 2.570 0.910 ;
        RECT 2.120 0.720 2.570 0.890 ;
        RECT 2.140 0.700 2.570 0.720 ;
        RECT 2.330 0.360 2.650 0.400 ;
        RECT 2.330 0.340 2.660 0.360 ;
        RECT 2.330 0.140 2.950 0.340 ;
        RECT 2.780 0.010 2.950 0.140 ;
        RECT 3.460 0.300 3.630 0.340 ;
        RECT 3.460 0.260 3.950 0.300 ;
        RECT 3.460 0.070 3.960 0.260 ;
        RECT 3.460 0.040 3.950 0.070 ;
        RECT 3.460 0.010 3.630 0.040 ;
        RECT 2.140 -0.100 2.570 -0.080 ;
        RECT 2.120 -0.270 2.570 -0.100 ;
        RECT 4.070 -0.230 4.300 -0.220 ;
        RECT 2.140 -0.290 2.570 -0.270 ;
        RECT 3.990 -0.400 4.320 -0.230 ;
        RECT 4.070 -0.410 4.300 -0.400 ;
        RECT 2.330 -0.630 2.650 -0.590 ;
        RECT 2.330 -0.650 2.660 -0.630 ;
        RECT 2.330 -0.850 2.950 -0.650 ;
        RECT 2.780 -0.980 2.950 -0.850 ;
        RECT 3.460 -0.690 3.630 -0.650 ;
        RECT 3.460 -0.730 3.950 -0.690 ;
        RECT 3.460 -0.920 3.960 -0.730 ;
        RECT 3.460 -0.950 3.950 -0.920 ;
        RECT 3.460 -0.980 3.630 -0.950 ;
        RECT 2.140 -1.090 2.570 -1.070 ;
        RECT 2.120 -1.260 2.570 -1.090 ;
        RECT 2.140 -1.280 2.570 -1.260 ;
      LAYER mcon ;
        RECT 2.570 4.080 2.740 4.250 ;
        RECT 3.660 4.090 3.830 4.260 ;
        RECT 2.140 3.580 2.310 3.750 ;
        RECT 4.510 3.520 4.680 3.690 ;
        RECT 2.580 3.090 2.750 3.260 ;
        RECT 3.670 3.100 3.840 3.270 ;
        RECT 2.120 2.660 2.290 2.830 ;
        RECT 2.580 2.100 2.750 2.270 ;
        RECT 3.670 2.110 3.840 2.280 ;
        RECT 2.100 1.670 2.270 1.840 ;
        RECT 2.390 1.170 2.560 1.340 ;
        RECT 3.690 1.070 3.860 1.240 ;
        RECT 2.390 0.180 2.560 0.350 ;
        RECT 3.690 0.080 3.860 0.250 ;
        RECT 4.100 -0.400 4.270 -0.230 ;
        RECT 2.390 -0.810 2.560 -0.640 ;
        RECT 3.690 -0.910 3.860 -0.740 ;
      LAYER met1 ;
        RECT 2.500 4.010 2.820 4.330 ;
        RECT 3.590 4.020 3.910 4.340 ;
        RECT 2.070 3.510 2.390 3.830 ;
        RECT 2.510 3.020 2.830 3.340 ;
        RECT 3.600 3.030 3.920 3.350 ;
        RECT 2.050 2.590 2.370 2.910 ;
        RECT 2.510 2.030 2.830 2.350 ;
        RECT 3.600 2.040 3.920 2.360 ;
        RECT 2.030 1.600 2.350 1.920 ;
        RECT 2.320 1.100 2.640 1.420 ;
        RECT 3.620 1.000 3.940 1.320 ;
        RECT 2.290 0.920 2.610 0.960 ;
        RECT 2.060 0.690 2.610 0.920 ;
        RECT 2.290 0.640 2.610 0.690 ;
        RECT 2.320 0.110 2.640 0.430 ;
        RECT 3.620 0.010 3.940 0.330 ;
        RECT 2.290 -0.070 2.610 -0.030 ;
        RECT 2.060 -0.300 2.610 -0.070 ;
        RECT 2.290 -0.350 2.610 -0.300 ;
        RECT 2.320 -0.880 2.640 -0.560 ;
        RECT 3.620 -0.980 3.940 -0.660 ;
        RECT 2.290 -1.060 2.610 -1.020 ;
        RECT 2.060 -1.290 2.610 -1.060 ;
        RECT 2.290 -1.340 2.610 -1.290 ;
      LAYER via ;
        RECT 2.530 4.040 2.790 4.300 ;
        RECT 3.620 4.050 3.880 4.310 ;
        RECT 2.100 3.540 2.360 3.800 ;
        RECT 2.540 3.050 2.800 3.310 ;
        RECT 3.630 3.060 3.890 3.320 ;
        RECT 2.080 2.620 2.340 2.880 ;
        RECT 2.540 2.060 2.800 2.320 ;
        RECT 3.630 2.070 3.890 2.330 ;
        RECT 2.060 1.630 2.320 1.890 ;
        RECT 2.350 1.130 2.610 1.390 ;
        RECT 3.650 1.030 3.910 1.290 ;
        RECT 2.320 0.670 2.580 0.930 ;
        RECT 2.350 0.140 2.610 0.400 ;
        RECT 3.650 0.040 3.910 0.300 ;
        RECT 2.320 -0.320 2.580 -0.060 ;
        RECT 2.350 -0.850 2.610 -0.590 ;
        RECT 3.650 -0.950 3.910 -0.690 ;
        RECT 2.320 -1.310 2.580 -1.050 ;
  END
END sky130_hilas_Trans4small

MACRO sky130_hilas_drainSelect01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_drainSelect01 ;
  ORIGIN -10.500 0.280 ;
  SIZE 5.720 BY 6.590 ;
  PIN DRAIN3
    ANTENNADIFFAREA 0.322600 ;
    PORT
      LAYER met2 ;
        RECT 12.250 2.680 12.570 2.700 ;
        RECT 14.660 2.680 14.980 2.730 ;
        RECT 10.500 2.580 11.070 2.590 ;
        RECT 10.500 2.570 11.770 2.580 ;
        RECT 12.250 2.570 14.980 2.680 ;
        RECT 10.500 2.490 14.980 2.570 ;
        RECT 10.500 2.440 12.570 2.490 ;
        RECT 10.500 2.410 12.500 2.440 ;
        RECT 14.660 2.410 14.980 2.490 ;
    END
  END DRAIN3
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 10.500 -0.280 13.920 6.310 ;
      LAYER met1 ;
        RECT 11.080 6.040 11.330 6.260 ;
        RECT 10.690 4.970 11.330 6.040 ;
        RECT 11.080 4.260 11.330 4.970 ;
        RECT 10.690 3.190 11.330 4.260 ;
        RECT 11.080 2.840 11.330 3.190 ;
        RECT 10.690 1.770 11.330 2.840 ;
        RECT 11.080 1.060 11.330 1.770 ;
        RECT 10.690 -0.010 11.330 1.060 ;
        RECT 11.080 -0.230 11.330 -0.010 ;
    END
  END VINJ
  PIN DRAIN_MUX
    USE ANALOG ;
    ANTENNADIFFAREA 0.846400 ;
    PORT
      LAYER met1 ;
        RECT 14.070 -0.230 14.300 6.260 ;
    END
  END DRAIN_MUX
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 15.420 6.040 15.610 6.260 ;
        RECT 15.420 5.550 15.890 6.040 ;
        RECT 15.420 5.290 15.610 5.550 ;
        RECT 15.380 5.000 15.610 5.290 ;
        RECT 15.420 4.230 15.610 5.000 ;
        RECT 15.380 3.940 15.610 4.230 ;
        RECT 15.420 3.680 15.610 3.940 ;
        RECT 15.420 3.190 15.890 3.680 ;
        RECT 15.420 2.840 15.610 3.190 ;
        RECT 15.420 2.350 15.890 2.840 ;
        RECT 15.420 2.090 15.610 2.350 ;
        RECT 15.380 1.800 15.610 2.090 ;
        RECT 15.420 1.030 15.610 1.800 ;
        RECT 15.380 0.740 15.610 1.030 ;
        RECT 15.420 0.480 15.610 0.740 ;
        RECT 15.420 -0.010 15.890 0.480 ;
        RECT 15.420 -0.230 15.610 -0.010 ;
    END
  END VGND
  PIN SELECT2
    ANTENNAGATEAREA 0.730000 ;
    PORT
      LAYER met2 ;
        RECT 15.740 4.070 16.080 4.130 ;
        RECT 15.740 3.830 16.220 4.070 ;
    END
  END SELECT2
  PIN SELECT1
    ANTENNAGATEAREA 0.730000 ;
    PORT
      LAYER met2 ;
        RECT 15.740 5.170 16.220 5.400 ;
        RECT 15.740 5.100 16.080 5.170 ;
    END
  END SELECT1
  PIN SELECT3
    ANTENNAGATEAREA 0.730000 ;
    PORT
      LAYER met2 ;
        RECT 15.740 1.970 16.220 2.200 ;
        RECT 15.740 1.900 16.080 1.970 ;
    END
  END SELECT3
  PIN SELECT4
    ANTENNAGATEAREA 0.730000 ;
    PORT
      LAYER met2 ;
        RECT 15.740 0.860 16.080 0.930 ;
        RECT 15.740 0.630 16.220 0.860 ;
    END
  END SELECT4
  OBS
      LAYER li1 ;
        RECT 10.720 5.090 10.890 5.980 ;
        RECT 11.120 5.000 11.290 5.930 ;
        RECT 14.810 5.860 15.050 5.890 ;
        RECT 11.820 5.690 12.780 5.860 ;
        RECT 13.230 5.690 14.570 5.860 ;
        RECT 14.810 5.690 15.380 5.860 ;
        RECT 12.100 5.680 12.270 5.690 ;
        RECT 14.810 5.650 15.050 5.690 ;
        RECT 15.690 5.560 15.860 5.980 ;
        RECT 12.300 5.240 12.640 5.420 ;
        RECT 15.760 5.340 15.930 5.380 ;
        RECT 15.400 5.240 15.590 5.260 ;
        RECT 11.820 5.070 14.570 5.240 ;
        RECT 15.030 5.070 15.590 5.240 ;
        RECT 15.400 5.030 15.590 5.070 ;
        RECT 15.760 5.170 15.990 5.340 ;
        RECT 15.760 4.820 15.930 5.170 ;
        RECT 10.720 3.250 10.890 4.140 ;
        RECT 11.120 3.300 11.290 4.230 ;
        RECT 15.400 4.160 15.590 4.200 ;
        RECT 11.820 3.990 14.570 4.160 ;
        RECT 15.030 3.990 15.590 4.160 ;
        RECT 12.300 3.810 12.640 3.990 ;
        RECT 15.400 3.970 15.590 3.990 ;
        RECT 15.760 4.060 15.930 4.410 ;
        RECT 15.760 3.890 15.990 4.060 ;
        RECT 15.760 3.850 15.930 3.890 ;
        RECT 12.100 3.540 12.270 3.550 ;
        RECT 14.810 3.540 15.050 3.580 ;
        RECT 11.820 3.370 12.780 3.540 ;
        RECT 13.230 3.370 14.570 3.540 ;
        RECT 14.810 3.370 15.380 3.540 ;
        RECT 14.810 3.340 15.050 3.370 ;
        RECT 15.690 3.250 15.860 3.670 ;
        RECT 10.720 1.890 10.890 2.780 ;
        RECT 11.120 1.800 11.290 2.730 ;
        RECT 14.810 2.660 15.050 2.690 ;
        RECT 11.820 2.490 12.780 2.660 ;
        RECT 13.230 2.490 14.570 2.660 ;
        RECT 14.810 2.490 15.380 2.660 ;
        RECT 12.100 2.480 12.270 2.490 ;
        RECT 14.810 2.450 15.050 2.490 ;
        RECT 15.690 2.360 15.860 2.780 ;
        RECT 12.300 2.040 12.640 2.220 ;
        RECT 15.760 2.140 15.930 2.180 ;
        RECT 15.400 2.040 15.590 2.060 ;
        RECT 11.820 1.870 14.570 2.040 ;
        RECT 15.030 1.870 15.590 2.040 ;
        RECT 15.400 1.830 15.590 1.870 ;
        RECT 15.760 1.970 15.990 2.140 ;
        RECT 15.760 1.620 15.930 1.970 ;
        RECT 10.720 0.050 10.890 0.940 ;
        RECT 11.120 0.100 11.290 1.030 ;
        RECT 15.400 0.960 15.590 1.000 ;
        RECT 11.820 0.790 14.570 0.960 ;
        RECT 15.030 0.790 15.590 0.960 ;
        RECT 12.300 0.610 12.640 0.790 ;
        RECT 15.400 0.770 15.590 0.790 ;
        RECT 15.760 0.860 15.930 1.210 ;
        RECT 15.760 0.690 15.990 0.860 ;
        RECT 15.760 0.650 15.930 0.690 ;
        RECT 12.100 0.340 12.270 0.350 ;
        RECT 14.810 0.340 15.050 0.380 ;
        RECT 11.820 0.170 12.780 0.340 ;
        RECT 13.230 0.170 14.570 0.340 ;
        RECT 14.810 0.170 15.380 0.340 ;
        RECT 14.810 0.140 15.050 0.170 ;
        RECT 15.690 0.050 15.860 0.470 ;
      LAYER mcon ;
        RECT 10.720 5.810 10.890 5.980 ;
        RECT 10.720 5.450 10.890 5.620 ;
        RECT 14.100 5.690 14.270 5.860 ;
        RECT 14.850 5.690 15.020 5.860 ;
        RECT 15.690 5.810 15.860 5.980 ;
        RECT 11.120 5.360 11.290 5.530 ;
        RECT 15.410 5.060 15.580 5.230 ;
        RECT 15.820 5.170 15.990 5.340 ;
        RECT 10.720 3.970 10.890 4.140 ;
        RECT 10.720 3.610 10.890 3.780 ;
        RECT 15.410 4.000 15.580 4.170 ;
        RECT 11.120 3.700 11.290 3.870 ;
        RECT 15.820 3.890 15.990 4.060 ;
        RECT 12.100 3.380 12.270 3.550 ;
        RECT 14.100 3.370 14.270 3.540 ;
        RECT 14.850 3.370 15.020 3.540 ;
        RECT 10.720 2.610 10.890 2.780 ;
        RECT 10.720 2.250 10.890 2.420 ;
        RECT 14.100 2.490 14.270 2.660 ;
        RECT 14.850 2.490 15.020 2.660 ;
        RECT 15.690 2.610 15.860 2.780 ;
        RECT 11.120 2.160 11.290 2.330 ;
        RECT 15.410 1.860 15.580 2.030 ;
        RECT 15.820 1.970 15.990 2.140 ;
        RECT 10.720 0.770 10.890 0.940 ;
        RECT 10.720 0.410 10.890 0.580 ;
        RECT 15.410 0.800 15.580 0.970 ;
        RECT 11.120 0.500 11.290 0.670 ;
        RECT 15.820 0.690 15.990 0.860 ;
        RECT 12.100 0.180 12.270 0.350 ;
        RECT 14.100 0.170 14.270 0.340 ;
        RECT 14.850 0.170 15.020 0.340 ;
      LAYER met1 ;
        RECT 12.230 5.880 12.570 5.930 ;
        RECT 12.010 5.860 12.570 5.880 ;
        RECT 14.660 5.900 15.030 5.920 ;
        RECT 12.010 5.690 12.690 5.860 ;
        RECT 12.010 5.650 12.570 5.690 ;
        RECT 12.230 5.610 12.570 5.650 ;
        RECT 14.660 5.640 15.080 5.900 ;
        RECT 14.660 5.630 15.030 5.640 ;
        RECT 15.750 5.110 16.070 5.390 ;
        RECT 15.750 3.840 16.070 4.120 ;
        RECT 12.230 3.580 12.570 3.620 ;
        RECT 12.010 3.540 12.570 3.580 ;
        RECT 14.660 3.590 15.030 3.600 ;
        RECT 12.010 3.370 12.690 3.540 ;
        RECT 12.010 3.350 12.570 3.370 ;
        RECT 12.230 3.300 12.570 3.350 ;
        RECT 14.660 3.330 15.080 3.590 ;
        RECT 14.660 3.310 15.030 3.330 ;
        RECT 12.230 2.680 12.570 2.730 ;
        RECT 12.010 2.660 12.570 2.680 ;
        RECT 14.660 2.700 15.030 2.720 ;
        RECT 12.010 2.490 12.690 2.660 ;
        RECT 12.010 2.450 12.570 2.490 ;
        RECT 12.230 2.410 12.570 2.450 ;
        RECT 14.660 2.440 15.080 2.700 ;
        RECT 14.660 2.430 15.030 2.440 ;
        RECT 15.750 1.910 16.070 2.190 ;
        RECT 15.750 0.640 16.070 0.920 ;
        RECT 12.230 0.380 12.570 0.420 ;
        RECT 12.010 0.340 12.570 0.380 ;
        RECT 14.660 0.390 15.030 0.400 ;
        RECT 12.010 0.170 12.690 0.340 ;
        RECT 12.010 0.150 12.570 0.170 ;
        RECT 12.230 0.100 12.570 0.150 ;
        RECT 14.660 0.130 15.080 0.390 ;
        RECT 14.660 0.110 15.030 0.130 ;
      LAYER via ;
        RECT 12.280 5.640 12.540 5.900 ;
        RECT 14.690 5.640 14.950 5.900 ;
        RECT 15.780 5.120 16.040 5.380 ;
        RECT 15.780 3.850 16.040 4.110 ;
        RECT 12.280 3.330 12.540 3.590 ;
        RECT 14.690 3.330 14.950 3.590 ;
        RECT 12.280 2.440 12.540 2.700 ;
        RECT 14.690 2.440 14.950 2.700 ;
        RECT 15.780 1.920 16.040 2.180 ;
        RECT 15.780 0.650 16.040 0.910 ;
        RECT 12.280 0.130 12.540 0.390 ;
        RECT 14.690 0.130 14.950 0.390 ;
      LAYER met2 ;
        RECT 12.250 5.880 12.570 5.900 ;
        RECT 14.660 5.880 14.980 5.930 ;
        RECT 12.250 5.850 14.980 5.880 ;
        RECT 10.500 5.690 14.980 5.850 ;
        RECT 10.500 5.670 12.570 5.690 ;
        RECT 12.250 5.640 12.570 5.670 ;
        RECT 14.660 5.610 14.980 5.690 ;
        RECT 12.250 3.540 12.570 3.590 ;
        RECT 14.660 3.540 14.980 3.620 ;
        RECT 12.250 3.530 14.980 3.540 ;
        RECT 10.500 3.370 14.980 3.530 ;
        RECT 12.250 3.350 14.980 3.370 ;
        RECT 12.250 3.330 12.570 3.350 ;
        RECT 14.660 3.300 14.980 3.350 ;
        RECT 12.250 0.340 12.570 0.390 ;
        RECT 14.660 0.340 14.980 0.420 ;
        RECT 12.250 0.320 14.980 0.340 ;
        RECT 10.500 0.150 14.980 0.320 ;
        RECT 12.250 0.130 12.570 0.150 ;
        RECT 14.660 0.100 14.980 0.150 ;
  END
END sky130_hilas_drainSelect01

MACRO sky130_hilas_VinjInv2
  CLASS BLOCK ;
  FOREIGN sky130_hilas_VinjInv2 ;
  ORIGIN 3.360 -1.440 ;
  SIZE 3.610 BY 1.640 ;
  OBS
      LAYER nwell ;
        RECT -3.360 1.440 -1.380 3.080 ;
      LAYER li1 ;
        RECT -2.740 2.650 -2.570 2.790 ;
        RECT -2.740 2.480 -2.550 2.650 ;
        RECT -2.740 2.380 -2.570 2.480 ;
        RECT -3.170 2.000 -3.000 2.100 ;
        RECT -3.190 1.830 -3.000 2.000 ;
        RECT -3.170 1.770 -3.000 1.830 ;
        RECT -2.750 2.040 -2.580 2.100 ;
        RECT -2.750 1.770 -2.500 2.040 ;
        RECT -2.010 2.020 -1.760 2.100 ;
        RECT -2.010 1.850 -0.710 2.020 ;
        RECT -0.150 2.010 0.020 2.640 ;
        RECT -2.740 1.750 -2.500 1.770 ;
        RECT -1.930 1.760 -1.760 1.850 ;
        RECT -0.230 1.840 0.100 2.010 ;
      LAYER mcon ;
        RECT -2.720 2.480 -2.550 2.650 ;
        RECT -0.150 2.120 0.020 2.290 ;
        RECT -2.710 1.800 -2.540 1.970 ;
        RECT -1.370 1.850 -1.200 2.020 ;
      LAYER met1 ;
        RECT -2.750 2.700 -2.530 3.040 ;
        RECT -2.750 2.440 -2.520 2.700 ;
        RECT -3.280 1.760 -2.970 2.110 ;
        RECT -2.750 2.040 -2.530 2.440 ;
        RECT -2.750 1.730 -2.500 2.040 ;
        RECT -1.450 1.800 -1.130 2.060 ;
        RECT -2.750 1.530 -2.530 1.730 ;
        RECT -0.180 1.530 0.050 3.040 ;
      LAYER via ;
        RECT -3.250 1.790 -2.990 2.050 ;
        RECT -1.420 1.800 -1.160 2.060 ;
      LAYER met2 ;
        RECT -3.360 2.470 0.250 2.650 ;
        RECT -3.280 1.950 -2.960 2.050 ;
        RECT -3.290 1.790 -2.960 1.950 ;
        RECT -1.450 1.980 -1.130 2.060 ;
        RECT -1.450 1.800 0.250 1.980 ;
  END
END sky130_hilas_VinjInv2

MACRO sky130_hilas_cellAttempt01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_cellAttempt01 ;
  ORIGIN 2.630 4.040 ;
  SIZE 10.070 BY 6.500 ;
  PIN VTUN
    ANTENNADIFFAREA 2.237600 ;
    PORT
      LAYER nwell ;
        RECT -2.630 -4.040 -0.900 2.450 ;
      LAYER met1 ;
        RECT -2.280 -4.040 -1.880 2.460 ;
    END
  END VTUN
  PIN VINJ
    ANTENNADIFFAREA 1.088000 ;
    PORT
      LAYER nwell ;
        RECT 4.880 -4.040 7.440 2.460 ;
      LAYER met1 ;
        RECT 6.920 1.750 7.080 2.450 ;
        RECT 6.810 1.200 7.080 1.750 ;
        RECT 6.810 1.150 7.090 1.200 ;
        RECT 6.920 1.060 7.090 1.150 ;
        RECT 6.920 0.590 7.080 1.060 ;
        RECT 6.920 0.500 7.090 0.590 ;
        RECT 6.810 0.450 7.090 0.500 ;
        RECT 6.810 -0.100 7.080 0.450 ;
        RECT 6.920 -1.490 7.080 -0.100 ;
        RECT 6.810 -2.040 7.080 -1.490 ;
        RECT 6.810 -2.090 7.090 -2.040 ;
        RECT 6.920 -2.180 7.090 -2.090 ;
        RECT 6.920 -2.640 7.080 -2.180 ;
        RECT 6.920 -2.730 7.090 -2.640 ;
        RECT 6.810 -2.780 7.090 -2.730 ;
        RECT 6.810 -3.330 7.080 -2.780 ;
        RECT 6.920 -4.030 7.080 -3.330 ;
    END
  END VINJ
  PIN COLSEL1
    ANTENNAGATEAREA 0.720000 ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met1 ;
        RECT 6.110 1.720 6.270 2.450 ;
        RECT 6.110 1.700 6.310 1.720 ;
        RECT 6.090 1.460 6.320 1.700 ;
        RECT 6.110 1.410 6.320 1.460 ;
        RECT 6.480 1.410 6.670 2.400 ;
        RECT 6.110 0.240 6.270 1.410 ;
        RECT 6.500 1.290 6.670 1.410 ;
        RECT 6.510 0.360 6.670 1.290 ;
        RECT 6.500 0.240 6.670 0.360 ;
        RECT 6.110 0.190 6.320 0.240 ;
        RECT 6.090 -0.050 6.320 0.190 ;
        RECT 6.110 -0.070 6.310 -0.050 ;
        RECT 6.110 -0.700 6.270 -0.070 ;
        RECT 6.480 -0.680 6.670 0.240 ;
        RECT 6.460 -0.700 6.700 -0.680 ;
        RECT 6.110 -0.890 6.700 -0.700 ;
        RECT 6.110 -1.520 6.270 -0.890 ;
        RECT 6.460 -0.910 6.700 -0.890 ;
        RECT 6.110 -1.540 6.310 -1.520 ;
        RECT 6.090 -1.780 6.320 -1.540 ;
        RECT 6.110 -1.830 6.320 -1.780 ;
        RECT 6.480 -1.830 6.670 -0.910 ;
        RECT 6.110 -2.990 6.270 -1.830 ;
        RECT 6.500 -1.950 6.670 -1.830 ;
        RECT 6.510 -2.870 6.670 -1.950 ;
        RECT 6.500 -2.990 6.670 -2.870 ;
        RECT 6.110 -3.040 6.320 -2.990 ;
        RECT 6.090 -3.280 6.320 -3.040 ;
        RECT 6.110 -3.300 6.310 -3.280 ;
        RECT 6.110 -4.030 6.270 -3.300 ;
        RECT 6.480 -3.980 6.670 -2.990 ;
    END
  END COLSEL1
  PIN GATE1
    ANTENNADIFFAREA 3.253900 ;
    PORT
      LAYER nwell ;
        RECT 1.120 -4.040 3.350 2.450 ;
      LAYER met1 ;
        RECT 1.770 0.310 2.150 2.460 ;
        RECT 1.760 -1.550 2.150 0.310 ;
        RECT 1.770 -4.040 2.150 -1.550 ;
    END
  END GATE1
  PIN ROW4
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 4.970 -2.870 5.280 -2.740 ;
        RECT -2.630 -3.050 7.440 -2.870 ;
        RECT 4.970 -3.070 5.280 -3.050 ;
    END
  END ROW4
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.120 -2.260 0.440 -2.250 ;
        RECT 4.050 -2.260 4.370 -2.200 ;
        RECT 0.120 -2.440 4.370 -2.260 ;
        RECT 0.120 -2.510 0.440 -2.440 ;
        RECT 4.050 -2.490 4.370 -2.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.090 1.070 4.330 2.460 ;
        RECT 4.070 0.410 4.340 1.070 ;
        RECT 4.090 -2.180 4.330 0.410 ;
        RECT 4.080 -2.500 4.340 -2.180 ;
        RECT 4.090 -4.040 4.330 -2.500 ;
      LAYER via ;
        RECT 4.080 -2.470 4.340 -2.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.160 1.050 0.400 2.460 ;
        RECT 0.150 0.390 0.410 1.050 ;
        RECT 0.160 -2.220 0.400 0.390 ;
        RECT 0.150 -2.540 0.410 -2.220 ;
        RECT 0.160 -4.040 0.400 -2.540 ;
      LAYER via ;
        RECT 0.150 -2.510 0.410 -2.250 ;
    END
  END VGND
  PIN DRAIN4
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 4.970 -3.300 5.280 -3.290 ;
        RECT -2.630 -3.470 7.440 -3.300 ;
        RECT 4.970 -3.480 7.440 -3.470 ;
        RECT 4.970 -3.620 5.280 -3.480 ;
    END
  END DRAIN4
  PIN DRAIN1
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 4.970 1.900 5.280 2.040 ;
        RECT -2.630 1.720 7.440 1.900 ;
        RECT 4.970 1.710 5.280 1.720 ;
    END
  END DRAIN1
  PIN ROW1
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 4.970 1.470 5.280 1.490 ;
        RECT 4.880 1.460 7.440 1.470 ;
        RECT -2.630 1.290 7.440 1.460 ;
        RECT -2.630 1.280 5.280 1.290 ;
        RECT 4.970 1.160 5.280 1.280 ;
    END
  END ROW1
  PIN ROW3
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 4.970 -1.770 5.280 -1.750 ;
        RECT -2.630 -1.950 7.440 -1.770 ;
        RECT 4.970 -2.080 5.280 -1.950 ;
    END
  END ROW3
  PIN DRAIN3
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 4.970 -1.340 5.280 -1.200 ;
        RECT -2.630 -1.520 7.440 -1.340 ;
        RECT 4.970 -1.530 5.280 -1.520 ;
    END
  END DRAIN3
  PIN DRAIN2
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 4.970 -0.070 5.280 -0.060 ;
        RECT -2.630 -0.250 7.440 -0.070 ;
        RECT 4.970 -0.390 5.280 -0.250 ;
    END
  END DRAIN2
  PIN ROW2
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 4.970 0.360 5.280 0.490 ;
        RECT -2.630 0.180 7.440 0.360 ;
        RECT 4.970 0.160 5.280 0.180 ;
    END
  END ROW2
  OBS
      LAYER li1 ;
        RECT 4.980 1.990 5.300 2.000 ;
        RECT 4.980 1.820 5.560 1.990 ;
        RECT 4.980 1.770 5.310 1.820 ;
        RECT 4.980 1.740 5.300 1.770 ;
        RECT 6.840 1.720 7.040 2.070 ;
        RECT 4.980 1.410 5.300 1.450 ;
        RECT 4.980 1.370 5.310 1.410 ;
        RECT 4.980 1.200 5.560 1.370 ;
        RECT 4.980 1.190 5.300 1.200 ;
        RECT 6.110 1.100 6.310 1.700 ;
        RECT 6.840 1.690 7.050 1.720 ;
        RECT 6.830 1.100 7.050 1.690 ;
        RECT 0.190 0.480 0.360 1.010 ;
        RECT 4.130 0.470 4.300 1.000 ;
        RECT 4.980 0.450 5.300 0.460 ;
        RECT 4.980 0.280 5.560 0.450 ;
        RECT 4.980 0.240 5.310 0.280 ;
        RECT 4.980 0.200 5.300 0.240 ;
        RECT 6.110 -0.050 6.310 0.550 ;
        RECT 6.830 -0.040 7.050 0.550 ;
        RECT 6.840 -0.070 7.050 -0.040 ;
        RECT 4.980 -0.120 5.300 -0.090 ;
        RECT 4.980 -0.170 5.310 -0.120 ;
        RECT -2.210 -1.020 -1.660 -0.590 ;
        RECT 0.200 -1.230 0.370 -0.220 ;
        RECT 4.980 -0.340 5.560 -0.170 ;
        RECT 4.980 -0.350 5.300 -0.340 ;
        RECT 1.820 -1.090 2.370 -0.660 ;
        RECT 4.130 -1.370 4.300 -0.360 ;
        RECT 6.840 -0.420 7.040 -0.070 ;
        RECT 6.230 -0.880 6.670 -0.710 ;
        RECT 4.980 -1.250 5.300 -1.240 ;
        RECT 4.980 -1.420 5.560 -1.250 ;
        RECT 4.980 -1.470 5.310 -1.420 ;
        RECT 4.980 -1.500 5.300 -1.470 ;
        RECT 6.840 -1.520 7.040 -1.170 ;
        RECT 4.980 -1.830 5.300 -1.790 ;
        RECT 4.980 -1.870 5.310 -1.830 ;
        RECT 4.980 -2.040 5.560 -1.870 ;
        RECT 4.980 -2.050 5.300 -2.040 ;
        RECT 6.110 -2.140 6.310 -1.540 ;
        RECT 6.840 -1.550 7.050 -1.520 ;
        RECT 6.830 -2.140 7.050 -1.550 ;
        RECT 4.980 -2.780 5.300 -2.770 ;
        RECT 4.980 -2.950 5.560 -2.780 ;
        RECT 4.980 -2.990 5.310 -2.950 ;
        RECT 4.980 -3.030 5.300 -2.990 ;
        RECT 6.110 -3.280 6.310 -2.680 ;
        RECT 6.830 -3.270 7.050 -2.680 ;
        RECT 6.840 -3.300 7.050 -3.270 ;
        RECT 4.980 -3.350 5.300 -3.320 ;
        RECT 4.980 -3.400 5.310 -3.350 ;
        RECT 4.980 -3.570 5.560 -3.400 ;
        RECT 4.980 -3.580 5.300 -3.570 ;
        RECT 6.840 -3.650 7.040 -3.300 ;
      LAYER mcon ;
        RECT 5.040 1.780 5.210 1.950 ;
        RECT 6.120 1.490 6.290 1.660 ;
        RECT 5.040 1.230 5.210 1.400 ;
        RECT 6.850 1.520 7.020 1.690 ;
        RECT 0.190 0.840 0.360 1.010 ;
        RECT 4.130 0.830 4.300 1.000 ;
        RECT 5.040 0.250 5.210 0.420 ;
        RECT 6.120 -0.010 6.290 0.160 ;
        RECT 6.850 -0.040 7.020 0.130 ;
        RECT 5.040 -0.300 5.210 -0.130 ;
        RECT -2.210 -0.940 -1.940 -0.670 ;
        RECT 0.200 -0.620 0.370 -0.450 ;
        RECT 0.200 -0.980 0.370 -0.810 ;
        RECT 1.820 -1.010 2.090 -0.740 ;
        RECT 4.130 -0.760 4.300 -0.590 ;
        RECT 6.490 -0.880 6.670 -0.710 ;
        RECT 4.130 -1.120 4.300 -0.950 ;
        RECT 5.040 -1.460 5.210 -1.290 ;
        RECT 6.120 -1.750 6.290 -1.580 ;
        RECT 5.040 -2.010 5.210 -1.840 ;
        RECT 6.850 -1.720 7.020 -1.550 ;
        RECT 5.040 -2.980 5.210 -2.810 ;
        RECT 6.120 -3.240 6.290 -3.070 ;
        RECT 6.850 -3.270 7.020 -3.100 ;
        RECT 5.040 -3.530 5.210 -3.360 ;
      LAYER met1 ;
        RECT 4.970 1.710 5.290 2.030 ;
        RECT 4.970 1.160 5.290 1.480 ;
        RECT 4.970 0.170 5.290 0.490 ;
        RECT 4.970 -0.380 5.290 -0.060 ;
        RECT 4.970 -1.530 5.290 -1.210 ;
        RECT 4.970 -2.080 5.290 -1.760 ;
        RECT 4.970 -3.060 5.290 -2.740 ;
        RECT 4.970 -3.610 5.290 -3.290 ;
      LAYER via ;
        RECT 5.000 1.740 5.260 2.000 ;
        RECT 5.000 1.190 5.260 1.450 ;
        RECT 5.000 0.200 5.260 0.460 ;
        RECT 5.000 -0.350 5.260 -0.090 ;
        RECT 5.000 -1.500 5.260 -1.240 ;
        RECT 5.000 -2.050 5.260 -1.790 ;
        RECT 5.000 -3.030 5.260 -2.770 ;
        RECT 5.000 -3.580 5.260 -3.320 ;
  END
END sky130_hilas_cellAttempt01

MACRO sky130_hilas_DAC5bit01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_DAC5bit01 ;
  ORIGIN -3.820 -5.240 ;
  SIZE 16.580 BY 5.990 ;
  PIN A0
    USE ANALOG ;
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER met2 ;
        RECT 12.080 6.230 12.400 6.260 ;
        RECT 3.820 6.030 12.400 6.230 ;
        RECT 12.080 6.000 12.400 6.030 ;
    END
  END A0
  PIN A1
    USE ANALOG ;
    ANTENNAGATEAREA 0.456300 ;
    PORT
      LAYER met2 ;
        RECT 15.410 10.910 15.730 11.230 ;
        RECT 15.530 7.350 15.680 10.910 ;
        RECT 3.820 7.150 15.690 7.350 ;
        RECT 3.820 7.140 3.960 7.150 ;
    END
  END A1
  PIN A2
    USE ANALOG ;
    ANTENNAGATEAREA 0.608400 ;
    PORT
      LAYER met2 ;
        RECT 13.800 10.930 14.120 11.230 ;
        RECT 13.800 10.910 14.130 10.930 ;
        RECT 13.930 8.330 14.130 10.910 ;
        RECT 3.820 8.120 14.130 8.330 ;
    END
  END A2
  PIN A3
    USE ANALOG ;
    ANTENNAGATEAREA 2.281500 ;
    PORT
      LAYER met2 ;
        RECT 12.190 10.900 12.510 11.220 ;
        RECT 7.310 10.660 7.630 10.810 ;
        RECT 7.300 10.490 7.630 10.660 ;
        RECT 3.820 10.200 5.880 10.260 ;
        RECT 7.300 10.200 7.520 10.490 ;
        RECT 12.220 10.210 12.470 10.900 ;
        RECT 12.220 10.200 12.500 10.210 ;
        RECT 3.820 10.050 12.500 10.200 ;
        RECT 4.080 9.870 4.280 10.050 ;
        RECT 5.720 9.900 12.500 10.050 ;
        RECT 4.030 9.550 4.350 9.870 ;
    END
  END A3
  PIN A4
    USE ANALOG ;
    ANTENNAGATEAREA 3.650400 ;
    PORT
      LAYER met2 ;
        RECT 5.760 11.210 6.080 11.220 ;
        RECT 8.960 11.210 9.280 11.220 ;
        RECT 10.570 11.210 10.890 11.230 ;
        RECT 3.820 11.020 10.890 11.210 ;
        RECT 3.820 11.000 4.370 11.020 ;
        RECT 4.050 10.860 4.370 11.000 ;
        RECT 5.760 10.900 6.080 11.020 ;
        RECT 8.960 10.900 9.280 11.020 ;
        RECT 10.570 10.910 10.890 11.020 ;
    END
  END A4
  PIN VPWR
    USE ANALOG ;
    ANTENNADIFFAREA 3.264300 ;
    PORT
      LAYER met2 ;
        RECT 16.530 10.930 17.690 11.210 ;
        RECT 16.650 10.750 16.960 10.930 ;
        RECT 17.280 10.920 17.690 10.930 ;
        RECT 17.320 10.750 17.630 10.920 ;
    END
  END VPWR
  PIN OUT
    USE ANALOG ;
    ANTENNADIFFAREA 3.264300 ;
    PORT
      LAYER met1 ;
        RECT 6.830 5.480 7.060 5.530 ;
        RECT 8.450 5.480 8.680 5.530 ;
        RECT 10.050 5.480 10.280 5.530 ;
        RECT 11.670 5.480 11.900 5.530 ;
        RECT 13.270 5.480 13.500 5.530 ;
        RECT 14.890 5.480 15.120 5.530 ;
        RECT 16.490 5.480 16.720 5.530 ;
        RECT 18.100 5.480 18.330 5.530 ;
        RECT 6.830 5.250 20.400 5.480 ;
        RECT 6.830 5.240 7.060 5.250 ;
        RECT 8.450 5.240 8.680 5.250 ;
        RECT 10.050 5.240 10.280 5.250 ;
        RECT 11.670 5.240 11.900 5.250 ;
        RECT 13.270 5.240 13.500 5.250 ;
        RECT 14.890 5.240 15.120 5.250 ;
        RECT 16.490 5.240 16.720 5.250 ;
        RECT 18.100 5.240 18.330 5.250 ;
    END
  END OUT
  OBS
      LAYER nwell ;
        RECT 4.190 5.270 20.290 10.920 ;
      LAYER li1 ;
        RECT 4.100 10.710 4.310 11.140 ;
        RECT 5.810 10.750 6.020 11.180 ;
        RECT 5.830 10.730 6.000 10.750 ;
        RECT 7.160 10.740 7.590 10.760 ;
        RECT 9.010 10.750 9.220 11.180 ;
        RECT 10.620 10.760 10.830 11.190 ;
        RECT 4.120 10.690 4.290 10.710 ;
        RECT 7.140 10.570 7.590 10.740 ;
        RECT 9.030 10.730 9.200 10.750 ;
        RECT 10.640 10.740 10.810 10.760 ;
        RECT 12.240 10.750 12.450 11.180 ;
        RECT 13.850 10.760 14.060 11.190 ;
        RECT 15.460 10.760 15.670 11.190 ;
        RECT 16.770 11.040 16.980 11.050 ;
        RECT 16.660 11.000 16.980 11.040 ;
        RECT 17.330 11.000 17.650 11.040 ;
        RECT 16.660 10.810 16.990 11.000 ;
        RECT 17.330 10.810 17.660 11.000 ;
        RECT 16.660 10.780 16.980 10.810 ;
        RECT 17.330 10.780 17.650 10.810 ;
        RECT 12.260 10.730 12.430 10.750 ;
        RECT 13.870 10.740 14.040 10.760 ;
        RECT 15.480 10.740 15.650 10.760 ;
        RECT 7.160 10.550 7.590 10.570 ;
        RECT 7.800 10.270 7.970 10.280 ;
        RECT 16.770 10.270 16.980 10.780 ;
        RECT 17.440 10.270 17.610 10.780 ;
        RECT 6.190 10.040 17.620 10.270 ;
        RECT 4.080 9.400 4.290 9.830 ;
        RECT 6.190 9.700 6.360 10.040 ;
        RECT 4.100 9.380 4.270 9.400 ;
        RECT 6.180 9.370 6.360 9.700 ;
        RECT 4.100 8.450 4.310 8.880 ;
        RECT 6.190 8.740 6.360 9.370 ;
        RECT 4.120 8.430 4.290 8.450 ;
        RECT 6.180 8.410 6.360 8.740 ;
        RECT 4.100 7.510 4.310 7.940 ;
        RECT 6.190 7.780 6.360 8.410 ;
        RECT 4.120 7.490 4.290 7.510 ;
        RECT 6.180 7.450 6.360 7.780 ;
        RECT 6.190 6.820 6.360 7.450 ;
        RECT 6.180 6.490 6.360 6.820 ;
        RECT 6.190 6.480 6.360 6.490 ;
        RECT 6.850 9.700 7.020 9.710 ;
        RECT 7.800 9.700 7.970 10.040 ;
        RECT 9.390 9.700 9.560 10.040 ;
        RECT 6.850 9.370 7.030 9.700 ;
        RECT 7.790 9.370 7.970 9.700 ;
        RECT 8.470 9.670 8.640 9.700 ;
        RECT 8.470 9.370 8.650 9.670 ;
        RECT 6.850 8.740 7.020 9.370 ;
        RECT 7.800 8.740 7.970 9.370 ;
        RECT 8.480 8.740 8.650 9.370 ;
        RECT 6.850 8.410 7.030 8.740 ;
        RECT 7.790 8.410 7.970 8.740 ;
        RECT 8.470 8.410 8.650 8.740 ;
        RECT 6.850 7.780 7.020 8.410 ;
        RECT 7.800 7.780 7.970 8.410 ;
        RECT 8.480 7.780 8.650 8.410 ;
        RECT 6.850 7.450 7.030 7.780 ;
        RECT 7.790 7.450 7.970 7.780 ;
        RECT 8.470 7.450 8.650 7.780 ;
        RECT 6.850 6.820 7.020 7.450 ;
        RECT 7.800 6.820 7.970 7.450 ;
        RECT 8.480 6.820 8.650 7.450 ;
        RECT 6.850 6.490 7.030 6.820 ;
        RECT 7.790 6.490 7.970 6.820 ;
        RECT 8.470 6.490 8.650 6.820 ;
        RECT 6.850 5.500 7.020 6.490 ;
        RECT 7.800 6.480 7.970 6.490 ;
        RECT 8.480 5.500 8.650 6.490 ;
        RECT 9.390 9.370 9.570 9.700 ;
        RECT 9.390 8.740 9.560 9.370 ;
        RECT 9.390 8.410 9.570 8.740 ;
        RECT 9.390 7.780 9.560 8.410 ;
        RECT 9.390 7.450 9.570 7.780 ;
        RECT 9.390 6.820 9.560 7.450 ;
        RECT 9.390 6.490 9.570 6.820 ;
        RECT 9.390 6.480 9.560 6.490 ;
        RECT 10.080 5.500 10.250 9.750 ;
        RECT 10.540 8.460 10.750 8.890 ;
        RECT 10.560 8.440 10.730 8.460 ;
        RECT 11.010 6.480 11.180 10.040 ;
        RECT 12.630 9.700 12.800 10.040 ;
        RECT 11.690 9.370 11.870 9.700 ;
        RECT 12.620 9.370 12.800 9.700 ;
        RECT 11.700 8.740 11.870 9.370 ;
        RECT 12.630 8.740 12.800 9.370 ;
        RECT 11.690 8.410 11.870 8.740 ;
        RECT 12.620 8.410 12.800 8.740 ;
        RECT 11.700 7.780 11.870 8.410 ;
        RECT 12.140 7.980 12.310 8.000 ;
        RECT 11.690 7.450 11.870 7.780 ;
        RECT 12.120 7.550 12.330 7.980 ;
        RECT 11.700 6.820 11.870 7.450 ;
        RECT 12.630 6.820 12.800 8.410 ;
        RECT 11.690 6.490 11.870 6.820 ;
        RECT 12.620 6.500 12.800 6.820 ;
        RECT 12.620 6.490 12.790 6.500 ;
        RECT 11.700 5.500 11.870 6.490 ;
        RECT 13.300 5.500 13.470 9.750 ;
        RECT 13.760 6.550 13.970 6.980 ;
        RECT 13.780 6.530 13.950 6.550 ;
        RECT 14.230 6.490 14.400 10.040 ;
        RECT 14.920 9.700 15.090 9.750 ;
        RECT 14.910 9.370 15.090 9.700 ;
        RECT 14.920 8.740 15.090 9.370 ;
        RECT 14.910 8.410 15.090 8.740 ;
        RECT 14.920 7.780 15.090 8.410 ;
        RECT 14.910 7.450 15.090 7.780 ;
        RECT 14.920 6.820 15.090 7.450 ;
        RECT 14.910 6.490 15.090 6.820 ;
        RECT 15.840 6.490 16.010 10.040 ;
        RECT 14.920 5.500 15.090 6.490 ;
        RECT 16.520 5.500 16.690 9.730 ;
        RECT 17.450 6.470 17.620 10.040 ;
        RECT 18.130 5.500 18.300 9.910 ;
        RECT 6.850 5.270 7.040 5.500 ;
        RECT 8.470 5.270 8.660 5.500 ;
        RECT 10.070 5.270 10.260 5.500 ;
        RECT 11.690 5.270 11.880 5.500 ;
        RECT 13.290 5.270 13.480 5.500 ;
        RECT 14.910 5.270 15.100 5.500 ;
        RECT 16.510 5.270 16.700 5.500 ;
        RECT 18.120 5.270 18.310 5.500 ;
        RECT 6.850 5.250 7.020 5.270 ;
        RECT 8.480 5.250 8.650 5.270 ;
        RECT 10.080 5.250 10.250 5.270 ;
        RECT 11.700 5.250 11.870 5.270 ;
        RECT 13.300 5.250 13.470 5.270 ;
        RECT 14.920 5.250 15.090 5.270 ;
        RECT 16.520 5.250 16.690 5.270 ;
        RECT 18.130 5.250 18.300 5.270 ;
      LAYER mcon ;
        RECT 16.720 10.820 16.890 10.990 ;
        RECT 17.390 10.820 17.560 10.990 ;
        RECT 12.140 7.830 12.310 8.000 ;
        RECT 6.860 5.300 7.030 5.470 ;
        RECT 8.480 5.300 8.650 5.470 ;
        RECT 10.080 5.300 10.250 5.470 ;
        RECT 11.700 5.300 11.870 5.470 ;
        RECT 13.300 5.300 13.470 5.470 ;
        RECT 14.920 5.300 15.090 5.470 ;
        RECT 16.520 5.300 16.690 5.470 ;
        RECT 18.130 5.300 18.300 5.470 ;
      LAYER met1 ;
        RECT 4.050 10.860 4.370 11.180 ;
        RECT 5.760 10.900 6.080 11.220 ;
        RECT 8.960 10.900 9.280 11.220 ;
        RECT 10.570 10.910 10.890 11.230 ;
        RECT 4.090 10.630 4.320 10.860 ;
        RECT 5.800 10.670 6.030 10.900 ;
        RECT 7.310 10.770 7.630 10.810 ;
        RECT 7.080 10.540 7.630 10.770 ;
        RECT 9.000 10.670 9.230 10.900 ;
        RECT 10.610 10.680 10.840 10.910 ;
        RECT 12.190 10.900 12.510 11.220 ;
        RECT 13.800 10.910 14.120 11.230 ;
        RECT 15.410 10.910 15.730 11.230 ;
        RECT 12.230 10.670 12.460 10.900 ;
        RECT 13.840 10.680 14.070 10.910 ;
        RECT 15.450 10.680 15.680 10.910 ;
        RECT 16.650 10.750 16.970 11.070 ;
        RECT 17.320 10.750 17.640 11.070 ;
        RECT 7.310 10.490 7.630 10.540 ;
        RECT 4.030 9.550 4.350 9.870 ;
        RECT 4.070 9.320 4.300 9.550 ;
        RECT 4.050 8.600 4.370 8.920 ;
        RECT 10.560 8.890 14.010 8.970 ;
        RECT 10.540 8.800 14.010 8.890 ;
        RECT 10.540 8.670 10.760 8.800 ;
        RECT 4.090 8.370 4.320 8.600 ;
        RECT 10.530 8.380 10.760 8.670 ;
        RECT 4.050 7.660 4.370 7.980 ;
        RECT 4.090 7.430 4.320 7.660 ;
        RECT 12.110 7.550 12.340 8.060 ;
        RECT 12.110 6.290 12.290 7.550 ;
        RECT 13.810 6.980 14.010 8.800 ;
        RECT 13.760 6.960 14.010 6.980 ;
        RECT 13.760 6.760 13.980 6.960 ;
        RECT 13.750 6.470 13.980 6.760 ;
        RECT 12.110 5.970 12.370 6.290 ;
      LAYER via ;
        RECT 4.080 10.890 4.340 11.150 ;
        RECT 5.790 10.930 6.050 11.190 ;
        RECT 8.990 10.930 9.250 11.190 ;
        RECT 10.600 10.940 10.860 11.200 ;
        RECT 12.220 10.930 12.480 11.190 ;
        RECT 7.340 10.520 7.600 10.780 ;
        RECT 13.830 10.940 14.090 11.200 ;
        RECT 15.440 10.940 15.700 11.200 ;
        RECT 16.680 10.780 16.940 11.040 ;
        RECT 17.350 10.780 17.610 11.040 ;
        RECT 4.060 9.580 4.320 9.840 ;
        RECT 4.080 8.630 4.340 8.890 ;
        RECT 4.080 7.690 4.340 7.950 ;
        RECT 12.110 6.000 12.370 6.260 ;
      LAYER met2 ;
        RECT 4.050 8.600 4.370 8.920 ;
        RECT 4.050 7.660 4.370 7.980 ;
  END
END sky130_hilas_DAC5bit01

MACRO sky130_hilas_VinjNOR3
  CLASS BLOCK ;
  FOREIGN sky130_hilas_VinjNOR3 ;
  ORIGIN 3.370 -1.440 ;
  SIZE 6.880 BY 1.640 ;
  OBS
      LAYER nwell ;
        RECT -3.360 1.440 0.080 3.080 ;
      LAYER li1 ;
        RECT -2.740 2.650 -2.570 2.790 ;
        RECT -2.010 2.670 -1.840 2.750 ;
        RECT -1.200 2.670 -1.030 2.750 ;
        RECT 0.340 2.710 0.510 2.830 ;
        RECT -2.740 2.480 -2.550 2.650 ;
        RECT -2.740 2.380 -2.570 2.480 ;
        RECT -2.010 2.100 -1.800 2.670 ;
        RECT -1.240 2.420 -1.030 2.670 ;
        RECT -0.640 2.490 -0.470 2.590 ;
        RECT 0.300 2.540 0.510 2.710 ;
        RECT 2.230 2.640 2.490 2.710 ;
        RECT 3.030 2.640 3.210 2.770 ;
        RECT 0.340 2.500 0.510 2.540 ;
        RECT -1.240 2.100 -1.070 2.420 ;
        RECT -0.670 2.320 -0.470 2.490 ;
        RECT -0.640 2.220 -0.470 2.320 ;
        RECT 0.900 2.460 1.770 2.630 ;
        RECT 2.230 2.460 3.210 2.640 ;
        RECT -3.170 2.000 -3.000 2.100 ;
        RECT -3.190 1.830 -3.000 2.000 ;
        RECT -3.170 1.770 -3.000 1.830 ;
        RECT -2.750 2.040 -2.580 2.100 ;
        RECT -2.750 1.770 -2.500 2.040 ;
        RECT -2.010 1.850 -1.760 2.100 ;
        RECT -2.740 1.750 -2.500 1.770 ;
        RECT -1.930 1.760 -1.760 1.850 ;
        RECT -1.280 1.850 -1.070 2.100 ;
        RECT 0.900 2.020 1.070 2.460 ;
        RECT 2.230 2.020 2.490 2.460 ;
        RECT 3.030 2.350 3.210 2.460 ;
        RECT -0.560 1.850 1.070 2.020 ;
        RECT 1.520 1.850 2.490 2.020 ;
        RECT 2.940 1.850 3.280 2.020 ;
        RECT -1.280 1.770 -1.110 1.850 ;
        RECT 0.210 1.810 0.380 1.850 ;
      LAYER mcon ;
        RECT -2.720 2.480 -2.550 2.650 ;
        RECT -2.710 1.800 -2.540 1.970 ;
        RECT 2.260 2.140 2.440 2.320 ;
      LAYER met1 ;
        RECT -2.750 2.700 -2.530 3.040 ;
        RECT -2.750 2.440 -2.520 2.700 ;
        RECT -3.280 1.760 -2.970 2.110 ;
        RECT -2.750 2.040 -2.530 2.440 ;
        RECT -0.730 2.280 -0.400 2.540 ;
        RECT 0.240 2.500 0.670 2.790 ;
        RECT -2.750 1.730 -2.500 2.040 ;
        RECT 0.110 1.750 0.500 2.020 ;
        RECT -2.750 1.530 -2.530 1.730 ;
        RECT 2.220 1.530 2.490 3.050 ;
        RECT 3.040 1.760 3.350 2.080 ;
      LAYER via ;
        RECT -3.250 1.790 -2.990 2.050 ;
        RECT -0.690 2.280 -0.430 2.540 ;
        RECT 0.300 2.530 0.560 2.790 ;
        RECT 0.170 1.750 0.430 2.010 ;
        RECT 3.070 1.790 3.330 2.050 ;
      LAYER met2 ;
        RECT -3.370 2.730 0.670 2.890 ;
        RECT -0.730 2.460 -0.400 2.540 ;
        RECT 0.250 2.500 0.670 2.730 ;
        RECT -1.000 2.440 -0.400 2.460 ;
        RECT -3.360 2.280 -0.400 2.440 ;
        RECT -3.280 1.950 -2.960 2.050 ;
        RECT -3.360 1.790 -2.960 1.950 ;
        RECT 0.130 1.930 0.500 2.010 ;
        RECT 0.130 1.920 1.160 1.930 ;
        RECT 3.040 1.920 3.350 2.080 ;
        RECT 0.130 1.750 3.510 1.920 ;
  END
END sky130_hilas_VinjNOR3

MACRO sky130_hilas_VinjDecode2to4
  CLASS BLOCK ;
  FOREIGN sky130_hilas_VinjDecode2to4 ;
  ORIGIN 6.370 -0.540 ;
  SIZE 12.950 BY 6.160 ;
  PIN OUTPUT00
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 3.200 5.550 3.570 5.630 ;
        RECT 3.200 5.540 4.230 5.550 ;
        RECT 6.110 5.540 6.420 5.700 ;
        RECT 3.200 5.370 6.580 5.540 ;
    END
  END OUTPUT00
  PIN OUTPUT01
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 3.200 4.040 3.570 4.120 ;
        RECT 3.200 4.030 4.230 4.040 ;
        RECT 6.110 4.030 6.420 4.190 ;
        RECT 3.200 3.860 6.580 4.030 ;
    END
  END OUTPUT01
  PIN OUTPUT10
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 3.200 2.530 3.570 2.610 ;
        RECT 3.200 2.520 4.230 2.530 ;
        RECT 6.110 2.520 6.420 2.680 ;
        RECT 3.200 2.350 6.580 2.520 ;
    END
  END OUTPUT10
  PIN OUTPUT11
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 3.200 1.030 3.570 1.110 ;
        RECT 3.200 1.020 4.230 1.030 ;
        RECT 6.110 1.020 6.420 1.180 ;
        RECT 3.200 0.850 6.580 1.020 ;
    END
  END OUTPUT11
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 5.290 0.630 5.560 6.670 ;
    END
    PORT
      LAYER met1 ;
        RECT -3.190 2.130 -2.960 6.660 ;
    END
  END VGND
  PIN VINJ
    ANTENNADIFFAREA 0.914000 ;
    PORT
      LAYER nwell ;
        RECT -0.290 0.540 3.150 6.700 ;
      LAYER met1 ;
        RECT 0.320 6.320 0.540 6.660 ;
        RECT 0.320 6.060 0.550 6.320 ;
        RECT 0.320 5.660 0.540 6.060 ;
        RECT 0.320 5.350 0.570 5.660 ;
        RECT 0.320 4.810 0.540 5.350 ;
        RECT 0.320 4.550 0.550 4.810 ;
        RECT 0.320 4.150 0.540 4.550 ;
        RECT 0.320 3.840 0.570 4.150 ;
        RECT 0.320 3.300 0.540 3.840 ;
        RECT 0.320 3.040 0.550 3.300 ;
        RECT 0.320 2.640 0.540 3.040 ;
        RECT 0.320 2.330 0.570 2.640 ;
        RECT 0.320 1.800 0.540 2.330 ;
        RECT 0.320 1.540 0.550 1.800 ;
        RECT 0.320 1.140 0.540 1.540 ;
        RECT 0.320 0.830 0.570 1.140 ;
        RECT 0.320 0.630 0.540 0.830 ;
    END
    PORT
      LAYER nwell ;
        RECT -6.370 2.040 -4.390 6.700 ;
      LAYER met1 ;
        RECT -5.760 6.320 -5.540 6.660 ;
        RECT -5.760 6.060 -5.530 6.320 ;
        RECT -5.760 5.660 -5.540 6.060 ;
        RECT -5.760 5.350 -5.510 5.660 ;
        RECT -5.760 4.810 -5.540 5.350 ;
        RECT -5.760 4.550 -5.530 4.810 ;
        RECT -5.760 4.150 -5.540 4.550 ;
        RECT -5.760 3.840 -5.510 4.150 ;
        RECT -5.760 3.300 -5.540 3.840 ;
        RECT -5.760 3.040 -5.530 3.300 ;
        RECT -5.760 2.640 -5.540 3.040 ;
        RECT -5.760 2.330 -5.510 2.640 ;
        RECT -5.760 2.130 -5.540 2.330 ;
    END
  END VINJ
  PIN IN2
    ANTENNAGATEAREA 0.642800 ;
    PORT
      LAYER met2 ;
        RECT -1.810 6.060 -1.480 6.120 ;
        RECT 2.340 6.080 2.670 6.160 ;
        RECT 2.070 6.060 2.670 6.080 ;
        RECT -1.810 5.900 2.670 6.060 ;
        RECT -1.810 5.850 -1.480 5.900 ;
        RECT -6.370 4.740 -1.580 4.760 ;
        RECT -6.370 4.580 -1.530 4.740 ;
        RECT -1.800 4.550 -1.530 4.580 ;
        RECT -1.800 4.410 -1.520 4.550 ;
        RECT -1.750 4.390 -1.520 4.410 ;
        RECT -1.830 3.040 -1.500 3.100 ;
        RECT 2.340 3.060 2.670 3.140 ;
        RECT 2.070 3.040 2.670 3.060 ;
        RECT -1.830 2.880 2.670 3.040 ;
        RECT -1.830 2.830 -1.500 2.880 ;
    END
  END IN2
  PIN IN1
    ANTENNAGATEAREA 0.673600 ;
    PORT
      LAYER met2 ;
        RECT -2.660 6.500 3.740 6.510 ;
        RECT -2.680 6.350 3.740 6.500 ;
        RECT -2.680 6.340 -2.410 6.350 ;
        RECT -2.710 6.270 -2.410 6.340 ;
        RECT -6.370 6.090 -2.410 6.270 ;
        RECT 3.320 6.120 3.740 6.350 ;
        RECT -2.710 6.010 -2.440 6.090 ;
        RECT -2.740 5.170 -2.410 5.230 ;
        RECT -2.740 5.010 -1.100 5.170 ;
        RECT -2.740 4.960 -2.410 5.010 ;
        RECT -1.260 5.000 -1.100 5.010 ;
        RECT -1.260 4.840 3.740 5.000 ;
        RECT 3.320 4.610 3.740 4.840 ;
    END
  END IN1
  PIN ENABLE
    PORT
      LAYER met2 ;
        RECT -6.370 3.070 -2.760 3.250 ;
    END
  END ENABLE
  OBS
      LAYER li1 ;
        RECT -5.750 6.270 -5.580 6.410 ;
        RECT 0.330 6.270 0.500 6.410 ;
        RECT 1.060 6.290 1.230 6.370 ;
        RECT 1.870 6.290 2.040 6.370 ;
        RECT 3.410 6.330 3.580 6.450 ;
        RECT -5.750 6.100 -5.560 6.270 ;
        RECT -5.750 6.000 -5.580 6.100 ;
        RECT -6.180 5.620 -6.010 5.720 ;
        RECT -6.200 5.450 -6.010 5.620 ;
        RECT -6.180 5.390 -6.010 5.450 ;
        RECT -5.760 5.660 -5.590 5.720 ;
        RECT -5.760 5.390 -5.510 5.660 ;
        RECT -5.020 5.640 -4.770 5.720 ;
        RECT -5.020 5.470 -3.720 5.640 ;
        RECT -3.160 5.630 -2.990 6.260 ;
        RECT 0.330 6.100 0.520 6.270 ;
        RECT 0.330 6.000 0.500 6.100 ;
        RECT 1.060 5.720 1.270 6.290 ;
        RECT 1.830 6.040 2.040 6.290 ;
        RECT 2.430 6.110 2.600 6.210 ;
        RECT 3.370 6.160 3.580 6.330 ;
        RECT 5.300 6.260 5.560 6.330 ;
        RECT 6.100 6.260 6.280 6.390 ;
        RECT 3.410 6.120 3.580 6.160 ;
        RECT 1.830 5.720 2.000 6.040 ;
        RECT 2.400 5.940 2.600 6.110 ;
        RECT 2.430 5.840 2.600 5.940 ;
        RECT 3.970 6.080 4.840 6.250 ;
        RECT 5.300 6.080 6.280 6.260 ;
        RECT -5.750 5.370 -5.510 5.390 ;
        RECT -4.940 5.380 -4.770 5.470 ;
        RECT -3.240 5.460 -2.910 5.630 ;
        RECT -0.100 5.620 0.070 5.720 ;
        RECT -0.120 5.450 0.070 5.620 ;
        RECT -0.100 5.390 0.070 5.450 ;
        RECT 0.320 5.660 0.490 5.720 ;
        RECT 0.320 5.390 0.570 5.660 ;
        RECT 1.060 5.470 1.310 5.720 ;
        RECT 0.330 5.370 0.570 5.390 ;
        RECT 1.140 5.380 1.310 5.470 ;
        RECT 1.790 5.470 2.000 5.720 ;
        RECT 3.970 5.640 4.140 6.080 ;
        RECT 5.300 5.640 5.560 6.080 ;
        RECT 6.100 5.970 6.280 6.080 ;
        RECT 2.510 5.470 4.140 5.640 ;
        RECT 4.590 5.470 5.560 5.640 ;
        RECT 6.010 5.470 6.350 5.640 ;
        RECT 1.790 5.390 1.960 5.470 ;
        RECT 3.280 5.430 3.450 5.470 ;
        RECT -5.750 4.760 -5.580 4.900 ;
        RECT 0.330 4.760 0.500 4.900 ;
        RECT 1.060 4.780 1.230 4.860 ;
        RECT 1.870 4.780 2.040 4.860 ;
        RECT 3.410 4.820 3.580 4.940 ;
        RECT -5.750 4.590 -5.560 4.760 ;
        RECT -5.750 4.490 -5.580 4.590 ;
        RECT -6.180 4.110 -6.010 4.210 ;
        RECT -6.200 3.940 -6.010 4.110 ;
        RECT -6.180 3.880 -6.010 3.940 ;
        RECT -5.760 4.150 -5.590 4.210 ;
        RECT -5.760 3.880 -5.510 4.150 ;
        RECT -5.020 4.130 -4.770 4.210 ;
        RECT -5.020 3.960 -3.720 4.130 ;
        RECT -3.160 4.120 -2.990 4.750 ;
        RECT 0.330 4.590 0.520 4.760 ;
        RECT 0.330 4.490 0.500 4.590 ;
        RECT 1.060 4.210 1.270 4.780 ;
        RECT 1.830 4.530 2.040 4.780 ;
        RECT 2.430 4.600 2.600 4.700 ;
        RECT 3.370 4.650 3.580 4.820 ;
        RECT 5.300 4.750 5.560 4.820 ;
        RECT 6.100 4.750 6.280 4.880 ;
        RECT 3.410 4.610 3.580 4.650 ;
        RECT 1.830 4.210 2.000 4.530 ;
        RECT 2.400 4.430 2.600 4.600 ;
        RECT 2.430 4.330 2.600 4.430 ;
        RECT 3.970 4.570 4.840 4.740 ;
        RECT 5.300 4.570 6.280 4.750 ;
        RECT -5.750 3.860 -5.510 3.880 ;
        RECT -4.940 3.870 -4.770 3.960 ;
        RECT -3.240 3.950 -2.910 4.120 ;
        RECT -0.100 4.110 0.070 4.210 ;
        RECT -0.120 3.940 0.070 4.110 ;
        RECT -0.100 3.880 0.070 3.940 ;
        RECT 0.320 4.150 0.490 4.210 ;
        RECT 0.320 3.880 0.570 4.150 ;
        RECT 1.060 3.960 1.310 4.210 ;
        RECT 0.330 3.860 0.570 3.880 ;
        RECT 1.140 3.870 1.310 3.960 ;
        RECT 1.790 3.960 2.000 4.210 ;
        RECT 3.970 4.130 4.140 4.570 ;
        RECT 5.300 4.130 5.560 4.570 ;
        RECT 6.100 4.460 6.280 4.570 ;
        RECT 2.510 3.960 4.140 4.130 ;
        RECT 4.590 3.960 5.560 4.130 ;
        RECT 6.010 3.960 6.350 4.130 ;
        RECT 1.790 3.880 1.960 3.960 ;
        RECT 3.280 3.920 3.450 3.960 ;
        RECT -5.750 3.250 -5.580 3.390 ;
        RECT 0.330 3.250 0.500 3.390 ;
        RECT 1.060 3.270 1.230 3.350 ;
        RECT 1.870 3.270 2.040 3.350 ;
        RECT 3.410 3.310 3.580 3.430 ;
        RECT -5.750 3.080 -5.560 3.250 ;
        RECT -5.750 2.980 -5.580 3.080 ;
        RECT -6.180 2.600 -6.010 2.700 ;
        RECT -6.200 2.430 -6.010 2.600 ;
        RECT -6.180 2.370 -6.010 2.430 ;
        RECT -5.760 2.640 -5.590 2.700 ;
        RECT -5.760 2.370 -5.510 2.640 ;
        RECT -5.020 2.620 -4.770 2.700 ;
        RECT -5.020 2.450 -3.720 2.620 ;
        RECT -3.160 2.610 -2.990 3.240 ;
        RECT 0.330 3.080 0.520 3.250 ;
        RECT 0.330 2.980 0.500 3.080 ;
        RECT 1.060 2.700 1.270 3.270 ;
        RECT 1.830 3.020 2.040 3.270 ;
        RECT 2.430 3.090 2.600 3.190 ;
        RECT 3.370 3.140 3.580 3.310 ;
        RECT 5.300 3.240 5.560 3.310 ;
        RECT 6.100 3.240 6.280 3.370 ;
        RECT 3.410 3.100 3.580 3.140 ;
        RECT 1.830 2.700 2.000 3.020 ;
        RECT 2.400 2.920 2.600 3.090 ;
        RECT 2.430 2.820 2.600 2.920 ;
        RECT 3.970 3.060 4.840 3.230 ;
        RECT 5.300 3.060 6.280 3.240 ;
        RECT -5.750 2.350 -5.510 2.370 ;
        RECT -4.940 2.360 -4.770 2.450 ;
        RECT -3.240 2.440 -2.910 2.610 ;
        RECT -0.100 2.600 0.070 2.700 ;
        RECT -0.120 2.430 0.070 2.600 ;
        RECT -0.100 2.370 0.070 2.430 ;
        RECT 0.320 2.640 0.490 2.700 ;
        RECT 0.320 2.370 0.570 2.640 ;
        RECT 1.060 2.450 1.310 2.700 ;
        RECT 0.330 2.350 0.570 2.370 ;
        RECT 1.140 2.360 1.310 2.450 ;
        RECT 1.790 2.450 2.000 2.700 ;
        RECT 3.970 2.620 4.140 3.060 ;
        RECT 5.300 2.620 5.560 3.060 ;
        RECT 6.100 2.950 6.280 3.060 ;
        RECT 2.510 2.450 4.140 2.620 ;
        RECT 4.590 2.450 5.560 2.620 ;
        RECT 6.010 2.450 6.350 2.620 ;
        RECT 1.790 2.370 1.960 2.450 ;
        RECT 3.280 2.410 3.450 2.450 ;
        RECT 0.330 1.750 0.500 1.890 ;
        RECT 1.060 1.770 1.230 1.850 ;
        RECT 1.870 1.770 2.040 1.850 ;
        RECT 3.410 1.810 3.580 1.930 ;
        RECT 0.330 1.580 0.520 1.750 ;
        RECT 0.330 1.480 0.500 1.580 ;
        RECT 1.060 1.200 1.270 1.770 ;
        RECT 1.830 1.520 2.040 1.770 ;
        RECT 2.430 1.590 2.600 1.690 ;
        RECT 3.370 1.640 3.580 1.810 ;
        RECT 5.300 1.740 5.560 1.810 ;
        RECT 6.100 1.740 6.280 1.870 ;
        RECT 3.410 1.600 3.580 1.640 ;
        RECT 1.830 1.200 2.000 1.520 ;
        RECT 2.400 1.420 2.600 1.590 ;
        RECT 2.430 1.320 2.600 1.420 ;
        RECT 3.970 1.560 4.840 1.730 ;
        RECT 5.300 1.560 6.280 1.740 ;
        RECT -0.100 1.100 0.070 1.200 ;
        RECT -0.120 0.930 0.070 1.100 ;
        RECT -0.100 0.870 0.070 0.930 ;
        RECT 0.320 1.140 0.490 1.200 ;
        RECT 0.320 0.870 0.570 1.140 ;
        RECT 1.060 0.950 1.310 1.200 ;
        RECT 0.330 0.850 0.570 0.870 ;
        RECT 1.140 0.860 1.310 0.950 ;
        RECT 1.790 0.950 2.000 1.200 ;
        RECT 3.970 1.120 4.140 1.560 ;
        RECT 5.300 1.120 5.560 1.560 ;
        RECT 6.100 1.450 6.280 1.560 ;
        RECT 2.510 0.950 4.140 1.120 ;
        RECT 4.590 0.950 5.560 1.120 ;
        RECT 6.010 0.950 6.350 1.120 ;
        RECT 1.790 0.870 1.960 0.950 ;
        RECT 3.280 0.910 3.450 0.950 ;
      LAYER mcon ;
        RECT -5.730 6.100 -5.560 6.270 ;
        RECT 0.350 6.100 0.520 6.270 ;
        RECT -3.160 5.740 -2.990 5.910 ;
        RECT -5.720 5.420 -5.550 5.590 ;
        RECT -4.380 5.470 -4.210 5.640 ;
        RECT 0.360 5.420 0.530 5.590 ;
        RECT 5.330 5.760 5.510 5.940 ;
        RECT -5.730 4.590 -5.560 4.760 ;
        RECT 0.350 4.590 0.520 4.760 ;
        RECT -3.160 4.230 -2.990 4.400 ;
        RECT -5.720 3.910 -5.550 4.080 ;
        RECT -4.380 3.960 -4.210 4.130 ;
        RECT 0.360 3.910 0.530 4.080 ;
        RECT 5.330 4.250 5.510 4.430 ;
        RECT -5.730 3.080 -5.560 3.250 ;
        RECT 0.350 3.080 0.520 3.250 ;
        RECT -3.160 2.720 -2.990 2.890 ;
        RECT -5.720 2.400 -5.550 2.570 ;
        RECT -4.380 2.450 -4.210 2.620 ;
        RECT 0.360 2.400 0.530 2.570 ;
        RECT 5.330 2.740 5.510 2.920 ;
        RECT 0.350 1.580 0.520 1.750 ;
        RECT 0.360 0.900 0.530 1.070 ;
        RECT 5.330 1.240 5.510 1.420 ;
      LAYER met1 ;
        RECT -2.700 6.310 -2.430 6.600 ;
        RECT -2.740 6.040 -2.410 6.310 ;
        RECT -6.290 5.380 -5.980 5.730 ;
        RECT -4.460 5.420 -4.140 5.680 ;
        RECT -2.700 5.260 -2.430 6.040 ;
        RECT -2.710 4.930 -2.430 5.260 ;
        RECT -2.700 4.900 -2.430 4.930 ;
        RECT -6.290 3.870 -5.980 4.220 ;
        RECT -4.460 3.910 -4.140 4.170 ;
        RECT -2.240 3.580 -1.970 5.700 ;
        RECT -1.780 4.710 -1.510 6.170 ;
        RECT 2.340 5.900 2.670 6.160 ;
        RECT 3.310 6.120 3.740 6.410 ;
        RECT -0.830 5.670 -0.540 5.720 ;
        RECT -0.850 5.320 -0.540 5.670 ;
        RECT -0.210 5.380 0.100 5.730 ;
        RECT 3.180 5.370 3.570 5.640 ;
        RECT 6.110 5.380 6.420 5.700 ;
        RECT -1.830 4.440 -1.500 4.710 ;
        RECT -2.250 3.250 -1.970 3.580 ;
        RECT -6.290 2.360 -5.980 2.710 ;
        RECT -4.460 2.400 -4.140 2.660 ;
        RECT -2.240 2.080 -1.970 3.250 ;
        RECT -1.780 3.130 -1.510 4.440 ;
        RECT -1.800 2.800 -1.510 3.130 ;
        RECT -1.780 2.780 -1.510 2.800 ;
        RECT -1.310 4.170 -1.040 4.230 ;
        RECT -1.310 3.840 -1.030 4.170 ;
        RECT -2.240 1.750 -1.940 2.080 ;
        RECT -2.240 1.700 -1.970 1.750 ;
        RECT -1.310 1.630 -1.040 3.840 ;
        RECT -1.330 1.300 -1.040 1.630 ;
        RECT -1.310 1.270 -1.040 1.300 ;
        RECT -0.830 2.670 -0.540 5.320 ;
        RECT 2.340 4.390 2.670 4.650 ;
        RECT 3.310 4.610 3.740 4.900 ;
        RECT -0.210 3.870 0.100 4.220 ;
        RECT 3.180 3.860 3.570 4.130 ;
        RECT 6.110 3.870 6.420 4.190 ;
        RECT 2.340 2.880 2.670 3.140 ;
        RECT 3.310 3.100 3.740 3.390 ;
        RECT -0.830 2.320 -0.530 2.670 ;
        RECT -0.210 2.360 0.100 2.710 ;
        RECT 3.180 2.350 3.570 2.620 ;
        RECT 6.110 2.360 6.420 2.680 ;
        RECT -0.830 0.780 -0.540 2.320 ;
        RECT 2.340 1.380 2.670 1.640 ;
        RECT 3.310 1.600 3.740 1.890 ;
        RECT -0.210 0.860 0.100 1.210 ;
        RECT 3.180 0.850 3.570 1.120 ;
        RECT 6.110 0.860 6.420 1.180 ;
      LAYER via ;
        RECT -2.710 6.040 -2.440 6.310 ;
        RECT -6.260 5.410 -6.000 5.670 ;
        RECT -4.430 5.420 -4.170 5.680 ;
        RECT -1.780 5.850 -1.510 6.120 ;
        RECT 2.380 5.900 2.640 6.160 ;
        RECT 3.370 6.150 3.630 6.410 ;
        RECT -2.710 4.960 -2.440 5.230 ;
        RECT -2.240 5.360 -1.970 5.630 ;
        RECT -6.260 3.900 -6.000 4.160 ;
        RECT -4.430 3.910 -4.170 4.170 ;
        RECT -0.850 5.350 -0.560 5.640 ;
        RECT -0.180 5.410 0.080 5.670 ;
        RECT 3.240 5.370 3.500 5.630 ;
        RECT 6.140 5.410 6.400 5.670 ;
        RECT -1.800 4.440 -1.530 4.710 ;
        RECT -2.250 3.280 -1.980 3.550 ;
        RECT -6.260 2.390 -6.000 2.650 ;
        RECT -4.430 2.400 -4.170 2.660 ;
        RECT -1.800 2.830 -1.530 3.100 ;
        RECT -1.300 3.870 -1.030 4.140 ;
        RECT 2.380 4.390 2.640 4.650 ;
        RECT 3.370 4.640 3.630 4.900 ;
        RECT -0.810 3.840 -0.550 4.100 ;
        RECT -0.180 3.900 0.080 4.160 ;
        RECT 3.240 3.860 3.500 4.120 ;
        RECT 6.140 3.900 6.400 4.160 ;
        RECT -2.210 1.780 -1.940 2.050 ;
        RECT -1.330 1.330 -1.060 1.600 ;
        RECT 2.380 2.880 2.640 3.140 ;
        RECT 3.370 3.130 3.630 3.390 ;
        RECT -0.820 2.350 -0.530 2.640 ;
        RECT -0.180 2.390 0.080 2.650 ;
        RECT 3.240 2.350 3.500 2.610 ;
        RECT 6.140 2.390 6.400 2.650 ;
        RECT 2.380 1.380 2.640 1.640 ;
        RECT 3.370 1.630 3.630 1.890 ;
        RECT -0.830 0.810 -0.540 1.100 ;
        RECT -0.180 0.890 0.080 1.150 ;
        RECT 3.240 0.850 3.500 1.110 ;
        RECT 6.140 0.890 6.400 1.150 ;
      LAYER met2 ;
        RECT -6.290 5.570 -5.970 5.670 ;
        RECT -6.300 5.410 -5.970 5.570 ;
        RECT -4.460 5.600 -4.140 5.680 ;
        RECT -2.270 5.600 -1.940 5.630 ;
        RECT -4.460 5.420 -1.920 5.600 ;
        RECT -2.270 5.410 -1.920 5.420 ;
        RECT -0.880 5.570 -0.530 5.640 ;
        RECT -0.210 5.570 0.110 5.670 ;
        RECT -0.880 5.410 0.110 5.570 ;
        RECT -2.270 5.360 -1.940 5.410 ;
        RECT -0.880 5.350 -0.530 5.410 ;
        RECT 2.340 4.570 2.670 4.650 ;
        RECT 2.070 4.550 2.670 4.570 ;
        RECT -1.250 4.390 2.670 4.550 ;
        RECT -6.290 4.060 -5.970 4.160 ;
        RECT -6.300 3.900 -5.970 4.060 ;
        RECT -4.460 4.090 -4.140 4.170 ;
        RECT -1.250 4.140 -1.090 4.390 ;
        RECT -1.330 4.090 -1.000 4.140 ;
        RECT -4.460 3.910 -1.000 4.090 ;
        RECT -1.330 3.870 -1.000 3.910 ;
        RECT -0.840 4.060 -0.520 4.100 ;
        RECT -0.210 4.060 0.110 4.160 ;
        RECT -0.840 3.900 0.110 4.060 ;
        RECT -0.840 3.840 -0.520 3.900 ;
        RECT -2.280 3.490 -1.950 3.550 ;
        RECT -2.280 3.330 3.740 3.490 ;
        RECT -2.280 3.280 -1.950 3.330 ;
        RECT 3.320 3.100 3.740 3.330 ;
        RECT -6.290 2.550 -5.970 2.650 ;
        RECT -6.300 2.390 -5.970 2.550 ;
        RECT -4.460 2.580 -4.140 2.660 ;
        RECT -0.850 2.580 -0.500 2.640 ;
        RECT -4.460 2.550 -0.360 2.580 ;
        RECT -0.210 2.550 0.110 2.650 ;
        RECT -4.460 2.400 0.110 2.550 ;
        RECT -0.850 2.390 0.110 2.400 ;
        RECT -0.850 2.350 -0.500 2.390 ;
        RECT -2.240 1.990 -1.910 2.050 ;
        RECT -2.240 1.830 3.740 1.990 ;
        RECT -2.240 1.780 -1.910 1.830 ;
        RECT -1.360 1.540 -1.030 1.600 ;
        RECT 2.340 1.560 2.670 1.640 ;
        RECT 3.320 1.600 3.740 1.830 ;
        RECT 2.070 1.540 2.670 1.560 ;
        RECT -1.360 1.380 2.670 1.540 ;
        RECT -1.360 1.330 -1.030 1.380 ;
        RECT -0.860 1.050 -0.510 1.100 ;
        RECT -0.210 1.050 0.110 1.150 ;
        RECT -0.860 0.890 0.110 1.050 ;
        RECT -0.860 0.810 -0.510 0.890 ;
  END
END sky130_hilas_VinjDecode2to4

MACRO sky130_hilas_capacitorSize04
  CLASS BLOCK ;
  FOREIGN sky130_hilas_capacitorSize04 ;
  ORIGIN -14.150 0.180 ;
  SIZE 5.780 BY 5.290 ;
  PIN CAP1TERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 19.110 3.650 19.770 4.310 ;
    END
  END CAP1TERM02
  PIN CAP2TERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 19.110 0.650 19.770 1.310 ;
    END
  END CAP2TERM02
  PIN CAP2TERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 14.270 1.050 14.930 1.310 ;
        RECT 16.710 1.050 17.160 1.060 ;
        RECT 14.270 0.650 17.210 1.050 ;
        RECT 14.720 0.640 17.210 0.650 ;
        RECT 16.690 0.560 17.210 0.640 ;
    END
  END CAP2TERM01
  PIN CAP1TERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 14.240 4.060 14.900 4.310 ;
        RECT 16.710 4.060 17.160 4.070 ;
        RECT 14.240 3.650 17.210 4.060 ;
        RECT 16.690 3.570 17.210 3.650 ;
    END
  END CAP1TERM01
  OBS
      LAYER met2 ;
        RECT 14.170 4.800 19.920 4.980 ;
        RECT 14.170 4.370 19.920 4.550 ;
        RECT 14.370 4.130 14.740 4.190 ;
        RECT 14.170 3.850 14.740 4.130 ;
        RECT 14.370 3.790 14.740 3.850 ;
        RECT 19.240 4.130 19.610 4.190 ;
        RECT 19.240 3.850 19.920 4.130 ;
        RECT 19.240 3.790 19.610 3.850 ;
        RECT 14.170 3.370 19.920 3.550 ;
        RECT 14.170 2.940 19.920 3.120 ;
        RECT 14.170 1.790 19.920 1.960 ;
        RECT 14.170 1.370 19.920 1.540 ;
        RECT 14.400 1.130 14.770 1.190 ;
        RECT 14.170 0.850 14.770 1.130 ;
        RECT 14.400 0.790 14.770 0.850 ;
        RECT 19.240 1.130 19.610 1.190 ;
        RECT 19.240 0.850 19.930 1.130 ;
        RECT 19.240 0.790 19.610 0.850 ;
        RECT 14.170 0.390 19.920 0.560 ;
        RECT 14.170 -0.050 19.920 0.120 ;
      LAYER via2 ;
        RECT 14.420 3.850 14.700 4.130 ;
        RECT 19.290 3.850 19.570 4.130 ;
        RECT 14.450 0.850 14.730 1.130 ;
        RECT 19.290 0.850 19.570 1.130 ;
      LAYER met3 ;
        RECT 15.860 4.340 18.160 5.110 ;
        RECT 14.150 3.590 14.940 4.340 ;
        RECT 15.860 3.590 19.810 4.340 ;
        RECT 15.860 2.830 18.160 3.590 ;
        RECT 14.180 0.590 14.970 1.340 ;
        RECT 15.860 1.330 18.160 2.100 ;
        RECT 19.020 1.330 19.810 1.340 ;
        RECT 15.860 0.600 19.810 1.330 ;
        RECT 15.860 -0.180 18.160 0.600 ;
        RECT 19.020 0.590 19.810 0.600 ;
      LAYER via3 ;
        RECT 14.340 3.740 14.770 4.220 ;
        RECT 19.210 3.740 19.640 4.220 ;
        RECT 14.370 0.740 14.800 1.220 ;
        RECT 19.210 0.740 19.640 1.220 ;
  END
END sky130_hilas_capacitorSize04

MACRO sky130_hilas_swc4x1cellOverlap2
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc4x1cellOverlap2 ;
  ORIGIN 1.910 3.870 ;
  SIZE 9.350 BY 6.160 ;
  OBS
      LAYER nwell ;
        RECT 4.880 2.230 7.440 2.290 ;
        RECT 0.880 -3.820 7.440 2.230 ;
        RECT 4.880 -3.870 7.440 -3.820 ;
      LAYER li1 ;
        RECT -0.850 1.020 -0.680 1.910 ;
        RECT 1.230 0.920 4.540 1.900 ;
        RECT 4.980 1.820 5.300 1.830 ;
        RECT 4.980 1.650 5.560 1.820 ;
        RECT 4.980 1.600 5.310 1.650 ;
        RECT 4.980 1.570 5.300 1.600 ;
        RECT 6.840 1.550 7.040 1.900 ;
        RECT 4.980 1.240 5.300 1.280 ;
        RECT 4.980 1.200 5.310 1.240 ;
        RECT 4.980 1.030 5.560 1.200 ;
        RECT 4.980 1.020 5.300 1.030 ;
        RECT 6.110 0.930 6.310 1.530 ;
        RECT 6.840 1.520 7.050 1.550 ;
        RECT 6.830 0.930 7.050 1.520 ;
        RECT -0.850 -0.500 -0.680 0.390 ;
        RECT 1.230 -0.550 4.540 0.430 ;
        RECT 4.980 0.390 5.300 0.400 ;
        RECT 4.980 0.220 5.560 0.390 ;
        RECT 4.980 0.180 5.310 0.220 ;
        RECT 4.980 0.140 5.300 0.180 ;
        RECT 6.110 -0.110 6.310 0.490 ;
        RECT 6.830 -0.100 7.050 0.490 ;
        RECT 6.840 -0.130 7.050 -0.100 ;
        RECT 4.980 -0.180 5.300 -0.150 ;
        RECT 4.980 -0.230 5.310 -0.180 ;
        RECT 4.980 -0.400 5.560 -0.230 ;
        RECT 4.980 -0.410 5.300 -0.400 ;
        RECT 6.840 -0.480 7.040 -0.130 ;
        RECT 6.230 -0.880 6.670 -0.710 ;
        RECT -0.850 -1.950 -0.680 -1.060 ;
        RECT 1.230 -2.020 4.540 -1.040 ;
        RECT 4.980 -1.190 5.300 -1.180 ;
        RECT 4.980 -1.360 5.560 -1.190 ;
        RECT 4.980 -1.410 5.310 -1.360 ;
        RECT 4.980 -1.440 5.300 -1.410 ;
        RECT 6.840 -1.460 7.040 -1.110 ;
        RECT 4.980 -1.770 5.300 -1.730 ;
        RECT 4.980 -1.810 5.310 -1.770 ;
        RECT 4.980 -1.980 5.560 -1.810 ;
        RECT 4.980 -1.990 5.300 -1.980 ;
        RECT 6.110 -2.080 6.310 -1.480 ;
        RECT 6.840 -1.490 7.050 -1.460 ;
        RECT 6.830 -2.080 7.050 -1.490 ;
        RECT -0.850 -3.490 -0.680 -2.600 ;
        RECT 1.230 -3.490 4.540 -2.510 ;
        RECT 4.980 -2.610 5.300 -2.600 ;
        RECT 4.980 -2.780 5.560 -2.610 ;
        RECT 4.980 -2.820 5.310 -2.780 ;
        RECT 4.980 -2.860 5.300 -2.820 ;
        RECT 6.110 -3.110 6.310 -2.510 ;
        RECT 6.830 -3.100 7.050 -2.510 ;
        RECT 6.840 -3.130 7.050 -3.100 ;
        RECT 4.980 -3.180 5.300 -3.150 ;
        RECT 4.980 -3.230 5.310 -3.180 ;
        RECT 4.980 -3.400 5.560 -3.230 ;
        RECT 4.980 -3.410 5.300 -3.400 ;
        RECT 6.840 -3.480 7.040 -3.130 ;
      LAYER mcon ;
        RECT -0.850 1.710 -0.680 1.880 ;
        RECT 2.800 1.670 2.970 1.840 ;
        RECT 5.040 1.610 5.210 1.780 ;
        RECT 6.120 1.320 6.290 1.490 ;
        RECT 2.800 0.980 2.970 1.150 ;
        RECT 5.040 1.060 5.210 1.230 ;
        RECT 6.850 1.350 7.020 1.520 ;
        RECT -0.850 0.190 -0.680 0.360 ;
        RECT 2.800 0.200 2.970 0.370 ;
        RECT 5.040 0.190 5.210 0.360 ;
        RECT 6.120 -0.070 6.290 0.100 ;
        RECT 6.850 -0.100 7.020 0.070 ;
        RECT 2.800 -0.490 2.970 -0.320 ;
        RECT 5.040 -0.360 5.210 -0.190 ;
        RECT 6.490 -0.880 6.670 -0.710 ;
        RECT -0.850 -1.260 -0.680 -1.090 ;
        RECT 2.800 -1.270 2.970 -1.100 ;
        RECT 5.040 -1.400 5.210 -1.230 ;
        RECT 6.120 -1.690 6.290 -1.520 ;
        RECT 2.800 -1.960 2.970 -1.790 ;
        RECT 5.040 -1.950 5.210 -1.780 ;
        RECT 6.850 -1.660 7.020 -1.490 ;
        RECT -0.850 -2.800 -0.680 -2.630 ;
        RECT 2.800 -2.740 2.970 -2.570 ;
        RECT 5.040 -2.810 5.210 -2.640 ;
        RECT 6.120 -3.070 6.290 -2.900 ;
        RECT 6.850 -3.100 7.020 -2.930 ;
        RECT 2.800 -3.430 2.970 -3.260 ;
        RECT 5.040 -3.360 5.210 -3.190 ;
      LAYER met1 ;
        RECT -0.900 -3.820 -0.630 2.230 ;
        RECT 2.760 1.260 3.000 1.900 ;
        RECT 4.970 1.540 5.290 1.860 ;
        RECT 6.110 1.550 6.270 2.280 ;
        RECT 6.110 1.530 6.310 1.550 ;
        RECT 2.770 1.000 3.000 1.260 ;
        RECT 2.770 0.780 3.010 1.000 ;
        RECT 4.970 0.990 5.290 1.310 ;
        RECT 6.090 1.290 6.320 1.530 ;
        RECT 6.110 1.240 6.320 1.290 ;
        RECT 6.480 1.240 6.670 2.230 ;
        RECT 6.920 1.580 7.080 2.280 ;
        RECT 2.760 -0.210 3.000 0.430 ;
        RECT 4.970 0.110 5.290 0.430 ;
        RECT 6.110 0.180 6.270 1.240 ;
        RECT 6.500 1.120 6.670 1.240 ;
        RECT 6.510 0.300 6.670 1.120 ;
        RECT 6.810 1.030 7.080 1.580 ;
        RECT 6.810 0.980 7.090 1.030 ;
        RECT 6.920 0.890 7.090 0.980 ;
        RECT 6.920 0.530 7.080 0.890 ;
        RECT 6.920 0.440 7.090 0.530 ;
        RECT 6.500 0.180 6.670 0.300 ;
        RECT 6.110 0.130 6.320 0.180 ;
        RECT 6.090 -0.110 6.320 0.130 ;
        RECT 2.770 -0.470 3.000 -0.210 ;
        RECT 4.970 -0.440 5.290 -0.120 ;
        RECT 6.110 -0.130 6.310 -0.110 ;
        RECT 2.770 -0.690 3.010 -0.470 ;
        RECT 2.760 -1.680 3.000 -1.040 ;
        RECT 4.970 -1.470 5.290 -1.150 ;
        RECT 6.110 -1.460 6.270 -0.130 ;
        RECT 6.480 -0.680 6.670 0.180 ;
        RECT 6.810 0.390 7.090 0.440 ;
        RECT 6.810 -0.160 7.080 0.390 ;
        RECT 6.460 -0.910 6.700 -0.680 ;
        RECT 6.110 -1.480 6.310 -1.460 ;
        RECT 2.770 -1.940 3.000 -1.680 ;
        RECT 2.770 -2.160 3.010 -1.940 ;
        RECT 4.970 -2.020 5.290 -1.700 ;
        RECT 6.090 -1.720 6.320 -1.480 ;
        RECT 6.110 -1.770 6.320 -1.720 ;
        RECT 6.480 -1.770 6.670 -0.910 ;
        RECT 6.920 -1.430 7.080 -0.160 ;
        RECT 2.760 -3.150 3.000 -2.510 ;
        RECT 4.970 -2.890 5.290 -2.570 ;
        RECT 6.110 -2.820 6.270 -1.770 ;
        RECT 6.500 -1.890 6.670 -1.770 ;
        RECT 6.510 -2.700 6.670 -1.890 ;
        RECT 6.810 -1.980 7.080 -1.430 ;
        RECT 6.810 -2.030 7.090 -1.980 ;
        RECT 6.920 -2.120 7.090 -2.030 ;
        RECT 6.920 -2.470 7.080 -2.120 ;
        RECT 6.920 -2.560 7.090 -2.470 ;
        RECT 6.500 -2.820 6.670 -2.700 ;
        RECT 6.110 -2.870 6.320 -2.820 ;
        RECT 6.090 -3.110 6.320 -2.870 ;
        RECT 2.770 -3.410 3.000 -3.150 ;
        RECT 2.770 -3.630 3.010 -3.410 ;
        RECT 4.970 -3.440 5.290 -3.120 ;
        RECT 6.110 -3.130 6.310 -3.110 ;
        RECT 6.110 -3.860 6.270 -3.130 ;
        RECT 6.480 -3.810 6.670 -2.820 ;
        RECT 6.810 -2.610 7.090 -2.560 ;
        RECT 6.810 -3.160 7.080 -2.610 ;
        RECT 6.920 -3.860 7.080 -3.160 ;
      LAYER via ;
        RECT 5.000 1.570 5.260 1.830 ;
        RECT 5.000 1.020 5.260 1.280 ;
        RECT 5.000 0.140 5.260 0.400 ;
        RECT 5.000 -0.410 5.260 -0.150 ;
        RECT 5.000 -1.440 5.260 -1.180 ;
        RECT 5.000 -1.990 5.260 -1.730 ;
        RECT 5.000 -2.860 5.260 -2.600 ;
        RECT 5.000 -3.410 5.260 -3.150 ;
      LAYER met2 ;
        RECT 4.970 1.730 5.280 1.870 ;
        RECT -1.910 1.550 7.440 1.730 ;
        RECT 4.970 1.540 5.280 1.550 ;
        RECT 4.970 1.300 5.280 1.320 ;
        RECT -1.910 1.120 7.440 1.300 ;
        RECT 4.970 0.990 5.280 1.120 ;
        RECT 4.970 0.300 5.280 0.430 ;
        RECT -1.910 0.120 7.440 0.300 ;
        RECT 4.970 0.100 5.280 0.120 ;
        RECT 4.970 -0.130 5.280 -0.120 ;
        RECT -1.910 -0.200 4.960 -0.130 ;
        RECT 4.970 -0.200 7.440 -0.130 ;
        RECT -1.910 -0.310 7.440 -0.200 ;
        RECT 4.970 -0.450 5.280 -0.310 ;
        RECT 4.970 -1.280 5.280 -1.140 ;
        RECT 4.970 -1.290 7.440 -1.280 ;
        RECT -1.910 -1.460 7.440 -1.290 ;
        RECT 4.970 -1.470 5.280 -1.460 ;
        RECT 4.970 -1.710 5.280 -1.690 ;
        RECT -1.910 -1.880 7.440 -1.710 ;
        RECT 4.880 -1.890 7.440 -1.880 ;
        RECT 4.970 -2.020 5.280 -1.890 ;
        RECT 4.970 -2.690 5.280 -2.570 ;
        RECT -1.910 -2.700 5.280 -2.690 ;
        RECT -1.910 -2.860 7.440 -2.700 ;
        RECT 4.880 -2.880 7.440 -2.860 ;
        RECT 4.970 -2.900 5.280 -2.880 ;
        RECT 4.970 -3.130 5.280 -3.120 ;
        RECT -1.910 -3.300 7.440 -3.130 ;
        RECT 4.970 -3.310 7.440 -3.300 ;
        RECT 4.970 -3.450 5.280 -3.310 ;
  END
END sky130_hilas_swc4x1cellOverlap2

MACRO sky130_hilas_TA2Cell_NoFG
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TA2Cell_NoFG ;
  ORIGIN 14.730 -1.350 ;
  SIZE 17.920 BY 6.150 ;
  PIN COLSEL1
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT -4.160 5.990 -3.970 7.450 ;
        RECT -4.160 5.960 -3.940 5.990 ;
        RECT -4.180 5.690 -3.930 5.960 ;
        RECT -4.170 5.680 -3.930 5.690 ;
        RECT -4.170 5.440 -3.940 5.680 ;
        RECT -4.130 3.410 -3.970 5.440 ;
        RECT -4.170 3.170 -3.940 3.410 ;
        RECT -4.170 3.160 -3.930 3.170 ;
        RECT -4.180 2.890 -3.930 3.160 ;
        RECT -4.160 2.860 -3.940 2.890 ;
        RECT -4.160 1.400 -3.970 2.860 ;
    END
  END COLSEL1
  PIN VIN12
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -2.260 1.670 -1.950 1.740 ;
        RECT -2.860 1.420 -1.950 1.670 ;
        RECT -2.260 1.410 -1.950 1.420 ;
    END
  END VIN12
  PIN VIN21
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -0.940 4.750 -0.630 4.790 ;
        RECT -1.030 4.740 -0.600 4.750 ;
        RECT -1.260 4.510 -0.160 4.740 ;
        RECT -0.940 4.460 -0.630 4.510 ;
    END
  END VIN21
  PIN VIN22
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -1.300 7.430 -1.050 7.440 ;
        RECT -0.700 7.430 -0.390 7.440 ;
        RECT -1.300 7.180 -0.390 7.430 ;
        RECT -0.700 7.110 -0.390 7.180 ;
    END
  END VIN22
  PIN OUTPUT1
    ANTENNADIFFAREA 0.308800 ;
    PORT
      LAYER met2 ;
        RECT 0.270 4.140 0.580 4.190 ;
        RECT 2.560 4.140 2.870 4.270 ;
        RECT 0.270 3.920 3.190 4.140 ;
        RECT 0.270 3.860 0.580 3.920 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    ANTENNADIFFAREA 0.308800 ;
    PORT
      LAYER met2 ;
        RECT 0.270 4.970 0.580 5.030 ;
        RECT 2.570 4.970 2.880 4.990 ;
        RECT 0.270 4.740 3.190 4.970 ;
        RECT 0.270 4.700 0.580 4.740 ;
        RECT 2.570 4.660 2.880 4.740 ;
    END
  END OUTPUT2
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 1.230 6.000 1.570 6.090 ;
        RECT -1.120 5.810 1.570 6.000 ;
        RECT -1.120 5.240 -0.930 5.810 ;
        RECT 1.230 5.760 1.570 5.810 ;
        RECT -11.910 5.050 -0.930 5.240 ;
        RECT -11.910 4.870 -11.720 5.050 ;
        RECT -11.930 3.880 -11.580 4.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.230 1.400 1.570 7.450 ;
      LAYER via ;
        RECT 1.270 5.790 1.530 6.050 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 1.920 7.270 3.190 7.450 ;
        RECT 1.910 1.400 3.190 7.270 ;
      LAYER met1 ;
        RECT 1.900 5.870 2.170 7.450 ;
        RECT 1.900 5.580 2.180 5.870 ;
        RECT 1.900 3.280 2.170 5.580 ;
        RECT 1.900 2.990 2.180 3.280 ;
        RECT 1.900 1.400 2.170 2.990 ;
    END
  END VPWR
  PIN DRAIN1
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT -5.680 6.950 -5.370 6.960 ;
        RECT -14.730 6.770 -3.200 6.950 ;
        RECT -5.680 6.630 -5.370 6.770 ;
    END
  END DRAIN1
  PIN DRAIN2
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT -5.680 2.080 -5.370 2.220 ;
        RECT -5.680 2.070 -3.200 2.080 ;
        RECT -14.730 1.920 -3.200 2.070 ;
        RECT -5.680 1.900 -3.200 1.920 ;
        RECT -5.680 1.890 -5.370 1.900 ;
    END
  END DRAIN2
  PIN VTUN
    ANTENNADIFFAREA 2.516100 ;
    PORT
      LAYER nwell ;
        RECT -14.720 6.700 -12.990 7.450 ;
        RECT -14.720 5.550 -12.980 6.700 ;
        RECT -14.710 3.310 -12.980 5.550 ;
        RECT -14.720 3.130 -12.980 3.310 ;
        RECT -14.720 1.410 -12.990 3.130 ;
      LAYER met1 ;
        RECT -14.380 1.400 -13.960 7.450 ;
    END
  END VTUN
  PIN GATE1
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT -10.960 5.060 -8.240 6.710 ;
        RECT -10.960 5.020 -8.250 5.060 ;
        RECT -10.960 3.690 -8.250 3.730 ;
        RECT -10.960 2.040 -8.240 3.690 ;
      LAYER met1 ;
        RECT -10.680 6.240 -10.450 7.450 ;
        RECT -10.680 5.450 -10.420 6.240 ;
        RECT -10.680 3.300 -10.450 5.450 ;
        RECT -10.680 2.510 -10.420 3.300 ;
        RECT -10.680 1.400 -10.450 2.510 ;
    END
  END GATE1
  PIN VINJ
    ANTENNADIFFAREA 1.574400 ;
    PORT
      LAYER nwell ;
        RECT -6.510 7.450 -3.200 7.500 ;
        RECT -6.510 7.440 -1.650 7.450 ;
        RECT -6.510 1.410 -0.090 7.440 ;
        RECT -6.510 1.350 -3.200 1.410 ;
        RECT -1.950 1.400 -0.090 1.410 ;
      LAYER met2 ;
        RECT -4.590 4.590 -4.270 4.850 ;
        RECT -4.550 4.570 -3.370 4.590 ;
        RECT -4.550 4.310 -3.330 4.570 ;
        RECT -4.550 4.250 -3.370 4.310 ;
        RECT -4.590 4.240 -3.370 4.250 ;
        RECT -4.590 3.990 -4.270 4.240 ;
    END
  END VINJ
  PIN VIN11
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -2.500 4.340 -2.190 4.390 ;
        RECT -2.820 4.110 -1.720 4.340 ;
        RECT -2.820 4.100 -2.160 4.110 ;
        RECT -2.500 4.060 -2.190 4.100 ;
    END
  END VIN11
  OBS
      LAYER li1 ;
        RECT -0.960 7.400 -0.790 7.450 ;
        RECT -0.960 7.140 -0.400 7.400 ;
        RECT 0.510 7.150 0.710 7.190 ;
        RECT -0.960 7.120 -0.790 7.140 ;
        RECT -5.610 6.870 -5.080 7.040 ;
        RECT -3.800 6.770 -3.600 7.120 ;
        RECT -3.800 6.740 -3.590 6.770 ;
        RECT -14.290 5.310 -13.740 5.740 ;
        RECT -10.660 5.500 -10.430 6.190 ;
        RECT -5.360 5.960 -5.190 6.480 ;
        RECT -5.520 5.700 -5.190 5.960 ;
        RECT -11.900 4.470 -11.440 4.880 ;
        RECT -5.360 4.790 -5.190 5.700 ;
        RECT -4.530 4.880 -4.360 6.490 ;
        RECT -3.810 6.160 -3.590 6.740 ;
        RECT -3.800 6.150 -3.590 6.160 ;
        RECT -4.160 5.980 -3.970 5.990 ;
        RECT -4.160 5.690 -3.960 5.980 ;
        RECT -4.170 5.360 -3.880 5.690 ;
        RECT -4.530 4.690 -4.350 4.880 ;
        RECT -11.900 4.290 -8.140 4.470 ;
        RECT -14.290 3.580 -13.740 4.010 ;
        RECT -11.900 3.870 -11.440 4.290 ;
        RECT -10.660 2.560 -10.430 3.290 ;
        RECT -5.360 3.200 -5.190 4.060 ;
        RECT -5.520 2.940 -5.190 3.200 ;
        RECT -5.360 2.370 -5.190 2.940 ;
        RECT -4.530 3.970 -4.350 4.160 ;
        RECT -4.530 2.360 -4.360 3.970 ;
        RECT -4.170 3.160 -3.880 3.490 ;
        RECT -4.160 2.870 -3.960 3.160 ;
        RECT -3.100 3.070 -2.920 6.980 ;
        RECT -2.290 5.190 -2.120 6.970 ;
        RECT -1.540 6.040 -1.360 6.970 ;
        RECT 0.280 6.890 0.710 7.150 ;
        RECT -0.810 6.710 -0.480 6.880 ;
        RECT 0.510 6.860 0.710 6.890 ;
        RECT -0.730 6.570 -0.480 6.710 ;
        RECT -0.730 6.310 -0.250 6.570 ;
        RECT 0.100 6.500 0.270 6.540 ;
        RECT 0.510 6.500 0.710 6.530 ;
        RECT -1.660 6.010 -1.340 6.040 ;
        RECT -1.660 5.820 -1.330 6.010 ;
        RECT -1.660 5.780 -1.340 5.820 ;
        RECT -2.370 5.130 -1.830 5.190 ;
        RECT -2.370 5.020 -1.820 5.130 ;
        RECT -2.010 4.900 -1.820 5.020 ;
        RECT -2.540 4.600 -2.370 4.760 ;
        RECT -2.540 4.430 -2.320 4.600 ;
        RECT -2.490 4.350 -2.320 4.430 ;
        RECT -2.490 4.310 -2.170 4.350 ;
        RECT -2.490 4.120 -2.160 4.310 ;
        RECT -2.490 4.090 -2.170 4.120 ;
        RECT -3.220 3.030 -2.900 3.070 ;
        RECT -4.160 2.860 -3.970 2.870 ;
        RECT -3.220 2.840 -2.890 3.030 ;
        RECT -3.220 2.810 -2.900 2.840 ;
        RECT -3.800 2.690 -3.590 2.700 ;
        RECT -3.810 2.110 -3.590 2.690 ;
        RECT -3.800 2.080 -3.590 2.110 ;
        RECT -5.610 1.810 -5.080 1.980 ;
        RECT -3.800 1.730 -3.600 2.080 ;
        RECT -3.100 1.880 -2.920 2.810 ;
        RECT -2.290 2.540 -2.120 3.920 ;
        RECT -2.290 2.280 -1.810 2.540 ;
        RECT -2.290 2.140 -2.040 2.280 ;
        RECT -2.370 1.970 -2.040 2.140 ;
        RECT -1.540 1.870 -1.360 5.780 ;
        RECT -0.730 4.930 -0.560 6.310 ;
        RECT 0.100 6.240 0.710 6.500 ;
        RECT 0.100 6.210 0.270 6.240 ;
        RECT 0.510 6.200 0.710 6.240 ;
        RECT 1.100 6.200 1.650 7.190 ;
        RECT 2.470 7.040 3.100 7.210 ;
        RECT 2.470 6.940 2.860 7.040 ;
        RECT 2.470 6.910 2.850 6.940 ;
        RECT 2.470 6.760 2.830 6.910 ;
        RECT 2.120 6.590 2.830 6.760 ;
        RECT 2.120 5.840 2.820 6.150 ;
        RECT 0.100 5.650 0.270 5.680 ;
        RECT 0.510 5.650 0.710 5.690 ;
        RECT 0.100 5.390 0.710 5.650 ;
        RECT 0.100 5.350 0.270 5.390 ;
        RECT 0.510 5.360 0.710 5.390 ;
        RECT 0.510 5.000 0.710 5.030 ;
        RECT -0.930 4.730 -0.610 4.760 ;
        RECT 0.280 4.740 0.710 5.000 ;
        RECT -0.930 4.540 -0.600 4.730 ;
        RECT 0.510 4.700 0.710 4.740 ;
        RECT 1.100 4.700 1.650 5.690 ;
        RECT 1.970 5.610 2.820 5.840 ;
        RECT 2.120 5.270 2.820 5.610 ;
        RECT 2.580 4.910 2.900 4.950 ;
        RECT 2.580 4.850 2.910 4.910 ;
        RECT 2.110 4.720 2.910 4.850 ;
        RECT 2.110 4.690 2.900 4.720 ;
        RECT 2.110 4.670 2.810 4.690 ;
        RECT -0.930 4.500 -0.610 4.540 ;
        RECT -0.930 4.420 -0.760 4.500 ;
        RECT -0.980 4.250 -0.760 4.420 ;
        RECT -0.980 4.090 -0.810 4.250 ;
        RECT 2.570 4.190 2.890 4.230 ;
        RECT 0.510 4.150 0.710 4.190 ;
        RECT -0.450 3.830 -0.260 3.950 ;
        RECT 0.280 3.890 0.710 4.150 ;
        RECT 0.510 3.860 0.710 3.890 ;
        RECT -0.810 3.720 -0.260 3.830 ;
        RECT -0.810 3.660 -0.270 3.720 ;
        RECT -0.730 1.880 -0.560 3.660 ;
        RECT 0.100 3.500 0.270 3.540 ;
        RECT 0.510 3.500 0.710 3.530 ;
        RECT 0.100 3.240 0.710 3.500 ;
        RECT 0.100 3.210 0.270 3.240 ;
        RECT 0.510 3.200 0.710 3.240 ;
        RECT 1.100 3.200 1.650 4.190 ;
        RECT 2.110 4.010 2.900 4.190 ;
        RECT 2.570 4.000 2.900 4.010 ;
        RECT 2.570 3.970 2.890 4.000 ;
        RECT 2.120 3.250 2.820 3.590 ;
        RECT 1.970 3.020 2.820 3.250 ;
        RECT 2.120 2.710 2.820 3.020 ;
        RECT 0.100 2.650 0.270 2.680 ;
        RECT 0.510 2.650 0.710 2.690 ;
        RECT 0.100 2.390 0.710 2.650 ;
        RECT 0.100 2.350 0.270 2.390 ;
        RECT 0.510 2.360 0.710 2.390 ;
        RECT 0.510 2.000 0.710 2.030 ;
        RECT 0.280 1.740 0.710 2.000 ;
        RECT -2.520 1.710 -2.350 1.730 ;
        RECT -2.520 1.450 -1.960 1.710 ;
        RECT 0.510 1.700 0.710 1.740 ;
        RECT 1.100 1.700 1.650 2.690 ;
        RECT 2.120 2.100 2.830 2.270 ;
        RECT 2.470 1.820 2.830 2.100 ;
        RECT 2.470 1.650 3.100 1.820 ;
        RECT -2.520 1.400 -2.350 1.450 ;
      LAYER mcon ;
        RECT -0.630 7.180 -0.460 7.350 ;
        RECT -3.790 6.570 -3.620 6.740 ;
        RECT -10.630 5.990 -10.460 6.160 ;
        RECT -14.290 5.390 -14.020 5.660 ;
        RECT -10.630 5.540 -10.460 5.710 ;
        RECT -5.460 5.740 -5.290 5.910 ;
        RECT -4.150 5.730 -3.970 5.920 ;
        RECT -11.870 4.620 -11.700 4.790 ;
        RECT -11.870 4.280 -11.700 4.450 ;
        RECT -14.290 3.660 -14.020 3.930 ;
        RECT -11.870 3.930 -11.700 4.100 ;
        RECT -10.630 3.040 -10.460 3.210 ;
        RECT -5.460 2.980 -5.290 3.150 ;
        RECT -10.630 2.590 -10.460 2.760 ;
        RECT -4.150 2.930 -3.970 3.120 ;
        RECT 0.340 6.930 0.510 7.100 ;
        RECT 1.320 6.610 1.490 6.780 ;
        RECT 2.590 6.950 2.760 7.120 ;
        RECT -0.480 6.350 -0.310 6.520 ;
        RECT -1.600 5.830 -1.430 6.000 ;
        RECT -2.000 4.930 -1.830 5.100 ;
        RECT -2.430 4.130 -2.260 4.300 ;
        RECT -3.160 2.850 -2.990 3.020 ;
        RECT -3.790 2.110 -3.620 2.280 ;
        RECT -2.040 2.330 -1.870 2.500 ;
        RECT 0.290 6.280 0.460 6.450 ;
        RECT 0.290 5.440 0.460 5.610 ;
        RECT 1.980 5.640 2.150 5.810 ;
        RECT 1.320 5.110 1.490 5.280 ;
        RECT 0.340 4.790 0.510 4.960 ;
        RECT -0.870 4.550 -0.700 4.720 ;
        RECT 2.640 4.730 2.810 4.900 ;
        RECT -0.440 3.750 -0.270 3.920 ;
        RECT 0.340 3.930 0.510 4.100 ;
        RECT 2.630 4.010 2.800 4.180 ;
        RECT 1.320 3.610 1.490 3.780 ;
        RECT 0.290 3.280 0.460 3.450 ;
        RECT 1.980 3.050 2.150 3.220 ;
        RECT 0.290 2.440 0.460 2.610 ;
        RECT 1.320 2.110 1.490 2.280 ;
        RECT 0.340 1.790 0.510 1.960 ;
        RECT 2.550 1.760 2.720 1.930 ;
        RECT -2.190 1.500 -2.020 1.670 ;
      LAYER met1 ;
        RECT -11.900 4.880 -11.670 7.450 ;
        RECT -5.680 6.630 -5.370 7.070 ;
        RECT -3.720 6.800 -3.440 7.450 ;
        RECT -0.710 7.110 -0.390 7.430 ;
        RECT 0.270 6.860 0.590 7.180 ;
        RECT 2.520 6.880 2.840 7.200 ;
        RECT -3.830 6.200 -3.440 6.800 ;
        RECT -0.560 6.280 -0.240 6.600 ;
        RECT 0.220 6.210 0.540 6.530 ;
        RECT -5.530 5.670 -5.210 5.990 ;
        RECT -4.560 4.880 -4.320 5.010 ;
        RECT -11.940 3.870 -11.560 4.880 ;
        RECT -4.560 4.560 -4.300 4.880 ;
        RECT -3.720 4.600 -3.440 6.200 ;
        RECT -1.670 5.750 -1.350 6.070 ;
        RECT -0.450 5.590 -0.240 5.700 ;
        RECT -0.470 5.270 -0.210 5.590 ;
        RECT 0.220 5.360 0.540 5.680 ;
        RECT -2.030 4.870 -1.800 5.160 ;
        RECT -3.720 4.280 -3.360 4.600 ;
        RECT -4.560 3.960 -4.300 4.280 ;
        RECT -11.900 1.400 -11.670 3.870 ;
        RECT -4.560 3.840 -4.320 3.960 ;
        RECT -5.530 2.910 -5.210 3.230 ;
        RECT -3.720 2.650 -3.440 4.280 ;
        RECT -2.500 4.060 -2.180 4.380 ;
        RECT -2.010 3.580 -1.800 4.870 ;
        RECT -0.940 4.470 -0.620 4.790 ;
        RECT -0.450 3.980 -0.240 5.270 ;
        RECT 0.270 4.710 0.590 5.030 ;
        RECT 2.570 4.660 2.890 4.980 ;
        RECT -0.470 3.690 -0.240 3.980 ;
        RECT 0.270 3.860 0.590 4.180 ;
        RECT 2.560 3.940 2.880 4.260 ;
        RECT -2.030 3.260 -1.770 3.580 ;
        RECT -2.010 3.150 -1.800 3.260 ;
        RECT 0.220 3.210 0.540 3.530 ;
        RECT -3.230 2.780 -2.910 3.100 ;
        RECT -5.680 1.780 -5.370 2.220 ;
        RECT -3.830 2.050 -3.440 2.650 ;
        RECT -2.120 2.250 -1.800 2.570 ;
        RECT 0.220 2.360 0.540 2.680 ;
        RECT -3.720 1.400 -3.440 2.050 ;
        RECT -2.270 1.420 -1.950 1.740 ;
        RECT 0.270 1.710 0.590 2.030 ;
        RECT 2.480 1.690 2.800 2.010 ;
      LAYER via ;
        RECT -5.650 6.660 -5.390 6.920 ;
        RECT -0.680 7.140 -0.420 7.400 ;
        RECT 0.300 6.890 0.560 7.150 ;
        RECT 2.550 6.910 2.810 7.170 ;
        RECT -0.530 6.310 -0.270 6.570 ;
        RECT 0.250 6.240 0.510 6.500 ;
        RECT -5.500 5.700 -5.240 5.960 ;
        RECT -11.900 3.910 -11.610 4.840 ;
        RECT -4.560 4.590 -4.300 4.850 ;
        RECT -1.640 5.780 -1.380 6.040 ;
        RECT -0.470 5.300 -0.210 5.560 ;
        RECT 0.250 5.390 0.510 5.650 ;
        RECT -3.620 4.310 -3.360 4.570 ;
        RECT -4.560 3.990 -4.300 4.250 ;
        RECT -5.500 2.940 -5.240 3.200 ;
        RECT -2.470 4.090 -2.210 4.350 ;
        RECT -0.910 4.500 -0.650 4.760 ;
        RECT 0.300 4.740 0.560 5.000 ;
        RECT 2.600 4.690 2.860 4.950 ;
        RECT 0.300 3.890 0.560 4.150 ;
        RECT 2.590 3.970 2.850 4.230 ;
        RECT -2.030 3.290 -1.770 3.550 ;
        RECT 0.250 3.240 0.510 3.500 ;
        RECT -3.200 2.810 -2.940 3.070 ;
        RECT -5.650 1.930 -5.390 2.190 ;
        RECT -2.090 2.280 -1.830 2.540 ;
        RECT 0.250 2.390 0.510 2.650 ;
        RECT 0.300 1.740 0.560 2.000 ;
        RECT 2.510 1.720 2.770 1.980 ;
        RECT -2.240 1.450 -1.980 1.710 ;
      LAYER met2 ;
        RECT 0.270 7.110 0.580 7.190 ;
        RECT 2.520 7.110 2.830 7.210 ;
        RECT 0.270 6.880 2.830 7.110 ;
        RECT 0.270 6.860 0.580 6.880 ;
        RECT -0.550 6.570 -0.240 6.610 ;
        RECT -0.730 6.460 0.010 6.570 ;
        RECT 0.220 6.460 0.530 6.540 ;
        RECT -0.730 6.320 0.530 6.460 ;
        RECT -0.550 6.280 0.530 6.320 ;
        RECT -0.240 6.250 0.530 6.280 ;
        RECT -0.240 6.200 0.010 6.250 ;
        RECT 0.220 6.210 0.530 6.250 ;
        RECT -5.530 5.930 -5.220 6.000 ;
        RECT -1.670 5.930 -1.360 6.070 ;
        RECT -5.530 5.740 -1.360 5.930 ;
        RECT -5.530 5.710 -1.620 5.740 ;
        RECT -5.530 5.670 -5.220 5.710 ;
        RECT 0.220 5.640 0.530 5.680 ;
        RECT -0.210 5.560 0.530 5.640 ;
        RECT -0.500 5.540 0.530 5.560 ;
        RECT -0.550 5.430 0.530 5.540 ;
        RECT -0.550 5.350 0.000 5.430 ;
        RECT 0.220 5.350 0.530 5.430 ;
        RECT -0.550 5.290 -0.080 5.350 ;
        RECT -2.110 3.470 -1.640 3.560 ;
        RECT -2.110 3.460 0.000 3.470 ;
        RECT 0.220 3.460 0.530 3.540 ;
        RECT -2.110 3.310 0.530 3.460 ;
        RECT -2.060 3.290 0.530 3.310 ;
        RECT -1.770 3.270 0.530 3.290 ;
        RECT -0.080 3.250 0.530 3.270 ;
        RECT -5.530 3.170 -5.220 3.240 ;
        RECT 0.220 3.210 0.530 3.250 ;
        RECT -3.340 3.170 -3.180 3.180 ;
        RECT -5.530 3.110 -3.180 3.170 ;
        RECT -5.530 2.960 -2.920 3.110 ;
        RECT -5.530 2.910 -5.220 2.960 ;
        RECT -3.340 2.780 -2.920 2.960 ;
        RECT -2.060 2.640 0.000 2.670 ;
        RECT 0.220 2.640 0.530 2.680 ;
        RECT -2.060 2.570 0.530 2.640 ;
        RECT -2.110 2.530 0.530 2.570 ;
        RECT -2.290 2.460 0.530 2.530 ;
        RECT -2.290 2.280 -1.740 2.460 ;
        RECT -0.080 2.430 0.530 2.460 ;
        RECT 0.220 2.350 0.530 2.430 ;
        RECT -2.110 2.240 -1.800 2.280 ;
        RECT 0.270 1.980 0.580 2.030 ;
        RECT 2.480 1.980 2.790 2.020 ;
        RECT 0.270 1.750 2.980 1.980 ;
        RECT 0.270 1.700 0.580 1.750 ;
        RECT 2.480 1.690 2.790 1.750 ;
  END
END sky130_hilas_TA2Cell_NoFG

MACRO sky130_hilas_FGBias2x1cell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_FGBias2x1cell ;
  ORIGIN 3.960 3.870 ;
  SIZE 11.530 BY 6.150 ;
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 2.516100 ;
    PORT
      LAYER nwell ;
        RECT -3.950 1.480 -2.220 2.230 ;
        RECT -3.950 0.330 -2.210 1.480 ;
        RECT -3.940 -1.910 -2.210 0.330 ;
        RECT -3.950 -2.090 -2.210 -1.910 ;
        RECT -3.950 -3.810 -2.220 -2.090 ;
      LAYER met1 ;
        RECT -3.610 -3.820 -3.190 2.230 ;
    END
  END VTUN
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT -1.130 -3.820 -0.900 2.230 ;
    END
  END VGND
  PIN GATE_CONTROL
    USE ANALOG ;
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT -0.190 -0.160 2.530 1.490 ;
        RECT -0.190 -0.200 2.520 -0.160 ;
        RECT -0.190 -1.530 2.520 -1.490 ;
        RECT -0.190 -3.180 2.530 -1.530 ;
      LAYER met1 ;
        RECT 0.090 1.020 0.320 2.230 ;
        RECT 0.090 0.230 0.350 1.020 ;
        RECT 0.090 -1.920 0.320 0.230 ;
        RECT 0.090 -2.710 0.350 -1.920 ;
        RECT 0.090 -3.820 0.320 -2.710 ;
    END
  END GATE_CONTROL
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 5.090 1.730 5.400 1.740 ;
        RECT -3.960 1.550 7.570 1.730 ;
        RECT 5.090 1.410 5.400 1.550 ;
    END
  END DRAIN1
  PIN DRAIN4
    USE ANALOG ;
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 5.090 -3.140 5.400 -3.000 ;
        RECT 5.090 -3.150 7.570 -3.140 ;
        RECT -3.960 -3.300 7.570 -3.150 ;
        RECT 5.090 -3.320 7.570 -3.300 ;
        RECT 5.090 -3.330 5.400 -3.320 ;
    END
  END DRAIN4
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 4.260 -3.870 7.570 2.280 ;
      LAYER met2 ;
        RECT 6.180 -0.630 6.500 -0.370 ;
        RECT 6.220 -0.650 7.400 -0.630 ;
        RECT 6.220 -0.910 7.440 -0.650 ;
        RECT 6.220 -0.970 7.400 -0.910 ;
        RECT 6.180 -0.980 7.400 -0.970 ;
        RECT 6.180 -1.230 6.500 -0.980 ;
    END
  END VINJ
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 5.240 0.710 5.550 0.780 ;
        RECT 5.240 0.490 7.570 0.710 ;
        RECT 5.240 0.450 5.550 0.490 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 5.240 -2.050 5.550 -1.980 ;
        RECT 5.240 -2.260 7.570 -2.050 ;
        RECT 5.240 -2.310 5.550 -2.260 ;
    END
  END OUTPUT2
  PIN GATECOL
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT 6.610 0.770 6.800 2.230 ;
        RECT 6.610 0.740 6.830 0.770 ;
        RECT 6.590 0.470 6.840 0.740 ;
        RECT 6.600 0.460 6.840 0.470 ;
        RECT 6.600 0.220 6.830 0.460 ;
        RECT 6.640 -1.810 6.800 0.220 ;
        RECT 6.600 -2.050 6.830 -1.810 ;
        RECT 6.600 -2.060 6.840 -2.050 ;
        RECT 6.590 -2.330 6.840 -2.060 ;
        RECT 6.610 -2.360 6.830 -2.330 ;
        RECT 6.610 -3.820 6.800 -2.360 ;
    END
  END GATECOL
  PIN VINJ
    ANTENNADIFFAREA 0.544000 ;
    PORT
      LAYER met1 ;
        RECT 7.050 1.580 7.330 2.230 ;
        RECT 6.940 0.980 7.330 1.580 ;
        RECT 7.050 -0.620 7.330 0.980 ;
        RECT 7.050 -0.940 7.410 -0.620 ;
        RECT 7.050 -2.570 7.330 -0.940 ;
        RECT 6.940 -3.170 7.330 -2.570 ;
        RECT 7.050 -3.820 7.330 -3.170 ;
      LAYER via ;
        RECT 7.150 -0.910 7.410 -0.650 ;
    END
  END VINJ
  OBS
      LAYER li1 ;
        RECT 5.160 1.650 5.690 1.820 ;
        RECT 6.970 1.550 7.170 1.900 ;
        RECT 6.970 1.520 7.180 1.550 ;
        RECT -3.520 0.090 -2.970 0.520 ;
        RECT 0.110 0.280 0.340 0.970 ;
        RECT 5.410 0.740 5.580 1.260 ;
        RECT 5.250 0.480 5.580 0.740 ;
        RECT -0.920 -0.740 -0.730 -0.340 ;
        RECT 5.410 -0.430 5.580 0.480 ;
        RECT 6.240 -0.340 6.410 1.270 ;
        RECT 6.960 0.940 7.180 1.520 ;
        RECT 6.970 0.930 7.180 0.940 ;
        RECT 6.610 0.760 6.800 0.770 ;
        RECT 6.610 0.470 6.810 0.760 ;
        RECT 6.600 0.140 6.890 0.470 ;
        RECT 6.240 -0.530 6.420 -0.340 ;
        RECT -1.110 -0.750 -0.730 -0.740 ;
        RECT -1.110 -0.930 2.630 -0.750 ;
        RECT -1.110 -0.970 -0.730 -0.930 ;
        RECT -3.520 -1.640 -2.970 -1.210 ;
        RECT -0.920 -1.350 -0.730 -0.970 ;
        RECT 0.110 -2.660 0.340 -1.930 ;
        RECT 5.410 -2.020 5.580 -1.160 ;
        RECT 5.250 -2.280 5.580 -2.020 ;
        RECT 5.410 -2.850 5.580 -2.280 ;
        RECT 6.240 -1.250 6.420 -1.060 ;
        RECT 6.240 -2.860 6.410 -1.250 ;
        RECT 6.600 -2.060 6.890 -1.730 ;
        RECT 6.610 -2.350 6.810 -2.060 ;
        RECT 6.610 -2.360 6.800 -2.350 ;
        RECT 6.970 -2.530 7.180 -2.520 ;
        RECT 6.960 -3.110 7.180 -2.530 ;
        RECT 6.970 -3.140 7.180 -3.110 ;
        RECT 5.160 -3.410 5.690 -3.240 ;
        RECT 6.970 -3.490 7.170 -3.140 ;
      LAYER mcon ;
        RECT 6.980 1.350 7.150 1.520 ;
        RECT 0.140 0.770 0.310 0.940 ;
        RECT -3.520 0.170 -3.250 0.440 ;
        RECT 0.140 0.320 0.310 0.490 ;
        RECT 5.310 0.520 5.480 0.690 ;
        RECT 6.620 0.510 6.800 0.700 ;
        RECT -1.100 -0.940 -0.930 -0.770 ;
        RECT -3.520 -1.560 -3.250 -1.290 ;
        RECT 0.140 -2.180 0.310 -2.010 ;
        RECT 5.310 -2.240 5.480 -2.070 ;
        RECT 0.140 -2.630 0.310 -2.460 ;
        RECT 6.620 -2.290 6.800 -2.100 ;
        RECT 6.980 -3.110 7.150 -2.940 ;
      LAYER met1 ;
        RECT 5.090 1.410 5.400 1.850 ;
        RECT 5.240 0.450 5.560 0.770 ;
        RECT 6.210 -0.340 6.450 -0.210 ;
        RECT 6.210 -0.660 6.470 -0.340 ;
        RECT 6.210 -1.260 6.470 -0.940 ;
        RECT 6.210 -1.380 6.450 -1.260 ;
        RECT 5.240 -2.310 5.560 -1.990 ;
        RECT 5.090 -3.440 5.400 -3.000 ;
      LAYER via ;
        RECT 5.120 1.440 5.380 1.700 ;
        RECT 5.270 0.480 5.530 0.740 ;
        RECT 6.210 -0.630 6.470 -0.370 ;
        RECT 6.210 -1.230 6.470 -0.970 ;
        RECT 5.270 -2.280 5.530 -2.020 ;
        RECT 5.120 -3.290 5.380 -3.030 ;
  END
END sky130_hilas_FGBias2x1cell

MACRO sky130_hilas_Tgate4Single01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_Tgate4Single01 ;
  ORIGIN 0.360 1.640 ;
  SIZE 4.760 BY 6.410 ;
  PIN VPWR
    USE ANALOG ;
    ANTENNADIFFAREA 0.966800 ;
    PORT
      LAYER nwell ;
        RECT -0.240 -1.640 2.520 4.770 ;
      LAYER met1 ;
        RECT 0.380 3.850 0.580 4.770 ;
        RECT 0.370 3.560 0.600 3.850 ;
        RECT 0.380 2.770 0.580 3.560 ;
        RECT 0.370 2.480 0.600 2.770 ;
        RECT 0.380 0.650 0.580 2.480 ;
        RECT 0.370 0.360 0.600 0.650 ;
        RECT 0.380 -0.430 0.580 0.360 ;
        RECT 0.370 -0.720 0.600 -0.430 ;
        RECT 0.380 -1.640 0.580 -0.720 ;
    END
  END VPWR
  PIN INPUT1_2
    USE ANALOG ;
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT 1.280 1.930 1.590 2.050 ;
        RECT 0.510 1.920 1.630 1.930 ;
        RECT 2.850 1.920 3.160 2.050 ;
        RECT -0.360 1.720 3.160 1.920 ;
        RECT 0.510 1.710 1.630 1.720 ;
    END
  END INPUT1_2
  PIN SELECT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT -0.070 2.900 0.250 2.990 ;
        RECT -0.360 2.700 0.250 2.900 ;
    END
  END SELECT2
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 3.890 3.850 4.080 4.770 ;
        RECT 3.870 3.560 4.100 3.850 ;
        RECT 3.890 2.770 4.080 3.560 ;
        RECT 3.870 2.480 4.100 2.770 ;
        RECT 3.890 0.650 4.080 2.480 ;
        RECT 3.870 0.360 4.100 0.650 ;
        RECT 3.890 -0.430 4.080 0.360 ;
        RECT 3.870 -0.720 4.100 -0.430 ;
        RECT 3.890 -1.640 4.080 -0.720 ;
    END
  END VGND
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.212400 ;
    PORT
      LAYER met2 ;
        RECT 2.200 2.900 2.520 2.920 ;
        RECT 3.210 2.900 3.530 2.930 ;
        RECT 2.150 2.700 4.400 2.900 ;
        RECT 2.200 2.660 2.520 2.700 ;
        RECT 3.210 2.670 3.530 2.700 ;
    END
  END OUTPUT2
  PIN OUTPUT4
    ANTENNADIFFAREA 0.212400 ;
    PORT
      LAYER met2 ;
        RECT 2.200 -0.300 2.520 -0.280 ;
        RECT 3.210 -0.300 3.530 -0.270 ;
        RECT 2.150 -0.500 4.400 -0.300 ;
        RECT 2.200 -0.540 2.520 -0.500 ;
        RECT 3.210 -0.530 3.530 -0.500 ;
    END
  END OUTPUT4
  PIN OUTPUT3
    ANTENNADIFFAREA 0.212400 ;
    PORT
      LAYER met2 ;
        RECT 2.200 0.430 2.520 0.470 ;
        RECT 3.210 0.430 3.530 0.460 ;
        RECT 2.150 0.230 4.400 0.430 ;
        RECT 2.200 0.210 2.520 0.230 ;
        RECT 3.210 0.200 3.530 0.230 ;
    END
  END OUTPUT3
  PIN OUTPUT1
    ANTENNADIFFAREA 0.212400 ;
    PORT
      LAYER met2 ;
        RECT 2.200 3.630 2.520 3.670 ;
        RECT 3.210 3.630 3.530 3.660 ;
        RECT 2.150 3.430 4.400 3.630 ;
        RECT 2.200 3.410 2.520 3.430 ;
        RECT 3.210 3.400 3.530 3.430 ;
    END
  END OUTPUT1
  PIN INPUT1_4
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT 1.280 -1.270 1.590 -1.150 ;
        RECT 0.510 -1.280 1.630 -1.270 ;
        RECT 2.850 -1.280 3.160 -1.150 ;
        RECT -0.360 -1.480 3.160 -1.280 ;
        RECT 0.510 -1.490 1.630 -1.480 ;
    END
  END INPUT1_4
  PIN SELECT4
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT -0.070 -0.300 0.250 -0.210 ;
        RECT -0.360 -0.500 0.250 -0.300 ;
    END
  END SELECT4
  PIN SELECT3
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT -0.360 0.230 0.250 0.430 ;
        RECT -0.070 0.140 0.250 0.230 ;
    END
  END SELECT3
  PIN INPUT1_3
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT 0.510 1.410 1.630 1.420 ;
        RECT -0.360 1.210 3.160 1.410 ;
        RECT 0.510 1.200 1.630 1.210 ;
        RECT 1.280 1.080 1.590 1.200 ;
        RECT 2.850 1.080 3.160 1.210 ;
    END
  END INPUT1_3
  PIN SELECT1
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT -0.360 3.430 0.250 3.630 ;
        RECT -0.070 3.340 0.250 3.430 ;
    END
  END SELECT1
  PIN INPUT1_1
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT 0.510 4.610 1.630 4.620 ;
        RECT -0.360 4.410 3.160 4.610 ;
        RECT 0.510 4.400 1.630 4.410 ;
        RECT 1.280 4.280 1.590 4.400 ;
        RECT 2.850 4.280 3.160 4.410 ;
    END
  END INPUT1_1
  OBS
      LAYER li1 ;
        RECT 1.290 4.550 1.610 4.580 ;
        RECT 2.860 4.550 3.180 4.580 ;
        RECT 0.070 4.210 0.240 4.490 ;
        RECT 1.290 4.360 1.620 4.550 ;
        RECT 2.300 4.410 2.490 4.430 ;
        RECT 1.290 4.320 1.610 4.360 ;
        RECT 0.070 4.170 0.280 4.210 ;
        RECT 0.070 4.150 0.300 4.170 ;
        RECT 1.420 4.160 1.590 4.320 ;
        RECT 2.030 4.240 2.490 4.410 ;
        RECT 2.860 4.360 3.190 4.550 ;
        RECT 3.430 4.410 3.620 4.440 ;
        RECT 2.860 4.320 3.180 4.360 ;
        RECT 2.280 4.230 2.490 4.240 ;
        RECT 2.300 4.200 2.490 4.230 ;
        RECT 2.920 4.160 3.090 4.320 ;
        RECT 3.430 4.240 3.870 4.410 ;
        RECT 3.430 4.210 3.620 4.240 ;
        RECT 0.070 4.130 0.330 4.150 ;
        RECT 0.070 4.080 0.410 4.130 ;
        RECT 0.070 4.020 0.560 4.080 ;
        RECT 0.070 3.990 0.580 4.020 ;
        RECT 0.110 3.960 0.580 3.990 ;
        RECT 0.240 3.910 0.580 3.960 ;
        RECT 0.360 3.900 0.580 3.910 ;
        RECT 0.370 3.870 0.580 3.900 ;
        RECT 0.390 3.790 0.580 3.870 ;
        RECT 1.750 3.790 2.080 3.910 ;
        RECT 4.150 3.820 4.320 4.500 ;
        RECT -0.100 3.740 0.070 3.760 ;
        RECT -0.120 3.310 0.090 3.740 ;
        RECT 0.390 3.620 0.910 3.790 ;
        RECT 0.390 3.590 0.580 3.620 ;
        RECT 1.260 3.610 3.160 3.790 ;
        RECT 3.890 3.780 4.320 3.820 ;
        RECT 3.540 3.620 4.320 3.780 ;
        RECT 3.540 3.610 4.080 3.620 ;
        RECT 3.890 3.590 4.080 3.610 ;
        RECT -0.120 2.590 0.090 3.020 ;
        RECT 0.390 2.710 0.580 2.740 ;
        RECT 3.890 2.720 4.080 2.740 ;
        RECT -0.100 2.570 0.070 2.590 ;
        RECT 0.390 2.540 0.910 2.710 ;
        RECT 1.260 2.540 3.160 2.720 ;
        RECT 3.540 2.710 4.080 2.720 ;
        RECT 3.540 2.550 4.320 2.710 ;
        RECT 0.390 2.460 0.580 2.540 ;
        RECT 0.370 2.430 0.580 2.460 ;
        RECT 0.360 2.420 0.580 2.430 ;
        RECT 1.750 2.420 2.080 2.540 ;
        RECT 3.890 2.510 4.320 2.550 ;
        RECT 0.240 2.370 0.580 2.420 ;
        RECT 0.110 2.340 0.580 2.370 ;
        RECT 0.070 2.310 0.580 2.340 ;
        RECT 0.070 2.250 0.560 2.310 ;
        RECT 0.070 2.200 0.410 2.250 ;
        RECT 0.070 2.180 0.330 2.200 ;
        RECT 0.070 2.160 0.300 2.180 ;
        RECT 0.070 2.120 0.280 2.160 ;
        RECT 0.070 1.840 0.240 2.120 ;
        RECT 1.420 2.010 1.590 2.170 ;
        RECT 2.300 2.100 2.490 2.130 ;
        RECT 2.280 2.090 2.490 2.100 ;
        RECT 1.290 1.970 1.610 2.010 ;
        RECT 1.290 1.780 1.620 1.970 ;
        RECT 2.030 1.920 2.490 2.090 ;
        RECT 2.920 2.010 3.090 2.170 ;
        RECT 3.430 2.090 3.620 2.120 ;
        RECT 2.300 1.900 2.490 1.920 ;
        RECT 2.860 1.970 3.180 2.010 ;
        RECT 2.860 1.780 3.190 1.970 ;
        RECT 3.430 1.920 3.870 2.090 ;
        RECT 3.430 1.890 3.620 1.920 ;
        RECT 4.150 1.830 4.320 2.510 ;
        RECT 1.290 1.750 1.610 1.780 ;
        RECT 2.860 1.750 3.180 1.780 ;
        RECT 1.290 1.350 1.610 1.380 ;
        RECT 2.860 1.350 3.180 1.380 ;
        RECT 0.070 1.010 0.240 1.290 ;
        RECT 1.290 1.160 1.620 1.350 ;
        RECT 2.300 1.210 2.490 1.230 ;
        RECT 1.290 1.120 1.610 1.160 ;
        RECT 0.070 0.970 0.280 1.010 ;
        RECT 0.070 0.950 0.300 0.970 ;
        RECT 1.420 0.960 1.590 1.120 ;
        RECT 2.030 1.040 2.490 1.210 ;
        RECT 2.860 1.160 3.190 1.350 ;
        RECT 3.430 1.210 3.620 1.240 ;
        RECT 2.860 1.120 3.180 1.160 ;
        RECT 2.280 1.030 2.490 1.040 ;
        RECT 2.300 1.000 2.490 1.030 ;
        RECT 2.920 0.960 3.090 1.120 ;
        RECT 3.430 1.040 3.870 1.210 ;
        RECT 3.430 1.010 3.620 1.040 ;
        RECT 0.070 0.930 0.330 0.950 ;
        RECT 0.070 0.880 0.410 0.930 ;
        RECT 0.070 0.820 0.560 0.880 ;
        RECT 0.070 0.790 0.580 0.820 ;
        RECT 0.110 0.760 0.580 0.790 ;
        RECT 0.240 0.710 0.580 0.760 ;
        RECT 0.360 0.700 0.580 0.710 ;
        RECT 0.370 0.670 0.580 0.700 ;
        RECT 0.390 0.590 0.580 0.670 ;
        RECT 1.750 0.590 2.080 0.710 ;
        RECT 4.150 0.620 4.320 1.300 ;
        RECT -0.100 0.540 0.070 0.560 ;
        RECT -0.120 0.110 0.090 0.540 ;
        RECT 0.390 0.420 0.910 0.590 ;
        RECT 0.390 0.390 0.580 0.420 ;
        RECT 1.260 0.410 3.160 0.590 ;
        RECT 3.890 0.580 4.320 0.620 ;
        RECT 3.540 0.420 4.320 0.580 ;
        RECT 3.540 0.410 4.080 0.420 ;
        RECT 3.890 0.390 4.080 0.410 ;
        RECT -0.120 -0.610 0.090 -0.180 ;
        RECT 0.390 -0.490 0.580 -0.460 ;
        RECT 3.890 -0.480 4.080 -0.460 ;
        RECT -0.100 -0.630 0.070 -0.610 ;
        RECT 0.390 -0.660 0.910 -0.490 ;
        RECT 1.260 -0.660 3.160 -0.480 ;
        RECT 3.540 -0.490 4.080 -0.480 ;
        RECT 3.540 -0.650 4.320 -0.490 ;
        RECT 0.390 -0.740 0.580 -0.660 ;
        RECT 0.370 -0.770 0.580 -0.740 ;
        RECT 0.360 -0.780 0.580 -0.770 ;
        RECT 1.750 -0.780 2.080 -0.660 ;
        RECT 3.890 -0.690 4.320 -0.650 ;
        RECT 0.240 -0.830 0.580 -0.780 ;
        RECT 0.110 -0.860 0.580 -0.830 ;
        RECT 0.070 -0.890 0.580 -0.860 ;
        RECT 0.070 -0.950 0.560 -0.890 ;
        RECT 0.070 -1.000 0.410 -0.950 ;
        RECT 0.070 -1.020 0.330 -1.000 ;
        RECT 0.070 -1.040 0.300 -1.020 ;
        RECT 0.070 -1.080 0.280 -1.040 ;
        RECT 0.070 -1.360 0.240 -1.080 ;
        RECT 1.420 -1.190 1.590 -1.030 ;
        RECT 2.300 -1.100 2.490 -1.070 ;
        RECT 2.280 -1.110 2.490 -1.100 ;
        RECT 1.290 -1.230 1.610 -1.190 ;
        RECT 1.290 -1.420 1.620 -1.230 ;
        RECT 2.030 -1.280 2.490 -1.110 ;
        RECT 2.920 -1.190 3.090 -1.030 ;
        RECT 3.430 -1.110 3.620 -1.080 ;
        RECT 2.300 -1.300 2.490 -1.280 ;
        RECT 2.860 -1.230 3.180 -1.190 ;
        RECT 2.860 -1.420 3.190 -1.230 ;
        RECT 3.430 -1.280 3.870 -1.110 ;
        RECT 3.430 -1.310 3.620 -1.280 ;
        RECT 4.150 -1.370 4.320 -0.690 ;
        RECT 1.290 -1.450 1.610 -1.420 ;
        RECT 2.860 -1.450 3.180 -1.420 ;
      LAYER mcon ;
        RECT 1.350 4.370 1.520 4.540 ;
        RECT 2.310 4.230 2.480 4.400 ;
        RECT 2.920 4.370 3.090 4.540 ;
        RECT 3.440 4.240 3.610 4.410 ;
        RECT -0.100 3.590 0.070 3.760 ;
        RECT 0.400 3.620 0.570 3.790 ;
        RECT 3.900 3.620 4.070 3.790 ;
        RECT 0.400 2.540 0.570 2.710 ;
        RECT 3.900 2.540 4.070 2.710 ;
        RECT 1.350 1.790 1.520 1.960 ;
        RECT 2.310 1.930 2.480 2.100 ;
        RECT 2.920 1.790 3.090 1.960 ;
        RECT 3.440 1.920 3.610 2.090 ;
        RECT 1.350 1.170 1.520 1.340 ;
        RECT 2.310 1.030 2.480 1.200 ;
        RECT 2.920 1.170 3.090 1.340 ;
        RECT 3.440 1.040 3.610 1.210 ;
        RECT -0.100 0.390 0.070 0.560 ;
        RECT 0.400 0.420 0.570 0.590 ;
        RECT 3.900 0.420 4.070 0.590 ;
        RECT 0.400 -0.660 0.570 -0.490 ;
        RECT 3.900 -0.660 4.070 -0.490 ;
        RECT 1.350 -1.410 1.520 -1.240 ;
        RECT 2.310 -1.270 2.480 -1.100 ;
        RECT 2.920 -1.410 3.090 -1.240 ;
        RECT 3.440 -1.280 3.610 -1.110 ;
      LAYER met1 ;
        RECT 1.280 4.290 1.600 4.610 ;
        RECT 2.280 4.170 2.510 4.460 ;
        RECT 2.850 4.290 3.170 4.610 ;
        RECT 3.410 4.180 3.640 4.470 ;
        RECT -0.130 3.630 0.100 3.820 ;
        RECT 2.300 3.700 2.490 4.170 ;
        RECT -0.130 3.530 0.220 3.630 ;
        RECT -0.120 3.310 0.220 3.530 ;
        RECT 2.230 3.380 2.490 3.700 ;
        RECT 3.410 3.690 3.600 4.180 ;
        RECT 3.230 3.440 3.600 3.690 ;
        RECT 3.230 3.370 3.500 3.440 ;
        RECT -0.120 2.800 0.220 3.020 ;
        RECT -0.130 2.700 0.220 2.800 ;
        RECT -0.130 2.510 0.100 2.700 ;
        RECT 2.230 2.630 2.490 2.950 ;
        RECT 3.230 2.890 3.500 2.960 ;
        RECT 3.230 2.640 3.600 2.890 ;
        RECT 2.300 2.160 2.490 2.630 ;
        RECT 1.280 1.720 1.600 2.040 ;
        RECT 2.280 1.870 2.510 2.160 ;
        RECT 3.410 2.150 3.600 2.640 ;
        RECT 2.850 1.720 3.170 2.040 ;
        RECT 3.410 1.860 3.640 2.150 ;
        RECT 1.280 1.090 1.600 1.410 ;
        RECT 2.280 0.970 2.510 1.260 ;
        RECT 2.850 1.090 3.170 1.410 ;
        RECT 3.410 0.980 3.640 1.270 ;
        RECT -0.130 0.430 0.100 0.620 ;
        RECT 2.300 0.500 2.490 0.970 ;
        RECT -0.130 0.330 0.220 0.430 ;
        RECT -0.120 0.110 0.220 0.330 ;
        RECT 2.230 0.180 2.490 0.500 ;
        RECT 3.410 0.490 3.600 0.980 ;
        RECT 3.230 0.240 3.600 0.490 ;
        RECT 3.230 0.170 3.500 0.240 ;
        RECT -0.120 -0.400 0.220 -0.180 ;
        RECT -0.130 -0.500 0.220 -0.400 ;
        RECT -0.130 -0.690 0.100 -0.500 ;
        RECT 2.230 -0.570 2.490 -0.250 ;
        RECT 3.230 -0.310 3.500 -0.240 ;
        RECT 3.230 -0.560 3.600 -0.310 ;
        RECT 2.300 -1.040 2.490 -0.570 ;
        RECT 1.280 -1.480 1.600 -1.160 ;
        RECT 2.280 -1.330 2.510 -1.040 ;
        RECT 3.410 -1.050 3.600 -0.560 ;
        RECT 2.850 -1.480 3.170 -1.160 ;
        RECT 3.410 -1.340 3.640 -1.050 ;
      LAYER via ;
        RECT 1.310 4.320 1.570 4.580 ;
        RECT 2.880 4.320 3.140 4.580 ;
        RECT -0.040 3.340 0.220 3.600 ;
        RECT 2.230 3.410 2.490 3.670 ;
        RECT 3.240 3.400 3.500 3.660 ;
        RECT -0.040 2.730 0.220 2.990 ;
        RECT 2.230 2.660 2.490 2.920 ;
        RECT 3.240 2.670 3.500 2.930 ;
        RECT 1.310 1.750 1.570 2.010 ;
        RECT 2.880 1.750 3.140 2.010 ;
        RECT 1.310 1.120 1.570 1.380 ;
        RECT 2.880 1.120 3.140 1.380 ;
        RECT -0.040 0.140 0.220 0.400 ;
        RECT 2.230 0.210 2.490 0.470 ;
        RECT 3.240 0.200 3.500 0.460 ;
        RECT -0.040 -0.470 0.220 -0.210 ;
        RECT 2.230 -0.540 2.490 -0.280 ;
        RECT 3.240 -0.530 3.500 -0.270 ;
        RECT 1.310 -1.450 1.570 -1.190 ;
        RECT 2.880 -1.450 3.140 -1.190 ;
  END
END sky130_hilas_Tgate4Single01

MACRO sky130_hilas_swc4x1BiasCell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc4x1BiasCell ;
  ORIGIN 2.640 4.000 ;
  SIZE 10.080 BY 6.500 ;
  PIN ROW1
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 4.970 1.510 5.280 1.530 ;
        RECT -2.630 1.330 7.440 1.510 ;
        RECT -2.630 1.320 5.280 1.330 ;
        RECT 4.970 1.200 5.280 1.320 ;
    END
  END ROW1
  PIN ROW2
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 4.970 0.420 5.280 0.550 ;
        RECT -2.630 0.240 7.440 0.420 ;
        RECT 4.970 0.220 5.280 0.240 ;
    END
  END ROW2
  PIN ROW3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -2.630 -1.870 -2.160 -1.710 ;
        RECT -2.620 -1.880 -2.160 -1.870 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.970 -1.730 5.280 -1.710 ;
        RECT -1.860 -1.900 7.440 -1.730 ;
        RECT 4.880 -1.910 7.440 -1.900 ;
        RECT 4.970 -2.040 5.280 -1.910 ;
    END
  END ROW3
  PIN ROW4
    USE ANALOG ;
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT -2.630 -2.700 5.000 -2.690 ;
        RECT -2.630 -2.830 5.280 -2.700 ;
        RECT -2.630 -2.860 7.440 -2.830 ;
        RECT 4.880 -3.010 7.440 -2.860 ;
        RECT 4.970 -3.030 5.280 -3.010 ;
    END
  END ROW4
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 2.243500 ;
    PORT
      LAYER nwell ;
        RECT -2.630 -4.000 -0.900 2.500 ;
      LAYER met1 ;
        RECT -2.280 -4.000 -1.880 2.500 ;
    END
  END VTUN
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 3.253900 ;
    PORT
      LAYER nwell ;
        RECT 1.120 -4.000 3.350 2.490 ;
      LAYER met1 ;
        RECT 1.770 0.310 2.150 2.500 ;
        RECT 1.760 -1.550 2.150 0.310 ;
        RECT 1.770 -4.000 2.150 -1.550 ;
    END
  END GATE1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 4.880 -4.000 7.440 2.500 ;
      LAYER met1 ;
        RECT 6.920 1.790 7.080 2.490 ;
        RECT 6.810 1.240 7.080 1.790 ;
        RECT 6.810 1.190 7.090 1.240 ;
        RECT 6.920 1.100 7.090 1.190 ;
        RECT 6.920 0.650 7.080 1.100 ;
        RECT 6.920 0.560 7.090 0.650 ;
        RECT 6.810 0.510 7.090 0.560 ;
        RECT 6.810 -0.040 7.080 0.510 ;
        RECT 6.920 -1.450 7.080 -0.040 ;
        RECT 6.810 -2.000 7.080 -1.450 ;
        RECT 6.810 -2.050 7.090 -2.000 ;
        RECT 6.920 -2.140 7.090 -2.050 ;
        RECT 6.920 -2.600 7.080 -2.140 ;
        RECT 6.920 -2.690 7.090 -2.600 ;
        RECT 6.810 -2.740 7.090 -2.690 ;
        RECT 6.810 -3.290 7.080 -2.740 ;
        RECT 6.920 -3.990 7.080 -3.290 ;
    END
  END VINJ
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 6.110 1.760 6.270 2.490 ;
        RECT 6.110 1.740 6.310 1.760 ;
        RECT 6.090 1.500 6.320 1.740 ;
        RECT 6.110 1.450 6.320 1.500 ;
        RECT 6.480 1.450 6.670 2.440 ;
        RECT 6.110 0.300 6.270 1.450 ;
        RECT 6.500 1.330 6.670 1.450 ;
        RECT 6.510 0.420 6.670 1.330 ;
        RECT 6.500 0.300 6.670 0.420 ;
        RECT 6.110 0.250 6.320 0.300 ;
        RECT 6.090 0.010 6.320 0.250 ;
        RECT 6.110 -0.010 6.310 0.010 ;
        RECT 6.110 -0.650 6.270 -0.010 ;
        RECT 6.480 -0.620 6.670 0.300 ;
        RECT 6.460 -0.650 6.700 -0.620 ;
        RECT 6.110 -0.820 6.700 -0.650 ;
        RECT 6.110 -1.480 6.270 -0.820 ;
        RECT 6.460 -0.850 6.700 -0.820 ;
        RECT 6.110 -1.500 6.310 -1.480 ;
        RECT 6.090 -1.740 6.320 -1.500 ;
        RECT 6.110 -1.790 6.320 -1.740 ;
        RECT 6.480 -1.790 6.670 -0.850 ;
        RECT 6.110 -2.950 6.270 -1.790 ;
        RECT 6.500 -1.910 6.670 -1.790 ;
        RECT 6.510 -2.830 6.670 -1.910 ;
        RECT 6.500 -2.950 6.670 -2.830 ;
        RECT 6.110 -3.000 6.320 -2.950 ;
        RECT 6.090 -3.240 6.320 -3.000 ;
        RECT 6.110 -3.260 6.310 -3.240 ;
        RECT 6.110 -3.990 6.270 -3.260 ;
        RECT 6.480 -3.940 6.670 -2.950 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT -0.100 -2.300 0.230 -2.270 ;
        RECT 3.930 -2.300 4.250 -2.240 ;
        RECT -0.100 -2.470 4.250 -2.300 ;
        RECT -0.100 -2.530 0.230 -2.470 ;
        RECT 3.930 -2.520 4.250 -2.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.960 -2.210 4.210 2.500 ;
        RECT 3.950 -2.240 4.230 -2.210 ;
        RECT 3.940 -2.520 4.240 -2.240 ;
        RECT 3.950 -2.540 4.230 -2.520 ;
        RECT 3.960 -4.000 4.210 -2.540 ;
      LAYER via ;
        RECT 3.960 -2.510 4.220 -2.250 ;
    END
    PORT
      LAYER met1 ;
        RECT -0.070 -2.240 0.200 2.500 ;
        RECT -0.090 -2.550 0.220 -2.240 ;
        RECT -0.070 -4.000 0.200 -2.550 ;
      LAYER via ;
        RECT -0.070 -2.530 0.200 -2.270 ;
    END
  END VGND
  PIN DRAIN3
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 4.970 -1.290 5.280 -1.160 ;
        RECT 4.850 -1.300 5.280 -1.290 ;
        RECT 4.850 -1.460 7.440 -1.300 ;
        RECT 4.970 -1.480 7.440 -1.460 ;
        RECT 4.970 -1.490 5.280 -1.480 ;
    END
  END DRAIN3
  PIN DRAIN4
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 4.970 -3.260 5.280 -3.250 ;
        RECT 4.970 -3.440 7.440 -3.260 ;
        RECT 4.970 -3.580 5.280 -3.440 ;
    END
  END DRAIN4
  PIN DRAIN1
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 4.970 1.940 5.280 2.080 ;
        RECT 4.970 1.760 7.440 1.940 ;
        RECT 4.970 1.750 5.280 1.760 ;
    END
  END DRAIN1
  PIN DRAIN2
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 4.970 -0.010 5.280 0.000 ;
        RECT 4.970 -0.170 7.440 -0.010 ;
        RECT 4.880 -0.190 7.440 -0.170 ;
        RECT 4.880 -0.310 5.280 -0.190 ;
        RECT 4.970 -0.330 5.280 -0.310 ;
    END
  END DRAIN2
  OBS
      LAYER li1 ;
        RECT 4.980 2.030 5.300 2.040 ;
        RECT 4.980 1.860 5.560 2.030 ;
        RECT 4.980 1.810 5.310 1.860 ;
        RECT 4.980 1.780 5.300 1.810 ;
        RECT 6.840 1.760 7.040 2.110 ;
        RECT 4.980 1.450 5.300 1.490 ;
        RECT 4.980 1.410 5.310 1.450 ;
        RECT 4.980 1.240 5.560 1.410 ;
        RECT 4.980 1.230 5.300 1.240 ;
        RECT 6.110 1.140 6.310 1.740 ;
        RECT 6.840 1.730 7.050 1.760 ;
        RECT 6.830 1.140 7.050 1.730 ;
        RECT -0.020 0.480 0.150 1.010 ;
        RECT 4.000 0.450 4.170 0.980 ;
        RECT 4.980 0.510 5.300 0.520 ;
        RECT 4.980 0.340 5.560 0.510 ;
        RECT 4.980 0.300 5.310 0.340 ;
        RECT 4.980 0.260 5.300 0.300 ;
        RECT 6.110 0.010 6.310 0.610 ;
        RECT 6.830 0.020 7.050 0.610 ;
        RECT 6.840 -0.010 7.050 0.020 ;
        RECT 4.980 -0.060 5.300 -0.030 ;
        RECT 4.980 -0.110 5.310 -0.060 ;
        RECT -2.210 -1.020 -1.660 -0.590 ;
        RECT -0.010 -1.450 0.160 -0.280 ;
        RECT 1.820 -1.090 2.370 -0.660 ;
        RECT 4.010 -1.410 4.180 -0.220 ;
        RECT 4.980 -0.280 5.560 -0.110 ;
        RECT 4.980 -0.290 5.300 -0.280 ;
        RECT 6.840 -0.360 7.040 -0.010 ;
        RECT 6.230 -0.820 6.670 -0.650 ;
        RECT 4.980 -1.210 5.300 -1.200 ;
        RECT 4.980 -1.380 5.560 -1.210 ;
        RECT 4.980 -1.430 5.310 -1.380 ;
        RECT 4.980 -1.460 5.300 -1.430 ;
        RECT 6.840 -1.480 7.040 -1.130 ;
        RECT 4.980 -1.790 5.300 -1.750 ;
        RECT 4.980 -1.830 5.310 -1.790 ;
        RECT 4.980 -2.000 5.560 -1.830 ;
        RECT 4.980 -2.010 5.300 -2.000 ;
        RECT 6.110 -2.100 6.310 -1.500 ;
        RECT 6.840 -1.510 7.050 -1.480 ;
        RECT 6.830 -2.100 7.050 -1.510 ;
        RECT 4.980 -2.740 5.300 -2.730 ;
        RECT 4.980 -2.910 5.560 -2.740 ;
        RECT 4.980 -2.950 5.310 -2.910 ;
        RECT 4.980 -2.990 5.300 -2.950 ;
        RECT 6.110 -3.240 6.310 -2.640 ;
        RECT 6.830 -3.230 7.050 -2.640 ;
        RECT 6.840 -3.260 7.050 -3.230 ;
        RECT 4.980 -3.310 5.300 -3.280 ;
        RECT 4.980 -3.360 5.310 -3.310 ;
        RECT 4.980 -3.530 5.560 -3.360 ;
        RECT 4.980 -3.540 5.300 -3.530 ;
        RECT 6.840 -3.610 7.040 -3.260 ;
      LAYER mcon ;
        RECT 5.040 1.820 5.210 1.990 ;
        RECT 6.120 1.530 6.290 1.700 ;
        RECT 5.040 1.270 5.210 1.440 ;
        RECT 6.850 1.560 7.020 1.730 ;
        RECT -0.020 0.840 0.150 1.010 ;
        RECT 4.000 0.810 4.170 0.980 ;
        RECT 5.040 0.310 5.210 0.480 ;
        RECT 6.120 0.050 6.290 0.220 ;
        RECT 6.850 0.020 7.020 0.190 ;
        RECT -0.010 -0.450 0.160 -0.280 ;
        RECT -2.210 -0.940 -1.940 -0.670 ;
        RECT 4.010 -0.390 4.180 -0.220 ;
        RECT 5.040 -0.240 5.210 -0.070 ;
        RECT -0.010 -1.090 0.160 -0.920 ;
        RECT 1.820 -1.010 2.090 -0.740 ;
        RECT 6.490 -0.820 6.670 -0.650 ;
        RECT 4.010 -1.050 4.180 -0.880 ;
        RECT 5.040 -1.420 5.210 -1.250 ;
        RECT 6.120 -1.710 6.290 -1.540 ;
        RECT 5.040 -1.970 5.210 -1.800 ;
        RECT 6.850 -1.680 7.020 -1.510 ;
        RECT 5.040 -2.940 5.210 -2.770 ;
        RECT 6.120 -3.200 6.290 -3.030 ;
        RECT 6.850 -3.230 7.020 -3.060 ;
        RECT 5.040 -3.490 5.210 -3.320 ;
      LAYER met1 ;
        RECT 4.970 1.750 5.290 2.070 ;
        RECT 4.970 1.200 5.290 1.520 ;
        RECT 4.970 0.230 5.290 0.550 ;
        RECT 4.970 -0.320 5.290 0.000 ;
        RECT 4.970 -1.490 5.290 -1.170 ;
        RECT 4.970 -2.040 5.290 -1.720 ;
        RECT 4.970 -3.020 5.290 -2.700 ;
        RECT 4.970 -3.570 5.290 -3.250 ;
      LAYER via ;
        RECT 5.000 1.780 5.260 2.040 ;
        RECT 5.000 1.230 5.260 1.490 ;
        RECT 5.000 0.260 5.260 0.520 ;
        RECT 5.000 -0.290 5.260 -0.030 ;
        RECT 5.000 -1.460 5.260 -1.200 ;
        RECT 5.000 -2.010 5.260 -1.750 ;
        RECT 5.000 -2.990 5.260 -2.730 ;
        RECT 5.000 -3.540 5.260 -3.280 ;
  END
END sky130_hilas_swc4x1BiasCell

MACRO sky130_hilas_capacitorSize03
  CLASS BLOCK ;
  FOREIGN sky130_hilas_capacitorSize03 ;
  ORIGIN -14.140 0.470 ;
  SIZE 5.790 BY 5.870 ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 19.100 2.160 19.760 2.820 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 16.710 4.060 17.160 4.070 ;
        RECT 16.690 3.570 17.210 4.060 ;
        RECT 14.250 2.720 14.910 2.780 ;
        RECT 16.720 2.730 17.160 3.570 ;
        RECT 15.300 2.720 16.310 2.730 ;
        RECT 16.710 2.720 17.170 2.730 ;
        RECT 14.250 2.220 17.170 2.720 ;
        RECT 14.250 2.210 15.660 2.220 ;
        RECT 14.250 2.120 14.910 2.210 ;
        RECT 16.710 1.560 17.170 2.220 ;
        RECT 16.710 1.050 17.190 1.560 ;
        RECT 16.690 0.560 17.210 1.050 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 14.140 4.800 19.920 4.980 ;
        RECT 14.140 4.370 19.920 4.550 ;
        RECT 14.170 3.370 19.920 3.550 ;
        RECT 14.170 2.940 19.920 3.120 ;
        RECT 14.380 2.600 14.750 2.660 ;
        RECT 14.160 2.320 14.750 2.600 ;
        RECT 14.380 2.260 14.750 2.320 ;
        RECT 19.230 2.640 19.600 2.700 ;
        RECT 19.230 2.360 19.930 2.640 ;
        RECT 19.230 2.300 19.600 2.360 ;
        RECT 14.170 1.790 19.920 1.960 ;
        RECT 14.170 1.370 19.920 1.540 ;
        RECT 14.170 0.390 19.920 0.560 ;
        RECT 14.170 -0.050 19.920 0.120 ;
      LAYER via2 ;
        RECT 14.430 2.320 14.710 2.600 ;
        RECT 19.280 2.360 19.560 2.640 ;
      LAYER met3 ;
        RECT 15.590 2.850 18.430 5.400 ;
        RECT 14.160 2.060 14.950 2.810 ;
        RECT 15.590 2.100 19.800 2.850 ;
        RECT 15.590 -0.470 18.430 2.100 ;
      LAYER via3 ;
        RECT 14.350 2.210 14.780 2.690 ;
        RECT 19.200 2.250 19.630 2.730 ;
  END
END sky130_hilas_capacitorSize03

MACRO sky130_hilas_FGtrans2x1cell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_FGtrans2x1cell ;
  ORIGIN 3.950 3.870 ;
  SIZE 11.520 BY 6.150 ;
  PIN COLSEL1
    USE ANALOG ;
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT 6.610 0.770 6.800 2.230 ;
        RECT 6.610 0.740 6.830 0.770 ;
        RECT 6.590 0.470 6.840 0.740 ;
        RECT 6.600 0.460 6.840 0.470 ;
        RECT 6.600 0.220 6.830 0.460 ;
        RECT 6.640 -1.810 6.800 0.220 ;
        RECT 6.600 -2.050 6.830 -1.810 ;
        RECT 6.600 -2.060 6.840 -2.050 ;
        RECT 6.590 -2.330 6.840 -2.060 ;
        RECT 6.610 -2.360 6.830 -2.330 ;
        RECT 6.610 -3.820 6.800 -2.360 ;
    END
  END COLSEL1
  PIN VINJ
    USE ANALOG ;
    ANTENNADIFFAREA 0.544000 ;
    PORT
      LAYER nwell ;
        RECT 4.260 -3.870 7.570 2.280 ;
      LAYER met1 ;
        RECT 7.050 1.580 7.210 2.230 ;
        RECT 6.940 1.030 7.210 1.580 ;
        RECT 6.940 0.980 7.220 1.030 ;
        RECT 7.050 0.890 7.220 0.980 ;
        RECT 7.050 -2.480 7.210 0.890 ;
        RECT 7.050 -2.570 7.220 -2.480 ;
        RECT 6.940 -2.620 7.220 -2.570 ;
        RECT 6.940 -3.170 7.210 -2.620 ;
        RECT 7.050 -3.820 7.210 -3.170 ;
    END
  END VINJ
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 4.840 1.740 5.160 1.750 ;
        RECT 4.840 1.730 5.400 1.740 ;
        RECT -3.950 1.550 7.570 1.730 ;
        RECT 5.090 1.410 5.400 1.550 ;
    END
  END DRAIN1
  PIN DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 5.090 -3.140 5.400 -3.000 ;
        RECT 5.090 -3.150 7.570 -3.140 ;
        RECT -3.950 -3.300 7.570 -3.150 ;
        RECT 5.090 -3.320 7.570 -3.300 ;
        RECT 5.090 -3.330 5.400 -3.320 ;
    END
  END DRAIN2
  PIN PROG
    USE ANALOG ;
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER met1 ;
        RECT 3.840 -0.490 4.050 2.230 ;
        RECT 3.840 -1.000 4.080 -0.490 ;
        RECT 3.840 -3.820 4.050 -1.000 ;
    END
  END PROG
  PIN RUN
    USE ANALOG ;
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER met1 ;
        RECT 2.790 -2.300 2.970 2.230 ;
        RECT 2.740 -2.640 3.030 -2.300 ;
        RECT 2.790 -3.820 2.970 -2.640 ;
    END
  END RUN
  PIN VIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.217200 ;
    PORT
      LAYER met1 ;
        RECT 4.720 -1.200 4.910 -1.070 ;
        RECT 4.700 -1.490 4.930 -1.200 ;
        RECT 4.720 -3.110 4.910 -1.490 ;
        RECT 4.680 -3.320 4.910 -3.110 ;
        RECT 4.680 -3.400 4.920 -3.320 ;
        RECT 4.690 -3.820 4.920 -3.400 ;
    END
  END VIN2
  PIN VIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.217200 ;
    PORT
      LAYER met1 ;
        RECT 4.720 1.860 4.930 2.230 ;
        RECT 4.710 1.570 4.940 1.860 ;
        RECT 4.720 -0.130 4.930 1.570 ;
        RECT 4.710 -0.420 4.940 -0.130 ;
        RECT 4.720 -0.560 4.930 -0.420 ;
    END
  END VIN1
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 0.434600 ;
    PORT
      LAYER met1 ;
        RECT 4.270 1.300 4.460 2.230 ;
        RECT 4.240 1.010 4.470 1.300 ;
        RECT 4.270 -1.020 4.460 1.010 ;
        RECT 4.240 -1.310 4.470 -1.020 ;
        RECT 4.270 -2.600 4.460 -1.310 ;
        RECT 4.250 -2.890 4.480 -2.600 ;
        RECT 4.270 -3.820 4.460 -2.890 ;
    END
  END GATE1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT -1.130 -3.820 -0.900 2.230 ;
    END
  END VGND
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 2.516100 ;
    PORT
      LAYER nwell ;
        RECT -3.950 1.480 -2.220 2.230 ;
        RECT -3.950 0.330 -2.210 1.480 ;
        RECT -3.940 -1.910 -2.210 0.330 ;
        RECT -3.950 -2.090 -2.210 -1.910 ;
        RECT -3.950 -3.810 -2.220 -2.090 ;
      LAYER met1 ;
        RECT -3.610 -3.820 -3.190 2.230 ;
    END
  END VTUN
  PIN COL1
    ANTENNADIFFAREA 1.030400 ;
    PORT
      LAYER met2 ;
        RECT 6.190 -0.690 6.510 -0.660 ;
        RECT -3.950 -0.920 6.510 -0.690 ;
    END
  END COL1
  PIN ROW1
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 5.480 0.190 5.790 0.210 ;
        RECT -3.950 0.000 5.790 0.190 ;
        RECT 5.480 -0.120 5.790 0.000 ;
    END
  END ROW1
  PIN ROW2
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 5.490 -1.670 5.800 -1.480 ;
        RECT -3.950 -1.810 5.800 -1.670 ;
        RECT -3.950 -1.860 5.770 -1.810 ;
    END
  END ROW2
  OBS
      LAYER nwell ;
        RECT -0.190 -0.160 2.530 1.490 ;
        RECT -0.180 -0.200 2.530 -0.160 ;
        RECT -0.180 -1.530 2.530 -1.490 ;
        RECT -0.190 -3.180 2.530 -1.530 ;
      LAYER li1 ;
        RECT 4.730 1.800 4.920 1.830 ;
        RECT 3.860 1.630 4.920 1.800 ;
        RECT 5.160 1.650 5.690 1.820 ;
        RECT 3.860 1.240 4.030 1.630 ;
        RECT 4.730 1.600 4.920 1.630 ;
        RECT 6.970 1.550 7.170 1.900 ;
        RECT 6.970 1.520 7.180 1.550 ;
        RECT 3.290 1.070 4.030 1.240 ;
        RECT 4.260 1.240 4.450 1.270 ;
        RECT 4.260 1.070 4.990 1.240 ;
        RECT 4.260 1.040 4.450 1.070 ;
        RECT -3.520 0.090 -2.970 0.520 ;
        RECT 2.000 0.450 2.230 0.970 ;
        RECT 2.000 0.280 4.990 0.450 ;
        RECT 5.410 0.170 5.580 1.260 ;
        RECT 5.410 0.130 5.810 0.170 ;
        RECT 5.410 -0.060 5.820 0.130 ;
        RECT 5.410 -0.090 5.810 -0.060 ;
        RECT 4.730 -0.340 4.920 -0.160 ;
        RECT -0.920 -0.740 -0.730 -0.340 ;
        RECT 3.300 -0.510 3.640 -0.340 ;
        RECT -1.110 -0.750 -0.730 -0.740 ;
        RECT -1.110 -0.930 2.630 -0.750 ;
        RECT -1.110 -0.970 -0.730 -0.930 ;
        RECT -3.520 -1.640 -2.970 -1.210 ;
        RECT -0.920 -1.350 -0.730 -0.970 ;
        RECT 3.380 -1.080 3.550 -0.510 ;
        RECT 3.860 -0.920 4.070 -0.490 ;
        RECT 4.640 -0.510 4.990 -0.340 ;
        RECT 5.410 -0.430 5.580 -0.090 ;
        RECT 6.240 -0.340 6.410 1.270 ;
        RECT 6.960 0.940 7.180 1.520 ;
        RECT 6.970 0.930 7.180 0.940 ;
        RECT 6.610 0.760 6.800 0.770 ;
        RECT 6.610 0.470 6.810 0.760 ;
        RECT 6.600 0.140 6.870 0.470 ;
        RECT 6.240 -0.530 6.420 -0.340 ;
        RECT 3.880 -0.940 4.050 -0.920 ;
        RECT 3.300 -1.110 3.640 -1.080 ;
        RECT 4.260 -1.100 4.450 -1.050 ;
        RECT 4.220 -1.110 4.450 -1.100 ;
        RECT 3.300 -1.250 4.450 -1.110 ;
        RECT 4.640 -1.250 4.990 -1.080 ;
        RECT 3.470 -1.280 4.450 -1.250 ;
        RECT 3.470 -1.310 4.310 -1.280 ;
        RECT 4.720 -1.460 4.910 -1.250 ;
        RECT 5.410 -1.520 5.580 -1.160 ;
        RECT 6.240 -1.250 6.420 -1.060 ;
        RECT 5.410 -1.560 5.820 -1.520 ;
        RECT 5.410 -1.750 5.830 -1.560 ;
        RECT 5.410 -1.780 5.820 -1.750 ;
        RECT 2.060 -1.970 4.990 -1.870 ;
        RECT 2.000 -2.040 4.990 -1.970 ;
        RECT 2.000 -2.660 2.230 -2.040 ;
        RECT 2.800 -2.360 2.970 -2.300 ;
        RECT 2.780 -2.570 2.990 -2.360 ;
        RECT 2.800 -2.640 2.970 -2.570 ;
        RECT 4.270 -2.660 4.460 -2.630 ;
        RECT 3.290 -2.830 4.100 -2.660 ;
        RECT 3.910 -3.170 4.100 -2.830 ;
        RECT 4.270 -2.830 4.990 -2.660 ;
        RECT 4.270 -2.860 4.460 -2.830 ;
        RECT 5.410 -2.850 5.580 -1.780 ;
        RECT 6.240 -2.860 6.410 -1.250 ;
        RECT 6.600 -2.060 6.870 -1.730 ;
        RECT 6.610 -2.350 6.810 -2.060 ;
        RECT 6.610 -2.360 6.800 -2.350 ;
        RECT 6.970 -2.530 7.180 -2.520 ;
        RECT 6.960 -3.110 7.180 -2.530 ;
        RECT 6.970 -3.140 7.180 -3.110 ;
        RECT 4.700 -3.170 4.890 -3.140 ;
        RECT 3.910 -3.350 4.890 -3.170 ;
        RECT 4.700 -3.370 4.890 -3.350 ;
        RECT 5.160 -3.410 5.690 -3.240 ;
        RECT 6.970 -3.490 7.170 -3.140 ;
      LAYER mcon ;
        RECT 4.740 1.630 4.910 1.800 ;
        RECT 6.980 1.350 7.150 1.520 ;
        RECT 4.270 1.070 4.440 1.240 ;
        RECT 2.030 0.770 2.200 0.940 ;
        RECT -3.520 0.170 -3.250 0.440 ;
        RECT 2.030 0.320 2.200 0.490 ;
        RECT 5.550 -0.050 5.720 0.120 ;
        RECT 4.740 -0.360 4.910 -0.190 ;
        RECT -1.100 -0.940 -0.930 -0.770 ;
        RECT -3.520 -1.560 -3.250 -1.290 ;
        RECT 6.620 0.510 6.800 0.700 ;
        RECT 4.270 -1.250 4.440 -1.080 ;
        RECT 4.730 -1.430 4.900 -1.260 ;
        RECT 5.560 -1.740 5.730 -1.570 ;
        RECT 2.030 -2.180 2.200 -2.010 ;
        RECT 2.030 -2.630 2.200 -2.460 ;
        RECT 4.280 -2.830 4.450 -2.660 ;
        RECT 6.620 -2.290 6.800 -2.100 ;
        RECT 6.980 -3.110 7.150 -2.940 ;
        RECT 4.710 -3.340 4.880 -3.170 ;
      LAYER met1 ;
        RECT 5.090 1.410 5.400 1.850 ;
        RECT 1.990 0.230 2.250 1.020 ;
        RECT 5.480 -0.120 5.800 0.200 ;
        RECT 6.210 -0.630 6.450 -0.210 ;
        RECT 6.210 -0.950 6.480 -0.630 ;
        RECT 6.210 -1.380 6.450 -0.950 ;
        RECT 5.490 -1.810 5.810 -1.490 ;
        RECT 1.990 -2.710 2.250 -1.920 ;
        RECT 5.090 -3.440 5.400 -3.000 ;
      LAYER via ;
        RECT 5.120 1.440 5.380 1.700 ;
        RECT 5.510 -0.090 5.770 0.170 ;
        RECT 6.220 -0.920 6.480 -0.660 ;
        RECT 5.520 -1.780 5.780 -1.520 ;
        RECT 5.120 -3.290 5.380 -3.030 ;
  END
END sky130_hilas_FGtrans2x1cell

MACRO sky130_hilas_WTA4Stage01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_WTA4Stage01 ;
  ORIGIN 11.210 0.610 ;
  SIZE 14.170 BY 6.500 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 2.510 1.160 2.840 1.250 ;
        RECT -7.420 1.090 -7.100 1.150 ;
        RECT -3.840 1.090 2.840 1.160 ;
        RECT -7.420 0.990 2.840 1.090 ;
        RECT -7.420 0.920 -3.070 0.990 ;
        RECT 2.510 0.960 2.840 0.990 ;
        RECT -7.420 0.870 -7.100 0.920 ;
        RECT -3.400 0.860 -3.070 0.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.570 1.270 2.800 5.620 ;
        RECT 2.530 1.260 2.810 1.270 ;
        RECT 2.530 0.940 2.830 1.260 ;
        RECT 2.570 -0.430 2.800 0.940 ;
      LAYER via ;
        RECT 2.540 0.970 2.810 1.240 ;
    END
  END VGND
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT -8.450 4.900 -8.140 4.920 ;
        RECT -0.650 4.900 -0.510 4.910 ;
        RECT -10.610 4.720 -0.500 4.900 ;
        RECT -8.450 4.710 -0.500 4.720 ;
        RECT -8.450 4.590 -8.140 4.710 ;
        RECT -0.650 4.570 -0.500 4.710 ;
        RECT -0.650 4.480 0.560 4.570 ;
        RECT -0.650 4.420 0.690 4.480 ;
        RECT -0.650 4.370 2.960 4.420 ;
        RECT 0.380 4.260 2.960 4.370 ;
        RECT 0.380 4.150 0.690 4.260 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT -8.450 3.810 -8.140 3.940 ;
        RECT -10.610 3.630 0.660 3.810 ;
        RECT -8.450 3.610 -8.140 3.630 ;
        RECT 0.380 3.600 0.660 3.630 ;
        RECT 0.380 3.490 0.690 3.600 ;
        RECT 0.380 3.330 2.960 3.490 ;
        RECT 0.380 3.270 0.690 3.330 ;
    END
  END OUTPUT2
  PIN OUTPUT3
    USE ANALOG ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 0.380 1.680 0.690 1.710 ;
        RECT -1.010 1.650 0.690 1.680 ;
        RECT -1.010 1.520 2.960 1.650 ;
        RECT -1.010 1.510 -0.550 1.520 ;
        RECT 0.380 1.490 2.960 1.520 ;
        RECT 0.380 1.380 0.690 1.490 ;
    END
  END OUTPUT3
  PIN OUTPUT4
    USE ANALOG ;
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 0.380 0.720 0.690 0.830 ;
        RECT 0.380 0.710 2.960 0.720 ;
        RECT -0.550 0.700 2.960 0.710 ;
        RECT -8.170 0.690 2.960 0.700 ;
        RECT -8.450 0.560 2.960 0.690 ;
        RECT -10.610 0.530 0.690 0.560 ;
        RECT -10.610 0.380 -8.050 0.530 ;
        RECT 0.380 0.500 0.690 0.530 ;
        RECT -8.450 0.360 -8.140 0.380 ;
    END
  END OUTPUT4
  PIN INPUT1
    USE ANALOG ;
    ANTENNAGATEAREA 0.118000 ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT -7.850 5.310 -7.530 5.330 ;
        RECT -7.850 5.120 0.070 5.310 ;
        RECT 0.230 5.120 0.540 5.160 ;
        RECT -7.850 5.100 0.540 5.120 ;
        RECT -7.850 5.070 -7.530 5.100 ;
        RECT -0.140 4.910 0.540 5.100 ;
        RECT 0.230 4.830 0.540 4.910 ;
        RECT -11.120 4.270 -10.970 4.690 ;
        RECT -7.870 4.270 -7.550 4.280 ;
        RECT -11.120 4.120 -7.550 4.270 ;
        RECT -7.990 4.020 -7.550 4.120 ;
    END
  END INPUT1
  PIN INPUT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.118000 ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT -11.140 3.520 -10.820 3.790 ;
        RECT -7.910 3.040 -7.680 3.050 ;
        RECT -7.910 3.010 -0.340 3.040 ;
        RECT -7.910 2.840 -0.280 3.010 ;
        RECT 0.230 2.840 0.540 2.920 ;
        RECT -11.160 2.740 -10.840 2.770 ;
        RECT -7.910 2.740 -7.670 2.840 ;
        RECT -11.160 2.560 -7.670 2.740 ;
        RECT -0.470 2.640 0.540 2.840 ;
        RECT 0.130 2.630 0.540 2.640 ;
        RECT 0.230 2.590 0.540 2.630 ;
        RECT -11.160 2.540 -7.750 2.560 ;
        RECT -11.160 2.510 -10.840 2.540 ;
    END
  END INPUT2
  PIN INPUT3
    USE ANALOG ;
    ANTENNAGATEAREA 0.118000 ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT -7.870 2.360 -7.550 2.400 ;
        RECT -7.870 2.340 -0.320 2.360 ;
        RECT 0.230 2.350 0.540 2.390 ;
        RECT 0.130 2.340 0.540 2.350 ;
        RECT -7.870 2.140 0.540 2.340 ;
        RECT -7.770 2.130 -7.450 2.140 ;
        RECT 0.230 2.060 0.540 2.140 ;
        RECT -11.180 1.180 -10.980 1.680 ;
        RECT -8.000 1.180 -7.680 1.220 ;
        RECT -11.180 0.980 -7.630 1.180 ;
        RECT -8.000 0.960 -7.680 0.980 ;
    END
  END INPUT3
  PIN INPUT4
    USE ANALOG ;
    ANTENNAGATEAREA 0.118000 ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT -11.210 0.440 -10.900 0.770 ;
        RECT 0.230 0.090 0.540 0.150 ;
        RECT -0.320 0.080 0.540 0.090 ;
        RECT -7.900 -0.140 0.540 0.080 ;
        RECT -7.900 -0.150 -0.310 -0.140 ;
        RECT -7.900 -0.160 -7.130 -0.150 ;
        RECT -11.160 -0.200 -10.850 -0.190 ;
        RECT -11.160 -0.330 -10.800 -0.200 ;
        RECT -7.900 -0.330 -7.660 -0.160 ;
        RECT 0.230 -0.180 0.540 -0.140 ;
        RECT -11.160 -0.520 -7.660 -0.330 ;
        RECT -11.030 -0.570 -7.660 -0.520 ;
    END
  END INPUT4
  PIN DRAIN1
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT -8.450 5.330 -8.140 5.470 ;
        RECT -11.160 5.150 -8.140 5.330 ;
        RECT -8.450 5.140 -8.140 5.150 ;
    END
  END DRAIN1
  PIN GATE1
    ANTENNADIFFAREA 3.253900 ;
    PORT
      LAYER nwell ;
        RECT -6.520 -0.610 -4.290 5.880 ;
      LAYER met1 ;
        RECT -5.320 3.700 -4.940 5.890 ;
        RECT -5.320 1.840 -4.930 3.700 ;
        RECT -5.320 -0.610 -4.940 1.840 ;
    END
  END GATE1
  PIN VTUN
    ANTENNADIFFAREA 2.243500 ;
    PORT
      LAYER nwell ;
        RECT -2.270 -0.610 -0.540 5.890 ;
      LAYER met1 ;
        RECT -1.290 -0.610 -0.890 5.890 ;
    END
  END VTUN
  PIN WTAMIDDLENODE
    ANTENNAGATEAREA 0.472000 ;
    ANTENNADIFFAREA 0.708000 ;
    PORT
      LAYER met1 ;
        RECT 1.310 -0.430 1.540 5.620 ;
    END
  END WTAMIDDLENODE
  PIN COLSEL1
    ANTENNAGATEAREA 0.720000 ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met1 ;
        RECT -9.840 4.840 -9.650 5.830 ;
        RECT -9.440 5.150 -9.280 5.880 ;
        RECT -9.480 5.130 -9.280 5.150 ;
        RECT -9.490 4.890 -9.260 5.130 ;
        RECT -9.490 4.840 -9.280 4.890 ;
        RECT -9.840 4.720 -9.670 4.840 ;
        RECT -9.840 3.810 -9.680 4.720 ;
        RECT -9.840 3.690 -9.670 3.810 ;
        RECT -9.440 3.690 -9.280 4.840 ;
        RECT -9.840 2.770 -9.650 3.690 ;
        RECT -9.490 3.640 -9.280 3.690 ;
        RECT -9.490 3.400 -9.260 3.640 ;
        RECT -9.480 3.380 -9.280 3.400 ;
        RECT -9.870 2.740 -9.630 2.770 ;
        RECT -9.440 2.740 -9.280 3.380 ;
        RECT -9.870 2.570 -9.280 2.740 ;
        RECT -9.870 2.540 -9.630 2.570 ;
        RECT -9.840 1.600 -9.650 2.540 ;
        RECT -9.440 1.910 -9.280 2.570 ;
        RECT -9.480 1.890 -9.280 1.910 ;
        RECT -9.490 1.650 -9.260 1.890 ;
        RECT -9.490 1.600 -9.280 1.650 ;
        RECT -9.840 1.480 -9.670 1.600 ;
        RECT -9.840 0.560 -9.680 1.480 ;
        RECT -9.840 0.440 -9.670 0.560 ;
        RECT -9.440 0.440 -9.280 1.600 ;
        RECT -9.840 -0.550 -9.650 0.440 ;
        RECT -9.490 0.390 -9.280 0.440 ;
        RECT -9.490 0.150 -9.260 0.390 ;
        RECT -9.480 0.130 -9.280 0.150 ;
        RECT -9.440 -0.600 -9.280 0.130 ;
    END
  END COLSEL1
  PIN VINJ
    ANTENNADIFFAREA 1.088000 ;
    PORT
      LAYER nwell ;
        RECT -10.610 5.620 -8.050 5.890 ;
        RECT -11.010 3.690 -8.050 5.620 ;
        RECT -11.120 2.540 -8.050 3.690 ;
        RECT -11.010 -0.420 -8.050 2.540 ;
        RECT -10.610 -0.610 -8.050 -0.420 ;
      LAYER met1 ;
        RECT -10.250 5.180 -10.090 5.880 ;
        RECT -10.250 4.630 -9.980 5.180 ;
        RECT -10.260 4.580 -9.980 4.630 ;
        RECT -10.260 4.490 -10.090 4.580 ;
        RECT -10.250 4.040 -10.090 4.490 ;
        RECT -10.260 3.950 -10.090 4.040 ;
        RECT -10.260 3.900 -9.980 3.950 ;
        RECT -10.250 3.350 -9.980 3.900 ;
        RECT -10.250 1.940 -10.090 3.350 ;
        RECT -10.250 1.390 -9.980 1.940 ;
        RECT -10.260 1.340 -9.980 1.390 ;
        RECT -10.260 1.250 -10.090 1.340 ;
        RECT -10.250 0.790 -10.090 1.250 ;
        RECT -10.260 0.700 -10.090 0.790 ;
        RECT -10.260 0.650 -9.980 0.700 ;
        RECT -10.250 0.100 -9.980 0.650 ;
        RECT -10.250 -0.600 -10.090 0.100 ;
    END
  END VINJ
  PIN DRAIN2
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT -8.450 3.380 -8.140 3.390 ;
        RECT -11.190 3.220 -8.140 3.380 ;
        RECT -11.190 3.200 -8.050 3.220 ;
        RECT -8.450 3.080 -8.050 3.200 ;
        RECT -8.450 3.060 -8.140 3.080 ;
    END
  END DRAIN2
  PIN DRAIN3
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT -8.450 2.100 -8.140 2.230 ;
        RECT -8.450 2.090 -8.020 2.100 ;
        RECT -11.160 1.930 -8.020 2.090 ;
        RECT -11.160 1.910 -8.140 1.930 ;
        RECT -8.450 1.900 -8.140 1.910 ;
    END
  END DRAIN3
  PIN DRAIN4
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT -8.450 0.130 -8.140 0.140 ;
        RECT -11.180 -0.050 -8.140 0.130 ;
        RECT -8.450 -0.190 -8.140 -0.050 ;
    END
  END DRAIN4
  OBS
      LAYER li1 ;
        RECT -10.210 5.150 -10.010 5.500 ;
        RECT -8.470 5.420 -8.150 5.430 ;
        RECT -8.730 5.250 -8.150 5.420 ;
        RECT -8.480 5.200 -8.150 5.250 ;
        RECT -8.470 5.170 -8.150 5.200 ;
        RECT -10.220 5.120 -10.010 5.150 ;
        RECT -10.220 4.530 -10.000 5.120 ;
        RECT -9.480 4.530 -9.280 5.130 ;
        RECT 0.240 5.100 0.560 5.130 ;
        RECT 0.240 4.930 2.030 5.100 ;
        RECT 0.240 4.910 0.570 4.930 ;
        RECT -8.470 4.840 -8.150 4.880 ;
        RECT 0.240 4.870 0.560 4.910 ;
        RECT -8.480 4.800 -8.150 4.840 ;
        RECT -8.730 4.630 -8.150 4.800 ;
        RECT 1.860 4.700 2.030 4.930 ;
        RECT -8.470 4.620 -8.150 4.630 ;
        RECT 0.710 4.450 1.050 4.700 ;
        RECT 1.220 4.530 1.550 4.700 ;
        RECT 1.770 4.530 2.110 4.700 ;
        RECT -10.220 3.410 -10.000 4.000 ;
        RECT -10.220 3.380 -10.010 3.410 ;
        RECT -9.480 3.400 -9.280 4.000 ;
        RECT -8.470 3.900 -8.150 3.910 ;
        RECT -8.730 3.730 -8.150 3.900 ;
        RECT -7.340 3.840 -7.170 4.370 ;
        RECT -3.320 3.870 -3.150 4.400 ;
        RECT 0.390 4.190 1.050 4.450 ;
        RECT 1.300 4.360 1.470 4.530 ;
        RECT 1.860 4.360 2.030 4.530 ;
        RECT 1.220 4.190 1.550 4.360 ;
        RECT 1.770 4.190 2.110 4.360 ;
        RECT 1.300 3.960 1.550 4.190 ;
        RECT 2.430 4.110 2.940 4.780 ;
        RECT -8.480 3.690 -8.150 3.730 ;
        RECT -8.470 3.650 -8.150 3.690 ;
        RECT 1.300 3.790 1.970 3.960 ;
        RECT 1.300 3.560 1.550 3.790 ;
        RECT -10.210 3.030 -10.010 3.380 ;
        RECT -8.470 3.330 -8.150 3.360 ;
        RECT -8.480 3.280 -8.150 3.330 ;
        RECT 0.390 3.300 1.050 3.560 ;
        RECT 1.220 3.390 1.550 3.560 ;
        RECT 1.770 3.390 2.110 3.560 ;
        RECT -8.730 3.110 -8.150 3.280 ;
        RECT -8.470 3.100 -8.150 3.110 ;
        RECT -9.840 2.570 -9.400 2.740 ;
        RECT -10.210 1.910 -10.010 2.260 ;
        RECT -8.470 2.180 -8.150 2.190 ;
        RECT -8.730 2.010 -8.150 2.180 ;
        RECT -8.480 1.960 -8.150 2.010 ;
        RECT -7.350 1.980 -7.180 3.170 ;
        RECT -5.540 2.300 -4.990 2.730 ;
        RECT -8.470 1.930 -8.150 1.960 ;
        RECT -3.330 1.940 -3.160 3.110 ;
        RECT 0.710 3.050 1.050 3.300 ;
        RECT 1.300 3.220 1.470 3.390 ;
        RECT 1.860 3.220 2.030 3.390 ;
        RECT 1.220 3.050 1.550 3.220 ;
        RECT 1.770 3.050 2.110 3.220 ;
        RECT 0.240 2.840 0.560 2.880 ;
        RECT 0.240 2.820 0.570 2.840 ;
        RECT 1.860 2.820 2.030 3.050 ;
        RECT 2.430 2.970 2.940 3.640 ;
        RECT -1.510 2.370 -0.960 2.800 ;
        RECT 0.240 2.650 2.030 2.820 ;
        RECT 0.240 2.620 0.560 2.650 ;
        RECT 0.240 2.330 0.560 2.360 ;
        RECT 0.240 2.160 2.030 2.330 ;
        RECT 0.240 2.140 0.570 2.160 ;
        RECT 0.240 2.100 0.560 2.140 ;
        RECT 1.860 1.930 2.030 2.160 ;
        RECT -10.220 1.880 -10.010 1.910 ;
        RECT -10.220 1.290 -10.000 1.880 ;
        RECT -9.480 1.290 -9.280 1.890 ;
        RECT 0.710 1.680 1.050 1.930 ;
        RECT 1.220 1.760 1.550 1.930 ;
        RECT 1.770 1.760 2.110 1.930 ;
        RECT -8.470 1.600 -8.150 1.640 ;
        RECT -8.480 1.560 -8.150 1.600 ;
        RECT -8.730 1.390 -8.150 1.560 ;
        RECT 0.390 1.420 1.050 1.680 ;
        RECT 1.300 1.590 1.470 1.760 ;
        RECT 1.860 1.590 2.030 1.760 ;
        RECT 1.220 1.420 1.550 1.590 ;
        RECT 1.770 1.420 2.110 1.590 ;
        RECT -8.470 1.380 -8.150 1.390 ;
        RECT 1.300 1.190 1.550 1.420 ;
        RECT 2.430 1.340 2.940 2.010 ;
        RECT 1.300 1.020 1.970 1.190 ;
        RECT 1.300 0.790 1.550 1.020 ;
        RECT -11.200 0.690 -10.880 0.730 ;
        RECT -11.200 0.500 -10.870 0.690 ;
        RECT -11.200 0.470 -10.880 0.500 ;
        RECT -11.150 -0.230 -10.970 0.470 ;
        RECT -10.220 0.160 -10.000 0.750 ;
        RECT -10.220 0.130 -10.010 0.160 ;
        RECT -9.480 0.150 -9.280 0.750 ;
        RECT -8.470 0.650 -8.150 0.660 ;
        RECT -8.730 0.480 -8.150 0.650 ;
        RECT 0.390 0.530 1.050 0.790 ;
        RECT 1.220 0.620 1.550 0.790 ;
        RECT 1.770 0.620 2.110 0.790 ;
        RECT -8.480 0.440 -8.150 0.480 ;
        RECT -8.470 0.400 -8.150 0.440 ;
        RECT 0.710 0.280 1.050 0.530 ;
        RECT 1.300 0.450 1.470 0.620 ;
        RECT 1.860 0.450 2.030 0.620 ;
        RECT 1.220 0.280 1.550 0.450 ;
        RECT 1.770 0.280 2.110 0.450 ;
        RECT -10.210 -0.220 -10.010 0.130 ;
        RECT -8.470 0.080 -8.150 0.110 ;
        RECT -8.480 0.030 -8.150 0.080 ;
        RECT -8.730 -0.140 -8.150 0.030 ;
        RECT -8.470 -0.150 -8.150 -0.140 ;
        RECT 0.240 0.070 0.560 0.110 ;
        RECT 0.240 0.050 0.570 0.070 ;
        RECT 1.860 0.050 2.030 0.280 ;
        RECT 2.430 0.200 2.940 0.870 ;
        RECT 0.240 -0.120 2.030 0.050 ;
        RECT 0.240 -0.150 0.560 -0.120 ;
        RECT -11.150 -0.270 -10.830 -0.230 ;
        RECT -11.150 -0.460 -10.820 -0.270 ;
        RECT -11.150 -0.490 -10.830 -0.460 ;
      LAYER mcon ;
        RECT -8.380 5.210 -8.210 5.380 ;
        RECT -10.190 4.950 -10.020 5.120 ;
        RECT -9.460 4.920 -9.290 5.090 ;
        RECT 0.300 4.920 0.470 5.090 ;
        RECT -8.380 4.660 -8.210 4.830 ;
        RECT -7.340 4.200 -7.170 4.370 ;
        RECT -10.190 3.410 -10.020 3.580 ;
        RECT -8.380 3.700 -8.210 3.870 ;
        RECT -3.320 4.230 -3.150 4.400 ;
        RECT 0.450 4.240 0.620 4.410 ;
        RECT 2.600 4.360 2.770 4.530 ;
        RECT 1.340 3.790 1.510 3.960 ;
        RECT -9.460 3.440 -9.290 3.610 ;
        RECT -8.380 3.150 -8.210 3.320 ;
        RECT 0.450 3.340 0.620 3.510 ;
        RECT -7.350 3.000 -7.180 3.170 ;
        RECT -3.330 2.940 -3.160 3.110 ;
        RECT 2.600 3.220 2.770 3.390 ;
        RECT -7.350 2.340 -7.180 2.510 ;
        RECT -8.380 1.970 -8.210 2.140 ;
        RECT -5.260 2.380 -4.990 2.650 ;
        RECT -3.330 2.300 -3.160 2.470 ;
        RECT -1.230 2.450 -0.960 2.720 ;
        RECT 0.300 2.660 0.470 2.830 ;
        RECT 0.300 2.150 0.470 2.320 ;
        RECT -10.190 1.710 -10.020 1.880 ;
        RECT -9.460 1.680 -9.290 1.850 ;
        RECT -8.380 1.420 -8.210 1.590 ;
        RECT 0.450 1.470 0.620 1.640 ;
        RECT 2.600 1.590 2.770 1.760 ;
        RECT 1.340 1.020 1.510 1.190 ;
        RECT -11.140 0.510 -10.970 0.680 ;
        RECT -10.190 0.160 -10.020 0.330 ;
        RECT -8.380 0.450 -8.210 0.620 ;
        RECT 0.450 0.570 0.620 0.740 ;
        RECT -9.460 0.190 -9.290 0.360 ;
        RECT 2.600 0.450 2.770 0.620 ;
        RECT -8.380 -0.100 -8.210 0.070 ;
        RECT 0.300 -0.110 0.470 0.060 ;
        RECT -11.090 -0.450 -10.920 -0.280 ;
      LAYER met1 ;
        RECT -8.460 5.140 -8.140 5.460 ;
        RECT -7.820 5.040 -7.560 5.360 ;
        RECT -8.460 4.590 -8.140 4.910 ;
        RECT -7.820 4.310 -7.610 5.040 ;
        RECT -7.840 3.990 -7.580 4.310 ;
        RECT -11.110 3.690 -10.850 3.810 ;
        RECT -11.120 3.490 -10.850 3.690 ;
        RECT -8.460 3.620 -8.140 3.940 ;
        RECT -11.120 2.800 -10.910 3.490 ;
        RECT -8.460 3.070 -8.140 3.390 ;
        RECT -11.130 2.480 -10.870 2.800 ;
        RECT -8.460 1.900 -8.140 2.220 ;
        RECT -7.840 2.110 -7.580 2.430 ;
        RECT -8.460 1.350 -8.140 1.670 ;
        RECT -7.840 1.250 -7.680 2.110 ;
        RECT -7.970 0.930 -7.680 1.250 ;
        RECT -7.380 1.180 -7.130 5.890 ;
        RECT -7.400 1.150 -7.120 1.180 ;
        RECT -3.370 1.150 -3.100 5.890 ;
        RECT 0.230 4.840 0.550 5.160 ;
        RECT 0.380 4.160 0.700 4.480 ;
        RECT 0.380 3.270 0.700 3.590 ;
        RECT 0.230 2.590 0.550 2.910 ;
        RECT 0.230 2.070 0.550 2.390 ;
        RECT 0.380 1.390 0.700 1.710 ;
        RECT -7.410 0.870 -7.110 1.150 ;
        RECT -7.400 0.850 -7.120 0.870 ;
        RECT -11.210 0.440 -10.890 0.760 ;
        RECT -8.460 0.370 -8.140 0.690 ;
        RECT -8.460 -0.180 -8.140 0.140 ;
        RECT -11.160 -0.520 -10.840 -0.200 ;
        RECT -7.380 -0.610 -7.130 0.850 ;
        RECT -3.390 0.840 -3.080 1.150 ;
        RECT -3.370 -0.610 -3.100 0.840 ;
        RECT 0.380 0.500 0.700 0.820 ;
        RECT 0.230 -0.180 0.550 0.140 ;
      LAYER via ;
        RECT -8.430 5.170 -8.170 5.430 ;
        RECT -7.820 5.070 -7.560 5.330 ;
        RECT -8.430 4.620 -8.170 4.880 ;
        RECT -7.840 4.020 -7.580 4.280 ;
        RECT -11.110 3.520 -10.850 3.780 ;
        RECT -8.430 3.650 -8.170 3.910 ;
        RECT -8.430 3.100 -8.170 3.360 ;
        RECT -11.130 2.510 -10.870 2.770 ;
        RECT -8.430 1.930 -8.170 2.190 ;
        RECT -7.840 2.140 -7.580 2.400 ;
        RECT -8.430 1.380 -8.170 1.640 ;
        RECT -7.970 0.960 -7.710 1.220 ;
        RECT 0.260 4.870 0.520 5.130 ;
        RECT 0.410 4.190 0.670 4.450 ;
        RECT 0.410 3.300 0.670 3.560 ;
        RECT 0.260 2.620 0.520 2.880 ;
        RECT 0.260 2.100 0.520 2.360 ;
        RECT 0.410 1.420 0.670 1.680 ;
        RECT -7.390 0.880 -7.130 1.140 ;
        RECT -3.370 0.860 -3.100 1.120 ;
        RECT -11.180 0.470 -10.920 0.730 ;
        RECT -8.430 0.400 -8.170 0.660 ;
        RECT -8.430 -0.150 -8.170 0.110 ;
        RECT -11.130 -0.490 -10.870 -0.230 ;
        RECT 0.410 0.530 0.670 0.790 ;
        RECT 0.260 -0.150 0.520 0.110 ;
      LAYER met2 ;
        RECT -8.450 1.660 -8.140 1.680 ;
        RECT -10.610 1.490 -1.310 1.660 ;
        RECT -10.610 1.480 -8.050 1.490 ;
        RECT -8.450 1.350 -8.140 1.480 ;
  END
END sky130_hilas_WTA4Stage01

MACRO sky130_hilas_TopProtectStructure
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TopProtectStructure ;
  ORIGIN 154.680 243.370 ;
  SIZE 372.850 BY 389.100 ;
  PIN IO07
    PORT
      LAYER met1 ;
        RECT 215.620 -58.690 216.210 -58.680 ;
        RECT 215.620 -62.290 218.170 -58.690 ;
        RECT 214.270 -62.580 218.170 -62.290 ;
    END
  END IO07
  PIN IO08
    PORT
      LAYER met1 ;
        RECT 216.920 -30.090 218.170 -30.080 ;
        RECT 215.620 -33.700 218.170 -30.090 ;
        RECT 214.270 -33.970 218.170 -33.700 ;
        RECT 214.270 -33.980 216.920 -33.970 ;
        RECT 214.270 -33.990 216.210 -33.980 ;
    END
  END IO08
  PIN IO09
    PORT
      LAYER met1 ;
        RECT 215.620 -5.110 218.150 -1.500 ;
        RECT 214.270 -5.390 218.150 -5.110 ;
        RECT 214.270 -5.400 216.210 -5.390 ;
    END
  END IO09
  PIN IO10
    PORT
      LAYER met1 ;
        RECT 216.920 27.100 218.170 27.110 ;
        RECT 216.200 27.090 218.170 27.100 ;
        RECT 215.620 23.480 218.170 27.090 ;
        RECT 214.270 23.220 218.170 23.480 ;
        RECT 214.270 23.210 216.920 23.220 ;
        RECT 214.270 23.190 216.210 23.210 ;
    END
  END IO10
  PIN IO11
    PORT
      LAYER met1 ;
        RECT 215.620 55.670 216.210 55.680 ;
        RECT 215.620 52.070 218.160 55.670 ;
        RECT 214.270 51.780 218.160 52.070 ;
    END
  END IO11
  PIN IO12
    PORT
      LAYER met1 ;
        RECT 215.620 80.660 218.160 84.270 ;
        RECT 214.270 80.380 218.160 80.660 ;
        RECT 214.270 80.370 216.210 80.380 ;
    END
  END IO12
  PIN IO13
    PORT
      LAYER met1 ;
        RECT 216.920 112.860 218.170 112.870 ;
        RECT 215.620 109.250 218.170 112.860 ;
        RECT 214.270 108.980 218.170 109.250 ;
        RECT 214.270 108.970 216.920 108.980 ;
        RECT 214.270 108.960 216.210 108.970 ;
    END
  END IO13
  PIN IO25
    PORT
      LAYER met1 ;
        RECT -153.430 113.570 -152.030 113.580 ;
        RECT -154.680 109.970 -152.030 113.570 ;
        RECT -154.680 109.680 -150.680 109.970 ;
    END
  END IO25
  PIN IO26
    PORT
      LAYER met1 ;
        RECT -154.670 81.380 -152.030 84.990 ;
        RECT -154.670 81.100 -150.680 81.380 ;
        RECT -153.430 81.090 -150.680 81.100 ;
    END
  END IO26
  PIN IO27
    PORT
      LAYER met1 ;
        RECT -153.430 56.390 -152.030 56.400 ;
        RECT -154.680 52.790 -152.030 56.390 ;
        RECT -154.680 52.500 -150.680 52.790 ;
    END
  END IO27
  PIN IO28
    PORT
      LAYER met1 ;
        RECT -153.420 27.800 -152.030 27.810 ;
        RECT -154.660 24.200 -152.030 27.800 ;
        RECT -154.660 23.910 -150.680 24.200 ;
    END
  END IO28
  PIN IO29
    PORT
      LAYER met1 ;
        RECT -154.670 -4.390 -152.030 -0.780 ;
        RECT -154.670 -4.670 -150.680 -4.390 ;
        RECT -153.430 -4.680 -150.680 -4.670 ;
    END
  END IO29
  PIN IO30
    PORT
      LAYER met1 ;
        RECT -153.430 -29.380 -152.030 -29.370 ;
        RECT -154.680 -32.980 -152.030 -29.380 ;
        RECT -154.680 -33.270 -150.680 -32.980 ;
    END
  END IO30
  PIN IO31
    PORT
      LAYER met1 ;
        RECT -153.430 -57.960 -152.620 -57.950 ;
        RECT -154.670 -61.570 -152.030 -57.960 ;
        RECT -154.670 -61.850 -150.680 -61.570 ;
        RECT -152.620 -61.860 -150.680 -61.850 ;
    END
  END IO31
  PIN IO32
    PORT
      LAYER met1 ;
        RECT -154.640 -86.550 -152.600 -86.540 ;
        RECT -154.640 -90.160 -152.030 -86.550 ;
        RECT -154.640 -90.430 -150.680 -90.160 ;
        RECT -153.410 -90.440 -150.680 -90.430 ;
        RECT -152.620 -90.450 -150.680 -90.440 ;
    END
  END IO32
  PIN IO33
    PORT
      LAYER met1 ;
        RECT -153.420 -115.150 -152.030 -115.140 ;
        RECT -154.660 -118.750 -152.030 -115.150 ;
        RECT -154.660 -119.040 -150.680 -118.750 ;
    END
  END IO33
  PIN IO34
    PORT
      LAYER met1 ;
        RECT -153.420 -143.740 -152.030 -143.730 ;
        RECT -154.670 -147.340 -152.030 -143.740 ;
        RECT -154.670 -147.630 -150.680 -147.340 ;
    END
  END IO34
  PIN IO35
    PORT
      LAYER met1 ;
        RECT -153.420 -172.330 -152.030 -172.320 ;
        RECT -154.670 -175.930 -152.030 -172.330 ;
        RECT -154.670 -176.220 -150.680 -175.930 ;
    END
  END IO35
  PIN IO36
    PORT
      LAYER met1 ;
        RECT -153.410 -200.920 -152.030 -200.910 ;
        RECT -154.660 -204.520 -152.030 -200.920 ;
        RECT -154.660 -204.810 -150.680 -204.520 ;
    END
  END IO36
  PIN IO37
    PORT
      LAYER met1 ;
        RECT -154.660 -233.110 -152.030 -229.500 ;
        RECT -154.660 -233.390 -150.680 -233.110 ;
        RECT -153.430 -233.400 -150.680 -233.390 ;
    END
  END IO37
  PIN VSSA1
    ANTENNADIFFAREA 1733.686401 ;
    PORT
      LAYER nwell ;
        RECT 3.820 126.200 6.040 127.890 ;
        RECT 36.080 112.300 39.470 113.050 ;
        RECT 36.070 108.730 39.480 112.300 ;
        RECT 36.070 107.390 39.470 108.730 ;
        RECT 36.080 106.270 39.470 107.390 ;
        RECT 36.080 102.700 39.480 106.270 ;
        RECT 36.090 100.980 39.470 102.700 ;
        RECT 36.050 93.000 39.490 99.490 ;
        RECT 36.080 83.670 37.810 90.170 ;
      LAYER met2 ;
        RECT 213.810 141.650 215.000 141.660 ;
        RECT -151.260 141.640 -53.000 141.650 ;
        RECT 2.430 141.640 215.000 141.650 ;
        RECT -151.390 140.370 215.000 141.640 ;
        RECT -151.390 140.250 202.560 140.370 ;
        RECT -151.390 138.730 -149.100 140.250 ;
        RECT -138.300 140.240 -137.370 140.250 ;
        RECT -109.710 140.240 -108.780 140.250 ;
        RECT -81.120 140.240 -80.190 140.250 ;
        RECT 2.900 140.240 3.830 140.250 ;
        RECT 31.490 140.240 32.420 140.250 ;
        RECT 60.080 140.240 61.010 140.250 ;
        RECT 88.670 140.240 89.600 140.250 ;
        RECT 117.260 140.240 118.190 140.250 ;
        RECT 145.850 140.240 146.780 140.250 ;
        RECT 174.440 140.240 175.370 140.250 ;
        RECT -138.050 139.130 -137.880 140.240 ;
        RECT -109.460 139.130 -109.290 140.240 ;
        RECT -80.870 139.130 -80.700 140.240 ;
        RECT 3.150 139.130 3.320 140.240 ;
        RECT 31.740 139.130 31.910 140.240 ;
        RECT 60.330 139.130 60.500 140.240 ;
        RECT 88.920 139.130 89.090 140.240 ;
        RECT 117.510 139.130 117.680 140.240 ;
        RECT 146.100 139.130 146.270 140.240 ;
        RECT 174.690 139.130 174.860 140.240 ;
        RECT -150.940 138.690 -149.100 138.730 ;
        RECT -150.500 130.560 -149.100 138.690 ;
        RECT -150.530 130.170 -149.100 130.560 ;
        RECT 212.840 139.050 215.000 140.370 ;
        RECT -150.530 103.370 -149.130 130.170 ;
        RECT 212.840 129.840 214.120 139.050 ;
        RECT 13.430 125.480 13.880 125.500 ;
        RECT 13.420 125.470 13.900 125.480 ;
        RECT 37.040 125.470 38.460 125.510 ;
        RECT 13.420 125.070 38.510 125.470 ;
        RECT 13.420 125.060 13.900 125.070 ;
        RECT 13.430 125.040 13.880 125.060 ;
        RECT 37.040 125.030 38.460 125.070 ;
        RECT -22.600 122.860 -22.290 123.070 ;
        RECT -21.170 122.860 -20.860 123.090 ;
        RECT -24.950 122.700 -20.030 122.860 ;
        RECT -26.760 122.530 -20.030 122.700 ;
        RECT 14.520 122.850 15.020 122.870 ;
        RECT 20.260 122.850 20.700 122.900 ;
        RECT 34.630 122.850 35.130 122.870 ;
        RECT -26.760 122.480 -20.020 122.530 ;
        RECT -26.760 122.370 -20.000 122.480 ;
        RECT 14.520 122.430 41.030 122.850 ;
        RECT 14.670 122.410 41.030 122.430 ;
        RECT 20.260 122.400 20.700 122.410 ;
        RECT 40.430 122.390 40.930 122.410 ;
        RECT -26.760 122.300 -24.490 122.370 ;
        RECT -52.870 122.090 -52.390 122.120 ;
        RECT -26.760 122.100 -26.360 122.300 ;
        RECT -23.390 122.160 -23.080 122.370 ;
        RECT -22.460 122.160 -22.150 122.370 ;
        RECT -21.760 122.160 -21.450 122.370 ;
        RECT -21.020 122.190 -20.000 122.370 ;
        RECT -7.910 122.190 -7.600 122.310 ;
        RECT 1.950 122.190 2.260 122.330 ;
        RECT -21.020 122.160 2.260 122.190 ;
        RECT -27.110 122.090 -26.360 122.100 ;
        RECT -52.870 121.710 -26.360 122.090 ;
        RECT -21.000 122.000 2.260 122.160 ;
        RECT -21.000 121.980 2.230 122.000 ;
        RECT -52.870 121.690 -52.390 121.710 ;
        RECT -27.110 121.700 -26.360 121.710 ;
        RECT -52.870 117.320 -52.330 117.350 ;
        RECT -52.870 117.300 -26.930 117.320 ;
        RECT -7.800 117.300 -7.400 117.310 ;
        RECT -52.870 116.950 -7.400 117.300 ;
        RECT -52.870 116.910 -26.930 116.950 ;
        RECT -7.800 116.920 -7.400 116.950 ;
        RECT -52.870 116.870 -52.330 116.910 ;
        RECT 50.900 107.350 51.220 107.500 ;
        RECT 34.710 107.200 51.220 107.350 ;
        RECT 34.710 107.050 35.030 107.200 ;
        RECT 40.510 107.050 40.830 107.200 ;
        RECT 34.780 103.860 35.100 103.910 ;
        RECT 34.780 103.610 40.800 103.860 ;
        RECT 40.480 103.540 40.800 103.610 ;
        RECT -150.530 102.860 -149.120 103.370 ;
        RECT -150.530 102.690 -148.010 102.860 ;
        RECT -150.530 102.440 -149.120 102.690 ;
        RECT 212.720 102.650 214.120 129.840 ;
        RECT -150.530 74.780 -149.130 102.440 ;
        RECT 212.710 102.140 214.120 102.650 ;
        RECT 211.600 101.970 214.120 102.140 ;
        RECT 212.710 101.720 214.120 101.970 ;
        RECT 40.480 101.320 40.800 101.330 ;
        RECT 50.920 101.320 51.250 101.460 ;
        RECT 40.480 101.160 51.250 101.320 ;
        RECT 40.480 101.150 41.170 101.160 ;
        RECT 40.480 101.030 40.800 101.150 ;
        RECT 30.780 94.780 31.100 94.840 ;
        RECT 34.710 94.780 35.030 94.790 ;
        RECT 40.510 94.780 40.830 94.790 ;
        RECT 44.440 94.780 44.760 94.840 ;
        RECT 30.780 94.600 44.760 94.780 ;
        RECT 30.780 94.550 31.100 94.600 ;
        RECT 34.710 94.530 35.030 94.600 ;
        RECT 40.510 94.530 40.830 94.600 ;
        RECT 44.440 94.550 44.760 94.600 ;
        RECT -9.920 89.350 -9.600 89.410 ;
        RECT -8.050 89.380 -7.760 89.400 ;
        RECT -9.920 89.340 -9.440 89.350 ;
        RECT -8.060 89.340 -7.740 89.380 ;
        RECT -9.920 89.150 -7.740 89.340 ;
        RECT -9.920 89.140 -9.440 89.150 ;
        RECT -9.920 89.090 -9.600 89.140 ;
        RECT -8.060 89.120 -7.740 89.150 ;
        RECT -8.050 89.100 -7.760 89.120 ;
        RECT 40.860 85.440 41.190 85.530 ;
        RECT 30.930 85.370 31.250 85.430 ;
        RECT 34.510 85.370 41.190 85.440 ;
        RECT 30.930 85.270 41.190 85.370 ;
        RECT 30.930 85.200 35.280 85.270 ;
        RECT 40.860 85.240 41.190 85.270 ;
        RECT 30.930 85.150 31.250 85.200 ;
        RECT 34.950 85.140 35.280 85.200 ;
        RECT 14.590 82.590 14.920 82.830 ;
        RECT 20.450 82.720 20.750 82.730 ;
        RECT 20.440 82.590 20.760 82.720 ;
        RECT 30.980 82.590 31.260 82.890 ;
        RECT 35.010 82.590 35.310 82.870 ;
        RECT 14.590 82.570 35.310 82.590 ;
        RECT 14.590 82.540 35.300 82.570 ;
        RECT 14.590 82.430 35.240 82.540 ;
        RECT 43.850 82.120 44.150 82.140 ;
        RECT 40.420 81.780 44.160 82.120 ;
        RECT 40.440 81.770 40.750 81.780 ;
        RECT -52.810 81.240 -52.350 81.250 ;
        RECT -52.810 80.820 15.040 81.240 ;
        RECT -52.810 80.800 -26.940 80.820 ;
        RECT -52.810 80.780 -52.350 80.800 ;
        RECT -3.890 80.320 -3.060 80.820 ;
        RECT 43.250 79.330 43.570 81.780 ;
        RECT 43.850 81.760 44.160 81.780 ;
        RECT 40.410 79.000 43.570 79.330 ;
        RECT -10.300 78.800 -10.010 78.820 ;
        RECT -8.070 78.800 -7.760 78.820 ;
        RECT -10.310 78.440 -7.760 78.800 ;
        RECT -10.300 78.420 -10.010 78.440 ;
        RECT -8.070 78.420 -7.760 78.440 ;
        RECT 43.250 77.960 43.570 79.000 ;
        RECT 40.410 77.640 43.570 77.960 ;
        RECT 40.440 77.630 40.750 77.640 ;
        RECT 41.540 77.630 41.850 77.640 ;
        RECT 42.640 77.630 42.950 77.640 ;
        RECT -150.530 74.270 -149.120 74.780 ;
        RECT -150.530 74.100 -148.010 74.270 ;
        RECT -150.530 73.850 -149.120 74.100 ;
        RECT 212.720 74.060 214.120 101.720 ;
        RECT -150.530 46.190 -149.130 73.850 ;
        RECT 212.710 73.550 214.120 74.060 ;
        RECT 211.600 73.380 214.120 73.550 ;
        RECT 212.710 73.130 214.120 73.380 ;
        RECT -150.530 45.680 -149.120 46.190 ;
        RECT -150.530 45.510 -148.010 45.680 ;
        RECT -150.530 45.260 -149.120 45.510 ;
        RECT 212.720 45.470 214.120 73.130 ;
        RECT -150.530 17.600 -149.130 45.260 ;
        RECT 212.710 44.960 214.120 45.470 ;
        RECT 211.600 44.790 214.120 44.960 ;
        RECT 212.710 44.540 214.120 44.790 ;
        RECT -150.530 17.090 -149.120 17.600 ;
        RECT -150.530 16.920 -148.010 17.090 ;
        RECT -150.530 16.670 -149.120 16.920 ;
        RECT 212.720 16.880 214.120 44.540 ;
        RECT -150.530 -10.990 -149.130 16.670 ;
        RECT 212.710 16.370 214.120 16.880 ;
        RECT 211.600 16.200 214.120 16.370 ;
        RECT 212.710 15.950 214.120 16.200 ;
        RECT -150.530 -11.500 -149.120 -10.990 ;
        RECT -150.530 -11.670 -148.010 -11.500 ;
        RECT -150.530 -11.920 -149.120 -11.670 ;
        RECT 212.720 -11.710 214.120 15.950 ;
        RECT -150.530 -39.580 -149.130 -11.920 ;
        RECT 212.710 -12.220 214.120 -11.710 ;
        RECT 211.600 -12.390 214.120 -12.220 ;
        RECT 212.710 -12.640 214.120 -12.390 ;
        RECT -150.530 -40.090 -149.120 -39.580 ;
        RECT -150.530 -40.260 -148.010 -40.090 ;
        RECT -150.530 -40.510 -149.120 -40.260 ;
        RECT 212.720 -40.300 214.120 -12.640 ;
        RECT -150.530 -68.170 -149.130 -40.510 ;
        RECT 212.710 -40.810 214.120 -40.300 ;
        RECT 211.600 -40.980 214.120 -40.810 ;
        RECT 212.710 -41.230 214.120 -40.980 ;
        RECT -150.530 -68.680 -149.120 -68.170 ;
        RECT -150.530 -68.850 -148.010 -68.680 ;
        RECT -150.530 -69.100 -149.120 -68.850 ;
        RECT 212.720 -68.890 214.120 -41.230 ;
        RECT -150.530 -96.760 -149.130 -69.100 ;
        RECT 212.710 -69.400 214.120 -68.890 ;
        RECT 211.600 -69.570 214.120 -69.400 ;
        RECT 212.710 -69.820 214.120 -69.570 ;
        RECT 212.720 -69.980 214.120 -69.820 ;
        RECT 212.720 -70.380 214.130 -69.980 ;
        RECT 212.740 -71.070 214.120 -70.380 ;
        RECT 212.730 -72.240 214.130 -71.070 ;
        RECT -150.530 -97.270 -149.120 -96.760 ;
        RECT -150.530 -97.440 -148.010 -97.270 ;
        RECT -150.530 -97.690 -149.120 -97.440 ;
        RECT -150.530 -125.350 -149.130 -97.690 ;
        RECT -150.530 -125.860 -149.120 -125.350 ;
        RECT -150.530 -126.030 -148.010 -125.860 ;
        RECT -150.530 -126.280 -149.120 -126.030 ;
        RECT -150.530 -153.940 -149.130 -126.280 ;
        RECT -150.530 -154.450 -149.120 -153.940 ;
        RECT -150.530 -154.620 -148.010 -154.450 ;
        RECT -150.530 -154.870 -149.120 -154.620 ;
        RECT -150.530 -182.530 -149.130 -154.870 ;
        RECT -150.530 -183.040 -149.120 -182.530 ;
        RECT -150.530 -183.210 -148.010 -183.040 ;
        RECT -150.530 -183.460 -149.120 -183.210 ;
        RECT -150.530 -211.120 -149.130 -183.460 ;
        RECT -150.530 -211.630 -149.120 -211.120 ;
        RECT -150.530 -211.800 -148.010 -211.630 ;
        RECT -150.530 -212.050 -149.120 -211.800 ;
        RECT -150.530 -239.710 -149.130 -212.050 ;
        RECT -150.530 -240.220 -149.120 -239.710 ;
        RECT -150.530 -240.390 -148.010 -240.220 ;
        RECT -150.530 -240.640 -149.120 -240.390 ;
        RECT -150.530 -243.040 -149.130 -240.640 ;
    END
  END VSSA1
  PIN ANALOG10
    PORT
      LAYER met1 ;
        RECT -131.060 143.740 -127.170 145.710 ;
        RECT -131.060 143.150 -127.160 143.740 ;
        RECT -131.060 141.800 -130.770 143.150 ;
    END
  END ANALOG10
  PIN ANALOG09
    PORT
      LAYER met1 ;
        RECT -102.470 143.740 -98.580 145.700 ;
        RECT -102.470 143.150 -98.570 143.740 ;
        RECT -102.470 141.800 -102.180 143.150 ;
    END
  END ANALOG09
  PIN ANALOG08
    PORT
      LAYER met1 ;
        RECT -73.880 143.740 -69.990 145.700 ;
        RECT -73.880 143.150 -69.980 143.740 ;
        RECT -73.880 141.800 -73.590 143.150 ;
    END
  END ANALOG08
  PIN ANALOG07
    PORT
      LAYER met1 ;
        RECT -31.980 143.760 -28.090 145.730 ;
        RECT -31.980 143.120 -29.570 143.760 ;
        RECT -31.960 141.770 -31.550 143.120 ;
    END
  END ANALOG07
  PIN ANALOG06
    PORT
      LAYER met1 ;
        RECT 10.140 143.740 14.030 145.710 ;
        RECT 10.140 143.150 14.040 143.740 ;
        RECT 10.140 141.800 10.430 143.150 ;
    END
  END ANALOG06
  PIN ANALOG05
    PORT
      LAYER met1 ;
        RECT 38.730 143.740 42.620 145.710 ;
        RECT 38.730 143.150 42.630 143.740 ;
        RECT 38.730 141.800 39.020 143.150 ;
    END
  END ANALOG05
  PIN ANALOG04
    PORT
      LAYER met1 ;
        RECT 67.330 143.740 71.220 145.710 ;
        RECT 67.320 143.150 71.220 143.740 ;
        RECT 67.320 141.800 67.610 143.150 ;
    END
  END ANALOG04
  PIN ANALOG03
    PORT
      LAYER met1 ;
        RECT 95.920 143.740 99.810 145.710 ;
        RECT 95.910 143.150 99.810 143.740 ;
        RECT 95.910 141.800 96.200 143.150 ;
    END
  END ANALOG03
  PIN ANALOG02
    PORT
      LAYER met1 ;
        RECT 124.510 144.540 128.400 145.710 ;
        RECT 124.500 143.740 128.390 144.540 ;
        RECT 124.500 143.150 128.400 143.740 ;
        RECT 124.500 141.800 124.790 143.150 ;
    END
  END ANALOG02
  PIN ANALOG01
    PORT
      LAYER met1 ;
        RECT 153.100 144.540 156.990 145.700 ;
        RECT 153.090 144.530 156.990 144.540 ;
        RECT 153.090 143.740 156.980 144.530 ;
        RECT 153.090 143.150 156.990 143.740 ;
        RECT 153.090 141.800 153.380 143.150 ;
    END
  END ANALOG01
  PIN ANALOG00
    PORT
      LAYER met1 ;
        RECT 181.690 143.740 185.580 145.700 ;
        RECT 181.680 143.150 185.580 143.740 ;
        RECT 181.680 141.800 181.970 143.150 ;
    END
  END ANALOG00
  PIN VDDA1
    ANTENNADIFFAREA 295.115784 ;
    PORT
      LAYER nwell ;
        RECT -123.900 134.780 -111.850 140.720 ;
        RECT -95.310 134.780 -83.260 140.720 ;
        RECT -66.720 134.780 -54.670 140.720 ;
        RECT 17.300 134.780 29.350 140.720 ;
        RECT 45.890 134.780 57.940 140.720 ;
        RECT 74.480 134.780 86.530 140.720 ;
        RECT 103.070 134.780 115.120 140.720 ;
        RECT 131.660 134.780 143.710 140.720 ;
        RECT 160.250 134.780 172.300 140.720 ;
        RECT 188.840 134.780 200.890 140.720 ;
        RECT -149.600 116.840 -143.660 128.890 ;
        RECT -23.810 124.410 -21.070 127.910 ;
        RECT -6.930 121.910 -2.930 127.900 ;
        RECT 17.170 102.830 19.670 116.940 ;
        RECT 207.250 116.120 213.190 128.170 ;
        RECT 26.290 109.970 29.600 113.100 ;
        RECT 22.190 107.070 29.600 109.970 ;
        RECT 45.950 113.050 49.260 113.100 ;
        RECT 45.950 113.040 50.600 113.050 ;
        RECT 22.190 103.380 29.610 107.070 ;
        RECT 26.300 100.920 29.610 103.380 ;
        RECT 45.950 100.970 51.110 113.040 ;
        RECT 45.950 100.920 49.260 100.970 ;
        RECT -149.600 88.250 -143.660 100.300 ;
        RECT 17.170 92.700 19.670 99.700 ;
        RECT 22.170 92.910 25.590 99.500 ;
        RECT 27.710 93.000 30.270 99.500 ;
        RECT 45.270 93.000 47.830 99.500 ;
        RECT 17.130 83.640 19.630 90.640 ;
        RECT 22.200 89.830 25.620 90.230 ;
        RECT 27.740 89.900 30.300 90.170 ;
        RECT 27.340 89.830 30.300 89.900 ;
        RECT 22.200 83.830 30.300 89.830 ;
        RECT 207.250 87.530 213.190 99.580 ;
        RECT 22.200 83.640 25.620 83.830 ;
        RECT 27.740 83.670 30.300 83.830 ;
        RECT -149.600 59.660 -143.660 71.710 ;
        RECT 207.250 58.940 213.190 70.990 ;
        RECT -149.600 31.070 -143.660 43.120 ;
        RECT 207.250 30.350 213.190 42.400 ;
        RECT -149.600 2.480 -143.660 14.530 ;
        RECT 207.250 1.760 213.190 13.810 ;
        RECT -149.600 -26.110 -143.660 -14.060 ;
        RECT 207.250 -26.830 213.190 -14.780 ;
        RECT -149.600 -54.700 -143.660 -42.650 ;
        RECT 207.250 -55.420 213.190 -43.370 ;
        RECT -149.600 -83.290 -143.660 -71.240 ;
        RECT -149.600 -111.880 -143.660 -99.830 ;
        RECT -149.600 -140.470 -143.660 -128.420 ;
        RECT -149.600 -169.060 -143.660 -157.010 ;
        RECT -149.600 -197.650 -143.660 -185.600 ;
        RECT -149.600 -226.240 -143.660 -214.190 ;
      LAYER met2 ;
        RECT -112.430 135.350 -111.790 138.360 ;
        RECT -83.840 135.350 -83.200 138.360 ;
        RECT -55.250 135.350 -54.610 138.360 ;
        RECT 28.770 135.350 29.410 138.360 ;
        RECT 57.360 135.350 58.000 138.360 ;
        RECT 85.950 135.350 86.590 138.360 ;
        RECT 114.540 135.350 115.180 138.360 ;
        RECT 143.130 135.350 143.770 138.360 ;
        RECT 171.720 135.350 172.360 138.360 ;
        RECT 200.310 135.350 200.950 138.360 ;
        RECT -138.770 135.280 207.830 135.350 ;
        RECT -144.230 133.950 207.830 135.280 ;
        RECT -144.230 133.880 -138.480 133.950 ;
        RECT -144.230 130.040 -142.830 133.880 ;
        RECT -113.330 133.820 -110.700 133.950 ;
        RECT -84.740 133.820 -82.110 133.950 ;
        RECT -56.150 133.820 -53.520 133.950 ;
        RECT 27.870 133.820 30.500 133.950 ;
        RECT 56.460 133.820 59.090 133.950 ;
        RECT 85.050 133.820 87.680 133.950 ;
        RECT 113.640 133.820 116.270 133.950 ;
        RECT 142.230 133.820 144.860 133.950 ;
        RECT 170.820 133.820 173.450 133.950 ;
        RECT 199.410 133.820 202.040 133.950 ;
        RECT -113.330 133.310 -110.780 133.820 ;
        RECT -84.740 133.310 -82.190 133.820 ;
        RECT -56.150 133.310 -53.600 133.820 ;
        RECT 27.870 133.310 30.420 133.820 ;
        RECT 56.460 133.310 59.010 133.820 ;
        RECT 85.050 133.310 87.600 133.820 ;
        RECT 113.640 133.310 116.190 133.820 ;
        RECT 142.230 133.310 144.780 133.820 ;
        RECT 170.820 133.310 173.370 133.820 ;
        RECT 199.410 133.310 201.960 133.820 ;
        RECT -113.330 133.240 -112.710 133.310 ;
        RECT -84.740 133.240 -84.120 133.310 ;
        RECT -56.150 133.240 -55.530 133.310 ;
        RECT 27.870 133.240 28.490 133.310 ;
        RECT 56.460 133.240 57.080 133.310 ;
        RECT 85.050 133.240 85.670 133.310 ;
        RECT 113.640 133.240 114.260 133.310 ;
        RECT 142.230 133.240 142.850 133.310 ;
        RECT 170.820 133.240 171.440 133.310 ;
        RECT 199.410 133.240 200.030 133.310 ;
        RECT -144.230 129.960 -142.700 130.040 ;
        RECT -144.230 128.950 -142.190 129.960 ;
        RECT 206.420 129.320 207.820 133.950 ;
        RECT 206.290 129.240 207.820 129.320 ;
        RECT -147.240 128.310 -142.190 128.950 ;
        RECT -144.230 128.030 -142.190 128.310 ;
        RECT 205.780 128.230 207.820 129.240 ;
        RECT -144.230 127.410 -142.120 128.030 ;
        RECT 205.780 127.590 210.830 128.230 ;
        RECT -144.230 101.450 -142.830 127.410 ;
        RECT 205.780 127.310 207.820 127.590 ;
        RECT -56.220 126.510 -55.600 126.530 ;
        RECT -56.220 126.500 -24.620 126.510 ;
        RECT -23.310 126.500 -22.990 126.700 ;
        RECT -22.580 126.500 -22.270 126.710 ;
        RECT -21.900 126.500 -21.580 126.710 ;
        RECT 205.710 126.690 207.820 127.310 ;
        RECT -21.240 126.500 -6.590 126.630 ;
        RECT -56.220 126.420 -6.590 126.500 ;
        RECT -56.220 126.250 -21.100 126.420 ;
        RECT -7.170 126.410 -6.420 126.420 ;
        RECT -56.220 126.140 -21.240 126.250 ;
        RECT -56.220 126.070 -55.600 126.140 ;
        RECT -27.100 126.110 -21.240 126.140 ;
        RECT -24.830 125.740 -21.240 126.110 ;
        RECT -7.170 126.110 -5.550 126.410 ;
        RECT -7.170 125.970 -6.930 126.110 ;
        RECT -5.850 126.050 -5.550 126.110 ;
        RECT -23.310 125.570 -22.990 125.740 ;
        RECT -22.580 125.540 -22.270 125.740 ;
        RECT -21.880 125.590 -21.560 125.740 ;
        RECT -7.190 125.640 -6.880 125.970 ;
        RECT -5.850 125.730 -5.520 126.050 ;
        RECT -5.830 125.720 -5.520 125.730 ;
        RECT 18.940 123.860 19.440 123.890 ;
        RECT 24.660 123.860 25.160 123.890 ;
        RECT 18.940 123.450 49.100 123.860 ;
        RECT 19.090 123.420 49.100 123.450 ;
        RECT -56.340 118.220 -55.720 118.310 ;
        RECT -56.340 118.100 -26.890 118.220 ;
        RECT -56.340 117.810 -24.300 118.100 ;
        RECT -56.340 117.720 -55.720 117.810 ;
        RECT -26.890 117.800 -24.300 117.810 ;
        RECT 26.490 112.910 26.810 113.030 ;
        RECT 48.760 112.910 49.080 113.030 ;
        RECT 26.490 112.730 49.080 112.910 ;
        RECT 47.870 110.190 48.190 110.450 ;
        RECT 47.910 110.170 49.090 110.190 ;
        RECT 47.910 109.910 49.130 110.170 ;
        RECT 47.910 109.850 49.090 109.910 ;
        RECT 47.870 109.840 49.090 109.850 ;
        RECT 47.870 109.590 48.190 109.840 ;
        RECT 26.540 106.850 26.860 106.970 ;
        RECT 48.740 106.850 49.060 106.970 ;
        RECT 26.540 106.670 49.060 106.850 ;
        RECT 47.870 104.160 48.190 104.420 ;
        RECT 47.910 104.140 49.090 104.160 ;
        RECT 47.910 103.880 49.130 104.140 ;
        RECT 47.910 103.820 49.090 103.880 ;
        RECT 47.870 103.810 49.090 103.820 ;
        RECT 47.870 103.560 48.190 103.810 ;
        RECT -144.230 101.370 -142.700 101.450 ;
        RECT -144.230 100.360 -142.190 101.370 ;
        RECT 206.420 100.730 207.820 126.690 ;
        RECT 206.290 100.650 207.820 100.730 ;
        RECT -147.240 99.720 -142.190 100.360 ;
        RECT -144.230 99.440 -142.190 99.720 ;
        RECT 205.780 99.640 207.820 100.650 ;
        RECT -144.230 98.820 -142.120 99.440 ;
        RECT 27.910 99.220 47.650 99.400 ;
        RECT 27.910 99.080 28.330 99.220 ;
        RECT 47.310 99.090 47.650 99.220 ;
        RECT 205.780 99.000 210.830 99.640 ;
        RECT -144.230 72.860 -142.830 98.820 ;
        RECT 205.780 98.720 207.820 99.000 ;
        RECT 205.710 98.100 207.820 98.720 ;
        RECT 19.020 83.290 19.350 83.310 ;
        RECT 19.010 83.210 19.360 83.290 ;
        RECT 24.760 83.210 25.080 83.270 ;
        RECT 19.010 83.050 25.080 83.210 ;
        RECT 19.010 82.980 19.360 83.050 ;
        RECT 24.760 83.000 25.080 83.050 ;
        RECT -56.240 82.220 -55.640 82.270 ;
        RECT -56.240 82.210 -26.900 82.220 ;
        RECT 18.400 82.210 18.840 82.220 ;
        RECT -56.240 82.200 18.840 82.210 ;
        RECT -56.240 81.790 18.860 82.200 ;
        RECT -56.240 81.780 -26.900 81.790 ;
        RECT 11.550 81.780 12.030 81.790 ;
        RECT 18.380 81.780 18.860 81.790 ;
        RECT -56.240 81.710 -55.640 81.780 ;
        RECT 18.400 81.770 18.840 81.780 ;
        RECT -144.230 72.780 -142.700 72.860 ;
        RECT -144.230 71.770 -142.190 72.780 ;
        RECT 206.420 72.140 207.820 98.100 ;
        RECT 206.290 72.060 207.820 72.140 ;
        RECT -147.240 71.130 -142.190 71.770 ;
        RECT -144.230 70.850 -142.190 71.130 ;
        RECT 205.780 71.050 207.820 72.060 ;
        RECT -144.230 70.230 -142.120 70.850 ;
        RECT 205.780 70.410 210.830 71.050 ;
        RECT -144.230 44.270 -142.830 70.230 ;
        RECT 205.780 70.130 207.820 70.410 ;
        RECT 205.710 69.510 207.820 70.130 ;
        RECT -144.230 44.190 -142.700 44.270 ;
        RECT -144.230 43.180 -142.190 44.190 ;
        RECT 206.420 43.550 207.820 69.510 ;
        RECT 206.290 43.470 207.820 43.550 ;
        RECT -147.240 42.540 -142.190 43.180 ;
        RECT -144.230 42.260 -142.190 42.540 ;
        RECT 205.780 42.460 207.820 43.470 ;
        RECT -144.230 41.640 -142.120 42.260 ;
        RECT 205.780 41.820 210.830 42.460 ;
        RECT -144.230 15.680 -142.830 41.640 ;
        RECT 205.780 41.540 207.820 41.820 ;
        RECT 205.710 40.920 207.820 41.540 ;
        RECT -144.230 15.600 -142.700 15.680 ;
        RECT -144.230 14.590 -142.190 15.600 ;
        RECT 206.420 14.960 207.820 40.920 ;
        RECT 206.290 14.880 207.820 14.960 ;
        RECT -147.240 13.950 -142.190 14.590 ;
        RECT -144.230 13.670 -142.190 13.950 ;
        RECT 205.780 13.870 207.820 14.880 ;
        RECT -144.230 13.050 -142.120 13.670 ;
        RECT 205.780 13.230 210.830 13.870 ;
        RECT -144.230 -12.910 -142.830 13.050 ;
        RECT 205.780 12.950 207.820 13.230 ;
        RECT 205.710 12.330 207.820 12.950 ;
        RECT -144.230 -12.990 -142.700 -12.910 ;
        RECT -144.230 -14.000 -142.190 -12.990 ;
        RECT 206.420 -13.630 207.820 12.330 ;
        RECT 206.290 -13.710 207.820 -13.630 ;
        RECT -147.240 -14.640 -142.190 -14.000 ;
        RECT -144.230 -14.920 -142.190 -14.640 ;
        RECT 205.780 -14.720 207.820 -13.710 ;
        RECT -144.230 -15.540 -142.120 -14.920 ;
        RECT 205.780 -15.360 210.830 -14.720 ;
        RECT -144.230 -41.500 -142.830 -15.540 ;
        RECT 205.780 -15.640 207.820 -15.360 ;
        RECT 205.710 -16.260 207.820 -15.640 ;
        RECT -144.230 -41.580 -142.700 -41.500 ;
        RECT -144.230 -42.590 -142.190 -41.580 ;
        RECT 206.420 -42.220 207.820 -16.260 ;
        RECT 206.290 -42.300 207.820 -42.220 ;
        RECT -147.240 -43.230 -142.190 -42.590 ;
        RECT -144.230 -43.510 -142.190 -43.230 ;
        RECT 205.780 -43.310 207.820 -42.300 ;
        RECT -144.230 -44.130 -142.120 -43.510 ;
        RECT 205.780 -43.950 210.830 -43.310 ;
        RECT -144.230 -70.090 -142.830 -44.130 ;
        RECT 205.780 -44.230 207.820 -43.950 ;
        RECT 205.710 -44.850 207.820 -44.230 ;
        RECT -144.230 -70.170 -142.700 -70.090 ;
        RECT -144.230 -71.180 -142.190 -70.170 ;
        RECT 206.420 -70.230 207.820 -44.850 ;
        RECT 206.400 -70.290 207.820 -70.230 ;
        RECT 206.400 -71.010 207.800 -70.290 ;
        RECT 206.390 -71.130 207.800 -71.010 ;
        RECT -147.240 -71.820 -142.190 -71.180 ;
        RECT -144.230 -72.100 -142.190 -71.820 ;
        RECT 206.380 -71.280 207.800 -71.130 ;
        RECT -144.230 -72.720 -142.120 -72.100 ;
        RECT 206.380 -72.180 207.790 -71.280 ;
        RECT -144.230 -98.680 -142.830 -72.720 ;
        RECT -144.230 -98.760 -142.700 -98.680 ;
        RECT -144.230 -99.770 -142.190 -98.760 ;
        RECT -147.240 -100.410 -142.190 -99.770 ;
        RECT -144.230 -100.690 -142.190 -100.410 ;
        RECT -144.230 -101.310 -142.120 -100.690 ;
        RECT -144.230 -127.270 -142.830 -101.310 ;
        RECT -144.230 -127.350 -142.700 -127.270 ;
        RECT -144.230 -128.360 -142.190 -127.350 ;
        RECT -147.240 -129.000 -142.190 -128.360 ;
        RECT -144.230 -129.280 -142.190 -129.000 ;
        RECT -144.230 -129.900 -142.120 -129.280 ;
        RECT -144.230 -155.860 -142.830 -129.900 ;
        RECT -144.230 -155.940 -142.700 -155.860 ;
        RECT -144.230 -156.950 -142.190 -155.940 ;
        RECT -147.240 -157.590 -142.190 -156.950 ;
        RECT -144.230 -157.870 -142.190 -157.590 ;
        RECT -144.230 -158.490 -142.120 -157.870 ;
        RECT -144.230 -184.450 -142.830 -158.490 ;
        RECT -144.230 -184.530 -142.700 -184.450 ;
        RECT -144.230 -185.540 -142.190 -184.530 ;
        RECT -147.240 -186.180 -142.190 -185.540 ;
        RECT -144.230 -186.460 -142.190 -186.180 ;
        RECT -144.230 -187.080 -142.120 -186.460 ;
        RECT -144.230 -213.040 -142.830 -187.080 ;
        RECT -144.230 -213.120 -142.700 -213.040 ;
        RECT -144.230 -214.130 -142.190 -213.120 ;
        RECT -147.240 -214.770 -142.190 -214.130 ;
        RECT -144.230 -215.050 -142.190 -214.770 ;
        RECT -144.230 -215.670 -142.120 -215.050 ;
        RECT -144.230 -243.370 -142.830 -215.670 ;
    END
  END VDDA1
  PIN LADATAOUT01
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 10.930 86.810 11.390 86.960 ;
        RECT 10.540 86.640 11.390 86.810 ;
        RECT 10.540 86.600 10.710 86.640 ;
        RECT 0.940 86.560 1.310 86.570 ;
        RECT 10.540 86.560 10.700 86.600 ;
        RECT 0.940 86.390 10.700 86.560 ;
        RECT 0.940 86.180 1.310 86.390 ;
        RECT 0.850 60.520 1.390 60.590 ;
        RECT -8.580 60.090 1.390 60.520 ;
        RECT -8.580 59.080 -6.600 60.090 ;
        RECT -8.630 58.420 -6.600 59.080 ;
        RECT -8.630 -236.590 -6.610 58.420 ;
        RECT -8.630 -238.150 -6.600 -236.590 ;
        RECT -8.630 -238.160 -6.610 -238.150 ;
    END
  END LADATAOUT01
  PIN LADATAOUT00
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 0.250 85.020 0.640 85.120 ;
        RECT 10.930 85.090 11.390 85.210 ;
        RECT 10.450 85.020 11.390 85.090 ;
        RECT 0.250 84.920 11.390 85.020 ;
        RECT 0.250 84.850 10.740 84.920 ;
        RECT 10.930 84.890 11.390 84.920 ;
        RECT 0.250 84.750 0.640 84.850 ;
        RECT 10.570 84.830 10.740 84.850 ;
        RECT 0.200 61.360 0.740 61.400 ;
        RECT -12.630 61.320 0.740 61.360 ;
        RECT -12.680 60.930 0.740 61.320 ;
        RECT -12.680 59.050 -10.670 60.930 ;
        RECT 0.200 60.900 0.740 60.930 ;
        RECT -12.700 58.390 -10.670 59.050 ;
        RECT -12.690 -238.160 -10.670 58.390 ;
    END
  END LADATAOUT00
  PIN LADATAOUT02
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 10.930 88.620 11.390 88.710 ;
        RECT 10.620 88.450 11.390 88.620 ;
        RECT 1.550 88.100 1.940 88.210 ;
        RECT 10.620 88.160 10.790 88.450 ;
        RECT 10.930 88.390 11.390 88.450 ;
        RECT 10.620 88.100 10.780 88.160 ;
        RECT 1.550 87.940 10.780 88.100 ;
        RECT 1.550 87.930 10.430 87.940 ;
        RECT 1.550 87.830 1.940 87.930 ;
        RECT 1.530 59.710 2.020 59.910 ;
        RECT -4.080 59.690 2.020 59.710 ;
        RECT -4.650 59.410 2.020 59.690 ;
        RECT -4.650 59.310 1.930 59.410 ;
        RECT -4.650 59.080 -2.670 59.310 ;
        RECT -4.670 58.420 -2.640 59.080 ;
        RECT -4.660 -236.600 -2.640 58.420 ;
        RECT -4.670 -238.160 -2.640 -236.600 ;
    END
  END LADATAOUT02
  PIN LADATAOUT03
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 10.930 90.380 11.390 90.460 ;
        RECT 10.680 90.140 11.390 90.380 ;
        RECT 10.680 90.110 11.060 90.140 ;
        RECT 10.680 89.890 10.960 90.110 ;
        RECT 2.210 89.670 2.620 89.770 ;
        RECT 10.680 89.670 10.950 89.890 ;
        RECT 2.210 89.500 10.950 89.670 ;
        RECT 2.210 89.410 2.620 89.500 ;
        RECT 10.680 89.490 10.850 89.500 ;
        RECT 1.360 59.080 2.010 59.090 ;
        RECT -0.670 58.450 2.010 59.080 ;
        RECT -0.670 58.420 1.360 58.450 ;
        RECT -0.660 -236.600 1.360 58.420 ;
        RECT -0.670 -238.160 1.360 -236.600 ;
    END
  END LADATAOUT03
  PIN LADATAOUT04
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 2.850 94.840 3.270 94.930 ;
        RECT 2.850 94.670 10.660 94.840 ;
        RECT 2.850 94.570 3.270 94.670 ;
        RECT 10.490 94.180 10.660 94.670 ;
        RECT 10.970 94.180 11.430 94.270 ;
        RECT 10.490 94.010 11.430 94.180 ;
        RECT 10.970 93.950 11.430 94.010 ;
        RECT 2.860 59.060 3.410 59.080 ;
        RECT 2.860 58.630 5.410 59.060 ;
        RECT 3.380 58.400 5.410 58.630 ;
        RECT 3.390 -238.160 5.410 58.400 ;
    END
  END LADATAOUT04
  PIN LADATAOUT05
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 3.460 96.320 3.850 96.400 ;
        RECT 3.460 96.150 10.640 96.320 ;
        RECT 3.460 96.070 3.850 96.150 ;
        RECT 10.490 96.080 10.640 96.150 ;
        RECT 10.490 95.970 10.660 96.080 ;
        RECT 10.970 95.970 11.430 96.020 ;
        RECT 10.490 95.800 11.430 95.970 ;
        RECT 10.970 95.700 11.430 95.800 ;
        RECT 3.470 59.310 9.450 59.650 ;
        RECT 7.420 59.050 9.460 59.310 ;
        RECT 7.410 58.430 9.460 59.050 ;
        RECT 7.400 58.390 9.460 58.430 ;
        RECT 7.400 -236.590 9.420 58.390 ;
        RECT 7.390 -238.150 9.420 -236.590 ;
        RECT 7.400 -238.160 9.420 -238.150 ;
    END
  END LADATAOUT05
  PIN LADATAOUT06
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 4.080 97.870 4.470 97.960 ;
        RECT 4.080 97.770 11.040 97.870 ;
        RECT 4.080 97.700 11.430 97.770 ;
        RECT 4.080 97.610 4.470 97.700 ;
        RECT 10.750 97.580 11.430 97.700 ;
        RECT 10.970 97.450 11.430 97.580 ;
        RECT 11.370 60.300 13.390 60.320 ;
        RECT 4.210 60.290 13.420 60.300 ;
        RECT 4.110 59.970 13.420 60.290 ;
        RECT 4.110 59.960 4.500 59.970 ;
        RECT 11.340 58.420 13.420 59.970 ;
        RECT 11.400 -238.160 13.420 58.420 ;
    END
  END LADATAOUT06
  PIN LADATAOUT07
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 4.720 99.460 5.090 99.580 ;
        RECT 10.970 99.460 11.430 99.520 ;
        RECT 4.720 99.290 11.430 99.460 ;
        RECT 4.720 99.180 5.090 99.290 ;
        RECT 10.970 99.200 11.430 99.290 ;
        RECT 4.760 60.600 17.500 60.930 ;
        RECT 15.450 59.300 17.480 60.600 ;
        RECT 15.450 59.010 17.490 59.300 ;
        RECT 15.460 58.430 17.490 59.010 ;
        RECT 15.460 58.400 17.510 58.430 ;
        RECT 15.490 -238.160 17.510 58.400 ;
    END
  END LADATAOUT07
  PIN LADATAOUT08
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 5.330 104.930 5.720 105.020 ;
        RECT 5.330 104.760 10.700 104.930 ;
        RECT 5.330 104.670 5.720 104.760 ;
        RECT 10.540 104.650 10.700 104.760 ;
        RECT 10.540 104.350 10.710 104.650 ;
        RECT 10.970 104.350 11.430 104.400 ;
        RECT 10.540 104.180 11.430 104.350 ;
        RECT 10.970 104.080 11.430 104.180 ;
        RECT 5.340 61.570 5.730 61.620 ;
        RECT 5.340 61.290 21.700 61.570 ;
        RECT 5.600 61.240 21.700 61.290 ;
        RECT 19.630 58.430 21.660 61.240 ;
        RECT 19.620 58.420 21.660 58.430 ;
        RECT 19.620 -236.600 21.640 58.420 ;
        RECT 19.610 -238.160 21.640 -236.600 ;
    END
  END LADATAOUT08
  PIN LADATAOUT09
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 5.890 106.500 6.310 106.590 ;
        RECT 5.890 106.330 10.790 106.500 ;
        RECT 5.890 106.240 6.310 106.330 ;
        RECT 10.620 106.150 10.790 106.330 ;
        RECT 10.620 105.980 11.430 106.150 ;
        RECT 10.970 105.830 11.430 105.980 ;
        RECT 5.920 62.180 6.310 62.190 ;
        RECT 5.920 61.860 25.610 62.180 ;
        RECT 6.020 61.850 25.610 61.860 ;
        RECT 23.620 59.140 25.610 61.850 ;
        RECT 23.610 58.390 25.640 59.140 ;
        RECT 23.620 -236.600 25.640 58.390 ;
        RECT 23.610 -238.160 25.640 -236.600 ;
    END
  END LADATAOUT09
  PIN LADATAOUT10
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 6.520 108.030 6.910 108.130 ;
        RECT 6.520 107.900 11.340 108.030 ;
        RECT 6.520 107.860 11.430 107.900 ;
        RECT 6.520 107.760 6.910 107.860 ;
        RECT 10.790 107.700 11.430 107.860 ;
        RECT 10.970 107.580 11.430 107.700 ;
        RECT 6.520 62.830 6.930 62.840 ;
        RECT 6.520 62.810 29.590 62.830 ;
        RECT 6.520 62.500 29.600 62.810 ;
        RECT 6.520 62.490 6.930 62.500 ;
        RECT 27.600 59.120 29.600 62.500 ;
        RECT 27.570 58.420 29.600 59.120 ;
        RECT 27.580 -236.600 29.600 58.420 ;
        RECT 27.570 -238.160 29.600 -236.600 ;
    END
  END LADATAOUT10
  PIN LADATAOUT11
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 7.130 109.600 7.520 109.710 ;
        RECT 10.970 109.600 11.430 109.650 ;
        RECT 7.130 109.430 11.430 109.600 ;
        RECT 7.130 109.330 7.520 109.430 ;
        RECT 10.970 109.330 11.430 109.430 ;
        RECT 7.100 63.450 7.510 63.460 ;
        RECT 7.090 63.120 33.610 63.450 ;
        RECT 7.100 63.100 7.510 63.120 ;
        RECT 31.700 59.050 33.610 63.120 ;
        RECT 31.620 58.400 33.650 59.050 ;
        RECT 31.630 -236.590 33.650 58.400 ;
        RECT 31.630 -238.150 33.660 -236.590 ;
        RECT 31.630 -238.160 33.650 -238.150 ;
    END
  END LADATAOUT11
  PIN LADATAOUT12
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 10.970 110.340 11.430 110.440 ;
        RECT 7.770 110.170 8.160 110.260 ;
        RECT 10.710 110.170 11.430 110.340 ;
        RECT 7.770 110.120 11.430 110.170 ;
        RECT 7.770 110.000 11.340 110.120 ;
        RECT 7.770 109.910 8.160 110.000 ;
        RECT 10.710 109.980 10.880 110.000 ;
        RECT 7.760 64.120 8.160 64.140 ;
        RECT 7.760 63.790 37.700 64.120 ;
        RECT 7.760 63.780 8.160 63.790 ;
        RECT 35.740 59.070 37.690 63.790 ;
        RECT 35.690 58.430 37.720 59.070 ;
        RECT 35.690 58.420 37.740 58.430 ;
        RECT 35.720 -238.160 37.740 58.420 ;
    END
  END LADATAOUT12
  PIN LADATAOUT13
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 10.970 112.060 11.430 112.190 ;
        RECT 10.540 111.890 11.430 112.060 ;
        RECT 8.410 111.770 8.800 111.870 ;
        RECT 10.540 111.770 10.710 111.890 ;
        RECT 10.970 111.870 11.430 111.890 ;
        RECT 8.410 111.600 10.710 111.770 ;
        RECT 8.410 111.500 8.800 111.600 ;
        RECT 8.350 64.760 8.770 64.770 ;
        RECT 8.350 64.430 41.710 64.760 ;
        RECT 8.350 64.420 8.770 64.430 ;
        RECT 39.720 59.070 41.710 64.430 ;
        RECT 39.720 58.420 41.750 59.070 ;
        RECT 39.730 -236.610 41.750 58.420 ;
        RECT 39.730 -238.160 41.760 -236.610 ;
        RECT 39.740 -238.170 41.760 -238.160 ;
    END
  END LADATAOUT13
  PIN LADATAOUT14
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 10.970 113.790 11.430 113.940 ;
        RECT 10.580 113.620 11.430 113.790 ;
        RECT 9.010 113.350 9.340 113.360 ;
        RECT 8.990 113.250 9.360 113.350 ;
        RECT 10.580 113.250 10.750 113.620 ;
        RECT 8.990 113.080 10.750 113.250 ;
        RECT 8.990 112.970 9.360 113.080 ;
        RECT 10.580 113.070 10.750 113.080 ;
        RECT 8.990 65.390 9.370 65.400 ;
        RECT 8.990 65.060 45.790 65.390 ;
        RECT 8.990 65.050 9.370 65.060 ;
        RECT 39.720 65.050 45.790 65.060 ;
        RECT 43.830 64.730 45.790 65.050 ;
        RECT 43.830 59.070 45.780 64.730 ;
        RECT 43.770 58.420 45.800 59.070 ;
        RECT 43.770 -236.600 45.790 58.420 ;
        RECT 43.770 -238.160 45.800 -236.600 ;
    END
  END LADATAOUT14
  PIN LADATAOUT15
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 10.970 115.620 11.430 115.690 ;
        RECT 10.580 115.450 11.430 115.620 ;
        RECT 9.610 114.890 10.000 114.980 ;
        RECT 10.580 114.890 10.750 115.450 ;
        RECT 10.970 115.370 11.430 115.450 ;
        RECT 9.610 114.720 10.760 114.890 ;
        RECT 9.590 66.010 10.010 66.020 ;
        RECT 9.590 65.760 49.860 66.010 ;
        RECT 9.590 65.680 49.870 65.760 ;
        RECT 9.590 65.670 10.010 65.680 ;
        RECT 43.830 65.660 49.870 65.680 ;
        RECT 47.930 65.160 49.870 65.660 ;
        RECT 47.930 59.090 49.860 65.160 ;
        RECT 47.840 58.430 49.870 59.090 ;
        RECT 47.840 58.310 49.880 58.430 ;
        RECT 47.860 -236.620 49.880 58.310 ;
        RECT 47.860 -238.160 49.890 -236.620 ;
        RECT 47.870 -238.180 49.890 -238.160 ;
    END
  END LADATAOUT15
  PIN LADATA16
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT 70.370 109.260 70.830 109.390 ;
        RECT 76.680 109.260 78.150 109.340 ;
        RECT 70.370 109.140 78.150 109.260 ;
        RECT 70.370 109.060 76.950 109.140 ;
        RECT 70.370 108.940 70.830 109.060 ;
        RECT 77.830 109.050 78.150 109.140 ;
        RECT 70.450 65.550 70.880 65.570 ;
        RECT 51.950 65.520 53.910 65.550 ;
        RECT 70.430 65.520 70.890 65.550 ;
        RECT 51.950 65.170 70.890 65.520 ;
        RECT 51.950 59.070 53.910 65.170 ;
        RECT 70.430 65.150 70.890 65.170 ;
        RECT 70.450 65.140 70.880 65.150 ;
        RECT 51.920 58.430 53.950 59.070 ;
        RECT 51.910 58.420 53.950 58.430 ;
        RECT 51.910 -238.160 53.930 58.420 ;
    END
  END LADATA16
  PIN LADATAOUT17
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT 71.380 108.610 71.740 108.710 ;
        RECT 77.830 108.610 78.150 108.700 ;
        RECT 71.380 108.410 78.150 108.610 ;
        RECT 71.380 108.290 71.740 108.410 ;
        RECT 71.350 64.740 71.780 64.760 ;
        RECT 71.340 64.730 71.790 64.740 ;
        RECT 55.880 64.350 71.790 64.730 ;
        RECT 55.880 59.050 57.840 64.350 ;
        RECT 71.350 64.330 71.780 64.350 ;
        RECT 55.870 58.400 57.900 59.050 ;
        RECT 55.880 -238.160 57.900 58.400 ;
    END
  END LADATAOUT17
  PIN LADATAOUT18
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT 72.300 106.350 72.690 106.370 ;
        RECT 72.290 106.240 72.700 106.350 ;
        RECT 72.290 106.140 76.950 106.240 ;
        RECT 72.290 106.040 78.150 106.140 ;
        RECT 72.290 105.940 72.700 106.040 ;
        RECT 76.720 105.940 78.150 106.040 ;
        RECT 72.300 105.920 72.690 105.940 ;
        RECT 77.830 105.850 78.150 105.940 ;
        RECT 72.270 63.910 72.720 63.920 ;
        RECT 60.030 63.530 72.720 63.910 ;
        RECT 60.030 59.070 62.010 63.530 ;
        RECT 59.990 58.420 62.020 59.070 ;
        RECT 60.000 -238.160 62.020 58.420 ;
    END
  END LADATAOUT18
  PIN LADATAOUT19
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT 73.120 105.650 73.520 105.660 ;
        RECT 73.100 105.590 73.540 105.650 ;
        RECT 73.100 105.410 76.950 105.590 ;
        RECT 77.830 105.410 78.150 105.500 ;
        RECT 73.100 105.390 78.150 105.410 ;
        RECT 73.120 105.380 73.520 105.390 ;
        RECT 76.600 105.210 78.150 105.390 ;
        RECT 73.110 63.120 73.530 63.150 ;
        RECT 64.140 62.740 73.530 63.120 ;
        RECT 64.140 59.040 66.120 62.740 ;
        RECT 73.110 62.710 73.530 62.740 ;
        RECT 64.130 58.390 66.160 59.040 ;
        RECT 64.130 -238.170 66.150 58.390 ;
    END
  END LADATAOUT19
  PIN LADATAOUT20
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER met2 ;
        RECT 75.220 68.010 75.480 68.330 ;
        RECT 75.250 59.950 75.450 68.010 ;
        RECT 69.210 59.750 75.450 59.950 ;
        RECT 69.210 59.070 69.410 59.750 ;
        RECT 68.120 58.430 70.150 59.070 ;
        RECT 68.120 58.420 70.160 58.430 ;
        RECT 68.140 -238.160 70.160 58.420 ;
    END
  END LADATAOUT20
  PIN LADATAOUT21
    ANTENNAGATEAREA 0.456300 ;
    PORT
      LAYER met2 ;
        RECT 76.370 71.610 76.570 71.620 ;
        RECT 80.130 71.610 80.450 71.660 ;
        RECT 76.370 71.460 80.450 71.610 ;
        RECT 76.370 59.890 76.570 71.460 ;
        RECT 80.130 71.340 80.450 71.460 ;
        RECT 76.360 59.750 76.570 59.890 ;
        RECT 76.370 59.540 76.570 59.750 ;
        RECT 74.140 59.340 76.570 59.540 ;
        RECT 74.140 59.070 74.340 59.340 ;
        RECT 72.140 58.770 74.340 59.070 ;
        RECT 72.140 58.420 74.170 58.770 ;
        RECT 72.150 -236.480 74.170 58.420 ;
        RECT 72.150 -238.140 74.190 -236.480 ;
    END
  END LADATAOUT21
  PIN LADATAOUT22
    ANTENNAGATEAREA 0.608400 ;
    PORT
      LAYER met2 ;
        RECT 77.340 70.050 80.150 70.060 ;
        RECT 77.340 69.860 80.450 70.050 ;
        RECT 77.340 59.070 77.550 69.860 ;
        RECT 80.130 69.730 80.450 69.860 ;
        RECT 76.220 58.430 78.250 59.070 ;
        RECT 76.220 58.420 78.260 58.430 ;
        RECT 76.240 -236.500 78.260 58.420 ;
        RECT 76.240 -238.160 78.270 -236.500 ;
    END
  END LADATAOUT22
  PIN LADATAOUT23
    ANTENNAGATEAREA 2.281500 ;
    PORT
      LAYER met2 ;
        RECT 79.120 68.400 79.430 68.430 ;
        RECT 80.120 68.400 80.440 68.440 ;
        RECT 79.120 68.150 80.440 68.400 ;
        RECT 79.120 63.450 79.420 68.150 ;
        RECT 80.120 68.120 80.440 68.150 ;
        RECT 79.710 63.450 80.030 63.560 ;
        RECT 79.120 63.240 80.030 63.450 ;
        RECT 79.120 63.230 79.880 63.240 ;
        RECT 79.120 61.810 79.420 63.230 ;
        RECT 79.120 61.650 79.480 61.810 ;
        RECT 78.770 60.210 79.090 60.280 ;
        RECT 79.270 60.210 79.480 61.650 ;
        RECT 78.770 60.010 79.480 60.210 ;
        RECT 78.770 59.960 79.090 60.010 ;
        RECT 79.270 58.980 79.480 60.010 ;
        RECT 80.400 58.980 82.430 59.070 ;
        RECT 79.270 58.770 82.430 58.980 ;
        RECT 80.400 58.420 82.430 58.770 ;
        RECT 80.410 -238.160 82.430 58.420 ;
    END
  END LADATAOUT23
  PIN LADATAOUT24
    ANTENNAGATEAREA 3.650400 ;
    PORT
      LAYER met2 ;
        RECT 80.130 66.500 80.450 66.820 ;
        RECT 80.240 65.210 80.430 66.500 ;
        RECT 80.120 64.890 80.440 65.210 ;
        RECT 80.240 62.010 80.430 64.890 ;
        RECT 80.120 61.690 80.440 62.010 ;
        RECT 80.240 60.300 80.430 61.690 ;
        RECT 80.080 59.980 80.430 60.300 ;
        RECT 80.220 59.770 80.430 59.980 ;
        RECT 80.220 59.750 85.240 59.770 ;
        RECT 80.240 59.580 85.240 59.750 ;
        RECT 85.050 59.120 85.240 59.580 ;
        RECT 85.050 59.050 86.080 59.120 ;
        RECT 84.380 58.430 86.410 59.050 ;
        RECT 84.380 58.400 86.430 58.430 ;
        RECT 84.410 -236.500 86.430 58.400 ;
        RECT 84.410 -238.160 86.440 -236.500 ;
    END
  END LADATAOUT24
  PIN LADATAIN00
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 85.000 39.040 85.110 ;
        RECT 38.730 84.990 41.310 85.000 ;
        RECT 44.520 84.990 44.840 85.040 ;
        RECT 37.800 84.980 44.840 84.990 ;
        RECT 30.180 84.970 44.840 84.980 ;
        RECT 29.900 84.840 44.840 84.970 ;
        RECT 27.740 84.810 39.040 84.840 ;
        RECT 41.230 84.830 44.840 84.840 ;
        RECT 27.740 84.660 30.300 84.810 ;
        RECT 38.730 84.780 39.040 84.810 ;
        RECT 44.520 84.780 44.840 84.830 ;
        RECT 29.900 84.640 30.210 84.660 ;
        RECT 44.500 76.860 90.290 76.870 ;
        RECT 44.500 76.370 90.500 76.860 ;
        RECT 88.490 59.070 90.500 76.370 ;
        RECT 88.430 58.550 90.500 59.070 ;
        RECT 88.430 58.430 90.460 58.550 ;
        RECT 88.420 58.420 90.460 58.430 ;
        RECT 88.420 -236.500 90.440 58.420 ;
        RECT 88.390 -238.160 90.440 -236.500 ;
    END
  END LADATAIN00
  PIN LADATAIN01
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 38.730 85.960 39.040 85.990 ;
        RECT 37.340 85.930 39.040 85.960 ;
        RECT 37.340 85.920 41.310 85.930 ;
        RECT 45.020 85.920 45.340 85.970 ;
        RECT 37.340 85.800 45.340 85.920 ;
        RECT 37.340 85.790 37.800 85.800 ;
        RECT 38.730 85.770 45.340 85.800 ;
        RECT 38.730 85.660 39.040 85.770 ;
        RECT 41.230 85.760 45.340 85.770 ;
        RECT 45.020 85.710 45.340 85.760 ;
        RECT 44.980 77.750 94.250 77.770 ;
        RECT 44.980 77.270 94.360 77.750 ;
        RECT 92.350 59.070 94.360 77.270 ;
        RECT 92.350 58.420 94.420 59.070 ;
        RECT 92.350 58.380 94.400 58.420 ;
        RECT 92.380 -236.500 94.400 58.380 ;
        RECT 92.370 -238.160 94.400 -236.500 ;
    END
  END LADATAIN01
  PIN LADATAIN02
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 29.900 88.090 30.210 88.220 ;
        RECT 27.740 87.910 39.010 88.090 ;
        RECT 29.900 87.890 30.210 87.910 ;
        RECT 38.730 87.880 39.010 87.910 ;
        RECT 38.730 87.770 39.040 87.880 ;
        RECT 38.730 87.760 41.310 87.770 ;
        RECT 45.490 87.760 45.810 87.810 ;
        RECT 38.730 87.610 45.810 87.760 ;
        RECT 38.730 87.550 39.040 87.610 ;
        RECT 41.230 87.600 45.810 87.610 ;
        RECT 45.490 87.550 45.810 87.600 ;
        RECT 96.430 78.670 98.440 78.690 ;
        RECT 45.450 78.170 98.440 78.670 ;
        RECT 96.430 59.050 98.440 78.170 ;
        RECT 96.430 58.400 98.470 59.050 ;
        RECT 96.430 -236.500 98.450 58.400 ;
        RECT 96.430 -238.160 98.470 -236.500 ;
    END
  END LADATAIN02
  PIN LADATAIN03
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 29.900 89.180 30.210 89.200 ;
        RECT 37.700 89.180 37.840 89.190 ;
        RECT 27.740 89.000 37.850 89.180 ;
        RECT 29.900 88.990 37.850 89.000 ;
        RECT 29.900 88.870 30.210 88.990 ;
        RECT 37.700 88.850 37.850 88.990 ;
        RECT 37.700 88.760 38.910 88.850 ;
        RECT 37.700 88.700 39.040 88.760 ;
        RECT 37.700 88.690 41.310 88.700 ;
        RECT 46.010 88.690 46.330 88.740 ;
        RECT 37.700 88.650 46.330 88.690 ;
        RECT 38.730 88.540 46.330 88.650 ;
        RECT 38.730 88.430 39.040 88.540 ;
        RECT 41.230 88.530 46.330 88.540 ;
        RECT 46.010 88.480 46.330 88.530 ;
        RECT 45.990 79.070 102.530 79.570 ;
        RECT 100.520 59.070 102.530 79.070 ;
        RECT 100.490 58.490 102.530 59.070 ;
        RECT 100.490 58.420 102.520 58.490 ;
        RECT 100.490 -236.500 102.510 58.420 ;
        RECT 100.490 -238.160 102.530 -236.500 ;
    END
  END LADATAIN03
  PIN VCCA
    ANTENNADIFFAREA 40.596500 ;
    PORT
      LAYER nwell ;
        RECT -10.540 110.420 -8.510 110.430 ;
        RECT -10.540 107.330 -7.970 110.420 ;
        RECT 11.530 102.830 13.300 116.940 ;
        RECT 53.110 100.970 54.390 113.050 ;
        RECT 77.660 104.070 80.420 110.480 ;
        RECT 11.530 92.700 13.300 99.700 ;
        RECT -12.370 87.500 -10.000 87.700 ;
        RECT -12.370 85.530 -9.440 87.500 ;
        RECT -12.370 84.830 -10.000 85.530 ;
        RECT 11.490 83.640 13.260 90.640 ;
        RECT 29.510 82.390 37.350 82.400 ;
        RECT 27.500 82.370 37.350 82.390 ;
        RECT 19.700 76.700 37.350 82.370 ;
        RECT 19.700 76.670 27.540 76.700 ;
        RECT 74.490 76.050 80.140 76.220 ;
        RECT -15.060 66.980 -11.140 72.680 ;
        RECT 74.490 60.120 81.490 76.050 ;
        RECT 80.130 60.110 81.490 60.120 ;
      LAYER met2 ;
        RECT 11.770 119.640 12.070 119.700 ;
        RECT 53.090 119.640 53.390 119.670 ;
        RECT 11.770 119.410 53.460 119.640 ;
        RECT 11.770 119.380 12.070 119.410 ;
        RECT 53.090 119.330 53.390 119.410 ;
        RECT 53.300 113.870 53.770 113.930 ;
        RECT 78.200 113.880 78.490 113.890 ;
        RECT 78.200 113.870 78.500 113.880 ;
        RECT 88.730 113.870 89.180 113.890 ;
        RECT 53.300 113.440 112.090 113.870 ;
        RECT 78.200 113.430 78.500 113.440 ;
        RECT 78.200 113.410 78.490 113.430 ;
        RECT -9.940 86.740 -9.620 86.790 ;
        RECT -8.480 86.740 -8.160 86.790 ;
        RECT -9.940 86.530 -8.160 86.740 ;
        RECT -9.940 86.470 -9.620 86.530 ;
        RECT -8.480 86.490 -8.160 86.530 ;
        RECT 109.550 84.210 114.080 84.290 ;
        RECT 88.860 84.190 114.150 84.210 ;
        RECT 67.960 83.550 68.520 83.620 ;
        RECT 80.680 83.550 81.360 83.610 ;
        RECT 88.210 83.550 114.150 84.190 ;
        RECT 67.960 83.140 114.150 83.550 ;
        RECT 67.960 83.090 68.520 83.140 ;
        RECT 80.680 83.080 81.360 83.140 ;
        RECT 88.210 83.060 114.150 83.140 ;
        RECT 88.210 83.040 88.870 83.060 ;
        RECT 109.550 83.040 114.080 83.060 ;
        RECT 30.210 81.410 30.520 81.440 ;
        RECT 31.300 81.410 31.610 81.420 ;
        RECT 35.250 81.410 35.560 81.420 ;
        RECT 36.340 81.410 36.650 81.440 ;
        RECT 20.400 81.380 20.710 81.410 ;
        RECT 21.490 81.380 21.800 81.390 ;
        RECT 25.440 81.380 25.750 81.390 ;
        RECT 26.530 81.380 26.840 81.410 ;
        RECT 20.400 81.080 23.350 81.380 ;
        RECT 21.490 81.060 21.800 81.080 ;
        RECT 22.600 81.040 23.350 81.080 ;
        RECT 22.970 80.910 23.350 81.040 ;
        RECT 23.000 80.040 23.350 80.910 ;
        RECT 20.400 79.710 23.350 80.040 ;
        RECT 23.000 77.270 23.350 79.710 ;
        RECT 20.410 77.260 23.350 77.270 ;
        RECT 20.400 76.950 23.350 77.260 ;
        RECT 23.890 81.080 26.840 81.380 ;
        RECT 30.210 81.110 33.160 81.410 ;
        RECT 31.300 81.090 31.610 81.110 ;
        RECT 23.890 81.040 24.640 81.080 ;
        RECT 25.440 81.060 25.750 81.080 ;
        RECT 32.410 81.070 33.160 81.110 ;
        RECT 23.890 80.910 24.270 81.040 ;
        RECT 32.780 80.940 33.160 81.070 ;
        RECT 23.890 80.040 24.240 80.910 ;
        RECT 32.810 80.070 33.160 80.940 ;
        RECT 23.890 79.710 26.840 80.040 ;
        RECT 30.210 79.740 33.160 80.070 ;
        RECT 23.890 77.270 24.240 79.710 ;
        RECT 32.810 77.300 33.160 79.740 ;
        RECT 30.220 77.290 33.160 77.300 ;
        RECT 23.890 77.260 26.830 77.270 ;
        RECT 23.890 76.950 26.840 77.260 ;
        RECT 30.210 76.980 33.160 77.290 ;
        RECT 33.700 81.110 36.650 81.410 ;
        RECT 33.700 81.070 34.450 81.110 ;
        RECT 35.250 81.090 35.560 81.110 ;
        RECT 33.700 80.940 34.080 81.070 ;
        RECT 33.700 80.070 34.050 80.940 ;
        RECT 33.700 79.740 36.650 80.070 ;
        RECT 33.700 77.300 34.050 79.740 ;
        RECT 33.700 77.290 36.640 77.300 ;
        RECT 33.700 76.980 36.650 77.290 ;
        RECT 30.210 76.970 32.930 76.980 ;
        RECT 33.930 76.970 36.650 76.980 ;
        RECT 30.210 76.960 30.520 76.970 ;
        RECT 31.300 76.960 31.610 76.970 ;
        RECT 35.250 76.960 35.560 76.970 ;
        RECT 36.340 76.960 36.650 76.970 ;
        RECT 20.400 76.940 23.120 76.950 ;
        RECT 24.120 76.940 26.840 76.950 ;
        RECT 20.400 76.930 20.710 76.940 ;
        RECT 21.490 76.930 21.800 76.940 ;
        RECT 25.440 76.930 25.750 76.940 ;
        RECT 26.530 76.930 26.840 76.940 ;
        RECT 23.090 76.260 33.990 76.290 ;
        RECT 23.080 76.010 33.990 76.260 ;
        RECT 23.080 75.980 23.420 76.010 ;
        RECT 23.820 76.000 24.160 76.010 ;
        RECT 32.890 75.980 33.230 76.010 ;
        RECT 80.140 73.560 80.430 73.620 ;
        RECT -14.860 73.460 -14.510 73.490 ;
        RECT -8.480 73.480 -8.150 73.520 ;
        RECT -8.490 73.460 -8.140 73.480 ;
        RECT -14.860 73.200 -4.830 73.460 ;
        RECT 79.970 73.250 80.430 73.560 ;
        RECT 80.140 73.210 80.430 73.250 ;
        RECT -14.820 73.170 -4.830 73.200 ;
        RECT -8.480 73.150 -8.150 73.170 ;
        RECT -5.130 71.090 -4.840 73.170 ;
        RECT 80.150 72.890 80.430 73.210 ;
        RECT 79.970 72.580 80.430 72.890 ;
        RECT 80.150 72.460 80.430 72.580 ;
        RECT 11.290 71.090 11.610 71.110 ;
        RECT 67.290 71.090 68.450 71.120 ;
        RECT -5.320 69.970 68.450 71.090 ;
        RECT 11.290 69.950 11.610 69.970 ;
        RECT 22.660 69.890 24.580 69.970 ;
        RECT 32.470 69.860 34.400 69.970 ;
        RECT 67.290 69.940 68.450 69.970 ;
        RECT 108.710 -79.140 113.310 -78.360 ;
        RECT 108.710 -80.820 207.860 -79.140 ;
        RECT 108.710 -82.110 207.990 -80.820 ;
        RECT 108.710 -82.930 113.310 -82.110 ;
    END
  END VCCA
  OBS
      LAYER nwell ;
        RECT -18.200 123.320 -8.510 127.920 ;
        RECT -1.370 127.900 1.340 127.940 ;
        RECT -1.380 126.250 1.340 127.900 ;
        RECT -1.370 124.910 1.340 124.950 ;
        RECT -18.800 121.930 -8.510 123.320 ;
        RECT -1.380 122.250 1.340 124.910 ;
        RECT 31.330 110.660 34.050 112.310 ;
        RECT 41.500 110.660 44.220 112.310 ;
        RECT 31.330 110.620 34.040 110.660 ;
        RECT 41.500 110.620 44.210 110.660 ;
        RECT 31.330 109.290 34.040 109.330 ;
        RECT 41.500 109.290 44.210 109.330 ;
        RECT 31.330 107.640 34.050 109.290 ;
        RECT 41.500 107.640 44.220 109.290 ;
        RECT 31.340 104.630 34.060 106.280 ;
        RECT 31.350 104.590 34.060 104.630 ;
        RECT 41.500 104.630 44.220 106.280 ;
        RECT 41.500 104.590 44.210 104.630 ;
        RECT 31.350 103.260 34.060 103.300 ;
        RECT 31.340 101.610 34.060 103.260 ;
        RECT 41.500 103.260 44.210 103.300 ;
        RECT 41.500 101.610 44.220 103.260 ;
        RECT 31.800 93.000 34.030 99.490 ;
        RECT 41.510 93.000 43.740 99.490 ;
        RECT 31.830 83.670 34.060 90.160 ;
      LAYER li1 ;
        RECT -131.040 141.800 -130.790 143.260 ;
        RECT -131.000 141.790 -130.830 141.800 ;
        RECT -124.360 141.770 -124.110 143.250 ;
        RECT -102.450 141.800 -102.200 143.260 ;
        RECT -102.410 141.790 -102.240 141.800 ;
        RECT -95.770 141.770 -95.520 143.250 ;
        RECT -73.860 141.800 -73.610 143.260 ;
        RECT -73.820 141.790 -73.650 141.800 ;
        RECT -67.180 141.770 -66.930 143.250 ;
        RECT -31.900 141.990 -31.680 143.110 ;
        RECT -31.950 141.800 -31.620 141.990 ;
        RECT -25.160 141.800 -24.920 143.150 ;
        RECT 10.160 141.800 10.410 143.260 ;
        RECT 10.200 141.790 10.370 141.800 ;
        RECT 16.840 141.770 17.090 143.250 ;
        RECT 38.750 141.800 39.000 143.260 ;
        RECT 38.790 141.790 38.960 141.800 ;
        RECT 45.430 141.770 45.680 143.250 ;
        RECT 67.340 141.800 67.590 143.260 ;
        RECT 67.380 141.790 67.550 141.800 ;
        RECT 74.020 141.770 74.270 143.250 ;
        RECT 95.930 141.800 96.180 143.260 ;
        RECT 95.970 141.790 96.140 141.800 ;
        RECT 102.610 141.770 102.860 143.250 ;
        RECT 124.520 141.800 124.770 143.260 ;
        RECT 124.560 141.790 124.730 141.800 ;
        RECT 131.200 141.770 131.450 143.250 ;
        RECT 153.110 141.800 153.360 143.260 ;
        RECT 153.150 141.790 153.320 141.800 ;
        RECT 159.790 141.770 160.040 143.250 ;
        RECT 181.700 141.800 181.950 143.260 ;
        RECT 181.740 141.790 181.910 141.800 ;
        RECT 188.380 141.770 188.630 143.250 ;
        RECT -138.220 141.050 -110.840 141.560 ;
        RECT -138.220 139.120 -137.420 141.050 ;
        RECT -136.840 140.600 -136.670 140.680 ;
        RECT -125.600 140.600 -125.370 140.690 ;
        RECT -136.840 140.590 -125.370 140.600 ;
        RECT -138.220 134.540 -137.710 139.120 ;
        RECT -136.850 135.120 -125.370 140.590 ;
        RECT -136.920 134.950 -125.370 135.120 ;
        RECT -136.850 134.890 -136.660 134.950 ;
        RECT -125.600 134.710 -125.370 134.950 ;
        RECT -136.970 134.540 -135.170 134.550 ;
        RECT -124.810 134.540 -124.300 141.050 ;
        RECT -123.540 140.160 -112.290 140.330 ;
        RECT -123.540 135.290 -123.370 140.160 ;
        RECT -122.980 139.830 -112.870 139.850 ;
        RECT -122.980 139.790 -112.850 139.830 ;
        RECT -123.030 139.620 -112.850 139.790 ;
        RECT -122.980 135.600 -112.850 139.620 ;
        RECT -112.460 138.400 -112.290 140.160 ;
        RECT -122.980 135.520 -112.870 135.600 ;
        RECT -123.550 135.220 -123.370 135.290 ;
        RECT -112.460 135.220 -111.850 138.400 ;
        RECT -123.550 135.050 -111.850 135.220 ;
        RECT -112.390 134.940 -111.850 135.050 ;
        RECT -111.390 134.700 -110.840 141.050 ;
        RECT -111.400 134.540 -110.840 134.700 ;
        RECT -138.220 134.200 -110.840 134.540 ;
        RECT -109.630 141.050 -82.250 141.560 ;
        RECT -109.630 139.120 -108.830 141.050 ;
        RECT -108.250 140.600 -108.080 140.680 ;
        RECT -97.010 140.600 -96.780 140.690 ;
        RECT -108.250 140.590 -96.780 140.600 ;
        RECT -109.630 134.540 -109.120 139.120 ;
        RECT -108.260 135.120 -96.780 140.590 ;
        RECT -108.330 134.950 -96.780 135.120 ;
        RECT -108.260 134.890 -108.070 134.950 ;
        RECT -97.010 134.710 -96.780 134.950 ;
        RECT -108.380 134.540 -106.580 134.550 ;
        RECT -96.220 134.540 -95.710 141.050 ;
        RECT -94.950 140.160 -83.700 140.330 ;
        RECT -94.950 135.290 -94.780 140.160 ;
        RECT -94.390 139.830 -84.280 139.850 ;
        RECT -94.390 139.790 -84.260 139.830 ;
        RECT -94.440 139.620 -84.260 139.790 ;
        RECT -94.390 135.600 -84.260 139.620 ;
        RECT -83.870 138.400 -83.700 140.160 ;
        RECT -94.390 135.520 -84.280 135.600 ;
        RECT -94.960 135.220 -94.780 135.290 ;
        RECT -83.870 135.220 -83.260 138.400 ;
        RECT -94.960 135.050 -83.260 135.220 ;
        RECT -83.800 134.940 -83.260 135.050 ;
        RECT -82.800 134.700 -82.250 141.050 ;
        RECT -82.810 134.540 -82.250 134.700 ;
        RECT -109.630 134.200 -82.250 134.540 ;
        RECT -81.040 141.050 -53.660 141.560 ;
        RECT -81.040 139.120 -80.240 141.050 ;
        RECT -79.660 140.600 -79.490 140.680 ;
        RECT -68.420 140.600 -68.190 140.690 ;
        RECT -79.660 140.590 -68.190 140.600 ;
        RECT -81.040 134.540 -80.530 139.120 ;
        RECT -79.670 135.120 -68.190 140.590 ;
        RECT -79.740 134.950 -68.190 135.120 ;
        RECT -79.670 134.890 -79.480 134.950 ;
        RECT -68.420 134.710 -68.190 134.950 ;
        RECT -79.790 134.540 -77.990 134.550 ;
        RECT -67.630 134.540 -67.120 141.050 ;
        RECT -66.360 140.160 -55.110 140.330 ;
        RECT -66.360 135.290 -66.190 140.160 ;
        RECT -65.800 139.830 -55.690 139.850 ;
        RECT -65.800 139.790 -55.670 139.830 ;
        RECT -65.850 139.620 -55.670 139.790 ;
        RECT -65.800 135.600 -55.670 139.620 ;
        RECT -55.280 138.400 -55.110 140.160 ;
        RECT -65.800 135.520 -55.690 135.600 ;
        RECT -66.370 135.220 -66.190 135.290 ;
        RECT -55.280 135.220 -54.670 138.400 ;
        RECT -66.370 135.050 -54.670 135.220 ;
        RECT -55.210 134.940 -54.670 135.050 ;
        RECT -54.210 134.700 -53.660 141.050 ;
        RECT -54.220 134.540 -53.660 134.700 ;
        RECT -81.040 134.200 -53.660 134.540 ;
        RECT -138.190 134.030 -110.840 134.200 ;
        RECT -109.600 134.030 -82.250 134.200 ;
        RECT -81.010 134.030 -53.660 134.200 ;
        RECT -52.660 141.330 2.080 141.600 ;
        RECT -52.660 141.200 -28.320 141.330 ;
        RECT -19.630 141.200 2.080 141.330 ;
        RECT -138.190 134.010 -137.500 134.030 ;
        RECT -136.990 134.020 -135.190 134.030 ;
        RECT -109.600 134.010 -108.910 134.030 ;
        RECT -108.400 134.020 -106.600 134.030 ;
        RECT -81.010 134.010 -80.320 134.030 ;
        RECT -79.810 134.020 -78.010 134.030 ;
        RECT -52.660 133.600 -52.490 141.200 ;
        RECT 1.910 134.120 2.080 141.200 ;
        RECT 2.980 141.050 30.360 141.560 ;
        RECT 2.980 139.120 3.780 141.050 ;
        RECT 4.360 140.600 4.530 140.680 ;
        RECT 15.600 140.600 15.830 140.690 ;
        RECT 4.360 140.590 15.830 140.600 ;
        RECT 2.980 134.540 3.490 139.120 ;
        RECT 4.350 135.120 15.830 140.590 ;
        RECT 4.280 134.950 15.830 135.120 ;
        RECT 4.350 134.890 4.540 134.950 ;
        RECT 15.600 134.710 15.830 134.950 ;
        RECT 4.230 134.540 6.030 134.550 ;
        RECT 16.390 134.540 16.900 141.050 ;
        RECT 17.660 140.160 28.910 140.330 ;
        RECT 17.660 135.290 17.830 140.160 ;
        RECT 18.220 139.830 28.330 139.850 ;
        RECT 18.220 139.790 28.350 139.830 ;
        RECT 18.170 139.620 28.350 139.790 ;
        RECT 18.220 135.600 28.350 139.620 ;
        RECT 28.740 138.400 28.910 140.160 ;
        RECT 18.220 135.520 28.330 135.600 ;
        RECT 17.650 135.220 17.830 135.290 ;
        RECT 28.740 135.220 29.350 138.400 ;
        RECT 17.650 135.050 29.350 135.220 ;
        RECT 28.810 134.940 29.350 135.050 ;
        RECT 29.810 134.700 30.360 141.050 ;
        RECT 29.800 134.540 30.360 134.700 ;
        RECT 2.980 134.200 30.360 134.540 ;
        RECT 31.570 141.050 58.950 141.560 ;
        RECT 31.570 139.120 32.370 141.050 ;
        RECT 32.950 140.600 33.120 140.680 ;
        RECT 44.190 140.600 44.420 140.690 ;
        RECT 32.950 140.590 44.420 140.600 ;
        RECT 31.570 134.540 32.080 139.120 ;
        RECT 32.940 135.120 44.420 140.590 ;
        RECT 32.870 134.950 44.420 135.120 ;
        RECT 32.940 134.890 33.130 134.950 ;
        RECT 44.190 134.710 44.420 134.950 ;
        RECT 32.820 134.540 34.620 134.550 ;
        RECT 44.980 134.540 45.490 141.050 ;
        RECT 46.250 140.160 57.500 140.330 ;
        RECT 46.250 135.290 46.420 140.160 ;
        RECT 46.810 139.830 56.920 139.850 ;
        RECT 46.810 139.790 56.940 139.830 ;
        RECT 46.760 139.620 56.940 139.790 ;
        RECT 46.810 135.600 56.940 139.620 ;
        RECT 57.330 138.400 57.500 140.160 ;
        RECT 46.810 135.520 56.920 135.600 ;
        RECT 46.240 135.220 46.420 135.290 ;
        RECT 57.330 135.220 57.940 138.400 ;
        RECT 46.240 135.050 57.940 135.220 ;
        RECT 57.400 134.940 57.940 135.050 ;
        RECT 58.400 134.700 58.950 141.050 ;
        RECT 58.390 134.540 58.950 134.700 ;
        RECT 31.570 134.200 58.950 134.540 ;
        RECT 60.160 141.050 87.540 141.560 ;
        RECT 60.160 139.120 60.960 141.050 ;
        RECT 61.540 140.600 61.710 140.680 ;
        RECT 72.780 140.600 73.010 140.690 ;
        RECT 61.540 140.590 73.010 140.600 ;
        RECT 60.160 134.540 60.670 139.120 ;
        RECT 61.530 135.120 73.010 140.590 ;
        RECT 61.460 134.950 73.010 135.120 ;
        RECT 61.530 134.890 61.720 134.950 ;
        RECT 72.780 134.710 73.010 134.950 ;
        RECT 61.410 134.540 63.210 134.550 ;
        RECT 73.570 134.540 74.080 141.050 ;
        RECT 74.840 140.160 86.090 140.330 ;
        RECT 74.840 135.290 75.010 140.160 ;
        RECT 75.400 139.830 85.510 139.850 ;
        RECT 75.400 139.790 85.530 139.830 ;
        RECT 75.350 139.620 85.530 139.790 ;
        RECT 75.400 135.600 85.530 139.620 ;
        RECT 85.920 138.400 86.090 140.160 ;
        RECT 75.400 135.520 85.510 135.600 ;
        RECT 74.830 135.220 75.010 135.290 ;
        RECT 85.920 135.220 86.530 138.400 ;
        RECT 74.830 135.050 86.530 135.220 ;
        RECT 85.990 134.940 86.530 135.050 ;
        RECT 86.990 134.700 87.540 141.050 ;
        RECT 86.980 134.540 87.540 134.700 ;
        RECT 60.160 134.200 87.540 134.540 ;
        RECT 88.750 141.050 116.130 141.560 ;
        RECT 88.750 139.120 89.550 141.050 ;
        RECT 90.130 140.600 90.300 140.680 ;
        RECT 101.370 140.600 101.600 140.690 ;
        RECT 90.130 140.590 101.600 140.600 ;
        RECT 88.750 134.540 89.260 139.120 ;
        RECT 90.120 135.120 101.600 140.590 ;
        RECT 90.050 134.950 101.600 135.120 ;
        RECT 90.120 134.890 90.310 134.950 ;
        RECT 101.370 134.710 101.600 134.950 ;
        RECT 90.000 134.540 91.800 134.550 ;
        RECT 102.160 134.540 102.670 141.050 ;
        RECT 103.430 140.160 114.680 140.330 ;
        RECT 103.430 135.290 103.600 140.160 ;
        RECT 103.990 139.830 114.100 139.850 ;
        RECT 103.990 139.790 114.120 139.830 ;
        RECT 103.940 139.620 114.120 139.790 ;
        RECT 103.990 135.600 114.120 139.620 ;
        RECT 114.510 138.400 114.680 140.160 ;
        RECT 103.990 135.520 114.100 135.600 ;
        RECT 103.420 135.220 103.600 135.290 ;
        RECT 114.510 135.220 115.120 138.400 ;
        RECT 103.420 135.050 115.120 135.220 ;
        RECT 114.580 134.940 115.120 135.050 ;
        RECT 115.580 134.700 116.130 141.050 ;
        RECT 115.570 134.540 116.130 134.700 ;
        RECT 88.750 134.200 116.130 134.540 ;
        RECT 117.340 141.050 144.720 141.560 ;
        RECT 117.340 139.120 118.140 141.050 ;
        RECT 118.720 140.600 118.890 140.680 ;
        RECT 129.960 140.600 130.190 140.690 ;
        RECT 118.720 140.590 130.190 140.600 ;
        RECT 117.340 134.540 117.850 139.120 ;
        RECT 118.710 135.120 130.190 140.590 ;
        RECT 118.640 134.950 130.190 135.120 ;
        RECT 118.710 134.890 118.900 134.950 ;
        RECT 129.960 134.710 130.190 134.950 ;
        RECT 118.590 134.540 120.390 134.550 ;
        RECT 130.750 134.540 131.260 141.050 ;
        RECT 132.020 140.160 143.270 140.330 ;
        RECT 132.020 135.290 132.190 140.160 ;
        RECT 132.580 139.830 142.690 139.850 ;
        RECT 132.580 139.790 142.710 139.830 ;
        RECT 132.530 139.620 142.710 139.790 ;
        RECT 132.580 135.600 142.710 139.620 ;
        RECT 143.100 138.400 143.270 140.160 ;
        RECT 132.580 135.520 142.690 135.600 ;
        RECT 132.010 135.220 132.190 135.290 ;
        RECT 143.100 135.220 143.710 138.400 ;
        RECT 132.010 135.050 143.710 135.220 ;
        RECT 143.170 134.940 143.710 135.050 ;
        RECT 144.170 134.700 144.720 141.050 ;
        RECT 144.160 134.540 144.720 134.700 ;
        RECT 117.340 134.200 144.720 134.540 ;
        RECT 145.930 141.050 173.310 141.560 ;
        RECT 145.930 139.120 146.730 141.050 ;
        RECT 147.310 140.600 147.480 140.680 ;
        RECT 158.550 140.600 158.780 140.690 ;
        RECT 147.310 140.590 158.780 140.600 ;
        RECT 145.930 134.540 146.440 139.120 ;
        RECT 147.300 135.120 158.780 140.590 ;
        RECT 147.230 134.950 158.780 135.120 ;
        RECT 147.300 134.890 147.490 134.950 ;
        RECT 158.550 134.710 158.780 134.950 ;
        RECT 147.180 134.540 148.980 134.550 ;
        RECT 159.340 134.540 159.850 141.050 ;
        RECT 160.610 140.160 171.860 140.330 ;
        RECT 160.610 135.290 160.780 140.160 ;
        RECT 161.170 139.830 171.280 139.850 ;
        RECT 161.170 139.790 171.300 139.830 ;
        RECT 161.120 139.620 171.300 139.790 ;
        RECT 161.170 135.600 171.300 139.620 ;
        RECT 171.690 138.400 171.860 140.160 ;
        RECT 161.170 135.520 171.280 135.600 ;
        RECT 160.600 135.220 160.780 135.290 ;
        RECT 171.690 135.220 172.300 138.400 ;
        RECT 160.600 135.050 172.300 135.220 ;
        RECT 171.760 134.940 172.300 135.050 ;
        RECT 172.760 134.700 173.310 141.050 ;
        RECT 172.750 134.540 173.310 134.700 ;
        RECT 145.930 134.200 173.310 134.540 ;
        RECT 174.520 141.050 201.900 141.560 ;
        RECT 174.520 139.120 175.320 141.050 ;
        RECT 175.900 140.600 176.070 140.680 ;
        RECT 187.140 140.600 187.370 140.690 ;
        RECT 175.900 140.590 187.370 140.600 ;
        RECT 174.520 134.540 175.030 139.120 ;
        RECT 175.890 135.120 187.370 140.590 ;
        RECT 175.820 134.950 187.370 135.120 ;
        RECT 175.890 134.890 176.080 134.950 ;
        RECT 187.140 134.710 187.370 134.950 ;
        RECT 175.770 134.540 177.570 134.550 ;
        RECT 187.930 134.540 188.440 141.050 ;
        RECT 189.200 140.160 200.450 140.330 ;
        RECT 189.200 135.290 189.370 140.160 ;
        RECT 189.760 139.830 199.870 139.850 ;
        RECT 189.760 139.790 199.890 139.830 ;
        RECT 189.710 139.620 199.890 139.790 ;
        RECT 189.760 135.600 199.890 139.620 ;
        RECT 200.280 138.400 200.450 140.160 ;
        RECT 189.760 135.520 199.870 135.600 ;
        RECT 189.190 135.220 189.370 135.290 ;
        RECT 200.280 135.220 200.890 138.400 ;
        RECT 189.190 135.050 200.890 135.220 ;
        RECT 200.350 134.940 200.890 135.050 ;
        RECT 201.350 134.700 201.900 141.050 ;
        RECT 201.340 134.540 201.900 134.700 ;
        RECT 174.520 134.200 201.900 134.540 ;
        RECT 3.010 134.030 30.360 134.200 ;
        RECT 31.600 134.030 58.950 134.200 ;
        RECT 60.190 134.030 87.540 134.200 ;
        RECT 88.780 134.030 116.130 134.200 ;
        RECT 117.370 134.030 144.720 134.200 ;
        RECT 145.960 134.030 173.310 134.200 ;
        RECT 174.550 134.030 201.900 134.200 ;
        RECT 3.010 134.010 3.700 134.030 ;
        RECT 4.210 134.020 6.010 134.030 ;
        RECT 31.600 134.010 32.290 134.030 ;
        RECT 32.800 134.020 34.600 134.030 ;
        RECT 60.190 134.010 60.880 134.030 ;
        RECT 61.390 134.020 63.190 134.030 ;
        RECT 88.780 134.010 89.470 134.030 ;
        RECT 89.980 134.020 91.780 134.030 ;
        RECT 117.370 134.010 118.060 134.030 ;
        RECT 118.570 134.020 120.370 134.030 ;
        RECT 145.960 134.010 146.650 134.030 ;
        RECT 147.160 134.020 148.960 134.030 ;
        RECT 174.550 134.010 175.240 134.030 ;
        RECT 175.750 134.020 177.550 134.030 ;
        RECT -26.220 133.260 -23.860 133.430 ;
        RECT -150.440 129.350 -142.910 129.900 ;
        RECT -152.130 116.380 -150.650 116.630 ;
        RECT -150.440 116.440 -149.930 129.350 ;
        RECT -143.580 129.340 -142.910 129.350 ;
        RECT -147.280 128.450 -143.820 128.890 ;
        RECT -149.210 128.350 -143.820 128.450 ;
        RECT -149.210 128.280 -143.930 128.350 ;
        RECT -149.210 117.370 -149.040 128.280 ;
        RECT -148.710 127.870 -144.480 127.890 ;
        RECT -148.730 117.760 -144.400 127.870 ;
        RECT -148.670 117.710 -148.500 117.760 ;
        RECT -144.100 117.370 -143.930 128.280 ;
        RECT -149.210 117.200 -143.930 117.370 ;
        RECT -144.170 117.190 -143.930 117.200 ;
        RECT -143.420 116.440 -142.910 129.340 ;
        RECT 206.500 128.630 214.030 129.180 ;
        RECT 206.500 128.620 207.170 128.630 ;
        RECT -23.850 127.630 -23.680 127.790 ;
        RECT -22.450 127.630 -22.280 127.790 ;
        RECT -23.850 127.490 -23.610 127.630 ;
        RECT -23.850 127.460 -22.810 127.490 ;
        RECT -22.450 127.480 -22.240 127.630 ;
        RECT -20.610 127.520 -19.940 127.690 ;
        RECT -22.450 127.460 -21.400 127.480 ;
        RECT -23.810 127.310 -22.810 127.460 ;
        RECT -22.410 127.310 -21.400 127.460 ;
        RECT -20.610 126.730 -19.940 126.900 ;
        RECT -22.600 126.630 -22.280 126.670 ;
        RECT -23.480 126.460 -21.400 126.630 ;
        RECT -6.590 126.590 -3.280 127.570 ;
        RECT 0.810 126.770 1.040 127.460 ;
        RECT 5.510 126.720 5.740 127.410 ;
        RECT -22.610 126.440 -22.280 126.460 ;
        RECT -22.600 126.410 -22.280 126.440 ;
        RECT -23.300 126.050 -21.480 126.220 ;
        RECT -22.600 125.810 -22.280 125.830 ;
        RECT -23.480 125.640 -21.400 125.810 ;
        RECT -20.690 125.800 -20.480 126.230 ;
        RECT -6.480 125.930 -6.310 126.280 ;
        RECT -5.760 126.010 -5.590 126.040 ;
        RECT -5.850 125.970 -5.530 126.010 ;
        RECT -5.080 126.000 -4.910 126.040 ;
        RECT -7.210 125.890 -6.310 125.930 ;
        RECT -20.670 125.780 -20.500 125.800 ;
        RECT -7.220 125.700 -6.310 125.890 ;
        RECT -5.860 125.780 -5.530 125.970 ;
        RECT -5.160 125.960 -4.840 126.000 ;
        RECT -5.850 125.750 -5.530 125.780 ;
        RECT -5.170 125.770 -4.840 125.960 ;
        RECT -5.760 125.710 -5.590 125.750 ;
        RECT -5.160 125.740 -4.840 125.770 ;
        RECT -5.080 125.710 -4.910 125.740 ;
        RECT -7.210 125.670 -6.310 125.700 ;
        RECT 2.020 125.690 2.190 125.710 ;
        RECT -22.610 125.600 -22.280 125.640 ;
        RECT -22.600 125.570 -22.280 125.600 ;
        RECT -20.610 125.300 -19.940 125.470 ;
        RECT -23.480 124.800 -22.810 124.970 ;
        RECT -22.080 124.800 -21.400 124.970 ;
        RECT -21.100 124.680 -20.910 124.740 ;
        RECT -21.100 124.510 -19.930 124.680 ;
        RECT -21.170 124.230 -21.000 124.260 ;
        RECT -21.170 124.200 -20.840 124.230 ;
        RECT -21.170 124.010 -20.830 124.200 ;
        RECT -21.170 123.970 -20.840 124.010 ;
        RECT -21.170 123.930 -21.000 123.970 ;
        RECT -22.420 123.850 -22.250 123.910 ;
        RECT -20.600 123.900 -19.930 124.070 ;
        RECT -23.480 123.680 -22.810 123.850 ;
        RECT -22.420 123.680 -21.400 123.850 ;
        RECT -22.420 123.580 -22.250 123.680 ;
        RECT -22.620 123.010 -22.300 123.030 ;
        RECT -21.190 123.010 -20.870 123.050 ;
        RECT -23.490 122.840 -19.910 123.010 ;
        RECT -22.630 122.800 -22.300 122.840 ;
        RECT -21.200 122.820 -20.870 122.840 ;
        RECT -22.620 122.770 -22.300 122.800 ;
        RECT -21.190 122.790 -20.870 122.820 ;
        RECT -23.410 122.410 -23.090 122.450 ;
        RECT -22.480 122.410 -22.160 122.450 ;
        RECT -21.780 122.410 -21.460 122.450 ;
        RECT -21.040 122.410 -20.720 122.450 ;
        RECT -23.420 122.340 -23.090 122.410 ;
        RECT -22.490 122.340 -22.160 122.410 ;
        RECT -21.790 122.340 -21.460 122.410 ;
        RECT -21.050 122.390 -20.720 122.410 ;
        RECT -20.330 122.400 -20.010 122.440 ;
        RECT -20.340 122.390 -20.010 122.400 ;
        RECT -21.050 122.340 -20.010 122.390 ;
        RECT -23.440 122.170 -20.010 122.340 ;
        RECT -18.340 122.230 -18.170 122.900 ;
        RECT -7.850 122.810 -7.680 125.460 ;
        RECT -6.480 125.270 -6.310 125.670 ;
        RECT -0.870 125.520 2.190 125.690 ;
        RECT 2.020 124.870 2.190 125.520 ;
        RECT -6.590 123.790 -3.280 124.770 ;
        RECT 2.020 124.700 3.290 124.870 ;
        RECT 0.810 123.780 1.040 124.470 ;
        RECT -7.850 122.270 -7.670 122.810 ;
        RECT -7.930 122.230 -7.610 122.270 ;
        RECT -6.590 122.240 -3.280 123.220 ;
        RECT 0.810 122.770 1.040 123.460 ;
        RECT 2.020 122.290 2.190 124.700 ;
        RECT 4.760 123.050 4.930 123.940 ;
        RECT 1.930 122.250 2.250 122.290 ;
        RECT -20.860 122.160 -20.010 122.170 ;
        RECT -7.940 122.040 -7.610 122.230 ;
        RECT 1.920 122.060 2.250 122.250 ;
        RECT -7.930 122.010 -7.610 122.040 ;
        RECT 1.930 122.030 2.250 122.060 ;
        RECT -7.900 118.450 -6.380 118.460 ;
        RECT -7.900 117.660 -6.350 118.450 ;
        RECT -150.440 115.930 -142.910 116.440 ;
        RECT 13.190 116.400 13.540 116.500 ;
        RECT 16.950 116.490 17.240 116.510 ;
        RECT 16.780 116.450 17.240 116.490 ;
        RECT 15.800 116.430 17.240 116.450 ;
        RECT 14.850 116.400 15.310 116.430 ;
        RECT 11.780 116.230 12.540 116.400 ;
        RECT 12.790 116.230 13.960 116.400 ;
        RECT 14.200 116.260 15.310 116.400 ;
        RECT 15.760 116.270 17.240 116.430 ;
        RECT 15.760 116.260 16.950 116.270 ;
        RECT 14.200 116.230 15.020 116.260 ;
        RECT 11.780 116.220 12.010 116.230 ;
        RECT -152.140 109.910 -150.680 109.950 ;
        RECT -152.140 109.740 -150.670 109.910 ;
        RECT -152.140 109.700 -150.680 109.740 ;
        RECT -150.440 103.320 -149.930 115.930 ;
        RECT -149.570 115.140 -143.590 115.370 ;
        RECT -149.480 104.080 -143.830 115.140 ;
        RECT -143.420 105.570 -142.910 115.930 ;
        RECT 11.740 115.780 12.010 116.220 ;
        RECT 14.760 116.090 15.020 116.230 ;
        RECT 13.220 115.780 13.550 116.040 ;
        RECT 14.760 115.920 15.940 116.090 ;
        RECT 14.760 115.780 15.020 115.920 ;
        RECT 11.190 115.640 11.360 115.700 ;
        RECT 11.160 115.420 11.380 115.640 ;
        RECT 11.710 115.600 12.040 115.780 ;
        RECT 12.290 115.610 14.450 115.780 ;
        RECT 14.690 115.610 15.020 115.780 ;
        RECT 14.850 115.560 15.020 115.610 ;
        RECT 15.310 115.420 15.520 115.750 ;
        RECT 15.760 115.480 15.940 115.920 ;
        RECT 17.570 115.820 17.740 116.580 ;
        RECT 17.940 116.430 18.390 116.580 ;
        RECT 17.940 116.260 18.540 116.430 ;
        RECT 19.000 116.250 19.330 116.420 ;
        RECT 17.360 115.810 17.740 115.820 ;
        RECT 17.360 115.750 17.830 115.810 ;
        RECT 19.080 115.790 19.260 116.250 ;
        RECT 16.490 115.640 17.830 115.750 ;
        RECT 16.490 115.580 17.750 115.640 ;
        RECT 18.300 115.620 19.260 115.790 ;
        RECT 206.500 115.720 207.010 128.620 ;
        RECT 207.410 127.730 210.870 128.170 ;
        RECT 207.410 127.630 212.800 127.730 ;
        RECT 207.520 127.560 212.800 127.630 ;
        RECT 207.520 116.650 207.690 127.560 ;
        RECT 208.070 127.150 212.300 127.170 ;
        RECT 207.990 117.040 212.320 127.150 ;
        RECT 212.090 116.990 212.260 117.040 ;
        RECT 212.630 116.650 212.800 127.560 ;
        RECT 207.520 116.480 212.800 116.650 ;
        RECT 207.520 116.470 207.760 116.480 ;
        RECT 213.520 115.720 214.030 128.630 ;
        RECT 17.360 115.530 17.750 115.580 ;
        RECT 11.190 115.370 11.360 115.420 ;
        RECT 13.190 114.650 13.540 114.750 ;
        RECT 16.950 114.740 17.240 114.760 ;
        RECT 16.780 114.700 17.240 114.740 ;
        RECT 15.800 114.680 17.240 114.700 ;
        RECT 14.850 114.650 15.310 114.680 ;
        RECT 11.780 114.480 12.540 114.650 ;
        RECT 12.790 114.480 13.960 114.650 ;
        RECT 14.200 114.510 15.310 114.650 ;
        RECT 15.760 114.520 17.240 114.680 ;
        RECT 15.760 114.510 16.950 114.520 ;
        RECT 14.200 114.480 15.020 114.510 ;
        RECT 11.780 114.470 12.010 114.480 ;
        RECT 11.740 114.030 12.010 114.470 ;
        RECT 14.760 114.340 15.020 114.480 ;
        RECT 13.220 114.030 13.550 114.290 ;
        RECT 14.760 114.170 15.940 114.340 ;
        RECT 14.760 114.030 15.020 114.170 ;
        RECT 11.190 113.890 11.360 113.950 ;
        RECT 11.160 113.670 11.380 113.890 ;
        RECT 11.710 113.850 12.040 114.030 ;
        RECT 12.290 113.860 14.450 114.030 ;
        RECT 14.690 113.860 15.020 114.030 ;
        RECT 14.850 113.810 15.020 113.860 ;
        RECT 15.310 113.670 15.520 114.000 ;
        RECT 15.760 113.730 15.940 114.170 ;
        RECT 17.570 114.070 17.740 114.830 ;
        RECT 17.940 114.680 18.390 114.830 ;
        RECT 17.940 114.510 18.540 114.680 ;
        RECT 19.000 114.500 19.330 114.670 ;
        RECT 40.070 114.500 40.740 115.370 ;
        RECT 52.350 114.520 54.450 115.370 ;
        RECT 206.500 115.210 214.030 115.720 ;
        RECT 214.240 115.660 215.720 115.910 ;
        RECT 17.360 114.060 17.740 114.070 ;
        RECT 17.360 114.000 17.830 114.060 ;
        RECT 19.080 114.040 19.260 114.500 ;
        RECT 16.490 113.890 17.830 114.000 ;
        RECT 16.490 113.830 17.750 113.890 ;
        RECT 18.300 113.870 19.260 114.040 ;
        RECT 17.360 113.780 17.750 113.830 ;
        RECT 11.190 113.620 11.360 113.670 ;
        RECT -9.700 113.130 -9.500 113.170 ;
        RECT -10.010 112.870 -9.500 113.130 ;
        RECT -9.700 112.840 -9.500 112.870 ;
        RECT -9.110 113.140 -8.910 113.170 ;
        RECT -9.110 113.100 -8.600 113.140 ;
        RECT -9.110 112.910 -8.590 113.100 ;
        RECT -9.110 112.880 -8.600 112.910 ;
        RECT 13.190 112.900 13.540 113.000 ;
        RECT 16.950 112.990 17.240 113.010 ;
        RECT 16.780 112.950 17.240 112.990 ;
        RECT 15.800 112.930 17.240 112.950 ;
        RECT 14.850 112.900 15.310 112.930 ;
        RECT -9.110 112.840 -8.910 112.880 ;
        RECT 11.780 112.730 12.540 112.900 ;
        RECT 12.790 112.730 13.960 112.900 ;
        RECT 14.200 112.760 15.310 112.900 ;
        RECT 15.760 112.770 17.240 112.930 ;
        RECT 15.760 112.760 16.950 112.770 ;
        RECT 14.200 112.730 15.020 112.760 ;
        RECT 11.780 112.720 12.010 112.730 ;
        RECT -10.280 112.630 -9.920 112.700 ;
        RECT -10.440 112.530 -9.920 112.630 ;
        RECT -8.410 112.590 -8.240 112.640 ;
        RECT -8.420 112.560 -8.240 112.590 ;
        RECT -8.420 112.550 -7.990 112.560 ;
        RECT -10.440 112.450 -10.070 112.530 ;
        RECT -10.440 112.400 -10.110 112.450 ;
        RECT -10.440 112.370 -10.120 112.400 ;
        RECT -8.420 112.320 -7.830 112.550 ;
        RECT -8.420 112.310 -7.990 112.320 ;
        RECT -8.420 112.280 -8.230 112.310 ;
        RECT 11.740 112.280 12.010 112.720 ;
        RECT 14.760 112.590 15.020 112.730 ;
        RECT 13.220 112.280 13.550 112.540 ;
        RECT 14.760 112.420 15.940 112.590 ;
        RECT 14.760 112.280 15.020 112.420 ;
        RECT -8.410 112.250 -8.230 112.280 ;
        RECT -9.690 112.140 -9.490 112.180 ;
        RECT -10.000 111.880 -9.490 112.140 ;
        RECT -9.690 111.850 -9.490 111.880 ;
        RECT -9.100 112.150 -8.900 112.180 ;
        RECT -9.100 112.110 -8.590 112.150 ;
        RECT 11.190 112.140 11.360 112.200 ;
        RECT -9.100 111.920 -8.580 112.110 ;
        RECT 11.160 111.920 11.380 112.140 ;
        RECT 11.710 112.100 12.040 112.280 ;
        RECT 12.290 112.110 14.450 112.280 ;
        RECT 14.690 112.110 15.020 112.280 ;
        RECT 14.850 112.060 15.020 112.110 ;
        RECT 15.310 111.920 15.520 112.250 ;
        RECT 15.760 111.980 15.940 112.420 ;
        RECT 17.570 112.320 17.740 113.080 ;
        RECT 17.940 112.930 18.390 113.080 ;
        RECT 50.240 113.000 50.410 113.050 ;
        RECT 17.940 112.760 18.540 112.930 ;
        RECT 19.000 112.750 19.330 112.920 ;
        RECT 17.360 112.310 17.740 112.320 ;
        RECT 17.360 112.250 17.830 112.310 ;
        RECT 19.080 112.290 19.260 112.750 ;
        RECT 50.240 112.740 50.800 113.000 ;
        RECT 51.710 112.750 51.910 112.790 ;
        RECT 50.240 112.720 50.410 112.740 ;
        RECT 26.690 112.370 26.890 112.720 ;
        RECT 28.170 112.470 28.700 112.640 ;
        RECT 28.940 112.620 29.130 112.650 ;
        RECT 28.940 112.450 30.000 112.620 ;
        RECT 46.850 112.470 47.380 112.640 ;
        RECT 28.940 112.420 29.130 112.450 ;
        RECT 16.490 112.140 17.830 112.250 ;
        RECT 16.490 112.080 17.750 112.140 ;
        RECT 18.300 112.120 19.260 112.290 ;
        RECT 26.680 112.340 26.890 112.370 ;
        RECT 17.360 112.030 17.750 112.080 ;
        RECT -9.100 111.890 -8.590 111.920 ;
        RECT -9.100 111.850 -8.900 111.890 ;
        RECT 11.190 111.870 11.360 111.920 ;
        RECT 26.680 111.760 26.900 112.340 ;
        RECT 26.680 111.750 26.890 111.760 ;
        RECT -10.460 111.540 -9.910 111.710 ;
        RECT 27.060 111.580 27.250 111.590 ;
        RECT -10.460 111.480 -10.130 111.540 ;
        RECT -10.460 111.450 -10.140 111.480 ;
        RECT -9.690 111.150 -9.490 111.190 ;
        RECT -10.000 110.890 -9.490 111.150 ;
        RECT -9.690 110.860 -9.490 110.890 ;
        RECT -9.100 111.160 -8.900 111.190 ;
        RECT -9.100 111.120 -8.590 111.160 ;
        RECT 13.190 111.150 13.540 111.250 ;
        RECT 16.950 111.240 17.240 111.260 ;
        RECT 16.780 111.200 17.240 111.240 ;
        RECT 15.800 111.180 17.240 111.200 ;
        RECT 14.850 111.150 15.310 111.180 ;
        RECT -9.100 110.930 -8.580 111.120 ;
        RECT 11.780 110.980 12.540 111.150 ;
        RECT 12.790 110.980 13.960 111.150 ;
        RECT 14.200 111.010 15.310 111.150 ;
        RECT 15.760 111.020 17.240 111.180 ;
        RECT 15.760 111.010 16.950 111.020 ;
        RECT 14.200 110.980 15.020 111.010 ;
        RECT 11.780 110.970 12.010 110.980 ;
        RECT -9.100 110.900 -8.590 110.930 ;
        RECT -9.100 110.860 -8.900 110.900 ;
        RECT -10.480 110.550 -9.910 110.720 ;
        RECT -10.480 110.490 -10.150 110.550 ;
        RECT 11.740 110.530 12.010 110.970 ;
        RECT 14.760 110.840 15.020 110.980 ;
        RECT 13.220 110.530 13.550 110.790 ;
        RECT 14.760 110.670 15.940 110.840 ;
        RECT 14.760 110.530 15.020 110.670 ;
        RECT -10.480 110.460 -10.160 110.490 ;
        RECT 11.190 110.390 11.360 110.450 ;
        RECT -10.190 110.180 -9.870 110.220 ;
        RECT -10.190 110.160 -9.860 110.180 ;
        RECT 11.160 110.170 11.380 110.390 ;
        RECT 11.710 110.350 12.040 110.530 ;
        RECT 12.290 110.360 14.450 110.530 ;
        RECT 14.690 110.360 15.020 110.530 ;
        RECT 14.850 110.310 15.020 110.360 ;
        RECT 15.310 110.170 15.520 110.500 ;
        RECT 15.760 110.230 15.940 110.670 ;
        RECT 17.570 110.570 17.740 111.330 ;
        RECT 17.940 111.180 18.390 111.330 ;
        RECT 27.050 111.290 27.250 111.580 ;
        RECT 17.940 111.010 18.540 111.180 ;
        RECT 19.000 111.000 19.330 111.170 ;
        RECT 17.360 110.560 17.740 110.570 ;
        RECT 17.360 110.500 17.830 110.560 ;
        RECT 19.080 110.540 19.260 111.000 ;
        RECT 26.990 110.960 27.260 111.290 ;
        RECT 16.490 110.390 17.830 110.500 ;
        RECT 16.490 110.330 17.750 110.390 ;
        RECT 18.300 110.370 19.260 110.540 ;
        RECT 27.450 110.480 27.620 112.090 ;
        RECT 28.280 110.990 28.450 112.080 ;
        RECT 29.410 112.060 29.600 112.090 ;
        RECT 28.870 111.890 29.600 112.060 ;
        RECT 29.830 112.060 30.000 112.450 ;
        RECT 48.660 112.370 48.860 112.720 ;
        RECT 48.660 112.340 48.870 112.370 ;
        RECT 29.830 111.890 30.570 112.060 ;
        RECT 29.410 111.860 29.600 111.890 ;
        RECT 31.630 111.270 31.860 111.790 ;
        RECT 28.870 111.100 31.860 111.270 ;
        RECT 28.050 110.950 28.450 110.990 ;
        RECT 28.040 110.760 28.450 110.950 ;
        RECT 36.830 110.910 37.380 111.340 ;
        RECT 38.170 110.910 38.720 111.340 ;
        RECT 41.800 111.100 42.030 111.790 ;
        RECT 47.100 111.560 47.270 112.080 ;
        RECT 46.940 111.300 47.270 111.560 ;
        RECT 28.050 110.730 28.450 110.760 ;
        RECT 17.360 110.280 17.750 110.330 ;
        RECT 27.440 110.290 27.620 110.480 ;
        RECT 28.280 110.390 28.450 110.730 ;
        RECT 28.940 110.480 29.130 110.660 ;
        RECT 28.870 110.310 29.220 110.480 ;
        RECT -10.190 109.960 -9.570 110.160 ;
        RECT -9.740 109.830 -9.570 109.960 ;
        RECT -9.060 110.120 -8.890 110.160 ;
        RECT 11.190 110.120 11.360 110.170 ;
        RECT -9.060 110.080 -8.570 110.120 ;
        RECT -9.060 109.890 -8.560 110.080 ;
        RECT 29.790 109.900 30.000 110.330 ;
        RECT 30.220 110.310 30.560 110.480 ;
        RECT -9.060 109.860 -8.570 109.890 ;
        RECT 29.810 109.880 29.980 109.900 ;
        RECT -9.060 109.830 -8.890 109.860 ;
        RECT -10.380 109.720 -9.950 109.740 ;
        RECT -10.400 109.550 -9.950 109.720 ;
        RECT 11.190 109.600 11.360 109.650 ;
        RECT -10.380 109.530 -9.950 109.550 ;
        RECT 11.160 109.380 11.380 109.600 ;
        RECT 11.190 109.320 11.360 109.380 ;
        RECT 11.710 109.240 12.040 109.420 ;
        RECT 14.850 109.410 15.020 109.460 ;
        RECT 12.290 109.240 14.450 109.410 ;
        RECT 14.690 109.240 15.020 109.410 ;
        RECT 15.310 109.270 15.520 109.600 ;
        RECT -10.190 109.190 -9.870 109.230 ;
        RECT -10.190 109.170 -9.860 109.190 ;
        RECT -10.190 108.970 -9.570 109.170 ;
        RECT -9.740 108.840 -9.570 108.970 ;
        RECT -9.060 109.130 -8.890 109.170 ;
        RECT -9.060 109.090 -8.570 109.130 ;
        RECT -9.060 108.900 -8.560 109.090 ;
        RECT -9.060 108.870 -8.570 108.900 ;
        RECT -9.060 108.840 -8.890 108.870 ;
        RECT 11.740 108.800 12.010 109.240 ;
        RECT 13.220 108.980 13.550 109.240 ;
        RECT 14.760 109.100 15.020 109.240 ;
        RECT 15.760 109.100 15.940 109.540 ;
        RECT 17.360 109.440 17.750 109.490 ;
        RECT 16.490 109.380 17.750 109.440 ;
        RECT 16.490 109.270 17.830 109.380 ;
        RECT 17.360 109.210 17.830 109.270 ;
        RECT 18.300 109.230 19.260 109.400 ;
        RECT 17.360 109.200 17.740 109.210 ;
        RECT 11.780 108.790 12.010 108.800 ;
        RECT 14.760 108.930 15.940 109.100 ;
        RECT 14.760 108.790 15.020 108.930 ;
        RECT -10.380 108.730 -9.950 108.750 ;
        RECT -10.400 108.560 -9.950 108.730 ;
        RECT 11.780 108.620 12.540 108.790 ;
        RECT 12.790 108.620 13.960 108.790 ;
        RECT 14.200 108.760 15.020 108.790 ;
        RECT 14.200 108.620 15.310 108.760 ;
        RECT -8.450 108.600 -8.220 108.610 ;
        RECT -10.380 108.540 -9.950 108.560 ;
        RECT -8.530 108.430 -8.200 108.600 ;
        RECT 13.190 108.520 13.540 108.620 ;
        RECT 14.850 108.590 15.310 108.620 ;
        RECT 15.760 108.750 16.950 108.760 ;
        RECT 15.760 108.590 17.240 108.750 ;
        RECT 15.800 108.570 17.240 108.590 ;
        RECT 16.780 108.530 17.240 108.570 ;
        RECT 16.950 108.510 17.240 108.530 ;
        RECT 17.570 108.440 17.740 109.200 ;
        RECT 19.080 108.770 19.260 109.230 ;
        RECT 20.250 109.220 20.420 109.640 ;
        RECT 21.060 109.520 21.300 109.550 ;
        RECT 20.730 109.350 21.300 109.520 ;
        RECT 21.540 109.350 22.880 109.520 ;
        RECT 23.330 109.350 24.290 109.520 ;
        RECT 21.060 109.310 21.300 109.350 ;
        RECT 23.840 109.340 24.010 109.350 ;
        RECT 20.180 109.000 20.350 109.040 ;
        RECT 20.120 108.830 20.350 109.000 ;
        RECT 17.940 108.590 18.540 108.760 ;
        RECT 19.000 108.600 19.330 108.770 ;
        RECT 17.940 108.440 18.390 108.590 ;
        RECT 20.180 108.480 20.350 108.830 ;
        RECT 20.520 108.900 20.710 108.920 ;
        RECT 23.470 108.900 23.810 109.080 ;
        RECT 20.520 108.730 21.080 108.900 ;
        RECT 21.540 108.730 24.290 108.900 ;
        RECT 20.520 108.690 20.710 108.730 ;
        RECT 24.820 108.660 24.990 109.590 ;
        RECT 25.220 108.750 25.390 109.640 ;
        RECT 27.440 109.570 27.620 109.760 ;
        RECT 26.990 108.760 27.260 109.090 ;
        RECT 27.050 108.470 27.250 108.760 ;
        RECT 27.060 108.460 27.250 108.470 ;
        RECT -8.450 108.420 -8.220 108.430 ;
        RECT 26.680 108.290 26.890 108.300 ;
        RECT -10.190 108.200 -9.870 108.240 ;
        RECT -10.190 108.180 -9.860 108.200 ;
        RECT -10.190 107.980 -9.570 108.180 ;
        RECT -9.740 107.850 -9.570 107.980 ;
        RECT -9.060 108.140 -8.890 108.180 ;
        RECT -9.060 108.100 -8.570 108.140 ;
        RECT -9.060 107.910 -8.560 108.100 ;
        RECT -9.060 107.880 -8.570 107.910 ;
        RECT -9.060 107.850 -8.890 107.880 ;
        RECT 11.190 107.850 11.360 107.900 ;
        RECT -10.380 107.740 -9.950 107.760 ;
        RECT -10.400 107.570 -9.950 107.740 ;
        RECT 11.160 107.630 11.380 107.850 ;
        RECT 11.190 107.570 11.360 107.630 ;
        RECT -10.380 107.550 -9.950 107.570 ;
        RECT 11.710 107.490 12.040 107.670 ;
        RECT 14.850 107.660 15.020 107.710 ;
        RECT 12.290 107.490 14.450 107.660 ;
        RECT 14.690 107.490 15.020 107.660 ;
        RECT 15.310 107.520 15.520 107.850 ;
        RECT 11.740 107.050 12.010 107.490 ;
        RECT 13.220 107.230 13.550 107.490 ;
        RECT 14.760 107.350 15.020 107.490 ;
        RECT 15.760 107.350 15.940 107.790 ;
        RECT 17.360 107.690 17.750 107.740 ;
        RECT 20.180 107.720 20.350 108.070 ;
        RECT 16.490 107.630 17.750 107.690 ;
        RECT 16.490 107.520 17.830 107.630 ;
        RECT 17.360 107.460 17.830 107.520 ;
        RECT 18.300 107.480 19.260 107.650 ;
        RECT 20.120 107.550 20.350 107.720 ;
        RECT 20.520 107.820 20.710 107.860 ;
        RECT 20.520 107.650 21.080 107.820 ;
        RECT 21.540 107.650 24.290 107.820 ;
        RECT 20.520 107.630 20.710 107.650 ;
        RECT 20.180 107.510 20.350 107.550 ;
        RECT 17.360 107.450 17.740 107.460 ;
        RECT 11.780 107.040 12.010 107.050 ;
        RECT 14.760 107.180 15.940 107.350 ;
        RECT 14.760 107.040 15.020 107.180 ;
        RECT 11.780 106.870 12.540 107.040 ;
        RECT 12.790 106.870 13.960 107.040 ;
        RECT 14.200 107.010 15.020 107.040 ;
        RECT 14.200 106.870 15.310 107.010 ;
        RECT 13.190 106.770 13.540 106.870 ;
        RECT 14.850 106.840 15.310 106.870 ;
        RECT 15.760 107.000 16.950 107.010 ;
        RECT 15.760 106.840 17.240 107.000 ;
        RECT 15.800 106.820 17.240 106.840 ;
        RECT 16.780 106.780 17.240 106.820 ;
        RECT 16.950 106.760 17.240 106.780 ;
        RECT 17.570 106.690 17.740 107.450 ;
        RECT 19.080 107.020 19.260 107.480 ;
        RECT 23.470 107.470 23.810 107.650 ;
        RECT 17.940 106.840 18.540 107.010 ;
        RECT 19.000 106.850 19.330 107.020 ;
        RECT 20.250 106.910 20.420 107.330 ;
        RECT 21.060 107.200 21.300 107.240 ;
        RECT 23.840 107.200 24.010 107.210 ;
        RECT 20.730 107.030 21.300 107.200 ;
        RECT 21.540 107.030 22.880 107.200 ;
        RECT 23.330 107.030 24.290 107.200 ;
        RECT 21.060 107.000 21.300 107.030 ;
        RECT 24.820 106.960 24.990 107.890 ;
        RECT 25.220 106.910 25.390 107.800 ;
        RECT 26.680 107.710 26.900 108.290 ;
        RECT 27.450 107.960 27.620 109.570 ;
        RECT 28.280 109.300 28.450 109.660 ;
        RECT 28.870 109.570 29.220 109.740 ;
        RECT 29.410 109.720 29.600 109.770 ;
        RECT 30.310 109.740 30.480 110.310 ;
        RECT 34.590 110.080 34.780 110.480 ;
        RECT 40.770 110.080 40.960 110.480 ;
        RECT 47.100 110.390 47.270 111.300 ;
        RECT 47.930 110.480 48.100 112.090 ;
        RECT 48.650 111.760 48.870 112.340 ;
        RECT 48.660 111.750 48.870 111.760 ;
        RECT 49.660 111.640 49.840 112.570 ;
        RECT 51.480 112.490 51.910 112.750 ;
        RECT 50.390 112.310 50.720 112.480 ;
        RECT 51.710 112.460 51.910 112.490 ;
        RECT 50.470 112.170 50.720 112.310 ;
        RECT 50.470 111.910 50.950 112.170 ;
        RECT 51.300 112.100 51.470 112.140 ;
        RECT 51.710 112.100 51.910 112.130 ;
        RECT 49.540 111.610 49.860 111.640 ;
        RECT 48.300 111.580 48.490 111.590 ;
        RECT 48.300 111.290 48.500 111.580 ;
        RECT 49.540 111.420 49.870 111.610 ;
        RECT 49.540 111.380 49.860 111.420 ;
        RECT 48.290 110.960 48.580 111.290 ;
        RECT 47.930 110.290 48.110 110.480 ;
        RECT 34.590 110.070 34.970 110.080 ;
        RECT 31.230 109.890 34.970 110.070 ;
        RECT 34.590 109.850 34.970 109.890 ;
        RECT 40.580 110.070 40.960 110.080 ;
        RECT 40.580 109.890 44.320 110.070 ;
        RECT 40.580 109.850 40.960 109.890 ;
        RECT 29.410 109.710 29.640 109.720 ;
        RECT 30.220 109.710 30.560 109.740 ;
        RECT 29.410 109.570 30.560 109.710 ;
        RECT 28.950 109.360 29.140 109.570 ;
        RECT 29.410 109.540 30.390 109.570 ;
        RECT 29.550 109.510 30.390 109.540 ;
        RECT 34.590 109.470 34.780 109.850 ;
        RECT 28.040 109.260 28.450 109.300 ;
        RECT 28.030 109.070 28.450 109.260 ;
        RECT 36.830 109.180 37.380 109.610 ;
        RECT 38.170 109.180 38.720 109.610 ;
        RECT 40.770 109.470 40.960 109.850 ;
        RECT 28.040 109.040 28.450 109.070 ;
        RECT 28.280 107.970 28.450 109.040 ;
        RECT 28.870 108.850 31.800 108.950 ;
        RECT 28.870 108.780 31.860 108.850 ;
        RECT 30.890 108.460 31.060 108.520 ;
        RECT 30.870 108.250 31.080 108.460 ;
        RECT 29.400 108.160 29.590 108.190 ;
        RECT 30.890 108.180 31.060 108.250 ;
        RECT 31.630 108.160 31.860 108.780 ;
        RECT 41.800 108.160 42.030 108.890 ;
        RECT 47.100 108.800 47.270 109.660 ;
        RECT 46.940 108.540 47.270 108.800 ;
        RECT 28.870 107.990 29.590 108.160 ;
        RECT 29.400 107.960 29.590 107.990 ;
        RECT 29.760 107.990 30.570 108.160 ;
        RECT 26.680 107.680 26.890 107.710 ;
        RECT 26.690 107.330 26.890 107.680 ;
        RECT 28.970 107.650 29.160 107.680 ;
        RECT 29.760 107.650 29.950 107.990 ;
        RECT 47.100 107.970 47.270 108.540 ;
        RECT 47.930 109.570 48.110 109.760 ;
        RECT 47.930 107.960 48.100 109.570 ;
        RECT 48.290 108.760 48.580 109.090 ;
        RECT 48.300 108.470 48.500 108.760 ;
        RECT 48.300 108.460 48.490 108.470 ;
        RECT 48.660 108.290 48.870 108.300 ;
        RECT 48.650 107.710 48.870 108.290 ;
        RECT 28.170 107.410 28.700 107.580 ;
        RECT 28.970 107.470 29.950 107.650 ;
        RECT 48.660 107.680 48.870 107.710 ;
        RECT 28.970 107.450 29.160 107.470 ;
        RECT 46.850 107.410 47.380 107.580 ;
        RECT 48.660 107.330 48.860 107.680 ;
        RECT 49.660 107.470 49.840 111.380 ;
        RECT 50.470 110.530 50.640 111.910 ;
        RECT 51.300 111.840 51.910 112.100 ;
        RECT 51.300 111.810 51.470 111.840 ;
        RECT 51.710 111.800 51.910 111.840 ;
        RECT 52.300 111.800 52.850 112.790 ;
        RECT 53.670 112.640 54.300 112.810 ;
        RECT 53.670 112.540 54.060 112.640 ;
        RECT 53.670 112.510 54.050 112.540 ;
        RECT 53.670 112.360 54.030 112.510 ;
        RECT 53.320 112.190 54.030 112.360 ;
        RECT 53.320 111.440 54.020 111.750 ;
        RECT 51.300 111.250 51.470 111.280 ;
        RECT 51.710 111.250 51.910 111.290 ;
        RECT 51.300 110.990 51.910 111.250 ;
        RECT 51.300 110.950 51.470 110.990 ;
        RECT 51.710 110.960 51.910 110.990 ;
        RECT 51.710 110.600 51.910 110.630 ;
        RECT 50.270 110.330 50.590 110.360 ;
        RECT 51.480 110.340 51.910 110.600 ;
        RECT 50.270 110.140 50.600 110.330 ;
        RECT 51.710 110.300 51.910 110.340 ;
        RECT 52.300 110.300 52.850 111.290 ;
        RECT 53.170 111.210 54.020 111.440 ;
        RECT 53.320 110.870 54.020 111.210 ;
        RECT 53.780 110.510 54.100 110.550 ;
        RECT 53.780 110.450 54.110 110.510 ;
        RECT 53.310 110.320 54.110 110.450 ;
        RECT 53.310 110.290 54.100 110.320 ;
        RECT 53.310 110.270 54.010 110.290 ;
        RECT 79.190 110.260 79.510 110.290 ;
        RECT 80.760 110.260 81.080 110.290 ;
        RECT 50.270 110.100 50.590 110.140 ;
        RECT 50.270 110.020 50.440 110.100 ;
        RECT 50.220 109.850 50.440 110.020 ;
        RECT 77.970 109.920 78.140 110.200 ;
        RECT 79.190 110.070 79.520 110.260 ;
        RECT 80.200 110.120 80.390 110.140 ;
        RECT 79.190 110.030 79.510 110.070 ;
        RECT 77.970 109.880 78.180 109.920 ;
        RECT 77.970 109.860 78.200 109.880 ;
        RECT 79.320 109.870 79.490 110.030 ;
        RECT 79.930 109.950 80.390 110.120 ;
        RECT 80.760 110.070 81.090 110.260 ;
        RECT 81.330 110.120 81.520 110.150 ;
        RECT 80.760 110.030 81.080 110.070 ;
        RECT 80.180 109.940 80.390 109.950 ;
        RECT 80.200 109.910 80.390 109.940 ;
        RECT 80.820 109.870 80.990 110.030 ;
        RECT 81.330 109.950 81.770 110.120 ;
        RECT 81.330 109.920 81.520 109.950 ;
        RECT 50.220 109.690 50.390 109.850 ;
        RECT 77.970 109.840 78.230 109.860 ;
        RECT 53.770 109.790 54.090 109.830 ;
        RECT 77.970 109.790 78.310 109.840 ;
        RECT 51.710 109.750 51.910 109.790 ;
        RECT 50.750 109.430 50.940 109.550 ;
        RECT 51.480 109.490 51.910 109.750 ;
        RECT 51.710 109.460 51.910 109.490 ;
        RECT 50.390 109.320 50.940 109.430 ;
        RECT 50.390 109.260 50.930 109.320 ;
        RECT 50.470 107.480 50.640 109.260 ;
        RECT 51.300 109.100 51.470 109.140 ;
        RECT 51.710 109.100 51.910 109.130 ;
        RECT 51.300 108.840 51.910 109.100 ;
        RECT 51.300 108.810 51.470 108.840 ;
        RECT 51.710 108.800 51.910 108.840 ;
        RECT 52.300 108.800 52.850 109.790 ;
        RECT 53.310 109.610 54.100 109.790 ;
        RECT 77.970 109.730 78.460 109.790 ;
        RECT 77.970 109.700 78.480 109.730 ;
        RECT 78.010 109.670 78.480 109.700 ;
        RECT 78.140 109.620 78.480 109.670 ;
        RECT 78.260 109.610 78.480 109.620 ;
        RECT 53.770 109.600 54.100 109.610 ;
        RECT 53.770 109.570 54.090 109.600 ;
        RECT 78.270 109.580 78.480 109.610 ;
        RECT 78.290 109.500 78.480 109.580 ;
        RECT 79.650 109.500 79.980 109.620 ;
        RECT 82.050 109.530 82.220 110.210 ;
        RECT 77.800 109.450 77.970 109.470 ;
        RECT 53.320 108.850 54.020 109.190 ;
        RECT 77.780 109.020 77.990 109.450 ;
        RECT 78.290 109.330 78.810 109.500 ;
        RECT 78.290 109.300 78.480 109.330 ;
        RECT 79.160 109.320 81.060 109.500 ;
        RECT 81.790 109.490 82.220 109.530 ;
        RECT 81.440 109.330 82.220 109.490 ;
        RECT 81.440 109.320 81.980 109.330 ;
        RECT 81.790 109.300 81.980 109.320 ;
        RECT 53.170 108.620 54.020 108.850 ;
        RECT 53.320 108.310 54.020 108.620 ;
        RECT 77.780 108.300 77.990 108.730 ;
        RECT 78.290 108.420 78.480 108.450 ;
        RECT 81.790 108.430 81.980 108.450 ;
        RECT 51.300 108.250 51.470 108.280 ;
        RECT 51.710 108.250 51.910 108.290 ;
        RECT 51.300 107.990 51.910 108.250 ;
        RECT 51.300 107.950 51.470 107.990 ;
        RECT 51.710 107.960 51.910 107.990 ;
        RECT 51.710 107.600 51.910 107.630 ;
        RECT 51.480 107.340 51.910 107.600 ;
        RECT 51.710 107.300 51.910 107.340 ;
        RECT 52.300 107.300 52.850 108.290 ;
        RECT 77.800 108.280 77.970 108.300 ;
        RECT 78.290 108.250 78.810 108.420 ;
        RECT 79.160 108.250 81.060 108.430 ;
        RECT 81.440 108.420 81.980 108.430 ;
        RECT 81.440 108.260 82.220 108.420 ;
        RECT 78.290 108.170 78.480 108.250 ;
        RECT 78.270 108.140 78.480 108.170 ;
        RECT 78.260 108.130 78.480 108.140 ;
        RECT 79.650 108.130 79.980 108.250 ;
        RECT 81.790 108.220 82.220 108.260 ;
        RECT 78.140 108.080 78.480 108.130 ;
        RECT 78.010 108.050 78.480 108.080 ;
        RECT 77.970 108.020 78.480 108.050 ;
        RECT 77.970 107.960 78.460 108.020 ;
        RECT 77.970 107.910 78.310 107.960 ;
        RECT 77.970 107.890 78.230 107.910 ;
        RECT 77.970 107.870 78.200 107.890 ;
        RECT 53.320 107.700 54.030 107.870 ;
        RECT 53.670 107.420 54.030 107.700 ;
        RECT 77.970 107.830 78.180 107.870 ;
        RECT 77.970 107.550 78.140 107.830 ;
        RECT 79.320 107.720 79.490 107.880 ;
        RECT 80.200 107.810 80.390 107.840 ;
        RECT 80.180 107.800 80.390 107.810 ;
        RECT 79.190 107.680 79.510 107.720 ;
        RECT 79.190 107.490 79.520 107.680 ;
        RECT 79.930 107.630 80.390 107.800 ;
        RECT 80.820 107.720 80.990 107.880 ;
        RECT 81.330 107.800 81.520 107.830 ;
        RECT 80.200 107.610 80.390 107.630 ;
        RECT 80.760 107.680 81.080 107.720 ;
        RECT 80.760 107.490 81.090 107.680 ;
        RECT 81.330 107.630 81.770 107.800 ;
        RECT 81.330 107.600 81.520 107.630 ;
        RECT 82.050 107.540 82.220 108.220 ;
        RECT 79.190 107.460 79.510 107.490 ;
        RECT 80.760 107.460 81.080 107.490 ;
        RECT 53.670 107.250 54.300 107.420 ;
        RECT 79.190 107.060 79.510 107.090 ;
        RECT 80.760 107.060 81.080 107.090 ;
        RECT 50.240 106.970 50.410 107.020 ;
        RECT 17.940 106.690 18.390 106.840 ;
        RECT 11.190 106.100 11.360 106.150 ;
        RECT 11.160 105.880 11.380 106.100 ;
        RECT 11.190 105.820 11.360 105.880 ;
        RECT 11.710 105.740 12.040 105.920 ;
        RECT 14.850 105.910 15.020 105.960 ;
        RECT 12.290 105.740 14.450 105.910 ;
        RECT 14.690 105.740 15.020 105.910 ;
        RECT 15.310 105.770 15.520 106.100 ;
        RECT -143.430 105.550 -142.910 105.570 ;
        RECT -149.480 104.070 -143.770 104.080 ;
        RECT -149.560 103.900 -143.770 104.070 ;
        RECT -149.470 103.890 -143.770 103.900 ;
        RECT -144.000 103.820 -143.830 103.890 ;
        RECT -143.430 103.770 -142.900 105.550 ;
        RECT 11.740 105.300 12.010 105.740 ;
        RECT 13.220 105.480 13.550 105.740 ;
        RECT 14.760 105.600 15.020 105.740 ;
        RECT 15.760 105.600 15.940 106.040 ;
        RECT 20.250 106.020 20.420 106.440 ;
        RECT 21.060 106.320 21.300 106.350 ;
        RECT 20.730 106.150 21.300 106.320 ;
        RECT 21.540 106.150 22.880 106.320 ;
        RECT 23.330 106.150 24.290 106.320 ;
        RECT 21.060 106.110 21.300 106.150 ;
        RECT 23.840 106.140 24.010 106.150 ;
        RECT 17.360 105.940 17.750 105.990 ;
        RECT 16.490 105.880 17.750 105.940 ;
        RECT 16.490 105.770 17.830 105.880 ;
        RECT 17.360 105.710 17.830 105.770 ;
        RECT 18.300 105.730 19.260 105.900 ;
        RECT 20.180 105.800 20.350 105.840 ;
        RECT 17.360 105.700 17.740 105.710 ;
        RECT 11.780 105.290 12.010 105.300 ;
        RECT 14.760 105.430 15.940 105.600 ;
        RECT 14.760 105.290 15.020 105.430 ;
        RECT 11.780 105.120 12.540 105.290 ;
        RECT 12.790 105.120 13.960 105.290 ;
        RECT 14.200 105.260 15.020 105.290 ;
        RECT 14.200 105.120 15.310 105.260 ;
        RECT 13.190 105.020 13.540 105.120 ;
        RECT 14.850 105.090 15.310 105.120 ;
        RECT 15.760 105.250 16.950 105.260 ;
        RECT 15.760 105.090 17.240 105.250 ;
        RECT 15.800 105.070 17.240 105.090 ;
        RECT 16.780 105.030 17.240 105.070 ;
        RECT 16.950 105.010 17.240 105.030 ;
        RECT 17.570 104.940 17.740 105.700 ;
        RECT 19.080 105.270 19.260 105.730 ;
        RECT 20.120 105.630 20.350 105.800 ;
        RECT 20.180 105.280 20.350 105.630 ;
        RECT 20.520 105.700 20.710 105.720 ;
        RECT 23.470 105.700 23.810 105.880 ;
        RECT 20.520 105.530 21.080 105.700 ;
        RECT 21.540 105.530 24.290 105.700 ;
        RECT 20.520 105.490 20.710 105.530 ;
        RECT 24.820 105.460 24.990 106.390 ;
        RECT 25.220 105.550 25.390 106.440 ;
        RECT 26.700 106.340 26.900 106.690 ;
        RECT 28.180 106.440 28.710 106.610 ;
        RECT 26.690 106.310 26.900 106.340 ;
        RECT 26.690 105.730 26.910 106.310 ;
        RECT 26.690 105.720 26.900 105.730 ;
        RECT 27.070 105.550 27.260 105.560 ;
        RECT 17.940 105.090 18.540 105.260 ;
        RECT 19.000 105.100 19.330 105.270 ;
        RECT 27.060 105.260 27.260 105.550 ;
        RECT 17.940 104.940 18.390 105.090 ;
        RECT 26.980 104.930 27.270 105.260 ;
        RECT 20.180 104.520 20.350 104.870 ;
        RECT 11.190 104.350 11.360 104.400 ;
        RECT 20.120 104.350 20.350 104.520 ;
        RECT 20.520 104.620 20.710 104.660 ;
        RECT 20.520 104.450 21.080 104.620 ;
        RECT 21.540 104.450 24.290 104.620 ;
        RECT 20.520 104.430 20.710 104.450 ;
        RECT 11.160 104.130 11.380 104.350 ;
        RECT 11.190 104.070 11.360 104.130 ;
        RECT 11.710 103.990 12.040 104.170 ;
        RECT 14.850 104.160 15.020 104.210 ;
        RECT 12.290 103.990 14.450 104.160 ;
        RECT 14.690 103.990 15.020 104.160 ;
        RECT 15.310 104.020 15.520 104.350 ;
        RECT 20.180 104.310 20.350 104.350 ;
        RECT -143.420 103.750 -142.900 103.770 ;
        RECT -150.440 103.030 -148.000 103.320 ;
        RECT -143.420 103.240 -142.910 103.750 ;
        RECT 11.740 103.550 12.010 103.990 ;
        RECT 13.220 103.730 13.550 103.990 ;
        RECT 14.760 103.850 15.020 103.990 ;
        RECT 15.760 103.850 15.940 104.290 ;
        RECT 23.470 104.270 23.810 104.450 ;
        RECT 17.360 104.190 17.750 104.240 ;
        RECT 16.490 104.130 17.750 104.190 ;
        RECT 16.490 104.020 17.830 104.130 ;
        RECT 17.360 103.960 17.830 104.020 ;
        RECT 18.300 103.980 19.260 104.150 ;
        RECT 17.360 103.950 17.740 103.960 ;
        RECT 11.780 103.540 12.010 103.550 ;
        RECT 14.760 103.680 15.940 103.850 ;
        RECT 14.760 103.540 15.020 103.680 ;
        RECT 11.780 103.370 12.540 103.540 ;
        RECT 12.790 103.370 13.960 103.540 ;
        RECT 14.200 103.510 15.020 103.540 ;
        RECT 14.200 103.370 15.310 103.510 ;
        RECT 13.190 103.270 13.540 103.370 ;
        RECT 14.850 103.340 15.310 103.370 ;
        RECT 15.760 103.500 16.950 103.510 ;
        RECT 15.760 103.340 17.240 103.500 ;
        RECT 15.800 103.320 17.240 103.340 ;
        RECT 16.780 103.280 17.240 103.320 ;
        RECT 16.950 103.260 17.240 103.280 ;
        RECT -143.420 103.030 -142.890 103.240 ;
        RECT 17.570 103.190 17.740 103.950 ;
        RECT 19.080 103.520 19.260 103.980 ;
        RECT 20.250 103.710 20.420 104.130 ;
        RECT 21.060 104.000 21.300 104.040 ;
        RECT 23.840 104.000 24.010 104.010 ;
        RECT 20.730 103.830 21.300 104.000 ;
        RECT 21.540 103.830 22.880 104.000 ;
        RECT 23.330 103.830 24.290 104.000 ;
        RECT 21.060 103.800 21.300 103.830 ;
        RECT 24.820 103.760 24.990 104.690 ;
        RECT 25.220 103.710 25.390 104.600 ;
        RECT 27.460 104.450 27.630 106.060 ;
        RECT 27.450 104.260 27.630 104.450 ;
        RECT 28.290 105.530 28.460 106.050 ;
        RECT 30.900 106.010 35.960 106.840 ;
        RECT 50.240 106.710 50.800 106.970 ;
        RECT 51.710 106.720 51.910 106.760 ;
        RECT 50.240 106.690 50.410 106.710 ;
        RECT 46.850 106.440 47.380 106.610 ;
        RECT 48.660 106.340 48.860 106.690 ;
        RECT 48.660 106.310 48.870 106.340 ;
        RECT 35.410 105.930 35.890 106.010 ;
        RECT 28.290 105.270 28.620 105.530 ;
        RECT 28.290 104.360 28.460 105.270 ;
        RECT 33.530 105.070 33.760 105.760 ;
        RECT 35.410 105.680 35.880 105.930 ;
        RECT 36.840 104.880 37.390 105.310 ;
        RECT 38.170 104.880 38.720 105.310 ;
        RECT 41.800 105.070 42.030 105.760 ;
        RECT 47.100 105.530 47.270 106.050 ;
        RECT 46.940 105.270 47.270 105.530 ;
        RECT 34.600 104.040 34.990 104.450 ;
        RECT 31.240 103.860 34.990 104.040 ;
        RECT 27.450 103.540 27.630 103.730 ;
        RECT 17.940 103.340 18.540 103.510 ;
        RECT 19.000 103.350 19.330 103.520 ;
        RECT 17.940 103.190 18.390 103.340 ;
        RECT -150.440 102.550 -142.890 103.030 ;
        RECT 26.980 102.730 27.270 103.060 ;
        RECT -150.440 102.520 -143.080 102.550 ;
        RECT 27.060 102.440 27.260 102.730 ;
        RECT 27.070 102.430 27.260 102.440 ;
        RECT 26.690 102.260 26.900 102.270 ;
        RECT 26.690 101.680 26.910 102.260 ;
        RECT 27.460 101.930 27.630 103.540 ;
        RECT 28.290 102.770 28.460 103.630 ;
        RECT 34.600 103.440 34.990 103.860 ;
        RECT 40.540 104.040 40.960 104.450 ;
        RECT 47.100 104.360 47.270 105.270 ;
        RECT 47.930 104.450 48.100 106.060 ;
        RECT 48.650 105.730 48.870 106.310 ;
        RECT 48.660 105.720 48.870 105.730 ;
        RECT 49.660 105.610 49.840 106.540 ;
        RECT 51.480 106.460 51.910 106.720 ;
        RECT 50.390 106.280 50.720 106.450 ;
        RECT 51.710 106.430 51.910 106.460 ;
        RECT 50.470 106.140 50.720 106.280 ;
        RECT 50.470 105.880 50.950 106.140 ;
        RECT 51.300 106.070 51.470 106.110 ;
        RECT 51.710 106.070 51.910 106.100 ;
        RECT 49.540 105.580 49.860 105.610 ;
        RECT 48.300 105.550 48.490 105.560 ;
        RECT 48.300 105.260 48.500 105.550 ;
        RECT 49.540 105.390 49.870 105.580 ;
        RECT 49.540 105.350 49.860 105.390 ;
        RECT 48.290 104.930 48.580 105.260 ;
        RECT 47.930 104.260 48.110 104.450 ;
        RECT 40.540 103.860 44.320 104.040 ;
        RECT 36.840 103.150 37.390 103.580 ;
        RECT 38.170 103.150 38.720 103.580 ;
        RECT 40.540 103.440 40.960 103.860 ;
        RECT 28.290 102.510 28.620 102.770 ;
        RECT 28.290 101.940 28.460 102.510 ;
        RECT 33.530 102.130 33.760 102.860 ;
        RECT 35.570 102.000 35.910 102.250 ;
        RECT 41.800 102.130 42.030 102.860 ;
        RECT 47.100 102.770 47.270 103.630 ;
        RECT 46.940 102.510 47.270 102.770 ;
        RECT 35.570 101.920 35.920 102.000 ;
        RECT 47.100 101.940 47.270 102.510 ;
        RECT 47.930 103.540 48.110 103.730 ;
        RECT 47.930 101.930 48.100 103.540 ;
        RECT 48.290 102.730 48.580 103.060 ;
        RECT 48.300 102.440 48.500 102.730 ;
        RECT 48.300 102.430 48.490 102.440 ;
        RECT 48.660 102.260 48.870 102.270 ;
        RECT 26.690 101.650 26.900 101.680 ;
        RECT -150.440 100.760 -142.910 101.310 ;
        RECT 26.700 101.300 26.900 101.650 ;
        RECT 28.180 101.380 28.710 101.550 ;
        RECT 30.870 101.070 35.920 101.920 ;
        RECT 48.650 101.680 48.870 102.260 ;
        RECT 48.660 101.650 48.870 101.680 ;
        RECT 46.850 101.380 47.380 101.550 ;
        RECT 48.660 101.300 48.860 101.650 ;
        RECT 49.660 101.440 49.840 105.350 ;
        RECT 50.470 104.500 50.640 105.880 ;
        RECT 51.300 105.810 51.910 106.070 ;
        RECT 51.300 105.780 51.470 105.810 ;
        RECT 51.710 105.770 51.910 105.810 ;
        RECT 52.300 105.770 52.850 106.760 ;
        RECT 53.670 106.610 54.300 106.780 ;
        RECT 77.970 106.720 78.140 107.000 ;
        RECT 79.190 106.870 79.520 107.060 ;
        RECT 80.200 106.920 80.390 106.940 ;
        RECT 79.190 106.830 79.510 106.870 ;
        RECT 77.970 106.680 78.180 106.720 ;
        RECT 77.970 106.660 78.200 106.680 ;
        RECT 79.320 106.670 79.490 106.830 ;
        RECT 79.930 106.750 80.390 106.920 ;
        RECT 80.760 106.870 81.090 107.060 ;
        RECT 81.330 106.920 81.520 106.950 ;
        RECT 80.760 106.830 81.080 106.870 ;
        RECT 80.180 106.740 80.390 106.750 ;
        RECT 80.200 106.710 80.390 106.740 ;
        RECT 80.820 106.670 80.990 106.830 ;
        RECT 81.330 106.750 81.770 106.920 ;
        RECT 81.330 106.720 81.520 106.750 ;
        RECT 77.970 106.640 78.230 106.660 ;
        RECT 53.670 106.510 54.060 106.610 ;
        RECT 77.970 106.590 78.310 106.640 ;
        RECT 77.970 106.530 78.460 106.590 ;
        RECT 53.670 106.480 54.050 106.510 ;
        RECT 77.970 106.500 78.480 106.530 ;
        RECT 53.670 106.330 54.030 106.480 ;
        RECT 78.010 106.470 78.480 106.500 ;
        RECT 78.140 106.420 78.480 106.470 ;
        RECT 78.260 106.410 78.480 106.420 ;
        RECT 78.270 106.380 78.480 106.410 ;
        RECT 53.320 106.160 54.030 106.330 ;
        RECT 78.290 106.300 78.480 106.380 ;
        RECT 79.650 106.300 79.980 106.420 ;
        RECT 82.050 106.330 82.220 107.010 ;
        RECT 77.800 106.250 77.970 106.270 ;
        RECT 77.780 105.820 77.990 106.250 ;
        RECT 78.290 106.130 78.810 106.300 ;
        RECT 78.290 106.100 78.480 106.130 ;
        RECT 79.160 106.120 81.060 106.300 ;
        RECT 81.790 106.290 82.220 106.330 ;
        RECT 81.440 106.130 82.220 106.290 ;
        RECT 81.440 106.120 81.980 106.130 ;
        RECT 81.790 106.100 81.980 106.120 ;
        RECT 53.320 105.410 54.020 105.720 ;
        RECT 51.300 105.220 51.470 105.250 ;
        RECT 51.710 105.220 51.910 105.260 ;
        RECT 51.300 104.960 51.910 105.220 ;
        RECT 51.300 104.920 51.470 104.960 ;
        RECT 51.710 104.930 51.910 104.960 ;
        RECT 51.710 104.570 51.910 104.600 ;
        RECT 50.270 104.300 50.590 104.330 ;
        RECT 51.480 104.310 51.910 104.570 ;
        RECT 50.270 104.110 50.600 104.300 ;
        RECT 51.710 104.270 51.910 104.310 ;
        RECT 52.300 104.270 52.850 105.260 ;
        RECT 53.170 105.180 54.020 105.410 ;
        RECT 53.320 104.840 54.020 105.180 ;
        RECT 77.780 105.100 77.990 105.530 ;
        RECT 78.290 105.220 78.480 105.250 ;
        RECT 81.790 105.230 81.980 105.250 ;
        RECT 77.800 105.080 77.970 105.100 ;
        RECT 78.290 105.050 78.810 105.220 ;
        RECT 79.160 105.050 81.060 105.230 ;
        RECT 81.440 105.220 81.980 105.230 ;
        RECT 81.440 105.060 82.220 105.220 ;
        RECT 78.290 104.970 78.480 105.050 ;
        RECT 78.270 104.940 78.480 104.970 ;
        RECT 78.260 104.930 78.480 104.940 ;
        RECT 79.650 104.930 79.980 105.050 ;
        RECT 81.790 105.020 82.220 105.060 ;
        RECT 78.140 104.880 78.480 104.930 ;
        RECT 78.010 104.850 78.480 104.880 ;
        RECT 77.970 104.820 78.480 104.850 ;
        RECT 77.970 104.760 78.460 104.820 ;
        RECT 77.970 104.710 78.310 104.760 ;
        RECT 77.970 104.690 78.230 104.710 ;
        RECT 77.970 104.670 78.200 104.690 ;
        RECT 77.970 104.630 78.180 104.670 ;
        RECT 53.780 104.480 54.100 104.520 ;
        RECT 53.780 104.420 54.110 104.480 ;
        RECT 53.310 104.290 54.110 104.420 ;
        RECT 77.970 104.350 78.140 104.630 ;
        RECT 79.320 104.520 79.490 104.680 ;
        RECT 80.200 104.610 80.390 104.640 ;
        RECT 80.180 104.600 80.390 104.610 ;
        RECT 79.190 104.480 79.510 104.520 ;
        RECT 79.190 104.290 79.520 104.480 ;
        RECT 79.930 104.430 80.390 104.600 ;
        RECT 80.820 104.520 80.990 104.680 ;
        RECT 81.330 104.600 81.520 104.630 ;
        RECT 80.200 104.410 80.390 104.430 ;
        RECT 80.760 104.480 81.080 104.520 ;
        RECT 80.760 104.290 81.090 104.480 ;
        RECT 81.330 104.430 81.770 104.600 ;
        RECT 81.330 104.400 81.520 104.430 ;
        RECT 82.050 104.340 82.220 105.020 ;
        RECT 206.500 104.850 207.010 115.210 ;
        RECT 207.180 114.420 213.160 114.650 ;
        RECT 206.500 104.830 207.020 104.850 ;
        RECT 53.310 104.260 54.100 104.290 ;
        RECT 79.190 104.260 79.510 104.290 ;
        RECT 80.760 104.260 81.080 104.290 ;
        RECT 53.310 104.240 54.010 104.260 ;
        RECT 50.270 104.070 50.590 104.110 ;
        RECT 50.270 103.990 50.440 104.070 ;
        RECT 50.220 103.820 50.440 103.990 ;
        RECT 50.220 103.660 50.390 103.820 ;
        RECT 53.770 103.760 54.090 103.800 ;
        RECT 51.710 103.720 51.910 103.760 ;
        RECT 50.750 103.400 50.940 103.520 ;
        RECT 51.480 103.460 51.910 103.720 ;
        RECT 51.710 103.430 51.910 103.460 ;
        RECT 50.390 103.290 50.940 103.400 ;
        RECT 50.390 103.230 50.930 103.290 ;
        RECT 50.470 101.450 50.640 103.230 ;
        RECT 51.300 103.070 51.470 103.110 ;
        RECT 51.710 103.070 51.910 103.100 ;
        RECT 51.300 102.810 51.910 103.070 ;
        RECT 51.300 102.780 51.470 102.810 ;
        RECT 51.710 102.770 51.910 102.810 ;
        RECT 52.300 102.770 52.850 103.760 ;
        RECT 53.310 103.580 54.100 103.760 ;
        RECT 53.770 103.570 54.100 103.580 ;
        RECT 53.770 103.540 54.090 103.570 ;
        RECT 53.320 102.820 54.020 103.160 ;
        RECT 206.490 103.050 207.020 104.830 ;
        RECT 207.420 103.360 213.070 114.420 ;
        RECT 207.360 103.350 213.070 103.360 ;
        RECT 207.360 103.180 213.150 103.350 ;
        RECT 207.360 103.170 213.060 103.180 ;
        RECT 207.420 103.100 207.590 103.170 ;
        RECT 206.490 103.030 207.010 103.050 ;
        RECT 53.170 102.590 54.020 102.820 ;
        RECT 53.320 102.280 54.020 102.590 ;
        RECT 206.500 102.520 207.010 103.030 ;
        RECT 213.520 102.600 214.030 115.210 ;
        RECT 214.270 109.190 215.730 109.230 ;
        RECT 214.260 109.020 215.730 109.190 ;
        RECT 214.270 108.980 215.730 109.020 ;
        RECT 206.480 102.310 207.010 102.520 ;
        RECT 211.590 102.310 214.030 102.600 ;
        RECT 51.300 102.220 51.470 102.250 ;
        RECT 51.710 102.220 51.910 102.260 ;
        RECT 51.300 101.960 51.910 102.220 ;
        RECT 51.300 101.920 51.470 101.960 ;
        RECT 51.710 101.930 51.910 101.960 ;
        RECT 51.710 101.570 51.910 101.600 ;
        RECT 51.480 101.310 51.910 101.570 ;
        RECT 51.710 101.270 51.910 101.310 ;
        RECT 52.300 101.270 52.850 102.260 ;
        RECT 53.320 101.670 54.030 101.840 ;
        RECT 206.480 101.830 214.030 102.310 ;
        RECT 206.670 101.800 214.030 101.830 ;
        RECT 53.670 101.390 54.030 101.670 ;
        RECT 53.670 101.220 54.300 101.390 ;
        RECT -152.130 87.790 -150.650 88.040 ;
        RECT -150.440 87.850 -149.930 100.760 ;
        RECT -143.580 100.750 -142.910 100.760 ;
        RECT -147.280 99.860 -143.820 100.300 ;
        RECT -149.210 99.760 -143.820 99.860 ;
        RECT -149.210 99.690 -143.930 99.760 ;
        RECT -149.210 88.780 -149.040 99.690 ;
        RECT -148.710 99.280 -144.480 99.300 ;
        RECT -148.730 89.170 -144.400 99.280 ;
        RECT -148.670 89.120 -148.500 89.170 ;
        RECT -144.100 88.780 -143.930 99.690 ;
        RECT -149.210 88.610 -143.930 88.780 ;
        RECT -144.170 88.600 -143.930 88.610 ;
        RECT -143.420 87.850 -142.910 100.750 ;
        RECT 206.500 100.040 214.030 100.590 ;
        RECT 206.500 100.030 207.170 100.040 ;
        RECT 11.190 99.470 11.360 99.520 ;
        RECT 11.160 99.250 11.380 99.470 ;
        RECT 11.190 99.190 11.360 99.250 ;
        RECT 11.710 99.110 12.040 99.290 ;
        RECT 14.850 99.280 15.020 99.330 ;
        RECT 12.290 99.110 14.450 99.280 ;
        RECT 14.690 99.110 15.020 99.280 ;
        RECT 15.310 99.140 15.520 99.470 ;
        RECT 11.740 98.670 12.010 99.110 ;
        RECT 13.220 98.850 13.550 99.110 ;
        RECT 14.760 98.970 15.020 99.110 ;
        RECT 15.760 98.970 15.940 99.410 ;
        RECT 17.360 99.310 17.750 99.360 ;
        RECT 16.490 99.250 17.750 99.310 ;
        RECT 16.490 99.140 17.830 99.250 ;
        RECT 17.360 99.080 17.830 99.140 ;
        RECT 18.300 99.100 19.260 99.270 ;
        RECT 17.360 99.070 17.740 99.080 ;
        RECT 11.780 98.660 12.010 98.670 ;
        RECT 14.760 98.800 15.940 98.970 ;
        RECT 14.760 98.660 15.020 98.800 ;
        RECT 11.780 98.490 12.540 98.660 ;
        RECT 12.790 98.490 13.960 98.660 ;
        RECT 14.200 98.630 15.020 98.660 ;
        RECT 14.200 98.490 15.310 98.630 ;
        RECT 13.190 98.390 13.540 98.490 ;
        RECT 14.850 98.460 15.310 98.490 ;
        RECT 15.760 98.620 16.950 98.630 ;
        RECT 15.760 98.460 17.240 98.620 ;
        RECT 15.800 98.440 17.240 98.460 ;
        RECT 16.780 98.400 17.240 98.440 ;
        RECT 16.950 98.380 17.240 98.400 ;
        RECT 17.570 98.310 17.740 99.070 ;
        RECT 19.080 98.640 19.260 99.100 ;
        RECT 20.230 98.750 20.400 99.170 ;
        RECT 21.040 99.050 21.280 99.080 ;
        RECT 20.710 98.880 21.280 99.050 ;
        RECT 21.520 98.880 22.860 99.050 ;
        RECT 23.310 98.880 24.270 99.050 ;
        RECT 21.040 98.840 21.280 98.880 ;
        RECT 23.820 98.870 23.990 98.880 ;
        RECT 17.940 98.460 18.540 98.630 ;
        RECT 19.000 98.470 19.330 98.640 ;
        RECT 20.160 98.530 20.330 98.570 ;
        RECT 17.940 98.310 18.390 98.460 ;
        RECT 20.100 98.360 20.330 98.530 ;
        RECT 20.160 98.010 20.330 98.360 ;
        RECT 20.500 98.430 20.690 98.450 ;
        RECT 23.450 98.430 23.790 98.610 ;
        RECT 20.500 98.260 21.060 98.430 ;
        RECT 21.520 98.260 24.270 98.430 ;
        RECT 20.500 98.220 20.690 98.260 ;
        RECT 24.800 98.190 24.970 99.120 ;
        RECT 25.200 98.280 25.370 99.170 ;
        RECT 28.110 98.760 28.310 99.110 ;
        RECT 29.850 99.030 30.170 99.040 ;
        RECT 29.590 98.860 30.170 99.030 ;
        RECT 29.840 98.810 30.170 98.860 ;
        RECT 29.850 98.780 30.170 98.810 ;
        RECT 45.370 99.030 45.690 99.040 ;
        RECT 45.370 98.860 45.950 99.030 ;
        RECT 45.370 98.810 45.700 98.860 ;
        RECT 45.370 98.780 45.690 98.810 ;
        RECT 28.100 98.730 28.310 98.760 ;
        RECT 47.230 98.760 47.430 99.110 ;
        RECT 28.100 98.140 28.320 98.730 ;
        RECT 28.840 98.140 29.040 98.740 ;
        RECT 29.850 98.450 30.170 98.490 ;
        RECT 29.840 98.410 30.170 98.450 ;
        RECT 29.590 98.240 30.170 98.410 ;
        RECT 29.850 98.230 30.170 98.240 ;
        RECT 45.370 98.450 45.690 98.490 ;
        RECT 45.370 98.410 45.700 98.450 ;
        RECT 45.370 98.240 45.950 98.410 ;
        RECT 45.370 98.230 45.690 98.240 ;
        RECT 46.500 98.140 46.700 98.740 ;
        RECT 47.230 98.730 47.440 98.760 ;
        RECT 47.220 98.140 47.440 98.730 ;
        RECT 11.190 97.720 11.360 97.770 ;
        RECT 11.160 97.500 11.380 97.720 ;
        RECT 11.190 97.440 11.360 97.500 ;
        RECT 11.710 97.360 12.040 97.540 ;
        RECT 14.850 97.530 15.020 97.580 ;
        RECT 12.290 97.360 14.450 97.530 ;
        RECT 14.690 97.360 15.020 97.530 ;
        RECT 15.310 97.390 15.520 97.720 ;
        RECT 11.740 96.920 12.010 97.360 ;
        RECT 13.220 97.100 13.550 97.360 ;
        RECT 14.760 97.220 15.020 97.360 ;
        RECT 15.760 97.220 15.940 97.660 ;
        RECT 17.360 97.560 17.750 97.610 ;
        RECT 16.490 97.500 17.750 97.560 ;
        RECT 16.490 97.390 17.830 97.500 ;
        RECT 17.360 97.330 17.830 97.390 ;
        RECT 18.300 97.350 19.260 97.520 ;
        RECT 17.360 97.320 17.740 97.330 ;
        RECT 11.780 96.910 12.010 96.920 ;
        RECT 14.760 97.050 15.940 97.220 ;
        RECT 14.760 96.910 15.020 97.050 ;
        RECT 11.780 96.740 12.540 96.910 ;
        RECT 12.790 96.740 13.960 96.910 ;
        RECT 14.200 96.880 15.020 96.910 ;
        RECT 14.200 96.740 15.310 96.880 ;
        RECT 13.190 96.640 13.540 96.740 ;
        RECT 14.850 96.710 15.310 96.740 ;
        RECT 15.760 96.870 16.950 96.880 ;
        RECT 15.760 96.710 17.240 96.870 ;
        RECT 15.800 96.690 17.240 96.710 ;
        RECT 16.780 96.650 17.240 96.690 ;
        RECT 16.950 96.630 17.240 96.650 ;
        RECT 17.570 96.560 17.740 97.320 ;
        RECT 19.080 96.890 19.260 97.350 ;
        RECT 20.160 97.250 20.330 97.600 ;
        RECT 20.100 97.080 20.330 97.250 ;
        RECT 20.500 97.350 20.690 97.390 ;
        RECT 20.500 97.180 21.060 97.350 ;
        RECT 21.520 97.180 24.270 97.350 ;
        RECT 20.500 97.160 20.690 97.180 ;
        RECT 20.160 97.040 20.330 97.080 ;
        RECT 23.450 97.000 23.790 97.180 ;
        RECT 17.940 96.710 18.540 96.880 ;
        RECT 19.000 96.720 19.330 96.890 ;
        RECT 17.940 96.560 18.390 96.710 ;
        RECT 20.230 96.440 20.400 96.860 ;
        RECT 21.040 96.730 21.280 96.770 ;
        RECT 23.820 96.730 23.990 96.740 ;
        RECT 20.710 96.560 21.280 96.730 ;
        RECT 21.520 96.560 22.860 96.730 ;
        RECT 23.310 96.560 24.270 96.730 ;
        RECT 21.040 96.530 21.280 96.560 ;
        RECT 24.800 96.490 24.970 97.420 ;
        RECT 25.200 96.440 25.370 97.330 ;
        RECT 28.100 97.000 28.320 97.590 ;
        RECT 28.100 96.970 28.310 97.000 ;
        RECT 28.840 96.990 29.040 97.590 ;
        RECT 30.850 97.510 31.020 98.040 ;
        RECT 34.790 97.520 34.960 98.050 ;
        RECT 40.580 97.520 40.750 98.050 ;
        RECT 44.520 97.510 44.690 98.040 ;
        RECT 29.850 97.490 30.170 97.500 ;
        RECT 29.590 97.320 30.170 97.490 ;
        RECT 29.840 97.280 30.170 97.320 ;
        RECT 29.850 97.240 30.170 97.280 ;
        RECT 45.370 97.490 45.690 97.500 ;
        RECT 45.370 97.320 45.950 97.490 ;
        RECT 45.370 97.280 45.700 97.320 ;
        RECT 45.370 97.240 45.690 97.280 ;
        RECT 46.500 96.990 46.700 97.590 ;
        RECT 47.220 97.000 47.440 97.590 ;
        RECT 28.110 96.620 28.310 96.970 ;
        RECT 47.230 96.970 47.440 97.000 ;
        RECT 29.850 96.920 30.170 96.950 ;
        RECT 29.840 96.870 30.170 96.920 ;
        RECT 29.590 96.700 30.170 96.870 ;
        RECT 45.370 96.920 45.690 96.950 ;
        RECT 45.370 96.870 45.700 96.920 ;
        RECT 29.850 96.690 30.170 96.700 ;
        RECT 28.480 96.160 28.920 96.330 ;
        RECT 11.190 95.970 11.360 96.020 ;
        RECT 11.160 95.750 11.380 95.970 ;
        RECT 11.190 95.690 11.360 95.750 ;
        RECT 11.710 95.610 12.040 95.790 ;
        RECT 14.850 95.780 15.020 95.830 ;
        RECT 12.290 95.610 14.450 95.780 ;
        RECT 14.690 95.610 15.020 95.780 ;
        RECT 15.310 95.640 15.520 95.970 ;
        RECT 11.740 95.170 12.010 95.610 ;
        RECT 13.220 95.350 13.550 95.610 ;
        RECT 14.760 95.470 15.020 95.610 ;
        RECT 15.760 95.470 15.940 95.910 ;
        RECT 17.360 95.810 17.750 95.860 ;
        RECT 16.490 95.750 17.750 95.810 ;
        RECT 16.490 95.640 17.830 95.750 ;
        RECT 17.360 95.580 17.830 95.640 ;
        RECT 18.300 95.600 19.260 95.770 ;
        RECT 17.360 95.570 17.740 95.580 ;
        RECT 11.780 95.160 12.010 95.170 ;
        RECT 14.760 95.300 15.940 95.470 ;
        RECT 14.760 95.160 15.020 95.300 ;
        RECT 11.780 94.990 12.540 95.160 ;
        RECT 12.790 94.990 13.960 95.160 ;
        RECT 14.200 95.130 15.020 95.160 ;
        RECT 14.200 94.990 15.310 95.130 ;
        RECT 13.190 94.890 13.540 94.990 ;
        RECT 14.850 94.960 15.310 94.990 ;
        RECT 15.760 95.120 16.950 95.130 ;
        RECT 15.760 94.960 17.240 95.120 ;
        RECT 15.800 94.940 17.240 94.960 ;
        RECT 16.780 94.900 17.240 94.940 ;
        RECT 16.950 94.880 17.240 94.900 ;
        RECT 17.570 94.810 17.740 95.570 ;
        RECT 19.080 95.140 19.260 95.600 ;
        RECT 20.230 95.550 20.400 95.970 ;
        RECT 21.040 95.850 21.280 95.880 ;
        RECT 20.710 95.680 21.280 95.850 ;
        RECT 21.520 95.680 22.860 95.850 ;
        RECT 23.310 95.680 24.270 95.850 ;
        RECT 21.040 95.640 21.280 95.680 ;
        RECT 23.820 95.670 23.990 95.680 ;
        RECT 20.160 95.330 20.330 95.370 ;
        RECT 20.100 95.160 20.330 95.330 ;
        RECT 17.940 94.960 18.540 95.130 ;
        RECT 19.000 94.970 19.330 95.140 ;
        RECT 17.940 94.810 18.390 94.960 ;
        RECT 20.160 94.810 20.330 95.160 ;
        RECT 20.500 95.230 20.690 95.250 ;
        RECT 23.450 95.230 23.790 95.410 ;
        RECT 20.500 95.060 21.060 95.230 ;
        RECT 21.520 95.060 24.270 95.230 ;
        RECT 20.500 95.020 20.690 95.060 ;
        RECT 24.800 94.990 24.970 95.920 ;
        RECT 25.200 95.080 25.370 95.970 ;
        RECT 28.110 95.520 28.310 95.870 ;
        RECT 29.850 95.790 30.170 95.800 ;
        RECT 29.590 95.620 30.170 95.790 ;
        RECT 30.850 95.670 31.020 96.680 ;
        RECT 32.780 95.950 33.330 96.380 ;
        RECT 34.780 95.810 34.950 96.820 ;
        RECT 36.810 96.020 37.360 96.450 ;
        RECT 38.180 96.020 38.730 96.450 ;
        RECT 40.590 95.810 40.760 96.820 ;
        RECT 45.370 96.700 45.950 96.870 ;
        RECT 45.370 96.690 45.690 96.700 ;
        RECT 42.210 95.950 42.760 96.380 ;
        RECT 44.520 95.670 44.690 96.680 ;
        RECT 47.230 96.620 47.430 96.970 ;
        RECT 46.620 96.160 47.060 96.330 ;
        RECT 45.370 95.790 45.690 95.800 ;
        RECT 29.840 95.570 30.170 95.620 ;
        RECT 29.850 95.540 30.170 95.570 ;
        RECT 45.370 95.620 45.950 95.790 ;
        RECT 45.370 95.570 45.700 95.620 ;
        RECT 45.370 95.540 45.690 95.570 ;
        RECT 28.100 95.490 28.310 95.520 ;
        RECT 47.230 95.520 47.430 95.870 ;
        RECT 28.100 94.900 28.320 95.490 ;
        RECT 28.840 94.900 29.040 95.500 ;
        RECT 29.850 95.210 30.170 95.250 ;
        RECT 29.840 95.170 30.170 95.210 ;
        RECT 29.590 95.000 30.170 95.170 ;
        RECT 29.850 94.990 30.170 95.000 ;
        RECT 45.370 95.210 45.690 95.250 ;
        RECT 45.370 95.170 45.700 95.210 ;
        RECT 45.370 95.000 45.950 95.170 ;
        RECT 45.370 94.990 45.690 95.000 ;
        RECT 46.500 94.900 46.700 95.500 ;
        RECT 47.230 95.490 47.440 95.520 ;
        RECT 47.220 94.900 47.440 95.490 ;
        RECT 11.190 94.220 11.360 94.270 ;
        RECT 11.160 94.000 11.380 94.220 ;
        RECT 11.190 93.940 11.360 94.000 ;
        RECT 11.710 93.860 12.040 94.040 ;
        RECT 14.850 94.030 15.020 94.080 ;
        RECT 12.290 93.860 14.450 94.030 ;
        RECT 14.690 93.860 15.020 94.030 ;
        RECT 15.310 93.890 15.520 94.220 ;
        RECT 11.740 93.420 12.010 93.860 ;
        RECT 13.220 93.600 13.550 93.860 ;
        RECT 14.760 93.720 15.020 93.860 ;
        RECT 15.760 93.720 15.940 94.160 ;
        RECT 17.360 94.060 17.750 94.110 ;
        RECT 16.490 94.000 17.750 94.060 ;
        RECT 20.160 94.050 20.330 94.400 ;
        RECT 16.490 93.890 17.830 94.000 ;
        RECT 17.360 93.830 17.830 93.890 ;
        RECT 18.300 93.850 19.260 94.020 ;
        RECT 20.100 93.880 20.330 94.050 ;
        RECT 20.500 94.150 20.690 94.190 ;
        RECT 20.500 93.980 21.060 94.150 ;
        RECT 21.520 93.980 24.270 94.150 ;
        RECT 20.500 93.960 20.690 93.980 ;
        RECT 17.360 93.820 17.740 93.830 ;
        RECT 11.780 93.410 12.010 93.420 ;
        RECT 14.760 93.550 15.940 93.720 ;
        RECT 14.760 93.410 15.020 93.550 ;
        RECT 11.780 93.240 12.540 93.410 ;
        RECT 12.790 93.240 13.960 93.410 ;
        RECT 14.200 93.380 15.020 93.410 ;
        RECT 14.200 93.240 15.310 93.380 ;
        RECT 13.190 93.140 13.540 93.240 ;
        RECT 14.850 93.210 15.310 93.240 ;
        RECT 15.760 93.370 16.950 93.380 ;
        RECT 15.760 93.210 17.240 93.370 ;
        RECT 15.800 93.190 17.240 93.210 ;
        RECT 16.780 93.150 17.240 93.190 ;
        RECT 16.950 93.130 17.240 93.150 ;
        RECT 17.570 93.060 17.740 93.820 ;
        RECT 19.080 93.390 19.260 93.850 ;
        RECT 20.160 93.840 20.330 93.880 ;
        RECT 23.450 93.800 23.790 93.980 ;
        RECT 17.940 93.210 18.540 93.380 ;
        RECT 19.000 93.220 19.330 93.390 ;
        RECT 20.230 93.240 20.400 93.660 ;
        RECT 21.040 93.530 21.280 93.570 ;
        RECT 23.820 93.530 23.990 93.540 ;
        RECT 20.710 93.360 21.280 93.530 ;
        RECT 21.520 93.360 22.860 93.530 ;
        RECT 23.310 93.360 24.270 93.530 ;
        RECT 21.040 93.330 21.280 93.360 ;
        RECT 24.800 93.290 24.970 94.220 ;
        RECT 25.200 93.240 25.370 94.130 ;
        RECT 28.100 93.770 28.320 94.360 ;
        RECT 28.100 93.740 28.310 93.770 ;
        RECT 28.840 93.760 29.040 94.360 ;
        RECT 29.850 94.260 30.170 94.270 ;
        RECT 29.590 94.090 30.170 94.260 ;
        RECT 29.840 94.050 30.170 94.090 ;
        RECT 29.850 94.010 30.170 94.050 ;
        RECT 45.370 94.260 45.690 94.270 ;
        RECT 45.370 94.090 45.950 94.260 ;
        RECT 45.370 94.050 45.700 94.090 ;
        RECT 45.370 94.010 45.690 94.050 ;
        RECT 46.500 93.760 46.700 94.360 ;
        RECT 47.220 93.770 47.440 94.360 ;
        RECT 28.110 93.390 28.310 93.740 ;
        RECT 47.230 93.740 47.440 93.770 ;
        RECT 29.850 93.690 30.170 93.720 ;
        RECT 29.840 93.640 30.170 93.690 ;
        RECT 29.590 93.470 30.170 93.640 ;
        RECT 29.850 93.460 30.170 93.470 ;
        RECT 45.370 93.690 45.690 93.720 ;
        RECT 45.370 93.640 45.700 93.690 ;
        RECT 45.370 93.470 45.950 93.640 ;
        RECT 45.370 93.460 45.690 93.470 ;
        RECT 47.230 93.390 47.430 93.740 ;
        RECT 17.940 93.060 18.390 93.210 ;
        RECT -12.140 90.110 -11.970 90.600 ;
        RECT -12.290 90.080 -11.970 90.110 ;
        RECT -11.590 90.110 -11.420 90.600 ;
        RECT -10.950 90.550 -10.780 90.600 ;
        RECT -10.400 90.550 -10.230 90.600 ;
        RECT -11.070 90.520 -10.750 90.550 ;
        RECT -10.420 90.520 -10.100 90.550 ;
        RECT -11.070 90.330 -10.740 90.520 ;
        RECT -10.420 90.330 -10.090 90.520 ;
        RECT 11.150 90.410 11.320 90.460 ;
        RECT -11.070 90.290 -10.750 90.330 ;
        RECT -10.420 90.290 -10.100 90.330 ;
        RECT -11.590 90.080 -11.270 90.110 ;
        RECT -12.290 89.890 -11.960 90.080 ;
        RECT -11.590 89.890 -11.260 90.080 ;
        RECT -12.290 89.850 -11.970 89.890 ;
        RECT -12.680 88.390 -12.510 88.410 ;
        RECT -12.700 87.960 -12.490 88.390 ;
        RECT -12.140 88.200 -11.970 89.850 ;
        RECT -11.590 89.850 -11.270 89.890 ;
        RECT -11.590 88.200 -11.420 89.850 ;
        RECT -10.950 88.200 -10.780 90.290 ;
        RECT -10.400 88.200 -10.230 90.290 ;
        RECT 11.120 90.190 11.340 90.410 ;
        RECT 11.150 90.130 11.320 90.190 ;
        RECT 11.670 90.050 12.000 90.230 ;
        RECT 14.810 90.220 14.980 90.270 ;
        RECT 12.250 90.050 14.410 90.220 ;
        RECT 14.650 90.050 14.980 90.220 ;
        RECT 15.270 90.080 15.480 90.410 ;
        RECT -9.850 88.840 -9.680 89.690 ;
        RECT 11.700 89.610 11.970 90.050 ;
        RECT 13.180 89.790 13.510 90.050 ;
        RECT 14.720 89.910 14.980 90.050 ;
        RECT 15.720 89.910 15.900 90.350 ;
        RECT 17.320 90.250 17.710 90.300 ;
        RECT 16.450 90.190 17.710 90.250 ;
        RECT 16.450 90.080 17.790 90.190 ;
        RECT 17.320 90.020 17.790 90.080 ;
        RECT 18.260 90.040 19.220 90.210 ;
        RECT 17.320 90.010 17.700 90.020 ;
        RECT 11.740 89.600 11.970 89.610 ;
        RECT 14.720 89.740 15.900 89.910 ;
        RECT 14.720 89.600 14.980 89.740 ;
        RECT 11.740 89.430 12.500 89.600 ;
        RECT 12.750 89.430 13.920 89.600 ;
        RECT 14.160 89.570 14.980 89.600 ;
        RECT 14.160 89.430 15.270 89.570 ;
        RECT 13.150 89.330 13.500 89.430 ;
        RECT 14.810 89.400 15.270 89.430 ;
        RECT 15.720 89.560 16.910 89.570 ;
        RECT 15.720 89.400 17.200 89.560 ;
        RECT 15.760 89.380 17.200 89.400 ;
        RECT 16.740 89.340 17.200 89.380 ;
        RECT 16.910 89.320 17.200 89.340 ;
        RECT 17.530 89.250 17.700 90.010 ;
        RECT 19.040 89.580 19.220 90.040 ;
        RECT 17.900 89.400 18.500 89.570 ;
        RECT 18.960 89.410 19.290 89.580 ;
        RECT 20.260 89.480 20.430 89.900 ;
        RECT 21.070 89.780 21.310 89.810 ;
        RECT 20.740 89.610 21.310 89.780 ;
        RECT 21.550 89.610 22.890 89.780 ;
        RECT 23.340 89.610 24.300 89.780 ;
        RECT 21.070 89.570 21.310 89.610 ;
        RECT 23.850 89.600 24.020 89.610 ;
        RECT 17.900 89.250 18.350 89.400 ;
        RECT 20.190 89.260 20.360 89.300 ;
        RECT 20.130 89.090 20.360 89.260 ;
        RECT 20.190 88.740 20.360 89.090 ;
        RECT 20.530 89.160 20.720 89.180 ;
        RECT 23.480 89.160 23.820 89.340 ;
        RECT 20.530 88.990 21.090 89.160 ;
        RECT 21.550 88.990 24.300 89.160 ;
        RECT 20.530 88.950 20.720 88.990 ;
        RECT 24.830 88.920 25.000 89.850 ;
        RECT 25.230 89.010 25.400 89.900 ;
        RECT 28.140 89.430 28.340 89.780 ;
        RECT 29.880 89.700 30.200 89.710 ;
        RECT 29.620 89.530 30.200 89.700 ;
        RECT 29.870 89.480 30.200 89.530 ;
        RECT 29.880 89.450 30.200 89.480 ;
        RECT 28.130 89.400 28.340 89.430 ;
        RECT 28.130 88.810 28.350 89.400 ;
        RECT 28.870 88.810 29.070 89.410 ;
        RECT 38.590 89.380 38.910 89.410 ;
        RECT 38.590 89.210 40.380 89.380 ;
        RECT 38.590 89.190 38.920 89.210 ;
        RECT 29.880 89.120 30.200 89.160 ;
        RECT 38.590 89.150 38.910 89.190 ;
        RECT 29.870 89.080 30.200 89.120 ;
        RECT 29.620 88.910 30.200 89.080 ;
        RECT 40.210 88.980 40.380 89.210 ;
        RECT 29.880 88.900 30.200 88.910 ;
        RECT 39.060 88.730 39.400 88.980 ;
        RECT 39.570 88.810 39.900 88.980 ;
        RECT 40.120 88.810 40.460 88.980 ;
        RECT 11.150 88.660 11.320 88.710 ;
        RECT 11.120 88.440 11.340 88.660 ;
        RECT 11.150 88.380 11.320 88.440 ;
        RECT 11.670 88.300 12.000 88.480 ;
        RECT 14.810 88.470 14.980 88.520 ;
        RECT 12.250 88.300 14.410 88.470 ;
        RECT 14.650 88.300 14.980 88.470 ;
        RECT 15.270 88.330 15.480 88.660 ;
        RECT -9.960 88.210 -9.530 88.230 ;
        RECT -9.960 88.040 -9.510 88.210 ;
        RECT -9.960 88.020 -9.530 88.040 ;
        RECT 11.700 87.860 11.970 88.300 ;
        RECT 13.180 88.040 13.510 88.300 ;
        RECT 14.720 88.160 14.980 88.300 ;
        RECT 15.720 88.160 15.900 88.600 ;
        RECT 17.320 88.500 17.710 88.550 ;
        RECT 16.450 88.440 17.710 88.500 ;
        RECT 16.450 88.330 17.790 88.440 ;
        RECT 17.320 88.270 17.790 88.330 ;
        RECT 18.260 88.290 19.220 88.460 ;
        RECT 17.320 88.260 17.700 88.270 ;
        RECT -150.440 87.340 -142.910 87.850 ;
        RECT 11.740 87.850 11.970 87.860 ;
        RECT 14.720 87.990 15.900 88.160 ;
        RECT 14.720 87.850 14.980 87.990 ;
        RECT -152.140 81.320 -150.680 81.360 ;
        RECT -152.140 81.150 -150.670 81.320 ;
        RECT -152.140 81.110 -150.680 81.150 ;
        RECT -150.440 74.730 -149.930 87.340 ;
        RECT -149.570 86.550 -143.590 86.780 ;
        RECT -149.480 75.490 -143.830 86.550 ;
        RECT -143.420 76.980 -142.910 87.340 ;
        RECT -12.690 87.320 -12.480 87.750 ;
        RECT -9.950 87.670 -9.520 87.690 ;
        RECT 11.740 87.680 12.500 87.850 ;
        RECT 12.750 87.680 13.920 87.850 ;
        RECT 14.160 87.820 14.980 87.850 ;
        RECT 14.160 87.680 15.270 87.820 ;
        RECT -12.670 87.300 -12.500 87.320 ;
        RECT -12.130 86.230 -11.960 87.550 ;
        RECT -12.260 86.200 -11.940 86.230 ;
        RECT -11.580 86.220 -11.410 87.560 ;
        RECT -12.260 86.010 -11.930 86.200 ;
        RECT -11.580 86.190 -11.250 86.220 ;
        RECT -12.260 85.970 -11.940 86.010 ;
        RECT -11.580 86.000 -11.240 86.190 ;
        RECT -12.130 85.060 -11.960 85.970 ;
        RECT -11.580 85.960 -11.250 86.000 ;
        RECT -11.580 85.060 -11.410 85.960 ;
        RECT -10.950 85.450 -10.780 87.550 ;
        RECT -11.090 85.420 -10.770 85.450 ;
        RECT -11.090 85.230 -10.760 85.420 ;
        RECT -10.400 85.390 -10.230 87.560 ;
        RECT -9.950 87.500 -9.500 87.670 ;
        RECT 13.150 87.580 13.500 87.680 ;
        RECT 14.810 87.650 15.270 87.680 ;
        RECT 15.720 87.810 16.910 87.820 ;
        RECT 15.720 87.650 17.200 87.810 ;
        RECT 15.760 87.630 17.200 87.650 ;
        RECT 16.740 87.590 17.200 87.630 ;
        RECT 16.910 87.570 17.200 87.590 ;
        RECT 17.530 87.500 17.700 88.260 ;
        RECT 19.040 87.830 19.220 88.290 ;
        RECT 20.190 87.980 20.360 88.330 ;
        RECT 17.900 87.650 18.500 87.820 ;
        RECT 18.960 87.660 19.290 87.830 ;
        RECT 20.130 87.810 20.360 87.980 ;
        RECT 20.530 88.080 20.720 88.120 ;
        RECT 20.530 87.910 21.090 88.080 ;
        RECT 21.550 87.910 24.300 88.080 ;
        RECT 20.530 87.890 20.720 87.910 ;
        RECT 20.190 87.770 20.360 87.810 ;
        RECT 23.480 87.730 23.820 87.910 ;
        RECT 17.900 87.500 18.350 87.650 ;
        RECT -9.950 87.480 -9.520 87.500 ;
        RECT 20.260 87.170 20.430 87.590 ;
        RECT 21.070 87.460 21.310 87.500 ;
        RECT 23.850 87.460 24.020 87.470 ;
        RECT 20.740 87.290 21.310 87.460 ;
        RECT 21.550 87.290 22.890 87.460 ;
        RECT 23.340 87.290 24.300 87.460 ;
        RECT 21.070 87.260 21.310 87.290 ;
        RECT 24.830 87.220 25.000 88.150 ;
        RECT 25.230 87.170 25.400 88.060 ;
        RECT 28.130 87.690 28.350 88.280 ;
        RECT 28.130 87.660 28.340 87.690 ;
        RECT 28.870 87.680 29.070 88.280 ;
        RECT 29.880 88.180 30.200 88.190 ;
        RECT 29.620 88.010 30.200 88.180 ;
        RECT 31.010 88.120 31.180 88.650 ;
        RECT 35.030 88.150 35.200 88.680 ;
        RECT 38.740 88.470 39.400 88.730 ;
        RECT 39.650 88.640 39.820 88.810 ;
        RECT 40.210 88.640 40.380 88.810 ;
        RECT 39.570 88.470 39.900 88.640 ;
        RECT 40.120 88.470 40.460 88.640 ;
        RECT 39.650 88.240 39.900 88.470 ;
        RECT 40.780 88.390 41.290 89.060 ;
        RECT 29.870 87.970 30.200 88.010 ;
        RECT 29.880 87.930 30.200 87.970 ;
        RECT 39.650 88.070 40.320 88.240 ;
        RECT 39.650 87.840 39.900 88.070 ;
        RECT 28.140 87.310 28.340 87.660 ;
        RECT 29.880 87.610 30.200 87.640 ;
        RECT 29.870 87.560 30.200 87.610 ;
        RECT 38.740 87.580 39.400 87.840 ;
        RECT 39.570 87.670 39.900 87.840 ;
        RECT 40.120 87.670 40.460 87.840 ;
        RECT 29.620 87.390 30.200 87.560 ;
        RECT 29.880 87.380 30.200 87.390 ;
        RECT -9.860 86.290 -9.690 86.960 ;
        RECT 11.150 86.910 11.320 86.960 ;
        RECT 11.120 86.690 11.340 86.910 ;
        RECT 11.150 86.630 11.320 86.690 ;
        RECT 11.670 86.550 12.000 86.730 ;
        RECT 14.810 86.720 14.980 86.770 ;
        RECT 12.250 86.550 14.410 86.720 ;
        RECT 14.650 86.550 14.980 86.720 ;
        RECT 15.270 86.580 15.480 86.910 ;
        RECT 28.510 86.850 28.950 87.020 ;
        RECT 11.700 86.110 11.970 86.550 ;
        RECT 13.180 86.290 13.510 86.550 ;
        RECT 14.720 86.410 14.980 86.550 ;
        RECT 15.720 86.410 15.900 86.850 ;
        RECT 17.320 86.750 17.710 86.800 ;
        RECT 16.450 86.690 17.710 86.750 ;
        RECT 16.450 86.580 17.790 86.690 ;
        RECT 17.320 86.520 17.790 86.580 ;
        RECT 18.260 86.540 19.220 86.710 ;
        RECT 17.320 86.510 17.700 86.520 ;
        RECT 11.740 86.100 11.970 86.110 ;
        RECT 14.720 86.240 15.900 86.410 ;
        RECT 14.720 86.100 14.980 86.240 ;
        RECT 11.740 85.930 12.500 86.100 ;
        RECT 12.750 85.930 13.920 86.100 ;
        RECT 14.160 86.070 14.980 86.100 ;
        RECT 14.160 85.930 15.270 86.070 ;
        RECT 13.150 85.830 13.500 85.930 ;
        RECT 14.810 85.900 15.270 85.930 ;
        RECT 15.720 86.060 16.910 86.070 ;
        RECT 15.720 85.900 17.200 86.060 ;
        RECT 15.760 85.880 17.200 85.900 ;
        RECT 16.740 85.840 17.200 85.880 ;
        RECT 16.910 85.820 17.200 85.840 ;
        RECT 17.530 85.750 17.700 86.510 ;
        RECT 19.040 86.080 19.220 86.540 ;
        RECT 20.260 86.280 20.430 86.700 ;
        RECT 21.070 86.580 21.310 86.610 ;
        RECT 20.740 86.410 21.310 86.580 ;
        RECT 21.550 86.410 22.890 86.580 ;
        RECT 23.340 86.410 24.300 86.580 ;
        RECT 21.070 86.370 21.310 86.410 ;
        RECT 23.850 86.400 24.020 86.410 ;
        RECT 17.900 85.900 18.500 86.070 ;
        RECT 18.960 85.910 19.290 86.080 ;
        RECT 20.190 86.060 20.360 86.100 ;
        RECT 17.900 85.750 18.350 85.900 ;
        RECT 20.130 85.890 20.360 86.060 ;
        RECT 20.190 85.540 20.360 85.890 ;
        RECT 20.530 85.960 20.720 85.980 ;
        RECT 23.480 85.960 23.820 86.140 ;
        RECT 20.530 85.790 21.090 85.960 ;
        RECT 21.550 85.790 24.300 85.960 ;
        RECT 20.530 85.750 20.720 85.790 ;
        RECT 24.830 85.720 25.000 86.650 ;
        RECT 25.230 85.810 25.400 86.700 ;
        RECT 28.140 86.190 28.340 86.540 ;
        RECT 29.880 86.460 30.200 86.470 ;
        RECT 29.620 86.290 30.200 86.460 ;
        RECT 29.870 86.240 30.200 86.290 ;
        RECT 31.000 86.260 31.170 87.450 ;
        RECT 32.810 86.580 33.360 87.010 ;
        RECT 29.880 86.210 30.200 86.240 ;
        RECT 35.020 86.220 35.190 87.390 ;
        RECT 39.060 87.330 39.400 87.580 ;
        RECT 39.650 87.500 39.820 87.670 ;
        RECT 40.210 87.500 40.380 87.670 ;
        RECT 39.570 87.330 39.900 87.500 ;
        RECT 40.120 87.330 40.460 87.500 ;
        RECT 38.590 87.120 38.910 87.160 ;
        RECT 38.590 87.100 38.920 87.120 ;
        RECT 40.210 87.100 40.380 87.330 ;
        RECT 40.780 87.250 41.290 87.920 ;
        RECT 36.840 86.650 37.390 87.080 ;
        RECT 38.590 86.930 40.380 87.100 ;
        RECT 206.500 87.130 207.010 100.030 ;
        RECT 207.410 99.140 210.870 99.580 ;
        RECT 207.410 99.040 212.800 99.140 ;
        RECT 207.520 98.970 212.800 99.040 ;
        RECT 207.520 88.060 207.690 98.970 ;
        RECT 208.070 98.560 212.300 98.580 ;
        RECT 207.990 88.450 212.320 98.560 ;
        RECT 212.090 88.400 212.260 88.450 ;
        RECT 212.630 88.060 212.800 98.970 ;
        RECT 207.520 87.890 212.800 88.060 ;
        RECT 207.520 87.880 207.760 87.890 ;
        RECT 213.520 87.130 214.030 100.040 ;
        RECT 38.590 86.900 38.910 86.930 ;
        RECT 38.590 86.610 38.910 86.640 ;
        RECT 206.500 86.620 214.030 87.130 ;
        RECT 214.240 87.070 215.720 87.320 ;
        RECT 38.590 86.440 40.380 86.610 ;
        RECT 38.590 86.420 38.920 86.440 ;
        RECT 38.590 86.380 38.910 86.420 ;
        RECT 40.210 86.210 40.380 86.440 ;
        RECT 28.130 86.160 28.340 86.190 ;
        RECT 28.130 85.570 28.350 86.160 ;
        RECT 28.870 85.570 29.070 86.170 ;
        RECT 39.060 85.960 39.400 86.210 ;
        RECT 39.570 86.040 39.900 86.210 ;
        RECT 40.120 86.040 40.460 86.210 ;
        RECT 29.880 85.880 30.200 85.920 ;
        RECT 29.870 85.840 30.200 85.880 ;
        RECT 29.620 85.670 30.200 85.840 ;
        RECT 38.740 85.700 39.400 85.960 ;
        RECT 39.650 85.870 39.820 86.040 ;
        RECT 40.210 85.870 40.380 86.040 ;
        RECT 39.570 85.700 39.900 85.870 ;
        RECT 40.120 85.700 40.460 85.870 ;
        RECT 29.880 85.660 30.200 85.670 ;
        RECT 39.650 85.470 39.900 85.700 ;
        RECT 40.780 85.620 41.290 86.290 ;
        RECT -10.400 85.360 -10.060 85.390 ;
        RECT -11.090 85.190 -10.770 85.230 ;
        RECT -10.950 85.060 -10.780 85.190 ;
        RECT -10.400 85.170 -10.050 85.360 ;
        RECT 39.650 85.300 40.320 85.470 ;
        RECT -10.400 85.130 -10.060 85.170 ;
        RECT 11.150 85.160 11.320 85.210 ;
        RECT -10.400 85.060 -10.230 85.130 ;
        RECT 11.120 84.940 11.340 85.160 ;
        RECT 11.150 84.880 11.320 84.940 ;
        RECT 11.670 84.800 12.000 84.980 ;
        RECT 14.810 84.970 14.980 85.020 ;
        RECT 12.250 84.800 14.410 84.970 ;
        RECT 14.650 84.800 14.980 84.970 ;
        RECT 15.270 84.830 15.480 85.160 ;
        RECT 11.700 84.360 11.970 84.800 ;
        RECT 13.180 84.540 13.510 84.800 ;
        RECT 14.720 84.660 14.980 84.800 ;
        RECT 15.720 84.660 15.900 85.100 ;
        RECT 17.320 85.000 17.710 85.050 ;
        RECT 16.450 84.940 17.710 85.000 ;
        RECT 16.450 84.830 17.790 84.940 ;
        RECT 17.320 84.770 17.790 84.830 ;
        RECT 18.260 84.790 19.220 84.960 ;
        RECT 17.320 84.760 17.700 84.770 ;
        RECT 11.740 84.350 11.970 84.360 ;
        RECT 14.720 84.490 15.900 84.660 ;
        RECT 14.720 84.350 14.980 84.490 ;
        RECT 11.740 84.180 12.500 84.350 ;
        RECT 12.750 84.180 13.920 84.350 ;
        RECT 14.160 84.320 14.980 84.350 ;
        RECT 14.160 84.180 15.270 84.320 ;
        RECT 13.150 84.080 13.500 84.180 ;
        RECT 14.810 84.150 15.270 84.180 ;
        RECT 15.720 84.310 16.910 84.320 ;
        RECT 15.720 84.150 17.200 84.310 ;
        RECT 15.760 84.130 17.200 84.150 ;
        RECT 16.740 84.090 17.200 84.130 ;
        RECT 16.910 84.070 17.200 84.090 ;
        RECT 17.530 84.000 17.700 84.760 ;
        RECT 19.040 84.330 19.220 84.790 ;
        RECT 20.190 84.780 20.360 85.130 ;
        RECT 39.650 85.070 39.900 85.300 ;
        RECT 27.150 84.970 27.470 85.010 ;
        RECT 20.130 84.610 20.360 84.780 ;
        RECT 20.530 84.880 20.720 84.920 ;
        RECT 20.530 84.710 21.090 84.880 ;
        RECT 21.550 84.710 24.300 84.880 ;
        RECT 20.530 84.690 20.720 84.710 ;
        RECT 20.190 84.570 20.360 84.610 ;
        RECT 23.480 84.530 23.820 84.710 ;
        RECT 17.900 84.150 18.500 84.320 ;
        RECT 18.960 84.160 19.290 84.330 ;
        RECT 17.900 84.000 18.350 84.150 ;
        RECT 20.260 83.970 20.430 84.390 ;
        RECT 21.070 84.260 21.310 84.300 ;
        RECT 23.850 84.260 24.020 84.270 ;
        RECT 20.740 84.090 21.310 84.260 ;
        RECT 21.550 84.090 22.890 84.260 ;
        RECT 23.340 84.090 24.300 84.260 ;
        RECT 21.070 84.060 21.310 84.090 ;
        RECT 24.830 84.020 25.000 84.950 ;
        RECT 25.230 83.970 25.400 84.860 ;
        RECT 27.150 84.780 27.480 84.970 ;
        RECT 27.150 84.750 27.470 84.780 ;
        RECT 27.200 84.050 27.380 84.750 ;
        RECT 28.130 84.440 28.350 85.030 ;
        RECT 28.130 84.410 28.340 84.440 ;
        RECT 28.870 84.430 29.070 85.030 ;
        RECT 29.880 84.930 30.200 84.940 ;
        RECT 29.620 84.760 30.200 84.930 ;
        RECT 38.740 84.810 39.400 85.070 ;
        RECT 39.570 84.900 39.900 85.070 ;
        RECT 40.120 84.900 40.460 85.070 ;
        RECT 29.870 84.720 30.200 84.760 ;
        RECT 29.880 84.680 30.200 84.720 ;
        RECT 39.060 84.560 39.400 84.810 ;
        RECT 39.650 84.730 39.820 84.900 ;
        RECT 40.210 84.730 40.380 84.900 ;
        RECT 39.570 84.560 39.900 84.730 ;
        RECT 40.120 84.560 40.460 84.730 ;
        RECT 28.140 84.060 28.340 84.410 ;
        RECT 29.880 84.360 30.200 84.390 ;
        RECT 29.870 84.310 30.200 84.360 ;
        RECT 29.620 84.140 30.200 84.310 ;
        RECT 29.880 84.130 30.200 84.140 ;
        RECT 38.590 84.350 38.910 84.390 ;
        RECT 38.590 84.330 38.920 84.350 ;
        RECT 40.210 84.330 40.380 84.560 ;
        RECT 40.780 84.480 41.290 85.150 ;
        RECT 38.590 84.160 40.380 84.330 ;
        RECT 38.590 84.130 38.910 84.160 ;
        RECT 27.200 84.010 27.520 84.050 ;
        RECT 27.200 83.820 27.530 84.010 ;
        RECT 27.200 83.790 27.520 83.820 ;
        RECT 19.940 82.050 20.110 82.140 ;
        RECT 19.860 82.010 20.180 82.050 ;
        RECT 19.860 81.820 20.190 82.010 ;
        RECT 19.860 81.790 20.180 81.820 ;
        RECT -14.330 79.930 -14.160 80.000 ;
        RECT -14.400 79.900 -14.080 79.930 ;
        RECT -14.410 79.710 -14.080 79.900 ;
        RECT -14.400 79.670 -14.080 79.710 ;
        RECT -14.330 77.160 -14.160 79.670 ;
        RECT -13.780 79.260 -13.610 80.000 ;
        RECT -13.230 79.940 -13.060 80.000 ;
        RECT -13.300 79.910 -12.980 79.940 ;
        RECT -13.310 79.720 -12.980 79.910 ;
        RECT -13.300 79.680 -12.980 79.720 ;
        RECT -13.850 79.230 -13.530 79.260 ;
        RECT -13.860 79.040 -13.530 79.230 ;
        RECT -13.850 79.000 -13.530 79.040 ;
        RECT -13.780 77.890 -13.610 79.000 ;
        RECT -13.850 77.860 -13.530 77.890 ;
        RECT -13.860 77.670 -13.530 77.860 ;
        RECT -13.850 77.630 -13.530 77.670 ;
        RECT -14.400 77.130 -14.080 77.160 ;
        RECT -143.430 76.960 -142.910 76.980 ;
        RECT -149.480 75.480 -143.770 75.490 ;
        RECT -149.560 75.310 -143.770 75.480 ;
        RECT -149.470 75.300 -143.770 75.310 ;
        RECT -144.000 75.230 -143.830 75.300 ;
        RECT -143.430 75.180 -142.900 76.960 ;
        RECT -14.410 76.940 -14.080 77.130 ;
        RECT -14.400 76.900 -14.080 76.940 ;
        RECT -14.330 75.820 -14.160 76.900 ;
        RECT -14.410 75.790 -14.090 75.820 ;
        RECT -14.420 75.600 -14.090 75.790 ;
        RECT -14.410 75.560 -14.090 75.600 ;
        RECT -143.420 75.160 -142.900 75.180 ;
        RECT -150.440 74.440 -148.000 74.730 ;
        RECT -143.420 74.650 -142.910 75.160 ;
        RECT -14.330 74.820 -14.160 75.560 ;
        RECT -13.780 75.120 -13.610 77.630 ;
        RECT -13.230 77.160 -13.060 79.680 ;
        RECT -12.680 79.260 -12.510 80.000 ;
        RECT -12.130 79.940 -11.960 80.000 ;
        RECT -12.210 79.910 -11.890 79.940 ;
        RECT -12.220 79.720 -11.890 79.910 ;
        RECT -12.210 79.680 -11.890 79.720 ;
        RECT -12.750 79.230 -12.430 79.260 ;
        RECT -12.760 79.040 -12.430 79.230 ;
        RECT -12.750 79.000 -12.430 79.040 ;
        RECT -12.680 77.890 -12.510 79.000 ;
        RECT -12.750 77.860 -12.430 77.890 ;
        RECT -12.760 77.670 -12.430 77.860 ;
        RECT -12.750 77.630 -12.430 77.670 ;
        RECT -13.300 77.130 -12.980 77.160 ;
        RECT -13.310 76.940 -12.980 77.130 ;
        RECT -13.300 76.900 -12.980 76.940 ;
        RECT -13.230 75.810 -13.060 76.900 ;
        RECT -13.300 75.780 -12.980 75.810 ;
        RECT -13.310 75.590 -12.980 75.780 ;
        RECT -13.300 75.550 -12.980 75.590 ;
        RECT -13.850 75.090 -13.530 75.120 ;
        RECT -13.860 74.900 -13.530 75.090 ;
        RECT -13.850 74.860 -13.530 74.900 ;
        RECT -13.780 74.820 -13.610 74.860 ;
        RECT -13.230 74.820 -13.060 75.550 ;
        RECT -12.680 75.110 -12.510 77.630 ;
        RECT -12.130 77.160 -11.960 79.680 ;
        RECT -11.580 79.260 -11.410 80.000 ;
        RECT -11.170 79.720 -10.660 80.400 ;
        RECT -3.900 79.900 -3.140 80.320 ;
        RECT -11.170 79.650 -10.650 79.720 ;
        RECT -11.160 79.390 -10.650 79.650 ;
        RECT -11.650 79.230 -11.330 79.260 ;
        RECT -11.660 79.040 -11.330 79.230 ;
        RECT -11.650 79.000 -11.330 79.040 ;
        RECT -11.580 77.890 -11.410 79.000 ;
        RECT -10.870 77.980 -10.700 79.200 ;
        RECT -3.880 79.110 -3.140 79.900 ;
        RECT 19.940 79.270 20.110 81.790 ;
        RECT 20.490 81.370 20.660 82.140 ;
        RECT 21.040 82.050 21.210 82.140 ;
        RECT 20.950 82.010 21.270 82.050 ;
        RECT 20.950 81.820 21.280 82.010 ;
        RECT 20.950 81.790 21.270 81.820 ;
        RECT 20.410 81.330 20.730 81.370 ;
        RECT 20.410 81.140 20.740 81.330 ;
        RECT 20.410 81.110 20.730 81.140 ;
        RECT 20.490 80.000 20.660 81.110 ;
        RECT 20.410 79.960 20.730 80.000 ;
        RECT 20.410 79.770 20.740 79.960 ;
        RECT 20.410 79.740 20.730 79.770 ;
        RECT 19.850 79.230 20.170 79.270 ;
        RECT 19.850 79.040 20.180 79.230 ;
        RECT 19.850 79.010 20.170 79.040 ;
        RECT 19.940 77.900 20.110 79.010 ;
        RECT -11.650 77.860 -11.330 77.890 ;
        RECT -11.660 77.670 -11.330 77.860 ;
        RECT -11.650 77.630 -11.330 77.670 ;
        RECT 19.850 77.860 20.170 77.900 ;
        RECT 19.850 77.670 20.180 77.860 ;
        RECT 19.850 77.640 20.170 77.670 ;
        RECT -12.210 77.130 -11.890 77.160 ;
        RECT -12.220 76.940 -11.890 77.130 ;
        RECT -12.210 76.900 -11.890 76.940 ;
        RECT -12.130 75.790 -11.960 76.900 ;
        RECT -12.210 75.760 -11.890 75.790 ;
        RECT -12.220 75.570 -11.890 75.760 ;
        RECT -12.210 75.530 -11.890 75.570 ;
        RECT -12.750 75.080 -12.430 75.110 ;
        RECT -12.760 74.890 -12.430 75.080 ;
        RECT -12.750 74.850 -12.430 74.890 ;
        RECT -12.680 74.820 -12.510 74.850 ;
        RECT -12.130 74.820 -11.960 75.530 ;
        RECT -11.580 75.110 -11.410 77.630 ;
        RECT 19.170 77.430 19.680 77.510 ;
        RECT 19.170 77.180 19.690 77.430 ;
        RECT 19.180 76.500 19.690 77.180 ;
        RECT 19.940 76.820 20.110 77.640 ;
        RECT 20.490 77.220 20.660 79.740 ;
        RECT 21.040 79.270 21.210 81.790 ;
        RECT 21.590 81.350 21.760 82.140 ;
        RECT 22.140 82.040 22.310 82.140 ;
        RECT 22.050 82.000 22.370 82.040 ;
        RECT 22.050 81.810 22.380 82.000 ;
        RECT 22.050 81.780 22.370 81.810 ;
        RECT 21.500 81.310 21.820 81.350 ;
        RECT 21.500 81.120 21.830 81.310 ;
        RECT 21.500 81.090 21.820 81.120 ;
        RECT 21.590 80.000 21.760 81.090 ;
        RECT 21.500 79.960 21.820 80.000 ;
        RECT 21.500 79.770 21.830 79.960 ;
        RECT 21.500 79.740 21.820 79.770 ;
        RECT 20.950 79.230 21.270 79.270 ;
        RECT 20.950 79.040 21.280 79.230 ;
        RECT 20.950 79.010 21.270 79.040 ;
        RECT 21.040 77.900 21.210 79.010 ;
        RECT 20.950 77.860 21.270 77.900 ;
        RECT 20.950 77.670 21.280 77.860 ;
        RECT 20.950 77.640 21.270 77.670 ;
        RECT 20.410 77.180 20.730 77.220 ;
        RECT 20.410 76.990 20.740 77.180 ;
        RECT 20.410 76.960 20.730 76.990 ;
        RECT 20.490 76.810 20.660 76.960 ;
        RECT 21.040 76.810 21.210 77.640 ;
        RECT 21.590 77.220 21.760 79.740 ;
        RECT 22.140 79.270 22.310 81.780 ;
        RECT 22.690 81.340 22.860 82.140 ;
        RECT 23.230 81.410 23.400 82.170 ;
        RECT 23.840 81.410 24.010 82.170 ;
        RECT 24.380 81.340 24.550 82.140 ;
        RECT 24.930 82.040 25.100 82.140 ;
        RECT 24.870 82.000 25.190 82.040 ;
        RECT 24.860 81.810 25.190 82.000 ;
        RECT 24.870 81.780 25.190 81.810 ;
        RECT 22.610 81.300 22.930 81.340 ;
        RECT 24.310 81.300 24.630 81.340 ;
        RECT 22.610 81.110 22.940 81.300 ;
        RECT 24.300 81.110 24.630 81.300 ;
        RECT 22.610 81.080 22.930 81.110 ;
        RECT 24.310 81.080 24.630 81.110 ;
        RECT 22.690 80.000 22.860 81.080 ;
        RECT 24.380 80.000 24.550 81.080 ;
        RECT 22.600 79.960 22.920 80.000 ;
        RECT 24.320 79.960 24.640 80.000 ;
        RECT 22.600 79.770 22.930 79.960 ;
        RECT 24.310 79.770 24.640 79.960 ;
        RECT 22.600 79.740 22.920 79.770 ;
        RECT 24.320 79.740 24.640 79.770 ;
        RECT 22.050 79.230 22.370 79.270 ;
        RECT 22.050 79.040 22.380 79.230 ;
        RECT 22.050 79.010 22.370 79.040 ;
        RECT 22.140 77.900 22.310 79.010 ;
        RECT 22.050 77.860 22.370 77.900 ;
        RECT 22.050 77.670 22.380 77.860 ;
        RECT 22.050 77.640 22.370 77.670 ;
        RECT 21.500 77.180 21.820 77.220 ;
        RECT 21.500 76.990 21.830 77.180 ;
        RECT 21.500 76.960 21.820 76.990 ;
        RECT 21.590 76.810 21.760 76.960 ;
        RECT 22.140 76.810 22.310 77.640 ;
        RECT 22.690 77.230 22.860 79.740 ;
        RECT 24.380 77.230 24.550 79.740 ;
        RECT 24.930 79.270 25.100 81.780 ;
        RECT 25.480 81.350 25.650 82.140 ;
        RECT 26.030 82.050 26.200 82.140 ;
        RECT 25.970 82.010 26.290 82.050 ;
        RECT 25.960 81.820 26.290 82.010 ;
        RECT 25.970 81.790 26.290 81.820 ;
        RECT 25.420 81.310 25.740 81.350 ;
        RECT 25.410 81.120 25.740 81.310 ;
        RECT 25.420 81.090 25.740 81.120 ;
        RECT 25.480 80.000 25.650 81.090 ;
        RECT 25.420 79.960 25.740 80.000 ;
        RECT 25.410 79.770 25.740 79.960 ;
        RECT 25.420 79.740 25.740 79.770 ;
        RECT 24.870 79.230 25.190 79.270 ;
        RECT 24.860 79.040 25.190 79.230 ;
        RECT 24.870 79.010 25.190 79.040 ;
        RECT 24.930 77.900 25.100 79.010 ;
        RECT 24.870 77.860 25.190 77.900 ;
        RECT 24.860 77.670 25.190 77.860 ;
        RECT 24.870 77.640 25.190 77.670 ;
        RECT 22.600 77.190 22.920 77.230 ;
        RECT 24.320 77.190 24.640 77.230 ;
        RECT 22.600 77.000 22.930 77.190 ;
        RECT 24.310 77.000 24.640 77.190 ;
        RECT 22.600 76.970 22.920 77.000 ;
        RECT 24.320 76.970 24.640 77.000 ;
        RECT 22.690 76.810 22.860 76.970 ;
        RECT 24.380 76.810 24.550 76.970 ;
        RECT 24.930 76.810 25.100 77.640 ;
        RECT 25.480 77.220 25.650 79.740 ;
        RECT 26.030 79.270 26.200 81.790 ;
        RECT 26.580 81.370 26.750 82.140 ;
        RECT 27.130 82.050 27.300 82.140 ;
        RECT 29.750 82.080 29.920 82.170 ;
        RECT 27.060 82.010 27.380 82.050 ;
        RECT 27.050 81.820 27.380 82.010 ;
        RECT 29.670 82.040 29.990 82.080 ;
        RECT 29.670 81.850 30.000 82.040 ;
        RECT 29.670 81.820 29.990 81.850 ;
        RECT 27.060 81.790 27.380 81.820 ;
        RECT 26.510 81.330 26.830 81.370 ;
        RECT 26.500 81.140 26.830 81.330 ;
        RECT 26.510 81.110 26.830 81.140 ;
        RECT 26.580 80.000 26.750 81.110 ;
        RECT 26.510 79.960 26.830 80.000 ;
        RECT 26.500 79.770 26.830 79.960 ;
        RECT 26.510 79.740 26.830 79.770 ;
        RECT 25.970 79.230 26.290 79.270 ;
        RECT 25.960 79.040 26.290 79.230 ;
        RECT 25.970 79.010 26.290 79.040 ;
        RECT 26.030 77.900 26.200 79.010 ;
        RECT 25.970 77.860 26.290 77.900 ;
        RECT 25.960 77.670 26.290 77.860 ;
        RECT 25.970 77.640 26.290 77.670 ;
        RECT 25.420 77.180 25.740 77.220 ;
        RECT 25.410 76.990 25.740 77.180 ;
        RECT 25.420 76.960 25.740 76.990 ;
        RECT 25.480 76.810 25.650 76.960 ;
        RECT 26.030 76.810 26.200 77.640 ;
        RECT 26.580 77.220 26.750 79.740 ;
        RECT 27.130 79.270 27.300 81.790 ;
        RECT 29.750 79.300 29.920 81.820 ;
        RECT 30.300 81.400 30.470 82.170 ;
        RECT 30.850 82.080 31.020 82.170 ;
        RECT 30.760 82.040 31.080 82.080 ;
        RECT 30.760 81.850 31.090 82.040 ;
        RECT 30.760 81.820 31.080 81.850 ;
        RECT 30.220 81.360 30.540 81.400 ;
        RECT 30.220 81.170 30.550 81.360 ;
        RECT 30.220 81.140 30.540 81.170 ;
        RECT 30.300 80.030 30.470 81.140 ;
        RECT 30.220 79.990 30.540 80.030 ;
        RECT 30.220 79.800 30.550 79.990 ;
        RECT 30.220 79.770 30.540 79.800 ;
        RECT 27.070 79.230 27.390 79.270 ;
        RECT 27.060 79.040 27.390 79.230 ;
        RECT 29.660 79.260 29.980 79.300 ;
        RECT 29.660 79.070 29.990 79.260 ;
        RECT 29.660 79.040 29.980 79.070 ;
        RECT 27.070 79.010 27.390 79.040 ;
        RECT 27.130 77.900 27.300 79.010 ;
        RECT 29.750 77.930 29.920 79.040 ;
        RECT 27.070 77.860 27.390 77.900 ;
        RECT 27.060 77.670 27.390 77.860 ;
        RECT 29.660 77.890 29.980 77.930 ;
        RECT 29.660 77.700 29.990 77.890 ;
        RECT 29.660 77.670 29.980 77.700 ;
        RECT 27.070 77.640 27.390 77.670 ;
        RECT 26.510 77.180 26.830 77.220 ;
        RECT 26.500 76.990 26.830 77.180 ;
        RECT 26.510 76.960 26.830 76.990 ;
        RECT 26.580 76.810 26.750 76.960 ;
        RECT 27.130 76.820 27.300 77.640 ;
        RECT 27.560 77.430 28.070 77.510 ;
        RECT 27.550 77.180 28.070 77.430 ;
        RECT 28.980 77.460 29.490 77.540 ;
        RECT 28.980 77.210 29.500 77.460 ;
        RECT 27.550 76.500 28.060 77.180 ;
        RECT 28.990 76.530 29.500 77.210 ;
        RECT 29.750 76.850 29.920 77.670 ;
        RECT 30.300 77.250 30.470 79.770 ;
        RECT 30.850 79.300 31.020 81.820 ;
        RECT 31.400 81.380 31.570 82.170 ;
        RECT 31.950 82.070 32.120 82.170 ;
        RECT 31.860 82.030 32.180 82.070 ;
        RECT 31.860 81.840 32.190 82.030 ;
        RECT 31.860 81.810 32.180 81.840 ;
        RECT 31.310 81.340 31.630 81.380 ;
        RECT 31.310 81.150 31.640 81.340 ;
        RECT 31.310 81.120 31.630 81.150 ;
        RECT 31.400 80.030 31.570 81.120 ;
        RECT 31.310 79.990 31.630 80.030 ;
        RECT 31.310 79.800 31.640 79.990 ;
        RECT 31.310 79.770 31.630 79.800 ;
        RECT 30.760 79.260 31.080 79.300 ;
        RECT 30.760 79.070 31.090 79.260 ;
        RECT 30.760 79.040 31.080 79.070 ;
        RECT 30.850 77.930 31.020 79.040 ;
        RECT 30.760 77.890 31.080 77.930 ;
        RECT 30.760 77.700 31.090 77.890 ;
        RECT 30.760 77.670 31.080 77.700 ;
        RECT 30.220 77.210 30.540 77.250 ;
        RECT 30.220 77.020 30.550 77.210 ;
        RECT 30.220 76.990 30.540 77.020 ;
        RECT 30.300 76.840 30.470 76.990 ;
        RECT 30.850 76.840 31.020 77.670 ;
        RECT 31.400 77.250 31.570 79.770 ;
        RECT 31.950 79.300 32.120 81.810 ;
        RECT 32.500 81.370 32.670 82.170 ;
        RECT 33.040 81.440 33.210 82.200 ;
        RECT 33.650 81.440 33.820 82.200 ;
        RECT 34.190 81.370 34.360 82.170 ;
        RECT 34.740 82.070 34.910 82.170 ;
        RECT 34.680 82.030 35.000 82.070 ;
        RECT 34.670 81.840 35.000 82.030 ;
        RECT 34.680 81.810 35.000 81.840 ;
        RECT 32.420 81.330 32.740 81.370 ;
        RECT 34.120 81.330 34.440 81.370 ;
        RECT 32.420 81.140 32.750 81.330 ;
        RECT 34.110 81.140 34.440 81.330 ;
        RECT 32.420 81.110 32.740 81.140 ;
        RECT 34.120 81.110 34.440 81.140 ;
        RECT 32.500 80.030 32.670 81.110 ;
        RECT 34.190 80.030 34.360 81.110 ;
        RECT 32.410 79.990 32.730 80.030 ;
        RECT 34.130 79.990 34.450 80.030 ;
        RECT 32.410 79.800 32.740 79.990 ;
        RECT 34.120 79.800 34.450 79.990 ;
        RECT 32.410 79.770 32.730 79.800 ;
        RECT 34.130 79.770 34.450 79.800 ;
        RECT 31.860 79.260 32.180 79.300 ;
        RECT 31.860 79.070 32.190 79.260 ;
        RECT 31.860 79.040 32.180 79.070 ;
        RECT 31.950 77.930 32.120 79.040 ;
        RECT 31.860 77.890 32.180 77.930 ;
        RECT 31.860 77.700 32.190 77.890 ;
        RECT 31.860 77.670 32.180 77.700 ;
        RECT 31.310 77.210 31.630 77.250 ;
        RECT 31.310 77.020 31.640 77.210 ;
        RECT 31.310 76.990 31.630 77.020 ;
        RECT 31.400 76.840 31.570 76.990 ;
        RECT 31.950 76.840 32.120 77.670 ;
        RECT 32.500 77.260 32.670 79.770 ;
        RECT 34.190 77.260 34.360 79.770 ;
        RECT 34.740 79.300 34.910 81.810 ;
        RECT 35.290 81.380 35.460 82.170 ;
        RECT 35.840 82.080 36.010 82.170 ;
        RECT 35.780 82.040 36.100 82.080 ;
        RECT 35.770 81.850 36.100 82.040 ;
        RECT 35.780 81.820 36.100 81.850 ;
        RECT 35.230 81.340 35.550 81.380 ;
        RECT 35.220 81.150 35.550 81.340 ;
        RECT 35.230 81.120 35.550 81.150 ;
        RECT 35.290 80.030 35.460 81.120 ;
        RECT 35.230 79.990 35.550 80.030 ;
        RECT 35.220 79.800 35.550 79.990 ;
        RECT 35.230 79.770 35.550 79.800 ;
        RECT 34.680 79.260 35.000 79.300 ;
        RECT 34.670 79.070 35.000 79.260 ;
        RECT 34.680 79.040 35.000 79.070 ;
        RECT 34.740 77.930 34.910 79.040 ;
        RECT 34.680 77.890 35.000 77.930 ;
        RECT 34.670 77.700 35.000 77.890 ;
        RECT 34.680 77.670 35.000 77.700 ;
        RECT 32.410 77.220 32.730 77.260 ;
        RECT 34.130 77.220 34.450 77.260 ;
        RECT 32.410 77.030 32.740 77.220 ;
        RECT 34.120 77.030 34.450 77.220 ;
        RECT 32.410 77.000 32.730 77.030 ;
        RECT 34.130 77.000 34.450 77.030 ;
        RECT 32.500 76.840 32.670 77.000 ;
        RECT 34.190 76.840 34.360 77.000 ;
        RECT 34.740 76.840 34.910 77.670 ;
        RECT 35.290 77.250 35.460 79.770 ;
        RECT 35.840 79.300 36.010 81.820 ;
        RECT 36.390 81.400 36.560 82.170 ;
        RECT 36.940 82.080 37.110 82.170 ;
        RECT 36.870 82.040 37.190 82.080 ;
        RECT 36.860 81.850 37.190 82.040 ;
        RECT 36.870 81.820 37.190 81.850 ;
        RECT 36.320 81.360 36.640 81.400 ;
        RECT 36.310 81.170 36.640 81.360 ;
        RECT 36.320 81.140 36.640 81.170 ;
        RECT 36.390 80.030 36.560 81.140 ;
        RECT 36.320 79.990 36.640 80.030 ;
        RECT 36.310 79.800 36.640 79.990 ;
        RECT 36.320 79.770 36.640 79.800 ;
        RECT 35.780 79.260 36.100 79.300 ;
        RECT 35.770 79.070 36.100 79.260 ;
        RECT 35.780 79.040 36.100 79.070 ;
        RECT 35.840 77.930 36.010 79.040 ;
        RECT 35.780 77.890 36.100 77.930 ;
        RECT 35.770 77.700 36.100 77.890 ;
        RECT 35.780 77.670 36.100 77.700 ;
        RECT 35.230 77.210 35.550 77.250 ;
        RECT 35.220 77.020 35.550 77.210 ;
        RECT 35.230 76.990 35.550 77.020 ;
        RECT 35.290 76.840 35.460 76.990 ;
        RECT 35.840 76.840 36.010 77.670 ;
        RECT 36.390 77.250 36.560 79.770 ;
        RECT 36.940 79.300 37.110 81.820 ;
        RECT 39.940 81.360 40.110 82.100 ;
        RECT 40.490 82.060 40.660 82.100 ;
        RECT 40.420 82.020 40.740 82.060 ;
        RECT 40.410 81.830 40.740 82.020 ;
        RECT 40.420 81.800 40.740 81.830 ;
        RECT 39.860 81.320 40.180 81.360 ;
        RECT 39.850 81.130 40.180 81.320 ;
        RECT 39.860 81.100 40.180 81.130 ;
        RECT 39.940 80.020 40.110 81.100 ;
        RECT 39.870 79.980 40.190 80.020 ;
        RECT 39.860 79.790 40.190 79.980 ;
        RECT 39.870 79.760 40.190 79.790 ;
        RECT 36.880 79.260 37.200 79.300 ;
        RECT 36.870 79.070 37.200 79.260 ;
        RECT 36.880 79.040 37.200 79.070 ;
        RECT 36.940 77.930 37.110 79.040 ;
        RECT 36.880 77.890 37.200 77.930 ;
        RECT 36.870 77.700 37.200 77.890 ;
        RECT 36.880 77.670 37.200 77.700 ;
        RECT 36.320 77.210 36.640 77.250 ;
        RECT 36.310 77.020 36.640 77.210 ;
        RECT 36.320 76.990 36.640 77.020 ;
        RECT 36.390 76.840 36.560 76.990 ;
        RECT 36.940 76.850 37.110 77.670 ;
        RECT 37.370 77.460 37.880 77.540 ;
        RECT 37.360 77.210 37.880 77.460 ;
        RECT 39.940 77.250 40.110 79.760 ;
        RECT 40.490 79.290 40.660 81.800 ;
        RECT 41.040 81.370 41.210 82.100 ;
        RECT 41.590 82.070 41.760 82.100 ;
        RECT 41.520 82.030 41.840 82.070 ;
        RECT 41.510 81.840 41.840 82.030 ;
        RECT 41.520 81.810 41.840 81.840 ;
        RECT 40.970 81.330 41.290 81.370 ;
        RECT 40.960 81.140 41.290 81.330 ;
        RECT 40.970 81.110 41.290 81.140 ;
        RECT 41.040 80.020 41.210 81.110 ;
        RECT 40.970 79.980 41.290 80.020 ;
        RECT 40.960 79.790 41.290 79.980 ;
        RECT 40.970 79.760 41.290 79.790 ;
        RECT 40.420 79.250 40.740 79.290 ;
        RECT 40.410 79.060 40.740 79.250 ;
        RECT 40.420 79.030 40.740 79.060 ;
        RECT 40.490 77.920 40.660 79.030 ;
        RECT 40.420 77.880 40.740 77.920 ;
        RECT 40.410 77.690 40.740 77.880 ;
        RECT 40.420 77.660 40.740 77.690 ;
        RECT 39.870 77.210 40.190 77.250 ;
        RECT 37.360 76.530 37.870 77.210 ;
        RECT 39.860 77.020 40.190 77.210 ;
        RECT 39.870 76.990 40.190 77.020 ;
        RECT 39.940 76.920 40.110 76.990 ;
        RECT 40.490 76.920 40.660 77.660 ;
        RECT 41.040 77.240 41.210 79.760 ;
        RECT 41.590 79.290 41.760 81.810 ;
        RECT 42.140 81.390 42.310 82.100 ;
        RECT 42.690 82.070 42.860 82.100 ;
        RECT 42.610 82.030 42.930 82.070 ;
        RECT 42.600 81.840 42.930 82.030 ;
        RECT 42.610 81.810 42.930 81.840 ;
        RECT 42.060 81.350 42.380 81.390 ;
        RECT 42.050 81.160 42.380 81.350 ;
        RECT 42.060 81.130 42.380 81.160 ;
        RECT 42.140 80.020 42.310 81.130 ;
        RECT 42.060 79.980 42.380 80.020 ;
        RECT 42.050 79.790 42.380 79.980 ;
        RECT 42.060 79.760 42.380 79.790 ;
        RECT 41.520 79.250 41.840 79.290 ;
        RECT 41.510 79.060 41.840 79.250 ;
        RECT 41.520 79.030 41.840 79.060 ;
        RECT 41.590 77.920 41.760 79.030 ;
        RECT 41.520 77.880 41.840 77.920 ;
        RECT 41.510 77.690 41.840 77.880 ;
        RECT 41.520 77.660 41.840 77.690 ;
        RECT 40.970 77.200 41.290 77.240 ;
        RECT 40.960 77.010 41.290 77.200 ;
        RECT 40.970 76.980 41.290 77.010 ;
        RECT 41.040 76.920 41.210 76.980 ;
        RECT 41.590 76.920 41.760 77.660 ;
        RECT 42.140 77.240 42.310 79.760 ;
        RECT 42.690 79.290 42.860 81.810 ;
        RECT 42.620 79.250 42.940 79.290 ;
        RECT 42.610 79.060 42.940 79.250 ;
        RECT 42.620 79.030 42.940 79.060 ;
        RECT 42.690 77.920 42.860 79.030 ;
        RECT 42.620 77.880 42.940 77.920 ;
        RECT 42.610 77.690 42.940 77.880 ;
        RECT 43.400 77.720 43.570 78.940 ;
        RECT 42.620 77.660 42.940 77.690 ;
        RECT 42.060 77.200 42.380 77.240 ;
        RECT 42.050 77.010 42.380 77.200 ;
        RECT 42.060 76.980 42.380 77.010 ;
        RECT 42.140 76.920 42.310 76.980 ;
        RECT 42.690 76.920 42.860 77.660 ;
        RECT 43.110 77.270 43.620 77.530 ;
        RECT 43.100 77.200 43.620 77.270 ;
        RECT 43.100 76.520 43.610 77.200 ;
        RECT 206.500 76.260 207.010 86.620 ;
        RECT 207.180 85.830 213.160 86.060 ;
        RECT 206.500 76.240 207.020 76.260 ;
        RECT -11.660 75.080 -11.340 75.110 ;
        RECT -11.670 74.890 -11.340 75.080 ;
        RECT -11.660 74.850 -11.340 74.890 ;
        RECT -11.580 74.820 -11.410 74.850 ;
        RECT -143.420 74.440 -142.890 74.650 ;
        RECT -150.440 73.960 -142.890 74.440 ;
        RECT 74.490 74.230 74.720 74.240 ;
        RECT 74.470 74.060 79.130 74.230 ;
        RECT 74.490 74.050 74.720 74.060 ;
        RECT -150.440 73.930 -143.080 73.960 ;
        RECT 80.030 73.580 80.220 73.590 ;
        RECT 75.690 73.540 79.490 73.550 ;
        RECT 80.000 73.540 80.260 73.580 ;
        RECT 75.690 73.380 80.260 73.540 ;
        RECT 79.260 73.370 80.260 73.380 ;
        RECT 79.260 72.910 79.490 73.370 ;
        RECT 80.000 73.260 80.260 73.370 ;
        RECT 80.030 72.910 80.220 72.920 ;
        RECT -150.440 72.170 -142.910 72.720 ;
        RECT -14.300 72.380 -14.130 72.540 ;
        RECT -14.360 72.350 -14.040 72.380 ;
        RECT -152.130 59.200 -150.650 59.450 ;
        RECT -150.440 59.260 -149.930 72.170 ;
        RECT -143.580 72.160 -142.910 72.170 ;
        RECT -14.370 72.160 -14.040 72.350 ;
        RECT -147.280 71.270 -143.820 71.710 ;
        RECT -149.210 71.170 -143.820 71.270 ;
        RECT -149.210 71.100 -143.930 71.170 ;
        RECT -149.210 60.190 -149.040 71.100 ;
        RECT -148.710 70.690 -144.480 70.710 ;
        RECT -148.730 60.580 -144.400 70.690 ;
        RECT -148.670 60.530 -148.500 60.580 ;
        RECT -144.100 60.190 -143.930 71.100 ;
        RECT -149.210 60.020 -143.930 60.190 ;
        RECT -144.170 60.010 -143.930 60.020 ;
        RECT -143.420 59.260 -142.910 72.160 ;
        RECT -14.360 72.120 -14.040 72.160 ;
        RECT -14.300 69.610 -14.130 72.120 ;
        RECT -13.750 71.710 -13.580 72.540 ;
        RECT -13.200 72.390 -13.030 72.540 ;
        RECT -13.260 72.360 -12.940 72.390 ;
        RECT -13.270 72.170 -12.940 72.360 ;
        RECT -13.260 72.130 -12.940 72.170 ;
        RECT -13.810 71.680 -13.490 71.710 ;
        RECT -13.820 71.490 -13.490 71.680 ;
        RECT -13.810 71.450 -13.490 71.490 ;
        RECT -13.750 70.340 -13.580 71.450 ;
        RECT -13.810 70.310 -13.490 70.340 ;
        RECT -13.820 70.120 -13.490 70.310 ;
        RECT -13.810 70.080 -13.490 70.120 ;
        RECT -14.360 69.580 -14.040 69.610 ;
        RECT -14.370 69.390 -14.040 69.580 ;
        RECT -14.360 69.350 -14.040 69.390 ;
        RECT -14.300 68.270 -14.130 69.350 ;
        RECT -14.370 68.240 -14.050 68.270 ;
        RECT -14.380 68.050 -14.050 68.240 ;
        RECT -14.370 68.010 -14.050 68.050 ;
        RECT -14.840 67.180 -14.670 67.940 ;
        RECT -14.300 67.210 -14.130 68.010 ;
        RECT -13.750 67.570 -13.580 70.080 ;
        RECT -13.200 69.610 -13.030 72.130 ;
        RECT -12.650 71.710 -12.480 72.540 ;
        RECT -12.100 72.390 -11.930 72.540 ;
        RECT -12.170 72.360 -11.850 72.390 ;
        RECT -12.180 72.170 -11.850 72.360 ;
        RECT -12.170 72.130 -11.850 72.170 ;
        RECT -12.710 71.680 -12.390 71.710 ;
        RECT -12.720 71.490 -12.390 71.680 ;
        RECT -12.710 71.450 -12.390 71.490 ;
        RECT -12.650 70.340 -12.480 71.450 ;
        RECT -12.710 70.310 -12.390 70.340 ;
        RECT -12.720 70.120 -12.390 70.310 ;
        RECT -12.710 70.080 -12.390 70.120 ;
        RECT -13.260 69.580 -12.940 69.610 ;
        RECT -13.270 69.390 -12.940 69.580 ;
        RECT -13.260 69.350 -12.940 69.390 ;
        RECT -13.200 68.260 -13.030 69.350 ;
        RECT -13.260 68.230 -12.940 68.260 ;
        RECT -13.270 68.040 -12.940 68.230 ;
        RECT -13.260 68.000 -12.940 68.040 ;
        RECT -13.810 67.540 -13.490 67.570 ;
        RECT -13.820 67.350 -13.490 67.540 ;
        RECT -13.810 67.310 -13.490 67.350 ;
        RECT -13.750 67.210 -13.580 67.310 ;
        RECT -13.200 67.210 -13.030 68.000 ;
        RECT -12.650 67.560 -12.480 70.080 ;
        RECT -12.100 69.610 -11.930 72.130 ;
        RECT -11.550 71.710 -11.380 72.530 ;
        RECT -11.130 72.170 -10.620 72.850 ;
        RECT 79.260 72.700 80.270 72.910 ;
        RECT 74.490 72.620 74.720 72.630 ;
        RECT 74.470 72.450 78.950 72.620 ;
        RECT 74.490 72.440 74.720 72.450 ;
        RECT -11.130 71.920 -10.610 72.170 ;
        RECT 79.260 71.940 79.490 72.700 ;
        RECT 80.000 72.590 80.260 72.700 ;
        RECT -11.120 71.840 -10.610 71.920 ;
        RECT 75.710 71.770 79.490 71.940 ;
        RECT -11.610 71.680 -11.290 71.710 ;
        RECT -11.620 71.490 -11.290 71.680 ;
        RECT -11.610 71.450 -11.290 71.490 ;
        RECT -11.550 70.340 -11.380 71.450 ;
        RECT -9.550 71.210 -7.160 71.580 ;
        RECT -11.610 70.310 -11.290 70.340 ;
        RECT -11.620 70.120 -11.290 70.310 ;
        RECT -11.610 70.080 -11.290 70.120 ;
        RECT -12.170 69.580 -11.850 69.610 ;
        RECT -12.180 69.390 -11.850 69.580 ;
        RECT -12.170 69.350 -11.850 69.390 ;
        RECT -12.100 68.240 -11.930 69.350 ;
        RECT -12.170 68.210 -11.850 68.240 ;
        RECT -12.180 68.020 -11.850 68.210 ;
        RECT -12.170 67.980 -11.850 68.020 ;
        RECT -12.710 67.530 -12.390 67.560 ;
        RECT -12.720 67.340 -12.390 67.530 ;
        RECT -12.710 67.300 -12.390 67.340 ;
        RECT -12.650 67.210 -12.480 67.300 ;
        RECT -12.100 67.210 -11.930 67.980 ;
        RECT -11.550 67.560 -11.380 70.080 ;
        RECT -9.500 67.950 -7.160 71.210 ;
        RECT 74.490 71.020 74.720 71.030 ;
        RECT 74.470 70.850 78.970 71.020 ;
        RECT 74.490 70.840 74.720 70.850 ;
        RECT 75.710 70.840 76.040 70.850 ;
        RECT 76.670 70.840 77.000 70.850 ;
        RECT 77.630 70.840 77.960 70.850 ;
        RECT 78.590 70.840 78.920 70.850 ;
        RECT 79.260 70.330 79.490 71.770 ;
        RECT 79.980 71.580 80.410 71.600 ;
        RECT 79.960 71.410 80.410 71.580 ;
        RECT 79.980 71.390 80.410 71.410 ;
        RECT 75.710 70.160 79.490 70.330 ;
        RECT 75.770 69.880 76.200 69.900 ;
        RECT 75.750 69.710 76.200 69.880 ;
        RECT 75.770 69.690 76.200 69.710 ;
        RECT 74.490 69.400 74.720 69.410 ;
        RECT 74.470 69.230 78.970 69.400 ;
        RECT 74.490 69.220 74.720 69.230 ;
        RECT 79.260 68.730 79.490 70.160 ;
        RECT 79.980 69.970 80.410 69.990 ;
        RECT 79.960 69.800 80.410 69.970 ;
        RECT 79.980 69.780 80.410 69.800 ;
        RECT 75.720 68.720 79.490 68.730 ;
        RECT 75.710 68.560 79.490 68.720 ;
        RECT 75.710 68.550 76.040 68.560 ;
        RECT 77.630 68.550 77.960 68.560 ;
        RECT 78.590 68.550 78.920 68.560 ;
        RECT 76.770 68.240 77.200 68.260 ;
        RECT 76.770 68.070 77.220 68.240 ;
        RECT 76.770 68.050 77.200 68.070 ;
        RECT -9.500 67.940 -7.170 67.950 ;
        RECT 74.490 67.800 74.720 67.810 ;
        RECT 74.470 67.630 78.920 67.800 ;
        RECT 74.490 67.620 74.720 67.630 ;
        RECT 75.710 67.620 76.040 67.630 ;
        RECT 76.670 67.620 77.000 67.630 ;
        RECT 77.630 67.620 77.960 67.630 ;
        RECT 78.590 67.620 78.920 67.630 ;
        RECT -11.620 67.530 -11.300 67.560 ;
        RECT -11.630 67.340 -11.300 67.530 ;
        RECT -11.620 67.300 -11.300 67.340 ;
        RECT -11.550 67.210 -11.380 67.300 ;
        RECT 79.260 67.110 79.490 68.560 ;
        RECT 79.970 68.360 80.400 68.380 ;
        RECT 79.950 68.190 80.400 68.360 ;
        RECT 79.970 68.170 80.400 68.190 ;
        RECT 75.700 66.940 79.490 67.110 ;
        RECT 77.680 66.660 78.110 66.680 ;
        RECT 77.660 66.490 78.110 66.660 ;
        RECT 77.680 66.470 78.110 66.490 ;
        RECT 74.490 66.180 74.720 66.190 ;
        RECT 74.470 66.010 78.970 66.180 ;
        RECT 74.490 66.000 74.720 66.010 ;
        RECT 75.710 65.490 76.040 65.500 ;
        RECT 76.670 65.490 77.000 65.500 ;
        RECT 77.630 65.490 77.960 65.500 ;
        RECT 78.590 65.490 78.920 65.500 ;
        RECT 79.260 65.490 79.490 66.940 ;
        RECT 79.980 66.740 80.410 66.760 ;
        RECT 79.960 66.570 80.410 66.740 ;
        RECT 79.980 66.550 80.410 66.570 ;
        RECT 75.700 65.320 79.490 65.490 ;
        RECT 74.490 64.580 74.720 64.590 ;
        RECT 74.470 64.570 78.890 64.580 ;
        RECT 74.470 64.410 78.920 64.570 ;
        RECT 74.490 64.400 74.720 64.410 ;
        RECT 75.710 64.400 76.040 64.410 ;
        RECT 76.670 64.400 77.000 64.410 ;
        RECT 77.630 64.400 77.960 64.410 ;
        RECT 78.590 64.400 78.920 64.410 ;
        RECT 79.260 63.900 79.490 65.320 ;
        RECT 79.970 65.130 80.400 65.150 ;
        RECT 79.950 64.960 80.400 65.130 ;
        RECT 79.970 64.940 80.400 64.960 ;
        RECT 75.700 63.730 79.500 63.900 ;
        RECT 75.710 63.720 76.040 63.730 ;
        RECT 76.670 63.720 77.000 63.730 ;
        RECT 77.630 63.720 77.960 63.730 ;
        RECT 78.590 63.720 78.920 63.730 ;
        RECT 74.490 62.950 74.720 62.970 ;
        RECT 75.710 62.950 76.040 62.960 ;
        RECT 76.670 62.950 77.000 62.960 ;
        RECT 77.630 62.950 77.960 62.960 ;
        RECT 78.590 62.950 78.920 62.960 ;
        RECT 74.470 62.780 78.930 62.950 ;
        RECT 79.260 62.290 79.490 63.730 ;
        RECT 79.770 63.090 79.980 63.520 ;
        RECT 79.790 63.070 79.960 63.090 ;
        RECT 75.700 62.120 79.490 62.290 ;
        RECT 75.710 62.110 76.040 62.120 ;
        RECT 76.670 62.110 77.000 62.120 ;
        RECT 77.630 62.110 77.960 62.120 ;
        RECT 78.590 62.110 78.920 62.120 ;
        RECT 79.970 61.930 80.400 61.950 ;
        RECT 79.950 61.760 80.400 61.930 ;
        RECT 79.970 61.740 80.400 61.760 ;
        RECT 80.680 60.950 81.050 75.820 ;
        RECT 206.490 74.460 207.020 76.240 ;
        RECT 207.420 74.770 213.070 85.830 ;
        RECT 207.360 74.760 213.070 74.770 ;
        RECT 207.360 74.590 213.150 74.760 ;
        RECT 207.360 74.580 213.060 74.590 ;
        RECT 207.420 74.510 207.590 74.580 ;
        RECT 206.490 74.440 207.010 74.460 ;
        RECT 206.500 73.930 207.010 74.440 ;
        RECT 213.520 74.010 214.030 86.620 ;
        RECT 214.270 80.600 215.730 80.640 ;
        RECT 214.260 80.430 215.730 80.600 ;
        RECT 214.270 80.390 215.730 80.430 ;
        RECT 206.480 73.720 207.010 73.930 ;
        RECT 211.590 73.720 214.030 74.010 ;
        RECT 206.480 73.240 214.030 73.720 ;
        RECT 206.670 73.210 214.030 73.240 ;
        RECT 206.500 71.450 214.030 72.000 ;
        RECT 206.500 71.440 207.170 71.450 ;
        RECT 80.680 60.700 81.060 60.950 ;
        RECT 76.730 60.220 77.160 60.240 ;
        RECT 77.670 60.220 78.100 60.240 ;
        RECT 79.930 60.220 80.360 60.240 ;
        RECT 76.710 60.050 77.160 60.220 ;
        RECT 77.650 60.050 78.100 60.220 ;
        RECT 78.620 60.200 79.050 60.220 ;
        RECT 76.730 60.030 77.160 60.050 ;
        RECT 77.670 60.030 78.100 60.050 ;
        RECT 78.600 60.030 79.050 60.200 ;
        RECT 79.910 60.050 80.360 60.220 ;
        RECT 79.930 60.030 80.360 60.050 ;
        RECT 78.620 60.010 79.050 60.030 ;
        RECT -150.440 58.750 -142.910 59.260 ;
        RECT -152.140 52.730 -150.680 52.770 ;
        RECT -152.140 52.560 -150.670 52.730 ;
        RECT -152.140 52.520 -150.680 52.560 ;
        RECT -150.440 46.140 -149.930 58.750 ;
        RECT -149.570 57.960 -143.590 58.190 ;
        RECT -149.480 46.900 -143.830 57.960 ;
        RECT -143.420 48.390 -142.910 58.750 ;
        RECT -143.430 48.370 -142.910 48.390 ;
        RECT 206.500 58.540 207.010 71.440 ;
        RECT 207.410 70.550 210.870 70.990 ;
        RECT 207.410 70.450 212.800 70.550 ;
        RECT 207.520 70.380 212.800 70.450 ;
        RECT 207.520 59.470 207.690 70.380 ;
        RECT 208.070 69.970 212.300 69.990 ;
        RECT 207.990 59.860 212.320 69.970 ;
        RECT 212.090 59.810 212.260 59.860 ;
        RECT 212.630 59.470 212.800 70.380 ;
        RECT 207.520 59.300 212.800 59.470 ;
        RECT 207.520 59.290 207.760 59.300 ;
        RECT 213.520 58.540 214.030 71.450 ;
        RECT 206.500 58.030 214.030 58.540 ;
        RECT 214.240 58.480 215.720 58.730 ;
        RECT -149.480 46.890 -143.770 46.900 ;
        RECT -149.560 46.720 -143.770 46.890 ;
        RECT -149.470 46.710 -143.770 46.720 ;
        RECT -144.000 46.640 -143.830 46.710 ;
        RECT -143.430 46.590 -142.900 48.370 ;
        RECT 206.500 47.670 207.010 58.030 ;
        RECT 207.180 57.240 213.160 57.470 ;
        RECT 206.500 47.650 207.020 47.670 ;
        RECT -143.420 46.570 -142.900 46.590 ;
        RECT -150.440 45.850 -148.000 46.140 ;
        RECT -143.420 46.060 -142.910 46.570 ;
        RECT -143.420 45.850 -142.890 46.060 ;
        RECT 206.490 45.870 207.020 47.650 ;
        RECT 207.420 46.180 213.070 57.240 ;
        RECT 207.360 46.170 213.070 46.180 ;
        RECT 207.360 46.000 213.150 46.170 ;
        RECT 207.360 45.990 213.060 46.000 ;
        RECT 207.420 45.920 207.590 45.990 ;
        RECT 206.490 45.850 207.010 45.870 ;
        RECT -150.440 45.370 -142.890 45.850 ;
        RECT -150.440 45.340 -143.080 45.370 ;
        RECT 206.500 45.340 207.010 45.850 ;
        RECT 213.520 45.420 214.030 58.030 ;
        RECT 214.270 52.010 215.730 52.050 ;
        RECT 214.260 51.840 215.730 52.010 ;
        RECT 214.270 51.800 215.730 51.840 ;
        RECT 206.480 45.130 207.010 45.340 ;
        RECT 211.590 45.130 214.030 45.420 ;
        RECT 206.480 44.650 214.030 45.130 ;
        RECT 206.670 44.620 214.030 44.650 ;
        RECT -150.440 43.580 -142.910 44.130 ;
        RECT -152.130 30.610 -150.650 30.860 ;
        RECT -150.440 30.670 -149.930 43.580 ;
        RECT -143.580 43.570 -142.910 43.580 ;
        RECT -147.280 42.680 -143.820 43.120 ;
        RECT -149.210 42.580 -143.820 42.680 ;
        RECT -149.210 42.510 -143.930 42.580 ;
        RECT -149.210 31.600 -149.040 42.510 ;
        RECT -148.710 42.100 -144.480 42.120 ;
        RECT -148.730 31.990 -144.400 42.100 ;
        RECT -148.670 31.940 -148.500 31.990 ;
        RECT -144.100 31.600 -143.930 42.510 ;
        RECT -149.210 31.430 -143.930 31.600 ;
        RECT -144.170 31.420 -143.930 31.430 ;
        RECT -143.420 30.670 -142.910 43.570 ;
        RECT -150.440 30.160 -142.910 30.670 ;
        RECT -152.140 24.140 -150.680 24.180 ;
        RECT -152.140 23.970 -150.670 24.140 ;
        RECT -152.140 23.930 -150.680 23.970 ;
        RECT -150.440 17.550 -149.930 30.160 ;
        RECT -149.570 29.370 -143.590 29.600 ;
        RECT -149.480 18.310 -143.830 29.370 ;
        RECT -143.420 19.800 -142.910 30.160 ;
        RECT -143.430 19.780 -142.910 19.800 ;
        RECT 206.500 42.860 214.030 43.410 ;
        RECT 206.500 42.850 207.170 42.860 ;
        RECT 206.500 29.950 207.010 42.850 ;
        RECT 207.410 41.960 210.870 42.400 ;
        RECT 207.410 41.860 212.800 41.960 ;
        RECT 207.520 41.790 212.800 41.860 ;
        RECT 207.520 30.880 207.690 41.790 ;
        RECT 208.070 41.380 212.300 41.400 ;
        RECT 207.990 31.270 212.320 41.380 ;
        RECT 212.090 31.220 212.260 31.270 ;
        RECT 212.630 30.880 212.800 41.790 ;
        RECT 207.520 30.710 212.800 30.880 ;
        RECT 207.520 30.700 207.760 30.710 ;
        RECT 213.520 29.950 214.030 42.860 ;
        RECT 206.500 29.440 214.030 29.950 ;
        RECT 214.240 29.890 215.720 30.140 ;
        RECT -149.480 18.300 -143.770 18.310 ;
        RECT -149.560 18.130 -143.770 18.300 ;
        RECT -149.470 18.120 -143.770 18.130 ;
        RECT -144.000 18.050 -143.830 18.120 ;
        RECT -143.430 18.000 -142.900 19.780 ;
        RECT 206.500 19.080 207.010 29.440 ;
        RECT 207.180 28.650 213.160 28.880 ;
        RECT 206.500 19.060 207.020 19.080 ;
        RECT -143.420 17.980 -142.900 18.000 ;
        RECT -150.440 17.260 -148.000 17.550 ;
        RECT -143.420 17.470 -142.910 17.980 ;
        RECT -143.420 17.260 -142.890 17.470 ;
        RECT 206.490 17.280 207.020 19.060 ;
        RECT 207.420 17.590 213.070 28.650 ;
        RECT 207.360 17.580 213.070 17.590 ;
        RECT 207.360 17.410 213.150 17.580 ;
        RECT 207.360 17.400 213.060 17.410 ;
        RECT 207.420 17.330 207.590 17.400 ;
        RECT 206.490 17.260 207.010 17.280 ;
        RECT -150.440 16.780 -142.890 17.260 ;
        RECT -150.440 16.750 -143.080 16.780 ;
        RECT 206.500 16.750 207.010 17.260 ;
        RECT 213.520 16.830 214.030 29.440 ;
        RECT 214.270 23.420 215.730 23.460 ;
        RECT 214.260 23.250 215.730 23.420 ;
        RECT 214.270 23.210 215.730 23.250 ;
        RECT 206.480 16.540 207.010 16.750 ;
        RECT 211.590 16.540 214.030 16.830 ;
        RECT 206.480 16.060 214.030 16.540 ;
        RECT 206.670 16.030 214.030 16.060 ;
        RECT -150.440 14.990 -142.910 15.540 ;
        RECT -152.130 2.020 -150.650 2.270 ;
        RECT -150.440 2.080 -149.930 14.990 ;
        RECT -143.580 14.980 -142.910 14.990 ;
        RECT -147.280 14.090 -143.820 14.530 ;
        RECT -149.210 13.990 -143.820 14.090 ;
        RECT -149.210 13.920 -143.930 13.990 ;
        RECT -149.210 3.010 -149.040 13.920 ;
        RECT -148.710 13.510 -144.480 13.530 ;
        RECT -148.730 3.400 -144.400 13.510 ;
        RECT -148.670 3.350 -148.500 3.400 ;
        RECT -144.100 3.010 -143.930 13.920 ;
        RECT -149.210 2.840 -143.930 3.010 ;
        RECT -144.170 2.830 -143.930 2.840 ;
        RECT -143.420 2.080 -142.910 14.980 ;
        RECT -150.440 1.570 -142.910 2.080 ;
        RECT -152.140 -4.450 -150.680 -4.410 ;
        RECT -152.140 -4.620 -150.670 -4.450 ;
        RECT -152.140 -4.660 -150.680 -4.620 ;
        RECT -150.440 -11.040 -149.930 1.570 ;
        RECT -149.570 0.780 -143.590 1.010 ;
        RECT -149.480 -10.280 -143.830 0.780 ;
        RECT -143.420 -8.790 -142.910 1.570 ;
        RECT -143.430 -8.810 -142.910 -8.790 ;
        RECT 206.500 14.270 214.030 14.820 ;
        RECT 206.500 14.260 207.170 14.270 ;
        RECT 206.500 1.360 207.010 14.260 ;
        RECT 207.410 13.370 210.870 13.810 ;
        RECT 207.410 13.270 212.800 13.370 ;
        RECT 207.520 13.200 212.800 13.270 ;
        RECT 207.520 2.290 207.690 13.200 ;
        RECT 208.070 12.790 212.300 12.810 ;
        RECT 207.990 2.680 212.320 12.790 ;
        RECT 212.090 2.630 212.260 2.680 ;
        RECT 212.630 2.290 212.800 13.200 ;
        RECT 207.520 2.120 212.800 2.290 ;
        RECT 207.520 2.110 207.760 2.120 ;
        RECT 213.520 1.360 214.030 14.270 ;
        RECT 206.500 0.850 214.030 1.360 ;
        RECT 214.240 1.300 215.720 1.550 ;
        RECT -149.480 -10.290 -143.770 -10.280 ;
        RECT -149.560 -10.460 -143.770 -10.290 ;
        RECT -149.470 -10.470 -143.770 -10.460 ;
        RECT -144.000 -10.540 -143.830 -10.470 ;
        RECT -143.430 -10.590 -142.900 -8.810 ;
        RECT 206.500 -9.510 207.010 0.850 ;
        RECT 207.180 0.060 213.160 0.290 ;
        RECT 206.500 -9.530 207.020 -9.510 ;
        RECT -143.420 -10.610 -142.900 -10.590 ;
        RECT -150.440 -11.330 -148.000 -11.040 ;
        RECT -143.420 -11.120 -142.910 -10.610 ;
        RECT -143.420 -11.330 -142.890 -11.120 ;
        RECT 206.490 -11.310 207.020 -9.530 ;
        RECT 207.420 -11.000 213.070 0.060 ;
        RECT 207.360 -11.010 213.070 -11.000 ;
        RECT 207.360 -11.180 213.150 -11.010 ;
        RECT 207.360 -11.190 213.060 -11.180 ;
        RECT 207.420 -11.260 207.590 -11.190 ;
        RECT 206.490 -11.330 207.010 -11.310 ;
        RECT -150.440 -11.810 -142.890 -11.330 ;
        RECT -150.440 -11.840 -143.080 -11.810 ;
        RECT 206.500 -11.840 207.010 -11.330 ;
        RECT 213.520 -11.760 214.030 0.850 ;
        RECT 214.270 -5.170 215.730 -5.130 ;
        RECT 214.260 -5.340 215.730 -5.170 ;
        RECT 214.270 -5.380 215.730 -5.340 ;
        RECT 206.480 -12.050 207.010 -11.840 ;
        RECT 211.590 -12.050 214.030 -11.760 ;
        RECT 206.480 -12.530 214.030 -12.050 ;
        RECT 206.670 -12.560 214.030 -12.530 ;
        RECT -150.440 -13.600 -142.910 -13.050 ;
        RECT -152.130 -26.570 -150.650 -26.320 ;
        RECT -150.440 -26.510 -149.930 -13.600 ;
        RECT -143.580 -13.610 -142.910 -13.600 ;
        RECT -147.280 -14.500 -143.820 -14.060 ;
        RECT -149.210 -14.600 -143.820 -14.500 ;
        RECT -149.210 -14.670 -143.930 -14.600 ;
        RECT -149.210 -25.580 -149.040 -14.670 ;
        RECT -148.710 -15.080 -144.480 -15.060 ;
        RECT -148.730 -25.190 -144.400 -15.080 ;
        RECT -148.670 -25.240 -148.500 -25.190 ;
        RECT -144.100 -25.580 -143.930 -14.670 ;
        RECT -149.210 -25.750 -143.930 -25.580 ;
        RECT -144.170 -25.760 -143.930 -25.750 ;
        RECT -143.420 -26.510 -142.910 -13.610 ;
        RECT -150.440 -27.020 -142.910 -26.510 ;
        RECT -152.140 -33.040 -150.680 -33.000 ;
        RECT -152.140 -33.210 -150.670 -33.040 ;
        RECT -152.140 -33.250 -150.680 -33.210 ;
        RECT -150.440 -39.630 -149.930 -27.020 ;
        RECT -149.570 -27.810 -143.590 -27.580 ;
        RECT -149.480 -38.870 -143.830 -27.810 ;
        RECT -143.420 -37.380 -142.910 -27.020 ;
        RECT -143.430 -37.400 -142.910 -37.380 ;
        RECT 206.500 -14.320 214.030 -13.770 ;
        RECT 206.500 -14.330 207.170 -14.320 ;
        RECT 206.500 -27.230 207.010 -14.330 ;
        RECT 207.410 -15.220 210.870 -14.780 ;
        RECT 207.410 -15.320 212.800 -15.220 ;
        RECT 207.520 -15.390 212.800 -15.320 ;
        RECT 207.520 -26.300 207.690 -15.390 ;
        RECT 208.070 -15.800 212.300 -15.780 ;
        RECT 207.990 -25.910 212.320 -15.800 ;
        RECT 212.090 -25.960 212.260 -25.910 ;
        RECT 212.630 -26.300 212.800 -15.390 ;
        RECT 207.520 -26.470 212.800 -26.300 ;
        RECT 207.520 -26.480 207.760 -26.470 ;
        RECT 213.520 -27.230 214.030 -14.320 ;
        RECT 206.500 -27.740 214.030 -27.230 ;
        RECT 214.240 -27.290 215.720 -27.040 ;
        RECT -149.480 -38.880 -143.770 -38.870 ;
        RECT -149.560 -39.050 -143.770 -38.880 ;
        RECT -149.470 -39.060 -143.770 -39.050 ;
        RECT -144.000 -39.130 -143.830 -39.060 ;
        RECT -143.430 -39.180 -142.900 -37.400 ;
        RECT 206.500 -38.100 207.010 -27.740 ;
        RECT 207.180 -28.530 213.160 -28.300 ;
        RECT 206.500 -38.120 207.020 -38.100 ;
        RECT -143.420 -39.200 -142.900 -39.180 ;
        RECT -150.440 -39.920 -148.000 -39.630 ;
        RECT -143.420 -39.710 -142.910 -39.200 ;
        RECT -143.420 -39.920 -142.890 -39.710 ;
        RECT 206.490 -39.900 207.020 -38.120 ;
        RECT 207.420 -39.590 213.070 -28.530 ;
        RECT 207.360 -39.600 213.070 -39.590 ;
        RECT 207.360 -39.770 213.150 -39.600 ;
        RECT 207.360 -39.780 213.060 -39.770 ;
        RECT 207.420 -39.850 207.590 -39.780 ;
        RECT 206.490 -39.920 207.010 -39.900 ;
        RECT -150.440 -40.400 -142.890 -39.920 ;
        RECT -150.440 -40.430 -143.080 -40.400 ;
        RECT 206.500 -40.430 207.010 -39.920 ;
        RECT 213.520 -40.350 214.030 -27.740 ;
        RECT 214.270 -33.760 215.730 -33.720 ;
        RECT 214.260 -33.930 215.730 -33.760 ;
        RECT 214.270 -33.970 215.730 -33.930 ;
        RECT 206.480 -40.640 207.010 -40.430 ;
        RECT 211.590 -40.640 214.030 -40.350 ;
        RECT 206.480 -41.120 214.030 -40.640 ;
        RECT 206.670 -41.150 214.030 -41.120 ;
        RECT -150.440 -42.190 -142.910 -41.640 ;
        RECT -152.130 -55.160 -150.650 -54.910 ;
        RECT -150.440 -55.100 -149.930 -42.190 ;
        RECT -143.580 -42.200 -142.910 -42.190 ;
        RECT -147.280 -43.090 -143.820 -42.650 ;
        RECT -149.210 -43.190 -143.820 -43.090 ;
        RECT -149.210 -43.260 -143.930 -43.190 ;
        RECT -149.210 -54.170 -149.040 -43.260 ;
        RECT -148.710 -43.670 -144.480 -43.650 ;
        RECT -148.730 -53.780 -144.400 -43.670 ;
        RECT -148.670 -53.830 -148.500 -53.780 ;
        RECT -144.100 -54.170 -143.930 -43.260 ;
        RECT -149.210 -54.340 -143.930 -54.170 ;
        RECT -144.170 -54.350 -143.930 -54.340 ;
        RECT -143.420 -55.100 -142.910 -42.200 ;
        RECT -150.440 -55.610 -142.910 -55.100 ;
        RECT -152.140 -61.630 -150.680 -61.590 ;
        RECT -152.140 -61.800 -150.670 -61.630 ;
        RECT -152.140 -61.840 -150.680 -61.800 ;
        RECT -150.440 -68.220 -149.930 -55.610 ;
        RECT -149.570 -56.400 -143.590 -56.170 ;
        RECT -149.480 -67.460 -143.830 -56.400 ;
        RECT -143.420 -65.970 -142.910 -55.610 ;
        RECT -143.430 -65.990 -142.910 -65.970 ;
        RECT 206.500 -42.910 214.030 -42.360 ;
        RECT 206.500 -42.920 207.170 -42.910 ;
        RECT 206.500 -55.820 207.010 -42.920 ;
        RECT 207.410 -43.810 210.870 -43.370 ;
        RECT 207.410 -43.910 212.800 -43.810 ;
        RECT 207.520 -43.980 212.800 -43.910 ;
        RECT 207.520 -54.890 207.690 -43.980 ;
        RECT 208.070 -44.390 212.300 -44.370 ;
        RECT 207.990 -54.500 212.320 -44.390 ;
        RECT 212.090 -54.550 212.260 -54.500 ;
        RECT 212.630 -54.890 212.800 -43.980 ;
        RECT 207.520 -55.060 212.800 -54.890 ;
        RECT 207.520 -55.070 207.760 -55.060 ;
        RECT 213.520 -55.820 214.030 -42.910 ;
        RECT 206.500 -56.330 214.030 -55.820 ;
        RECT 214.240 -55.880 215.720 -55.630 ;
        RECT -149.480 -67.470 -143.770 -67.460 ;
        RECT -149.560 -67.640 -143.770 -67.470 ;
        RECT -149.470 -67.650 -143.770 -67.640 ;
        RECT -144.000 -67.720 -143.830 -67.650 ;
        RECT -143.430 -67.770 -142.900 -65.990 ;
        RECT 206.500 -66.690 207.010 -56.330 ;
        RECT 207.180 -57.120 213.160 -56.890 ;
        RECT 206.500 -66.710 207.020 -66.690 ;
        RECT -143.420 -67.790 -142.900 -67.770 ;
        RECT -150.440 -68.510 -148.000 -68.220 ;
        RECT -143.420 -68.300 -142.910 -67.790 ;
        RECT -143.420 -68.510 -142.890 -68.300 ;
        RECT 206.490 -68.490 207.020 -66.710 ;
        RECT 207.420 -68.180 213.070 -57.120 ;
        RECT 207.360 -68.190 213.070 -68.180 ;
        RECT 207.360 -68.360 213.150 -68.190 ;
        RECT 207.360 -68.370 213.060 -68.360 ;
        RECT 207.420 -68.440 207.590 -68.370 ;
        RECT 206.490 -68.510 207.010 -68.490 ;
        RECT -150.440 -68.990 -142.890 -68.510 ;
        RECT -150.440 -69.020 -143.080 -68.990 ;
        RECT 206.500 -69.020 207.010 -68.510 ;
        RECT 213.520 -68.940 214.030 -56.330 ;
        RECT 214.270 -62.350 215.730 -62.310 ;
        RECT 214.260 -62.520 215.730 -62.350 ;
        RECT 214.270 -62.560 215.730 -62.520 ;
        RECT 206.480 -69.230 207.010 -69.020 ;
        RECT 211.590 -69.230 214.030 -68.940 ;
        RECT 206.480 -69.710 214.030 -69.230 ;
        RECT 206.670 -69.740 214.030 -69.710 ;
        RECT -150.440 -70.780 -142.910 -70.230 ;
        RECT -152.130 -83.750 -150.650 -83.500 ;
        RECT -150.440 -83.690 -149.930 -70.780 ;
        RECT -143.580 -70.790 -142.910 -70.780 ;
        RECT -147.280 -71.680 -143.820 -71.240 ;
        RECT -149.210 -71.780 -143.820 -71.680 ;
        RECT -149.210 -71.850 -143.930 -71.780 ;
        RECT -149.210 -82.760 -149.040 -71.850 ;
        RECT -148.710 -72.260 -144.480 -72.240 ;
        RECT -148.730 -82.370 -144.400 -72.260 ;
        RECT -148.670 -82.420 -148.500 -82.370 ;
        RECT -144.100 -82.760 -143.930 -71.850 ;
        RECT -149.210 -82.930 -143.930 -82.760 ;
        RECT -144.170 -82.940 -143.930 -82.930 ;
        RECT -143.420 -83.690 -142.910 -70.790 ;
        RECT -150.440 -84.200 -142.910 -83.690 ;
        RECT -152.140 -90.220 -150.680 -90.180 ;
        RECT -152.140 -90.390 -150.670 -90.220 ;
        RECT -152.140 -90.430 -150.680 -90.390 ;
        RECT -150.440 -96.810 -149.930 -84.200 ;
        RECT -149.570 -84.990 -143.590 -84.760 ;
        RECT -149.480 -96.050 -143.830 -84.990 ;
        RECT -143.420 -94.560 -142.910 -84.200 ;
        RECT -143.430 -94.580 -142.910 -94.560 ;
        RECT -149.480 -96.060 -143.770 -96.050 ;
        RECT -149.560 -96.230 -143.770 -96.060 ;
        RECT -149.470 -96.240 -143.770 -96.230 ;
        RECT -144.000 -96.310 -143.830 -96.240 ;
        RECT -143.430 -96.360 -142.900 -94.580 ;
        RECT -143.420 -96.380 -142.900 -96.360 ;
        RECT -150.440 -97.100 -148.000 -96.810 ;
        RECT -143.420 -96.890 -142.910 -96.380 ;
        RECT -143.420 -97.100 -142.890 -96.890 ;
        RECT -150.440 -97.580 -142.890 -97.100 ;
        RECT -150.440 -97.610 -143.080 -97.580 ;
        RECT -150.440 -99.370 -142.910 -98.820 ;
        RECT -152.130 -112.340 -150.650 -112.090 ;
        RECT -150.440 -112.280 -149.930 -99.370 ;
        RECT -143.580 -99.380 -142.910 -99.370 ;
        RECT -147.280 -100.270 -143.820 -99.830 ;
        RECT -149.210 -100.370 -143.820 -100.270 ;
        RECT -149.210 -100.440 -143.930 -100.370 ;
        RECT -149.210 -111.350 -149.040 -100.440 ;
        RECT -148.710 -100.850 -144.480 -100.830 ;
        RECT -148.730 -110.960 -144.400 -100.850 ;
        RECT -148.670 -111.010 -148.500 -110.960 ;
        RECT -144.100 -111.350 -143.930 -100.440 ;
        RECT -149.210 -111.520 -143.930 -111.350 ;
        RECT -144.170 -111.530 -143.930 -111.520 ;
        RECT -143.420 -112.280 -142.910 -99.380 ;
        RECT -150.440 -112.790 -142.910 -112.280 ;
        RECT -152.140 -118.810 -150.680 -118.770 ;
        RECT -152.140 -118.980 -150.670 -118.810 ;
        RECT -152.140 -119.020 -150.680 -118.980 ;
        RECT -150.440 -125.400 -149.930 -112.790 ;
        RECT -149.570 -113.580 -143.590 -113.350 ;
        RECT -149.480 -124.640 -143.830 -113.580 ;
        RECT -143.420 -123.150 -142.910 -112.790 ;
        RECT -143.430 -123.170 -142.910 -123.150 ;
        RECT -149.480 -124.650 -143.770 -124.640 ;
        RECT -149.560 -124.820 -143.770 -124.650 ;
        RECT -149.470 -124.830 -143.770 -124.820 ;
        RECT -144.000 -124.900 -143.830 -124.830 ;
        RECT -143.430 -124.950 -142.900 -123.170 ;
        RECT -143.420 -124.970 -142.900 -124.950 ;
        RECT -150.440 -125.690 -148.000 -125.400 ;
        RECT -143.420 -125.480 -142.910 -124.970 ;
        RECT -143.420 -125.690 -142.890 -125.480 ;
        RECT -150.440 -126.170 -142.890 -125.690 ;
        RECT -150.440 -126.200 -143.080 -126.170 ;
        RECT -150.440 -127.960 -142.910 -127.410 ;
        RECT -152.130 -140.930 -150.650 -140.680 ;
        RECT -150.440 -140.870 -149.930 -127.960 ;
        RECT -143.580 -127.970 -142.910 -127.960 ;
        RECT -147.280 -128.860 -143.820 -128.420 ;
        RECT -149.210 -128.960 -143.820 -128.860 ;
        RECT -149.210 -129.030 -143.930 -128.960 ;
        RECT -149.210 -139.940 -149.040 -129.030 ;
        RECT -148.710 -129.440 -144.480 -129.420 ;
        RECT -148.730 -139.550 -144.400 -129.440 ;
        RECT -148.670 -139.600 -148.500 -139.550 ;
        RECT -144.100 -139.940 -143.930 -129.030 ;
        RECT -149.210 -140.110 -143.930 -139.940 ;
        RECT -144.170 -140.120 -143.930 -140.110 ;
        RECT -143.420 -140.870 -142.910 -127.970 ;
        RECT -150.440 -141.380 -142.910 -140.870 ;
        RECT -152.140 -147.400 -150.680 -147.360 ;
        RECT -152.140 -147.570 -150.670 -147.400 ;
        RECT -152.140 -147.610 -150.680 -147.570 ;
        RECT -150.440 -153.990 -149.930 -141.380 ;
        RECT -149.570 -142.170 -143.590 -141.940 ;
        RECT -149.480 -153.230 -143.830 -142.170 ;
        RECT -143.420 -151.740 -142.910 -141.380 ;
        RECT -143.430 -151.760 -142.910 -151.740 ;
        RECT -149.480 -153.240 -143.770 -153.230 ;
        RECT -149.560 -153.410 -143.770 -153.240 ;
        RECT -149.470 -153.420 -143.770 -153.410 ;
        RECT -144.000 -153.490 -143.830 -153.420 ;
        RECT -143.430 -153.540 -142.900 -151.760 ;
        RECT -143.420 -153.560 -142.900 -153.540 ;
        RECT -150.440 -154.280 -148.000 -153.990 ;
        RECT -143.420 -154.070 -142.910 -153.560 ;
        RECT -143.420 -154.280 -142.890 -154.070 ;
        RECT -150.440 -154.760 -142.890 -154.280 ;
        RECT -150.440 -154.790 -143.080 -154.760 ;
        RECT -150.440 -156.550 -142.910 -156.000 ;
        RECT -152.130 -169.520 -150.650 -169.270 ;
        RECT -150.440 -169.460 -149.930 -156.550 ;
        RECT -143.580 -156.560 -142.910 -156.550 ;
        RECT -147.280 -157.450 -143.820 -157.010 ;
        RECT -149.210 -157.550 -143.820 -157.450 ;
        RECT -149.210 -157.620 -143.930 -157.550 ;
        RECT -149.210 -168.530 -149.040 -157.620 ;
        RECT -148.710 -158.030 -144.480 -158.010 ;
        RECT -148.730 -168.140 -144.400 -158.030 ;
        RECT -148.670 -168.190 -148.500 -168.140 ;
        RECT -144.100 -168.530 -143.930 -157.620 ;
        RECT -149.210 -168.700 -143.930 -168.530 ;
        RECT -144.170 -168.710 -143.930 -168.700 ;
        RECT -143.420 -169.460 -142.910 -156.560 ;
        RECT -150.440 -169.970 -142.910 -169.460 ;
        RECT -152.140 -175.990 -150.680 -175.950 ;
        RECT -152.140 -176.160 -150.670 -175.990 ;
        RECT -152.140 -176.200 -150.680 -176.160 ;
        RECT -150.440 -182.580 -149.930 -169.970 ;
        RECT -149.570 -170.760 -143.590 -170.530 ;
        RECT -149.480 -181.820 -143.830 -170.760 ;
        RECT -143.420 -180.330 -142.910 -169.970 ;
        RECT -143.430 -180.350 -142.910 -180.330 ;
        RECT -149.480 -181.830 -143.770 -181.820 ;
        RECT -149.560 -182.000 -143.770 -181.830 ;
        RECT -149.470 -182.010 -143.770 -182.000 ;
        RECT -144.000 -182.080 -143.830 -182.010 ;
        RECT -143.430 -182.130 -142.900 -180.350 ;
        RECT -143.420 -182.150 -142.900 -182.130 ;
        RECT -150.440 -182.870 -148.000 -182.580 ;
        RECT -143.420 -182.660 -142.910 -182.150 ;
        RECT -143.420 -182.870 -142.890 -182.660 ;
        RECT -150.440 -183.350 -142.890 -182.870 ;
        RECT -150.440 -183.380 -143.080 -183.350 ;
        RECT -150.440 -185.140 -142.910 -184.590 ;
        RECT -152.130 -198.110 -150.650 -197.860 ;
        RECT -150.440 -198.050 -149.930 -185.140 ;
        RECT -143.580 -185.150 -142.910 -185.140 ;
        RECT -147.280 -186.040 -143.820 -185.600 ;
        RECT -149.210 -186.140 -143.820 -186.040 ;
        RECT -149.210 -186.210 -143.930 -186.140 ;
        RECT -149.210 -197.120 -149.040 -186.210 ;
        RECT -148.710 -186.620 -144.480 -186.600 ;
        RECT -148.730 -196.730 -144.400 -186.620 ;
        RECT -148.670 -196.780 -148.500 -196.730 ;
        RECT -144.100 -197.120 -143.930 -186.210 ;
        RECT -149.210 -197.290 -143.930 -197.120 ;
        RECT -144.170 -197.300 -143.930 -197.290 ;
        RECT -143.420 -198.050 -142.910 -185.150 ;
        RECT -150.440 -198.560 -142.910 -198.050 ;
        RECT -152.140 -204.580 -150.680 -204.540 ;
        RECT -152.140 -204.750 -150.670 -204.580 ;
        RECT -152.140 -204.790 -150.680 -204.750 ;
        RECT -150.440 -211.170 -149.930 -198.560 ;
        RECT -149.570 -199.350 -143.590 -199.120 ;
        RECT -149.480 -210.410 -143.830 -199.350 ;
        RECT -143.420 -208.920 -142.910 -198.560 ;
        RECT -143.430 -208.940 -142.910 -208.920 ;
        RECT -149.480 -210.420 -143.770 -210.410 ;
        RECT -149.560 -210.590 -143.770 -210.420 ;
        RECT -149.470 -210.600 -143.770 -210.590 ;
        RECT -144.000 -210.670 -143.830 -210.600 ;
        RECT -143.430 -210.720 -142.900 -208.940 ;
        RECT -143.420 -210.740 -142.900 -210.720 ;
        RECT -150.440 -211.460 -148.000 -211.170 ;
        RECT -143.420 -211.250 -142.910 -210.740 ;
        RECT -143.420 -211.460 -142.890 -211.250 ;
        RECT -150.440 -211.940 -142.890 -211.460 ;
        RECT -150.440 -211.970 -143.080 -211.940 ;
        RECT -150.440 -213.730 -142.910 -213.180 ;
        RECT -152.130 -226.700 -150.650 -226.450 ;
        RECT -150.440 -226.640 -149.930 -213.730 ;
        RECT -143.580 -213.740 -142.910 -213.730 ;
        RECT -147.280 -214.630 -143.820 -214.190 ;
        RECT -149.210 -214.730 -143.820 -214.630 ;
        RECT -149.210 -214.800 -143.930 -214.730 ;
        RECT -149.210 -225.710 -149.040 -214.800 ;
        RECT -148.710 -215.210 -144.480 -215.190 ;
        RECT -148.730 -225.320 -144.400 -215.210 ;
        RECT -148.670 -225.370 -148.500 -225.320 ;
        RECT -144.100 -225.710 -143.930 -214.800 ;
        RECT -149.210 -225.880 -143.930 -225.710 ;
        RECT -144.170 -225.890 -143.930 -225.880 ;
        RECT -143.420 -226.640 -142.910 -213.740 ;
        RECT -150.440 -227.150 -142.910 -226.640 ;
        RECT -152.140 -233.170 -150.680 -233.130 ;
        RECT -152.140 -233.340 -150.670 -233.170 ;
        RECT -152.140 -233.380 -150.680 -233.340 ;
        RECT -150.440 -239.760 -149.930 -227.150 ;
        RECT -149.570 -227.940 -143.590 -227.710 ;
        RECT -149.480 -239.000 -143.830 -227.940 ;
        RECT -143.420 -237.510 -142.910 -227.150 ;
        RECT -143.430 -237.530 -142.910 -237.510 ;
        RECT -149.480 -239.010 -143.770 -239.000 ;
        RECT -149.560 -239.180 -143.770 -239.010 ;
        RECT -149.470 -239.190 -143.770 -239.180 ;
        RECT -144.000 -239.260 -143.830 -239.190 ;
        RECT -143.430 -239.310 -142.900 -237.530 ;
        RECT -143.420 -239.330 -142.900 -239.310 ;
        RECT -150.440 -240.050 -148.000 -239.760 ;
        RECT -143.420 -239.840 -142.910 -239.330 ;
        RECT -143.420 -240.050 -142.890 -239.840 ;
        RECT -150.440 -240.530 -142.890 -240.050 ;
        RECT -150.440 -240.560 -143.080 -240.530 ;
      LAYER mcon ;
        RECT -131.000 142.740 -130.830 142.910 ;
        RECT -131.000 142.380 -130.830 142.550 ;
        RECT -131.000 142.010 -130.830 142.180 ;
        RECT -124.320 143.060 -124.150 143.230 ;
        RECT -124.320 142.700 -124.150 142.870 ;
        RECT -124.320 142.340 -124.150 142.510 ;
        RECT -124.320 141.980 -124.150 142.150 ;
        RECT -102.410 142.740 -102.240 142.910 ;
        RECT -102.410 142.380 -102.240 142.550 ;
        RECT -102.410 142.010 -102.240 142.180 ;
        RECT -95.730 143.060 -95.560 143.230 ;
        RECT -95.730 142.700 -95.560 142.870 ;
        RECT -95.730 142.340 -95.560 142.510 ;
        RECT -95.730 141.980 -95.560 142.150 ;
        RECT -73.820 142.740 -73.650 142.910 ;
        RECT -73.820 142.380 -73.650 142.550 ;
        RECT -73.820 142.010 -73.650 142.180 ;
        RECT -67.140 143.060 -66.970 143.230 ;
        RECT -67.140 142.700 -66.970 142.870 ;
        RECT -67.140 142.340 -66.970 142.510 ;
        RECT -67.140 141.980 -66.970 142.150 ;
        RECT -31.870 142.910 -31.700 143.080 ;
        RECT -31.870 142.550 -31.700 142.720 ;
        RECT -31.870 142.190 -31.700 142.360 ;
        RECT -31.870 141.830 -31.700 142.000 ;
        RECT -25.120 142.740 -24.950 142.910 ;
        RECT -25.120 142.380 -24.950 142.550 ;
        RECT -25.120 142.020 -24.950 142.190 ;
        RECT 10.200 142.740 10.370 142.910 ;
        RECT 10.200 142.380 10.370 142.550 ;
        RECT 10.200 142.010 10.370 142.180 ;
        RECT 16.880 143.060 17.050 143.230 ;
        RECT 16.880 142.700 17.050 142.870 ;
        RECT 16.880 142.340 17.050 142.510 ;
        RECT 16.880 141.980 17.050 142.150 ;
        RECT 38.790 142.740 38.960 142.910 ;
        RECT 38.790 142.380 38.960 142.550 ;
        RECT 38.790 142.010 38.960 142.180 ;
        RECT 45.470 143.060 45.640 143.230 ;
        RECT 45.470 142.700 45.640 142.870 ;
        RECT 45.470 142.340 45.640 142.510 ;
        RECT 45.470 141.980 45.640 142.150 ;
        RECT 67.380 142.740 67.550 142.910 ;
        RECT 67.380 142.380 67.550 142.550 ;
        RECT 67.380 142.010 67.550 142.180 ;
        RECT 74.060 143.060 74.230 143.230 ;
        RECT 74.060 142.700 74.230 142.870 ;
        RECT 74.060 142.340 74.230 142.510 ;
        RECT 74.060 141.980 74.230 142.150 ;
        RECT 95.970 142.740 96.140 142.910 ;
        RECT 95.970 142.380 96.140 142.550 ;
        RECT 95.970 142.010 96.140 142.180 ;
        RECT 102.650 143.060 102.820 143.230 ;
        RECT 102.650 142.700 102.820 142.870 ;
        RECT 102.650 142.340 102.820 142.510 ;
        RECT 102.650 141.980 102.820 142.150 ;
        RECT 124.560 142.740 124.730 142.910 ;
        RECT 124.560 142.380 124.730 142.550 ;
        RECT 124.560 142.010 124.730 142.180 ;
        RECT 131.240 143.060 131.410 143.230 ;
        RECT 131.240 142.700 131.410 142.870 ;
        RECT 131.240 142.340 131.410 142.510 ;
        RECT 131.240 141.980 131.410 142.150 ;
        RECT 153.150 142.740 153.320 142.910 ;
        RECT 153.150 142.380 153.320 142.550 ;
        RECT 153.150 142.010 153.320 142.180 ;
        RECT 159.830 143.060 160.000 143.230 ;
        RECT 159.830 142.700 160.000 142.870 ;
        RECT 159.830 142.340 160.000 142.510 ;
        RECT 159.830 141.980 160.000 142.150 ;
        RECT 181.740 142.740 181.910 142.910 ;
        RECT 181.740 142.380 181.910 142.550 ;
        RECT 181.740 142.010 181.910 142.180 ;
        RECT 188.420 143.060 188.590 143.230 ;
        RECT 188.420 142.700 188.590 142.870 ;
        RECT 188.420 142.340 188.590 142.510 ;
        RECT 188.420 141.980 188.590 142.150 ;
        RECT -138.140 141.390 -136.280 141.400 ;
        RECT -138.140 141.220 -136.270 141.390 ;
        RECT -114.780 141.210 -111.620 141.390 ;
        RECT -138.100 139.130 -137.920 141.030 ;
        RECT -137.700 139.120 -137.520 141.030 ;
        RECT -136.510 140.090 -125.530 140.260 ;
        RECT -136.510 139.470 -125.530 139.640 ;
        RECT -136.500 138.850 -125.520 139.020 ;
        RECT -136.480 138.270 -125.500 138.440 ;
        RECT -136.470 137.680 -125.490 137.850 ;
        RECT -136.470 137.080 -125.490 137.250 ;
        RECT -136.520 136.480 -125.540 136.650 ;
        RECT -136.510 135.870 -125.530 136.040 ;
        RECT -136.520 135.270 -125.540 135.440 ;
        RECT -122.780 139.330 -113.330 139.500 ;
        RECT -122.790 138.580 -113.400 138.750 ;
        RECT -122.760 137.860 -113.360 138.030 ;
        RECT -122.750 137.200 -113.380 137.370 ;
        RECT -122.760 136.550 -113.310 136.720 ;
        RECT -122.750 135.910 -113.360 136.080 ;
        RECT -111.210 140.230 -111.010 141.160 ;
        RECT -112.280 134.990 -111.930 138.290 ;
        RECT -109.550 141.390 -107.690 141.400 ;
        RECT -109.550 141.220 -107.680 141.390 ;
        RECT -86.190 141.210 -83.030 141.390 ;
        RECT -109.510 139.130 -109.330 141.030 ;
        RECT -109.110 139.120 -108.930 141.030 ;
        RECT -107.920 140.090 -96.940 140.260 ;
        RECT -107.920 139.470 -96.940 139.640 ;
        RECT -107.910 138.850 -96.930 139.020 ;
        RECT -107.890 138.270 -96.910 138.440 ;
        RECT -107.880 137.680 -96.900 137.850 ;
        RECT -107.880 137.080 -96.900 137.250 ;
        RECT -107.930 136.480 -96.950 136.650 ;
        RECT -107.920 135.870 -96.940 136.040 ;
        RECT -107.930 135.270 -96.950 135.440 ;
        RECT -94.190 139.330 -84.740 139.500 ;
        RECT -94.200 138.580 -84.810 138.750 ;
        RECT -94.170 137.860 -84.770 138.030 ;
        RECT -94.160 137.200 -84.790 137.370 ;
        RECT -94.170 136.550 -84.720 136.720 ;
        RECT -94.160 135.910 -84.770 136.080 ;
        RECT -82.620 140.230 -82.420 141.160 ;
        RECT -83.690 134.990 -83.340 138.290 ;
        RECT -80.960 141.390 -79.100 141.400 ;
        RECT -80.960 141.220 -79.090 141.390 ;
        RECT -57.600 141.210 -54.440 141.390 ;
        RECT -80.920 139.130 -80.740 141.030 ;
        RECT -80.520 139.120 -80.340 141.030 ;
        RECT -79.330 140.090 -68.350 140.260 ;
        RECT -79.330 139.470 -68.350 139.640 ;
        RECT -79.320 138.850 -68.340 139.020 ;
        RECT -79.300 138.270 -68.320 138.440 ;
        RECT -79.290 137.680 -68.310 137.850 ;
        RECT -79.290 137.080 -68.310 137.250 ;
        RECT -79.340 136.480 -68.360 136.650 ;
        RECT -79.330 135.870 -68.350 136.040 ;
        RECT -79.340 135.270 -68.360 135.440 ;
        RECT -65.600 139.330 -56.150 139.500 ;
        RECT -65.610 138.580 -56.220 138.750 ;
        RECT -65.580 137.860 -56.180 138.030 ;
        RECT -65.570 137.200 -56.200 137.370 ;
        RECT -65.580 136.550 -56.130 136.720 ;
        RECT -65.570 135.910 -56.180 136.080 ;
        RECT -54.030 140.230 -53.830 141.160 ;
        RECT -55.100 134.990 -54.750 138.290 ;
        RECT -52.320 141.220 -28.420 141.390 ;
        RECT -19.540 141.220 1.630 141.390 ;
        RECT 3.060 141.390 4.920 141.400 ;
        RECT 3.060 141.220 4.930 141.390 ;
        RECT 26.420 141.210 29.580 141.390 ;
        RECT 3.100 139.130 3.280 141.030 ;
        RECT 3.500 139.120 3.680 141.030 ;
        RECT 4.690 140.090 15.670 140.260 ;
        RECT 4.690 139.470 15.670 139.640 ;
        RECT 4.700 138.850 15.680 139.020 ;
        RECT 4.720 138.270 15.700 138.440 ;
        RECT 4.730 137.680 15.710 137.850 ;
        RECT 4.730 137.080 15.710 137.250 ;
        RECT 4.680 136.480 15.660 136.650 ;
        RECT 4.690 135.870 15.670 136.040 ;
        RECT 4.680 135.270 15.660 135.440 ;
        RECT 18.420 139.330 27.870 139.500 ;
        RECT 18.410 138.580 27.800 138.750 ;
        RECT 18.440 137.860 27.840 138.030 ;
        RECT 18.450 137.200 27.820 137.370 ;
        RECT 18.440 136.550 27.890 136.720 ;
        RECT 18.450 135.910 27.840 136.080 ;
        RECT 29.990 140.230 30.190 141.160 ;
        RECT 28.920 134.990 29.270 138.290 ;
        RECT 31.650 141.390 33.510 141.400 ;
        RECT 31.650 141.220 33.520 141.390 ;
        RECT 55.010 141.210 58.170 141.390 ;
        RECT 31.690 139.130 31.870 141.030 ;
        RECT 32.090 139.120 32.270 141.030 ;
        RECT 33.280 140.090 44.260 140.260 ;
        RECT 33.280 139.470 44.260 139.640 ;
        RECT 33.290 138.850 44.270 139.020 ;
        RECT 33.310 138.270 44.290 138.440 ;
        RECT 33.320 137.680 44.300 137.850 ;
        RECT 33.320 137.080 44.300 137.250 ;
        RECT 33.270 136.480 44.250 136.650 ;
        RECT 33.280 135.870 44.260 136.040 ;
        RECT 33.270 135.270 44.250 135.440 ;
        RECT 47.010 139.330 56.460 139.500 ;
        RECT 47.000 138.580 56.390 138.750 ;
        RECT 47.030 137.860 56.430 138.030 ;
        RECT 47.040 137.200 56.410 137.370 ;
        RECT 47.030 136.550 56.480 136.720 ;
        RECT 47.040 135.910 56.430 136.080 ;
        RECT 58.580 140.230 58.780 141.160 ;
        RECT 57.510 134.990 57.860 138.290 ;
        RECT 60.240 141.390 62.100 141.400 ;
        RECT 60.240 141.220 62.110 141.390 ;
        RECT 83.600 141.210 86.760 141.390 ;
        RECT 60.280 139.130 60.460 141.030 ;
        RECT 60.680 139.120 60.860 141.030 ;
        RECT 61.870 140.090 72.850 140.260 ;
        RECT 61.870 139.470 72.850 139.640 ;
        RECT 61.880 138.850 72.860 139.020 ;
        RECT 61.900 138.270 72.880 138.440 ;
        RECT 61.910 137.680 72.890 137.850 ;
        RECT 61.910 137.080 72.890 137.250 ;
        RECT 61.860 136.480 72.840 136.650 ;
        RECT 61.870 135.870 72.850 136.040 ;
        RECT 61.860 135.270 72.840 135.440 ;
        RECT 75.600 139.330 85.050 139.500 ;
        RECT 75.590 138.580 84.980 138.750 ;
        RECT 75.620 137.860 85.020 138.030 ;
        RECT 75.630 137.200 85.000 137.370 ;
        RECT 75.620 136.550 85.070 136.720 ;
        RECT 75.630 135.910 85.020 136.080 ;
        RECT 87.170 140.230 87.370 141.160 ;
        RECT 86.100 134.990 86.450 138.290 ;
        RECT 88.830 141.390 90.690 141.400 ;
        RECT 88.830 141.220 90.700 141.390 ;
        RECT 112.190 141.210 115.350 141.390 ;
        RECT 88.870 139.130 89.050 141.030 ;
        RECT 89.270 139.120 89.450 141.030 ;
        RECT 90.460 140.090 101.440 140.260 ;
        RECT 90.460 139.470 101.440 139.640 ;
        RECT 90.470 138.850 101.450 139.020 ;
        RECT 90.490 138.270 101.470 138.440 ;
        RECT 90.500 137.680 101.480 137.850 ;
        RECT 90.500 137.080 101.480 137.250 ;
        RECT 90.450 136.480 101.430 136.650 ;
        RECT 90.460 135.870 101.440 136.040 ;
        RECT 90.450 135.270 101.430 135.440 ;
        RECT 104.190 139.330 113.640 139.500 ;
        RECT 104.180 138.580 113.570 138.750 ;
        RECT 104.210 137.860 113.610 138.030 ;
        RECT 104.220 137.200 113.590 137.370 ;
        RECT 104.210 136.550 113.660 136.720 ;
        RECT 104.220 135.910 113.610 136.080 ;
        RECT 115.760 140.230 115.960 141.160 ;
        RECT 114.690 134.990 115.040 138.290 ;
        RECT 117.420 141.390 119.280 141.400 ;
        RECT 117.420 141.220 119.290 141.390 ;
        RECT 140.780 141.210 143.940 141.390 ;
        RECT 117.460 139.130 117.640 141.030 ;
        RECT 117.860 139.120 118.040 141.030 ;
        RECT 119.050 140.090 130.030 140.260 ;
        RECT 119.050 139.470 130.030 139.640 ;
        RECT 119.060 138.850 130.040 139.020 ;
        RECT 119.080 138.270 130.060 138.440 ;
        RECT 119.090 137.680 130.070 137.850 ;
        RECT 119.090 137.080 130.070 137.250 ;
        RECT 119.040 136.480 130.020 136.650 ;
        RECT 119.050 135.870 130.030 136.040 ;
        RECT 119.040 135.270 130.020 135.440 ;
        RECT 132.780 139.330 142.230 139.500 ;
        RECT 132.770 138.580 142.160 138.750 ;
        RECT 132.800 137.860 142.200 138.030 ;
        RECT 132.810 137.200 142.180 137.370 ;
        RECT 132.800 136.550 142.250 136.720 ;
        RECT 132.810 135.910 142.200 136.080 ;
        RECT 144.350 140.230 144.550 141.160 ;
        RECT 143.280 134.990 143.630 138.290 ;
        RECT 146.010 141.390 147.870 141.400 ;
        RECT 146.010 141.220 147.880 141.390 ;
        RECT 169.370 141.210 172.530 141.390 ;
        RECT 146.050 139.130 146.230 141.030 ;
        RECT 146.450 139.120 146.630 141.030 ;
        RECT 147.640 140.090 158.620 140.260 ;
        RECT 147.640 139.470 158.620 139.640 ;
        RECT 147.650 138.850 158.630 139.020 ;
        RECT 147.670 138.270 158.650 138.440 ;
        RECT 147.680 137.680 158.660 137.850 ;
        RECT 147.680 137.080 158.660 137.250 ;
        RECT 147.630 136.480 158.610 136.650 ;
        RECT 147.640 135.870 158.620 136.040 ;
        RECT 147.630 135.270 158.610 135.440 ;
        RECT 161.370 139.330 170.820 139.500 ;
        RECT 161.360 138.580 170.750 138.750 ;
        RECT 161.390 137.860 170.790 138.030 ;
        RECT 161.400 137.200 170.770 137.370 ;
        RECT 161.390 136.550 170.840 136.720 ;
        RECT 161.400 135.910 170.790 136.080 ;
        RECT 172.940 140.230 173.140 141.160 ;
        RECT 171.870 134.990 172.220 138.290 ;
        RECT 174.600 141.390 176.460 141.400 ;
        RECT 174.600 141.220 176.470 141.390 ;
        RECT 197.960 141.210 201.120 141.390 ;
        RECT 174.640 139.130 174.820 141.030 ;
        RECT 175.040 139.120 175.220 141.030 ;
        RECT 176.230 140.090 187.210 140.260 ;
        RECT 176.230 139.470 187.210 139.640 ;
        RECT 176.240 138.850 187.220 139.020 ;
        RECT 176.260 138.270 187.240 138.440 ;
        RECT 176.270 137.680 187.250 137.850 ;
        RECT 176.270 137.080 187.250 137.250 ;
        RECT 176.220 136.480 187.200 136.650 ;
        RECT 176.230 135.870 187.210 136.040 ;
        RECT 176.220 135.270 187.200 135.440 ;
        RECT 189.960 139.330 199.410 139.500 ;
        RECT 189.950 138.580 199.340 138.750 ;
        RECT 189.980 137.860 199.380 138.030 ;
        RECT 189.990 137.200 199.360 137.370 ;
        RECT 189.980 136.550 199.430 136.720 ;
        RECT 189.990 135.910 199.380 136.080 ;
        RECT 201.530 140.230 201.730 141.160 ;
        RECT 200.460 134.990 200.810 138.290 ;
        RECT -25.850 133.260 -25.680 133.430 ;
        RECT -25.480 133.260 -25.310 133.430 ;
        RECT -25.120 133.260 -24.950 133.430 ;
        RECT -24.760 133.260 -24.590 133.430 ;
        RECT -24.400 133.260 -24.220 133.430 ;
        RECT -24.030 133.260 -23.860 133.430 ;
        RECT -150.040 129.530 -149.110 129.730 ;
        RECT -150.270 125.960 -150.090 129.120 ;
        RECT -147.170 128.460 -143.870 128.810 ;
        RECT -152.110 116.420 -151.940 116.590 ;
        RECT -151.750 116.420 -151.580 116.590 ;
        RECT -151.390 116.420 -151.220 116.590 ;
        RECT -151.030 116.420 -150.860 116.590 ;
        RECT -148.380 117.960 -148.210 127.410 ;
        RECT -147.630 117.950 -147.460 127.340 ;
        RECT -146.910 117.980 -146.740 127.380 ;
        RECT -146.250 117.990 -146.080 127.360 ;
        RECT -145.600 117.980 -145.430 127.430 ;
        RECT -144.960 117.990 -144.790 127.380 ;
        RECT 212.700 128.810 213.630 129.010 ;
        RECT -23.230 127.310 -23.060 127.480 ;
        RECT -20.360 127.520 -20.190 127.690 ;
        RECT -21.820 127.310 -21.650 127.480 ;
        RECT -5.020 127.340 -4.850 127.510 ;
        RECT -20.360 126.730 -20.190 126.900 ;
        RECT -5.020 126.650 -4.850 126.820 ;
        RECT 0.840 127.250 1.010 127.420 ;
        RECT 0.840 126.800 1.010 126.970 ;
        RECT 5.540 127.200 5.710 127.370 ;
        RECT 5.540 126.750 5.710 126.920 ;
        RECT -23.230 126.460 -23.060 126.630 ;
        RECT -22.510 126.450 -22.340 126.620 ;
        RECT -21.820 126.460 -21.650 126.630 ;
        RECT -23.050 126.050 -22.880 126.220 ;
        RECT -21.990 126.050 -21.820 126.220 ;
        RECT -23.230 125.640 -23.060 125.810 ;
        RECT -22.510 125.610 -22.340 125.780 ;
        RECT -21.820 125.640 -21.650 125.810 ;
        RECT -7.120 125.710 -6.950 125.880 ;
        RECT -5.760 125.790 -5.590 125.960 ;
        RECT -5.070 125.780 -4.900 125.950 ;
        RECT -20.360 125.300 -20.190 125.470 ;
        RECT -23.230 124.800 -23.060 124.970 ;
        RECT -21.820 124.800 -21.650 124.970 ;
        RECT -21.090 124.540 -20.920 124.710 ;
        RECT -21.100 124.020 -20.930 124.190 ;
        RECT -20.350 123.900 -20.180 124.070 ;
        RECT -23.230 123.680 -23.060 123.850 ;
        RECT -21.820 123.680 -21.650 123.850 ;
        RECT -22.530 122.810 -22.360 122.980 ;
        RECT -21.100 122.830 -20.930 123.000 ;
        RECT -18.340 122.480 -18.170 122.650 ;
        RECT -23.320 122.230 -23.150 122.400 ;
        RECT -22.390 122.230 -22.220 122.400 ;
        RECT -21.690 122.230 -21.520 122.400 ;
        RECT -20.950 122.230 -20.780 122.400 ;
        RECT -20.240 122.220 -20.070 122.390 ;
        RECT -5.020 124.540 -4.850 124.710 ;
        RECT -5.020 123.850 -4.850 124.020 ;
        RECT 0.840 124.260 1.010 124.430 ;
        RECT 0.840 123.810 1.010 123.980 ;
        RECT 0.840 123.250 1.010 123.420 ;
        RECT -5.020 122.990 -4.850 123.160 ;
        RECT 0.840 122.800 1.010 122.970 ;
        RECT -5.020 122.300 -4.850 122.470 ;
        RECT 4.760 123.740 4.930 123.910 ;
        RECT -7.840 122.050 -7.670 122.220 ;
        RECT 2.020 122.070 2.190 122.240 ;
        RECT -7.830 117.690 -7.400 118.430 ;
        RECT 13.270 116.270 13.480 116.480 ;
        RECT 17.010 116.290 17.180 116.460 ;
        RECT -151.790 109.740 -151.620 109.910 ;
        RECT -151.430 109.740 -151.260 109.910 ;
        RECT -151.060 109.740 -150.890 109.910 ;
        RECT -150.270 104.460 -150.100 104.470 ;
        RECT -150.280 102.600 -150.100 104.460 ;
        RECT -149.140 104.230 -148.970 115.210 ;
        RECT -148.520 104.230 -148.350 115.210 ;
        RECT -147.900 104.240 -147.730 115.220 ;
        RECT -147.320 104.260 -147.150 115.240 ;
        RECT -146.730 104.270 -146.560 115.250 ;
        RECT -146.130 104.270 -145.960 115.250 ;
        RECT -145.530 104.220 -145.360 115.200 ;
        RECT -144.920 104.230 -144.750 115.210 ;
        RECT -144.320 104.220 -144.150 115.200 ;
        RECT 11.800 115.900 11.970 116.070 ;
        RECT 18.050 116.330 18.220 116.500 ;
        RECT 19.090 115.990 19.260 116.160 ;
        RECT 19.090 115.630 19.260 115.800 ;
        RECT 207.460 127.740 210.760 128.090 ;
        RECT 208.380 117.270 208.550 126.660 ;
        RECT 209.020 117.260 209.190 126.710 ;
        RECT 209.670 117.270 209.840 126.640 ;
        RECT 210.330 117.260 210.500 126.660 ;
        RECT 211.050 117.230 211.220 126.620 ;
        RECT 211.800 117.240 211.970 126.690 ;
        RECT 213.680 125.240 213.860 128.400 ;
        RECT 13.270 114.520 13.480 114.730 ;
        RECT 17.010 114.540 17.180 114.710 ;
        RECT 11.800 114.150 11.970 114.320 ;
        RECT 18.050 114.580 18.220 114.750 ;
        RECT 40.460 114.530 40.720 115.350 ;
        RECT 52.410 114.560 52.730 115.350 ;
        RECT 214.450 115.700 214.620 115.870 ;
        RECT 214.810 115.700 214.980 115.870 ;
        RECT 215.170 115.700 215.340 115.870 ;
        RECT 215.530 115.700 215.700 115.870 ;
        RECT 19.090 114.240 19.260 114.410 ;
        RECT 19.090 113.880 19.260 114.050 ;
        RECT -9.950 112.910 -9.780 113.080 ;
        RECT -8.860 112.920 -8.690 113.090 ;
        RECT 13.270 112.770 13.480 112.980 ;
        RECT 17.010 112.790 17.180 112.960 ;
        RECT -10.380 112.410 -10.210 112.580 ;
        RECT -8.010 112.350 -7.840 112.520 ;
        RECT 11.800 112.400 11.970 112.570 ;
        RECT -9.940 111.920 -9.770 112.090 ;
        RECT -8.850 111.930 -8.680 112.100 ;
        RECT 18.050 112.830 18.220 113.000 ;
        RECT 50.570 112.780 50.740 112.950 ;
        RECT 19.090 112.490 19.260 112.660 ;
        RECT 28.520 112.470 28.700 112.640 ;
        RECT 28.950 112.450 29.120 112.620 ;
        RECT 19.090 112.130 19.260 112.300 ;
        RECT 26.710 112.170 26.880 112.340 ;
        RECT -10.400 111.490 -10.230 111.660 ;
        RECT 27.060 111.330 27.240 111.520 ;
        RECT -9.940 110.930 -9.770 111.100 ;
        RECT -8.850 110.940 -8.680 111.110 ;
        RECT 13.270 111.020 13.480 111.230 ;
        RECT 17.010 111.040 17.180 111.210 ;
        RECT -10.420 110.500 -10.250 110.670 ;
        RECT 11.800 110.650 11.970 110.820 ;
        RECT 18.050 111.080 18.220 111.250 ;
        RECT 19.090 110.740 19.260 110.910 ;
        RECT 19.090 110.380 19.260 110.550 ;
        RECT 29.420 111.890 29.590 112.060 ;
        RECT 48.670 112.170 48.840 112.340 ;
        RECT 31.660 111.590 31.830 111.760 ;
        RECT 41.830 111.590 42.000 111.760 ;
        RECT 31.660 111.140 31.830 111.310 ;
        RECT 28.140 110.770 28.310 110.940 ;
        RECT 37.110 110.990 37.380 111.260 ;
        RECT 38.170 110.990 38.440 111.260 ;
        RECT 41.830 111.140 42.000 111.310 ;
        RECT 47.000 111.340 47.170 111.510 ;
        RECT 28.950 110.460 29.120 110.630 ;
        RECT -10.130 110.000 -9.960 110.170 ;
        RECT -8.830 109.900 -8.660 110.070 ;
        RECT -10.130 109.010 -9.960 109.180 ;
        RECT -8.830 108.910 -8.660 109.080 ;
        RECT 11.800 108.950 11.970 109.120 ;
        RECT 20.250 109.470 20.420 109.640 ;
        RECT 19.090 109.220 19.260 109.390 ;
        RECT 21.090 109.350 21.260 109.520 ;
        RECT 21.840 109.350 22.010 109.520 ;
        RECT -8.420 108.430 -8.250 108.600 ;
        RECT 13.270 108.540 13.480 108.750 ;
        RECT 17.010 108.560 17.180 108.730 ;
        RECT 19.090 108.860 19.260 109.030 ;
        RECT 18.050 108.520 18.220 108.690 ;
        RECT 24.820 109.020 24.990 109.190 ;
        RECT 20.530 108.720 20.700 108.890 ;
        RECT 25.220 109.470 25.390 109.640 ;
        RECT 51.540 112.530 51.710 112.700 ;
        RECT 52.520 112.210 52.690 112.380 ;
        RECT 53.790 112.550 53.960 112.720 ;
        RECT 50.720 111.950 50.890 112.120 ;
        RECT 48.310 111.330 48.490 111.520 ;
        RECT 49.600 111.430 49.770 111.600 ;
        RECT 34.790 109.880 34.960 110.050 ;
        RECT 40.590 109.880 40.760 110.050 ;
        RECT 25.220 109.110 25.390 109.280 ;
        RECT 27.060 108.530 27.240 108.720 ;
        RECT -10.130 108.020 -9.960 108.190 ;
        RECT -8.830 107.920 -8.660 108.090 ;
        RECT 11.800 107.200 11.970 107.370 ;
        RECT 19.090 107.470 19.260 107.640 ;
        RECT 20.530 107.660 20.700 107.830 ;
        RECT 29.420 109.570 29.590 109.740 ;
        RECT 28.960 109.390 29.130 109.560 ;
        RECT 28.130 109.080 28.300 109.250 ;
        RECT 37.110 109.260 37.380 109.530 ;
        RECT 38.170 109.260 38.440 109.530 ;
        RECT 31.660 108.640 31.830 108.810 ;
        RECT 31.660 108.190 31.830 108.360 ;
        RECT 41.830 108.640 42.000 108.810 ;
        RECT 47.000 108.580 47.170 108.750 ;
        RECT 41.830 108.190 42.000 108.360 ;
        RECT 29.410 107.990 29.580 108.160 ;
        RECT 13.270 106.790 13.480 107.000 ;
        RECT 17.010 106.810 17.180 106.980 ;
        RECT 24.820 107.360 24.990 107.530 ;
        RECT 19.090 107.110 19.260 107.280 ;
        RECT 18.050 106.770 18.220 106.940 ;
        RECT 21.090 107.030 21.260 107.200 ;
        RECT 21.840 107.030 22.010 107.200 ;
        RECT 23.840 107.040 24.010 107.210 ;
        RECT 25.220 107.630 25.390 107.800 ;
        RECT 26.710 107.710 26.880 107.880 ;
        RECT 25.220 107.270 25.390 107.440 ;
        RECT 48.310 108.530 48.490 108.720 ;
        RECT 48.670 107.710 48.840 107.880 ;
        RECT 28.520 107.410 28.700 107.580 ;
        RECT 28.980 107.480 29.150 107.650 ;
        RECT 51.490 111.880 51.660 112.050 ;
        RECT 51.490 111.040 51.660 111.210 ;
        RECT 53.180 111.240 53.350 111.410 ;
        RECT 52.520 110.710 52.690 110.880 ;
        RECT 51.540 110.390 51.710 110.560 ;
        RECT 50.330 110.150 50.500 110.320 ;
        RECT 53.840 110.330 54.010 110.500 ;
        RECT 79.250 110.080 79.420 110.250 ;
        RECT 80.210 109.940 80.380 110.110 ;
        RECT 80.820 110.080 80.990 110.250 ;
        RECT 81.340 109.950 81.510 110.120 ;
        RECT 50.760 109.350 50.930 109.520 ;
        RECT 51.540 109.530 51.710 109.700 ;
        RECT 53.830 109.610 54.000 109.780 ;
        RECT 52.520 109.210 52.690 109.380 ;
        RECT 51.490 108.880 51.660 109.050 ;
        RECT 77.800 109.300 77.970 109.470 ;
        RECT 78.300 109.330 78.470 109.500 ;
        RECT 81.800 109.330 81.970 109.500 ;
        RECT 53.180 108.650 53.350 108.820 ;
        RECT 51.490 108.040 51.660 108.210 ;
        RECT 78.300 108.250 78.470 108.420 ;
        RECT 81.800 108.250 81.970 108.420 ;
        RECT 52.520 107.710 52.690 107.880 ;
        RECT 51.540 107.390 51.710 107.560 ;
        RECT 53.750 107.360 53.920 107.530 ;
        RECT 79.250 107.500 79.420 107.670 ;
        RECT 80.210 107.640 80.380 107.810 ;
        RECT 80.820 107.500 80.990 107.670 ;
        RECT 81.340 107.630 81.510 107.800 ;
        RECT 20.250 106.270 20.420 106.440 ;
        RECT 11.800 105.450 11.970 105.620 ;
        RECT 21.090 106.150 21.260 106.320 ;
        RECT 21.840 106.150 22.010 106.320 ;
        RECT 19.090 105.720 19.260 105.890 ;
        RECT 13.270 105.040 13.480 105.250 ;
        RECT 17.010 105.060 17.180 105.230 ;
        RECT 19.090 105.360 19.260 105.530 ;
        RECT 24.820 105.820 24.990 105.990 ;
        RECT 20.530 105.520 20.700 105.690 ;
        RECT 25.220 106.270 25.390 106.440 ;
        RECT 28.530 106.440 28.710 106.610 ;
        RECT 25.220 105.910 25.390 106.080 ;
        RECT 26.720 106.140 26.890 106.310 ;
        RECT 27.070 105.300 27.250 105.490 ;
        RECT 18.050 105.020 18.220 105.190 ;
        RECT 20.530 104.460 20.700 104.630 ;
        RECT -149.910 103.040 -148.000 103.220 ;
        RECT 11.800 103.700 11.970 103.870 ;
        RECT 24.820 104.160 24.990 104.330 ;
        RECT 19.090 103.970 19.260 104.140 ;
        RECT 13.270 103.290 13.480 103.500 ;
        RECT 17.010 103.310 17.180 103.480 ;
        RECT 19.090 103.610 19.260 103.780 ;
        RECT 21.090 103.830 21.260 104.000 ;
        RECT 21.840 103.830 22.010 104.000 ;
        RECT 23.840 103.840 24.010 104.010 ;
        RECT 25.220 104.430 25.390 104.600 ;
        RECT 50.570 106.750 50.740 106.920 ;
        RECT 48.670 106.140 48.840 106.310 ;
        RECT 33.560 105.560 33.730 105.730 ;
        RECT 35.650 105.720 35.820 105.890 ;
        RECT 28.390 105.310 28.560 105.480 ;
        RECT 41.830 105.560 42.000 105.730 ;
        RECT 33.560 105.110 33.730 105.280 ;
        RECT 37.120 104.960 37.390 105.230 ;
        RECT 38.170 104.960 38.440 105.230 ;
        RECT 41.830 105.110 42.000 105.280 ;
        RECT 47.000 105.310 47.170 105.480 ;
        RECT 25.220 104.070 25.390 104.240 ;
        RECT 34.800 104.210 34.970 104.380 ;
        RECT 34.800 103.850 34.970 104.020 ;
        RECT 18.050 103.270 18.220 103.440 ;
        RECT -149.910 102.640 -148.010 102.820 ;
        RECT 27.070 102.500 27.250 102.690 ;
        RECT 34.810 103.490 34.980 103.660 ;
        RECT 40.590 104.210 40.760 104.380 ;
        RECT 51.540 106.500 51.710 106.670 ;
        RECT 52.520 106.180 52.690 106.350 ;
        RECT 53.790 106.520 53.960 106.690 ;
        RECT 79.250 106.880 79.420 107.050 ;
        RECT 80.210 106.740 80.380 106.910 ;
        RECT 80.820 106.880 80.990 107.050 ;
        RECT 81.340 106.750 81.510 106.920 ;
        RECT 50.720 105.920 50.890 106.090 ;
        RECT 48.310 105.300 48.490 105.490 ;
        RECT 49.600 105.400 49.770 105.570 ;
        RECT 40.590 103.850 40.760 104.020 ;
        RECT 37.120 103.230 37.390 103.500 ;
        RECT 38.170 103.230 38.440 103.500 ;
        RECT 40.590 103.490 40.760 103.660 ;
        RECT 28.390 102.550 28.560 102.720 ;
        RECT 33.560 102.610 33.730 102.780 ;
        RECT 33.560 102.160 33.730 102.330 ;
        RECT 41.830 102.610 42.000 102.780 ;
        RECT 47.000 102.550 47.170 102.720 ;
        RECT 35.680 102.030 35.850 102.200 ;
        RECT 41.830 102.160 42.000 102.330 ;
        RECT 48.310 102.500 48.490 102.690 ;
        RECT 26.720 101.680 26.890 101.850 ;
        RECT 28.530 101.380 28.710 101.550 ;
        RECT -150.040 100.940 -149.110 101.140 ;
        RECT 48.670 101.680 48.840 101.850 ;
        RECT 51.490 105.850 51.660 106.020 ;
        RECT 77.800 106.100 77.970 106.270 ;
        RECT 78.300 106.130 78.470 106.300 ;
        RECT 81.800 106.130 81.970 106.300 ;
        RECT 51.490 105.010 51.660 105.180 ;
        RECT 53.180 105.210 53.350 105.380 ;
        RECT 52.520 104.680 52.690 104.850 ;
        RECT 78.300 105.050 78.470 105.220 ;
        RECT 81.800 105.050 81.970 105.220 ;
        RECT 51.540 104.360 51.710 104.530 ;
        RECT 50.330 104.120 50.500 104.290 ;
        RECT 53.840 104.300 54.010 104.470 ;
        RECT 79.250 104.300 79.420 104.470 ;
        RECT 80.210 104.440 80.380 104.610 ;
        RECT 80.820 104.300 80.990 104.470 ;
        RECT 81.340 104.430 81.510 104.600 ;
        RECT 50.760 103.320 50.930 103.490 ;
        RECT 51.540 103.500 51.710 103.670 ;
        RECT 53.830 103.580 54.000 103.750 ;
        RECT 52.520 103.180 52.690 103.350 ;
        RECT 51.490 102.850 51.660 103.020 ;
        RECT 207.740 103.500 207.910 114.480 ;
        RECT 208.340 103.510 208.510 114.490 ;
        RECT 208.950 103.500 209.120 114.480 ;
        RECT 209.550 103.550 209.720 114.530 ;
        RECT 210.150 103.550 210.320 114.530 ;
        RECT 210.740 103.540 210.910 114.520 ;
        RECT 211.320 103.520 211.490 114.500 ;
        RECT 211.940 103.510 212.110 114.490 ;
        RECT 212.560 103.510 212.730 114.490 ;
        RECT 214.480 109.020 214.650 109.190 ;
        RECT 214.850 109.020 215.020 109.190 ;
        RECT 215.210 109.020 215.380 109.190 ;
        RECT 53.180 102.620 53.350 102.790 ;
        RECT 213.690 103.740 213.860 103.750 ;
        RECT 211.590 102.320 213.500 102.500 ;
        RECT 51.490 102.010 51.660 102.180 ;
        RECT 52.520 101.680 52.690 101.850 ;
        RECT 211.600 101.920 213.500 102.100 ;
        RECT 213.690 101.880 213.870 103.740 ;
        RECT 51.540 101.360 51.710 101.530 ;
        RECT 53.750 101.330 53.920 101.500 ;
        RECT -150.270 97.370 -150.090 100.530 ;
        RECT -147.170 99.870 -143.870 100.220 ;
        RECT -152.110 87.830 -151.940 88.000 ;
        RECT -151.750 87.830 -151.580 88.000 ;
        RECT -151.390 87.830 -151.220 88.000 ;
        RECT -151.030 87.830 -150.860 88.000 ;
        RECT -148.380 89.370 -148.210 98.820 ;
        RECT -147.630 89.360 -147.460 98.750 ;
        RECT -146.910 89.390 -146.740 98.790 ;
        RECT -146.250 89.400 -146.080 98.770 ;
        RECT -145.600 89.390 -145.430 98.840 ;
        RECT -144.960 89.400 -144.790 98.790 ;
        RECT 212.700 100.220 213.630 100.420 ;
        RECT 11.800 98.820 11.970 98.990 ;
        RECT 19.090 99.090 19.260 99.260 ;
        RECT 13.270 98.410 13.480 98.620 ;
        RECT 17.010 98.430 17.180 98.600 ;
        RECT 19.090 98.730 19.260 98.900 ;
        RECT 20.230 99.000 20.400 99.170 ;
        RECT 21.070 98.880 21.240 99.050 ;
        RECT 21.820 98.880 21.990 99.050 ;
        RECT 18.050 98.390 18.220 98.560 ;
        RECT 24.800 98.550 24.970 98.720 ;
        RECT 20.510 98.250 20.680 98.420 ;
        RECT 25.200 99.000 25.370 99.170 ;
        RECT 25.200 98.640 25.370 98.810 ;
        RECT 29.940 98.820 30.110 98.990 ;
        RECT 45.430 98.820 45.600 98.990 ;
        RECT 28.130 98.560 28.300 98.730 ;
        RECT 28.860 98.530 29.030 98.700 ;
        RECT 46.510 98.530 46.680 98.700 ;
        RECT 29.940 98.270 30.110 98.440 ;
        RECT 45.430 98.270 45.600 98.440 ;
        RECT 47.240 98.560 47.410 98.730 ;
        RECT 30.850 97.870 31.020 98.040 ;
        RECT 11.800 97.070 11.970 97.240 ;
        RECT 19.090 97.340 19.260 97.510 ;
        RECT 13.270 96.660 13.480 96.870 ;
        RECT 17.010 96.680 17.180 96.850 ;
        RECT 19.090 96.980 19.260 97.150 ;
        RECT 20.510 97.190 20.680 97.360 ;
        RECT 24.800 96.890 24.970 97.060 ;
        RECT 18.050 96.640 18.220 96.810 ;
        RECT 21.070 96.560 21.240 96.730 ;
        RECT 21.820 96.560 21.990 96.730 ;
        RECT 23.820 96.570 23.990 96.740 ;
        RECT 25.200 97.160 25.370 97.330 ;
        RECT 28.130 97.000 28.300 97.170 ;
        RECT 34.790 97.880 34.960 98.050 ;
        RECT 40.580 97.880 40.750 98.050 ;
        RECT 44.520 97.870 44.690 98.040 ;
        RECT 29.940 97.290 30.110 97.460 ;
        RECT 45.430 97.290 45.600 97.460 ;
        RECT 28.860 97.030 29.030 97.200 ;
        RECT 46.510 97.030 46.680 97.200 ;
        RECT 47.240 97.000 47.410 97.170 ;
        RECT 25.200 96.800 25.370 96.970 ;
        RECT 29.940 96.740 30.110 96.910 ;
        RECT 30.850 96.280 31.020 96.450 ;
        RECT 34.780 96.420 34.950 96.590 ;
        RECT 45.430 96.740 45.600 96.910 ;
        RECT 11.800 95.320 11.970 95.490 ;
        RECT 20.230 95.800 20.400 95.970 ;
        RECT 19.090 95.590 19.260 95.760 ;
        RECT 13.270 94.910 13.480 95.120 ;
        RECT 17.010 94.930 17.180 95.100 ;
        RECT 21.070 95.680 21.240 95.850 ;
        RECT 21.820 95.680 21.990 95.850 ;
        RECT 19.090 95.230 19.260 95.400 ;
        RECT 18.050 94.890 18.220 95.060 ;
        RECT 24.800 95.350 24.970 95.520 ;
        RECT 20.510 95.050 20.680 95.220 ;
        RECT 25.200 95.800 25.370 95.970 ;
        RECT 30.850 95.920 31.020 96.090 ;
        RECT 33.060 96.030 33.330 96.300 ;
        RECT 34.780 96.060 34.950 96.230 ;
        RECT 25.200 95.440 25.370 95.610 ;
        RECT 29.940 95.580 30.110 95.750 ;
        RECT 37.090 96.100 37.360 96.370 ;
        RECT 38.180 96.100 38.450 96.370 ;
        RECT 40.590 96.420 40.760 96.590 ;
        RECT 40.590 96.060 40.760 96.230 ;
        RECT 42.210 96.030 42.480 96.300 ;
        RECT 44.520 96.280 44.690 96.450 ;
        RECT 46.880 96.160 47.060 96.330 ;
        RECT 44.520 95.920 44.690 96.090 ;
        RECT 45.430 95.580 45.600 95.750 ;
        RECT 28.130 95.320 28.300 95.490 ;
        RECT 28.860 95.290 29.030 95.460 ;
        RECT 46.510 95.290 46.680 95.460 ;
        RECT 29.940 95.030 30.110 95.200 ;
        RECT 45.430 95.030 45.600 95.200 ;
        RECT 47.240 95.320 47.410 95.490 ;
        RECT 11.800 93.570 11.970 93.740 ;
        RECT 19.090 93.840 19.260 94.010 ;
        RECT 20.510 93.990 20.680 94.160 ;
        RECT 13.270 93.160 13.480 93.370 ;
        RECT 17.010 93.180 17.180 93.350 ;
        RECT 24.800 93.690 24.970 93.860 ;
        RECT 19.090 93.480 19.260 93.650 ;
        RECT 18.050 93.140 18.220 93.310 ;
        RECT 21.070 93.360 21.240 93.530 ;
        RECT 21.820 93.360 21.990 93.530 ;
        RECT 23.820 93.370 23.990 93.540 ;
        RECT 25.200 93.960 25.370 94.130 ;
        RECT 25.200 93.600 25.370 93.770 ;
        RECT 28.130 93.770 28.300 93.940 ;
        RECT 29.940 94.060 30.110 94.230 ;
        RECT 45.430 94.060 45.600 94.230 ;
        RECT 28.860 93.800 29.030 93.970 ;
        RECT 46.510 93.800 46.680 93.970 ;
        RECT 47.240 93.770 47.410 93.940 ;
        RECT 29.940 93.510 30.110 93.680 ;
        RECT 45.430 93.510 45.600 93.680 ;
        RECT -11.010 90.340 -10.840 90.510 ;
        RECT -10.360 90.340 -10.190 90.510 ;
        RECT -12.230 89.900 -12.060 90.070 ;
        RECT -11.530 89.900 -11.360 90.070 ;
        RECT -12.680 88.240 -12.510 88.410 ;
        RECT 11.760 89.760 11.930 89.930 ;
        RECT 19.050 90.030 19.220 90.200 ;
        RECT -9.850 89.520 -9.680 89.690 ;
        RECT 13.230 89.350 13.440 89.560 ;
        RECT 16.970 89.370 17.140 89.540 ;
        RECT 19.050 89.670 19.220 89.840 ;
        RECT 20.260 89.730 20.430 89.900 ;
        RECT 18.010 89.330 18.180 89.500 ;
        RECT 21.100 89.610 21.270 89.780 ;
        RECT 21.850 89.610 22.020 89.780 ;
        RECT 24.830 89.280 25.000 89.450 ;
        RECT 20.540 88.980 20.710 89.150 ;
        RECT 25.230 89.730 25.400 89.900 ;
        RECT 25.230 89.370 25.400 89.540 ;
        RECT 29.970 89.490 30.140 89.660 ;
        RECT 28.160 89.230 28.330 89.400 ;
        RECT 28.890 89.200 29.060 89.370 ;
        RECT 38.650 89.200 38.820 89.370 ;
        RECT 29.970 88.940 30.140 89.110 ;
        RECT -9.680 88.040 -9.510 88.210 ;
        RECT 11.760 88.010 11.930 88.180 ;
        RECT 31.010 88.480 31.180 88.650 ;
        RECT 19.050 88.280 19.220 88.450 ;
        RECT -151.790 81.150 -151.620 81.320 ;
        RECT -151.430 81.150 -151.260 81.320 ;
        RECT -151.060 81.150 -150.890 81.320 ;
        RECT -150.270 75.870 -150.100 75.880 ;
        RECT -150.280 74.010 -150.100 75.870 ;
        RECT -149.140 75.640 -148.970 86.620 ;
        RECT -148.520 75.640 -148.350 86.620 ;
        RECT -147.900 75.650 -147.730 86.630 ;
        RECT -147.320 75.670 -147.150 86.650 ;
        RECT -146.730 75.680 -146.560 86.660 ;
        RECT -146.130 75.680 -145.960 86.660 ;
        RECT -145.530 75.630 -145.360 86.610 ;
        RECT -144.920 75.640 -144.750 86.620 ;
        RECT -144.320 75.630 -144.150 86.610 ;
        RECT -12.200 86.020 -12.030 86.190 ;
        RECT -11.510 86.010 -11.340 86.180 ;
        RECT -11.030 85.240 -10.860 85.410 ;
        RECT -9.670 87.500 -9.500 87.670 ;
        RECT 13.230 87.600 13.440 87.810 ;
        RECT 16.970 87.620 17.140 87.790 ;
        RECT 19.050 87.920 19.220 88.090 ;
        RECT 18.010 87.580 18.180 87.750 ;
        RECT 20.540 87.920 20.710 88.090 ;
        RECT 24.830 87.620 25.000 87.790 ;
        RECT 21.100 87.290 21.270 87.460 ;
        RECT 21.850 87.290 22.020 87.460 ;
        RECT 23.850 87.300 24.020 87.470 ;
        RECT 25.230 87.890 25.400 88.060 ;
        RECT 25.230 87.530 25.400 87.700 ;
        RECT 28.160 87.690 28.330 87.860 ;
        RECT 29.970 87.980 30.140 88.150 ;
        RECT 35.030 88.510 35.200 88.680 ;
        RECT 38.800 88.520 38.970 88.690 ;
        RECT 40.950 88.640 41.120 88.810 ;
        RECT 39.690 88.070 39.860 88.240 ;
        RECT 28.890 87.720 29.060 87.890 ;
        RECT 29.970 87.430 30.140 87.600 ;
        RECT 38.800 87.620 38.970 87.790 ;
        RECT 31.000 87.280 31.170 87.450 ;
        RECT -9.860 86.540 -9.690 86.710 ;
        RECT 11.760 86.260 11.930 86.430 ;
        RECT 35.020 87.220 35.190 87.390 ;
        RECT 40.950 87.500 41.120 87.670 ;
        RECT 19.050 86.530 19.220 86.700 ;
        RECT 13.230 85.850 13.440 86.060 ;
        RECT 16.970 85.870 17.140 86.040 ;
        RECT 19.050 86.170 19.220 86.340 ;
        RECT 20.260 86.530 20.430 86.700 ;
        RECT 21.100 86.410 21.270 86.580 ;
        RECT 21.850 86.410 22.020 86.580 ;
        RECT 18.010 85.830 18.180 86.000 ;
        RECT 24.830 86.080 25.000 86.250 ;
        RECT 20.540 85.780 20.710 85.950 ;
        RECT 25.230 86.530 25.400 86.700 ;
        RECT 31.000 86.620 31.170 86.790 ;
        RECT 25.230 86.170 25.400 86.340 ;
        RECT 29.970 86.250 30.140 86.420 ;
        RECT 33.090 86.660 33.360 86.930 ;
        RECT 35.020 86.580 35.190 86.750 ;
        RECT 37.120 86.730 37.390 87.000 ;
        RECT 38.650 86.940 38.820 87.110 ;
        RECT 207.460 99.150 210.760 99.500 ;
        RECT 208.380 88.680 208.550 98.070 ;
        RECT 209.020 88.670 209.190 98.120 ;
        RECT 209.670 88.680 209.840 98.050 ;
        RECT 210.330 88.670 210.500 98.070 ;
        RECT 211.050 88.640 211.220 98.030 ;
        RECT 211.800 88.650 211.970 98.100 ;
        RECT 213.680 96.650 213.860 99.810 ;
        RECT 214.450 87.110 214.620 87.280 ;
        RECT 214.810 87.110 214.980 87.280 ;
        RECT 215.170 87.110 215.340 87.280 ;
        RECT 215.530 87.110 215.700 87.280 ;
        RECT 38.650 86.430 38.820 86.600 ;
        RECT 28.160 85.990 28.330 86.160 ;
        RECT 28.890 85.960 29.060 86.130 ;
        RECT 29.970 85.700 30.140 85.870 ;
        RECT 38.800 85.750 38.970 85.920 ;
        RECT 40.950 85.870 41.120 86.040 ;
        RECT -10.320 85.180 -10.150 85.350 ;
        RECT 39.690 85.300 39.860 85.470 ;
        RECT 11.760 84.510 11.930 84.680 ;
        RECT 19.050 84.780 19.220 84.950 ;
        RECT 13.230 84.100 13.440 84.310 ;
        RECT 16.970 84.120 17.140 84.290 ;
        RECT 20.540 84.720 20.710 84.890 ;
        RECT 19.050 84.420 19.220 84.590 ;
        RECT 24.830 84.420 25.000 84.590 ;
        RECT 18.010 84.080 18.180 84.250 ;
        RECT 21.100 84.090 21.270 84.260 ;
        RECT 21.850 84.090 22.020 84.260 ;
        RECT 23.850 84.100 24.020 84.270 ;
        RECT 25.230 84.690 25.400 84.860 ;
        RECT 27.210 84.790 27.380 84.960 ;
        RECT 25.230 84.330 25.400 84.500 ;
        RECT 28.160 84.440 28.330 84.610 ;
        RECT 29.970 84.730 30.140 84.900 ;
        RECT 38.800 84.850 38.970 85.020 ;
        RECT 28.890 84.470 29.060 84.640 ;
        RECT 40.950 84.730 41.120 84.900 ;
        RECT 29.970 84.180 30.140 84.350 ;
        RECT 38.650 84.170 38.820 84.340 ;
        RECT 27.260 83.830 27.430 84.000 ;
        RECT 19.920 81.830 20.090 82.000 ;
        RECT -11.000 80.160 -10.830 80.330 ;
        RECT -14.310 79.720 -14.140 79.890 ;
        RECT -13.210 79.730 -13.040 79.900 ;
        RECT -13.760 79.050 -13.590 79.220 ;
        RECT -13.760 77.680 -13.590 77.850 ;
        RECT -14.310 76.950 -14.140 77.120 ;
        RECT -14.320 75.610 -14.150 75.780 ;
        RECT -149.910 74.450 -148.000 74.630 ;
        RECT -12.120 79.730 -11.950 79.900 ;
        RECT -12.660 79.050 -12.490 79.220 ;
        RECT -12.660 77.680 -12.490 77.850 ;
        RECT -13.210 76.950 -13.040 77.120 ;
        RECT -13.210 75.600 -13.040 75.770 ;
        RECT -13.760 74.910 -13.590 75.080 ;
        RECT -3.680 79.980 -3.510 80.320 ;
        RECT -3.310 79.980 -3.140 80.320 ;
        RECT -10.990 79.690 -10.820 79.860 ;
        RECT -11.560 79.050 -11.390 79.220 ;
        RECT -10.870 79.030 -10.700 79.200 ;
        RECT 21.010 81.830 21.180 82.000 ;
        RECT 20.470 81.150 20.640 81.320 ;
        RECT 20.470 79.780 20.640 79.950 ;
        RECT 19.910 79.050 20.080 79.220 ;
        RECT -10.870 78.340 -10.700 78.510 ;
        RECT -11.560 77.680 -11.390 77.850 ;
        RECT 19.910 77.680 20.080 77.850 ;
        RECT -12.120 76.950 -11.950 77.120 ;
        RECT -12.120 75.580 -11.950 75.750 ;
        RECT -12.660 74.900 -12.490 75.070 ;
        RECT 19.340 77.040 19.510 77.210 ;
        RECT 22.110 81.820 22.280 81.990 ;
        RECT 21.560 81.130 21.730 81.300 ;
        RECT 21.560 79.780 21.730 79.950 ;
        RECT 21.010 79.050 21.180 79.220 ;
        RECT 21.010 77.680 21.180 77.850 ;
        RECT 20.470 77.000 20.640 77.170 ;
        RECT 23.230 82.000 23.400 82.170 ;
        RECT 23.230 81.640 23.400 81.810 ;
        RECT 23.840 82.000 24.010 82.170 ;
        RECT 23.840 81.640 24.010 81.810 ;
        RECT 24.960 81.820 25.130 81.990 ;
        RECT 22.670 81.120 22.840 81.290 ;
        RECT 24.400 81.120 24.570 81.290 ;
        RECT 22.660 79.780 22.830 79.950 ;
        RECT 24.410 79.780 24.580 79.950 ;
        RECT 22.110 79.050 22.280 79.220 ;
        RECT 22.110 77.680 22.280 77.850 ;
        RECT 21.560 77.000 21.730 77.170 ;
        RECT 26.060 81.830 26.230 82.000 ;
        RECT 25.510 81.130 25.680 81.300 ;
        RECT 25.510 79.780 25.680 79.950 ;
        RECT 24.960 79.050 25.130 79.220 ;
        RECT 24.960 77.680 25.130 77.850 ;
        RECT 22.660 77.010 22.830 77.180 ;
        RECT 24.410 77.010 24.580 77.180 ;
        RECT 27.150 81.830 27.320 82.000 ;
        RECT 29.730 81.860 29.900 82.030 ;
        RECT 26.600 81.150 26.770 81.320 ;
        RECT 26.600 79.780 26.770 79.950 ;
        RECT 26.060 79.050 26.230 79.220 ;
        RECT 26.060 77.680 26.230 77.850 ;
        RECT 25.510 77.000 25.680 77.170 ;
        RECT 30.820 81.860 30.990 82.030 ;
        RECT 30.280 81.180 30.450 81.350 ;
        RECT 30.280 79.810 30.450 79.980 ;
        RECT 27.160 79.050 27.330 79.220 ;
        RECT 29.720 79.080 29.890 79.250 ;
        RECT 27.160 77.680 27.330 77.850 ;
        RECT 29.720 77.710 29.890 77.880 ;
        RECT 26.600 77.000 26.770 77.170 ;
        RECT 27.730 77.040 27.900 77.210 ;
        RECT 19.350 76.570 19.520 76.740 ;
        RECT 27.720 76.570 27.890 76.740 ;
        RECT 29.150 77.070 29.320 77.240 ;
        RECT 31.920 81.850 32.090 82.020 ;
        RECT 31.370 81.160 31.540 81.330 ;
        RECT 31.370 79.810 31.540 79.980 ;
        RECT 30.820 79.080 30.990 79.250 ;
        RECT 30.820 77.710 30.990 77.880 ;
        RECT 30.280 77.030 30.450 77.200 ;
        RECT 33.040 82.030 33.210 82.200 ;
        RECT 33.040 81.670 33.210 81.840 ;
        RECT 33.650 82.030 33.820 82.200 ;
        RECT 33.650 81.670 33.820 81.840 ;
        RECT 34.770 81.850 34.940 82.020 ;
        RECT 32.480 81.150 32.650 81.320 ;
        RECT 34.210 81.150 34.380 81.320 ;
        RECT 32.470 79.810 32.640 79.980 ;
        RECT 34.220 79.810 34.390 79.980 ;
        RECT 31.920 79.080 32.090 79.250 ;
        RECT 31.920 77.710 32.090 77.880 ;
        RECT 31.370 77.030 31.540 77.200 ;
        RECT 35.870 81.860 36.040 82.030 ;
        RECT 35.320 81.160 35.490 81.330 ;
        RECT 35.320 79.810 35.490 79.980 ;
        RECT 34.770 79.080 34.940 79.250 ;
        RECT 34.770 77.710 34.940 77.880 ;
        RECT 32.470 77.040 32.640 77.210 ;
        RECT 34.220 77.040 34.390 77.210 ;
        RECT 36.960 81.860 37.130 82.030 ;
        RECT 36.410 81.180 36.580 81.350 ;
        RECT 36.410 79.810 36.580 79.980 ;
        RECT 35.870 79.080 36.040 79.250 ;
        RECT 35.870 77.710 36.040 77.880 ;
        RECT 35.320 77.030 35.490 77.200 ;
        RECT 40.510 81.840 40.680 82.010 ;
        RECT 39.950 81.140 40.120 81.310 ;
        RECT 39.960 79.800 40.130 79.970 ;
        RECT 36.970 79.080 37.140 79.250 ;
        RECT 36.970 77.710 37.140 77.880 ;
        RECT 36.410 77.030 36.580 77.200 ;
        RECT 41.610 81.850 41.780 82.020 ;
        RECT 41.060 81.150 41.230 81.320 ;
        RECT 41.060 79.800 41.230 79.970 ;
        RECT 40.510 79.070 40.680 79.240 ;
        RECT 40.510 77.700 40.680 77.870 ;
        RECT 37.540 77.070 37.710 77.240 ;
        RECT 29.160 76.600 29.330 76.770 ;
        RECT 39.960 77.030 40.130 77.200 ;
        RECT 42.700 81.850 42.870 82.020 ;
        RECT 42.150 81.170 42.320 81.340 ;
        RECT 42.150 79.800 42.320 79.970 ;
        RECT 41.610 79.070 41.780 79.240 ;
        RECT 41.610 77.700 41.780 77.870 ;
        RECT 41.060 77.020 41.230 77.190 ;
        RECT 42.710 79.070 42.880 79.240 ;
        RECT 43.400 78.770 43.570 78.940 ;
        RECT 43.400 78.410 43.570 78.580 ;
        RECT 42.710 77.700 42.880 77.870 ;
        RECT 42.150 77.020 42.320 77.190 ;
        RECT 43.280 77.060 43.450 77.230 ;
        RECT 37.530 76.600 37.700 76.770 ;
        RECT 43.270 76.590 43.440 76.760 ;
        RECT -11.570 74.900 -11.400 75.070 ;
        RECT -149.910 74.050 -148.010 74.230 ;
        RECT 74.520 74.060 74.690 74.230 ;
        RECT 80.040 73.320 80.210 73.490 ;
        RECT -150.040 72.350 -149.110 72.550 ;
        RECT -10.960 72.610 -10.790 72.780 ;
        RECT -14.270 72.170 -14.100 72.340 ;
        RECT -150.270 68.780 -150.090 71.940 ;
        RECT -147.170 71.280 -143.870 71.630 ;
        RECT -152.110 59.240 -151.940 59.410 ;
        RECT -151.750 59.240 -151.580 59.410 ;
        RECT -151.390 59.240 -151.220 59.410 ;
        RECT -151.030 59.240 -150.860 59.410 ;
        RECT -148.380 60.780 -148.210 70.230 ;
        RECT -147.630 60.770 -147.460 70.160 ;
        RECT -146.910 60.800 -146.740 70.200 ;
        RECT -146.250 60.810 -146.080 70.180 ;
        RECT -145.600 60.800 -145.430 70.250 ;
        RECT -144.960 60.810 -144.790 70.200 ;
        RECT -13.170 72.180 -13.000 72.350 ;
        RECT -13.720 71.500 -13.550 71.670 ;
        RECT -13.720 70.130 -13.550 70.300 ;
        RECT -14.270 69.400 -14.100 69.570 ;
        RECT -14.280 68.060 -14.110 68.230 ;
        RECT -14.840 67.540 -14.670 67.710 ;
        RECT -12.080 72.180 -11.910 72.350 ;
        RECT -12.620 71.500 -12.450 71.670 ;
        RECT -12.620 70.130 -12.450 70.300 ;
        RECT -13.170 69.400 -13.000 69.570 ;
        RECT -13.170 68.050 -13.000 68.220 ;
        RECT -13.720 67.360 -13.550 67.530 ;
        RECT 74.520 72.450 74.690 72.620 ;
        RECT -10.950 72.140 -10.780 72.310 ;
        RECT 80.040 72.650 80.210 72.820 ;
        RECT -11.520 71.500 -11.350 71.670 ;
        RECT -11.520 70.130 -11.350 70.300 ;
        RECT -12.080 69.400 -11.910 69.570 ;
        RECT -12.080 68.030 -11.910 68.200 ;
        RECT -12.620 67.350 -12.450 67.520 ;
        RECT -9.490 68.010 -9.320 71.530 ;
        RECT -9.130 68.010 -8.960 71.530 ;
        RECT -8.770 68.010 -8.600 71.530 ;
        RECT -8.080 68.010 -7.910 71.530 ;
        RECT -7.720 68.010 -7.550 71.530 ;
        RECT -7.360 68.010 -7.190 71.530 ;
        RECT 74.520 70.850 74.690 71.020 ;
        RECT 74.520 69.230 74.690 69.400 ;
        RECT 77.050 68.070 77.220 68.240 ;
        RECT 74.520 67.630 74.690 67.800 ;
        RECT -11.530 67.350 -11.360 67.520 ;
        RECT 74.520 66.010 74.690 66.180 ;
        RECT 74.520 64.410 74.690 64.580 ;
        RECT 74.520 62.790 74.690 62.960 ;
        RECT 80.880 60.800 81.050 75.750 ;
        RECT 207.740 74.910 207.910 85.890 ;
        RECT 208.340 74.920 208.510 85.900 ;
        RECT 208.950 74.910 209.120 85.890 ;
        RECT 209.550 74.960 209.720 85.940 ;
        RECT 210.150 74.960 210.320 85.940 ;
        RECT 210.740 74.950 210.910 85.930 ;
        RECT 211.320 74.930 211.490 85.910 ;
        RECT 211.940 74.920 212.110 85.900 ;
        RECT 212.560 74.920 212.730 85.900 ;
        RECT 214.480 80.430 214.650 80.600 ;
        RECT 214.850 80.430 215.020 80.600 ;
        RECT 215.210 80.430 215.380 80.600 ;
        RECT 213.690 75.150 213.860 75.160 ;
        RECT 211.590 73.730 213.500 73.910 ;
        RECT 211.600 73.330 213.500 73.510 ;
        RECT 213.690 73.290 213.870 75.150 ;
        RECT 212.700 71.630 213.630 71.830 ;
        RECT -151.790 52.560 -151.620 52.730 ;
        RECT -151.430 52.560 -151.260 52.730 ;
        RECT -151.060 52.560 -150.890 52.730 ;
        RECT -150.270 47.280 -150.100 47.290 ;
        RECT -150.280 45.420 -150.100 47.280 ;
        RECT -149.140 47.050 -148.970 58.030 ;
        RECT -148.520 47.050 -148.350 58.030 ;
        RECT -147.900 47.060 -147.730 58.040 ;
        RECT -147.320 47.080 -147.150 58.060 ;
        RECT -146.730 47.090 -146.560 58.070 ;
        RECT -146.130 47.090 -145.960 58.070 ;
        RECT -145.530 47.040 -145.360 58.020 ;
        RECT -144.920 47.050 -144.750 58.030 ;
        RECT -144.320 47.040 -144.150 58.020 ;
        RECT 207.460 70.560 210.760 70.910 ;
        RECT 208.380 60.090 208.550 69.480 ;
        RECT 209.020 60.080 209.190 69.530 ;
        RECT 209.670 60.090 209.840 69.460 ;
        RECT 210.330 60.080 210.500 69.480 ;
        RECT 211.050 60.050 211.220 69.440 ;
        RECT 211.800 60.060 211.970 69.510 ;
        RECT 213.680 68.060 213.860 71.220 ;
        RECT 214.450 58.520 214.620 58.690 ;
        RECT 214.810 58.520 214.980 58.690 ;
        RECT 215.170 58.520 215.340 58.690 ;
        RECT 215.530 58.520 215.700 58.690 ;
        RECT -149.910 45.860 -148.000 46.040 ;
        RECT 207.740 46.320 207.910 57.300 ;
        RECT 208.340 46.330 208.510 57.310 ;
        RECT 208.950 46.320 209.120 57.300 ;
        RECT 209.550 46.370 209.720 57.350 ;
        RECT 210.150 46.370 210.320 57.350 ;
        RECT 210.740 46.360 210.910 57.340 ;
        RECT 211.320 46.340 211.490 57.320 ;
        RECT 211.940 46.330 212.110 57.310 ;
        RECT 212.560 46.330 212.730 57.310 ;
        RECT 214.480 51.840 214.650 52.010 ;
        RECT 214.850 51.840 215.020 52.010 ;
        RECT 215.210 51.840 215.380 52.010 ;
        RECT -149.910 45.460 -148.010 45.640 ;
        RECT 213.690 46.560 213.860 46.570 ;
        RECT 211.590 45.140 213.500 45.320 ;
        RECT 211.600 44.740 213.500 44.920 ;
        RECT 213.690 44.700 213.870 46.560 ;
        RECT -150.040 43.760 -149.110 43.960 ;
        RECT -150.270 40.190 -150.090 43.350 ;
        RECT -147.170 42.690 -143.870 43.040 ;
        RECT -152.110 30.650 -151.940 30.820 ;
        RECT -151.750 30.650 -151.580 30.820 ;
        RECT -151.390 30.650 -151.220 30.820 ;
        RECT -151.030 30.650 -150.860 30.820 ;
        RECT -148.380 32.190 -148.210 41.640 ;
        RECT -147.630 32.180 -147.460 41.570 ;
        RECT -146.910 32.210 -146.740 41.610 ;
        RECT -146.250 32.220 -146.080 41.590 ;
        RECT -145.600 32.210 -145.430 41.660 ;
        RECT -144.960 32.220 -144.790 41.610 ;
        RECT -151.790 23.970 -151.620 24.140 ;
        RECT -151.430 23.970 -151.260 24.140 ;
        RECT -151.060 23.970 -150.890 24.140 ;
        RECT -150.270 18.690 -150.100 18.700 ;
        RECT -150.280 16.830 -150.100 18.690 ;
        RECT -149.140 18.460 -148.970 29.440 ;
        RECT -148.520 18.460 -148.350 29.440 ;
        RECT -147.900 18.470 -147.730 29.450 ;
        RECT -147.320 18.490 -147.150 29.470 ;
        RECT -146.730 18.500 -146.560 29.480 ;
        RECT -146.130 18.500 -145.960 29.480 ;
        RECT -145.530 18.450 -145.360 29.430 ;
        RECT -144.920 18.460 -144.750 29.440 ;
        RECT -144.320 18.450 -144.150 29.430 ;
        RECT 212.700 43.040 213.630 43.240 ;
        RECT 207.460 41.970 210.760 42.320 ;
        RECT 208.380 31.500 208.550 40.890 ;
        RECT 209.020 31.490 209.190 40.940 ;
        RECT 209.670 31.500 209.840 40.870 ;
        RECT 210.330 31.490 210.500 40.890 ;
        RECT 211.050 31.460 211.220 40.850 ;
        RECT 211.800 31.470 211.970 40.920 ;
        RECT 213.680 39.470 213.860 42.630 ;
        RECT 214.450 29.930 214.620 30.100 ;
        RECT 214.810 29.930 214.980 30.100 ;
        RECT 215.170 29.930 215.340 30.100 ;
        RECT 215.530 29.930 215.700 30.100 ;
        RECT -149.910 17.270 -148.000 17.450 ;
        RECT 207.740 17.730 207.910 28.710 ;
        RECT 208.340 17.740 208.510 28.720 ;
        RECT 208.950 17.730 209.120 28.710 ;
        RECT 209.550 17.780 209.720 28.760 ;
        RECT 210.150 17.780 210.320 28.760 ;
        RECT 210.740 17.770 210.910 28.750 ;
        RECT 211.320 17.750 211.490 28.730 ;
        RECT 211.940 17.740 212.110 28.720 ;
        RECT 212.560 17.740 212.730 28.720 ;
        RECT 214.480 23.250 214.650 23.420 ;
        RECT 214.850 23.250 215.020 23.420 ;
        RECT 215.210 23.250 215.380 23.420 ;
        RECT -149.910 16.870 -148.010 17.050 ;
        RECT 213.690 17.970 213.860 17.980 ;
        RECT 211.590 16.550 213.500 16.730 ;
        RECT 211.600 16.150 213.500 16.330 ;
        RECT 213.690 16.110 213.870 17.970 ;
        RECT -150.040 15.170 -149.110 15.370 ;
        RECT -150.270 11.600 -150.090 14.760 ;
        RECT -147.170 14.100 -143.870 14.450 ;
        RECT -152.110 2.060 -151.940 2.230 ;
        RECT -151.750 2.060 -151.580 2.230 ;
        RECT -151.390 2.060 -151.220 2.230 ;
        RECT -151.030 2.060 -150.860 2.230 ;
        RECT -148.380 3.600 -148.210 13.050 ;
        RECT -147.630 3.590 -147.460 12.980 ;
        RECT -146.910 3.620 -146.740 13.020 ;
        RECT -146.250 3.630 -146.080 13.000 ;
        RECT -145.600 3.620 -145.430 13.070 ;
        RECT -144.960 3.630 -144.790 13.020 ;
        RECT -151.790 -4.620 -151.620 -4.450 ;
        RECT -151.430 -4.620 -151.260 -4.450 ;
        RECT -151.060 -4.620 -150.890 -4.450 ;
        RECT -150.270 -9.900 -150.100 -9.890 ;
        RECT -150.280 -11.760 -150.100 -9.900 ;
        RECT -149.140 -10.130 -148.970 0.850 ;
        RECT -148.520 -10.130 -148.350 0.850 ;
        RECT -147.900 -10.120 -147.730 0.860 ;
        RECT -147.320 -10.100 -147.150 0.880 ;
        RECT -146.730 -10.090 -146.560 0.890 ;
        RECT -146.130 -10.090 -145.960 0.890 ;
        RECT -145.530 -10.140 -145.360 0.840 ;
        RECT -144.920 -10.130 -144.750 0.850 ;
        RECT -144.320 -10.140 -144.150 0.840 ;
        RECT 212.700 14.450 213.630 14.650 ;
        RECT 207.460 13.380 210.760 13.730 ;
        RECT 208.380 2.910 208.550 12.300 ;
        RECT 209.020 2.900 209.190 12.350 ;
        RECT 209.670 2.910 209.840 12.280 ;
        RECT 210.330 2.900 210.500 12.300 ;
        RECT 211.050 2.870 211.220 12.260 ;
        RECT 211.800 2.880 211.970 12.330 ;
        RECT 213.680 10.880 213.860 14.040 ;
        RECT 214.450 1.340 214.620 1.510 ;
        RECT 214.810 1.340 214.980 1.510 ;
        RECT 215.170 1.340 215.340 1.510 ;
        RECT 215.530 1.340 215.700 1.510 ;
        RECT -149.910 -11.320 -148.000 -11.140 ;
        RECT 207.740 -10.860 207.910 0.120 ;
        RECT 208.340 -10.850 208.510 0.130 ;
        RECT 208.950 -10.860 209.120 0.120 ;
        RECT 209.550 -10.810 209.720 0.170 ;
        RECT 210.150 -10.810 210.320 0.170 ;
        RECT 210.740 -10.820 210.910 0.160 ;
        RECT 211.320 -10.840 211.490 0.140 ;
        RECT 211.940 -10.850 212.110 0.130 ;
        RECT 212.560 -10.850 212.730 0.130 ;
        RECT 214.480 -5.340 214.650 -5.170 ;
        RECT 214.850 -5.340 215.020 -5.170 ;
        RECT 215.210 -5.340 215.380 -5.170 ;
        RECT -149.910 -11.720 -148.010 -11.540 ;
        RECT 213.690 -10.620 213.860 -10.610 ;
        RECT 211.590 -12.040 213.500 -11.860 ;
        RECT 211.600 -12.440 213.500 -12.260 ;
        RECT 213.690 -12.480 213.870 -10.620 ;
        RECT -150.040 -13.420 -149.110 -13.220 ;
        RECT -150.270 -16.990 -150.090 -13.830 ;
        RECT -147.170 -14.490 -143.870 -14.140 ;
        RECT -152.110 -26.530 -151.940 -26.360 ;
        RECT -151.750 -26.530 -151.580 -26.360 ;
        RECT -151.390 -26.530 -151.220 -26.360 ;
        RECT -151.030 -26.530 -150.860 -26.360 ;
        RECT -148.380 -24.990 -148.210 -15.540 ;
        RECT -147.630 -25.000 -147.460 -15.610 ;
        RECT -146.910 -24.970 -146.740 -15.570 ;
        RECT -146.250 -24.960 -146.080 -15.590 ;
        RECT -145.600 -24.970 -145.430 -15.520 ;
        RECT -144.960 -24.960 -144.790 -15.570 ;
        RECT -151.790 -33.210 -151.620 -33.040 ;
        RECT -151.430 -33.210 -151.260 -33.040 ;
        RECT -151.060 -33.210 -150.890 -33.040 ;
        RECT -150.270 -38.490 -150.100 -38.480 ;
        RECT -150.280 -40.350 -150.100 -38.490 ;
        RECT -149.140 -38.720 -148.970 -27.740 ;
        RECT -148.520 -38.720 -148.350 -27.740 ;
        RECT -147.900 -38.710 -147.730 -27.730 ;
        RECT -147.320 -38.690 -147.150 -27.710 ;
        RECT -146.730 -38.680 -146.560 -27.700 ;
        RECT -146.130 -38.680 -145.960 -27.700 ;
        RECT -145.530 -38.730 -145.360 -27.750 ;
        RECT -144.920 -38.720 -144.750 -27.740 ;
        RECT -144.320 -38.730 -144.150 -27.750 ;
        RECT 212.700 -14.140 213.630 -13.940 ;
        RECT 207.460 -15.210 210.760 -14.860 ;
        RECT 208.380 -25.680 208.550 -16.290 ;
        RECT 209.020 -25.690 209.190 -16.240 ;
        RECT 209.670 -25.680 209.840 -16.310 ;
        RECT 210.330 -25.690 210.500 -16.290 ;
        RECT 211.050 -25.720 211.220 -16.330 ;
        RECT 211.800 -25.710 211.970 -16.260 ;
        RECT 213.680 -17.710 213.860 -14.550 ;
        RECT 214.450 -27.250 214.620 -27.080 ;
        RECT 214.810 -27.250 214.980 -27.080 ;
        RECT 215.170 -27.250 215.340 -27.080 ;
        RECT 215.530 -27.250 215.700 -27.080 ;
        RECT -149.910 -39.910 -148.000 -39.730 ;
        RECT 207.740 -39.450 207.910 -28.470 ;
        RECT 208.340 -39.440 208.510 -28.460 ;
        RECT 208.950 -39.450 209.120 -28.470 ;
        RECT 209.550 -39.400 209.720 -28.420 ;
        RECT 210.150 -39.400 210.320 -28.420 ;
        RECT 210.740 -39.410 210.910 -28.430 ;
        RECT 211.320 -39.430 211.490 -28.450 ;
        RECT 211.940 -39.440 212.110 -28.460 ;
        RECT 212.560 -39.440 212.730 -28.460 ;
        RECT 214.480 -33.930 214.650 -33.760 ;
        RECT 214.850 -33.930 215.020 -33.760 ;
        RECT 215.210 -33.930 215.380 -33.760 ;
        RECT -149.910 -40.310 -148.010 -40.130 ;
        RECT 213.690 -39.210 213.860 -39.200 ;
        RECT 211.590 -40.630 213.500 -40.450 ;
        RECT 211.600 -41.030 213.500 -40.850 ;
        RECT 213.690 -41.070 213.870 -39.210 ;
        RECT -150.040 -42.010 -149.110 -41.810 ;
        RECT -150.270 -45.580 -150.090 -42.420 ;
        RECT -147.170 -43.080 -143.870 -42.730 ;
        RECT -152.110 -55.120 -151.940 -54.950 ;
        RECT -151.750 -55.120 -151.580 -54.950 ;
        RECT -151.390 -55.120 -151.220 -54.950 ;
        RECT -151.030 -55.120 -150.860 -54.950 ;
        RECT -148.380 -53.580 -148.210 -44.130 ;
        RECT -147.630 -53.590 -147.460 -44.200 ;
        RECT -146.910 -53.560 -146.740 -44.160 ;
        RECT -146.250 -53.550 -146.080 -44.180 ;
        RECT -145.600 -53.560 -145.430 -44.110 ;
        RECT -144.960 -53.550 -144.790 -44.160 ;
        RECT -151.790 -61.800 -151.620 -61.630 ;
        RECT -151.430 -61.800 -151.260 -61.630 ;
        RECT -151.060 -61.800 -150.890 -61.630 ;
        RECT -150.270 -67.080 -150.100 -67.070 ;
        RECT -150.280 -68.940 -150.100 -67.080 ;
        RECT -149.140 -67.310 -148.970 -56.330 ;
        RECT -148.520 -67.310 -148.350 -56.330 ;
        RECT -147.900 -67.300 -147.730 -56.320 ;
        RECT -147.320 -67.280 -147.150 -56.300 ;
        RECT -146.730 -67.270 -146.560 -56.290 ;
        RECT -146.130 -67.270 -145.960 -56.290 ;
        RECT -145.530 -67.320 -145.360 -56.340 ;
        RECT -144.920 -67.310 -144.750 -56.330 ;
        RECT -144.320 -67.320 -144.150 -56.340 ;
        RECT 212.700 -42.730 213.630 -42.530 ;
        RECT 207.460 -43.800 210.760 -43.450 ;
        RECT 208.380 -54.270 208.550 -44.880 ;
        RECT 209.020 -54.280 209.190 -44.830 ;
        RECT 209.670 -54.270 209.840 -44.900 ;
        RECT 210.330 -54.280 210.500 -44.880 ;
        RECT 211.050 -54.310 211.220 -44.920 ;
        RECT 211.800 -54.300 211.970 -44.850 ;
        RECT 213.680 -46.300 213.860 -43.140 ;
        RECT 214.450 -55.840 214.620 -55.670 ;
        RECT 214.810 -55.840 214.980 -55.670 ;
        RECT 215.170 -55.840 215.340 -55.670 ;
        RECT 215.530 -55.840 215.700 -55.670 ;
        RECT -149.910 -68.500 -148.000 -68.320 ;
        RECT 207.740 -68.040 207.910 -57.060 ;
        RECT 208.340 -68.030 208.510 -57.050 ;
        RECT 208.950 -68.040 209.120 -57.060 ;
        RECT 209.550 -67.990 209.720 -57.010 ;
        RECT 210.150 -67.990 210.320 -57.010 ;
        RECT 210.740 -68.000 210.910 -57.020 ;
        RECT 211.320 -68.020 211.490 -57.040 ;
        RECT 211.940 -68.030 212.110 -57.050 ;
        RECT 212.560 -68.030 212.730 -57.050 ;
        RECT 214.480 -62.520 214.650 -62.350 ;
        RECT 214.850 -62.520 215.020 -62.350 ;
        RECT 215.210 -62.520 215.380 -62.350 ;
        RECT -149.910 -68.900 -148.010 -68.720 ;
        RECT 213.690 -67.800 213.860 -67.790 ;
        RECT 211.590 -69.220 213.500 -69.040 ;
        RECT 211.600 -69.620 213.500 -69.440 ;
        RECT 213.690 -69.660 213.870 -67.800 ;
        RECT -150.040 -70.600 -149.110 -70.400 ;
        RECT -150.270 -74.170 -150.090 -71.010 ;
        RECT -147.170 -71.670 -143.870 -71.320 ;
        RECT -152.110 -83.710 -151.940 -83.540 ;
        RECT -151.750 -83.710 -151.580 -83.540 ;
        RECT -151.390 -83.710 -151.220 -83.540 ;
        RECT -151.030 -83.710 -150.860 -83.540 ;
        RECT -148.380 -82.170 -148.210 -72.720 ;
        RECT -147.630 -82.180 -147.460 -72.790 ;
        RECT -146.910 -82.150 -146.740 -72.750 ;
        RECT -146.250 -82.140 -146.080 -72.770 ;
        RECT -145.600 -82.150 -145.430 -72.700 ;
        RECT -144.960 -82.140 -144.790 -72.750 ;
        RECT -151.790 -90.390 -151.620 -90.220 ;
        RECT -151.430 -90.390 -151.260 -90.220 ;
        RECT -151.060 -90.390 -150.890 -90.220 ;
        RECT -150.270 -95.670 -150.100 -95.660 ;
        RECT -150.280 -97.530 -150.100 -95.670 ;
        RECT -149.140 -95.900 -148.970 -84.920 ;
        RECT -148.520 -95.900 -148.350 -84.920 ;
        RECT -147.900 -95.890 -147.730 -84.910 ;
        RECT -147.320 -95.870 -147.150 -84.890 ;
        RECT -146.730 -95.860 -146.560 -84.880 ;
        RECT -146.130 -95.860 -145.960 -84.880 ;
        RECT -145.530 -95.910 -145.360 -84.930 ;
        RECT -144.920 -95.900 -144.750 -84.920 ;
        RECT -144.320 -95.910 -144.150 -84.930 ;
        RECT -149.910 -97.090 -148.000 -96.910 ;
        RECT -149.910 -97.490 -148.010 -97.310 ;
        RECT -150.040 -99.190 -149.110 -98.990 ;
        RECT -150.270 -102.760 -150.090 -99.600 ;
        RECT -147.170 -100.260 -143.870 -99.910 ;
        RECT -152.110 -112.300 -151.940 -112.130 ;
        RECT -151.750 -112.300 -151.580 -112.130 ;
        RECT -151.390 -112.300 -151.220 -112.130 ;
        RECT -151.030 -112.300 -150.860 -112.130 ;
        RECT -148.380 -110.760 -148.210 -101.310 ;
        RECT -147.630 -110.770 -147.460 -101.380 ;
        RECT -146.910 -110.740 -146.740 -101.340 ;
        RECT -146.250 -110.730 -146.080 -101.360 ;
        RECT -145.600 -110.740 -145.430 -101.290 ;
        RECT -144.960 -110.730 -144.790 -101.340 ;
        RECT -151.790 -118.980 -151.620 -118.810 ;
        RECT -151.430 -118.980 -151.260 -118.810 ;
        RECT -151.060 -118.980 -150.890 -118.810 ;
        RECT -150.270 -124.260 -150.100 -124.250 ;
        RECT -150.280 -126.120 -150.100 -124.260 ;
        RECT -149.140 -124.490 -148.970 -113.510 ;
        RECT -148.520 -124.490 -148.350 -113.510 ;
        RECT -147.900 -124.480 -147.730 -113.500 ;
        RECT -147.320 -124.460 -147.150 -113.480 ;
        RECT -146.730 -124.450 -146.560 -113.470 ;
        RECT -146.130 -124.450 -145.960 -113.470 ;
        RECT -145.530 -124.500 -145.360 -113.520 ;
        RECT -144.920 -124.490 -144.750 -113.510 ;
        RECT -144.320 -124.500 -144.150 -113.520 ;
        RECT -149.910 -125.680 -148.000 -125.500 ;
        RECT -149.910 -126.080 -148.010 -125.900 ;
        RECT -150.040 -127.780 -149.110 -127.580 ;
        RECT -150.270 -131.350 -150.090 -128.190 ;
        RECT -147.170 -128.850 -143.870 -128.500 ;
        RECT -152.110 -140.890 -151.940 -140.720 ;
        RECT -151.750 -140.890 -151.580 -140.720 ;
        RECT -151.390 -140.890 -151.220 -140.720 ;
        RECT -151.030 -140.890 -150.860 -140.720 ;
        RECT -148.380 -139.350 -148.210 -129.900 ;
        RECT -147.630 -139.360 -147.460 -129.970 ;
        RECT -146.910 -139.330 -146.740 -129.930 ;
        RECT -146.250 -139.320 -146.080 -129.950 ;
        RECT -145.600 -139.330 -145.430 -129.880 ;
        RECT -144.960 -139.320 -144.790 -129.930 ;
        RECT -151.790 -147.570 -151.620 -147.400 ;
        RECT -151.430 -147.570 -151.260 -147.400 ;
        RECT -151.060 -147.570 -150.890 -147.400 ;
        RECT -150.270 -152.850 -150.100 -152.840 ;
        RECT -150.280 -154.710 -150.100 -152.850 ;
        RECT -149.140 -153.080 -148.970 -142.100 ;
        RECT -148.520 -153.080 -148.350 -142.100 ;
        RECT -147.900 -153.070 -147.730 -142.090 ;
        RECT -147.320 -153.050 -147.150 -142.070 ;
        RECT -146.730 -153.040 -146.560 -142.060 ;
        RECT -146.130 -153.040 -145.960 -142.060 ;
        RECT -145.530 -153.090 -145.360 -142.110 ;
        RECT -144.920 -153.080 -144.750 -142.100 ;
        RECT -144.320 -153.090 -144.150 -142.110 ;
        RECT -149.910 -154.270 -148.000 -154.090 ;
        RECT -149.910 -154.670 -148.010 -154.490 ;
        RECT -150.040 -156.370 -149.110 -156.170 ;
        RECT -150.270 -159.940 -150.090 -156.780 ;
        RECT -147.170 -157.440 -143.870 -157.090 ;
        RECT -152.110 -169.480 -151.940 -169.310 ;
        RECT -151.750 -169.480 -151.580 -169.310 ;
        RECT -151.390 -169.480 -151.220 -169.310 ;
        RECT -151.030 -169.480 -150.860 -169.310 ;
        RECT -148.380 -167.940 -148.210 -158.490 ;
        RECT -147.630 -167.950 -147.460 -158.560 ;
        RECT -146.910 -167.920 -146.740 -158.520 ;
        RECT -146.250 -167.910 -146.080 -158.540 ;
        RECT -145.600 -167.920 -145.430 -158.470 ;
        RECT -144.960 -167.910 -144.790 -158.520 ;
        RECT -151.790 -176.160 -151.620 -175.990 ;
        RECT -151.430 -176.160 -151.260 -175.990 ;
        RECT -151.060 -176.160 -150.890 -175.990 ;
        RECT -150.270 -181.440 -150.100 -181.430 ;
        RECT -150.280 -183.300 -150.100 -181.440 ;
        RECT -149.140 -181.670 -148.970 -170.690 ;
        RECT -148.520 -181.670 -148.350 -170.690 ;
        RECT -147.900 -181.660 -147.730 -170.680 ;
        RECT -147.320 -181.640 -147.150 -170.660 ;
        RECT -146.730 -181.630 -146.560 -170.650 ;
        RECT -146.130 -181.630 -145.960 -170.650 ;
        RECT -145.530 -181.680 -145.360 -170.700 ;
        RECT -144.920 -181.670 -144.750 -170.690 ;
        RECT -144.320 -181.680 -144.150 -170.700 ;
        RECT -149.910 -182.860 -148.000 -182.680 ;
        RECT -149.910 -183.260 -148.010 -183.080 ;
        RECT -150.040 -184.960 -149.110 -184.760 ;
        RECT -150.270 -188.530 -150.090 -185.370 ;
        RECT -147.170 -186.030 -143.870 -185.680 ;
        RECT -152.110 -198.070 -151.940 -197.900 ;
        RECT -151.750 -198.070 -151.580 -197.900 ;
        RECT -151.390 -198.070 -151.220 -197.900 ;
        RECT -151.030 -198.070 -150.860 -197.900 ;
        RECT -148.380 -196.530 -148.210 -187.080 ;
        RECT -147.630 -196.540 -147.460 -187.150 ;
        RECT -146.910 -196.510 -146.740 -187.110 ;
        RECT -146.250 -196.500 -146.080 -187.130 ;
        RECT -145.600 -196.510 -145.430 -187.060 ;
        RECT -144.960 -196.500 -144.790 -187.110 ;
        RECT -151.790 -204.750 -151.620 -204.580 ;
        RECT -151.430 -204.750 -151.260 -204.580 ;
        RECT -151.060 -204.750 -150.890 -204.580 ;
        RECT -150.270 -210.030 -150.100 -210.020 ;
        RECT -150.280 -211.890 -150.100 -210.030 ;
        RECT -149.140 -210.260 -148.970 -199.280 ;
        RECT -148.520 -210.260 -148.350 -199.280 ;
        RECT -147.900 -210.250 -147.730 -199.270 ;
        RECT -147.320 -210.230 -147.150 -199.250 ;
        RECT -146.730 -210.220 -146.560 -199.240 ;
        RECT -146.130 -210.220 -145.960 -199.240 ;
        RECT -145.530 -210.270 -145.360 -199.290 ;
        RECT -144.920 -210.260 -144.750 -199.280 ;
        RECT -144.320 -210.270 -144.150 -199.290 ;
        RECT -149.910 -211.450 -148.000 -211.270 ;
        RECT -149.910 -211.850 -148.010 -211.670 ;
        RECT -150.040 -213.550 -149.110 -213.350 ;
        RECT -150.270 -217.120 -150.090 -213.960 ;
        RECT -147.170 -214.620 -143.870 -214.270 ;
        RECT -152.110 -226.660 -151.940 -226.490 ;
        RECT -151.750 -226.660 -151.580 -226.490 ;
        RECT -151.390 -226.660 -151.220 -226.490 ;
        RECT -151.030 -226.660 -150.860 -226.490 ;
        RECT -148.380 -225.120 -148.210 -215.670 ;
        RECT -147.630 -225.130 -147.460 -215.740 ;
        RECT -146.910 -225.100 -146.740 -215.700 ;
        RECT -146.250 -225.090 -146.080 -215.720 ;
        RECT -145.600 -225.100 -145.430 -215.650 ;
        RECT -144.960 -225.090 -144.790 -215.700 ;
        RECT -151.790 -233.340 -151.620 -233.170 ;
        RECT -151.430 -233.340 -151.260 -233.170 ;
        RECT -151.060 -233.340 -150.890 -233.170 ;
        RECT -150.270 -238.620 -150.100 -238.610 ;
        RECT -150.280 -240.480 -150.100 -238.620 ;
        RECT -149.140 -238.850 -148.970 -227.870 ;
        RECT -148.520 -238.850 -148.350 -227.870 ;
        RECT -147.900 -238.840 -147.730 -227.860 ;
        RECT -147.320 -238.820 -147.150 -227.840 ;
        RECT -146.730 -238.810 -146.560 -227.830 ;
        RECT -146.130 -238.810 -145.960 -227.830 ;
        RECT -145.530 -238.860 -145.360 -227.880 ;
        RECT -144.920 -238.850 -144.750 -227.870 ;
        RECT -144.320 -238.860 -144.150 -227.880 ;
        RECT -149.910 -240.040 -148.000 -239.860 ;
        RECT -149.910 -240.440 -148.010 -240.260 ;
      LAYER met1 ;
        RECT -124.420 143.120 -124.070 143.280 ;
        RECT -95.830 143.120 -95.480 143.280 ;
        RECT -67.240 143.120 -66.890 143.280 ;
        RECT -124.430 142.170 -124.060 143.120 ;
        RECT -95.840 142.170 -95.470 143.120 ;
        RECT -67.250 142.170 -66.880 143.120 ;
        RECT -25.230 142.460 -24.820 143.230 ;
        RECT 16.780 143.120 17.130 143.280 ;
        RECT 45.370 143.120 45.720 143.280 ;
        RECT 73.960 143.120 74.310 143.280 ;
        RECT 102.550 143.120 102.900 143.280 ;
        RECT 131.140 143.120 131.490 143.280 ;
        RECT 159.730 143.120 160.080 143.280 ;
        RECT 188.320 143.120 188.670 143.280 ;
        RECT -25.500 142.190 -24.820 142.460 ;
        RECT -124.780 141.800 -122.310 142.170 ;
        RECT -96.190 141.800 -93.720 142.170 ;
        RECT -67.600 141.800 -65.130 142.170 ;
        RECT -138.330 141.000 -135.960 141.630 ;
        RECT -138.300 139.040 -137.350 141.000 ;
        RECT -136.600 140.980 -136.020 141.000 ;
        RECT -126.220 140.340 -122.310 141.800 ;
        RECT -114.990 141.150 -110.860 141.550 ;
        RECT -114.990 141.060 -110.850 141.150 ;
        RECT -135.930 140.330 -122.310 140.340 ;
        RECT -138.070 133.370 -137.350 139.040 ;
        RECT -136.600 139.770 -122.310 140.330 ;
        RECT -111.380 140.160 -110.850 141.060 ;
        RECT -109.740 141.000 -107.370 141.630 ;
        RECT -136.600 135.470 -113.250 139.770 ;
        RECT -109.710 139.040 -108.760 141.000 ;
        RECT -108.010 140.980 -107.430 141.000 ;
        RECT -97.630 140.340 -93.720 141.800 ;
        RECT -86.400 141.150 -82.270 141.550 ;
        RECT -86.400 141.060 -82.260 141.150 ;
        RECT -107.340 140.330 -93.720 140.340 ;
        RECT -112.480 138.350 -111.910 138.360 ;
        RECT -136.600 135.190 -122.310 135.470 ;
        RECT -126.220 133.640 -122.310 135.190 ;
        RECT -112.480 134.930 -111.860 138.350 ;
        RECT -112.480 134.920 -111.910 134.930 ;
        RECT -126.240 132.100 -122.290 133.640 ;
        RECT -113.310 133.290 -112.750 133.790 ;
        RECT -109.480 133.370 -108.760 139.040 ;
        RECT -108.010 139.770 -93.720 140.330 ;
        RECT -82.790 140.160 -82.260 141.060 ;
        RECT -81.150 141.000 -78.780 141.630 ;
        RECT -108.010 135.470 -84.660 139.770 ;
        RECT -81.120 139.040 -80.170 141.000 ;
        RECT -79.420 140.980 -78.840 141.000 ;
        RECT -69.040 140.340 -65.130 141.800 ;
        RECT -25.500 141.760 -23.810 142.190 ;
        RECT 16.770 142.170 17.140 143.120 ;
        RECT 45.360 142.170 45.730 143.120 ;
        RECT 73.950 142.170 74.320 143.120 ;
        RECT 102.540 142.170 102.910 143.120 ;
        RECT 131.130 142.170 131.500 143.120 ;
        RECT 159.720 142.170 160.090 143.120 ;
        RECT 188.310 142.170 188.680 143.120 ;
        RECT 16.420 141.800 18.890 142.170 ;
        RECT 45.010 141.800 47.480 142.170 ;
        RECT 73.600 141.800 76.070 142.170 ;
        RECT 102.190 141.800 104.660 142.170 ;
        RECT 130.780 141.800 133.250 142.170 ;
        RECT 159.370 141.800 161.840 142.170 ;
        RECT 187.960 141.800 190.430 142.170 ;
        RECT -52.710 141.580 -28.340 141.600 ;
        RECT -57.810 141.150 -53.680 141.550 ;
        RECT -52.770 141.190 -28.340 141.580 ;
        RECT -57.810 141.060 -53.670 141.150 ;
        RECT -78.750 140.330 -65.130 140.340 ;
        RECT -83.890 138.350 -83.320 138.360 ;
        RECT -108.010 135.190 -93.720 135.470 ;
        RECT -97.630 133.640 -93.720 135.190 ;
        RECT -83.890 134.930 -83.270 138.350 ;
        RECT -83.890 134.920 -83.320 134.930 ;
        RECT -113.300 133.070 -112.750 133.290 ;
        RECT -97.650 132.870 -93.700 133.640 ;
        RECT -84.720 133.290 -84.160 133.790 ;
        RECT -80.890 133.370 -80.170 139.040 ;
        RECT -79.420 139.770 -65.130 140.330 ;
        RECT -54.200 140.160 -53.670 141.060 ;
        RECT -79.420 135.470 -56.070 139.770 ;
        RECT -55.300 138.350 -54.730 138.360 ;
        RECT -79.420 135.190 -65.130 135.470 ;
        RECT -69.040 133.640 -65.130 135.190 ;
        RECT -55.300 134.930 -54.680 138.350 ;
        RECT -55.300 134.920 -54.730 134.930 ;
        RECT -84.710 133.070 -84.160 133.290 ;
        RECT -97.640 132.100 -93.690 132.870 ;
        RECT -69.060 132.100 -65.110 133.640 ;
        RECT -56.130 133.290 -55.570 133.790 ;
        RECT -56.120 133.120 -55.570 133.290 ;
        RECT -56.170 133.070 -55.570 133.120 ;
        RECT -150.030 129.880 -149.040 129.890 ;
        RECT -150.430 129.360 -149.040 129.880 ;
        RECT -150.430 125.750 -149.940 129.360 ;
        RECT -147.230 128.830 -143.810 128.880 ;
        RECT -147.240 128.260 -143.800 128.830 ;
        RECT -148.650 118.430 -144.350 127.490 ;
        RECT -142.670 127.440 -141.950 127.990 ;
        RECT -142.670 127.430 -142.170 127.440 ;
        RECT -125.540 122.220 -122.310 132.100 ;
        RECT -96.950 125.630 -93.720 132.100 ;
        RECT -68.360 129.920 -65.130 132.100 ;
        RECT -68.790 127.180 -64.960 129.920 ;
        RECT -56.170 126.560 -55.650 133.070 ;
        RECT -56.230 126.050 -55.580 126.560 ;
        RECT -97.110 122.740 -93.610 125.630 ;
        RECT -127.710 118.600 -122.310 122.220 ;
        RECT -140.150 118.520 -136.760 118.590 ;
        RECT -142.520 118.440 -141.750 118.450 ;
        RECT -141.120 118.440 -136.760 118.520 ;
        RECT -142.520 118.430 -136.760 118.440 ;
        RECT -151.050 116.680 -136.760 118.430 ;
        RECT -127.710 118.420 -124.770 118.600 ;
        RECT -56.170 118.370 -55.650 126.050 ;
        RECT -52.770 122.140 -52.360 141.190 ;
        RECT -26.170 133.690 -23.810 141.760 ;
        RECT -19.540 141.590 1.820 141.600 ;
        RECT -19.600 141.200 1.820 141.590 ;
        RECT -19.600 141.190 1.660 141.200 ;
        RECT 2.870 141.000 5.240 141.630 ;
        RECT 2.900 139.040 3.850 141.000 ;
        RECT 4.600 140.980 5.180 141.000 ;
        RECT 14.980 140.340 18.890 141.800 ;
        RECT 26.210 141.150 30.340 141.550 ;
        RECT 26.210 141.060 30.350 141.150 ;
        RECT 5.270 140.330 18.890 140.340 ;
        RECT -26.290 132.100 -23.810 133.690 ;
        RECT 3.130 133.370 3.850 139.040 ;
        RECT 4.600 139.770 18.890 140.330 ;
        RECT 29.820 140.160 30.350 141.060 ;
        RECT 31.460 141.000 33.830 141.630 ;
        RECT 4.600 135.470 27.950 139.770 ;
        RECT 31.490 139.040 32.440 141.000 ;
        RECT 33.190 140.980 33.770 141.000 ;
        RECT 43.570 140.340 47.480 141.800 ;
        RECT 54.800 141.150 58.930 141.550 ;
        RECT 54.800 141.060 58.940 141.150 ;
        RECT 33.860 140.330 47.480 140.340 ;
        RECT 28.720 138.350 29.290 138.360 ;
        RECT 4.600 135.190 18.890 135.470 ;
        RECT 14.980 133.640 18.890 135.190 ;
        RECT 28.720 134.930 29.340 138.350 ;
        RECT 28.720 134.920 29.290 134.930 ;
        RECT 14.960 132.110 18.910 133.640 ;
        RECT 27.890 133.400 28.450 133.790 ;
        RECT 27.300 133.260 28.450 133.400 ;
        RECT -25.660 131.350 -24.500 132.100 ;
        RECT -25.660 130.220 1.700 131.350 ;
        RECT -25.660 130.020 1.890 130.220 ;
        RECT 0.370 129.630 1.700 130.020 ;
        RECT 0.360 129.180 1.700 129.630 ;
        RECT -25.740 128.340 -25.240 128.820 ;
        RECT 0.360 128.760 13.880 129.180 ;
        RECT 15.660 129.110 18.890 132.110 ;
        RECT 27.280 131.300 28.460 133.260 ;
        RECT 26.480 130.390 28.460 131.300 ;
        RECT 26.480 130.210 28.290 130.390 ;
        RECT 31.720 130.250 32.440 139.040 ;
        RECT 33.190 139.770 47.480 140.330 ;
        RECT 58.410 140.160 58.940 141.060 ;
        RECT 60.050 141.000 62.420 141.630 ;
        RECT 33.190 135.470 56.540 139.770 ;
        RECT 60.080 139.040 61.030 141.000 ;
        RECT 61.780 140.980 62.360 141.000 ;
        RECT 72.160 140.340 76.070 141.800 ;
        RECT 83.390 141.150 87.520 141.550 ;
        RECT 83.390 141.060 87.530 141.150 ;
        RECT 62.450 140.330 76.070 140.340 ;
        RECT 57.310 138.350 57.880 138.360 ;
        RECT 33.190 135.190 47.480 135.470 ;
        RECT 43.570 133.640 47.480 135.190 ;
        RECT 57.310 134.930 57.930 138.350 ;
        RECT 57.310 134.920 57.880 134.930 ;
        RECT 43.550 132.100 47.500 133.640 ;
        RECT 56.480 133.290 57.040 133.790 ;
        RECT 56.490 133.070 57.040 133.290 ;
        RECT 52.430 132.350 52.770 132.490 ;
        RECT 60.310 132.350 61.030 139.040 ;
        RECT 61.780 139.770 76.070 140.330 ;
        RECT 87.000 140.160 87.530 141.060 ;
        RECT 88.640 141.000 91.010 141.630 ;
        RECT 61.780 135.470 85.130 139.770 ;
        RECT 88.670 139.040 89.620 141.000 ;
        RECT 90.370 140.980 90.950 141.000 ;
        RECT 100.750 140.340 104.660 141.800 ;
        RECT 111.980 141.150 116.110 141.550 ;
        RECT 111.980 141.060 116.120 141.150 ;
        RECT 91.040 140.330 104.660 140.340 ;
        RECT 85.900 138.350 86.470 138.360 ;
        RECT 61.780 135.190 76.070 135.470 ;
        RECT 72.160 133.640 76.070 135.190 ;
        RECT 85.900 134.930 86.520 138.350 ;
        RECT 85.900 134.920 86.470 134.930 ;
        RECT 15.670 129.090 18.860 129.110 ;
        RECT 0.360 128.620 1.700 128.760 ;
        RECT -52.890 121.670 -52.360 122.140 ;
        RECT -56.370 117.640 -55.650 118.370 ;
        RECT -152.000 116.670 -136.760 116.680 ;
        RECT -152.160 116.320 -136.760 116.670 ;
        RECT -152.000 116.310 -136.760 116.320 ;
        RECT -151.050 115.960 -136.760 116.310 ;
        RECT -150.680 114.520 -136.760 115.960 ;
        RECT -149.220 104.810 -144.070 114.520 ;
        RECT -142.520 114.500 -141.120 114.520 ;
        RECT -150.510 104.720 -149.880 104.780 ;
        RECT -150.510 104.140 -149.860 104.720 ;
        RECT -149.210 104.140 -144.070 104.810 ;
        RECT -150.510 103.390 -149.880 104.140 ;
        RECT -150.510 102.670 -142.250 103.390 ;
        RECT -150.510 102.440 -147.920 102.670 ;
        RECT -150.510 102.410 -149.880 102.440 ;
        RECT -150.030 101.290 -149.040 101.300 ;
        RECT -150.430 100.770 -149.040 101.290 ;
        RECT -150.430 97.160 -149.940 100.770 ;
        RECT -147.230 100.240 -143.810 100.290 ;
        RECT -147.240 99.670 -143.800 100.240 ;
        RECT -148.650 89.840 -144.350 98.900 ;
        RECT -142.670 98.850 -141.950 99.400 ;
        RECT -142.670 98.840 -142.170 98.850 ;
        RECT -142.520 89.840 -141.120 89.860 ;
        RECT -130.980 89.840 -128.720 89.880 ;
        RECT -151.050 88.090 -128.720 89.840 ;
        RECT -152.000 88.080 -128.720 88.090 ;
        RECT -152.160 87.730 -128.720 88.080 ;
        RECT -152.000 87.720 -128.720 87.730 ;
        RECT -151.050 87.370 -128.720 87.720 ;
        RECT -150.680 86.610 -128.720 87.370 ;
        RECT -150.680 85.930 -141.120 86.610 ;
        RECT -130.980 86.570 -128.720 86.610 ;
        RECT -149.220 76.220 -144.070 85.930 ;
        RECT -142.520 85.920 -141.120 85.930 ;
        RECT -142.520 85.910 -141.750 85.920 ;
        RECT -56.170 82.290 -55.650 117.640 ;
        RECT -52.770 117.420 -52.360 121.670 ;
        RECT -25.640 125.380 -25.250 128.340 ;
        RECT -5.050 128.020 -2.280 128.260 ;
        RECT -23.270 127.560 -23.010 127.760 ;
        RECT -20.410 127.720 -20.150 127.810 ;
        RECT -23.330 127.250 -22.950 127.560 ;
        RECT -21.920 127.250 -20.890 127.560 ;
        RECT -20.420 127.490 -20.130 127.720 ;
        RECT -23.280 126.460 -23.020 126.730 ;
        RECT -22.590 126.460 -22.270 126.700 ;
        RECT -21.870 126.460 -21.610 126.740 ;
        RECT -23.320 125.800 -21.570 126.460 ;
        RECT -23.280 125.540 -23.020 125.800 ;
        RECT -22.590 125.540 -22.270 125.800 ;
        RECT -21.850 125.560 -21.590 125.800 ;
        RECT -25.640 124.890 -25.170 125.380 ;
        RECT -25.640 124.880 -25.190 124.890 ;
        RECT -52.910 116.830 -52.290 117.420 ;
        RECT -56.250 81.690 -55.620 82.290 ;
        RECT -52.770 81.270 -52.360 116.830 ;
        RECT -52.820 80.770 -52.340 81.270 ;
        RECT -150.510 76.130 -149.880 76.190 ;
        RECT -150.510 75.550 -149.860 76.130 ;
        RECT -149.210 75.550 -144.070 76.220 ;
        RECT -150.510 74.800 -149.880 75.550 ;
        RECT -150.510 74.080 -142.250 74.800 ;
        RECT -150.510 73.850 -147.920 74.080 ;
        RECT -150.510 73.820 -149.880 73.850 ;
        RECT -150.030 72.700 -149.040 72.710 ;
        RECT -150.430 72.180 -149.040 72.700 ;
        RECT -150.430 68.570 -149.940 72.180 ;
        RECT -147.230 71.650 -143.810 71.700 ;
        RECT -147.240 71.080 -143.800 71.650 ;
        RECT -148.650 61.250 -144.350 70.310 ;
        RECT -142.670 70.260 -141.950 70.810 ;
        RECT -142.670 70.250 -142.170 70.260 ;
        RECT -25.640 66.770 -25.250 124.880 ;
        RECT -23.260 124.510 -23.030 125.030 ;
        RECT -23.280 124.190 -23.020 124.510 ;
        RECT -24.230 123.740 -23.970 124.060 ;
        RECT -24.220 121.520 -23.980 123.740 ;
        RECT -23.260 123.620 -23.030 124.190 ;
        RECT -21.850 123.620 -21.620 125.030 ;
        RECT -21.130 124.480 -20.890 127.250 ;
        RECT -5.050 126.930 -4.810 128.020 ;
        RECT -20.470 126.800 -20.080 126.930 ;
        RECT -20.470 126.510 -20.050 126.800 ;
        RECT -5.050 126.670 -4.820 126.930 ;
        RECT -20.750 125.950 -20.430 126.270 ;
        RECT -20.700 125.720 -20.470 125.950 ;
        RECT -20.280 125.570 -20.050 126.510 ;
        RECT -5.060 126.450 -4.820 126.670 ;
        RECT -7.200 125.640 -6.880 125.960 ;
        RECT -5.840 125.720 -5.520 126.040 ;
        RECT -5.150 125.710 -4.830 126.030 ;
        RECT -20.410 125.500 -20.050 125.570 ;
        RECT -20.470 125.390 -20.050 125.500 ;
        RECT -20.470 125.270 -20.080 125.390 ;
        RECT -21.170 123.940 -20.850 124.260 ;
        RECT -20.410 124.100 -20.140 125.270 ;
        RECT -5.050 124.130 -4.810 124.770 ;
        RECT -20.410 123.870 -20.080 124.100 ;
        RECT -5.050 123.870 -4.820 124.130 ;
        RECT -5.060 123.220 -4.820 123.870 ;
        RECT -22.610 122.740 -22.290 123.060 ;
        RECT -21.180 122.760 -20.860 123.080 ;
        RECT -23.400 122.160 -23.080 122.480 ;
        RECT -22.470 122.160 -22.150 122.480 ;
        RECT -21.770 122.160 -21.450 122.480 ;
        RECT -21.030 122.160 -20.710 122.480 ;
        RECT -20.320 122.150 -20.000 122.470 ;
        RECT -24.310 121.040 -23.890 121.520 ;
        RECT -18.420 120.280 -18.130 122.970 ;
        RECT -5.060 122.580 -4.810 123.220 ;
        RECT -7.920 121.980 -7.600 122.300 ;
        RECT -18.440 119.610 -18.030 120.280 ;
        RECT -5.060 118.920 -4.820 122.580 ;
        RECT -5.110 118.580 -4.770 118.920 ;
        RECT -7.860 118.480 -7.370 118.490 ;
        RECT -11.790 109.790 -11.560 113.270 ;
        RECT -11.120 112.650 -10.900 113.270 ;
        RECT -10.020 112.840 -9.700 113.160 ;
        RECT -8.930 112.850 -8.610 113.170 ;
        RECT -11.150 112.330 -10.890 112.650 ;
        RECT -10.450 112.340 -10.130 112.660 ;
        RECT -11.120 111.730 -10.900 112.330 ;
        RECT -10.010 111.850 -9.690 112.170 ;
        RECT -8.920 111.860 -8.600 112.180 ;
        RECT -11.180 111.410 -10.900 111.730 ;
        RECT -10.470 111.420 -10.150 111.740 ;
        RECT -11.120 110.810 -10.900 111.410 ;
        RECT -10.010 110.860 -9.690 111.180 ;
        RECT -8.920 110.870 -8.600 111.190 ;
        RECT -11.170 110.490 -10.900 110.810 ;
        RECT -11.820 109.470 -11.560 109.790 ;
        RECT -11.790 108.830 -11.560 109.470 ;
        RECT -11.860 108.510 -11.560 108.830 ;
        RECT -11.790 107.870 -11.560 108.510 ;
        RECT -11.820 107.550 -11.560 107.870 ;
        RECT -11.790 92.800 -11.560 107.550 ;
        RECT -11.120 92.800 -10.900 110.490 ;
        RECT -10.490 110.430 -10.170 110.750 ;
        RECT -10.200 109.930 -9.880 110.250 ;
        RECT -8.900 109.830 -8.580 110.150 ;
        RECT -10.230 109.750 -9.910 109.790 ;
        RECT -10.460 109.520 -9.910 109.750 ;
        RECT -10.230 109.470 -9.910 109.520 ;
        RECT -10.200 108.940 -9.880 109.260 ;
        RECT -8.900 108.840 -8.580 109.160 ;
        RECT -10.230 108.760 -9.910 108.800 ;
        RECT -10.460 108.530 -9.910 108.760 ;
        RECT -8.430 108.630 -8.210 117.540 ;
        RECT -7.870 117.330 -7.360 118.480 ;
        RECT -2.520 117.550 -2.280 128.020 ;
        RECT 0.790 127.690 3.820 127.960 ;
        RECT 0.790 126.710 1.060 127.690 ;
        RECT 0.800 124.500 1.060 124.520 ;
        RECT 0.760 118.520 1.070 124.500 ;
        RECT 1.940 122.000 2.260 122.320 ;
        RECT 0.680 118.150 1.070 118.520 ;
        RECT 3.550 118.010 3.820 127.690 ;
        RECT 5.500 126.670 5.760 128.760 ;
        RECT 13.460 125.510 13.880 128.760 ;
        RECT 17.270 126.270 17.690 129.090 ;
        RECT 17.270 125.790 17.740 126.270 ;
        RECT 13.420 125.030 13.900 125.510 ;
        RECT 4.730 123.960 4.960 124.130 ;
        RECT 4.720 122.090 4.970 123.960 ;
        RECT 18.970 123.420 19.410 123.920 ;
        RECT 24.690 123.420 25.130 123.920 ;
        RECT 14.550 122.400 14.990 122.900 ;
        RECT 4.720 121.910 4.980 122.090 ;
        RECT 4.720 119.010 4.970 121.910 ;
        RECT 11.760 119.660 12.080 119.710 ;
        RECT 11.670 119.370 12.080 119.660 ;
        RECT 4.680 118.650 5.010 119.010 ;
        RECT 3.510 117.700 3.850 118.010 ;
        RECT -7.920 117.230 -7.360 117.330 ;
        RECT -2.570 117.230 -2.230 117.550 ;
        RECT -8.030 116.830 -7.360 117.230 ;
        RECT 11.670 116.940 11.910 119.370 ;
        RECT 14.610 116.940 14.920 122.400 ;
        RECT -8.030 116.800 -7.370 116.830 ;
        RECT -8.030 112.580 -7.810 116.800 ;
        RECT 11.670 115.870 12.010 116.940 ;
        RECT 13.190 116.230 13.540 116.520 ;
        RECT 13.190 116.210 13.390 116.230 ;
        RECT 11.030 115.370 11.440 115.700 ;
        RECT -6.810 114.680 -6.460 115.140 ;
        RECT 9.620 114.700 9.990 115.010 ;
        RECT -7.410 114.320 -7.160 114.440 ;
        RECT -7.440 113.860 -7.120 114.320 ;
        RECT -8.040 112.290 -7.810 112.580 ;
        RECT -10.230 108.480 -9.910 108.530 ;
        RECT -8.480 108.400 -8.190 108.630 ;
        RECT -10.200 107.950 -9.880 108.270 ;
        RECT -8.900 107.850 -8.580 108.170 ;
        RECT -10.230 107.770 -9.910 107.810 ;
        RECT -10.460 107.540 -9.910 107.770 ;
        RECT -10.230 107.490 -9.910 107.540 ;
        RECT -11.900 92.270 -11.560 92.800 ;
        RECT -11.240 92.270 -10.900 92.800 ;
        RECT -13.210 91.530 -12.980 91.600 ;
        RECT -13.250 91.270 -12.930 91.530 ;
        RECT -13.700 91.160 -13.470 91.200 ;
        RECT -13.740 90.840 -13.470 91.160 ;
        RECT -23.050 89.600 -22.330 90.300 ;
        RECT -23.040 84.450 -22.380 89.600 ;
        RECT -13.700 87.320 -13.470 90.840 ;
        RECT -13.210 88.800 -12.980 91.270 ;
        RECT -11.790 91.180 -11.560 92.270 ;
        RECT -11.120 91.540 -10.900 92.270 ;
        RECT -9.360 91.560 -9.090 91.600 ;
        RECT -11.140 91.220 -10.880 91.540 ;
        RECT -9.380 91.230 -9.090 91.560 ;
        RECT -11.800 90.860 -11.540 91.180 ;
        RECT -11.080 90.260 -10.760 90.580 ;
        RECT -10.430 90.260 -10.110 90.580 ;
        RECT -12.300 89.820 -11.980 90.140 ;
        RECT -11.600 89.820 -11.280 90.140 ;
        RECT -9.910 88.810 -9.620 89.720 ;
        RECT -13.210 88.790 -12.480 88.800 ;
        RECT -13.210 88.470 -12.460 88.790 ;
        RECT -13.210 88.430 -12.480 88.470 ;
        RECT -13.700 87.250 -13.440 87.320 ;
        RECT -13.720 87.240 -13.440 87.250 ;
        RECT -13.750 86.930 -13.430 87.240 ;
        RECT -17.850 85.070 -17.420 85.500 ;
        RECT -23.040 83.730 -22.300 84.450 ;
        RECT -17.800 79.260 -17.430 85.070 ;
        RECT -13.210 80.930 -12.980 88.430 ;
        RECT -12.710 88.180 -12.480 88.430 ;
        RECT -10.000 88.240 -9.680 88.280 ;
        RECT -9.360 88.260 -9.090 91.230 ;
        RECT -9.480 88.240 -9.090 88.260 ;
        RECT -12.710 87.960 -12.490 88.180 ;
        RECT -10.000 88.010 -9.090 88.240 ;
        RECT -8.880 91.160 -8.640 91.200 ;
        RECT -8.880 90.840 -8.620 91.160 ;
        RECT -10.000 87.960 -9.680 88.010 ;
        RECT -12.690 87.530 -12.470 87.750 ;
        RECT -12.700 87.240 -12.470 87.530 ;
        RECT -9.990 87.700 -9.670 87.740 ;
        RECT -8.880 87.700 -8.640 90.840 ;
        RECT -9.990 87.470 -8.640 87.700 ;
        RECT -9.990 87.420 -9.670 87.470 ;
        RECT -12.720 86.920 -12.460 87.240 ;
        RECT -9.920 86.790 -9.650 86.970 ;
        RECT -9.940 86.470 -9.620 86.790 ;
        RECT -9.920 86.300 -9.650 86.470 ;
        RECT -12.270 85.940 -11.950 86.260 ;
        RECT -11.580 85.930 -11.260 86.250 ;
        RECT -11.100 85.160 -10.780 85.480 ;
        RECT -10.390 85.100 -10.070 85.420 ;
        RECT -13.210 80.700 -10.760 80.930 ;
        RECT -11.080 80.080 -10.760 80.700 ;
        RECT -14.390 79.640 -14.070 79.960 ;
        RECT -13.290 79.650 -12.970 79.970 ;
        RECT -12.200 79.650 -11.880 79.970 ;
        RECT -11.070 79.610 -10.750 79.930 ;
        RECT -17.840 78.830 -17.410 79.260 ;
        RECT -13.840 78.970 -13.520 79.290 ;
        RECT -12.740 78.970 -12.420 79.290 ;
        RECT -11.640 78.970 -11.320 79.290 ;
        RECT -10.930 78.800 -10.640 79.230 ;
        RECT -10.320 78.800 -9.990 78.830 ;
        RECT -10.930 78.780 -9.990 78.800 ;
        RECT -10.920 78.480 -9.990 78.780 ;
        RECT -10.920 77.950 -10.640 78.480 ;
        RECT -10.320 78.410 -9.990 78.480 ;
        RECT -10.910 77.920 -10.640 77.950 ;
        RECT -13.840 77.600 -13.520 77.920 ;
        RECT -12.740 77.600 -12.420 77.920 ;
        RECT -11.640 77.600 -11.320 77.920 ;
        RECT -14.390 76.870 -14.070 77.190 ;
        RECT -13.290 76.870 -12.970 77.190 ;
        RECT -12.200 76.870 -11.880 77.190 ;
        RECT -14.400 75.530 -14.080 75.850 ;
        RECT -13.290 75.520 -12.970 75.840 ;
        RECT -12.200 75.500 -11.880 75.820 ;
        RECT -13.840 74.830 -13.520 75.150 ;
        RECT -12.740 74.820 -12.420 75.140 ;
        RECT -11.650 74.820 -11.330 75.140 ;
        RECT -14.830 73.170 -14.540 73.520 ;
        RECT -14.820 67.880 -14.560 73.170 ;
        RECT -11.040 72.530 -10.720 72.850 ;
        RECT -8.880 72.810 -8.640 87.470 ;
        RECT -8.430 86.800 -8.210 108.400 ;
        RECT -8.030 89.410 -7.810 112.290 ;
        RECT -7.410 113.070 -7.160 113.860 ;
        RECT -7.410 112.750 -7.120 113.070 ;
        RECT -7.410 112.150 -7.160 112.750 ;
        RECT -7.410 111.830 -7.120 112.150 ;
        RECT -7.410 111.230 -7.160 111.830 ;
        RECT -7.410 110.910 -7.150 111.230 ;
        RECT -7.410 90.560 -7.160 110.910 ;
        RECT -6.790 110.140 -6.530 114.680 ;
        RECT 8.980 112.980 9.370 113.350 ;
        RECT 8.400 111.490 8.790 111.880 ;
        RECT -6.790 109.820 -6.510 110.140 ;
        RECT 7.760 109.900 8.150 110.280 ;
        RECT 7.790 109.890 8.130 109.900 ;
        RECT -6.790 109.180 -6.530 109.820 ;
        RECT 7.150 109.700 7.490 109.710 ;
        RECT 7.140 109.310 7.500 109.700 ;
        RECT -6.790 108.860 -6.500 109.180 ;
        RECT -6.790 108.220 -6.530 108.860 ;
        RECT -6.790 107.900 -6.510 108.220 ;
        RECT -7.410 90.540 -7.150 90.560 ;
        RECT -7.420 90.260 -7.140 90.540 ;
        RECT -7.410 90.240 -7.150 90.260 ;
        RECT -8.070 89.090 -7.750 89.410 ;
        RECT -8.470 86.480 -8.190 86.800 ;
        RECT -8.430 73.510 -8.210 86.480 ;
        RECT -8.030 81.270 -7.810 89.090 ;
        RECT -8.030 80.790 -7.740 81.270 ;
        RECT -8.030 78.830 -7.810 80.790 ;
        RECT -8.050 78.410 -7.790 78.830 ;
        RECT -8.030 73.790 -7.810 78.410 ;
        RECT -7.410 75.170 -7.160 90.240 ;
        RECT -6.790 86.230 -6.530 107.900 ;
        RECT 6.530 107.750 6.890 108.140 ;
        RECT 5.880 106.210 6.290 106.610 ;
        RECT 5.350 104.650 5.710 105.040 ;
        RECT 4.770 99.590 5.100 99.610 ;
        RECT 4.710 99.170 5.100 99.590 ;
        RECT 4.140 97.980 4.470 98.000 ;
        RECT 4.090 97.590 4.480 97.980 ;
        RECT 3.520 96.430 3.850 96.440 ;
        RECT 3.490 96.040 3.850 96.430 ;
        RECT 2.870 94.560 3.260 94.960 ;
        RECT 2.200 89.390 2.630 89.790 ;
        RECT 1.540 87.820 1.950 88.220 ;
        RECT -6.800 85.910 -6.490 86.230 ;
        RECT 0.930 86.180 1.320 86.580 ;
        RECT -7.450 74.770 -7.150 75.170 ;
        RECT -8.030 73.650 -7.790 73.790 ;
        RECT -8.470 73.160 -8.160 73.510 ;
        RECT -8.020 73.020 -7.790 73.650 ;
        RECT -14.350 72.090 -14.030 72.410 ;
        RECT -13.250 72.100 -12.930 72.420 ;
        RECT -12.160 72.100 -11.840 72.420 ;
        RECT -11.030 72.060 -10.710 72.380 ;
        RECT -9.670 72.250 -8.640 72.810 ;
        RECT -8.030 72.990 -7.790 73.020 ;
        RECT -9.670 72.140 -8.880 72.250 ;
        RECT -13.800 71.420 -13.480 71.740 ;
        RECT -12.700 71.420 -12.380 71.740 ;
        RECT -11.600 71.420 -11.280 71.740 ;
        RECT -8.030 71.600 -7.810 72.990 ;
        RECT -13.800 70.050 -13.480 70.370 ;
        RECT -12.700 70.050 -12.380 70.370 ;
        RECT -11.600 70.050 -11.280 70.370 ;
        RECT -14.350 69.320 -14.030 69.640 ;
        RECT -13.250 69.320 -12.930 69.640 ;
        RECT -12.160 69.320 -11.840 69.640 ;
        RECT -14.360 67.980 -14.040 68.300 ;
        RECT -13.250 67.970 -12.930 68.290 ;
        RECT -12.160 67.950 -11.840 68.270 ;
        RECT -9.560 67.920 -7.140 71.600 ;
        RECT -14.870 67.070 -14.560 67.880 ;
        RECT -6.790 67.630 -6.530 85.910 ;
        RECT 0.240 84.740 0.650 85.130 ;
        RECT -3.970 79.590 -3.040 81.240 ;
        RECT -3.880 79.110 -3.140 79.590 ;
        RECT -13.800 67.280 -13.480 67.600 ;
        RECT -12.700 67.270 -12.380 67.590 ;
        RECT -11.610 67.270 -11.290 67.590 ;
        RECT -6.880 67.220 -6.530 67.630 ;
        RECT -14.820 66.870 -14.560 67.070 ;
        RECT -25.810 66.250 -25.250 66.770 ;
        RECT 0.300 61.400 0.630 84.740 ;
        RECT 0.250 61.390 0.680 61.400 ;
        RECT -142.520 61.250 -141.750 61.270 ;
        RECT -127.070 61.250 -124.840 61.330 ;
        RECT -151.050 59.500 -124.840 61.250 ;
        RECT 0.220 60.930 0.710 61.390 ;
        RECT 0.250 60.910 0.680 60.930 ;
        RECT 0.950 60.610 1.280 86.180 ;
        RECT 0.860 60.120 1.350 60.610 ;
        RECT 1.600 59.900 1.930 87.820 ;
        RECT -152.000 59.490 -124.840 59.500 ;
        RECT -152.160 59.140 -124.840 59.490 ;
        RECT 1.570 59.440 1.970 59.900 ;
        RECT -152.000 59.130 -124.840 59.140 ;
        RECT -151.050 58.780 -124.840 59.130 ;
        RECT -150.680 58.020 -124.840 58.780 ;
        RECT 1.360 58.950 1.940 59.060 ;
        RECT 2.270 58.950 2.600 89.390 ;
        RECT 2.910 63.530 3.240 94.560 ;
        RECT 2.910 59.070 3.230 63.530 ;
        RECT 3.520 59.680 3.850 96.040 ;
        RECT 4.140 59.930 4.470 97.590 ;
        RECT 4.770 60.960 5.100 99.170 ;
        RECT 5.370 61.260 5.700 104.650 ;
        RECT 5.950 61.830 6.280 106.210 ;
        RECT 6.560 62.860 6.890 107.750 ;
        RECT 7.150 63.470 7.480 109.310 ;
        RECT 7.790 64.140 8.120 109.890 ;
        RECT 8.410 64.790 8.740 111.490 ;
        RECT 9.010 65.420 9.340 112.980 ;
        RECT 9.640 66.030 9.970 114.700 ;
        RECT 11.030 113.620 11.440 113.950 ;
        RECT 11.030 111.870 11.440 112.200 ;
        RECT 11.030 110.120 11.440 110.450 ;
        RECT 11.030 109.320 11.440 109.650 ;
        RECT 11.030 107.570 11.440 107.900 ;
        RECT 11.030 105.820 11.440 106.150 ;
        RECT 11.030 104.070 11.440 104.400 ;
        RECT 11.770 103.790 12.010 115.870 ;
        RECT 14.610 115.800 15.020 116.940 ;
        RECT 16.930 116.510 17.240 116.520 ;
        RECT 16.930 116.240 17.250 116.510 ;
        RECT 17.970 116.280 18.290 116.580 ;
        RECT 16.950 116.230 17.240 116.240 ;
        RECT 13.190 114.480 13.540 114.770 ;
        RECT 13.190 114.460 13.390 114.480 ;
        RECT 13.190 112.730 13.540 113.020 ;
        RECT 13.190 112.710 13.390 112.730 ;
        RECT 13.190 110.980 13.540 111.270 ;
        RECT 13.190 110.960 13.390 110.980 ;
        RECT 13.190 108.790 13.390 108.810 ;
        RECT 13.190 108.500 13.540 108.790 ;
        RECT 13.190 107.040 13.390 107.060 ;
        RECT 13.190 106.750 13.540 107.040 ;
        RECT 13.190 105.290 13.390 105.310 ;
        RECT 13.190 105.000 13.540 105.290 ;
        RECT 14.710 103.860 15.020 115.800 ;
        RECT 15.270 115.480 15.550 115.810 ;
        RECT 16.930 114.760 17.240 114.770 ;
        RECT 16.930 114.490 17.250 114.760 ;
        RECT 17.970 114.530 18.290 114.830 ;
        RECT 16.950 114.480 17.240 114.490 ;
        RECT 15.270 113.730 15.550 114.060 ;
        RECT 16.930 113.010 17.240 113.020 ;
        RECT 16.930 112.740 17.250 113.010 ;
        RECT 17.970 112.780 18.290 113.080 ;
        RECT 16.950 112.730 17.240 112.740 ;
        RECT 15.270 111.980 15.550 112.310 ;
        RECT 16.930 111.260 17.240 111.270 ;
        RECT 16.930 110.990 17.250 111.260 ;
        RECT 17.970 111.030 18.290 111.330 ;
        RECT 16.950 110.980 17.240 110.990 ;
        RECT 15.270 110.230 15.550 110.560 ;
        RECT 15.270 109.210 15.550 109.540 ;
        RECT 16.950 108.780 17.240 108.790 ;
        RECT 16.930 108.510 17.250 108.780 ;
        RECT 16.930 108.500 17.240 108.510 ;
        RECT 17.970 108.440 18.290 108.740 ;
        RECT 15.270 107.460 15.550 107.790 ;
        RECT 16.950 107.030 17.240 107.040 ;
        RECT 16.930 106.760 17.250 107.030 ;
        RECT 16.930 106.750 17.240 106.760 ;
        RECT 17.970 106.690 18.290 106.990 ;
        RECT 15.270 105.710 15.550 106.040 ;
        RECT 16.950 105.280 17.240 105.290 ;
        RECT 16.930 105.010 17.250 105.280 ;
        RECT 16.930 105.000 17.240 105.010 ;
        RECT 17.970 104.940 18.290 105.240 ;
        RECT 15.270 103.960 15.550 104.290 ;
        RECT 11.670 102.830 12.010 103.790 ;
        RECT 13.190 103.540 13.390 103.560 ;
        RECT 13.190 103.250 13.540 103.540 ;
        RECT 14.610 102.830 15.020 103.860 ;
        RECT 16.950 103.530 17.240 103.540 ;
        RECT 16.930 103.260 17.250 103.530 ;
        RECT 16.930 103.250 17.240 103.260 ;
        RECT 17.970 103.190 18.290 103.490 ;
        RECT 11.670 99.700 11.910 102.830 ;
        RECT 14.610 99.700 14.920 102.830 ;
        RECT 11.030 99.190 11.440 99.520 ;
        RECT 11.670 99.420 12.010 99.700 ;
        RECT 11.030 97.440 11.440 97.770 ;
        RECT 11.030 95.690 11.440 96.020 ;
        RECT 11.030 93.940 11.440 94.270 ;
        RECT 11.770 93.660 12.010 99.420 ;
        RECT 14.610 99.350 15.020 99.700 ;
        RECT 13.190 98.660 13.390 98.680 ;
        RECT 13.190 98.370 13.540 98.660 ;
        RECT 13.190 96.910 13.390 96.930 ;
        RECT 13.190 96.620 13.540 96.910 ;
        RECT 13.190 95.160 13.390 95.180 ;
        RECT 13.190 94.870 13.540 95.160 ;
        RECT 14.710 93.730 15.020 99.350 ;
        RECT 15.270 99.080 15.550 99.410 ;
        RECT 16.950 98.650 17.240 98.660 ;
        RECT 16.930 98.380 17.250 98.650 ;
        RECT 16.930 98.370 17.240 98.380 ;
        RECT 17.970 98.310 18.290 98.610 ;
        RECT 15.270 97.330 15.550 97.660 ;
        RECT 16.950 96.900 17.240 96.910 ;
        RECT 16.930 96.630 17.250 96.900 ;
        RECT 16.930 96.620 17.240 96.630 ;
        RECT 17.970 96.560 18.290 96.860 ;
        RECT 15.270 95.580 15.550 95.910 ;
        RECT 16.950 95.150 17.240 95.160 ;
        RECT 16.930 94.880 17.250 95.150 ;
        RECT 16.930 94.870 17.240 94.880 ;
        RECT 17.970 94.810 18.290 95.110 ;
        RECT 15.270 93.830 15.550 94.160 ;
        RECT 10.990 90.130 11.400 90.460 ;
        RECT 11.670 89.890 12.010 93.660 ;
        RECT 13.190 93.410 13.390 93.430 ;
        RECT 13.190 93.120 13.540 93.410 ;
        RECT 14.610 89.890 15.020 93.730 ;
        RECT 16.950 93.400 17.240 93.410 ;
        RECT 16.930 93.130 17.250 93.400 ;
        RECT 16.930 93.120 17.240 93.130 ;
        RECT 17.970 93.060 18.290 93.360 ;
        RECT 19.040 90.640 19.330 123.420 ;
        RECT 20.230 122.430 20.730 122.870 ;
        RECT 20.500 109.700 20.690 122.430 ;
        RECT 20.220 109.210 20.690 109.700 ;
        RECT 21.080 109.560 21.450 109.580 ;
        RECT 21.030 109.300 21.450 109.560 ;
        RECT 21.080 109.290 21.450 109.300 ;
        RECT 20.040 108.770 20.360 109.050 ;
        RECT 20.500 108.950 20.690 109.210 ;
        RECT 20.500 108.660 20.730 108.950 ;
        RECT 20.500 107.890 20.690 108.660 ;
        RECT 20.040 107.500 20.360 107.780 ;
        RECT 20.500 107.600 20.730 107.890 ;
        RECT 20.500 107.340 20.690 107.600 ;
        RECT 20.220 106.850 20.690 107.340 ;
        RECT 21.080 107.250 21.450 107.260 ;
        RECT 21.030 106.990 21.450 107.250 ;
        RECT 21.080 106.970 21.450 106.990 ;
        RECT 20.500 106.500 20.690 106.850 ;
        RECT 20.220 106.010 20.690 106.500 ;
        RECT 21.080 106.360 21.450 106.380 ;
        RECT 21.030 106.100 21.450 106.360 ;
        RECT 21.080 106.090 21.450 106.100 ;
        RECT 20.040 105.570 20.360 105.850 ;
        RECT 20.500 105.750 20.690 106.010 ;
        RECT 20.500 105.460 20.730 105.750 ;
        RECT 20.500 104.690 20.690 105.460 ;
        RECT 20.040 104.300 20.360 104.580 ;
        RECT 20.500 104.400 20.730 104.690 ;
        RECT 20.500 104.140 20.690 104.400 ;
        RECT 20.220 103.650 20.690 104.140 ;
        RECT 21.080 104.050 21.450 104.060 ;
        RECT 21.030 103.790 21.450 104.050 ;
        RECT 21.080 103.770 21.450 103.790 ;
        RECT 20.500 99.880 20.690 103.650 ;
        RECT 21.810 99.980 22.040 109.920 ;
        RECT 24.780 109.700 25.030 123.420 ;
        RECT 26.480 123.380 27.210 130.210 ;
        RECT 31.630 130.100 32.610 130.250 ;
        RECT 26.640 113.030 26.810 123.380 ;
        RECT 31.640 122.850 32.610 130.100 ;
        RECT 44.250 129.110 47.480 132.100 ;
        RECT 52.430 131.630 61.030 132.350 ;
        RECT 72.140 132.100 76.090 133.640 ;
        RECT 85.070 133.290 85.630 133.790 ;
        RECT 85.080 133.070 85.630 133.290 ;
        RECT 81.770 132.720 81.960 132.730 ;
        RECT 88.900 132.720 89.620 139.040 ;
        RECT 90.370 139.770 104.660 140.330 ;
        RECT 115.590 140.160 116.120 141.060 ;
        RECT 117.230 141.000 119.600 141.630 ;
        RECT 90.370 135.470 113.720 139.770 ;
        RECT 117.260 139.040 118.210 141.000 ;
        RECT 118.960 140.980 119.540 141.000 ;
        RECT 129.340 140.340 133.250 141.800 ;
        RECT 140.570 141.150 144.700 141.550 ;
        RECT 140.570 141.060 144.710 141.150 ;
        RECT 119.630 140.330 133.250 140.340 ;
        RECT 114.490 138.350 115.060 138.360 ;
        RECT 90.370 135.190 104.660 135.470 ;
        RECT 100.750 133.640 104.660 135.190 ;
        RECT 114.490 134.930 115.110 138.350 ;
        RECT 114.490 134.920 115.060 134.930 ;
        RECT 81.770 132.370 89.620 132.720 ;
        RECT 44.260 129.080 47.450 129.110 ;
        RECT 37.030 125.010 38.500 125.540 ;
        RECT 31.620 122.380 32.630 122.850 ;
        RECT 34.660 122.400 35.100 122.900 ;
        RECT 28.860 118.650 29.200 118.940 ;
        RECT 28.910 118.620 29.170 118.650 ;
        RECT 27.030 115.090 27.290 115.410 ;
        RECT 26.490 112.730 26.810 113.030 ;
        RECT 26.650 112.400 26.810 112.730 ;
        RECT 26.650 111.850 26.920 112.400 ;
        RECT 26.640 111.800 26.920 111.850 ;
        RECT 26.640 111.710 26.810 111.800 ;
        RECT 23.540 109.540 23.880 109.590 ;
        RECT 23.540 109.520 24.100 109.540 ;
        RECT 23.420 109.350 24.100 109.520 ;
        RECT 23.540 109.310 24.100 109.350 ;
        RECT 23.540 109.270 23.880 109.310 ;
        RECT 24.780 108.630 25.420 109.700 ;
        RECT 24.780 107.920 25.030 108.630 ;
        RECT 26.650 108.340 26.810 111.710 ;
        RECT 27.060 111.590 27.250 115.090 ;
        RECT 28.930 112.680 29.140 118.620 ;
        RECT 32.500 118.020 32.760 118.030 ;
        RECT 32.480 117.720 32.780 118.020 ;
        RECT 32.500 117.710 32.760 117.720 ;
        RECT 29.330 116.690 29.670 117.010 ;
        RECT 28.460 112.230 28.770 112.670 ;
        RECT 28.920 112.390 29.150 112.680 ;
        RECT 27.030 111.560 27.250 111.590 ;
        RECT 27.020 111.290 27.270 111.560 ;
        RECT 27.020 111.280 27.260 111.290 ;
        RECT 27.030 111.040 27.260 111.280 ;
        RECT 27.060 109.010 27.220 111.040 ;
        RECT 28.060 110.700 28.380 111.020 ;
        RECT 28.930 110.690 29.140 112.390 ;
        RECT 29.400 112.120 29.590 116.690 ;
        RECT 29.770 114.600 30.060 114.920 ;
        RECT 29.390 111.830 29.620 112.120 ;
        RECT 27.410 110.190 27.650 110.610 ;
        RECT 28.920 110.400 29.150 110.690 ;
        RECT 28.930 110.260 29.140 110.400 ;
        RECT 27.380 109.870 27.650 110.190 ;
        RECT 27.410 109.440 27.650 109.870 ;
        RECT 29.400 109.800 29.590 111.830 ;
        RECT 29.810 110.330 30.020 114.600 ;
        RECT 30.810 114.120 31.150 114.440 ;
        RECT 29.780 109.820 30.020 110.330 ;
        RECT 28.950 109.620 29.140 109.750 ;
        RECT 28.930 109.330 29.160 109.620 ;
        RECT 29.390 109.510 29.620 109.800 ;
        RECT 28.050 109.010 28.370 109.330 ;
        RECT 27.030 108.770 27.260 109.010 ;
        RECT 27.020 108.760 27.260 108.770 ;
        RECT 27.020 108.490 27.270 108.760 ;
        RECT 27.030 108.460 27.250 108.490 ;
        RECT 26.640 108.250 26.810 108.340 ;
        RECT 26.640 108.200 26.920 108.250 ;
        RECT 23.540 107.240 23.880 107.280 ;
        RECT 23.540 107.200 24.100 107.240 ;
        RECT 23.420 107.030 24.100 107.200 ;
        RECT 23.540 107.010 24.100 107.030 ;
        RECT 23.540 106.960 23.880 107.010 ;
        RECT 24.780 106.850 25.420 107.920 ;
        RECT 26.650 107.650 26.920 108.200 ;
        RECT 26.650 107.020 26.810 107.650 ;
        RECT 27.060 107.020 27.250 108.460 ;
        RECT 28.460 107.380 28.770 107.820 ;
        RECT 28.950 107.710 29.140 109.330 ;
        RECT 29.400 108.220 29.590 109.510 ;
        RECT 29.380 107.930 29.610 108.220 ;
        RECT 28.950 107.500 29.180 107.710 ;
        RECT 28.940 107.420 29.180 107.500 ;
        RECT 26.540 106.970 26.820 107.020 ;
        RECT 27.060 107.000 27.260 107.020 ;
        RECT 28.940 107.000 29.170 107.420 ;
        RECT 29.400 107.000 29.590 107.930 ;
        RECT 29.810 107.000 30.020 109.820 ;
        RECT 30.890 108.520 31.070 114.120 ;
        RECT 31.610 111.050 31.870 111.840 ;
        RECT 30.830 108.180 31.120 108.520 ;
        RECT 30.890 107.000 31.070 108.180 ;
        RECT 31.610 108.110 31.870 108.900 ;
        RECT 32.530 107.480 32.730 117.710 ;
        RECT 32.510 107.350 32.730 107.480 ;
        RECT 34.760 107.350 34.990 122.400 ;
        RECT 35.660 118.630 35.940 118.950 ;
        RECT 35.220 117.720 35.500 118.040 ;
        RECT 32.460 107.020 32.790 107.350 ;
        RECT 34.710 107.050 35.030 107.350 ;
        RECT 24.780 106.500 25.030 106.850 ;
        RECT 26.540 106.690 26.860 106.970 ;
        RECT 23.540 106.340 23.880 106.390 ;
        RECT 23.540 106.320 24.100 106.340 ;
        RECT 23.420 106.150 24.100 106.320 ;
        RECT 23.540 106.110 24.100 106.150 ;
        RECT 23.540 106.070 23.880 106.110 ;
        RECT 24.780 105.430 25.420 106.500 ;
        RECT 26.540 106.370 26.820 106.690 ;
        RECT 26.540 105.770 26.930 106.370 ;
        RECT 24.780 104.720 25.030 105.430 ;
        RECT 23.540 104.040 23.880 104.080 ;
        RECT 23.540 104.000 24.100 104.040 ;
        RECT 23.420 103.830 24.100 104.000 ;
        RECT 23.540 103.810 24.100 103.830 ;
        RECT 23.540 103.760 23.880 103.810 ;
        RECT 24.780 103.650 25.420 104.720 ;
        RECT 24.780 99.990 25.030 103.650 ;
        RECT 20.480 99.380 20.690 99.880 ;
        RECT 21.790 99.570 22.040 99.980 ;
        RECT 24.760 99.570 25.030 99.990 ;
        RECT 26.540 102.220 26.820 105.770 ;
        RECT 27.070 105.560 27.260 107.000 ;
        RECT 28.470 106.200 28.780 106.640 ;
        RECT 33.550 105.810 33.780 107.020 ;
        RECT 34.760 107.000 35.000 107.050 ;
        RECT 34.770 106.050 35.000 107.000 ;
        RECT 35.250 106.180 35.470 117.720 ;
        RECT 35.240 106.110 35.470 106.180 ;
        RECT 27.040 105.530 27.260 105.560 ;
        RECT 27.030 105.260 27.280 105.530 ;
        RECT 27.030 105.250 27.270 105.260 ;
        RECT 27.040 105.010 27.270 105.250 ;
        RECT 28.310 105.240 28.630 105.560 ;
        RECT 33.520 105.020 33.780 105.810 ;
        RECT 34.760 105.800 35.000 106.050 ;
        RECT 27.070 102.980 27.230 105.010 ;
        RECT 27.420 104.450 27.660 104.580 ;
        RECT 27.400 104.130 27.660 104.450 ;
        RECT 27.400 103.530 27.660 103.850 ;
        RECT 27.420 103.410 27.660 103.530 ;
        RECT 27.040 102.740 27.270 102.980 ;
        RECT 33.550 102.870 33.780 105.020 ;
        RECT 27.030 102.730 27.270 102.740 ;
        RECT 27.030 102.460 27.280 102.730 ;
        RECT 28.310 102.480 28.630 102.800 ;
        RECT 27.040 102.430 27.260 102.460 ;
        RECT 26.540 101.620 26.930 102.220 ;
        RECT 26.540 100.140 26.820 101.620 ;
        RECT 27.070 100.560 27.260 102.430 ;
        RECT 33.520 102.080 33.780 102.870 ;
        RECT 28.470 101.350 28.780 101.790 ;
        RECT 29.070 100.720 29.460 100.740 ;
        RECT 29.060 100.630 29.460 100.720 ;
        RECT 28.910 100.620 29.460 100.630 ;
        RECT 27.070 100.370 28.670 100.560 ;
        RECT 26.540 99.860 28.260 100.140 ;
        RECT 28.060 99.630 28.260 99.860 ;
        RECT 20.480 99.230 20.670 99.380 ;
        RECT 20.200 98.740 20.670 99.230 ;
        RECT 21.060 99.090 21.430 99.110 ;
        RECT 21.010 98.830 21.430 99.090 ;
        RECT 21.060 98.820 21.430 98.830 ;
        RECT 20.020 98.300 20.340 98.580 ;
        RECT 20.480 98.480 20.670 98.740 ;
        RECT 20.480 98.190 20.710 98.480 ;
        RECT 20.480 97.420 20.670 98.190 ;
        RECT 20.020 97.030 20.340 97.310 ;
        RECT 20.480 97.130 20.710 97.420 ;
        RECT 20.480 96.870 20.670 97.130 ;
        RECT 20.200 96.380 20.670 96.870 ;
        RECT 21.060 96.780 21.430 96.790 ;
        RECT 21.010 96.520 21.430 96.780 ;
        RECT 21.060 96.500 21.430 96.520 ;
        RECT 20.480 96.030 20.670 96.380 ;
        RECT 20.200 95.540 20.670 96.030 ;
        RECT 21.060 95.890 21.430 95.910 ;
        RECT 21.010 95.630 21.430 95.890 ;
        RECT 21.060 95.620 21.430 95.630 ;
        RECT 20.020 95.100 20.340 95.380 ;
        RECT 20.480 95.280 20.670 95.540 ;
        RECT 20.480 94.990 20.710 95.280 ;
        RECT 20.480 94.220 20.670 94.990 ;
        RECT 20.020 93.830 20.340 94.110 ;
        RECT 20.480 93.930 20.710 94.220 ;
        RECT 20.480 93.710 20.670 93.930 ;
        RECT 21.790 93.750 22.020 99.570 ;
        RECT 24.760 99.230 25.010 99.570 ;
        RECT 28.070 99.370 28.230 99.630 ;
        RECT 27.920 99.230 28.230 99.370 ;
        RECT 23.520 99.070 23.860 99.120 ;
        RECT 23.520 99.050 24.080 99.070 ;
        RECT 23.400 98.880 24.080 99.050 ;
        RECT 23.520 98.840 24.080 98.880 ;
        RECT 23.520 98.800 23.860 98.840 ;
        RECT 24.760 98.160 25.400 99.230 ;
        RECT 27.910 99.080 28.230 99.230 ;
        RECT 28.070 98.790 28.230 99.080 ;
        RECT 28.070 98.240 28.340 98.790 ;
        RECT 28.060 98.190 28.340 98.240 ;
        RECT 28.480 98.450 28.670 100.370 ;
        RECT 28.880 100.380 29.460 100.620 ;
        RECT 28.880 100.360 29.450 100.380 ;
        RECT 28.880 100.350 29.070 100.360 ;
        RECT 28.880 99.510 29.050 100.350 ;
        RECT 33.550 100.290 33.780 102.080 ;
        RECT 34.770 103.910 35.000 105.800 ;
        RECT 35.230 105.510 35.430 106.110 ;
        RECT 35.680 105.970 35.910 118.630 ;
        RECT 37.050 112.900 37.470 125.010 ;
        RECT 38.080 112.900 38.500 125.010 ;
        RECT 40.460 122.360 40.900 122.860 ;
        RECT 40.560 115.380 40.790 122.360 ;
        RECT 44.980 117.110 46.260 129.080 ;
        RECT 48.740 123.890 49.020 124.010 ;
        RECT 48.740 123.390 49.070 123.890 ;
        RECT 44.980 117.030 46.280 117.110 ;
        RECT 44.970 116.730 46.280 117.030 ;
        RECT 41.750 116.080 42.050 116.400 ;
        RECT 40.430 115.370 40.790 115.380 ;
        RECT 40.400 114.480 40.790 115.370 ;
        RECT 37.050 112.760 38.500 112.900 ;
        RECT 37.050 107.020 37.470 112.760 ;
        RECT 38.080 107.020 38.500 112.760 ;
        RECT 40.560 107.350 40.790 114.480 ;
        RECT 41.780 111.840 42.010 116.080 ;
        RECT 48.060 115.530 48.490 115.870 ;
        RECT 46.780 112.230 47.090 112.670 ;
        RECT 41.780 111.050 42.040 111.840 ;
        RECT 48.300 111.590 48.490 115.530 ;
        RECT 48.740 113.030 49.020 123.390 ;
        RECT 50.440 118.630 50.700 118.950 ;
        RECT 49.550 117.760 49.810 118.080 ;
        RECT 49.580 114.040 49.770 117.760 ;
        RECT 50.460 114.040 50.680 118.630 ;
        RECT 52.430 115.410 52.770 131.630 ;
        RECT 72.840 130.230 76.070 132.100 ;
        RECT 81.770 130.430 81.960 132.370 ;
        RECT 100.730 132.180 104.680 133.640 ;
        RECT 113.660 133.290 114.220 133.790 ;
        RECT 117.490 133.370 118.210 139.040 ;
        RECT 118.960 139.770 133.250 140.330 ;
        RECT 144.180 140.160 144.710 141.060 ;
        RECT 145.820 141.000 148.190 141.630 ;
        RECT 118.960 135.470 142.310 139.770 ;
        RECT 145.850 139.040 146.800 141.000 ;
        RECT 147.550 140.980 148.130 141.000 ;
        RECT 157.930 140.340 161.840 141.800 ;
        RECT 169.160 141.150 173.290 141.550 ;
        RECT 169.160 141.060 173.300 141.150 ;
        RECT 148.220 140.330 161.840 140.340 ;
        RECT 143.080 138.350 143.650 138.360 ;
        RECT 118.960 135.190 133.250 135.470 ;
        RECT 129.340 133.640 133.250 135.190 ;
        RECT 143.080 134.930 143.700 138.350 ;
        RECT 143.080 134.920 143.650 134.930 ;
        RECT 113.670 133.070 114.220 133.290 ;
        RECT 129.320 132.870 133.270 133.640 ;
        RECT 142.250 133.290 142.810 133.790 ;
        RECT 146.080 133.370 146.800 139.040 ;
        RECT 147.550 139.770 161.840 140.330 ;
        RECT 172.770 140.160 173.300 141.060 ;
        RECT 174.410 141.000 176.780 141.630 ;
        RECT 147.550 135.470 170.900 139.770 ;
        RECT 174.440 139.040 175.390 141.000 ;
        RECT 176.140 140.980 176.720 141.000 ;
        RECT 186.520 140.340 190.430 141.800 ;
        RECT 197.750 141.150 201.880 141.550 ;
        RECT 197.750 141.060 201.890 141.150 ;
        RECT 176.810 140.330 190.430 140.340 ;
        RECT 171.670 138.350 172.240 138.360 ;
        RECT 147.550 135.190 161.840 135.470 ;
        RECT 157.930 133.640 161.840 135.190 ;
        RECT 171.670 134.930 172.290 138.350 ;
        RECT 171.670 134.920 172.240 134.930 ;
        RECT 142.260 133.070 142.810 133.290 ;
        RECT 100.670 132.100 104.680 132.180 ;
        RECT 129.330 132.100 133.280 132.870 ;
        RECT 157.910 132.100 161.860 133.640 ;
        RECT 170.840 133.290 171.400 133.790 ;
        RECT 174.670 133.370 175.390 139.040 ;
        RECT 176.140 139.770 190.430 140.330 ;
        RECT 201.360 140.160 201.890 141.060 ;
        RECT 176.140 135.470 199.490 139.770 ;
        RECT 200.260 138.350 200.830 138.360 ;
        RECT 176.140 135.190 190.430 135.470 ;
        RECT 186.520 133.640 190.430 135.190 ;
        RECT 200.260 134.930 200.880 138.350 ;
        RECT 200.260 134.920 200.830 134.930 ;
        RECT 170.850 133.070 171.400 133.290 ;
        RECT 186.500 132.100 190.450 133.640 ;
        RECT 199.430 133.290 199.990 133.790 ;
        RECT 199.440 133.070 199.990 133.290 ;
        RECT 100.670 131.900 104.660 132.100 ;
        RECT 100.650 131.700 104.660 131.900 ;
        RECT 81.770 130.240 81.980 130.430 ;
        RECT 72.830 129.110 76.070 130.230 ;
        RECT 56.930 128.170 57.300 128.180 ;
        RECT 56.880 127.720 57.380 128.170 ;
        RECT 53.080 119.310 53.400 119.680 ;
        RECT 52.380 115.330 52.770 115.410 ;
        RECT 52.370 114.560 52.770 115.330 ;
        RECT 52.380 114.490 52.770 114.560 ;
        RECT 49.410 113.350 50.090 114.040 ;
        RECT 50.450 113.350 51.130 114.040 ;
        RECT 48.740 112.730 49.080 113.030 ;
        RECT 48.740 112.400 49.020 112.730 ;
        RECT 50.490 112.710 50.810 113.030 ;
        RECT 51.470 112.460 51.790 112.780 ;
        RECT 48.630 111.800 49.020 112.400 ;
        RECT 50.640 111.880 50.960 112.200 ;
        RECT 51.420 111.810 51.740 112.130 ;
        RECT 46.930 111.270 47.250 111.590 ;
        RECT 48.300 111.560 48.520 111.590 ;
        RECT 48.280 111.290 48.530 111.560 ;
        RECT 48.290 111.280 48.530 111.290 ;
        RECT 41.780 108.900 42.010 111.050 ;
        RECT 48.290 111.040 48.520 111.280 ;
        RECT 47.900 110.480 48.140 110.610 ;
        RECT 47.900 110.160 48.160 110.480 ;
        RECT 47.900 109.560 48.160 109.880 ;
        RECT 47.900 109.440 48.140 109.560 ;
        RECT 48.330 109.010 48.490 111.040 ;
        RECT 48.740 110.200 49.020 111.800 ;
        RECT 49.530 111.350 49.850 111.670 ;
        RECT 50.750 111.190 50.960 111.300 ;
        RECT 50.730 110.870 50.990 111.190 ;
        RECT 51.420 110.960 51.740 111.280 ;
        RECT 48.740 109.880 49.100 110.200 ;
        RECT 50.260 110.070 50.580 110.390 ;
        RECT 41.780 108.110 42.040 108.900 ;
        RECT 46.930 108.510 47.250 108.830 ;
        RECT 48.290 108.770 48.520 109.010 ;
        RECT 48.290 108.760 48.530 108.770 ;
        RECT 48.280 108.490 48.530 108.760 ;
        RECT 48.300 108.460 48.520 108.490 ;
        RECT 40.510 107.050 40.830 107.350 ;
        RECT 37.050 107.000 38.500 107.020 ;
        RECT 35.570 105.660 35.910 105.970 ;
        RECT 37.060 106.860 38.500 107.000 ;
        RECT 35.570 105.650 35.890 105.660 ;
        RECT 35.240 105.480 35.470 105.510 ;
        RECT 34.770 103.610 35.100 103.910 ;
        RECT 34.770 103.440 35.020 103.610 ;
        RECT 34.770 100.320 35.000 103.440 ;
        RECT 35.250 102.280 35.470 105.480 ;
        RECT 35.250 101.970 35.920 102.280 ;
        RECT 35.600 101.960 35.920 101.970 ;
        RECT 37.060 100.980 37.480 106.860 ;
        RECT 33.030 100.220 33.780 100.290 ;
        RECT 33.000 100.060 33.780 100.220 ;
        RECT 34.750 100.260 35.000 100.320 ;
        RECT 38.080 100.390 38.500 106.860 ;
        RECT 40.560 103.860 40.790 107.050 ;
        RECT 41.780 105.810 42.010 108.110 ;
        RECT 46.780 107.380 47.090 107.820 ;
        RECT 46.780 106.200 47.090 106.640 ;
        RECT 41.780 105.020 42.040 105.810 ;
        RECT 48.300 105.560 48.490 108.460 ;
        RECT 48.740 108.250 49.020 109.880 ;
        RECT 50.750 109.580 50.960 110.870 ;
        RECT 51.470 110.310 51.790 110.630 ;
        RECT 50.730 109.290 50.960 109.580 ;
        RECT 51.470 109.460 51.790 109.780 ;
        RECT 51.420 108.810 51.740 109.130 ;
        RECT 48.630 107.650 49.020 108.250 ;
        RECT 51.420 107.960 51.740 108.280 ;
        RECT 48.740 106.970 49.020 107.650 ;
        RECT 50.900 107.200 51.220 107.500 ;
        RECT 51.470 107.310 51.790 107.630 ;
        RECT 52.430 107.200 52.770 114.490 ;
        RECT 53.100 113.930 53.370 119.310 ;
        RECT 53.100 113.430 53.780 113.930 ;
        RECT 53.100 113.050 53.370 113.430 ;
        RECT 53.090 112.900 53.370 113.050 ;
        RECT 50.900 107.170 51.330 107.200 ;
        RECT 51.930 107.170 52.770 107.200 ;
        RECT 50.900 107.140 52.770 107.170 ;
        RECT 51.050 107.090 52.770 107.140 ;
        RECT 51.080 107.060 52.770 107.090 ;
        RECT 51.110 107.040 52.770 107.060 ;
        RECT 51.180 107.030 52.140 107.040 ;
        RECT 48.740 106.670 49.060 106.970 ;
        RECT 50.490 106.680 50.810 107.000 ;
        RECT 48.740 106.370 49.020 106.670 ;
        RECT 51.470 106.430 51.790 106.750 ;
        RECT 48.630 105.770 49.020 106.370 ;
        RECT 50.640 105.850 50.960 106.170 ;
        RECT 51.420 105.780 51.740 106.100 ;
        RECT 46.930 105.240 47.250 105.560 ;
        RECT 48.300 105.530 48.520 105.560 ;
        RECT 48.280 105.260 48.530 105.530 ;
        RECT 48.290 105.250 48.530 105.260 ;
        RECT 40.480 103.540 40.800 103.860 ;
        RECT 40.560 101.330 40.790 103.540 ;
        RECT 41.780 102.870 42.010 105.020 ;
        RECT 48.290 105.010 48.520 105.250 ;
        RECT 47.900 104.450 48.140 104.580 ;
        RECT 47.900 104.130 48.160 104.450 ;
        RECT 47.900 103.530 48.160 103.850 ;
        RECT 47.900 103.410 48.140 103.530 ;
        RECT 48.330 102.980 48.490 105.010 ;
        RECT 48.740 104.170 49.020 105.770 ;
        RECT 49.530 105.320 49.850 105.640 ;
        RECT 50.750 105.160 50.960 105.270 ;
        RECT 50.730 104.840 50.990 105.160 ;
        RECT 51.420 104.930 51.740 105.250 ;
        RECT 48.740 103.850 49.100 104.170 ;
        RECT 50.260 104.040 50.580 104.360 ;
        RECT 41.780 102.080 42.040 102.870 ;
        RECT 46.930 102.480 47.250 102.800 ;
        RECT 48.290 102.740 48.520 102.980 ;
        RECT 48.290 102.730 48.530 102.740 ;
        RECT 48.280 102.460 48.530 102.730 ;
        RECT 48.300 102.430 48.520 102.460 ;
        RECT 40.480 101.030 40.800 101.330 ;
        RECT 33.000 99.610 33.410 100.060 ;
        RECT 28.880 98.760 29.040 99.510 ;
        RECT 28.840 98.740 29.040 98.760 ;
        RECT 29.860 98.750 30.180 99.070 ;
        RECT 28.830 98.500 29.060 98.740 ;
        RECT 28.830 98.450 29.040 98.500 ;
        RECT 28.480 98.330 28.650 98.450 ;
        RECT 24.760 97.450 25.010 98.160 ;
        RECT 28.060 98.100 28.230 98.190 ;
        RECT 28.070 97.630 28.230 98.100 ;
        RECT 28.060 97.540 28.230 97.630 ;
        RECT 28.060 97.490 28.340 97.540 ;
        RECT 23.520 96.770 23.860 96.810 ;
        RECT 23.520 96.730 24.080 96.770 ;
        RECT 23.400 96.560 24.080 96.730 ;
        RECT 23.520 96.540 24.080 96.560 ;
        RECT 23.520 96.490 23.860 96.540 ;
        RECT 24.760 96.380 25.400 97.450 ;
        RECT 28.070 96.940 28.340 97.490 ;
        RECT 28.480 97.400 28.640 98.330 ;
        RECT 28.480 97.280 28.650 97.400 ;
        RECT 28.880 97.280 29.040 98.450 ;
        RECT 29.860 98.200 30.180 98.520 ;
        RECT 30.820 98.110 31.060 99.500 ;
        RECT 24.760 96.030 25.010 96.380 ;
        RECT 23.520 95.870 23.860 95.920 ;
        RECT 23.520 95.850 24.080 95.870 ;
        RECT 23.400 95.680 24.080 95.850 ;
        RECT 23.520 95.640 24.080 95.680 ;
        RECT 23.520 95.600 23.860 95.640 ;
        RECT 24.760 94.960 25.400 96.030 ;
        RECT 28.070 95.550 28.230 96.940 ;
        RECT 28.480 96.360 28.670 97.280 ;
        RECT 28.830 97.230 29.040 97.280 ;
        RECT 28.830 96.990 29.060 97.230 ;
        RECT 29.860 97.210 30.180 97.530 ;
        RECT 30.810 97.450 31.080 98.110 ;
        RECT 28.840 96.970 29.040 96.990 ;
        RECT 28.450 96.340 28.690 96.360 ;
        RECT 28.880 96.340 29.040 96.970 ;
        RECT 29.860 96.660 30.180 96.980 ;
        RECT 28.450 96.150 29.040 96.340 ;
        RECT 28.450 96.130 28.690 96.150 ;
        RECT 28.070 95.000 28.340 95.550 ;
        RECT 24.760 94.250 25.010 94.960 ;
        RECT 28.060 94.950 28.340 95.000 ;
        RECT 28.480 95.210 28.670 96.130 ;
        RECT 28.880 95.520 29.040 96.150 ;
        RECT 28.840 95.500 29.040 95.520 ;
        RECT 29.860 95.510 30.180 95.830 ;
        RECT 28.830 95.260 29.060 95.500 ;
        RECT 28.830 95.210 29.040 95.260 ;
        RECT 28.480 95.090 28.650 95.210 ;
        RECT 28.060 94.860 28.230 94.950 ;
        RECT 28.070 94.400 28.230 94.860 ;
        RECT 28.060 94.310 28.230 94.400 ;
        RECT 28.060 94.260 28.340 94.310 ;
        RECT 20.480 93.670 20.690 93.710 ;
        RECT 20.200 93.180 20.690 93.670 ;
        RECT 21.060 93.580 21.430 93.590 ;
        RECT 21.010 93.320 21.430 93.580 ;
        RECT 21.060 93.300 21.430 93.320 ;
        RECT 20.480 92.960 20.690 93.180 ;
        RECT 21.790 92.960 22.040 93.750 ;
        RECT 23.520 93.570 23.860 93.610 ;
        RECT 23.520 93.530 24.080 93.570 ;
        RECT 23.400 93.360 24.080 93.530 ;
        RECT 23.520 93.340 24.080 93.360 ;
        RECT 23.520 93.290 23.860 93.340 ;
        RECT 24.760 93.180 25.400 94.250 ;
        RECT 28.070 93.710 28.340 94.260 ;
        RECT 28.480 94.170 28.640 95.090 ;
        RECT 28.480 94.050 28.650 94.170 ;
        RECT 28.880 94.050 29.040 95.210 ;
        RECT 29.860 94.960 30.180 95.280 ;
        RECT 30.820 94.860 31.060 97.450 ;
        RECT 33.000 97.350 33.380 99.610 ;
        RECT 34.750 98.090 34.990 100.260 ;
        RECT 38.080 100.210 38.510 100.390 ;
        RECT 38.080 99.820 38.520 100.210 ;
        RECT 40.560 100.000 40.790 101.030 ;
        RECT 38.110 99.610 38.520 99.820 ;
        RECT 37.030 99.130 37.430 99.500 ;
        RECT 38.110 99.130 38.510 99.610 ;
        RECT 37.030 98.910 38.510 99.130 ;
        RECT 34.740 97.430 35.000 98.090 ;
        RECT 33.000 95.490 33.390 97.350 ;
        RECT 30.810 94.540 31.070 94.860 ;
        RECT 24.760 92.960 25.030 93.180 ;
        RECT 28.070 93.010 28.260 93.710 ;
        RECT 28.480 93.060 28.670 94.050 ;
        RECT 28.830 94.000 29.040 94.050 ;
        RECT 28.830 93.760 29.060 94.000 ;
        RECT 29.860 93.980 30.180 94.300 ;
        RECT 30.820 93.860 31.060 94.540 ;
        RECT 33.000 94.000 33.380 95.490 ;
        RECT 34.750 94.820 34.990 97.430 ;
        RECT 34.740 94.500 35.000 94.820 ;
        RECT 28.840 93.740 29.040 93.760 ;
        RECT 28.880 93.010 29.040 93.740 ;
        RECT 29.860 93.430 30.180 93.750 ;
        RECT 15.230 90.020 15.510 90.350 ;
        RECT 11.730 89.650 12.010 89.890 ;
        RECT 10.990 88.380 11.400 88.710 ;
        RECT 10.990 86.630 11.400 86.960 ;
        RECT 10.990 84.880 11.400 85.210 ;
        RECT 11.730 83.890 11.970 89.650 ;
        RECT 14.670 89.620 15.020 89.890 ;
        RECT 19.000 89.890 19.330 90.640 ;
        RECT 20.500 90.180 20.690 92.960 ;
        RECT 21.810 92.670 22.040 92.960 ;
        RECT 21.720 92.190 22.050 92.670 ;
        RECT 21.810 90.180 22.040 92.190 ;
        RECT 24.780 90.180 25.030 92.960 ;
        RECT 20.500 89.960 20.700 90.180 ;
        RECT 13.150 89.600 13.350 89.620 ;
        RECT 13.150 89.310 13.500 89.600 ;
        RECT 13.150 87.850 13.350 87.870 ;
        RECT 13.150 87.560 13.500 87.850 ;
        RECT 13.150 86.100 13.350 86.120 ;
        RECT 13.150 85.810 13.500 86.100 ;
        RECT 13.150 84.350 13.350 84.370 ;
        RECT 13.150 84.060 13.500 84.350 ;
        RECT 14.670 83.960 14.980 89.620 ;
        RECT 16.910 89.590 17.200 89.600 ;
        RECT 16.890 89.320 17.210 89.590 ;
        RECT 16.890 89.310 17.200 89.320 ;
        RECT 17.930 89.250 18.250 89.550 ;
        RECT 15.230 88.270 15.510 88.600 ;
        RECT 16.910 87.840 17.200 87.850 ;
        RECT 16.890 87.570 17.210 87.840 ;
        RECT 16.890 87.560 17.200 87.570 ;
        RECT 17.930 87.500 18.250 87.800 ;
        RECT 15.230 86.520 15.510 86.850 ;
        RECT 16.910 86.090 17.200 86.100 ;
        RECT 16.890 85.820 17.210 86.090 ;
        RECT 16.890 85.810 17.200 85.820 ;
        RECT 17.930 85.750 18.250 86.050 ;
        RECT 15.230 84.770 15.510 85.100 ;
        RECT 16.910 84.340 17.200 84.350 ;
        RECT 16.890 84.070 17.210 84.340 ;
        RECT 16.890 84.060 17.200 84.070 ;
        RECT 17.930 84.000 18.250 84.300 ;
        RECT 11.670 83.640 11.970 83.890 ;
        RECT 14.610 83.640 14.980 83.960 ;
        RECT 19.000 83.940 19.290 89.890 ;
        RECT 20.230 89.470 20.700 89.960 ;
        RECT 21.090 89.820 21.460 89.840 ;
        RECT 21.040 89.560 21.460 89.820 ;
        RECT 21.810 89.580 22.050 90.180 ;
        RECT 24.780 89.960 25.040 90.180 ;
        RECT 23.550 89.800 23.890 89.850 ;
        RECT 23.550 89.780 24.110 89.800 ;
        RECT 24.780 89.790 25.430 89.960 ;
        RECT 23.430 89.610 24.110 89.780 ;
        RECT 21.090 89.550 21.460 89.560 ;
        RECT 20.050 89.030 20.370 89.310 ;
        RECT 20.510 89.210 20.700 89.470 ;
        RECT 20.510 88.920 20.740 89.210 ;
        RECT 20.510 88.150 20.700 88.920 ;
        RECT 20.050 87.760 20.370 88.040 ;
        RECT 20.510 87.860 20.740 88.150 ;
        RECT 20.510 87.600 20.700 87.860 ;
        RECT 20.230 87.110 20.700 87.600 ;
        RECT 21.090 87.510 21.460 87.520 ;
        RECT 21.040 87.250 21.460 87.510 ;
        RECT 21.090 87.230 21.460 87.250 ;
        RECT 20.510 86.760 20.700 87.110 ;
        RECT 20.230 86.270 20.700 86.760 ;
        RECT 21.090 86.620 21.460 86.640 ;
        RECT 21.040 86.360 21.460 86.620 ;
        RECT 21.090 86.350 21.460 86.360 ;
        RECT 20.050 85.830 20.370 86.110 ;
        RECT 20.510 86.010 20.700 86.270 ;
        RECT 20.510 85.720 20.740 86.010 ;
        RECT 20.510 84.950 20.700 85.720 ;
        RECT 20.050 84.560 20.370 84.840 ;
        RECT 20.510 84.660 20.740 84.950 ;
        RECT 20.510 84.400 20.700 84.660 ;
        RECT 19.000 83.640 19.330 83.940 ;
        RECT 20.230 83.910 20.700 84.400 ;
        RECT 21.090 84.310 21.460 84.320 ;
        RECT 21.040 84.050 21.460 84.310 ;
        RECT 21.090 84.030 21.460 84.050 ;
        RECT 20.500 83.690 20.700 83.910 ;
        RECT 21.820 83.690 22.050 89.580 ;
        RECT 23.550 89.570 24.110 89.610 ;
        RECT 23.550 89.530 23.890 89.570 ;
        RECT 24.790 88.890 25.430 89.790 ;
        RECT 28.100 89.460 28.260 93.010 ;
        RECT 30.820 93.000 31.090 93.860 ;
        RECT 33.000 93.000 33.410 94.000 ;
        RECT 34.750 93.860 34.990 94.500 ;
        RECT 37.030 94.020 37.430 98.910 ;
        RECT 34.750 93.000 35.020 93.860 ;
        RECT 37.030 93.000 37.460 94.020 ;
        RECT 38.110 93.000 38.510 98.910 ;
        RECT 40.550 98.090 40.790 100.000 ;
        RECT 41.780 100.310 42.010 102.080 ;
        RECT 46.780 101.350 47.090 101.790 ;
        RECT 41.780 99.930 42.540 100.310 ;
        RECT 48.300 100.180 48.490 102.430 ;
        RECT 48.740 102.220 49.020 103.850 ;
        RECT 50.750 103.550 50.960 104.840 ;
        RECT 51.470 104.280 51.790 104.600 ;
        RECT 50.730 103.260 50.960 103.550 ;
        RECT 51.470 103.430 51.790 103.750 ;
        RECT 51.420 102.780 51.740 103.100 ;
        RECT 48.630 101.620 49.020 102.220 ;
        RECT 51.420 101.930 51.740 102.250 ;
        RECT 40.540 97.430 40.800 98.090 ;
        RECT 40.550 94.820 40.790 97.430 ;
        RECT 42.160 97.350 42.540 99.930 ;
        RECT 46.470 99.810 46.750 100.130 ;
        RECT 46.900 99.990 48.490 100.180 ;
        RECT 44.480 98.110 44.720 99.500 ;
        RECT 45.360 98.750 45.680 99.070 ;
        RECT 46.500 98.760 46.660 99.810 ;
        RECT 46.900 99.660 47.090 99.990 ;
        RECT 48.740 99.800 49.020 101.620 ;
        RECT 50.920 101.170 51.250 101.460 ;
        RECT 51.470 101.280 51.790 101.600 ;
        RECT 52.430 101.170 52.770 107.040 ;
        RECT 53.100 111.470 53.370 112.900 ;
        RECT 53.720 112.480 54.040 112.800 ;
        RECT 53.100 111.180 53.380 111.470 ;
        RECT 53.100 108.880 53.370 111.180 ;
        RECT 53.770 110.260 54.090 110.580 ;
        RECT 53.760 109.540 54.080 109.860 ;
        RECT 53.100 108.590 53.380 108.880 ;
        RECT 53.100 107.020 53.370 108.590 ;
        RECT 53.680 107.290 54.000 107.610 ;
        RECT 53.090 106.870 53.370 107.020 ;
        RECT 50.910 101.140 51.330 101.170 ;
        RECT 51.930 101.140 52.770 101.170 ;
        RECT 50.910 101.030 52.770 101.140 ;
        RECT 51.190 101.000 52.090 101.030 ;
        RECT 52.430 100.970 52.770 101.030 ;
        RECT 53.100 105.440 53.370 106.870 ;
        RECT 53.720 106.450 54.040 106.770 ;
        RECT 53.100 105.150 53.380 105.440 ;
        RECT 53.100 102.850 53.370 105.150 ;
        RECT 53.770 104.230 54.090 104.550 ;
        RECT 53.760 103.510 54.080 103.830 ;
        RECT 53.100 102.560 53.380 102.850 ;
        RECT 53.100 100.970 53.370 102.560 ;
        RECT 53.680 101.260 54.000 101.580 ;
        RECT 56.930 100.810 57.300 127.720 ;
        RECT 57.720 124.270 58.180 124.700 ;
        RECT 56.900 100.350 57.350 100.810 ;
        RECT 56.930 100.310 57.300 100.350 ;
        RECT 57.740 100.220 58.110 124.270 ;
        RECT 58.490 119.560 58.940 119.990 ;
        RECT 47.350 99.790 49.020 99.800 ;
        RECT 46.870 99.550 47.090 99.660 ;
        RECT 46.500 98.740 46.700 98.760 ;
        RECT 45.360 98.200 45.680 98.520 ;
        RECT 46.480 98.500 46.710 98.740 ;
        RECT 46.500 98.450 46.710 98.500 ;
        RECT 46.870 98.450 47.060 99.550 ;
        RECT 47.310 99.520 49.020 99.790 ;
        RECT 57.710 99.760 58.150 100.220 ;
        RECT 57.740 99.710 58.110 99.760 ;
        RECT 47.310 99.380 47.470 99.520 ;
        RECT 47.310 99.100 47.640 99.380 ;
        RECT 47.310 98.790 47.470 99.100 ;
        RECT 44.460 97.450 44.730 98.110 ;
        RECT 42.150 95.490 42.540 97.350 ;
        RECT 40.540 94.500 40.800 94.820 ;
        RECT 40.550 93.860 40.790 94.500 ;
        RECT 40.550 93.000 40.820 93.860 ;
        RECT 42.160 93.000 42.540 95.490 ;
        RECT 44.480 94.860 44.720 97.450 ;
        RECT 45.360 97.210 45.680 97.530 ;
        RECT 46.500 97.280 46.660 98.450 ;
        RECT 46.890 98.330 47.060 98.450 ;
        RECT 46.900 97.400 47.060 98.330 ;
        RECT 47.200 98.240 47.470 98.790 ;
        RECT 47.200 98.190 47.480 98.240 ;
        RECT 47.310 98.100 47.480 98.190 ;
        RECT 47.310 97.630 47.470 98.100 ;
        RECT 58.510 97.870 58.880 119.560 ;
        RECT 65.060 118.510 65.640 119.070 ;
        RECT 61.850 116.940 62.410 117.590 ;
        RECT 62.800 117.430 63.360 118.010 ;
        RECT 63.880 117.890 64.440 118.480 ;
        RECT 59.380 114.480 59.810 114.920 ;
        RECT 58.480 97.860 58.880 97.870 ;
        RECT 47.310 97.540 47.480 97.630 ;
        RECT 46.890 97.280 47.060 97.400 ;
        RECT 46.500 97.230 46.710 97.280 ;
        RECT 46.480 96.990 46.710 97.230 ;
        RECT 45.360 96.660 45.680 96.980 ;
        RECT 46.500 96.970 46.700 96.990 ;
        RECT 46.500 96.340 46.660 96.970 ;
        RECT 46.870 96.360 47.060 97.280 ;
        RECT 47.200 97.490 47.480 97.540 ;
        RECT 47.200 96.940 47.470 97.490 ;
        RECT 58.470 97.440 58.890 97.860 ;
        RECT 58.510 97.430 58.880 97.440 ;
        RECT 46.850 96.340 47.090 96.360 ;
        RECT 46.500 96.150 47.090 96.340 ;
        RECT 45.360 95.510 45.680 95.830 ;
        RECT 46.500 95.520 46.660 96.150 ;
        RECT 46.850 96.130 47.090 96.150 ;
        RECT 46.500 95.500 46.700 95.520 ;
        RECT 45.360 94.960 45.680 95.280 ;
        RECT 46.480 95.260 46.710 95.500 ;
        RECT 46.500 95.210 46.710 95.260 ;
        RECT 46.870 95.210 47.060 96.130 ;
        RECT 47.310 95.550 47.470 96.940 ;
        RECT 44.470 94.540 44.730 94.860 ;
        RECT 44.480 93.000 44.720 94.540 ;
        RECT 45.360 93.980 45.680 94.300 ;
        RECT 46.500 94.050 46.660 95.210 ;
        RECT 46.890 95.090 47.060 95.210 ;
        RECT 46.900 94.170 47.060 95.090 ;
        RECT 47.200 95.000 47.470 95.550 ;
        RECT 47.200 94.950 47.480 95.000 ;
        RECT 47.310 94.860 47.480 94.950 ;
        RECT 47.310 94.400 47.470 94.860 ;
        RECT 47.310 94.310 47.480 94.400 ;
        RECT 46.890 94.050 47.060 94.170 ;
        RECT 46.500 94.000 46.710 94.050 ;
        RECT 46.480 93.760 46.710 94.000 ;
        RECT 45.360 93.430 45.680 93.750 ;
        RECT 46.500 93.740 46.700 93.760 ;
        RECT 46.500 93.010 46.660 93.740 ;
        RECT 46.870 93.060 47.060 94.050 ;
        RECT 47.200 94.260 47.480 94.310 ;
        RECT 47.200 93.710 47.470 94.260 ;
        RECT 47.310 93.010 47.470 93.710 ;
        RECT 30.850 90.170 31.090 93.000 ;
        RECT 28.100 88.910 28.370 89.460 ;
        RECT 24.790 88.180 25.040 88.890 ;
        RECT 28.090 88.860 28.370 88.910 ;
        RECT 28.510 89.120 28.700 90.110 ;
        RECT 28.910 89.430 29.070 90.160 ;
        RECT 30.850 90.140 31.220 90.170 ;
        RECT 30.830 89.890 31.220 90.140 ;
        RECT 28.870 89.410 29.070 89.430 ;
        RECT 29.890 89.420 30.210 89.740 ;
        RECT 28.860 89.170 29.090 89.410 ;
        RECT 30.530 89.320 30.790 89.640 ;
        RECT 28.860 89.120 29.070 89.170 ;
        RECT 28.510 89.000 28.680 89.120 ;
        RECT 26.130 88.460 26.450 88.800 ;
        RECT 28.090 88.770 28.260 88.860 ;
        RECT 23.550 87.500 23.890 87.540 ;
        RECT 23.550 87.460 24.110 87.500 ;
        RECT 23.430 87.290 24.110 87.460 ;
        RECT 23.550 87.270 24.110 87.290 ;
        RECT 23.550 87.220 23.890 87.270 ;
        RECT 24.790 87.110 25.430 88.180 ;
        RECT 24.790 86.760 25.040 87.110 ;
        RECT 23.550 86.600 23.890 86.650 ;
        RECT 23.550 86.580 24.110 86.600 ;
        RECT 23.430 86.410 24.110 86.580 ;
        RECT 23.550 86.370 24.110 86.410 ;
        RECT 23.550 86.330 23.890 86.370 ;
        RECT 24.790 85.690 25.430 86.760 ;
        RECT 24.790 84.980 25.040 85.690 ;
        RECT 23.550 84.300 23.890 84.340 ;
        RECT 23.550 84.260 24.110 84.300 ;
        RECT 23.430 84.090 24.110 84.260 ;
        RECT 23.550 84.070 24.110 84.090 ;
        RECT 23.550 84.020 23.890 84.070 ;
        RECT 24.790 84.010 25.430 84.980 ;
        RECT 24.780 83.910 25.430 84.010 ;
        RECT 24.780 83.690 25.040 83.910 ;
        RECT 26.210 83.700 26.420 88.460 ;
        RECT 28.100 88.320 28.260 88.770 ;
        RECT 28.090 88.230 28.260 88.320 ;
        RECT 28.090 88.180 28.370 88.230 ;
        RECT 27.240 87.970 27.500 88.090 ;
        RECT 27.230 87.770 27.500 87.970 ;
        RECT 27.230 87.080 27.440 87.770 ;
        RECT 28.100 87.630 28.370 88.180 ;
        RECT 28.510 88.090 28.670 89.000 ;
        RECT 28.510 87.970 28.680 88.090 ;
        RECT 28.910 87.970 29.070 89.120 ;
        RECT 29.890 88.870 30.210 89.190 ;
        RECT 30.530 88.590 30.740 89.320 ;
        RECT 30.510 88.270 30.770 88.590 ;
        RECT 27.220 87.020 27.480 87.080 ;
        RECT 27.220 86.770 27.860 87.020 ;
        RECT 27.220 86.760 27.480 86.770 ;
        RECT 26.750 85.670 27.090 86.010 ;
        RECT 26.790 85.650 27.010 85.670 ;
        RECT 11.670 71.260 11.910 83.640 ;
        RECT 14.610 82.810 14.920 83.640 ;
        RECT 19.040 83.320 19.330 83.640 ;
        RECT 19.540 83.340 19.880 83.660 ;
        RECT 19.010 82.970 19.360 83.320 ;
        RECT 14.570 82.480 14.940 82.810 ;
        RECT 19.040 82.510 19.330 82.970 ;
        RECT 19.540 82.730 19.790 83.340 ;
        RECT 20.500 82.750 20.690 83.690 ;
        RECT 24.780 83.280 25.030 83.690 ;
        RECT 26.180 83.380 26.460 83.700 ;
        RECT 26.790 83.370 26.990 85.650 ;
        RECT 27.140 84.720 27.460 85.040 ;
        RECT 27.250 84.080 27.440 84.190 ;
        RECT 27.190 83.760 27.510 84.080 ;
        RECT 24.750 82.990 25.090 83.280 ;
        RECT 26.750 83.050 27.030 83.370 ;
        RECT 27.210 83.360 27.490 83.760 ;
        RECT 14.610 81.270 14.920 82.480 ;
        RECT 18.470 82.230 19.330 82.510 ;
        RECT 18.390 82.220 19.330 82.230 ;
        RECT 19.490 82.620 19.790 82.730 ;
        RECT 18.390 81.750 18.850 82.220 ;
        RECT 14.560 80.790 14.980 81.270 ;
        RECT 19.490 81.110 19.680 82.620 ;
        RECT 20.440 82.430 20.760 82.750 ;
        RECT 23.120 82.410 23.380 82.480 ;
        RECT 23.860 82.410 24.120 82.480 ;
        RECT 19.850 81.760 20.170 82.080 ;
        RECT 20.940 81.760 21.260 82.080 ;
        RECT 22.040 81.750 22.360 82.070 ;
        RECT 19.050 80.790 19.680 81.110 ;
        RECT 20.400 81.080 20.720 81.400 ;
        RECT 23.120 81.380 24.120 82.410 ;
        RECT 27.680 82.140 27.860 86.770 ;
        RECT 28.100 86.220 28.260 87.630 ;
        RECT 28.510 87.050 28.700 87.970 ;
        RECT 28.860 87.920 29.070 87.970 ;
        RECT 28.860 87.680 29.090 87.920 ;
        RECT 29.890 87.900 30.210 88.220 ;
        RECT 28.870 87.660 29.070 87.680 ;
        RECT 28.480 87.020 28.720 87.050 ;
        RECT 28.910 87.020 29.070 87.660 ;
        RECT 29.890 87.350 30.210 87.670 ;
        RECT 28.480 86.850 29.070 87.020 ;
        RECT 28.480 86.820 28.720 86.850 ;
        RECT 28.100 85.670 28.370 86.220 ;
        RECT 28.090 85.620 28.370 85.670 ;
        RECT 28.510 85.880 28.700 86.820 ;
        RECT 28.910 86.190 29.070 86.850 ;
        RECT 28.870 86.170 29.070 86.190 ;
        RECT 29.890 86.180 30.210 86.500 ;
        RECT 30.510 86.390 30.770 86.710 ;
        RECT 28.860 85.930 29.090 86.170 ;
        RECT 28.860 85.880 29.070 85.930 ;
        RECT 28.510 85.760 28.680 85.880 ;
        RECT 28.090 85.530 28.260 85.620 ;
        RECT 28.100 85.070 28.260 85.530 ;
        RECT 28.090 84.980 28.260 85.070 ;
        RECT 28.090 84.930 28.370 84.980 ;
        RECT 28.100 84.380 28.370 84.930 ;
        RECT 28.510 84.840 28.670 85.760 ;
        RECT 28.510 84.720 28.680 84.840 ;
        RECT 28.910 84.720 29.070 85.880 ;
        RECT 29.890 85.630 30.210 85.950 ;
        RECT 30.510 85.530 30.670 86.390 ;
        RECT 30.380 85.210 30.670 85.530 ;
        RECT 30.970 85.460 31.220 89.890 ;
        RECT 33.030 87.980 33.410 93.000 ;
        RECT 34.780 90.170 35.020 93.000 ;
        RECT 34.780 89.850 35.250 90.170 ;
        RECT 33.030 86.120 33.420 87.980 ;
        RECT 30.950 85.430 31.230 85.460 ;
        RECT 30.940 85.150 31.240 85.430 ;
        RECT 30.950 85.130 31.230 85.150 ;
        RECT 28.100 83.680 28.260 84.380 ;
        RECT 28.510 83.730 28.700 84.720 ;
        RECT 28.860 84.670 29.070 84.720 ;
        RECT 28.860 84.430 29.090 84.670 ;
        RECT 29.890 84.650 30.210 84.970 ;
        RECT 28.870 84.410 29.070 84.430 ;
        RECT 28.910 83.680 29.070 84.410 ;
        RECT 29.890 84.100 30.210 84.420 ;
        RECT 29.000 83.300 29.260 83.330 ;
        RECT 28.980 83.000 29.280 83.300 ;
        RECT 29.000 82.990 29.260 83.000 ;
        RECT 24.880 81.750 25.200 82.070 ;
        RECT 25.980 81.760 26.300 82.080 ;
        RECT 27.070 81.760 27.390 82.080 ;
        RECT 27.680 81.840 28.160 82.140 ;
        RECT 29.010 82.070 29.230 82.990 ;
        RECT 30.970 82.860 31.220 85.130 ;
        RECT 33.030 83.670 33.410 86.120 ;
        RECT 34.980 85.430 35.250 89.850 ;
        RECT 34.960 85.120 35.270 85.430 ;
        RECT 34.980 82.880 35.250 85.120 ;
        RECT 37.060 83.670 37.460 93.000 ;
        RECT 40.580 91.350 40.820 93.000 ;
        RECT 59.390 92.690 59.760 114.480 ;
        RECT 59.350 92.180 59.840 92.690 ;
        RECT 59.390 92.150 59.760 92.180 ;
        RECT 40.580 91.110 41.160 91.350 ;
        RECT 38.580 89.120 38.900 89.440 ;
        RECT 38.730 88.440 39.050 88.760 ;
        RECT 38.730 87.550 39.050 87.870 ;
        RECT 38.580 86.870 38.900 87.190 ;
        RECT 38.580 86.350 38.900 86.670 ;
        RECT 38.730 85.670 39.050 85.990 ;
        RECT 38.730 84.780 39.050 85.100 ;
        RECT 38.580 84.100 38.900 84.420 ;
        RECT 39.660 83.850 39.890 89.900 ;
        RECT 40.920 89.770 41.160 91.110 ;
        RECT 40.920 85.550 41.150 89.770 ;
        RECT 46.040 88.710 46.300 88.770 ;
        RECT 46.030 88.450 46.300 88.710 ;
        RECT 45.520 87.520 45.780 87.840 ;
        RECT 45.050 85.680 45.310 86.000 ;
        RECT 40.880 85.540 41.160 85.550 ;
        RECT 40.880 85.220 41.180 85.540 ;
        RECT 37.800 83.310 38.230 83.710 ;
        RECT 30.960 82.600 31.280 82.860 ;
        RECT 34.980 82.570 35.330 82.880 ;
        RECT 32.930 82.330 33.190 82.510 ;
        RECT 33.670 82.330 33.930 82.510 ;
        RECT 27.760 81.730 28.160 81.840 ;
        RECT 28.950 81.670 29.290 82.070 ;
        RECT 29.660 81.790 29.980 82.110 ;
        RECT 30.750 81.790 31.070 82.110 ;
        RECT 31.850 81.780 32.170 82.100 ;
        RECT 29.010 81.590 29.230 81.670 ;
        RECT 21.490 81.060 21.810 81.380 ;
        RECT 22.880 81.370 23.380 81.380 ;
        RECT 22.600 81.060 23.380 81.370 ;
        RECT 22.600 81.050 22.920 81.060 ;
        RECT 19.050 80.690 19.490 80.790 ;
        RECT 23.120 80.040 23.380 81.060 ;
        RECT 22.880 80.030 23.380 80.040 ;
        RECT 20.400 79.710 20.720 80.030 ;
        RECT 21.490 79.710 21.810 80.030 ;
        RECT 22.590 79.720 23.380 80.030 ;
        RECT 22.590 79.710 22.910 79.720 ;
        RECT 19.840 78.980 20.160 79.300 ;
        RECT 20.940 78.980 21.260 79.300 ;
        RECT 22.040 78.980 22.360 79.300 ;
        RECT 19.840 77.610 20.160 77.930 ;
        RECT 20.940 77.610 21.260 77.930 ;
        RECT 22.040 77.610 22.360 77.930 ;
        RECT 19.270 77.260 19.590 77.290 ;
        RECT 23.120 77.270 23.380 79.720 ;
        RECT 22.880 77.260 23.380 77.270 ;
        RECT 19.260 76.970 19.590 77.260 ;
        RECT 19.260 76.820 19.580 76.970 ;
        RECT 20.400 76.930 20.720 77.250 ;
        RECT 21.490 76.930 21.810 77.250 ;
        RECT 22.590 76.950 23.380 77.260 ;
        RECT 22.590 76.940 22.910 76.950 ;
        RECT 19.260 76.500 19.600 76.820 ;
        RECT 19.260 75.510 19.580 76.500 ;
        RECT 23.120 76.290 23.380 76.950 ;
        RECT 23.860 81.370 24.360 81.380 ;
        RECT 23.860 81.060 24.640 81.370 ;
        RECT 25.430 81.060 25.750 81.380 ;
        RECT 26.520 81.080 26.840 81.400 ;
        RECT 30.210 81.110 30.530 81.430 ;
        RECT 31.300 81.090 31.620 81.410 ;
        RECT 32.930 81.400 33.930 82.330 ;
        RECT 34.690 81.780 35.010 82.100 ;
        RECT 35.790 81.790 36.110 82.110 ;
        RECT 36.880 81.790 37.200 82.110 ;
        RECT 37.840 81.520 38.190 83.310 ;
        RECT 39.660 82.750 39.880 83.850 ;
        RECT 40.920 83.350 41.150 85.220 ;
        RECT 44.550 84.750 44.810 85.070 ;
        RECT 40.920 83.120 44.130 83.350 ;
        RECT 40.920 83.110 41.150 83.120 ;
        RECT 39.370 82.510 39.880 82.750 ;
        RECT 32.410 81.080 33.190 81.400 ;
        RECT 23.860 80.030 24.120 81.060 ;
        RECT 24.320 81.050 24.640 81.060 ;
        RECT 32.930 80.060 33.190 81.080 ;
        RECT 23.860 79.710 24.650 80.030 ;
        RECT 25.430 79.710 25.750 80.030 ;
        RECT 26.520 79.710 26.840 80.030 ;
        RECT 30.210 79.740 30.530 80.060 ;
        RECT 31.300 79.740 31.620 80.060 ;
        RECT 32.400 79.740 33.190 80.060 ;
        RECT 23.860 77.260 24.120 79.710 ;
        RECT 24.880 78.980 25.200 79.300 ;
        RECT 25.980 78.980 26.300 79.300 ;
        RECT 27.080 78.980 27.400 79.300 ;
        RECT 29.650 79.010 29.970 79.330 ;
        RECT 30.750 79.010 31.070 79.330 ;
        RECT 31.850 79.010 32.170 79.330 ;
        RECT 24.880 77.610 25.200 77.930 ;
        RECT 25.980 77.610 26.300 77.930 ;
        RECT 27.080 77.610 27.400 77.930 ;
        RECT 29.650 77.640 29.970 77.960 ;
        RECT 30.750 77.640 31.070 77.960 ;
        RECT 31.850 77.640 32.170 77.960 ;
        RECT 27.650 77.280 27.970 77.290 ;
        RECT 23.860 76.940 24.650 77.260 ;
        RECT 23.860 76.310 24.120 76.940 ;
        RECT 25.430 76.930 25.750 77.250 ;
        RECT 26.520 76.930 26.840 77.250 ;
        RECT 23.110 75.950 23.390 76.290 ;
        RECT 23.850 75.970 24.130 76.310 ;
        RECT 19.140 74.910 19.680 75.510 ;
        RECT 23.120 74.540 23.380 75.950 ;
        RECT 23.860 74.540 24.120 75.970 ;
        RECT 11.270 69.940 11.920 71.260 ;
        RECT 23.120 71.110 24.120 74.540 ;
        RECT 27.630 74.490 27.970 77.280 ;
        RECT 29.080 77.270 29.400 77.320 ;
        RECT 32.930 77.290 33.190 79.740 ;
        RECT 29.060 76.850 29.400 77.270 ;
        RECT 30.210 76.960 30.530 77.280 ;
        RECT 31.300 76.960 31.620 77.280 ;
        RECT 32.400 76.970 33.190 77.290 ;
        RECT 29.060 76.530 29.410 76.850 ;
        RECT 27.570 73.970 28.030 74.490 ;
        RECT 29.060 73.600 29.400 76.530 ;
        RECT 32.930 76.290 33.190 76.970 ;
        RECT 33.670 81.080 34.450 81.400 ;
        RECT 35.240 81.090 35.560 81.410 ;
        RECT 36.330 81.110 36.650 81.430 ;
        RECT 39.370 81.260 39.600 82.510 ;
        RECT 43.900 82.150 44.130 83.120 ;
        RECT 40.430 81.770 40.750 82.090 ;
        RECT 41.530 81.780 41.850 82.100 ;
        RECT 42.620 81.780 42.940 82.100 ;
        RECT 43.850 81.750 44.160 82.150 ;
        RECT 33.670 80.050 33.930 81.080 ;
        RECT 39.260 80.820 39.720 81.260 ;
        RECT 39.870 81.070 40.190 81.390 ;
        RECT 40.980 81.080 41.300 81.400 ;
        RECT 42.070 81.100 42.390 81.420 ;
        RECT 34.140 80.050 34.460 80.060 ;
        RECT 33.670 79.740 34.460 80.050 ;
        RECT 35.240 79.740 35.560 80.060 ;
        RECT 36.330 79.740 36.650 80.060 ;
        RECT 33.670 79.730 34.170 79.740 ;
        RECT 39.880 79.730 40.200 80.050 ;
        RECT 40.980 79.730 41.300 80.050 ;
        RECT 42.070 79.730 42.390 80.050 ;
        RECT 33.670 77.290 33.930 79.730 ;
        RECT 34.690 79.010 35.010 79.330 ;
        RECT 35.790 79.010 36.110 79.330 ;
        RECT 36.890 79.010 37.210 79.330 ;
        RECT 40.430 79.000 40.750 79.320 ;
        RECT 41.530 79.000 41.850 79.320 ;
        RECT 42.630 79.000 42.950 79.320 ;
        RECT 43.360 78.970 43.630 79.000 ;
        RECT 43.350 78.440 43.630 78.970 ;
        RECT 43.900 78.580 44.130 81.750 ;
        RECT 43.770 78.440 44.130 78.580 ;
        RECT 43.350 78.140 44.130 78.440 ;
        RECT 43.340 78.130 44.130 78.140 ;
        RECT 43.340 78.120 44.110 78.130 ;
        RECT 34.690 77.640 35.010 77.960 ;
        RECT 35.790 77.640 36.110 77.960 ;
        RECT 36.890 77.640 37.210 77.960 ;
        RECT 40.430 77.630 40.750 77.950 ;
        RECT 41.530 77.630 41.850 77.950 ;
        RECT 42.630 77.630 42.950 77.950 ;
        RECT 43.340 77.690 43.630 78.120 ;
        RECT 33.670 76.970 34.460 77.290 ;
        RECT 32.920 75.950 33.200 76.290 ;
        RECT 32.930 74.770 33.190 75.950 ;
        RECT 33.670 74.770 33.930 76.970 ;
        RECT 35.240 76.960 35.560 77.280 ;
        RECT 36.330 76.960 36.650 77.280 ;
        RECT 37.460 77.000 37.780 77.320 ;
        RECT 37.480 76.850 37.750 77.000 ;
        RECT 39.880 76.960 40.200 77.280 ;
        RECT 40.980 76.950 41.300 77.270 ;
        RECT 42.070 76.950 42.390 77.270 ;
        RECT 43.200 76.990 43.520 77.310 ;
        RECT 44.550 76.910 44.800 84.750 ;
        RECT 45.050 77.810 45.300 85.680 ;
        RECT 45.530 78.720 45.780 87.520 ;
        RECT 46.030 79.610 46.280 88.450 ;
        RECT 61.870 81.110 62.370 116.940 ;
        RECT 62.800 86.390 63.300 117.430 ;
        RECT 63.930 91.620 64.430 117.890 ;
        RECT 65.060 96.790 65.560 118.510 ;
        RECT 73.920 116.910 75.200 129.110 ;
        RECT 73.910 115.570 75.200 116.910 ;
        RECT 73.920 115.080 75.200 115.570 ;
        RECT 78.280 113.900 78.480 113.930 ;
        RECT 78.190 113.400 78.500 113.900 ;
        RECT 74.370 112.130 74.720 112.610 ;
        RECT 70.380 108.930 70.850 109.420 ;
        RECT 65.010 96.230 65.560 96.790 ;
        RECT 63.920 91.060 64.440 91.620 ;
        RECT 62.790 85.870 63.310 86.390 ;
        RECT 61.710 80.540 62.370 81.110 ;
        RECT 45.980 79.030 46.350 79.610 ;
        RECT 45.450 78.140 45.820 78.720 ;
        RECT 44.960 77.230 45.330 77.810 ;
        RECT 37.450 76.530 37.770 76.850 ;
        RECT 43.190 76.690 43.510 76.840 ;
        RECT 28.970 73.080 29.490 73.600 ;
        RECT 32.930 71.170 33.930 74.770 ;
        RECT 37.480 72.720 37.750 76.530 ;
        RECT 43.190 76.520 43.550 76.690 ;
        RECT 37.370 72.160 37.860 72.720 ;
        RECT 32.930 71.130 34.950 71.170 ;
        RECT 22.640 71.070 24.570 71.110 ;
        RECT 22.100 69.880 24.570 71.070 ;
        RECT 9.620 65.650 9.990 66.030 ;
        RECT 8.970 65.030 9.360 65.420 ;
        RECT 8.370 64.400 8.750 64.790 ;
        RECT 7.780 63.770 8.130 64.140 ;
        RECT 7.140 63.090 7.500 63.470 ;
        RECT 6.550 62.850 6.890 62.860 ;
        RECT 6.530 62.480 6.910 62.850 ;
        RECT 6.550 62.470 6.880 62.480 ;
        RECT 4.770 60.630 5.120 60.960 ;
        RECT 4.790 60.570 5.120 60.630 ;
        RECT 3.500 59.350 3.850 59.680 ;
        RECT 3.500 59.280 3.830 59.350 ;
        RECT 1.360 58.620 2.600 58.950 ;
        RECT 2.890 58.650 3.330 59.070 ;
        RECT 1.360 58.510 1.940 58.620 ;
        RECT 22.100 58.390 23.040 69.880 ;
        RECT 32.450 69.850 34.950 71.130 ;
        RECT 34.060 59.850 34.950 69.850 ;
        RECT 43.220 66.700 43.550 76.520 ;
        RECT 44.490 76.340 44.840 76.910 ;
        RECT 61.870 72.230 62.370 80.540 ;
        RECT 62.800 73.140 63.300 85.870 ;
        RECT 63.930 74.010 64.430 91.060 ;
        RECT 65.060 75.520 65.560 96.230 ;
        RECT 67.950 83.080 68.530 83.640 ;
        RECT 67.980 83.070 68.490 83.080 ;
        RECT 65.060 74.960 65.620 75.520 ;
        RECT 65.060 74.830 65.560 74.960 ;
        RECT 67.980 71.200 68.480 83.070 ;
        RECT 67.350 69.920 68.480 71.200 ;
        RECT 43.160 66.310 43.590 66.700 ;
        RECT 70.430 65.580 70.830 108.930 ;
        RECT 71.350 108.320 71.770 108.680 ;
        RECT 70.420 65.120 70.890 65.580 ;
        RECT 71.360 64.780 71.750 108.320 ;
        RECT 72.270 105.930 72.720 106.360 ;
        RECT 71.330 64.310 71.790 64.780 ;
        RECT 72.290 63.960 72.680 105.930 ;
        RECT 73.130 105.670 73.510 105.680 ;
        RECT 73.110 105.370 73.530 105.670 ;
        RECT 72.270 63.500 72.740 63.960 ;
        RECT 73.130 63.160 73.510 105.370 ;
        RECT 74.470 82.140 74.700 112.130 ;
        RECT 78.280 109.560 78.480 113.400 ;
        RECT 79.180 110.000 79.500 110.320 ;
        RECT 80.180 109.880 80.410 110.170 ;
        RECT 80.750 110.000 81.070 110.320 ;
        RECT 81.310 109.890 81.540 110.180 ;
        RECT 77.770 109.340 78.000 109.530 ;
        RECT 77.770 109.240 78.120 109.340 ;
        RECT 78.270 109.270 78.500 109.560 ;
        RECT 80.200 109.410 80.390 109.880 ;
        RECT 77.780 109.020 78.120 109.240 ;
        RECT 77.780 108.510 78.120 108.730 ;
        RECT 77.770 108.410 78.120 108.510 ;
        RECT 78.280 108.480 78.480 109.270 ;
        RECT 80.130 109.090 80.390 109.410 ;
        RECT 81.310 109.400 81.500 109.890 ;
        RECT 81.790 109.560 81.980 130.240 ;
        RECT 100.470 128.000 104.820 131.700 ;
        RECT 130.020 127.520 133.250 132.100 ;
        RECT 129.720 123.470 133.270 127.520 ;
        RECT 158.610 121.890 161.840 132.100 ;
        RECT 85.130 121.580 85.950 121.670 ;
        RECT 85.070 120.890 85.950 121.580 ;
        RECT 81.130 109.150 81.500 109.400 ;
        RECT 81.770 109.270 82.000 109.560 ;
        RECT 81.130 109.080 81.400 109.150 ;
        RECT 77.770 108.220 78.000 108.410 ;
        RECT 78.270 108.190 78.500 108.480 ;
        RECT 80.130 108.340 80.390 108.660 ;
        RECT 81.130 108.600 81.400 108.670 ;
        RECT 81.130 108.350 81.500 108.600 ;
        RECT 81.790 108.480 81.980 109.270 ;
        RECT 78.280 106.360 78.480 108.190 ;
        RECT 80.200 107.870 80.390 108.340 ;
        RECT 79.180 107.430 79.500 107.750 ;
        RECT 80.180 107.580 80.410 107.870 ;
        RECT 81.310 107.860 81.500 108.350 ;
        RECT 81.770 108.190 82.000 108.480 ;
        RECT 80.750 107.430 81.070 107.750 ;
        RECT 81.310 107.570 81.540 107.860 ;
        RECT 79.180 106.800 79.500 107.120 ;
        RECT 80.180 106.680 80.410 106.970 ;
        RECT 80.750 106.800 81.070 107.120 ;
        RECT 81.310 106.690 81.540 106.980 ;
        RECT 77.770 106.140 78.000 106.330 ;
        RECT 77.770 106.040 78.120 106.140 ;
        RECT 78.270 106.070 78.500 106.360 ;
        RECT 80.200 106.210 80.390 106.680 ;
        RECT 77.780 105.820 78.120 106.040 ;
        RECT 77.780 105.310 78.120 105.530 ;
        RECT 77.770 105.210 78.120 105.310 ;
        RECT 78.280 105.280 78.480 106.070 ;
        RECT 80.130 105.890 80.390 106.210 ;
        RECT 81.310 106.200 81.500 106.690 ;
        RECT 81.790 106.360 81.980 108.190 ;
        RECT 81.130 105.950 81.500 106.200 ;
        RECT 81.770 106.070 82.000 106.360 ;
        RECT 81.130 105.880 81.400 105.950 ;
        RECT 77.770 105.020 78.000 105.210 ;
        RECT 78.270 104.990 78.500 105.280 ;
        RECT 80.130 105.140 80.390 105.460 ;
        RECT 81.130 105.400 81.400 105.470 ;
        RECT 81.130 105.150 81.500 105.400 ;
        RECT 81.790 105.280 81.980 106.070 ;
        RECT 78.280 104.070 78.480 104.990 ;
        RECT 80.200 104.670 80.390 105.140 ;
        RECT 79.180 104.230 79.500 104.550 ;
        RECT 80.180 104.380 80.410 104.670 ;
        RECT 81.310 104.660 81.500 105.150 ;
        RECT 81.770 104.990 82.000 105.280 ;
        RECT 80.750 104.230 81.070 104.550 ;
        RECT 81.310 104.370 81.540 104.660 ;
        RECT 81.790 104.070 81.980 104.990 ;
        RECT 85.070 101.890 85.780 120.890 ;
        RECT 158.410 119.360 162.000 121.890 ;
        RECT 187.200 118.400 190.430 132.100 ;
        RECT 212.630 129.160 213.620 129.170 ;
        RECT 212.630 128.640 214.020 129.160 ;
        RECT 207.400 128.110 210.820 128.160 ;
        RECT 207.390 127.540 210.830 128.110 ;
        RECT 205.540 126.720 206.260 127.270 ;
        RECT 205.760 126.710 206.260 126.720 ;
        RECT 186.890 114.780 190.650 118.400 ;
        RECT 201.240 117.750 204.650 118.030 ;
        RECT 201.240 117.730 205.360 117.750 ;
        RECT 201.240 117.710 206.110 117.730 ;
        RECT 207.940 117.710 212.240 126.770 ;
        RECT 213.530 125.030 214.020 128.640 ;
        RECT 201.240 115.960 214.640 117.710 ;
        RECT 201.240 115.950 215.590 115.960 ;
        RECT 201.240 115.600 215.750 115.950 ;
        RECT 201.240 115.590 215.590 115.600 ;
        RECT 201.240 115.240 214.640 115.590 ;
        RECT 84.940 101.100 85.780 101.890 ;
        RECT 109.560 84.320 113.980 114.430 ;
        RECT 201.240 113.990 214.270 115.240 ;
        RECT 204.650 113.800 214.270 113.990 ;
        RECT 204.650 113.790 206.110 113.800 ;
        RECT 205.340 113.780 206.110 113.790 ;
        RECT 207.660 104.090 212.810 113.800 ;
        RECT 207.660 103.420 212.800 104.090 ;
        RECT 213.470 104.000 214.100 104.060 ;
        RECT 213.450 103.420 214.100 104.000 ;
        RECT 213.470 102.670 214.100 103.420 ;
        RECT 205.840 101.950 214.100 102.670 ;
        RECT 211.510 101.720 214.100 101.950 ;
        RECT 213.470 101.690 214.100 101.720 ;
        RECT 212.630 100.570 213.620 100.580 ;
        RECT 212.630 100.050 214.020 100.570 ;
        RECT 207.400 99.520 210.820 99.570 ;
        RECT 207.390 98.950 210.830 99.520 ;
        RECT 205.540 98.130 206.260 98.680 ;
        RECT 205.760 98.120 206.260 98.130 ;
        RECT 192.830 89.120 195.150 89.200 ;
        RECT 204.640 89.140 205.340 89.150 ;
        RECT 204.640 89.120 206.110 89.140 ;
        RECT 207.940 89.120 212.240 98.180 ;
        RECT 213.530 96.440 214.020 100.050 ;
        RECT 192.830 87.370 214.640 89.120 ;
        RECT 192.830 87.360 215.590 87.370 ;
        RECT 192.830 87.010 215.750 87.360 ;
        RECT 192.830 87.000 215.590 87.010 ;
        RECT 192.830 86.650 214.640 87.000 ;
        RECT 192.830 85.890 214.270 86.650 ;
        RECT 192.830 85.830 195.150 85.890 ;
        RECT 204.640 85.210 214.270 85.890 ;
        RECT 204.640 85.190 206.110 85.210 ;
        RECT 80.660 83.060 81.380 83.630 ;
        RECT 74.470 81.910 74.710 82.140 ;
        RECT 74.470 74.260 74.700 81.910 ;
        RECT 80.720 76.050 81.230 83.060 ;
        RECT 109.530 83.000 114.000 84.320 ;
        RECT 80.580 76.000 81.230 76.050 ;
        RECT 80.570 75.820 81.230 76.000 ;
        RECT 80.540 75.810 81.230 75.820 ;
        RECT 80.540 75.440 81.140 75.810 ;
        RECT 74.460 74.030 74.750 74.260 ;
        RECT 74.470 72.650 74.700 74.030 ;
        RECT 80.540 73.570 81.120 75.440 ;
        RECT 79.970 73.250 81.120 73.570 ;
        RECT 80.190 72.900 81.120 73.250 ;
        RECT 74.460 72.420 74.750 72.650 ;
        RECT 79.970 72.580 81.120 72.900 ;
        RECT 74.470 71.050 74.700 72.420 ;
        RECT 80.540 71.800 81.120 72.580 ;
        RECT 80.130 71.610 80.450 71.660 ;
        RECT 79.900 71.380 80.450 71.610 ;
        RECT 80.130 71.340 80.450 71.380 ;
        RECT 80.590 71.200 81.120 71.800 ;
        RECT 80.550 71.190 81.120 71.200 ;
        RECT 74.460 70.820 74.750 71.050 ;
        RECT 74.470 69.430 74.700 70.820 ;
        RECT 80.540 70.190 81.120 71.190 ;
        RECT 80.130 70.000 80.450 70.050 ;
        RECT 76.180 69.910 78.190 69.940 ;
        RECT 75.690 69.740 78.190 69.910 ;
        RECT 79.900 69.770 80.450 70.000 ;
        RECT 75.690 69.690 76.200 69.740 ;
        RECT 75.690 69.680 75.980 69.690 ;
        RECT 74.460 69.200 74.750 69.430 ;
        RECT 74.470 67.830 74.700 69.200 ;
        RECT 75.190 68.220 75.510 68.300 ;
        RECT 76.770 68.220 77.280 68.270 ;
        RECT 75.190 68.040 77.280 68.220 ;
        RECT 74.460 67.600 74.750 67.830 ;
        RECT 74.470 66.210 74.700 67.600 ;
        RECT 78.020 66.690 78.190 69.740 ;
        RECT 80.130 69.730 80.450 69.770 ;
        RECT 80.590 69.590 81.120 70.190 ;
        RECT 80.540 68.580 81.120 69.590 ;
        RECT 80.120 68.390 80.440 68.440 ;
        RECT 79.890 68.160 80.440 68.390 ;
        RECT 80.120 68.120 80.440 68.160 ;
        RECT 80.580 67.980 81.120 68.580 ;
        RECT 80.540 66.960 81.120 67.980 ;
        RECT 80.130 66.770 80.450 66.820 ;
        RECT 77.600 66.490 78.190 66.690 ;
        RECT 79.900 66.540 80.450 66.770 ;
        RECT 80.130 66.500 80.450 66.540 ;
        RECT 77.600 66.470 78.110 66.490 ;
        RECT 77.600 66.460 77.890 66.470 ;
        RECT 80.590 66.360 81.120 66.960 ;
        RECT 74.460 65.980 74.750 66.210 ;
        RECT 74.470 64.610 74.700 65.980 ;
        RECT 80.540 65.350 81.120 66.360 ;
        RECT 80.120 65.160 80.440 65.210 ;
        RECT 79.890 64.930 80.440 65.160 ;
        RECT 80.120 64.890 80.440 64.930 ;
        RECT 80.580 64.750 81.120 65.350 ;
        RECT 74.460 64.380 74.750 64.610 ;
        RECT 73.100 62.700 73.540 63.160 ;
        RECT 74.470 62.990 74.700 64.380 ;
        RECT 79.710 63.240 80.030 63.560 ;
        RECT 79.760 63.010 79.990 63.240 ;
        RECT 74.460 62.760 74.750 62.990 ;
        RECT 80.540 62.880 81.120 64.750 ;
        RECT 80.120 61.960 80.440 62.010 ;
        RECT 79.890 61.730 80.440 61.960 ;
        RECT 80.120 61.690 80.440 61.730 ;
        RECT 80.580 60.670 81.120 62.880 ;
        RECT 76.880 60.250 77.200 60.300 ;
        RECT 77.820 60.250 78.140 60.300 ;
        RECT 76.650 60.020 77.200 60.250 ;
        RECT 77.590 60.020 78.140 60.250 ;
        RECT 78.770 60.230 79.090 60.280 ;
        RECT 80.080 60.250 80.400 60.300 ;
        RECT 76.880 59.980 77.200 60.020 ;
        RECT 77.820 59.980 78.140 60.020 ;
        RECT 78.540 60.000 79.090 60.230 ;
        RECT 79.850 60.020 80.400 60.250 ;
        RECT 78.770 59.960 79.090 60.000 ;
        RECT 80.080 59.980 80.400 60.020 ;
        RECT 34.060 59.120 34.980 59.850 ;
        RECT 34.030 58.390 34.950 59.120 ;
        RECT -150.680 57.340 -141.110 58.020 ;
        RECT -127.070 57.870 -124.840 58.020 ;
        RECT -149.220 47.630 -144.070 57.340 ;
        RECT -142.520 57.320 -141.110 57.340 ;
        RECT -141.750 57.310 -141.110 57.320 ;
        RECT -150.510 47.540 -149.880 47.600 ;
        RECT -150.510 46.960 -149.860 47.540 ;
        RECT -149.210 46.960 -144.070 47.630 ;
        RECT -150.510 46.210 -149.880 46.960 ;
        RECT -150.510 45.490 -142.250 46.210 ;
        RECT -150.510 45.260 -147.920 45.490 ;
        RECT -150.510 45.230 -149.880 45.260 ;
        RECT -150.030 44.110 -149.040 44.120 ;
        RECT -150.430 43.590 -149.040 44.110 ;
        RECT -150.430 39.980 -149.940 43.590 ;
        RECT -147.230 43.060 -143.810 43.110 ;
        RECT -147.240 42.490 -143.800 43.060 ;
        RECT -148.650 32.660 -144.350 41.720 ;
        RECT -142.670 41.670 -141.950 42.220 ;
        RECT -142.670 41.660 -142.170 41.670 ;
        RECT -142.520 32.670 -141.750 32.680 ;
        RECT -142.520 32.660 -141.120 32.670 ;
        RECT -122.560 32.660 -120.150 32.760 ;
        RECT -151.050 30.910 -120.150 32.660 ;
        RECT -152.000 30.900 -120.150 30.910 ;
        RECT -152.160 30.550 -120.150 30.900 ;
        RECT -152.000 30.540 -120.150 30.550 ;
        RECT -151.050 30.190 -120.150 30.540 ;
        RECT -150.680 29.430 -120.150 30.190 ;
        RECT -150.680 28.750 -141.120 29.430 ;
        RECT -122.560 29.330 -120.150 29.430 ;
        RECT -149.220 19.040 -144.070 28.750 ;
        RECT -142.520 28.730 -141.120 28.750 ;
        RECT -150.510 18.950 -149.880 19.010 ;
        RECT -150.510 18.370 -149.860 18.950 ;
        RECT -149.210 18.370 -144.070 19.040 ;
        RECT -150.510 17.620 -149.880 18.370 ;
        RECT -150.510 16.900 -142.250 17.620 ;
        RECT -150.510 16.670 -147.920 16.900 ;
        RECT -150.510 16.640 -149.880 16.670 ;
        RECT -150.030 15.520 -149.040 15.530 ;
        RECT -150.430 15.000 -149.040 15.520 ;
        RECT -150.430 11.390 -149.940 15.000 ;
        RECT -147.230 14.470 -143.810 14.520 ;
        RECT -147.240 13.900 -143.800 14.470 ;
        RECT -148.650 4.070 -144.350 13.130 ;
        RECT -142.670 13.080 -141.950 13.630 ;
        RECT -142.670 13.070 -142.170 13.080 ;
        RECT -142.520 4.070 -141.110 4.090 ;
        RECT -118.000 4.070 -115.730 4.140 ;
        RECT -151.050 2.320 -115.730 4.070 ;
        RECT -152.000 2.310 -115.730 2.320 ;
        RECT -152.160 1.960 -115.730 2.310 ;
        RECT -152.000 1.950 -115.730 1.960 ;
        RECT -151.050 1.600 -115.730 1.950 ;
        RECT -150.680 0.840 -115.730 1.600 ;
        RECT -150.680 0.160 -141.110 0.840 ;
        RECT -118.000 0.740 -115.730 0.840 ;
        RECT -149.220 -9.550 -144.070 0.160 ;
        RECT -142.520 0.150 -141.110 0.160 ;
        RECT -142.520 0.140 -141.750 0.150 ;
        RECT -150.510 -9.640 -149.880 -9.580 ;
        RECT -150.510 -10.220 -149.860 -9.640 ;
        RECT -149.210 -10.220 -144.070 -9.550 ;
        RECT -150.510 -10.970 -149.880 -10.220 ;
        RECT -150.510 -11.690 -142.250 -10.970 ;
        RECT -150.510 -11.920 -147.920 -11.690 ;
        RECT -150.510 -11.950 -149.880 -11.920 ;
        RECT -150.030 -13.070 -149.040 -13.060 ;
        RECT -150.430 -13.590 -149.040 -13.070 ;
        RECT -150.430 -17.200 -149.940 -13.590 ;
        RECT -147.230 -14.120 -143.810 -14.070 ;
        RECT -147.240 -14.690 -143.800 -14.120 ;
        RECT -148.650 -24.520 -144.350 -15.460 ;
        RECT -142.670 -15.510 -141.950 -14.960 ;
        RECT -142.670 -15.520 -142.170 -15.510 ;
        RECT -142.520 -24.520 -141.120 -24.500 ;
        RECT -113.640 -24.520 -111.390 -24.460 ;
        RECT -151.050 -26.270 -111.390 -24.520 ;
        RECT -152.000 -26.280 -111.390 -26.270 ;
        RECT -152.160 -26.630 -111.390 -26.280 ;
        RECT -152.000 -26.640 -111.390 -26.630 ;
        RECT -151.050 -26.990 -111.390 -26.640 ;
        RECT -150.680 -27.750 -111.390 -26.990 ;
        RECT -150.680 -28.430 -141.120 -27.750 ;
        RECT -113.640 -27.830 -111.390 -27.750 ;
        RECT -149.220 -38.140 -144.070 -28.430 ;
        RECT -142.520 -28.440 -141.120 -28.430 ;
        RECT -142.520 -28.450 -141.750 -28.440 ;
        RECT -150.510 -38.230 -149.880 -38.170 ;
        RECT -150.510 -38.810 -149.860 -38.230 ;
        RECT -149.210 -38.810 -144.070 -38.140 ;
        RECT -150.510 -39.560 -149.880 -38.810 ;
        RECT -150.510 -40.280 -142.250 -39.560 ;
        RECT -150.510 -40.510 -147.920 -40.280 ;
        RECT -150.510 -40.540 -149.880 -40.510 ;
        RECT -150.030 -41.660 -149.040 -41.650 ;
        RECT -150.430 -42.180 -149.040 -41.660 ;
        RECT -150.430 -45.790 -149.940 -42.180 ;
        RECT -147.230 -42.710 -143.810 -42.660 ;
        RECT -147.240 -43.280 -143.800 -42.710 ;
        RECT -148.650 -53.110 -144.350 -44.050 ;
        RECT -142.670 -44.100 -141.950 -43.550 ;
        RECT -142.670 -44.110 -142.170 -44.100 ;
        RECT -142.520 -53.110 -141.120 -53.090 ;
        RECT -109.320 -53.110 -107.070 -53.000 ;
        RECT -151.050 -54.860 -106.920 -53.110 ;
        RECT -152.000 -54.870 -106.920 -54.860 ;
        RECT -152.160 -55.220 -106.920 -54.870 ;
        RECT -152.000 -55.230 -106.920 -55.220 ;
        RECT -151.050 -55.580 -106.920 -55.230 ;
        RECT -150.680 -56.340 -106.920 -55.580 ;
        RECT -150.680 -57.020 -141.120 -56.340 ;
        RECT -109.320 -56.450 -107.070 -56.340 ;
        RECT -149.220 -66.730 -144.070 -57.020 ;
        RECT -142.520 -57.030 -141.120 -57.020 ;
        RECT -142.520 -57.040 -141.750 -57.030 ;
        RECT -150.510 -66.820 -149.880 -66.760 ;
        RECT -150.510 -67.400 -149.860 -66.820 ;
        RECT -149.210 -67.400 -144.070 -66.730 ;
        RECT -150.510 -68.150 -149.880 -67.400 ;
        RECT -150.510 -68.870 -142.250 -68.150 ;
        RECT -150.510 -69.100 -147.920 -68.870 ;
        RECT -150.510 -69.130 -149.880 -69.100 ;
        RECT -150.030 -70.250 -149.040 -70.240 ;
        RECT -150.430 -70.770 -149.040 -70.250 ;
        RECT -150.430 -74.380 -149.940 -70.770 ;
        RECT -147.230 -71.300 -143.810 -71.250 ;
        RECT -147.240 -71.870 -143.800 -71.300 ;
        RECT -148.650 -81.700 -144.350 -72.640 ;
        RECT -142.670 -72.690 -141.950 -72.140 ;
        RECT -142.670 -72.700 -142.170 -72.690 ;
        RECT 109.560 -78.300 113.980 83.000 ;
        RECT 207.660 75.500 212.810 85.210 ;
        RECT 207.660 74.830 212.800 75.500 ;
        RECT 213.470 75.410 214.100 75.470 ;
        RECT 213.450 74.830 214.100 75.410 ;
        RECT 213.470 74.080 214.100 74.830 ;
        RECT 205.840 73.360 214.100 74.080 ;
        RECT 211.510 73.130 214.100 73.360 ;
        RECT 213.470 73.100 214.100 73.130 ;
        RECT 212.630 71.980 213.620 71.990 ;
        RECT 212.630 71.460 214.020 71.980 ;
        RECT 207.400 70.930 210.820 70.980 ;
        RECT 207.390 70.360 210.830 70.930 ;
        RECT 205.540 69.540 206.260 70.090 ;
        RECT 205.760 69.530 206.260 69.540 ;
        RECT 188.660 60.530 191.020 60.660 ;
        RECT 204.660 60.550 205.360 60.560 ;
        RECT 204.660 60.530 206.110 60.550 ;
        RECT 207.940 60.530 212.240 69.590 ;
        RECT 213.530 67.850 214.020 71.460 ;
        RECT 188.660 58.780 214.640 60.530 ;
        RECT 188.660 58.770 215.590 58.780 ;
        RECT 188.660 58.420 215.750 58.770 ;
        RECT 188.660 58.410 215.590 58.420 ;
        RECT 188.660 58.060 214.640 58.410 ;
        RECT 188.660 57.300 214.270 58.060 ;
        RECT 188.660 57.200 191.020 57.300 ;
        RECT 204.660 56.620 214.270 57.300 ;
        RECT 204.660 56.600 206.110 56.620 ;
        RECT 207.660 46.910 212.810 56.620 ;
        RECT 207.660 46.240 212.800 46.910 ;
        RECT 213.470 46.820 214.100 46.880 ;
        RECT 213.450 46.240 214.100 46.820 ;
        RECT 213.470 45.490 214.100 46.240 ;
        RECT 205.840 44.770 214.100 45.490 ;
        RECT 211.510 44.540 214.100 44.770 ;
        RECT 213.470 44.510 214.100 44.540 ;
        RECT 212.630 43.390 213.620 43.400 ;
        RECT 212.630 42.870 214.020 43.390 ;
        RECT 207.400 42.340 210.820 42.390 ;
        RECT 207.390 41.770 210.830 42.340 ;
        RECT 205.540 40.950 206.260 41.500 ;
        RECT 205.760 40.940 206.260 40.950 ;
        RECT 184.650 31.940 186.930 32.100 ;
        RECT 204.640 31.960 205.340 31.970 ;
        RECT 204.640 31.940 206.110 31.960 ;
        RECT 207.940 31.940 212.240 41.000 ;
        RECT 213.530 39.260 214.020 42.870 ;
        RECT 184.650 30.190 214.640 31.940 ;
        RECT 184.650 30.180 215.590 30.190 ;
        RECT 184.650 29.830 215.750 30.180 ;
        RECT 184.650 29.820 215.590 29.830 ;
        RECT 184.650 29.470 214.640 29.820 ;
        RECT 184.650 28.710 214.270 29.470 ;
        RECT 184.650 28.600 186.930 28.710 ;
        RECT 204.640 28.030 214.270 28.710 ;
        RECT 204.640 28.010 206.110 28.030 ;
        RECT 207.660 18.320 212.810 28.030 ;
        RECT 207.660 17.650 212.800 18.320 ;
        RECT 213.470 18.230 214.100 18.290 ;
        RECT 213.450 17.650 214.100 18.230 ;
        RECT 213.470 16.900 214.100 17.650 ;
        RECT 205.840 16.180 214.100 16.900 ;
        RECT 211.510 15.950 214.100 16.180 ;
        RECT 213.470 15.920 214.100 15.950 ;
        RECT 212.630 14.800 213.620 14.810 ;
        RECT 212.630 14.280 214.020 14.800 ;
        RECT 207.400 13.750 210.820 13.800 ;
        RECT 207.390 13.180 210.830 13.750 ;
        RECT 205.540 12.360 206.260 12.910 ;
        RECT 205.760 12.350 206.260 12.360 ;
        RECT 180.350 3.350 182.770 3.470 ;
        RECT 204.640 3.350 206.110 3.370 ;
        RECT 207.940 3.350 212.240 12.410 ;
        RECT 213.530 10.670 214.020 14.280 ;
        RECT 180.350 1.600 214.640 3.350 ;
        RECT 180.350 1.590 215.590 1.600 ;
        RECT 180.350 1.240 215.750 1.590 ;
        RECT 180.350 1.230 215.590 1.240 ;
        RECT 180.350 0.880 214.640 1.230 ;
        RECT 180.350 0.120 214.270 0.880 ;
        RECT 180.350 -0.040 182.770 0.120 ;
        RECT 204.640 -0.560 214.270 0.120 ;
        RECT 204.640 -0.580 206.110 -0.560 ;
        RECT 204.640 -0.590 205.340 -0.580 ;
        RECT 207.660 -10.270 212.810 -0.560 ;
        RECT 207.660 -10.940 212.800 -10.270 ;
        RECT 213.470 -10.360 214.100 -10.300 ;
        RECT 213.450 -10.940 214.100 -10.360 ;
        RECT 213.470 -11.690 214.100 -10.940 ;
        RECT 205.840 -12.410 214.100 -11.690 ;
        RECT 211.510 -12.640 214.100 -12.410 ;
        RECT 213.470 -12.670 214.100 -12.640 ;
        RECT 212.630 -13.790 213.620 -13.780 ;
        RECT 212.630 -14.310 214.020 -13.790 ;
        RECT 207.400 -14.840 210.820 -14.790 ;
        RECT 207.390 -15.410 210.830 -14.840 ;
        RECT 205.540 -16.230 206.260 -15.680 ;
        RECT 205.760 -16.240 206.260 -16.230 ;
        RECT 176.460 -25.240 178.730 -25.130 ;
        RECT 204.650 -25.220 205.350 -25.210 ;
        RECT 204.650 -25.240 206.110 -25.220 ;
        RECT 207.940 -25.240 212.240 -16.180 ;
        RECT 213.530 -17.920 214.020 -14.310 ;
        RECT 176.460 -26.990 214.640 -25.240 ;
        RECT 176.460 -27.000 215.590 -26.990 ;
        RECT 176.460 -27.350 215.750 -27.000 ;
        RECT 176.460 -27.360 215.590 -27.350 ;
        RECT 176.460 -27.710 214.640 -27.360 ;
        RECT 176.460 -28.470 214.270 -27.710 ;
        RECT 176.460 -28.600 178.730 -28.470 ;
        RECT 204.650 -29.150 214.270 -28.470 ;
        RECT 204.650 -29.170 206.110 -29.150 ;
        RECT 207.660 -38.860 212.810 -29.150 ;
        RECT 207.660 -39.530 212.800 -38.860 ;
        RECT 213.470 -38.950 214.100 -38.890 ;
        RECT 213.450 -39.530 214.100 -38.950 ;
        RECT 213.470 -40.280 214.100 -39.530 ;
        RECT 205.840 -41.000 214.100 -40.280 ;
        RECT 211.510 -41.230 214.100 -41.000 ;
        RECT 213.470 -41.260 214.100 -41.230 ;
        RECT 212.630 -42.380 213.620 -42.370 ;
        RECT 212.630 -42.900 214.020 -42.380 ;
        RECT 207.400 -43.430 210.820 -43.380 ;
        RECT 207.390 -44.000 210.830 -43.430 ;
        RECT 205.540 -44.820 206.260 -44.270 ;
        RECT 205.760 -44.830 206.260 -44.820 ;
        RECT 172.060 -53.830 174.360 -53.750 ;
        RECT 204.650 -53.830 206.110 -53.810 ;
        RECT 207.940 -53.830 212.240 -44.770 ;
        RECT 213.530 -46.510 214.020 -42.900 ;
        RECT 172.060 -55.580 214.640 -53.830 ;
        RECT 172.060 -55.590 215.590 -55.580 ;
        RECT 172.060 -55.940 215.750 -55.590 ;
        RECT 172.060 -55.950 215.590 -55.940 ;
        RECT 172.060 -56.300 214.640 -55.950 ;
        RECT 172.060 -57.060 214.270 -56.300 ;
        RECT 172.060 -57.160 174.360 -57.060 ;
        RECT 204.650 -57.740 214.270 -57.060 ;
        RECT 204.650 -57.760 206.110 -57.740 ;
        RECT 204.650 -57.770 205.350 -57.760 ;
        RECT 207.660 -67.450 212.810 -57.740 ;
        RECT 207.660 -68.120 212.800 -67.450 ;
        RECT 213.470 -67.540 214.100 -67.480 ;
        RECT 213.450 -68.120 214.100 -67.540 ;
        RECT 213.470 -68.870 214.100 -68.120 ;
        RECT 205.840 -69.590 214.100 -68.870 ;
        RECT 211.510 -69.820 214.100 -69.590 ;
        RECT 213.470 -69.850 214.100 -69.820 ;
        RECT -142.520 -81.690 -141.750 -81.680 ;
        RECT -142.520 -81.700 -141.120 -81.690 ;
        RECT -105.260 -81.700 -102.850 -81.600 ;
        RECT -151.050 -83.450 -102.850 -81.700 ;
        RECT 108.640 -82.040 113.980 -78.300 ;
        RECT 108.640 -83.000 113.400 -82.040 ;
        RECT -152.000 -83.460 -102.850 -83.450 ;
        RECT -152.160 -83.810 -102.850 -83.460 ;
        RECT -152.000 -83.820 -102.850 -83.810 ;
        RECT -151.050 -84.170 -102.850 -83.820 ;
        RECT -150.680 -84.930 -102.850 -84.170 ;
        RECT -150.680 -85.610 -141.120 -84.930 ;
        RECT -105.260 -85.110 -102.850 -84.930 ;
        RECT -149.220 -95.320 -144.070 -85.610 ;
        RECT -142.520 -85.630 -141.120 -85.610 ;
        RECT -150.510 -95.410 -149.880 -95.350 ;
        RECT -150.510 -95.990 -149.860 -95.410 ;
        RECT -149.210 -95.990 -144.070 -95.320 ;
        RECT -150.510 -96.740 -149.880 -95.990 ;
        RECT -150.510 -97.460 -142.250 -96.740 ;
        RECT -150.510 -97.690 -147.920 -97.460 ;
        RECT -150.510 -97.720 -149.880 -97.690 ;
        RECT -150.030 -98.840 -149.040 -98.830 ;
        RECT -150.430 -99.360 -149.040 -98.840 ;
        RECT -150.430 -102.970 -149.940 -99.360 ;
        RECT -147.230 -99.890 -143.810 -99.840 ;
        RECT -147.240 -100.460 -143.800 -99.890 ;
        RECT -148.650 -110.290 -144.350 -101.230 ;
        RECT -142.670 -101.280 -141.950 -100.730 ;
        RECT -142.670 -101.290 -142.170 -101.280 ;
        RECT -142.520 -110.280 -141.750 -110.270 ;
        RECT -142.520 -110.290 -141.120 -110.280 ;
        RECT -100.980 -110.290 -98.520 -110.220 ;
        RECT -151.050 -112.040 -98.520 -110.290 ;
        RECT -152.000 -112.050 -98.520 -112.040 ;
        RECT -152.160 -112.400 -98.520 -112.050 ;
        RECT -152.000 -112.410 -98.520 -112.400 ;
        RECT -151.050 -112.760 -98.520 -112.410 ;
        RECT -150.680 -113.520 -98.520 -112.760 ;
        RECT -150.680 -114.200 -141.120 -113.520 ;
        RECT -100.980 -113.570 -98.520 -113.520 ;
        RECT -149.220 -123.910 -144.070 -114.200 ;
        RECT -142.520 -114.220 -141.120 -114.200 ;
        RECT -150.510 -124.000 -149.880 -123.940 ;
        RECT -150.510 -124.580 -149.860 -124.000 ;
        RECT -149.210 -124.580 -144.070 -123.910 ;
        RECT -150.510 -125.330 -149.880 -124.580 ;
        RECT -150.510 -126.050 -142.250 -125.330 ;
        RECT -150.510 -126.280 -147.920 -126.050 ;
        RECT -150.510 -126.310 -149.880 -126.280 ;
        RECT -150.030 -127.430 -149.040 -127.420 ;
        RECT -150.430 -127.950 -149.040 -127.430 ;
        RECT -150.430 -131.560 -149.940 -127.950 ;
        RECT -147.230 -128.480 -143.810 -128.430 ;
        RECT -147.240 -129.050 -143.800 -128.480 ;
        RECT -148.650 -138.880 -144.350 -129.820 ;
        RECT -142.670 -129.870 -141.950 -129.320 ;
        RECT -142.670 -129.880 -142.170 -129.870 ;
        RECT -141.770 -138.860 -141.130 -138.850 ;
        RECT -142.520 -138.880 -141.130 -138.860 ;
        RECT -96.610 -138.880 -94.210 -138.740 ;
        RECT -151.050 -140.630 -94.210 -138.880 ;
        RECT -152.000 -140.640 -94.210 -140.630 ;
        RECT -152.160 -140.990 -94.210 -140.640 ;
        RECT -152.000 -141.000 -94.210 -140.990 ;
        RECT -151.050 -141.350 -94.210 -141.000 ;
        RECT -150.680 -142.110 -94.210 -141.350 ;
        RECT -150.680 -142.790 -141.130 -142.110 ;
        RECT -96.610 -142.210 -94.210 -142.110 ;
        RECT -149.220 -152.500 -144.070 -142.790 ;
        RECT -142.520 -142.810 -141.750 -142.790 ;
        RECT -150.510 -152.590 -149.880 -152.530 ;
        RECT -150.510 -153.170 -149.860 -152.590 ;
        RECT -149.210 -153.170 -144.070 -152.500 ;
        RECT -150.510 -153.920 -149.880 -153.170 ;
        RECT -150.510 -154.640 -142.250 -153.920 ;
        RECT -150.510 -154.870 -147.920 -154.640 ;
        RECT -150.510 -154.900 -149.880 -154.870 ;
        RECT -150.030 -156.020 -149.040 -156.010 ;
        RECT -150.430 -156.540 -149.040 -156.020 ;
        RECT -150.430 -160.150 -149.940 -156.540 ;
        RECT -147.230 -157.070 -143.810 -157.020 ;
        RECT -147.240 -157.640 -143.800 -157.070 ;
        RECT -148.650 -167.470 -144.350 -158.410 ;
        RECT -142.670 -158.460 -141.950 -157.910 ;
        RECT -142.670 -158.470 -142.170 -158.460 ;
        RECT -142.520 -167.470 -141.130 -167.450 ;
        RECT -92.670 -167.470 -90.180 -167.390 ;
        RECT -151.050 -169.220 -90.180 -167.470 ;
        RECT -152.000 -169.230 -90.180 -169.220 ;
        RECT -152.160 -169.580 -90.180 -169.230 ;
        RECT -152.000 -169.590 -90.180 -169.580 ;
        RECT -151.050 -169.940 -90.180 -169.590 ;
        RECT -150.680 -170.700 -90.180 -169.940 ;
        RECT -150.680 -171.380 -141.130 -170.700 ;
        RECT -92.670 -170.890 -90.180 -170.700 ;
        RECT -149.220 -181.090 -144.070 -171.380 ;
        RECT -142.520 -171.390 -141.130 -171.380 ;
        RECT -142.520 -171.400 -141.750 -171.390 ;
        RECT -150.510 -181.180 -149.880 -181.120 ;
        RECT -150.510 -181.760 -149.860 -181.180 ;
        RECT -149.210 -181.760 -144.070 -181.090 ;
        RECT -150.510 -182.510 -149.880 -181.760 ;
        RECT -150.510 -183.230 -142.250 -182.510 ;
        RECT -150.510 -183.460 -147.920 -183.230 ;
        RECT -150.510 -183.490 -149.880 -183.460 ;
        RECT -150.030 -184.610 -149.040 -184.600 ;
        RECT -150.430 -185.130 -149.040 -184.610 ;
        RECT -150.430 -188.740 -149.940 -185.130 ;
        RECT -147.230 -185.660 -143.810 -185.610 ;
        RECT -147.240 -186.230 -143.800 -185.660 ;
        RECT -148.650 -196.060 -144.350 -187.000 ;
        RECT -142.670 -187.050 -141.950 -186.500 ;
        RECT -142.670 -187.060 -142.170 -187.050 ;
        RECT -142.520 -196.050 -141.750 -196.040 ;
        RECT -142.520 -196.060 -141.110 -196.050 ;
        RECT -88.200 -196.060 -85.850 -195.960 ;
        RECT -151.050 -197.810 -85.850 -196.060 ;
        RECT -152.000 -197.820 -85.850 -197.810 ;
        RECT -152.160 -198.170 -85.850 -197.820 ;
        RECT -152.000 -198.180 -85.850 -198.170 ;
        RECT -151.050 -198.530 -85.850 -198.180 ;
        RECT -150.680 -199.290 -85.850 -198.530 ;
        RECT -150.680 -199.970 -141.110 -199.290 ;
        RECT -88.200 -199.420 -85.850 -199.290 ;
        RECT -149.220 -209.680 -144.070 -199.970 ;
        RECT -142.520 -199.990 -141.110 -199.970 ;
        RECT -150.510 -209.770 -149.880 -209.710 ;
        RECT -150.510 -210.350 -149.860 -209.770 ;
        RECT -149.210 -210.350 -144.070 -209.680 ;
        RECT -150.510 -211.100 -149.880 -210.350 ;
        RECT -150.510 -211.820 -142.250 -211.100 ;
        RECT -150.510 -212.050 -147.920 -211.820 ;
        RECT -150.510 -212.080 -149.880 -212.050 ;
        RECT -150.030 -213.200 -149.040 -213.190 ;
        RECT -150.430 -213.720 -149.040 -213.200 ;
        RECT -150.430 -217.330 -149.940 -213.720 ;
        RECT -147.230 -214.250 -143.810 -214.200 ;
        RECT -147.240 -214.820 -143.800 -214.250 ;
        RECT -148.650 -224.650 -144.350 -215.590 ;
        RECT -142.670 -215.640 -141.950 -215.090 ;
        RECT -142.670 -215.650 -142.170 -215.640 ;
        RECT -141.750 -224.630 -141.110 -224.620 ;
        RECT -142.520 -224.650 -141.110 -224.630 ;
        RECT -84.200 -224.650 -81.490 -224.590 ;
        RECT -151.050 -226.400 -81.490 -224.650 ;
        RECT -152.000 -226.410 -81.490 -226.400 ;
        RECT -152.160 -226.760 -81.490 -226.410 ;
        RECT -152.000 -226.770 -81.490 -226.760 ;
        RECT -151.050 -227.120 -81.490 -226.770 ;
        RECT -150.680 -227.880 -81.490 -227.120 ;
        RECT -150.680 -228.560 -141.110 -227.880 ;
        RECT -84.200 -228.000 -81.490 -227.880 ;
        RECT -149.220 -238.270 -144.070 -228.560 ;
        RECT -142.520 -228.580 -141.750 -228.560 ;
        RECT -150.510 -238.360 -149.880 -238.300 ;
        RECT -150.510 -238.940 -149.860 -238.360 ;
        RECT -149.210 -238.940 -144.070 -238.270 ;
        RECT -150.510 -239.690 -149.880 -238.940 ;
        RECT -150.510 -240.410 -142.250 -239.690 ;
        RECT -150.510 -240.640 -147.920 -240.410 ;
        RECT -150.510 -240.670 -149.880 -240.640 ;
      LAYER via ;
        RECT -138.110 141.150 -136.080 141.480 ;
        RECT -138.170 140.290 -137.470 140.910 ;
        RECT -114.720 141.150 -111.730 141.500 ;
        RECT -109.520 141.150 -107.490 141.480 ;
        RECT -111.290 140.350 -110.940 141.110 ;
        RECT -109.580 140.290 -108.880 140.910 ;
        RECT -86.130 141.150 -83.140 141.500 ;
        RECT -80.930 141.150 -78.900 141.480 ;
        RECT -112.320 135.060 -111.900 138.230 ;
        RECT -113.290 133.240 -112.770 133.760 ;
        RECT -82.700 140.350 -82.350 141.110 ;
        RECT -80.990 140.290 -80.290 140.910 ;
        RECT -57.540 141.150 -54.550 141.500 ;
        RECT -52.220 141.280 -28.420 141.540 ;
        RECT -83.730 135.060 -83.310 138.230 ;
        RECT -84.700 133.240 -84.180 133.760 ;
        RECT -54.110 140.350 -53.760 141.110 ;
        RECT -55.140 135.060 -54.720 138.230 ;
        RECT -56.110 133.240 -55.590 133.760 ;
        RECT -149.990 129.450 -149.230 129.800 ;
        RECT -150.380 126.020 -150.030 129.010 ;
        RECT -147.110 128.420 -143.940 128.840 ;
        RECT -142.640 127.450 -142.120 127.970 ;
        RECT -68.360 127.360 -65.130 129.610 ;
        RECT -56.170 126.080 -55.650 126.450 ;
        RECT -96.950 122.870 -93.720 125.120 ;
        RECT -127.370 118.600 -125.120 121.830 ;
        RECT -138.900 115.200 -137.040 118.430 ;
        RECT -19.540 141.280 1.320 141.540 ;
        RECT 3.090 141.150 5.120 141.480 ;
        RECT 3.030 140.290 3.730 140.910 ;
        RECT 26.480 141.150 29.470 141.500 ;
        RECT 31.680 141.150 33.710 141.480 ;
        RECT 29.910 140.350 30.260 141.110 ;
        RECT 31.620 140.290 32.320 140.910 ;
        RECT 55.070 141.150 58.060 141.500 ;
        RECT 60.270 141.150 62.300 141.480 ;
        RECT 28.880 135.060 29.300 138.230 ;
        RECT 27.910 133.240 28.430 133.760 ;
        RECT -25.690 128.390 -25.300 128.780 ;
        RECT 58.500 140.350 58.850 141.110 ;
        RECT 60.210 140.290 60.910 140.910 ;
        RECT 83.660 141.150 86.650 141.500 ;
        RECT 88.860 141.150 90.890 141.480 ;
        RECT 57.470 135.060 57.890 138.230 ;
        RECT 56.500 133.240 57.020 133.760 ;
        RECT 87.090 140.350 87.440 141.110 ;
        RECT 88.800 140.290 89.500 140.910 ;
        RECT 112.250 141.150 115.240 141.500 ;
        RECT 117.450 141.150 119.480 141.480 ;
        RECT 86.060 135.060 86.480 138.230 ;
        RECT -52.830 121.700 -52.420 122.110 ;
        RECT -56.310 117.760 -55.790 118.280 ;
        RECT -150.360 102.630 -150.030 104.660 ;
        RECT -149.790 102.570 -149.170 103.270 ;
        RECT -149.990 100.860 -149.230 101.210 ;
        RECT -150.380 97.430 -150.030 100.420 ;
        RECT -147.110 99.830 -143.940 100.250 ;
        RECT -142.640 98.860 -142.120 99.380 ;
        RECT -130.850 86.610 -128.770 89.840 ;
        RECT -23.270 127.470 -23.010 127.730 ;
        RECT -20.410 127.520 -20.150 127.780 ;
        RECT -23.280 126.440 -23.020 126.700 ;
        RECT -22.560 126.410 -22.300 126.670 ;
        RECT -21.870 126.450 -21.610 126.710 ;
        RECT -23.280 125.990 -23.020 126.250 ;
        RECT -21.870 126.010 -21.610 126.270 ;
        RECT -23.280 125.570 -23.020 125.830 ;
        RECT -22.560 125.570 -22.300 125.830 ;
        RECT -21.850 125.590 -21.590 125.850 ;
        RECT -25.610 124.940 -25.220 125.330 ;
        RECT -52.780 116.910 -52.370 117.320 ;
        RECT -56.210 81.740 -55.690 82.260 ;
        RECT -52.780 80.800 -52.370 81.240 ;
        RECT -150.360 74.040 -150.030 76.070 ;
        RECT -149.790 73.980 -149.170 74.680 ;
        RECT -149.990 72.270 -149.230 72.620 ;
        RECT -150.380 68.840 -150.030 71.830 ;
        RECT -147.110 71.240 -143.940 71.660 ;
        RECT -142.640 70.270 -142.120 70.790 ;
        RECT -23.280 124.220 -23.020 124.480 ;
        RECT -24.230 123.770 -23.970 124.030 ;
        RECT -20.720 125.980 -20.460 126.240 ;
        RECT -7.170 125.670 -6.910 125.930 ;
        RECT -5.810 125.750 -5.550 126.010 ;
        RECT -5.120 125.740 -4.860 126.000 ;
        RECT -21.140 123.970 -20.880 124.230 ;
        RECT -22.580 122.770 -22.320 123.030 ;
        RECT -21.150 122.790 -20.890 123.050 ;
        RECT -23.370 122.190 -23.110 122.450 ;
        RECT -22.440 122.190 -22.180 122.450 ;
        RECT -21.740 122.190 -21.480 122.450 ;
        RECT -21.000 122.190 -20.740 122.450 ;
        RECT -20.290 122.180 -20.030 122.440 ;
        RECT -24.310 121.070 -23.890 121.490 ;
        RECT -7.890 122.010 -7.630 122.270 ;
        RECT -18.360 119.670 -18.070 120.250 ;
        RECT -5.070 118.610 -4.810 118.870 ;
        RECT -9.990 112.870 -9.730 113.130 ;
        RECT -8.900 112.880 -8.640 113.140 ;
        RECT -11.150 112.360 -10.890 112.620 ;
        RECT -10.420 112.370 -10.160 112.630 ;
        RECT -9.980 111.880 -9.720 112.140 ;
        RECT -8.890 111.890 -8.630 112.150 ;
        RECT -11.180 111.440 -10.920 111.700 ;
        RECT -10.440 111.450 -10.180 111.710 ;
        RECT -9.980 110.890 -9.720 111.150 ;
        RECT -8.890 110.900 -8.630 111.160 ;
        RECT -11.170 110.520 -10.910 110.780 ;
        RECT -11.820 109.500 -11.560 109.760 ;
        RECT -11.860 108.540 -11.600 108.800 ;
        RECT -11.820 107.580 -11.560 107.840 ;
        RECT -10.460 110.460 -10.200 110.720 ;
        RECT -10.170 109.960 -9.910 110.220 ;
        RECT -8.870 109.860 -8.610 110.120 ;
        RECT -10.200 109.500 -9.940 109.760 ;
        RECT -10.170 108.970 -9.910 109.230 ;
        RECT -8.870 108.870 -8.610 109.130 ;
        RECT -10.200 108.510 -9.940 108.770 ;
        RECT 1.970 122.030 2.230 122.290 ;
        RECT 0.720 118.180 1.030 118.490 ;
        RECT 17.300 125.820 17.720 126.240 ;
        RECT 13.450 125.060 13.870 125.480 ;
        RECT 18.970 123.450 19.410 123.890 ;
        RECT 24.690 123.450 25.130 123.890 ;
        RECT 26.510 123.420 26.950 123.860 ;
        RECT 14.550 122.430 14.990 122.870 ;
        RECT 11.790 119.410 12.050 119.670 ;
        RECT 4.720 118.720 4.980 118.980 ;
        RECT 3.550 117.730 3.820 117.990 ;
        RECT -7.780 116.950 -7.430 117.300 ;
        RECT -2.530 117.260 -2.270 117.520 ;
        RECT 13.240 116.240 13.500 116.500 ;
        RECT 11.140 115.400 11.400 115.660 ;
        RECT -6.760 114.710 -6.500 115.100 ;
        RECT 9.640 114.720 9.970 114.980 ;
        RECT -7.400 113.890 -7.140 114.290 ;
        RECT -10.170 107.980 -9.910 108.240 ;
        RECT -8.870 107.880 -8.610 108.140 ;
        RECT -10.200 107.520 -9.940 107.780 ;
        RECT -11.860 92.300 -11.600 92.770 ;
        RECT -11.220 92.300 -10.960 92.770 ;
        RECT -13.220 91.270 -12.960 91.530 ;
        RECT -13.740 90.870 -13.480 91.130 ;
        RECT -23.020 89.620 -22.360 90.280 ;
        RECT -11.140 91.250 -10.880 91.510 ;
        RECT -9.380 91.260 -9.110 91.530 ;
        RECT -11.800 90.890 -11.540 91.150 ;
        RECT -11.050 90.290 -10.790 90.550 ;
        RECT -10.400 90.290 -10.140 90.550 ;
        RECT -12.270 89.850 -12.010 90.110 ;
        RECT -11.570 89.850 -11.310 90.110 ;
        RECT -9.890 89.120 -9.630 89.380 ;
        RECT -12.720 88.500 -12.460 88.760 ;
        RECT -13.720 86.960 -13.460 87.220 ;
        RECT -17.810 85.100 -17.440 85.470 ;
        RECT -22.980 83.760 -22.320 84.420 ;
        RECT -9.970 87.990 -9.710 88.250 ;
        RECT -8.880 90.870 -8.620 91.130 ;
        RECT -9.960 87.450 -9.700 87.710 ;
        RECT -12.720 86.950 -12.460 87.210 ;
        RECT -9.910 86.500 -9.650 86.760 ;
        RECT -12.240 85.970 -11.980 86.230 ;
        RECT -11.550 85.960 -11.290 86.220 ;
        RECT -11.070 85.190 -10.810 85.450 ;
        RECT -10.360 85.130 -10.100 85.390 ;
        RECT -11.050 80.110 -10.790 80.370 ;
        RECT -14.360 79.670 -14.100 79.930 ;
        RECT -13.260 79.680 -13.000 79.940 ;
        RECT -12.170 79.680 -11.910 79.940 ;
        RECT -11.040 79.640 -10.780 79.900 ;
        RECT -17.820 78.860 -17.450 79.230 ;
        RECT -13.810 79.000 -13.550 79.260 ;
        RECT -12.710 79.000 -12.450 79.260 ;
        RECT -11.610 79.000 -11.350 79.260 ;
        RECT -10.280 78.440 -10.020 78.800 ;
        RECT -13.810 77.630 -13.550 77.890 ;
        RECT -12.710 77.630 -12.450 77.890 ;
        RECT -11.610 77.630 -11.350 77.890 ;
        RECT -14.360 76.900 -14.100 77.160 ;
        RECT -13.260 76.900 -13.000 77.160 ;
        RECT -12.170 76.900 -11.910 77.160 ;
        RECT -14.370 75.560 -14.110 75.820 ;
        RECT -13.260 75.550 -13.000 75.810 ;
        RECT -12.170 75.530 -11.910 75.790 ;
        RECT -13.810 74.860 -13.550 75.120 ;
        RECT -12.710 74.850 -12.450 75.110 ;
        RECT -11.620 74.850 -11.360 75.110 ;
        RECT -14.830 73.200 -14.540 73.490 ;
        RECT -11.010 72.560 -10.750 72.820 ;
        RECT -7.380 112.780 -7.120 113.040 ;
        RECT -7.380 111.860 -7.120 112.120 ;
        RECT -7.410 110.940 -7.150 111.200 ;
        RECT 9.010 113.000 9.340 113.330 ;
        RECT 8.440 111.520 8.770 111.850 ;
        RECT -6.770 109.850 -6.510 110.110 ;
        RECT 7.800 109.920 8.130 110.250 ;
        RECT 7.160 109.350 7.490 109.680 ;
        RECT -6.760 108.890 -6.500 109.150 ;
        RECT -6.770 107.930 -6.510 108.190 ;
        RECT -7.410 90.270 -7.150 90.530 ;
        RECT -8.030 89.120 -7.770 89.380 ;
        RECT -8.450 86.510 -8.190 86.770 ;
        RECT -8.010 80.820 -7.750 81.240 ;
        RECT -8.050 78.440 -7.790 78.800 ;
        RECT 6.550 107.780 6.880 108.110 ;
        RECT 5.920 106.250 6.250 106.580 ;
        RECT 5.360 104.680 5.690 105.010 ;
        RECT 4.740 99.210 5.070 99.540 ;
        RECT 4.110 97.620 4.440 97.950 ;
        RECT 3.490 96.070 3.820 96.400 ;
        RECT 2.890 94.590 3.220 94.920 ;
        RECT 2.250 89.420 2.580 89.750 ;
        RECT 1.580 87.850 1.910 88.180 ;
        RECT -6.770 85.940 -6.510 86.200 ;
        RECT 0.960 86.210 1.290 86.540 ;
        RECT -7.430 74.810 -7.170 75.140 ;
        RECT -8.460 73.190 -8.170 73.480 ;
        RECT -14.320 72.120 -14.060 72.380 ;
        RECT -13.220 72.130 -12.960 72.390 ;
        RECT -12.130 72.130 -11.870 72.390 ;
        RECT -11.000 72.090 -10.740 72.350 ;
        RECT -9.620 72.180 -9.020 72.780 ;
        RECT -13.770 71.450 -13.510 71.710 ;
        RECT -12.670 71.450 -12.410 71.710 ;
        RECT -11.570 71.450 -11.310 71.710 ;
        RECT -13.770 70.080 -13.510 70.340 ;
        RECT -12.670 70.080 -12.410 70.340 ;
        RECT -11.570 70.080 -11.310 70.340 ;
        RECT -14.320 69.350 -14.060 69.610 ;
        RECT -13.220 69.350 -12.960 69.610 ;
        RECT -12.130 69.350 -11.870 69.610 ;
        RECT -14.330 68.010 -14.070 68.270 ;
        RECT -13.220 68.000 -12.960 68.260 ;
        RECT -12.130 67.980 -11.870 68.240 ;
        RECT 0.280 84.770 0.610 85.100 ;
        RECT -3.760 80.410 -3.180 81.120 ;
        RECT -13.770 67.310 -13.510 67.570 ;
        RECT -12.670 67.300 -12.410 67.560 ;
        RECT -11.580 67.300 -11.320 67.560 ;
        RECT -6.840 67.250 -6.580 67.590 ;
        RECT -25.750 66.310 -25.360 66.700 ;
        RECT -126.950 58.020 -124.870 61.250 ;
        RECT 0.250 60.940 0.680 61.370 ;
        RECT 0.900 60.150 1.330 60.580 ;
        RECT 1.570 59.470 1.970 59.870 ;
        RECT 1.400 58.530 1.910 59.040 ;
        RECT 11.140 113.650 11.400 113.910 ;
        RECT 11.140 111.900 11.400 112.160 ;
        RECT 11.140 110.150 11.400 110.410 ;
        RECT 11.140 109.360 11.400 109.620 ;
        RECT 11.140 107.610 11.400 107.870 ;
        RECT 11.140 105.860 11.400 106.120 ;
        RECT 11.140 104.110 11.400 104.370 ;
        RECT 16.960 116.250 17.220 116.510 ;
        RECT 18.000 116.290 18.260 116.550 ;
        RECT 13.240 114.490 13.500 114.750 ;
        RECT 13.240 112.740 13.500 113.000 ;
        RECT 13.240 110.990 13.500 111.250 ;
        RECT 13.240 108.520 13.500 108.780 ;
        RECT 13.240 106.770 13.500 107.030 ;
        RECT 13.240 105.020 13.500 105.280 ;
        RECT 15.280 115.520 15.540 115.780 ;
        RECT 16.960 114.500 17.220 114.760 ;
        RECT 18.000 114.540 18.260 114.800 ;
        RECT 15.280 113.770 15.540 114.030 ;
        RECT 16.960 112.750 17.220 113.010 ;
        RECT 18.000 112.790 18.260 113.050 ;
        RECT 15.280 112.020 15.540 112.280 ;
        RECT 16.960 111.000 17.220 111.260 ;
        RECT 18.000 111.040 18.260 111.300 ;
        RECT 15.280 110.270 15.540 110.530 ;
        RECT 15.280 109.240 15.540 109.500 ;
        RECT 16.960 108.510 17.220 108.770 ;
        RECT 18.000 108.470 18.260 108.730 ;
        RECT 15.280 107.490 15.540 107.750 ;
        RECT 16.960 106.760 17.220 107.020 ;
        RECT 18.000 106.720 18.260 106.980 ;
        RECT 15.280 105.740 15.540 106.000 ;
        RECT 16.960 105.010 17.220 105.270 ;
        RECT 18.000 104.970 18.260 105.230 ;
        RECT 15.280 103.990 15.540 104.250 ;
        RECT 13.240 103.270 13.500 103.530 ;
        RECT 16.960 103.260 17.220 103.520 ;
        RECT 18.000 103.220 18.260 103.480 ;
        RECT 11.140 99.230 11.400 99.490 ;
        RECT 11.140 97.480 11.400 97.740 ;
        RECT 11.140 95.730 11.400 95.990 ;
        RECT 11.140 93.980 11.400 94.240 ;
        RECT 13.240 98.390 13.500 98.650 ;
        RECT 13.240 96.640 13.500 96.900 ;
        RECT 13.240 94.890 13.500 95.150 ;
        RECT 15.280 99.110 15.540 99.370 ;
        RECT 16.960 98.380 17.220 98.640 ;
        RECT 18.000 98.340 18.260 98.600 ;
        RECT 15.280 97.360 15.540 97.620 ;
        RECT 16.960 96.630 17.220 96.890 ;
        RECT 18.000 96.590 18.260 96.850 ;
        RECT 15.280 95.610 15.540 95.870 ;
        RECT 16.960 94.880 17.220 95.140 ;
        RECT 18.000 94.840 18.260 95.100 ;
        RECT 15.280 93.860 15.540 94.120 ;
        RECT 11.100 90.170 11.360 90.430 ;
        RECT 13.240 93.140 13.500 93.400 ;
        RECT 16.960 93.130 17.220 93.390 ;
        RECT 18.000 93.090 18.260 93.350 ;
        RECT 20.260 122.430 20.700 122.870 ;
        RECT 21.160 109.300 21.420 109.560 ;
        RECT 20.070 108.780 20.330 109.040 ;
        RECT 20.070 107.510 20.330 107.770 ;
        RECT 21.160 106.990 21.420 107.250 ;
        RECT 21.160 106.100 21.420 106.360 ;
        RECT 20.070 105.580 20.330 105.840 ;
        RECT 20.070 104.310 20.330 104.570 ;
        RECT 21.160 103.790 21.420 104.050 ;
        RECT 85.090 133.240 85.610 133.760 ;
        RECT 115.680 140.350 116.030 141.110 ;
        RECT 117.390 140.290 118.090 140.910 ;
        RECT 140.840 141.150 143.830 141.500 ;
        RECT 146.040 141.150 148.070 141.480 ;
        RECT 114.650 135.060 115.070 138.230 ;
        RECT 37.070 125.060 38.420 125.480 ;
        RECT 31.650 122.420 32.600 122.830 ;
        RECT 34.660 122.430 35.100 122.870 ;
        RECT 28.910 118.650 29.170 118.910 ;
        RECT 27.030 115.120 27.290 115.380 ;
        RECT 26.520 112.750 26.780 113.010 ;
        RECT 23.570 109.300 23.830 109.560 ;
        RECT 32.500 117.740 32.760 118.000 ;
        RECT 29.370 116.720 29.630 116.980 ;
        RECT 28.480 112.260 28.740 112.520 ;
        RECT 28.090 110.730 28.350 110.990 ;
        RECT 29.790 114.630 30.050 114.890 ;
        RECT 27.380 109.900 27.640 110.160 ;
        RECT 30.850 114.150 31.110 114.410 ;
        RECT 28.080 109.040 28.340 109.300 ;
        RECT 23.570 106.990 23.830 107.250 ;
        RECT 28.480 107.530 28.740 107.790 ;
        RECT 35.670 118.660 35.930 118.920 ;
        RECT 35.230 117.750 35.490 118.010 ;
        RECT 32.490 107.050 32.760 107.320 ;
        RECT 34.740 107.070 35.000 107.330 ;
        RECT 26.570 106.700 26.830 106.960 ;
        RECT 23.570 106.100 23.830 106.360 ;
        RECT 23.570 103.790 23.830 104.050 ;
        RECT 28.490 106.230 28.750 106.490 ;
        RECT 28.340 105.270 28.600 105.530 ;
        RECT 27.400 104.160 27.660 104.420 ;
        RECT 27.400 103.560 27.660 103.820 ;
        RECT 28.340 102.510 28.600 102.770 ;
        RECT 28.490 101.500 28.750 101.760 ;
        RECT 21.140 98.830 21.400 99.090 ;
        RECT 20.050 98.310 20.310 98.570 ;
        RECT 20.050 97.040 20.310 97.300 ;
        RECT 21.140 96.520 21.400 96.780 ;
        RECT 21.140 95.630 21.400 95.890 ;
        RECT 20.050 95.110 20.310 95.370 ;
        RECT 20.050 93.840 20.310 94.100 ;
        RECT 23.550 98.830 23.810 99.090 ;
        RECT 27.950 99.100 28.210 99.360 ;
        RECT 29.130 100.410 29.410 100.690 ;
        RECT 40.460 122.390 40.900 122.830 ;
        RECT 48.790 123.420 49.070 123.860 ;
        RECT 45.010 116.760 46.230 117.020 ;
        RECT 41.770 116.110 42.030 116.370 ;
        RECT 48.100 115.570 48.360 115.830 ;
        RECT 46.810 112.260 47.070 112.520 ;
        RECT 50.440 118.660 50.700 118.920 ;
        RECT 49.550 117.790 49.810 118.050 ;
        RECT 113.680 133.240 114.200 133.760 ;
        RECT 144.270 140.350 144.620 141.110 ;
        RECT 145.980 140.290 146.680 140.910 ;
        RECT 169.430 141.150 172.420 141.500 ;
        RECT 174.630 141.150 176.660 141.480 ;
        RECT 143.240 135.060 143.660 138.230 ;
        RECT 142.270 133.240 142.790 133.760 ;
        RECT 172.860 140.350 173.210 141.110 ;
        RECT 174.570 140.290 175.270 140.910 ;
        RECT 198.020 141.150 201.010 141.500 ;
        RECT 171.830 135.060 172.250 138.230 ;
        RECT 170.860 133.240 171.380 133.760 ;
        RECT 201.450 140.350 201.800 141.110 ;
        RECT 200.420 135.060 200.840 138.230 ;
        RECT 199.450 133.240 199.970 133.760 ;
        RECT 56.960 127.760 57.330 128.130 ;
        RECT 53.110 119.370 53.370 119.640 ;
        RECT 49.550 113.580 49.810 113.840 ;
        RECT 50.570 113.590 50.830 113.850 ;
        RECT 48.790 112.750 49.050 113.010 ;
        RECT 50.520 112.740 50.780 113.000 ;
        RECT 51.500 112.490 51.760 112.750 ;
        RECT 50.670 111.910 50.930 112.170 ;
        RECT 51.450 111.840 51.710 112.100 ;
        RECT 46.960 111.300 47.220 111.560 ;
        RECT 47.900 110.190 48.160 110.450 ;
        RECT 47.900 109.590 48.160 109.850 ;
        RECT 49.560 111.380 49.820 111.640 ;
        RECT 50.730 110.900 50.990 111.160 ;
        RECT 51.450 110.990 51.710 111.250 ;
        RECT 48.840 109.910 49.100 110.170 ;
        RECT 50.290 110.100 50.550 110.360 ;
        RECT 46.960 108.540 47.220 108.800 ;
        RECT 40.540 107.070 40.800 107.330 ;
        RECT 35.600 105.680 35.860 105.940 ;
        RECT 34.810 103.630 35.070 103.890 ;
        RECT 35.630 101.990 35.890 102.250 ;
        RECT 46.810 107.530 47.070 107.790 ;
        RECT 46.810 106.230 47.070 106.490 ;
        RECT 51.500 110.340 51.760 110.600 ;
        RECT 51.500 109.490 51.760 109.750 ;
        RECT 51.450 108.840 51.710 109.100 ;
        RECT 51.450 107.990 51.710 108.250 ;
        RECT 50.930 107.220 51.190 107.480 ;
        RECT 51.500 107.340 51.760 107.600 ;
        RECT 53.320 113.470 53.750 113.900 ;
        RECT 48.770 106.690 49.030 106.950 ;
        RECT 50.520 106.710 50.780 106.970 ;
        RECT 51.500 106.460 51.760 106.720 ;
        RECT 50.670 105.880 50.930 106.140 ;
        RECT 51.450 105.810 51.710 106.070 ;
        RECT 46.960 105.270 47.220 105.530 ;
        RECT 40.510 103.570 40.770 103.830 ;
        RECT 47.900 104.160 48.160 104.420 ;
        RECT 47.900 103.560 48.160 103.820 ;
        RECT 49.560 105.350 49.820 105.610 ;
        RECT 50.730 104.870 50.990 105.130 ;
        RECT 51.450 104.960 51.710 105.220 ;
        RECT 48.840 103.880 49.100 104.140 ;
        RECT 50.290 104.070 50.550 104.330 ;
        RECT 46.960 102.510 47.220 102.770 ;
        RECT 40.510 101.050 40.770 101.310 ;
        RECT 29.890 98.780 30.150 99.040 ;
        RECT 23.550 96.520 23.810 96.780 ;
        RECT 29.890 98.230 30.150 98.490 ;
        RECT 23.550 95.630 23.810 95.890 ;
        RECT 29.890 97.240 30.150 97.500 ;
        RECT 29.890 96.690 30.150 96.950 ;
        RECT 29.890 95.540 30.150 95.800 ;
        RECT 21.140 93.320 21.400 93.580 ;
        RECT 23.550 93.320 23.810 93.580 ;
        RECT 29.890 94.990 30.150 95.250 ;
        RECT 30.810 94.570 31.070 94.830 ;
        RECT 29.890 94.010 30.150 94.270 ;
        RECT 34.740 94.530 35.000 94.790 ;
        RECT 29.890 93.460 30.150 93.720 ;
        RECT 15.240 90.050 15.500 90.310 ;
        RECT 11.100 88.420 11.360 88.680 ;
        RECT 11.100 86.670 11.360 86.930 ;
        RECT 11.100 84.920 11.360 85.180 ;
        RECT 21.760 92.220 22.020 92.630 ;
        RECT 13.200 89.330 13.460 89.590 ;
        RECT 13.200 87.580 13.460 87.840 ;
        RECT 13.200 85.830 13.460 86.090 ;
        RECT 13.200 84.080 13.460 84.340 ;
        RECT 16.920 89.320 17.180 89.580 ;
        RECT 17.960 89.280 18.220 89.540 ;
        RECT 15.240 88.300 15.500 88.560 ;
        RECT 16.920 87.570 17.180 87.830 ;
        RECT 17.960 87.530 18.220 87.790 ;
        RECT 15.240 86.550 15.500 86.810 ;
        RECT 16.920 85.820 17.180 86.080 ;
        RECT 17.960 85.780 18.220 86.040 ;
        RECT 15.240 84.800 15.500 85.060 ;
        RECT 16.920 84.070 17.180 84.330 ;
        RECT 17.960 84.030 18.220 84.290 ;
        RECT 21.170 89.560 21.430 89.820 ;
        RECT 20.080 89.040 20.340 89.300 ;
        RECT 20.080 87.770 20.340 88.030 ;
        RECT 21.170 87.250 21.430 87.510 ;
        RECT 21.170 86.360 21.430 86.620 ;
        RECT 20.080 85.840 20.340 86.100 ;
        RECT 20.080 84.570 20.340 84.830 ;
        RECT 21.170 84.050 21.430 84.310 ;
        RECT 23.580 89.560 23.840 89.820 ;
        RECT 46.810 101.500 47.070 101.760 ;
        RECT 51.500 104.310 51.760 104.570 ;
        RECT 51.500 103.460 51.760 103.720 ;
        RECT 51.450 102.810 51.710 103.070 ;
        RECT 51.450 101.960 51.710 102.220 ;
        RECT 46.480 99.840 46.740 100.100 ;
        RECT 45.390 98.780 45.650 99.040 ;
        RECT 50.950 101.180 51.220 101.440 ;
        RECT 51.500 101.310 51.760 101.570 ;
        RECT 53.750 112.510 54.010 112.770 ;
        RECT 53.800 110.290 54.060 110.550 ;
        RECT 53.790 109.570 54.050 109.830 ;
        RECT 53.710 107.320 53.970 107.580 ;
        RECT 53.750 106.480 54.010 106.740 ;
        RECT 53.800 104.260 54.060 104.520 ;
        RECT 53.790 103.540 54.050 103.800 ;
        RECT 53.710 101.290 53.970 101.550 ;
        RECT 57.780 124.300 58.150 124.670 ;
        RECT 56.970 100.390 57.340 100.760 ;
        RECT 58.550 119.590 58.920 119.960 ;
        RECT 45.390 98.230 45.650 98.490 ;
        RECT 57.740 99.800 58.110 100.170 ;
        RECT 47.350 99.110 47.610 99.370 ;
        RECT 40.540 94.530 40.800 94.790 ;
        RECT 45.390 97.240 45.650 97.500 ;
        RECT 65.100 118.540 65.600 119.040 ;
        RECT 61.880 116.980 62.380 117.480 ;
        RECT 62.830 117.470 63.330 117.970 ;
        RECT 63.910 117.940 64.410 118.440 ;
        RECT 59.430 114.520 59.800 114.890 ;
        RECT 45.390 96.690 45.650 96.950 ;
        RECT 58.480 97.470 58.850 97.840 ;
        RECT 45.390 95.540 45.650 95.800 ;
        RECT 45.390 94.990 45.650 95.250 ;
        RECT 44.470 94.570 44.730 94.830 ;
        RECT 45.390 94.010 45.650 94.270 ;
        RECT 45.390 93.460 45.650 93.720 ;
        RECT 29.920 89.450 30.180 89.710 ;
        RECT 30.530 89.350 30.790 89.610 ;
        RECT 26.160 88.500 26.420 88.760 ;
        RECT 23.580 87.250 23.840 87.510 ;
        RECT 23.580 86.360 23.840 86.620 ;
        RECT 23.580 84.050 23.840 84.310 ;
        RECT 27.240 87.800 27.500 88.060 ;
        RECT 29.920 88.900 30.180 89.160 ;
        RECT 30.510 88.300 30.770 88.560 ;
        RECT 27.220 86.790 27.480 87.050 ;
        RECT 26.790 85.720 27.050 85.980 ;
        RECT 19.580 83.370 19.840 83.630 ;
        RECT 19.040 83.000 19.330 83.290 ;
        RECT 14.600 82.490 14.910 82.800 ;
        RECT 26.190 83.410 26.450 83.670 ;
        RECT 27.170 84.750 27.430 85.010 ;
        RECT 27.220 83.790 27.480 84.050 ;
        RECT 27.220 83.400 27.480 83.660 ;
        RECT 24.790 83.000 25.050 83.260 ;
        RECT 26.760 83.080 27.020 83.340 ;
        RECT 18.410 81.780 18.830 82.200 ;
        RECT 14.560 80.820 14.980 81.240 ;
        RECT 20.470 82.460 20.730 82.720 ;
        RECT 19.880 81.790 20.140 82.050 ;
        RECT 20.970 81.790 21.230 82.050 ;
        RECT 22.070 81.780 22.330 82.040 ;
        RECT 29.920 87.930 30.180 88.190 ;
        RECT 29.920 87.380 30.180 87.640 ;
        RECT 29.920 86.210 30.180 86.470 ;
        RECT 30.510 86.420 30.770 86.680 ;
        RECT 29.920 85.660 30.180 85.920 ;
        RECT 30.380 85.240 30.640 85.500 ;
        RECT 30.960 85.160 31.220 85.420 ;
        RECT 29.920 84.680 30.180 84.940 ;
        RECT 29.920 84.130 30.180 84.390 ;
        RECT 29.000 83.020 29.260 83.280 ;
        RECT 24.910 81.780 25.170 82.040 ;
        RECT 26.010 81.790 26.270 82.050 ;
        RECT 27.100 81.790 27.360 82.050 ;
        RECT 27.800 81.770 28.130 82.100 ;
        RECT 34.980 85.140 35.250 85.400 ;
        RECT 59.410 92.220 59.780 92.630 ;
        RECT 38.610 89.150 38.870 89.410 ;
        RECT 38.760 88.470 39.020 88.730 ;
        RECT 38.760 87.580 39.020 87.840 ;
        RECT 38.610 86.900 38.870 87.160 ;
        RECT 38.610 86.380 38.870 86.640 ;
        RECT 38.760 85.700 39.020 85.960 ;
        RECT 38.760 84.810 39.020 85.070 ;
        RECT 38.610 84.130 38.870 84.390 ;
        RECT 46.040 88.480 46.300 88.740 ;
        RECT 45.520 87.550 45.780 87.810 ;
        RECT 45.050 85.710 45.310 85.970 ;
        RECT 40.890 85.250 41.160 85.520 ;
        RECT 37.840 83.330 38.190 83.680 ;
        RECT 30.990 82.600 31.250 82.860 ;
        RECT 35.030 82.570 35.300 82.840 ;
        RECT 28.950 81.700 29.290 82.040 ;
        RECT 29.690 81.820 29.950 82.080 ;
        RECT 30.780 81.820 31.040 82.080 ;
        RECT 31.880 81.810 32.140 82.070 ;
        RECT 20.430 81.110 20.690 81.370 ;
        RECT 21.520 81.090 21.780 81.350 ;
        RECT 22.630 81.080 22.890 81.340 ;
        RECT 19.090 80.730 19.410 81.050 ;
        RECT 20.430 79.740 20.690 80.000 ;
        RECT 21.520 79.740 21.780 80.000 ;
        RECT 22.620 79.740 22.880 80.000 ;
        RECT 19.870 79.010 20.130 79.270 ;
        RECT 20.970 79.010 21.230 79.270 ;
        RECT 22.070 79.010 22.330 79.270 ;
        RECT 19.870 77.640 20.130 77.900 ;
        RECT 20.970 77.640 21.230 77.900 ;
        RECT 22.070 77.640 22.330 77.900 ;
        RECT 19.300 77.000 19.560 77.260 ;
        RECT 20.430 76.960 20.690 77.220 ;
        RECT 21.520 76.960 21.780 77.220 ;
        RECT 22.620 76.970 22.880 77.230 ;
        RECT 19.310 76.530 19.570 76.790 ;
        RECT 24.350 81.080 24.610 81.340 ;
        RECT 25.460 81.090 25.720 81.350 ;
        RECT 26.550 81.110 26.810 81.370 ;
        RECT 30.240 81.140 30.500 81.400 ;
        RECT 34.720 81.810 34.980 82.070 ;
        RECT 35.820 81.820 36.080 82.080 ;
        RECT 36.910 81.820 37.170 82.080 ;
        RECT 44.550 84.780 44.810 85.040 ;
        RECT 37.880 81.560 38.140 81.880 ;
        RECT 31.330 81.120 31.590 81.380 ;
        RECT 32.440 81.110 32.700 81.370 ;
        RECT 24.360 79.740 24.620 80.000 ;
        RECT 25.460 79.740 25.720 80.000 ;
        RECT 26.550 79.740 26.810 80.000 ;
        RECT 30.240 79.770 30.500 80.030 ;
        RECT 31.330 79.770 31.590 80.030 ;
        RECT 32.430 79.770 32.690 80.030 ;
        RECT 24.910 79.010 25.170 79.270 ;
        RECT 26.010 79.010 26.270 79.270 ;
        RECT 27.110 79.010 27.370 79.270 ;
        RECT 29.680 79.040 29.940 79.300 ;
        RECT 30.780 79.040 31.040 79.300 ;
        RECT 31.880 79.040 32.140 79.300 ;
        RECT 24.910 77.640 25.170 77.900 ;
        RECT 26.010 77.640 26.270 77.900 ;
        RECT 27.110 77.640 27.370 77.900 ;
        RECT 29.680 77.670 29.940 77.930 ;
        RECT 30.780 77.670 31.040 77.930 ;
        RECT 31.880 77.670 32.140 77.930 ;
        RECT 24.360 76.970 24.620 77.230 ;
        RECT 25.460 76.960 25.720 77.220 ;
        RECT 26.550 76.960 26.810 77.220 ;
        RECT 27.680 77.000 27.940 77.260 ;
        RECT 27.670 76.530 27.930 76.790 ;
        RECT 23.110 75.980 23.390 76.260 ;
        RECT 23.850 76.000 24.130 76.280 ;
        RECT 19.190 74.950 19.650 75.410 ;
        RECT 29.110 77.030 29.370 77.290 ;
        RECT 30.240 76.990 30.500 77.250 ;
        RECT 31.330 76.990 31.590 77.250 ;
        RECT 32.430 77.000 32.690 77.260 ;
        RECT 29.120 76.560 29.380 76.820 ;
        RECT 27.570 74.000 28.030 74.460 ;
        RECT 34.160 81.110 34.420 81.370 ;
        RECT 35.270 81.120 35.530 81.380 ;
        RECT 36.360 81.140 36.620 81.400 ;
        RECT 40.460 81.800 40.720 82.060 ;
        RECT 41.560 81.810 41.820 82.070 ;
        RECT 42.650 81.810 42.910 82.070 ;
        RECT 43.870 81.780 44.130 82.120 ;
        RECT 39.300 80.850 39.680 81.230 ;
        RECT 39.900 81.100 40.160 81.360 ;
        RECT 41.010 81.110 41.270 81.370 ;
        RECT 42.100 81.130 42.360 81.390 ;
        RECT 34.170 79.770 34.430 80.030 ;
        RECT 35.270 79.770 35.530 80.030 ;
        RECT 36.360 79.770 36.620 80.030 ;
        RECT 39.910 79.760 40.170 80.020 ;
        RECT 41.010 79.760 41.270 80.020 ;
        RECT 42.100 79.760 42.360 80.020 ;
        RECT 34.720 79.040 34.980 79.300 ;
        RECT 35.820 79.040 36.080 79.300 ;
        RECT 36.920 79.040 37.180 79.300 ;
        RECT 40.460 79.030 40.720 79.290 ;
        RECT 41.560 79.030 41.820 79.290 ;
        RECT 42.660 79.030 42.920 79.290 ;
        RECT 34.720 77.670 34.980 77.930 ;
        RECT 35.820 77.670 36.080 77.930 ;
        RECT 36.920 77.670 37.180 77.930 ;
        RECT 40.460 77.660 40.720 77.920 ;
        RECT 41.560 77.660 41.820 77.920 ;
        RECT 42.660 77.660 42.920 77.920 ;
        RECT 34.170 77.000 34.430 77.260 ;
        RECT 35.270 76.990 35.530 77.250 ;
        RECT 32.920 75.980 33.200 76.260 ;
        RECT 36.360 76.990 36.620 77.250 ;
        RECT 37.490 77.030 37.750 77.290 ;
        RECT 39.910 76.990 40.170 77.250 ;
        RECT 41.010 76.980 41.270 77.240 ;
        RECT 42.100 76.980 42.360 77.240 ;
        RECT 43.230 77.020 43.490 77.280 ;
        RECT 73.910 115.600 75.190 116.880 ;
        RECT 78.230 113.440 78.490 113.870 ;
        RECT 74.400 112.160 74.660 112.580 ;
        RECT 70.400 108.960 70.800 109.360 ;
        RECT 65.010 96.260 65.510 96.760 ;
        RECT 63.930 91.070 64.430 91.540 ;
        RECT 62.800 85.880 63.300 86.380 ;
        RECT 61.750 80.580 62.250 81.080 ;
        RECT 46.020 79.070 46.280 79.570 ;
        RECT 45.480 78.170 45.740 78.670 ;
        RECT 45.010 77.270 45.270 77.770 ;
        RECT 37.480 76.560 37.740 76.820 ;
        RECT 43.220 76.550 43.480 76.810 ;
        RECT 29.000 73.110 29.460 73.570 ;
        RECT 37.390 72.200 37.850 72.660 ;
        RECT 11.320 69.970 11.580 71.090 ;
        RECT 23.430 71.030 24.550 71.050 ;
        RECT 22.690 69.930 24.550 71.030 ;
        RECT 22.690 69.910 23.810 69.930 ;
        RECT 32.500 69.880 34.360 71.070 ;
        RECT 9.640 65.680 9.970 66.010 ;
        RECT 9.020 65.060 9.350 65.390 ;
        RECT 8.390 64.430 8.720 64.760 ;
        RECT 7.790 63.800 8.120 64.130 ;
        RECT 7.150 63.120 7.480 63.450 ;
        RECT 6.550 62.500 6.880 62.830 ;
        RECT 5.950 61.860 6.280 62.190 ;
        RECT 5.370 61.290 5.700 61.620 ;
        RECT 4.790 60.600 5.120 60.930 ;
        RECT 4.140 59.960 4.470 60.290 ;
        RECT 3.500 59.310 3.830 59.650 ;
        RECT 2.920 58.670 3.290 59.040 ;
        RECT 44.530 76.370 44.790 76.870 ;
        RECT 67.990 83.100 68.490 83.600 ;
        RECT 65.120 74.990 65.620 75.490 ;
        RECT 63.930 74.040 64.430 74.500 ;
        RECT 62.800 73.170 63.300 73.630 ;
        RECT 61.870 72.260 62.370 72.720 ;
        RECT 67.410 69.970 68.350 71.090 ;
        RECT 43.200 66.340 43.530 66.670 ;
        RECT 71.380 108.320 71.740 108.680 ;
        RECT 70.460 65.150 70.860 65.550 ;
        RECT 72.300 105.950 72.690 106.340 ;
        RECT 71.370 64.350 71.760 64.740 ;
        RECT 73.130 105.390 73.510 105.650 ;
        RECT 72.300 63.530 72.690 63.920 ;
        RECT 79.210 110.030 79.470 110.290 ;
        RECT 80.780 110.030 81.040 110.290 ;
        RECT 77.860 109.050 78.120 109.310 ;
        RECT 101.430 128.670 104.660 130.730 ;
        RECT 130.020 123.780 132.080 127.080 ;
        RECT 85.180 120.930 85.890 121.640 ;
        RECT 77.860 108.440 78.120 108.700 ;
        RECT 80.130 109.120 80.390 109.380 ;
        RECT 81.140 109.110 81.400 109.370 ;
        RECT 80.130 108.370 80.390 108.630 ;
        RECT 81.140 108.380 81.400 108.640 ;
        RECT 79.210 107.460 79.470 107.720 ;
        RECT 80.780 107.460 81.040 107.720 ;
        RECT 79.210 106.830 79.470 107.090 ;
        RECT 80.780 106.830 81.040 107.090 ;
        RECT 77.860 105.850 78.120 106.110 ;
        RECT 77.860 105.240 78.120 105.500 ;
        RECT 80.130 105.920 80.390 106.180 ;
        RECT 81.140 105.910 81.400 106.170 ;
        RECT 80.130 105.170 80.390 105.430 ;
        RECT 81.140 105.180 81.400 105.440 ;
        RECT 79.210 104.260 79.470 104.520 ;
        RECT 80.780 104.260 81.040 104.520 ;
        RECT 158.610 119.530 161.840 121.590 ;
        RECT 212.820 128.730 213.580 129.080 ;
        RECT 207.530 127.700 210.700 128.120 ;
        RECT 205.710 126.730 206.230 127.250 ;
        RECT 187.200 115.120 190.430 117.170 ;
        RECT 213.620 125.300 213.970 128.290 ;
        RECT 201.540 114.480 203.530 117.710 ;
        RECT 84.990 101.140 85.700 101.850 ;
        RECT 109.800 113.500 112.020 113.820 ;
        RECT 212.760 101.850 213.380 102.550 ;
        RECT 213.620 101.910 213.950 103.940 ;
        RECT 212.820 100.140 213.580 100.490 ;
        RECT 207.530 99.110 210.700 99.530 ;
        RECT 205.710 98.140 206.230 98.660 ;
        RECT 213.620 96.710 213.970 99.700 ;
        RECT 192.990 85.890 195.080 89.120 ;
        RECT 80.790 83.090 81.300 83.600 ;
        RECT 109.640 83.110 113.920 84.200 ;
        RECT 80.000 73.280 80.260 73.540 ;
        RECT 80.000 72.610 80.260 72.870 ;
        RECT 80.160 71.370 80.420 71.630 ;
        RECT 75.220 68.040 75.480 68.300 ;
        RECT 80.160 69.760 80.420 70.020 ;
        RECT 80.150 68.150 80.410 68.410 ;
        RECT 80.160 66.530 80.420 66.790 ;
        RECT 80.150 64.920 80.410 65.180 ;
        RECT 73.120 62.740 73.500 63.120 ;
        RECT 79.740 63.270 80.000 63.530 ;
        RECT 80.150 61.720 80.410 61.980 ;
        RECT 76.910 60.010 77.170 60.270 ;
        RECT 77.850 60.010 78.110 60.270 ;
        RECT 78.800 59.990 79.060 60.250 ;
        RECT 80.110 60.010 80.370 60.270 ;
        RECT -150.360 45.450 -150.030 47.480 ;
        RECT -149.790 45.390 -149.170 46.090 ;
        RECT -149.990 43.680 -149.230 44.030 ;
        RECT -150.380 40.250 -150.030 43.240 ;
        RECT -147.110 42.650 -143.940 43.070 ;
        RECT -142.640 41.680 -142.120 42.200 ;
        RECT -122.320 29.430 -120.240 32.660 ;
        RECT -150.360 16.860 -150.030 18.890 ;
        RECT -149.790 16.800 -149.170 17.500 ;
        RECT -149.990 15.090 -149.230 15.440 ;
        RECT -150.380 11.660 -150.030 14.650 ;
        RECT -147.110 14.060 -143.940 14.480 ;
        RECT -142.640 13.090 -142.120 13.610 ;
        RECT -117.910 0.840 -115.830 4.070 ;
        RECT -150.360 -11.730 -150.030 -9.700 ;
        RECT -149.790 -11.790 -149.170 -11.090 ;
        RECT -149.990 -13.500 -149.230 -13.150 ;
        RECT -150.380 -16.930 -150.030 -13.940 ;
        RECT -147.110 -14.530 -143.940 -14.110 ;
        RECT -142.640 -15.500 -142.120 -14.980 ;
        RECT -113.570 -27.750 -111.490 -24.520 ;
        RECT -150.360 -40.320 -150.030 -38.290 ;
        RECT -149.790 -40.380 -149.170 -39.680 ;
        RECT -149.990 -42.090 -149.230 -41.740 ;
        RECT -150.380 -45.520 -150.030 -42.530 ;
        RECT -147.110 -43.120 -143.940 -42.700 ;
        RECT -142.640 -44.090 -142.120 -43.570 ;
        RECT -150.360 -68.910 -150.030 -66.880 ;
        RECT -149.790 -68.970 -149.170 -68.270 ;
        RECT -149.990 -70.680 -149.230 -70.330 ;
        RECT -150.380 -74.110 -150.030 -71.120 ;
        RECT -147.110 -71.710 -143.940 -71.290 ;
        RECT -142.640 -72.680 -142.120 -72.160 ;
        RECT 212.760 73.260 213.380 73.960 ;
        RECT 213.620 73.320 213.950 75.350 ;
        RECT 212.820 71.550 213.580 71.900 ;
        RECT 207.530 70.520 210.700 70.940 ;
        RECT 205.710 69.550 206.230 70.070 ;
        RECT 213.620 68.120 213.970 71.110 ;
        RECT 188.740 57.300 190.830 60.530 ;
        RECT 212.760 44.670 213.380 45.370 ;
        RECT 213.620 44.730 213.950 46.760 ;
        RECT 212.820 42.960 213.580 43.310 ;
        RECT 207.530 41.930 210.700 42.350 ;
        RECT 205.710 40.960 206.230 41.480 ;
        RECT 213.620 39.530 213.970 42.520 ;
        RECT 184.760 28.710 186.850 31.940 ;
        RECT 212.760 16.080 213.380 16.780 ;
        RECT 213.620 16.140 213.950 18.170 ;
        RECT 212.820 14.370 213.580 14.720 ;
        RECT 207.530 13.340 210.700 13.760 ;
        RECT 205.710 12.370 206.230 12.890 ;
        RECT 213.620 10.940 213.970 13.930 ;
        RECT 180.510 0.120 182.600 3.350 ;
        RECT 212.760 -12.510 213.380 -11.810 ;
        RECT 213.620 -12.450 213.950 -10.420 ;
        RECT 212.820 -14.220 213.580 -13.870 ;
        RECT 207.530 -15.250 210.700 -14.830 ;
        RECT 205.710 -16.220 206.230 -15.700 ;
        RECT 213.620 -17.650 213.970 -14.660 ;
        RECT 176.570 -28.470 178.660 -25.240 ;
        RECT 212.760 -41.100 213.380 -40.400 ;
        RECT 213.620 -41.040 213.950 -39.010 ;
        RECT 212.820 -42.810 213.580 -42.460 ;
        RECT 207.530 -43.840 210.700 -43.420 ;
        RECT 205.710 -44.810 206.230 -44.290 ;
        RECT 213.620 -46.240 213.970 -43.250 ;
        RECT 212.760 -69.690 213.380 -68.990 ;
        RECT 213.620 -69.630 213.950 -67.600 ;
        RECT -105.030 -84.930 -102.950 -81.700 ;
        RECT 108.820 -82.830 113.240 -78.410 ;
        RECT -150.360 -97.500 -150.030 -95.470 ;
        RECT -149.790 -97.560 -149.170 -96.860 ;
        RECT -149.990 -99.270 -149.230 -98.920 ;
        RECT -150.380 -102.700 -150.030 -99.710 ;
        RECT -147.110 -100.300 -143.940 -99.880 ;
        RECT -142.640 -101.270 -142.120 -100.750 ;
        RECT -150.360 -126.090 -150.030 -124.060 ;
        RECT -149.790 -126.150 -149.170 -125.450 ;
        RECT -149.990 -127.860 -149.230 -127.510 ;
        RECT -150.380 -131.290 -150.030 -128.300 ;
        RECT -147.110 -128.890 -143.940 -128.470 ;
        RECT -142.640 -129.860 -142.120 -129.340 ;
        RECT -96.410 -142.110 -94.330 -138.880 ;
        RECT -150.360 -154.680 -150.030 -152.650 ;
        RECT -149.790 -154.740 -149.170 -154.040 ;
        RECT -149.990 -156.450 -149.230 -156.100 ;
        RECT -150.380 -159.880 -150.030 -156.890 ;
        RECT -147.110 -157.480 -143.940 -157.060 ;
        RECT -142.640 -158.450 -142.120 -157.930 ;
        RECT -92.440 -170.700 -90.360 -167.470 ;
        RECT -150.360 -183.270 -150.030 -181.240 ;
        RECT -149.790 -183.330 -149.170 -182.630 ;
        RECT -149.990 -185.040 -149.230 -184.690 ;
        RECT -150.380 -188.470 -150.030 -185.480 ;
        RECT -147.110 -186.070 -143.940 -185.650 ;
        RECT -142.640 -187.040 -142.120 -186.520 ;
        RECT -88.000 -199.290 -85.920 -196.060 ;
        RECT -150.360 -211.860 -150.030 -209.830 ;
        RECT -149.790 -211.920 -149.170 -211.220 ;
        RECT -149.990 -213.630 -149.230 -213.280 ;
        RECT -150.380 -217.060 -150.030 -214.070 ;
        RECT -147.110 -214.660 -143.940 -214.240 ;
        RECT -142.640 -215.630 -142.120 -215.110 ;
        RECT -83.700 -227.880 -81.620 -224.650 ;
        RECT -150.360 -240.450 -150.030 -238.420 ;
        RECT -149.790 -240.510 -149.170 -239.810 ;
      LAYER met2 ;
        RECT -68.920 129.870 -64.830 130.120 ;
        RECT -26.950 129.870 -26.270 129.920 ;
        RECT -68.920 128.700 -26.270 129.870 ;
        RECT 87.770 129.440 88.630 129.480 ;
        RECT 100.280 129.440 105.080 131.530 ;
        RECT -25.720 128.700 -25.270 128.800 ;
        RECT -68.920 128.470 -25.270 128.700 ;
        RECT -68.920 127.620 -26.270 128.470 ;
        RECT -25.720 128.370 -25.270 128.470 ;
        RECT 56.900 128.130 57.360 128.150 ;
        RECT 87.770 128.130 105.130 129.440 ;
        RECT -20.440 127.730 -20.120 127.780 ;
        RECT 56.900 127.760 105.130 128.130 ;
        RECT 56.900 127.740 57.360 127.760 ;
        RECT -68.920 127.020 -64.830 127.620 ;
        RECT -26.950 127.600 -26.270 127.620 ;
        RECT -23.300 127.490 -20.120 127.730 ;
        RECT -23.300 127.470 -22.980 127.490 ;
        RECT 87.770 127.380 105.130 127.760 ;
        RECT -20.750 125.950 -20.430 126.270 ;
        RECT 17.280 126.240 17.730 126.260 ;
        RECT 17.270 126.180 17.750 126.240 ;
        RECT -5.120 126.040 17.750 126.180 ;
        RECT -97.040 125.380 -93.660 125.490 ;
        RECT -26.950 125.380 -26.270 125.390 ;
        RECT -97.450 124.510 -26.270 125.380 ;
        RECT -25.620 124.900 -25.190 125.370 ;
        RECT -20.730 124.910 -20.460 125.950 ;
        RECT -5.140 125.880 17.750 126.040 ;
        RECT -5.140 125.720 -4.820 125.880 ;
        RECT 17.270 125.820 17.750 125.880 ;
        RECT 17.280 125.800 17.730 125.820 ;
        RECT -5.140 125.710 -4.830 125.720 ;
        RECT -23.250 124.900 -20.460 124.910 ;
        RECT -25.620 124.890 -20.460 124.900 ;
        RECT -25.530 124.680 -20.460 124.890 ;
        RECT 87.770 125.310 88.630 125.350 ;
        RECT 129.870 125.310 133.180 127.370 ;
        RECT -25.530 124.670 -20.980 124.680 ;
        RECT 57.730 124.670 58.170 124.690 ;
        RECT 87.770 124.670 133.500 125.310 ;
        RECT -97.450 124.480 -23.290 124.510 ;
        RECT -97.450 124.220 -22.990 124.480 ;
        RECT 57.730 124.300 133.500 124.670 ;
        RECT 57.730 124.280 58.170 124.300 ;
        RECT -97.450 124.190 -23.290 124.220 ;
        RECT -97.450 123.130 -26.270 124.190 ;
        RECT -21.170 124.030 -20.860 124.260 ;
        RECT -24.260 123.930 -20.860 124.030 ;
        RECT -24.260 123.800 -20.880 123.930 ;
        RECT -24.260 123.770 -23.940 123.800 ;
        RECT 87.770 123.250 133.500 124.300 ;
        RECT -97.040 122.810 -93.660 123.130 ;
        RECT -26.950 123.070 -26.270 123.130 ;
        RECT -127.580 120.890 -124.940 122.070 ;
        RECT 85.150 121.490 85.920 121.640 ;
        RECT -24.340 121.070 85.920 121.490 ;
        RECT 85.150 120.930 85.920 121.070 ;
        RECT 87.740 121.230 88.600 121.260 ;
        RECT 158.260 121.230 162.190 121.680 ;
        RECT -27.400 120.890 -26.720 120.920 ;
        RECT -127.660 120.250 -26.720 120.890 ;
        RECT -18.480 120.250 -18.010 120.270 ;
        RECT -127.660 119.670 -18.010 120.250 ;
        RECT -127.660 119.430 -26.680 119.670 ;
        RECT -18.480 119.650 -18.010 119.670 ;
        RECT 58.510 119.960 58.930 119.980 ;
        RECT 87.740 119.960 162.190 121.230 ;
        RECT 58.510 119.590 162.190 119.960 ;
        RECT 58.510 119.570 58.930 119.590 ;
        RECT -127.660 118.640 -26.720 119.430 ;
        RECT 87.740 119.170 162.190 119.590 ;
        RECT 87.740 119.160 88.600 119.170 ;
        RECT 158.260 119.160 162.190 119.170 ;
        RECT 4.690 118.980 5.000 119.000 ;
        RECT -139.810 116.550 -136.920 118.510 ;
        RECT -127.580 118.470 -124.940 118.640 ;
        RECT -27.400 118.600 -26.720 118.640 ;
        RECT -5.100 118.900 -4.780 118.910 ;
        RECT 4.690 118.900 5.010 118.980 ;
        RECT 28.870 118.910 29.190 118.930 ;
        RECT 28.870 118.900 29.200 118.910 ;
        RECT 35.640 118.900 35.960 118.930 ;
        RECT 50.410 118.900 50.730 118.920 ;
        RECT 65.070 118.900 65.630 119.040 ;
        RECT -5.100 118.670 65.630 118.900 ;
        RECT -5.100 118.590 -4.780 118.670 ;
        RECT 4.690 118.660 5.000 118.670 ;
        RECT 28.870 118.650 29.200 118.670 ;
        RECT 35.640 118.650 35.960 118.670 ;
        RECT 50.410 118.660 50.730 118.670 ;
        RECT 65.070 118.530 65.630 118.670 ;
        RECT 0.690 118.450 1.060 118.510 ;
        RECT 63.890 118.450 64.430 118.470 ;
        RECT 0.690 118.220 64.430 118.450 ;
        RECT 0.690 118.160 1.060 118.220 ;
        RECT 32.490 118.000 32.770 118.010 ;
        RECT 3.520 117.990 3.830 118.000 ;
        RECT 32.470 117.990 32.790 118.000 ;
        RECT 35.200 117.990 35.520 118.020 ;
        RECT 49.520 117.990 49.840 118.050 ;
        RECT 62.810 117.990 63.350 118.000 ;
        RECT 3.520 117.760 63.350 117.990 ;
        RECT 63.890 117.910 64.430 118.220 ;
        RECT 3.520 117.730 3.850 117.760 ;
        RECT 32.470 117.740 32.790 117.760 ;
        RECT 35.200 117.740 35.520 117.760 ;
        RECT 32.490 117.730 32.770 117.740 ;
        RECT 3.520 117.710 3.830 117.730 ;
        RECT -2.560 117.530 -2.240 117.540 ;
        RECT 61.870 117.530 62.400 117.560 ;
        RECT -2.560 117.300 62.400 117.530 ;
        RECT 62.810 117.440 63.350 117.760 ;
        RECT -2.560 117.240 -2.240 117.300 ;
        RECT 29.340 116.950 29.660 116.990 ;
        RECT 44.990 116.950 46.270 117.050 ;
        RECT 61.870 116.950 62.400 117.300 ;
        RECT 29.340 116.740 46.270 116.950 ;
        RECT 187.060 116.890 190.560 117.430 ;
        RECT 29.340 116.710 29.660 116.740 ;
        RECT -27.720 116.550 -26.450 116.560 ;
        RECT -139.840 115.100 -26.450 116.550 ;
        RECT 13.240 115.730 13.500 116.530 ;
        RECT 16.940 116.510 17.260 116.520 ;
        RECT 16.930 116.500 17.260 116.510 ;
        RECT 17.970 116.500 18.290 116.550 ;
        RECT 16.930 116.300 22.250 116.500 ;
        RECT 41.760 116.370 42.040 116.390 ;
        RECT 16.930 116.250 17.260 116.300 ;
        RECT 17.970 116.290 18.290 116.300 ;
        RECT 16.940 116.230 17.260 116.250 ;
        RECT 22.050 115.800 22.250 116.300 ;
        RECT 41.740 116.340 42.060 116.370 ;
        RECT 73.880 116.340 75.220 116.880 ;
        RECT 88.580 116.870 190.650 116.890 ;
        RECT 41.740 116.130 75.220 116.340 ;
        RECT 41.740 116.110 42.060 116.130 ;
        RECT 41.760 116.090 42.040 116.110 ;
        RECT 48.070 115.800 48.380 115.860 ;
        RECT 15.240 115.730 15.580 115.790 ;
        RECT 13.140 115.510 15.580 115.730 ;
        RECT 22.050 115.600 48.380 115.800 ;
        RECT 73.880 115.600 75.220 116.130 ;
        RECT 48.070 115.540 48.380 115.600 ;
        RECT 27.000 115.330 27.320 115.380 ;
        RECT 22.000 115.130 27.370 115.330 ;
        RECT -16.370 115.100 -16.070 115.110 ;
        RECT -6.780 115.100 -6.490 115.120 ;
        RECT -139.840 114.710 -6.460 115.100 ;
        RECT -139.840 114.690 -26.450 114.710 ;
        RECT -6.780 114.690 -6.490 114.710 ;
        RECT -27.720 114.680 -26.450 114.690 ;
        RECT -7.420 114.290 -7.130 114.310 ;
        RECT -19.870 113.890 -7.110 114.290 ;
        RECT 13.240 113.980 13.500 114.780 ;
        RECT 16.940 114.760 17.260 114.770 ;
        RECT 16.930 114.750 17.260 114.760 ;
        RECT 17.970 114.750 18.290 114.800 ;
        RECT 22.000 114.750 22.200 115.130 ;
        RECT 27.000 115.120 27.320 115.130 ;
        RECT 29.760 114.890 30.070 114.900 ;
        RECT 59.390 114.890 59.820 114.910 ;
        RECT 87.740 114.890 190.650 116.870 ;
        RECT 29.760 114.860 30.080 114.890 ;
        RECT 16.930 114.550 22.200 114.750 ;
        RECT 22.510 114.660 30.080 114.860 ;
        RECT 16.930 114.500 17.260 114.550 ;
        RECT 17.970 114.540 18.290 114.550 ;
        RECT 16.940 114.480 17.260 114.500 ;
        RECT 15.240 113.980 15.580 114.040 ;
        RECT -130.950 112.070 -27.430 112.110 ;
        RECT -130.950 111.200 -26.160 112.070 ;
        RECT -19.870 111.200 -19.470 113.890 ;
        RECT -7.420 113.880 -7.130 113.890 ;
        RECT 13.140 113.760 15.580 113.980 ;
        RECT -16.070 113.210 -15.700 113.220 ;
        RECT -17.860 112.980 -15.700 113.210 ;
        RECT -10.020 113.080 -9.710 113.170 ;
        RECT -10.610 112.980 -9.710 113.080 ;
        RECT -17.860 112.910 -9.710 112.980 ;
        RECT -17.860 112.850 -10.440 112.910 ;
        RECT -17.860 112.150 -17.240 112.850 ;
        RECT -16.070 112.810 -10.440 112.850 ;
        RECT -10.020 112.840 -9.710 112.910 ;
        RECT -8.930 113.090 -8.620 113.180 ;
        RECT -8.930 112.990 -8.470 113.090 ;
        RECT -7.410 112.990 -7.090 113.040 ;
        RECT -8.930 112.850 -7.030 112.990 ;
        RECT -8.630 112.820 -7.030 112.850 ;
        RECT -7.410 112.780 -7.090 112.820 ;
        RECT -11.180 112.570 -10.860 112.620 ;
        RECT -10.450 112.570 -10.140 112.670 ;
        RECT -11.180 112.400 -10.140 112.570 ;
        RECT -11.180 112.360 -10.860 112.400 ;
        RECT -10.450 112.340 -10.140 112.400 ;
        RECT 13.240 112.230 13.500 113.030 ;
        RECT 16.940 113.010 17.260 113.020 ;
        RECT 16.930 113.000 17.260 113.010 ;
        RECT 17.970 113.000 18.290 113.050 ;
        RECT 22.510 113.000 22.710 114.660 ;
        RECT 29.760 114.630 30.080 114.660 ;
        RECT 59.390 114.840 190.650 114.890 ;
        RECT 59.390 114.770 88.600 114.840 ;
        RECT 29.760 114.620 30.070 114.630 ;
        RECT 59.390 114.520 88.490 114.770 ;
        RECT 59.390 114.490 59.800 114.520 ;
        RECT 30.820 114.380 31.140 114.420 ;
        RECT 16.930 112.800 22.710 113.000 ;
        RECT 23.060 114.180 31.220 114.380 ;
        RECT 16.930 112.750 17.260 112.800 ;
        RECT 17.970 112.790 18.290 112.800 ;
        RECT 16.940 112.730 17.260 112.750 ;
        RECT 15.240 112.230 15.580 112.290 ;
        RECT -16.070 112.150 -15.700 112.190 ;
        RECT -130.950 110.800 -19.470 111.200 ;
        RECT -18.390 112.060 -15.700 112.150 ;
        RECT -10.010 112.090 -9.700 112.180 ;
        RECT -10.540 112.060 -9.700 112.090 ;
        RECT -18.390 111.920 -9.700 112.060 ;
        RECT -18.390 111.890 -10.440 111.920 ;
        RECT -18.390 111.780 -15.700 111.890 ;
        RECT -10.010 111.850 -9.700 111.920 ;
        RECT -8.920 112.100 -8.610 112.190 ;
        RECT -8.920 112.070 -8.460 112.100 ;
        RECT -7.410 112.070 -7.090 112.120 ;
        RECT -8.920 111.900 -7.030 112.070 ;
        RECT 13.140 112.010 15.580 112.230 ;
        RECT -8.920 111.860 -8.610 111.900 ;
        RECT -7.410 111.860 -7.090 111.900 ;
        RECT -18.390 111.670 -17.240 111.780 ;
        RECT -18.390 111.220 -17.280 111.670 ;
        RECT -11.210 111.650 -10.890 111.700 ;
        RECT -10.470 111.650 -10.160 111.750 ;
        RECT -11.210 111.480 -10.160 111.650 ;
        RECT -11.210 111.440 -10.890 111.480 ;
        RECT -10.470 111.420 -10.160 111.480 ;
        RECT -16.070 111.220 -15.700 111.260 ;
        RECT -18.390 111.140 -15.700 111.220 ;
        RECT -18.390 111.110 -10.440 111.140 ;
        RECT -18.390 111.100 -10.400 111.110 ;
        RECT -10.010 111.100 -9.700 111.190 ;
        RECT -18.390 110.970 -9.700 111.100 ;
        RECT -18.390 110.850 -15.700 110.970 ;
        RECT -10.540 110.930 -9.700 110.970 ;
        RECT -10.010 110.860 -9.700 110.930 ;
        RECT -8.920 111.150 -8.610 111.200 ;
        RECT -7.440 111.150 -7.120 111.200 ;
        RECT -8.920 110.980 -7.030 111.150 ;
        RECT -8.920 110.940 -8.460 110.980 ;
        RECT -7.440 110.940 -7.120 110.980 ;
        RECT -8.920 110.870 -8.610 110.940 ;
        RECT -18.390 110.810 -17.490 110.850 ;
        RECT -130.950 110.190 -26.160 110.800 ;
        RECT -130.950 110.030 -27.430 110.190 ;
        RECT -130.950 89.920 -128.870 110.030 ;
        RECT -126.790 107.140 -26.950 107.230 ;
        RECT -126.790 106.260 -25.730 107.140 ;
        RECT -18.390 106.260 -18.020 110.810 ;
        RECT -11.200 110.730 -10.880 110.780 ;
        RECT -10.490 110.730 -10.180 110.760 ;
        RECT -11.200 110.560 -10.180 110.730 ;
        RECT -11.200 110.520 -10.880 110.560 ;
        RECT -10.490 110.430 -10.180 110.560 ;
        RECT 13.240 110.480 13.500 111.280 ;
        RECT 16.940 111.260 17.260 111.270 ;
        RECT 16.930 111.250 17.260 111.260 ;
        RECT 17.970 111.250 18.290 111.300 ;
        RECT 23.060 111.250 23.260 114.180 ;
        RECT 30.820 114.140 31.140 114.180 ;
        RECT 49.460 113.580 50.040 114.020 ;
        RECT 49.460 113.390 50.100 113.580 ;
        RECT 49.860 113.030 50.100 113.390 ;
        RECT 50.480 113.380 51.060 114.010 ;
        RECT 50.500 113.030 50.810 113.040 ;
        RECT 49.860 112.780 50.810 113.030 ;
        RECT 198.760 112.820 204.470 118.460 ;
        RECT 50.500 112.710 50.810 112.780 ;
        RECT 51.470 112.710 51.780 112.790 ;
        RECT 53.720 112.710 54.030 112.810 ;
        RECT 198.320 112.780 204.470 112.820 ;
        RECT 88.580 112.770 204.470 112.780 ;
        RECT 88.230 112.760 204.470 112.770 ;
        RECT 28.700 112.560 29.020 112.570 ;
        RECT 16.930 111.050 23.260 111.250 ;
        RECT 26.210 112.550 26.500 112.560 ;
        RECT 28.460 112.550 29.020 112.560 ;
        RECT 46.780 112.550 47.090 112.560 ;
        RECT 26.210 112.370 49.260 112.550 ;
        RECT 51.470 112.480 54.030 112.710 ;
        RECT 74.380 112.580 74.680 112.600 ;
        RECT 87.670 112.580 204.470 112.760 ;
        RECT 51.470 112.460 51.780 112.480 ;
        RECT 16.930 111.000 17.260 111.050 ;
        RECT 17.970 111.040 18.290 111.050 ;
        RECT 16.940 110.980 17.260 111.000 ;
        RECT 15.240 110.480 15.580 110.540 ;
        RECT 13.140 110.260 15.580 110.480 ;
        RECT -10.200 110.150 -9.890 110.260 ;
        RECT -10.540 110.140 -9.890 110.150 ;
        RECT -16.910 110.120 -9.890 110.140 ;
        RECT -126.790 105.890 -18.020 106.260 ;
        RECT -17.200 109.960 -9.890 110.120 ;
        RECT -17.200 109.950 -10.420 109.960 ;
        RECT -17.200 109.770 -15.700 109.950 ;
        RECT -10.200 109.930 -9.890 109.960 ;
        RECT -8.900 110.080 -8.590 110.160 ;
        RECT -6.800 110.080 -6.480 110.110 ;
        RECT -8.900 109.880 -6.380 110.080 ;
        RECT -8.900 109.830 -8.590 109.880 ;
        RECT -6.800 109.850 -6.480 109.880 ;
        RECT -17.200 109.180 -16.540 109.770 ;
        RECT -16.070 109.730 -15.700 109.770 ;
        RECT -11.850 109.720 -11.530 109.760 ;
        RECT -10.230 109.730 -9.910 109.790 ;
        RECT -10.540 109.720 -9.910 109.730 ;
        RECT -11.850 109.540 -9.910 109.720 ;
        RECT -11.850 109.530 -10.420 109.540 ;
        RECT -11.850 109.500 -11.530 109.530 ;
        RECT -10.230 109.470 -9.910 109.540 ;
        RECT 21.130 109.540 21.450 109.590 ;
        RECT 23.540 109.540 23.860 109.560 ;
        RECT 26.210 109.540 26.390 112.370 ;
        RECT 28.460 112.230 28.770 112.370 ;
        RECT 46.780 112.230 47.090 112.370 ;
        RECT 74.370 112.320 204.470 112.580 ;
        RECT 50.650 112.170 50.960 112.210 ;
        RECT 50.470 112.060 51.190 112.170 ;
        RECT 74.370 112.160 204.310 112.320 ;
        RECT 74.380 112.140 74.680 112.160 ;
        RECT 51.420 112.060 51.730 112.140 ;
        RECT 50.470 111.920 51.730 112.060 ;
        RECT 50.650 111.880 51.730 111.920 ;
        RECT 50.920 111.850 51.730 111.880 ;
        RECT 50.920 111.810 51.190 111.850 ;
        RECT 51.420 111.810 51.730 111.850 ;
        RECT 87.670 111.820 204.310 112.160 ;
        RECT 46.930 111.530 47.240 111.600 ;
        RECT 49.530 111.530 49.840 111.670 ;
        RECT 46.930 111.340 49.840 111.530 ;
        RECT 46.930 111.310 49.530 111.340 ;
        RECT 46.930 111.270 47.240 111.310 ;
        RECT 50.990 111.240 51.190 111.250 ;
        RECT 51.420 111.240 51.730 111.280 ;
        RECT 50.990 111.160 51.730 111.240 ;
        RECT 50.700 111.140 51.730 111.160 ;
        RECT 50.650 111.030 51.730 111.140 ;
        RECT 28.070 111.010 28.380 111.030 ;
        RECT 37.800 111.010 45.790 111.020 ;
        RECT 28.070 110.820 45.790 111.010 ;
        RECT 50.650 110.900 51.210 111.030 ;
        RECT 51.420 110.950 51.730 111.030 ;
        RECT 50.650 110.890 51.120 110.900 ;
        RECT 28.070 110.700 28.380 110.820 ;
        RECT 27.350 110.130 27.670 110.160 ;
        RECT 44.390 110.140 44.610 110.150 ;
        RECT 37.810 110.130 44.640 110.140 ;
        RECT 27.350 109.900 44.640 110.130 ;
        RECT 45.570 110.100 45.790 110.820 ;
        RECT 51.470 110.570 51.780 110.630 ;
        RECT 53.770 110.570 54.080 110.590 ;
        RECT 50.560 110.390 51.160 110.510 ;
        RECT 50.260 110.350 51.160 110.390 ;
        RECT 49.940 110.110 51.160 110.350 ;
        RECT 51.470 110.340 59.390 110.570 ;
        RECT 59.760 110.340 68.910 110.570 ;
        RECT 87.730 110.420 204.310 111.820 ;
        RECT 87.730 110.390 88.630 110.420 ;
        RECT 51.470 110.300 51.780 110.340 ;
        RECT 53.770 110.260 54.080 110.340 ;
        RECT 37.810 109.890 44.640 109.900 ;
        RECT 13.140 109.290 15.580 109.510 ;
        RECT -17.200 109.160 -10.420 109.180 ;
        RECT -10.200 109.160 -9.890 109.270 ;
        RECT -17.200 108.990 -9.890 109.160 ;
        RECT -17.200 108.810 -15.700 108.990 ;
        RECT -10.540 108.970 -9.890 108.990 ;
        RECT -10.200 108.940 -9.890 108.970 ;
        RECT -8.900 109.120 -8.590 109.170 ;
        RECT -6.790 109.120 -6.470 109.150 ;
        RECT -8.900 108.920 -6.380 109.120 ;
        RECT -8.900 108.840 -8.590 108.920 ;
        RECT -6.790 108.890 -6.470 108.920 ;
        RECT -17.200 108.800 -16.530 108.810 ;
        RECT -17.200 108.760 -16.540 108.800 ;
        RECT -16.070 108.770 -15.700 108.810 ;
        RECT -11.890 108.760 -11.570 108.800 ;
        RECT -126.790 105.260 -25.730 105.890 ;
        RECT -126.790 105.150 -26.950 105.260 ;
        RECT -131.020 86.550 -128.680 89.920 ;
        RECT -130.950 85.680 -128.870 86.550 ;
        RECT -126.790 61.320 -124.710 105.150 ;
        RECT -127.010 57.910 -124.710 61.320 ;
        RECT -126.790 57.580 -124.710 57.910 ;
        RECT -122.450 102.390 -26.950 102.410 ;
        RECT -122.450 101.500 -25.790 102.390 ;
        RECT -17.200 101.500 -16.830 108.760 ;
        RECT -11.890 108.740 -10.420 108.760 ;
        RECT -10.230 108.740 -9.910 108.800 ;
        RECT -11.890 108.570 -9.910 108.740 ;
        RECT -11.890 108.540 -11.570 108.570 ;
        RECT -10.540 108.550 -9.910 108.570 ;
        RECT -10.230 108.480 -9.910 108.550 ;
        RECT 13.240 108.490 13.500 109.290 ;
        RECT 15.240 109.230 15.580 109.290 ;
        RECT 21.130 109.370 26.390 109.540 ;
        RECT 21.130 109.350 23.860 109.370 ;
        RECT 21.130 109.270 21.450 109.350 ;
        RECT 23.540 109.300 23.860 109.350 ;
        RECT 28.060 109.150 28.370 109.340 ;
        RECT 37.810 109.150 41.320 109.160 ;
        RECT 16.940 108.770 17.260 108.790 ;
        RECT 16.930 108.720 17.260 108.770 ;
        RECT 19.780 108.760 20.370 109.060 ;
        RECT 28.060 109.010 41.320 109.150 ;
        RECT 28.090 108.970 41.320 109.010 ;
        RECT 28.090 108.960 37.810 108.970 ;
        RECT 19.780 108.740 20.130 108.760 ;
        RECT 17.970 108.720 18.290 108.730 ;
        RECT 19.780 108.720 19.980 108.740 ;
        RECT 16.930 108.520 19.980 108.720 ;
        RECT 16.930 108.510 17.260 108.520 ;
        RECT 16.940 108.500 17.260 108.510 ;
        RECT 17.970 108.470 18.290 108.520 ;
        RECT 41.090 108.370 41.320 108.970 ;
        RECT 44.350 108.720 44.640 109.890 ;
        RECT 45.540 110.060 45.790 110.100 ;
        RECT 50.260 110.060 51.160 110.110 ;
        RECT 45.540 109.420 45.800 110.060 ;
        RECT 50.560 109.950 51.160 110.060 ;
        RECT 68.620 110.240 68.910 110.340 ;
        RECT 78.410 110.320 79.530 110.330 ;
        RECT 76.600 110.240 81.060 110.320 ;
        RECT 68.620 110.120 81.060 110.240 ;
        RECT 68.620 110.040 76.950 110.120 ;
        RECT 78.410 110.110 79.530 110.120 ;
        RECT 68.620 110.030 68.910 110.040 ;
        RECT 79.180 109.990 79.490 110.110 ;
        RECT 80.750 109.990 81.060 110.120 ;
        RECT 51.470 109.740 51.780 109.790 ;
        RECT 53.760 109.740 54.070 109.870 ;
        RECT 51.470 109.520 59.390 109.740 ;
        RECT 59.760 109.520 67.970 109.740 ;
        RECT 51.470 109.460 51.780 109.520 ;
        RECT 45.540 109.210 49.670 109.420 ;
        RECT 49.460 109.070 49.670 109.210 ;
        RECT 51.420 109.070 51.730 109.140 ;
        RECT 49.460 108.860 51.730 109.070 ;
        RECT 51.120 108.850 51.730 108.860 ;
        RECT 46.930 108.770 47.240 108.840 ;
        RECT 51.420 108.810 51.730 108.850 ;
        RECT 46.930 108.720 49.260 108.770 ;
        RECT 44.350 108.560 49.260 108.720 ;
        RECT 44.350 108.500 47.240 108.560 ;
        RECT 44.350 108.490 44.640 108.500 ;
        RECT -122.450 101.130 -16.830 101.500 ;
        RECT -16.070 108.170 -10.420 108.220 ;
        RECT -10.200 108.170 -9.890 108.280 ;
        RECT 41.090 108.220 41.310 108.370 ;
        RECT 51.420 108.270 51.730 108.280 ;
        RECT 45.460 108.220 51.730 108.270 ;
        RECT -16.070 108.030 -9.890 108.170 ;
        RECT -122.450 100.510 -25.790 101.130 ;
        RECT -122.450 100.330 -26.950 100.510 ;
        RECT -122.450 32.840 -120.370 100.330 ;
        RECT -117.910 97.570 -26.950 97.710 ;
        RECT -117.910 96.660 -25.730 97.570 ;
        RECT -16.070 96.660 -15.700 108.030 ;
        RECT -10.540 107.980 -9.890 108.030 ;
        RECT -10.200 107.950 -9.890 107.980 ;
        RECT -8.900 108.160 -8.590 108.180 ;
        RECT -6.800 108.160 -6.480 108.190 ;
        RECT -8.900 107.960 -6.380 108.160 ;
        RECT 41.090 108.060 51.730 108.220 ;
        RECT 41.090 108.000 45.850 108.060 ;
        RECT 51.120 108.030 51.730 108.060 ;
        RECT -8.900 107.850 -8.590 107.960 ;
        RECT -6.800 107.930 -6.480 107.960 ;
        RECT 51.420 107.950 51.730 108.030 ;
        RECT -11.850 107.800 -11.530 107.840 ;
        RECT -11.850 107.750 -10.420 107.800 ;
        RECT -10.230 107.750 -9.910 107.810 ;
        RECT -11.850 107.610 -9.910 107.750 ;
        RECT -11.850 107.580 -11.530 107.610 ;
        RECT -10.540 107.560 -9.910 107.610 ;
        RECT -10.230 107.490 -9.910 107.560 ;
        RECT 13.140 107.540 15.580 107.760 ;
        RECT 20.030 107.720 20.370 107.790 ;
        RECT 13.240 106.740 13.500 107.540 ;
        RECT 15.240 107.480 15.580 107.540 ;
        RECT 19.730 107.490 20.370 107.720 ;
        RECT 28.460 107.680 28.770 107.820 ;
        RECT 26.290 107.670 28.770 107.680 ;
        RECT 46.780 107.680 47.090 107.820 ;
        RECT 46.780 107.670 49.260 107.680 ;
        RECT 25.770 107.520 49.260 107.670 ;
        RECT 67.750 107.640 67.970 109.520 ;
        RECT 80.100 109.340 80.420 109.380 ;
        RECT 81.110 109.340 81.430 109.370 ;
        RECT 80.050 109.140 83.820 109.340 ;
        RECT 80.100 109.120 80.420 109.140 ;
        RECT 81.110 109.110 81.430 109.140 ;
        RECT 82.100 109.060 83.810 109.140 ;
        RECT 80.100 108.610 80.420 108.630 ;
        RECT 81.110 108.610 81.430 108.640 ;
        RECT 83.610 108.610 83.810 109.060 ;
        RECT 80.050 108.410 83.810 108.610 ;
        RECT 80.100 108.370 80.420 108.410 ;
        RECT 81.110 108.380 81.430 108.410 ;
        RECT 79.180 107.640 79.490 107.760 ;
        RECT 67.750 107.630 69.350 107.640 ;
        RECT 78.410 107.630 79.530 107.640 ;
        RECT 80.750 107.630 81.060 107.760 ;
        RECT 25.770 107.500 28.770 107.520 ;
        RECT 25.770 107.490 26.500 107.500 ;
        RECT 28.460 107.490 28.770 107.500 ;
        RECT 46.780 107.500 49.260 107.520 ;
        RECT 51.470 107.580 51.780 107.630 ;
        RECT 53.680 107.580 53.990 107.620 ;
        RECT 46.780 107.490 47.090 107.500 ;
        RECT 16.940 107.020 17.260 107.040 ;
        RECT 16.930 106.970 17.260 107.020 ;
        RECT 17.970 106.970 18.290 106.980 ;
        RECT 19.730 106.970 19.930 107.490 ;
        RECT 25.770 107.280 25.950 107.490 ;
        RECT 51.470 107.350 54.180 107.580 ;
        RECT 67.750 107.430 81.060 107.630 ;
        RECT 67.750 107.420 69.350 107.430 ;
        RECT 78.410 107.420 79.530 107.430 ;
        RECT 83.610 107.360 83.810 108.410 ;
        RECT 192.980 108.040 195.070 108.220 ;
        RECT 88.580 108.030 195.070 108.040 ;
        RECT 87.700 107.360 195.070 108.030 ;
        RECT 32.470 107.330 32.780 107.340 ;
        RECT 16.930 106.770 19.930 106.970 ;
        RECT 21.130 107.200 21.450 107.280 ;
        RECT 23.610 107.250 25.950 107.280 ;
        RECT 32.460 107.270 32.790 107.330 ;
        RECT 51.470 107.300 51.780 107.350 ;
        RECT 53.680 107.290 53.990 107.350 ;
        RECT 23.540 107.200 25.950 107.250 ;
        RECT 32.110 107.220 32.790 107.270 ;
        RECT 21.130 107.120 25.950 107.200 ;
        RECT 21.130 107.010 23.860 107.120 ;
        RECT 24.340 107.110 25.950 107.120 ;
        RECT 25.040 107.100 25.950 107.110 ;
        RECT 21.130 106.960 21.450 107.010 ;
        RECT 23.540 106.990 23.860 107.010 ;
        RECT 28.880 107.050 32.790 107.220 ;
        RECT 54.940 107.060 59.390 107.220 ;
        RECT 28.880 107.000 32.780 107.050 ;
        RECT 54.910 107.020 59.390 107.060 ;
        RECT 59.760 107.120 76.950 107.220 ;
        RECT 78.410 107.120 79.530 107.130 ;
        RECT 59.760 107.020 81.060 107.120 ;
        RECT 49.500 107.000 50.060 107.020 ;
        RECT 50.500 107.000 50.810 107.010 ;
        RECT 16.930 106.760 17.260 106.770 ;
        RECT 16.940 106.750 17.260 106.760 ;
        RECT 17.970 106.720 18.290 106.770 ;
        RECT 49.500 106.750 50.810 107.000 ;
        RECT 28.470 106.520 28.780 106.530 ;
        RECT 46.780 106.520 47.090 106.530 ;
        RECT 21.130 106.340 21.450 106.390 ;
        RECT 23.540 106.340 23.860 106.360 ;
        RECT 21.130 106.320 23.860 106.340 ;
        RECT 25.870 106.340 49.260 106.520 ;
        RECT 49.500 106.480 50.060 106.750 ;
        RECT 50.500 106.680 50.810 106.750 ;
        RECT 51.470 106.680 51.780 106.760 ;
        RECT 53.720 106.680 54.030 106.780 ;
        RECT 51.470 106.450 54.030 106.680 ;
        RECT 51.470 106.430 51.780 106.450 ;
        RECT 25.870 106.320 26.050 106.340 ;
        RECT 21.130 106.160 26.050 106.320 ;
        RECT 28.470 106.200 28.780 106.340 ;
        RECT 46.780 106.200 47.090 106.340 ;
        RECT 21.130 106.150 23.860 106.160 ;
        RECT 21.130 106.070 21.450 106.150 ;
        RECT 23.540 106.100 23.860 106.150 ;
        RECT 50.650 106.140 50.960 106.180 ;
        RECT 50.470 106.030 51.190 106.140 ;
        RECT 51.420 106.030 51.730 106.110 ;
        RECT 13.140 105.790 15.580 106.010 ;
        RECT 35.580 105.940 35.890 105.980 ;
        RECT 35.200 105.920 36.040 105.940 ;
        RECT 19.890 105.850 20.370 105.860 ;
        RECT 13.240 104.990 13.500 105.790 ;
        RECT 15.240 105.730 15.580 105.790 ;
        RECT 19.760 105.560 20.370 105.850 ;
        RECT 35.200 105.740 37.830 105.920 ;
        RECT 50.470 105.890 51.730 106.030 ;
        RECT 50.650 105.850 51.730 105.890 ;
        RECT 50.920 105.820 51.730 105.850 ;
        RECT 50.920 105.780 51.190 105.820 ;
        RECT 51.420 105.780 51.730 105.820 ;
        RECT 35.580 105.650 35.890 105.740 ;
        RECT 19.760 105.410 20.080 105.560 ;
        RECT 28.320 105.500 28.630 105.570 ;
        RECT 26.300 105.490 28.630 105.500 ;
        RECT 46.930 105.500 47.240 105.570 ;
        RECT 49.530 105.500 49.840 105.640 ;
        RECT 16.940 105.270 17.260 105.290 ;
        RECT 16.930 105.220 17.260 105.270 ;
        RECT 17.970 105.220 18.290 105.230 ;
        RECT 19.760 105.220 19.960 105.410 ;
        RECT 26.300 105.280 45.790 105.490 ;
        RECT 27.610 105.270 45.790 105.280 ;
        RECT 28.320 105.240 28.630 105.270 ;
        RECT 16.930 105.020 19.960 105.220 ;
        RECT 16.930 105.010 17.260 105.020 ;
        RECT 16.940 105.000 17.260 105.010 ;
        RECT 17.970 104.970 18.290 105.020 ;
        RECT 20.030 104.520 20.370 104.590 ;
        RECT 19.890 104.470 20.370 104.520 ;
        RECT 19.690 104.290 20.370 104.470 ;
        RECT 27.370 104.300 44.610 104.520 ;
        RECT 13.140 104.040 15.580 104.260 ;
        RECT 13.240 103.240 13.500 104.040 ;
        RECT 15.240 103.980 15.580 104.040 ;
        RECT 16.940 103.520 17.260 103.540 ;
        RECT 16.930 103.470 17.260 103.520 ;
        RECT 17.970 103.470 18.290 103.480 ;
        RECT 19.690 103.470 19.870 104.290 ;
        RECT 27.370 104.160 27.690 104.300 ;
        RECT 21.130 104.000 21.450 104.080 ;
        RECT 23.540 104.020 23.860 104.050 ;
        RECT 23.540 104.000 26.150 104.020 ;
        RECT 21.130 103.840 26.150 104.000 ;
        RECT 21.130 103.810 23.860 103.840 ;
        RECT 21.130 103.760 21.450 103.810 ;
        RECT 23.540 103.790 23.860 103.810 ;
        RECT 16.930 103.270 19.880 103.470 ;
        RECT 16.930 103.260 17.260 103.270 ;
        RECT 16.940 103.250 17.260 103.260 ;
        RECT 17.970 103.220 18.290 103.270 ;
        RECT 25.970 101.650 26.150 103.840 ;
        RECT 27.390 103.820 27.650 104.160 ;
        RECT 27.370 103.560 27.690 103.820 ;
        RECT 28.320 102.740 28.630 102.810 ;
        RECT 26.300 102.530 41.310 102.740 ;
        RECT 27.610 102.520 41.310 102.530 ;
        RECT 28.320 102.480 28.630 102.520 ;
        RECT 35.610 102.230 35.920 102.290 ;
        RECT 35.150 102.220 35.920 102.230 ;
        RECT 35.150 102.210 36.040 102.220 ;
        RECT 35.150 102.000 37.830 102.210 ;
        RECT 41.090 102.190 41.310 102.520 ;
        RECT 44.390 102.690 44.610 104.300 ;
        RECT 45.570 104.070 45.790 105.270 ;
        RECT 46.930 105.310 49.840 105.500 ;
        RECT 46.930 105.280 49.530 105.310 ;
        RECT 46.930 105.240 47.240 105.280 ;
        RECT 50.990 105.210 51.190 105.220 ;
        RECT 51.420 105.210 51.730 105.250 ;
        RECT 50.990 105.130 51.730 105.210 ;
        RECT 50.700 105.110 51.730 105.130 ;
        RECT 50.650 105.000 51.730 105.110 ;
        RECT 50.650 104.870 51.210 105.000 ;
        RECT 51.420 104.920 51.730 105.000 ;
        RECT 50.650 104.860 51.120 104.870 ;
        RECT 51.470 104.540 51.780 104.600 ;
        RECT 53.770 104.540 54.080 104.560 ;
        RECT 54.910 104.540 55.140 107.020 ;
        RECT 76.650 106.920 81.060 107.020 ;
        RECT 78.410 106.910 79.530 106.920 ;
        RECT 79.180 106.790 79.490 106.910 ;
        RECT 80.750 106.790 81.060 106.920 ;
        RECT 83.610 106.930 195.070 107.360 ;
        RECT 83.610 106.240 83.810 106.930 ;
        RECT 80.100 106.140 80.420 106.180 ;
        RECT 81.110 106.140 81.430 106.170 ;
        RECT 82.100 106.140 83.810 106.240 ;
        RECT 80.050 105.940 83.810 106.140 ;
        RECT 87.700 105.950 195.070 106.930 ;
        RECT 87.700 105.940 88.600 105.950 ;
        RECT 80.100 105.920 80.420 105.940 ;
        RECT 81.110 105.910 81.430 105.940 ;
        RECT 83.610 105.590 83.810 105.940 ;
        RECT 80.100 105.410 80.420 105.430 ;
        RECT 81.110 105.410 81.430 105.440 ;
        RECT 82.100 105.410 83.810 105.590 ;
        RECT 80.050 105.270 83.810 105.410 ;
        RECT 80.050 105.210 83.800 105.270 ;
        RECT 80.100 105.170 80.420 105.210 ;
        RECT 81.110 105.180 81.430 105.210 ;
        RECT 50.540 104.360 51.160 104.460 ;
        RECT 50.260 104.320 51.160 104.360 ;
        RECT 49.940 104.080 51.160 104.320 ;
        RECT 51.470 104.310 55.140 104.540 ;
        RECT 55.750 104.410 59.390 104.610 ;
        RECT 59.760 104.430 76.950 104.610 ;
        RECT 79.180 104.440 79.490 104.560 ;
        RECT 78.410 104.430 79.530 104.440 ;
        RECT 80.750 104.430 81.060 104.560 ;
        RECT 59.760 104.410 81.060 104.430 ;
        RECT 51.470 104.270 51.780 104.310 ;
        RECT 53.770 104.230 54.080 104.310 ;
        RECT 45.540 104.030 45.790 104.070 ;
        RECT 50.260 104.030 51.160 104.080 ;
        RECT 45.540 103.390 45.800 104.030 ;
        RECT 50.540 103.930 51.160 104.030 ;
        RECT 51.470 103.710 51.780 103.760 ;
        RECT 53.760 103.710 54.070 103.840 ;
        RECT 55.750 103.710 55.950 104.410 ;
        RECT 76.690 104.230 81.060 104.410 ;
        RECT 78.410 104.220 79.530 104.230 ;
        RECT 51.470 103.560 55.950 103.710 ;
        RECT 51.470 103.490 55.920 103.560 ;
        RECT 51.470 103.430 51.780 103.490 ;
        RECT 45.540 103.180 49.670 103.390 ;
        RECT 49.460 103.040 49.670 103.180 ;
        RECT 51.420 103.040 51.730 103.110 ;
        RECT 49.460 102.830 51.730 103.040 ;
        RECT 51.120 102.820 51.730 102.830 ;
        RECT 46.930 102.740 47.240 102.810 ;
        RECT 51.420 102.780 51.730 102.820 ;
        RECT 46.930 102.690 49.260 102.740 ;
        RECT 44.390 102.530 49.260 102.690 ;
        RECT 87.700 102.640 88.600 102.650 ;
        RECT 44.390 102.470 47.240 102.530 ;
        RECT 51.420 102.240 51.730 102.250 ;
        RECT 45.460 102.190 51.730 102.240 ;
        RECT 41.090 102.030 51.730 102.190 ;
        RECT 35.150 101.980 36.040 102.000 ;
        RECT 35.610 101.960 35.920 101.980 ;
        RECT 41.090 101.970 45.850 102.030 ;
        RECT 51.120 102.000 51.730 102.030 ;
        RECT 51.420 101.920 51.730 102.000 ;
        RECT 28.470 101.650 28.780 101.790 ;
        RECT 25.970 101.640 28.780 101.650 ;
        RECT 46.780 101.650 47.090 101.790 ;
        RECT 84.960 101.730 85.740 101.880 ;
        RECT 87.700 101.730 190.930 102.640 ;
        RECT 46.780 101.640 49.260 101.650 ;
        RECT 25.970 101.490 49.260 101.640 ;
        RECT 25.970 101.470 28.780 101.490 ;
        RECT 28.470 101.460 28.780 101.470 ;
        RECT 46.780 101.470 49.260 101.490 ;
        RECT 51.470 101.550 51.780 101.600 ;
        RECT 53.680 101.550 53.990 101.590 ;
        RECT 46.780 101.460 47.090 101.470 ;
        RECT 51.470 101.320 54.180 101.550 ;
        RECT 51.470 101.270 51.780 101.320 ;
        RECT 53.680 101.260 53.990 101.320 ;
        RECT 84.960 101.260 190.930 101.730 ;
        RECT 84.960 101.110 85.740 101.260 ;
        RECT 29.110 100.710 29.430 100.720 ;
        RECT 56.920 100.710 57.380 100.780 ;
        RECT 29.110 100.430 57.380 100.710 ;
        RECT 87.700 100.560 190.930 101.260 ;
        RECT 88.580 100.550 190.930 100.560 ;
        RECT 29.110 100.380 29.430 100.430 ;
        RECT 56.920 100.370 57.380 100.430 ;
        RECT 57.710 100.110 58.140 100.190 ;
        RECT 46.450 99.850 58.140 100.110 ;
        RECT 46.450 99.840 46.770 99.850 ;
        RECT 57.710 99.780 58.140 99.850 ;
        RECT 13.140 99.160 15.580 99.380 ;
        RECT 13.240 98.360 13.500 99.160 ;
        RECT 15.240 99.100 15.580 99.160 ;
        RECT 21.110 99.070 21.430 99.120 ;
        RECT 23.520 99.070 23.840 99.090 ;
        RECT 21.110 99.050 25.590 99.070 ;
        RECT 25.890 99.050 26.070 99.060 ;
        RECT 21.110 98.940 26.070 99.050 ;
        RECT 29.870 98.940 30.180 99.080 ;
        RECT 45.360 98.940 45.670 99.080 ;
        RECT 21.110 98.900 47.830 98.940 ;
        RECT 21.110 98.880 23.840 98.900 ;
        RECT 21.110 98.800 21.430 98.880 ;
        RECT 23.520 98.830 23.840 98.880 ;
        RECT 25.550 98.870 47.830 98.900 ;
        RECT 25.890 98.760 47.830 98.870 ;
        RECT 29.870 98.750 30.180 98.760 ;
        RECT 45.360 98.750 45.670 98.760 ;
        RECT 16.940 98.640 17.260 98.660 ;
        RECT 16.930 98.590 17.260 98.640 ;
        RECT 17.970 98.590 18.290 98.600 ;
        RECT 16.930 98.390 20.350 98.590 ;
        RECT 47.680 98.560 48.240 98.740 ;
        RECT 29.870 98.510 30.180 98.530 ;
        RECT 45.360 98.510 45.670 98.530 ;
        RECT 16.930 98.380 17.260 98.390 ;
        RECT 16.940 98.370 17.260 98.380 ;
        RECT 17.970 98.340 18.290 98.390 ;
        RECT 19.870 98.360 20.350 98.390 ;
        RECT 20.010 98.290 20.350 98.360 ;
        RECT 27.710 98.500 30.270 98.510 ;
        RECT 45.270 98.500 47.830 98.510 ;
        RECT 27.710 98.330 47.830 98.500 ;
        RECT 29.870 98.320 45.670 98.330 ;
        RECT 29.870 98.200 30.180 98.320 ;
        RECT 45.360 98.200 45.670 98.320 ;
        RECT 58.450 97.740 58.890 97.860 ;
        RECT 13.140 97.410 15.580 97.630 ;
        RECT 58.320 97.560 58.890 97.740 ;
        RECT -117.910 96.290 -15.700 96.660 ;
        RECT 13.240 96.610 13.500 97.410 ;
        RECT 15.240 97.350 15.580 97.410 ;
        RECT 29.870 97.400 30.180 97.530 ;
        RECT 45.360 97.400 45.670 97.530 ;
        RECT 58.440 97.460 58.890 97.560 ;
        RECT 87.700 97.760 88.600 97.770 ;
        RECT 58.440 97.400 58.840 97.460 ;
        RECT 20.010 97.250 20.350 97.320 ;
        RECT 19.870 97.200 20.350 97.250 ;
        RECT 27.710 97.220 58.840 97.400 ;
        RECT 29.870 97.200 30.180 97.220 ;
        RECT 45.360 97.200 45.670 97.220 ;
        RECT 19.670 97.190 20.350 97.200 ;
        RECT 19.650 97.020 20.350 97.190 ;
        RECT 16.940 96.890 17.260 96.910 ;
        RECT 16.930 96.840 17.260 96.890 ;
        RECT 17.970 96.840 18.290 96.850 ;
        RECT 19.650 96.840 19.850 97.020 ;
        RECT 29.870 96.970 30.180 96.980 ;
        RECT 45.360 96.970 45.670 96.980 ;
        RECT 16.930 96.640 19.850 96.840 ;
        RECT 25.630 96.810 47.830 96.970 ;
        RECT 21.110 96.730 21.430 96.810 ;
        RECT 23.590 96.790 47.830 96.810 ;
        RECT 23.590 96.780 25.810 96.790 ;
        RECT 23.520 96.730 25.810 96.780 ;
        RECT 21.110 96.650 25.810 96.730 ;
        RECT 29.870 96.650 30.180 96.790 ;
        RECT 45.360 96.650 45.670 96.790 ;
        RECT 64.980 96.740 65.580 96.800 ;
        RECT 87.700 96.740 186.850 97.760 ;
        RECT 16.930 96.630 17.260 96.640 ;
        RECT 16.940 96.620 17.260 96.630 ;
        RECT 17.970 96.590 18.290 96.640 ;
        RECT 21.110 96.540 23.840 96.650 ;
        RECT 24.320 96.640 25.810 96.650 ;
        RECT 25.020 96.630 25.810 96.640 ;
        RECT 21.110 96.490 21.430 96.540 ;
        RECT 23.520 96.520 23.840 96.540 ;
        RECT -117.910 95.690 -25.730 96.290 ;
        RECT 64.980 96.270 186.850 96.740 ;
        RECT 64.980 96.220 65.580 96.270 ;
        RECT -117.910 95.630 -26.950 95.690 ;
        RECT 13.140 95.660 15.580 95.880 ;
        RECT -122.660 29.240 -120.090 32.840 ;
        RECT -122.450 29.200 -120.370 29.240 ;
        RECT -117.910 4.220 -115.830 95.630 ;
        RECT 13.240 94.860 13.500 95.660 ;
        RECT 15.240 95.600 15.580 95.660 ;
        RECT 21.110 95.870 21.430 95.920 ;
        RECT 23.520 95.870 23.840 95.890 ;
        RECT 21.110 95.850 23.840 95.870 ;
        RECT 21.110 95.840 25.830 95.850 ;
        RECT 21.110 95.700 25.840 95.840 ;
        RECT 29.870 95.700 30.180 95.840 ;
        RECT 45.360 95.700 45.670 95.840 ;
        RECT 21.110 95.690 47.830 95.700 ;
        RECT 21.110 95.680 23.840 95.690 ;
        RECT 21.110 95.600 21.430 95.680 ;
        RECT 23.520 95.630 23.840 95.680 ;
        RECT 25.660 95.520 47.830 95.690 ;
        RECT 87.700 95.680 186.850 96.270 ;
        RECT 88.580 95.670 186.850 95.680 ;
        RECT 29.870 95.510 30.180 95.520 ;
        RECT 45.360 95.510 45.670 95.520 ;
        RECT 19.870 95.370 20.350 95.390 ;
        RECT 16.940 95.140 17.260 95.160 ;
        RECT 16.930 95.090 17.260 95.140 ;
        RECT 17.970 95.090 18.290 95.100 ;
        RECT 19.600 95.090 20.350 95.370 ;
        RECT 29.870 95.270 30.180 95.290 ;
        RECT 45.360 95.270 45.670 95.290 ;
        RECT 27.710 95.090 47.830 95.270 ;
        RECT 16.930 95.040 20.090 95.090 ;
        RECT 16.930 94.890 19.950 95.040 ;
        RECT 29.870 94.960 30.180 95.090 ;
        RECT 45.360 94.960 45.670 95.090 ;
        RECT 16.930 94.880 17.260 94.890 ;
        RECT 16.940 94.870 17.260 94.880 ;
        RECT 17.970 94.840 18.290 94.890 ;
        RECT 29.870 94.170 30.180 94.300 ;
        RECT 45.360 94.170 45.670 94.300 ;
        RECT 13.140 93.910 15.580 94.130 ;
        RECT 20.010 94.050 20.350 94.120 ;
        RECT -113.560 93.350 -26.950 93.450 ;
        RECT -113.560 92.510 -25.790 93.350 ;
        RECT 13.240 93.110 13.500 93.910 ;
        RECT 15.240 93.850 15.580 93.910 ;
        RECT 19.640 93.820 20.350 94.050 ;
        RECT 27.710 93.990 47.830 94.170 ;
        RECT 29.870 93.970 30.180 93.990 ;
        RECT 45.360 93.970 45.670 93.990 ;
        RECT 16.940 93.390 17.260 93.410 ;
        RECT 16.930 93.340 17.260 93.390 ;
        RECT 17.970 93.340 18.290 93.350 ;
        RECT 19.640 93.340 19.840 93.820 ;
        RECT 29.870 93.740 30.180 93.750 ;
        RECT 45.360 93.740 45.670 93.750 ;
        RECT 16.930 93.140 19.840 93.340 ;
        RECT 21.110 93.530 21.430 93.610 ;
        RECT 23.520 93.550 23.840 93.580 ;
        RECT 25.630 93.570 47.830 93.740 ;
        RECT 25.630 93.560 30.180 93.570 ;
        RECT 25.640 93.550 25.820 93.560 ;
        RECT 23.520 93.530 25.820 93.550 ;
        RECT 21.110 93.370 25.820 93.530 ;
        RECT 29.870 93.420 30.180 93.560 ;
        RECT 45.360 93.560 47.830 93.570 ;
        RECT 45.360 93.420 45.670 93.560 ;
        RECT 21.110 93.340 23.840 93.370 ;
        RECT 21.110 93.290 21.430 93.340 ;
        RECT 23.520 93.320 23.840 93.340 ;
        RECT 16.930 93.130 17.260 93.140 ;
        RECT 16.940 93.120 17.260 93.130 ;
        RECT 17.970 93.090 18.290 93.140 ;
        RECT -11.890 92.770 -11.580 92.790 ;
        RECT -11.230 92.770 -10.920 92.790 ;
        RECT -113.560 92.140 -17.360 92.510 ;
        RECT -11.890 92.300 -4.570 92.770 ;
        RECT -11.890 92.280 -11.580 92.300 ;
        RECT -11.230 92.280 -10.920 92.300 ;
        RECT -113.560 91.470 -25.790 92.140 ;
        RECT -113.560 91.370 -26.950 91.470 ;
        RECT -118.070 0.650 -115.680 4.220 ;
        RECT -117.910 0.120 -115.830 0.650 ;
        RECT -113.560 -24.390 -111.480 91.370 ;
        RECT -17.730 90.790 -17.360 92.140 ;
        RECT -5.040 91.620 -4.570 92.300 ;
        RECT 21.730 92.630 22.040 92.650 ;
        RECT 59.370 92.630 59.820 92.660 ;
        RECT 21.730 92.220 59.820 92.630 ;
        RECT 21.730 92.200 22.040 92.220 ;
        RECT 59.370 92.200 59.820 92.220 ;
        RECT 87.730 92.560 88.630 92.590 ;
        RECT 87.730 91.620 182.760 92.560 ;
        RECT -13.220 91.490 -12.960 91.560 ;
        RECT -11.170 91.490 -10.850 91.510 ;
        RECT -9.410 91.490 -9.080 91.530 ;
        RECT -13.220 91.300 -9.080 91.490 ;
        RECT -13.220 91.240 -12.960 91.300 ;
        RECT -11.170 91.250 -10.850 91.300 ;
        RECT -9.410 91.260 -9.080 91.300 ;
        RECT -5.040 91.150 182.760 91.620 ;
        RECT -13.770 91.090 -13.450 91.130 ;
        RECT -11.830 91.090 -11.510 91.150 ;
        RECT -8.910 91.090 -8.590 91.130 ;
        RECT -13.770 90.900 -8.590 91.090 ;
        RECT 63.890 91.030 64.460 91.150 ;
        RECT -13.770 90.870 -13.450 90.900 ;
        RECT -11.830 90.890 -11.510 90.900 ;
        RECT -8.910 90.870 -8.590 90.900 ;
        RECT -17.730 90.780 -15.700 90.790 ;
        RECT -17.730 90.600 -15.480 90.780 ;
        RECT -17.730 90.540 -14.080 90.600 ;
        RECT -11.080 90.540 -10.770 90.580 ;
        RECT -17.730 90.420 -10.770 90.540 ;
        RECT -16.070 90.380 -10.770 90.420 ;
        RECT -15.700 90.320 -10.770 90.380 ;
        RECT -23.070 90.130 -22.300 90.320 ;
        RECT -11.080 90.250 -10.770 90.320 ;
        RECT -10.430 90.510 -10.120 90.580 ;
        RECT -7.430 90.530 -7.130 90.550 ;
        RECT -7.440 90.510 -7.120 90.530 ;
        RECT -10.430 90.300 -7.120 90.510 ;
        RECT 87.730 90.500 182.760 91.150 ;
        RECT 88.580 90.470 182.760 90.500 ;
        RECT -10.430 90.250 -10.120 90.300 ;
        RECT -9.660 90.290 -7.120 90.300 ;
        RECT -16.070 90.130 -15.680 90.150 ;
        RECT -23.070 90.090 -15.680 90.130 ;
        RECT -12.300 90.090 -11.990 90.140 ;
        RECT -23.070 89.880 -11.990 90.090 ;
        RECT -23.070 89.760 -15.690 89.880 ;
        RECT -12.300 89.810 -11.990 89.880 ;
        RECT -11.600 90.070 -11.290 90.140 ;
        RECT -9.660 90.070 -9.440 90.290 ;
        RECT -7.440 90.270 -7.120 90.290 ;
        RECT -7.430 90.250 -7.130 90.270 ;
        RECT 13.100 90.100 15.540 90.320 ;
        RECT -11.600 89.850 -9.440 90.070 ;
        RECT -11.600 89.810 -11.290 89.850 ;
        RECT -23.070 89.580 -22.300 89.760 ;
        RECT -16.070 89.740 -15.700 89.760 ;
        RECT -109.220 89.250 -26.950 89.380 ;
        RECT 13.200 89.300 13.460 90.100 ;
        RECT 15.200 90.040 15.540 90.100 ;
        RECT 21.140 89.800 21.460 89.850 ;
        RECT 23.550 89.800 23.870 89.820 ;
        RECT 21.140 89.790 25.620 89.800 ;
        RECT 21.140 89.630 25.750 89.790 ;
        RECT 21.140 89.610 23.870 89.630 ;
        RECT 25.440 89.610 25.750 89.630 ;
        RECT 29.900 89.610 30.210 89.750 ;
        RECT 16.900 89.580 17.220 89.600 ;
        RECT 16.890 89.530 17.220 89.580 ;
        RECT 17.930 89.530 18.250 89.540 ;
        RECT 21.140 89.530 21.460 89.610 ;
        RECT 23.550 89.560 23.870 89.610 ;
        RECT 16.890 89.330 19.970 89.530 ;
        RECT 25.570 89.430 30.210 89.610 ;
        RECT 29.900 89.420 30.210 89.430 ;
        RECT 30.500 89.590 30.820 89.610 ;
        RECT 30.500 89.400 38.420 89.590 ;
        RECT 38.580 89.400 38.890 89.440 ;
        RECT 30.500 89.380 38.890 89.400 ;
        RECT 30.500 89.350 30.820 89.380 ;
        RECT 16.890 89.320 17.220 89.330 ;
        RECT 16.900 89.310 17.220 89.320 ;
        RECT 17.930 89.280 18.250 89.330 ;
        RECT 19.770 89.320 19.970 89.330 ;
        RECT -109.220 88.480 -25.730 89.250 ;
        RECT 19.770 89.090 20.380 89.320 ;
        RECT 38.210 89.190 38.890 89.380 ;
        RECT 38.580 89.110 38.890 89.190 ;
        RECT 20.040 89.020 20.380 89.090 ;
        RECT 27.230 88.950 27.380 88.970 ;
        RECT 26.210 88.800 27.380 88.950 ;
        RECT -12.750 88.740 -12.430 88.760 ;
        RECT -12.970 88.520 -12.430 88.740 ;
        RECT -12.750 88.500 -12.430 88.520 ;
        RECT -109.220 88.110 -21.010 88.480 ;
        RECT 13.100 88.350 15.540 88.570 ;
        RECT 26.150 88.470 26.430 88.800 ;
        RECT 27.230 88.550 27.380 88.800 ;
        RECT 30.480 88.550 30.800 88.560 ;
        RECT 27.230 88.400 30.800 88.550 ;
        RECT -10.000 88.160 -9.680 88.280 ;
        RECT -109.220 87.370 -25.730 88.110 ;
        RECT -109.220 87.300 -26.950 87.370 ;
        RECT -113.740 -27.910 -111.290 -24.390 ;
        RECT -113.560 -28.030 -111.480 -27.910 ;
        RECT -109.220 -52.900 -107.140 87.300 ;
        RECT -21.380 86.450 -21.010 88.110 ;
        RECT -12.970 87.960 -9.680 88.160 ;
        RECT -12.970 87.950 -9.990 87.960 ;
        RECT -12.970 87.740 -9.990 87.760 ;
        RECT -12.970 87.550 -9.670 87.740 ;
        RECT 13.200 87.550 13.460 88.350 ;
        RECT 15.200 88.290 15.540 88.350 ;
        RECT 30.360 88.300 30.800 88.400 ;
        RECT 20.040 87.980 20.380 88.050 ;
        RECT 19.900 87.940 20.380 87.980 ;
        RECT 16.900 87.830 17.220 87.850 ;
        RECT 16.890 87.780 17.220 87.830 ;
        RECT 17.930 87.780 18.250 87.790 ;
        RECT 19.760 87.780 20.380 87.940 ;
        RECT 27.210 87.800 27.530 88.070 ;
        RECT 16.890 87.750 20.380 87.780 ;
        RECT 16.890 87.580 20.080 87.750 ;
        RECT 29.900 87.660 30.210 87.670 ;
        RECT 16.890 87.570 17.220 87.580 ;
        RECT 16.900 87.560 17.220 87.570 ;
        RECT -9.990 87.420 -9.670 87.550 ;
        RECT 17.930 87.530 18.250 87.580 ;
        RECT 25.550 87.540 30.210 87.660 ;
        RECT 21.140 87.460 21.460 87.540 ;
        RECT 23.620 87.510 30.210 87.540 ;
        RECT 88.580 87.510 178.630 87.520 ;
        RECT 23.550 87.500 30.210 87.510 ;
        RECT 23.550 87.480 30.300 87.500 ;
        RECT 23.550 87.460 25.730 87.480 ;
        RECT 21.140 87.380 25.730 87.460 ;
        RECT 21.140 87.270 23.870 87.380 ;
        RECT 24.350 87.370 25.730 87.380 ;
        RECT 25.050 87.360 25.730 87.370 ;
        RECT -13.740 87.220 -13.450 87.230 ;
        RECT 21.140 87.220 21.460 87.270 ;
        RECT 23.550 87.250 23.870 87.270 ;
        RECT 25.410 87.330 25.730 87.360 ;
        RECT 29.900 87.360 30.300 87.480 ;
        RECT 29.900 87.340 30.210 87.360 ;
        RECT 25.410 87.250 25.590 87.330 ;
        RECT 30.440 87.320 30.670 87.330 ;
        RECT 30.440 87.290 38.010 87.320 ;
        RECT -13.750 87.200 -13.430 87.220 ;
        RECT -12.750 87.200 -12.430 87.210 ;
        RECT -13.750 86.980 -12.430 87.200 ;
        RECT 30.440 87.120 38.070 87.290 ;
        RECT 38.580 87.120 38.890 87.200 ;
        RECT -13.750 86.960 -13.430 86.980 ;
        RECT -13.740 86.940 -13.450 86.960 ;
        RECT -12.750 86.950 -12.430 86.980 ;
        RECT 27.190 87.020 27.510 87.050 ;
        RECT 30.440 87.020 30.680 87.120 ;
        RECT 27.190 86.840 30.680 87.020 ;
        RECT 37.880 86.920 38.890 87.120 ;
        RECT 38.480 86.910 38.890 86.920 ;
        RECT 38.580 86.870 38.890 86.910 ;
        RECT 27.190 86.820 30.600 86.840 ;
        RECT 13.100 86.600 15.540 86.820 ;
        RECT 27.190 86.790 27.510 86.820 ;
        RECT -21.380 86.270 -15.430 86.450 ;
        RECT -21.380 86.200 -15.360 86.270 ;
        RECT -13.970 86.200 -12.700 86.210 ;
        RECT -12.270 86.200 -11.960 86.260 ;
        RECT -21.380 86.080 -11.960 86.200 ;
        RECT -16.070 86.040 -11.960 86.080 ;
        RECT -15.710 85.990 -11.960 86.040 ;
        RECT -12.270 85.930 -11.960 85.990 ;
        RECT -11.580 86.180 -11.270 86.250 ;
        RECT -6.790 86.200 -6.500 86.220 ;
        RECT -11.580 86.170 -9.440 86.180 ;
        RECT -6.800 86.170 -6.480 86.200 ;
        RECT -11.580 85.970 -6.480 86.170 ;
        RECT -11.580 85.920 -11.270 85.970 ;
        RECT -9.650 85.960 -6.480 85.970 ;
        RECT -17.840 85.470 -17.430 85.490 ;
        RECT -16.070 85.470 -14.080 85.490 ;
        RECT -17.840 85.430 -14.080 85.470 ;
        RECT -11.100 85.430 -10.790 85.480 ;
        RECT -105.060 85.160 -26.950 85.230 ;
        RECT -17.840 85.210 -10.790 85.430 ;
        RECT -105.060 84.340 -25.730 85.160 ;
        RECT -17.840 85.100 -15.690 85.210 ;
        RECT -11.100 85.150 -10.790 85.210 ;
        RECT -10.390 85.350 -10.080 85.420 ;
        RECT -9.650 85.350 -9.440 85.960 ;
        RECT -6.800 85.940 -6.480 85.960 ;
        RECT -6.790 85.920 -6.500 85.940 ;
        RECT 13.200 85.800 13.460 86.600 ;
        RECT 15.200 86.540 15.540 86.600 ;
        RECT 21.140 86.600 21.460 86.650 ;
        RECT 30.480 86.640 30.800 86.680 ;
        RECT 30.480 86.620 38.030 86.640 ;
        RECT 38.580 86.630 38.890 86.670 ;
        RECT 38.480 86.620 38.890 86.630 ;
        RECT 23.550 86.600 23.870 86.620 ;
        RECT 21.140 86.580 23.870 86.600 ;
        RECT 21.140 86.420 25.660 86.580 ;
        RECT 21.140 86.410 23.870 86.420 ;
        RECT 21.140 86.330 21.460 86.410 ;
        RECT 23.550 86.360 23.870 86.410 ;
        RECT 25.480 86.370 25.660 86.420 ;
        RECT 29.900 86.380 30.210 86.510 ;
        RECT 30.480 86.420 38.890 86.620 ;
        RECT 30.580 86.410 30.900 86.420 ;
        RECT 29.900 86.370 30.330 86.380 ;
        RECT 25.480 86.210 30.330 86.370 ;
        RECT 38.580 86.340 38.890 86.420 ;
        RECT 62.770 86.380 63.320 86.390 ;
        RECT 62.770 86.360 63.330 86.380 ;
        RECT 87.700 86.360 178.630 87.510 ;
        RECT 25.480 86.190 30.210 86.210 ;
        RECT 29.900 86.180 30.210 86.190 ;
        RECT 16.900 86.080 17.220 86.100 ;
        RECT 16.890 86.030 17.220 86.080 ;
        RECT 17.930 86.030 18.250 86.040 ;
        RECT 19.900 86.030 20.380 86.120 ;
        RECT 16.890 85.830 20.380 86.030 ;
        RECT 16.890 85.820 17.220 85.830 ;
        RECT 16.900 85.810 17.220 85.820 ;
        RECT 17.930 85.780 18.250 85.830 ;
        RECT 19.840 85.820 20.380 85.830 ;
        RECT 26.760 85.960 27.080 86.000 ;
        RECT 19.840 85.740 20.130 85.820 ;
        RECT 26.760 85.680 27.370 85.960 ;
        RECT 29.900 85.940 30.210 85.960 ;
        RECT 27.740 85.770 37.040 85.940 ;
        RECT 62.770 85.890 178.630 86.360 ;
        RECT 62.770 85.880 63.330 85.890 ;
        RECT 62.770 85.860 63.320 85.880 ;
        RECT 27.740 85.760 30.300 85.770 ;
        RECT -10.390 85.140 -9.440 85.350 ;
        RECT 27.170 85.460 27.370 85.680 ;
        RECT 29.900 85.630 30.210 85.760 ;
        RECT 30.350 85.460 30.670 85.500 ;
        RECT 27.170 85.260 30.720 85.460 ;
        RECT 87.700 85.430 178.630 85.890 ;
        RECT 87.700 85.420 88.600 85.430 ;
        RECT 30.350 85.240 30.670 85.260 ;
        RECT -17.840 85.080 -17.430 85.100 ;
        RECT -16.070 85.080 -15.700 85.100 ;
        RECT -10.390 85.090 -10.080 85.140 ;
        RECT 13.100 84.850 15.540 85.070 ;
        RECT 19.820 84.860 20.120 84.900 ;
        RECT -23.070 84.340 -22.270 84.480 ;
        RECT -105.060 83.840 -22.270 84.340 ;
        RECT 13.200 84.050 13.460 84.850 ;
        RECT 15.200 84.790 15.540 84.850 ;
        RECT 19.810 84.850 20.120 84.860 ;
        RECT 19.810 84.550 20.380 84.850 ;
        RECT 27.140 84.720 27.450 85.050 ;
        RECT 16.900 84.330 17.220 84.350 ;
        RECT 16.890 84.280 17.220 84.330 ;
        RECT 17.930 84.280 18.250 84.290 ;
        RECT 19.810 84.280 20.010 84.550 ;
        RECT 29.900 84.410 30.210 84.420 ;
        RECT 16.890 84.080 20.010 84.280 ;
        RECT 21.140 84.260 21.460 84.340 ;
        RECT 23.550 84.280 23.870 84.310 ;
        RECT 25.720 84.280 30.210 84.410 ;
        RECT 38.580 84.370 38.890 84.430 ;
        RECT 38.030 84.360 38.890 84.370 ;
        RECT 23.550 84.260 30.210 84.280 ;
        RECT 21.140 84.230 30.210 84.260 ;
        RECT 21.140 84.100 25.900 84.230 ;
        RECT 16.890 84.070 17.220 84.080 ;
        RECT 16.900 84.060 17.220 84.070 ;
        RECT 17.930 84.030 18.250 84.080 ;
        RECT 21.140 84.070 23.870 84.100 ;
        RECT 29.900 84.090 30.210 84.230 ;
        RECT 30.450 84.140 38.890 84.360 ;
        RECT 30.450 84.130 38.040 84.140 ;
        RECT 30.450 84.120 31.220 84.130 ;
        RECT 21.140 84.020 21.460 84.070 ;
        RECT 23.550 84.050 23.870 84.070 ;
        RECT 27.190 84.080 27.500 84.090 ;
        RECT -105.060 83.280 -25.730 83.840 ;
        RECT -23.070 83.710 -22.270 83.840 ;
        RECT 27.190 83.950 27.550 84.080 ;
        RECT 30.450 83.950 30.690 84.120 ;
        RECT 38.580 84.100 38.890 84.140 ;
        RECT 27.190 83.710 30.690 83.950 ;
        RECT 19.550 83.580 19.870 83.630 ;
        RECT 26.160 83.580 26.480 83.680 ;
        RECT 19.550 83.420 26.480 83.580 ;
        RECT 19.550 83.370 19.870 83.420 ;
        RECT 26.160 83.400 26.480 83.420 ;
        RECT 27.190 83.580 27.510 83.710 ;
        RECT 37.810 83.580 38.220 83.690 ;
        RECT 27.190 83.420 38.220 83.580 ;
        RECT 27.190 83.390 27.510 83.420 ;
        RECT 26.750 83.340 27.030 83.350 ;
        RECT -105.060 83.150 -26.950 83.280 ;
        RECT 26.730 83.250 27.050 83.340 ;
        RECT 37.810 83.320 38.220 83.420 ;
        RECT 28.970 83.250 29.290 83.280 ;
        RECT -109.470 -56.630 -106.870 -52.900 ;
        RECT -109.220 -56.960 -107.140 -56.630 ;
        RECT -105.060 -81.530 -102.980 83.150 ;
        RECT 26.700 83.090 29.290 83.250 ;
        RECT 26.730 83.080 27.050 83.090 ;
        RECT 26.750 83.070 27.030 83.080 ;
        RECT 28.970 83.020 29.290 83.090 ;
        RECT 28.990 83.010 29.270 83.020 ;
        RECT 27.770 82.100 28.150 82.130 ;
        RECT 29.120 82.120 32.180 82.130 ;
        RECT 19.310 82.090 22.370 82.100 ;
        RECT 19.220 81.760 22.370 82.090 ;
        RECT 24.870 81.760 28.150 82.100 ;
        RECT 29.030 82.040 32.180 82.120 ;
        RECT 19.220 81.080 19.540 81.760 ;
        RECT 22.040 81.750 22.350 81.760 ;
        RECT 24.890 81.750 25.200 81.760 ;
        RECT 19.070 80.700 19.540 81.080 ;
        RECT -100.810 80.010 -26.950 80.080 ;
        RECT -11.070 80.070 -10.460 80.400 ;
        RECT -100.810 79.230 -25.790 80.010 ;
        RECT -13.280 79.960 -12.970 79.970 ;
        RECT -12.190 79.960 -11.880 79.970 ;
        RECT -14.600 79.950 -11.880 79.960 ;
        RECT -14.830 79.640 -11.880 79.950 ;
        RECT -14.830 79.630 -11.890 79.640 ;
        RECT -17.830 79.230 -17.420 79.250 ;
        RECT -100.810 78.860 -17.420 79.230 ;
        RECT -100.810 78.130 -25.790 78.860 ;
        RECT -17.830 78.840 -17.420 78.860 ;
        RECT -100.810 78.000 -26.950 78.130 ;
        RECT -105.480 -85.200 -102.770 -81.530 ;
        RECT -105.060 -85.920 -102.980 -85.200 ;
        RECT -100.810 -110.150 -98.730 78.000 ;
        RECT -14.830 77.190 -14.480 79.630 ;
        RECT -11.060 79.580 -10.460 80.070 ;
        RECT 19.220 79.310 19.540 80.700 ;
        RECT 27.700 81.740 28.150 81.760 ;
        RECT 28.920 81.790 32.180 82.040 ;
        RECT 34.680 82.120 37.740 82.130 ;
        RECT 34.680 81.900 37.830 82.120 ;
        RECT 88.900 82.000 174.390 82.010 ;
        RECT 34.680 81.790 38.170 81.900 ;
        RECT 27.700 79.310 28.020 81.740 ;
        RECT 28.920 81.700 29.350 81.790 ;
        RECT 31.850 81.780 32.160 81.790 ;
        RECT 34.700 81.780 35.010 81.790 ;
        RECT -13.830 79.280 -13.520 79.290 ;
        RECT -12.730 79.280 -12.420 79.290 ;
        RECT -11.630 79.280 -11.320 79.290 ;
        RECT -13.860 78.960 -10.700 79.280 ;
        RECT -11.020 77.920 -10.700 78.960 ;
        RECT -13.860 77.590 -10.700 77.920 ;
        RECT 19.220 78.980 22.380 79.310 ;
        RECT 24.860 78.980 28.020 79.310 ;
        RECT 19.220 77.940 19.540 78.980 ;
        RECT 27.700 77.940 28.020 78.980 ;
        RECT 19.220 77.620 22.380 77.940 ;
        RECT 24.860 77.620 28.020 77.940 ;
        RECT 29.030 79.340 29.350 81.700 ;
        RECT 37.510 81.540 38.170 81.790 ;
        RECT 37.510 79.340 37.830 81.540 ;
        RECT 40.990 81.400 41.300 81.410 ;
        RECT 42.080 81.400 42.390 81.430 ;
        RECT 39.440 81.250 42.390 81.400 ;
        RECT 39.260 81.100 42.390 81.250 ;
        RECT 39.260 81.060 40.190 81.100 ;
        RECT 40.990 81.080 41.300 81.100 ;
        RECT 61.720 81.060 62.320 81.110 ;
        RECT 88.130 81.060 174.390 82.000 ;
        RECT 39.260 80.930 39.820 81.060 ;
        RECT 39.260 80.820 39.790 80.930 ;
        RECT 29.030 79.010 32.190 79.340 ;
        RECT 34.670 79.010 37.830 79.340 ;
        RECT 29.030 77.970 29.350 79.010 ;
        RECT 37.510 77.970 37.830 79.010 ;
        RECT 29.030 77.650 32.190 77.970 ;
        RECT 34.670 77.650 37.830 77.970 ;
        RECT 39.440 80.060 39.790 80.820 ;
        RECT 61.720 80.590 174.390 81.060 ;
        RECT 61.720 80.550 62.320 80.590 ;
        RECT 39.440 79.730 42.390 80.060 ;
        RECT 88.130 79.920 174.390 80.590 ;
        RECT 88.150 79.910 88.920 79.920 ;
        RECT 29.650 77.640 29.960 77.650 ;
        RECT 30.750 77.640 31.060 77.650 ;
        RECT 31.850 77.640 32.160 77.650 ;
        RECT 34.700 77.640 35.010 77.650 ;
        RECT 35.800 77.640 36.110 77.650 ;
        RECT 36.900 77.640 37.210 77.650 ;
        RECT 19.840 77.610 20.150 77.620 ;
        RECT 20.940 77.610 21.250 77.620 ;
        RECT 22.040 77.610 22.350 77.620 ;
        RECT 24.890 77.610 25.200 77.620 ;
        RECT 25.990 77.610 26.300 77.620 ;
        RECT 27.090 77.610 27.400 77.620 ;
        RECT -14.830 76.860 -11.880 77.190 ;
        RECT -14.830 75.990 -14.480 76.860 ;
        RECT -14.830 75.860 -14.450 75.990 ;
        RECT -16.110 75.840 -15.740 75.850 ;
        RECT -14.830 75.840 -14.080 75.860 ;
        RECT -17.430 75.820 -14.080 75.840 ;
        RECT -13.280 75.820 -12.970 75.840 ;
        RECT -96.550 75.720 -26.950 75.820 ;
        RECT -96.550 75.020 -25.730 75.720 ;
        RECT -17.430 75.520 -11.880 75.820 ;
        RECT -17.430 75.460 -14.820 75.520 ;
        RECT -13.280 75.510 -12.970 75.520 ;
        RECT -12.190 75.490 -11.880 75.520 ;
        RECT -17.430 75.020 -17.050 75.460 ;
        RECT -16.110 75.440 -15.740 75.460 ;
        RECT -13.830 75.140 -13.520 75.150 ;
        RECT -11.020 75.140 -10.700 77.590 ;
        RECT 18.980 76.830 19.580 77.320 ;
        RECT 27.660 76.830 28.260 77.320 ;
        RECT 18.980 76.500 19.590 76.830 ;
        RECT 27.650 76.500 28.260 76.830 ;
        RECT 28.790 76.860 29.390 77.350 ;
        RECT 37.470 76.860 38.070 77.350 ;
        RECT 39.440 77.290 39.790 79.730 ;
        RECT 39.440 77.280 42.380 77.290 ;
        RECT 39.440 76.970 42.390 77.280 ;
        RECT 39.670 76.960 42.390 76.970 ;
        RECT 40.990 76.950 41.300 76.960 ;
        RECT 42.080 76.950 42.390 76.960 ;
        RECT 28.790 76.530 29.400 76.860 ;
        RECT 37.460 76.530 38.070 76.860 ;
        RECT 43.210 76.850 43.810 77.340 ;
        RECT 43.200 76.520 43.810 76.850 ;
        RECT 19.160 75.470 19.660 75.480 ;
        RECT 65.090 75.470 65.650 75.490 ;
        RECT -7.440 75.140 -7.160 75.150 ;
        RECT -96.550 74.640 -17.050 75.020 ;
        RECT -13.850 74.810 -7.140 75.140 ;
        RECT 19.160 75.010 65.650 75.470 ;
        RECT 19.160 74.950 19.680 75.010 ;
        RECT 65.090 74.990 65.650 75.010 ;
        RECT 19.160 74.930 19.660 74.950 ;
        RECT -13.850 74.800 -10.790 74.810 ;
        RECT -7.440 74.790 -7.160 74.810 ;
        RECT -96.550 73.840 -25.730 74.640 ;
        RECT 27.470 74.100 64.550 74.560 ;
        RECT 27.540 74.000 28.060 74.100 ;
        RECT 63.900 74.040 64.460 74.100 ;
        RECT -96.550 73.740 -26.950 73.840 ;
        RECT -101.140 -113.630 -98.400 -110.150 ;
        RECT -100.810 -114.440 -98.730 -113.630 ;
        RECT -96.550 -138.440 -94.470 73.740 ;
        RECT 28.910 73.580 63.460 73.650 ;
        RECT 28.900 73.190 63.460 73.580 ;
        RECT 28.900 73.060 29.550 73.190 ;
        RECT 62.770 73.170 63.330 73.190 ;
        RECT -11.030 72.830 -10.420 72.850 ;
        RECT -11.030 72.520 -8.680 72.830 ;
        RECT -11.020 72.490 -8.680 72.520 ;
        RECT 37.350 72.710 37.870 72.730 ;
        RECT 61.840 72.710 62.400 72.720 ;
        RECT -13.240 72.410 -12.930 72.420 ;
        RECT -12.150 72.410 -11.840 72.420 ;
        RECT -14.560 72.400 -11.840 72.410 ;
        RECT -14.790 72.090 -11.840 72.400 ;
        RECT -11.020 72.250 -8.640 72.490 ;
        RECT 37.350 72.250 62.490 72.710 ;
        RECT -11.020 72.230 -8.680 72.250 ;
        RECT -14.790 72.080 -11.850 72.090 ;
        RECT -92.400 70.700 -26.950 70.780 ;
        RECT -92.400 69.790 -25.730 70.700 ;
        RECT -92.400 69.410 -17.030 69.790 ;
        RECT -92.400 68.820 -25.730 69.410 ;
        RECT -92.400 68.700 -26.950 68.820 ;
        RECT -96.770 -142.490 -93.980 -138.440 ;
        RECT -96.550 -142.770 -94.470 -142.490 ;
        RECT -92.400 -167.220 -90.320 68.700 ;
        RECT -17.410 68.560 -17.030 69.410 ;
        RECT -14.790 69.640 -14.440 72.080 ;
        RECT -11.020 72.030 -10.420 72.230 ;
        RECT -9.650 72.160 -8.990 72.230 ;
        RECT 37.350 72.200 37.880 72.250 ;
        RECT -9.620 72.150 -9.020 72.160 ;
        RECT 37.350 72.150 37.870 72.200 ;
        RECT -13.790 71.730 -13.480 71.740 ;
        RECT -12.690 71.730 -12.380 71.740 ;
        RECT -11.590 71.730 -11.280 71.740 ;
        RECT -13.820 71.410 -10.660 71.730 ;
        RECT -10.980 70.370 -10.660 71.410 ;
        RECT -13.820 70.040 -10.660 70.370 ;
        RECT -14.790 69.310 -11.840 69.640 ;
        RECT -16.110 68.560 -15.740 68.570 ;
        RECT -14.790 68.560 -14.440 69.310 ;
        RECT -17.410 68.440 -14.440 68.560 ;
        RECT -17.410 68.310 -14.410 68.440 ;
        RECT -17.410 68.270 -14.040 68.310 ;
        RECT -13.240 68.270 -12.930 68.290 ;
        RECT -17.410 68.180 -11.840 68.270 ;
        RECT -16.110 68.160 -15.740 68.180 ;
        RECT -14.790 67.970 -11.840 68.180 ;
        RECT -13.240 67.960 -12.930 67.970 ;
        RECT -12.150 67.940 -11.840 67.970 ;
        RECT -13.790 67.590 -13.480 67.600 ;
        RECT -10.980 67.590 -10.660 70.040 ;
        RECT -6.860 67.590 -6.550 67.610 ;
        RECT -13.810 67.250 -6.550 67.590 ;
        RECT -6.860 67.230 -6.550 67.250 ;
        RECT -25.790 66.640 -25.290 66.750 ;
        RECT 43.180 66.670 43.570 66.680 ;
        RECT 43.170 66.640 43.570 66.670 ;
        RECT -25.790 66.360 43.570 66.640 ;
        RECT -25.790 66.280 -25.290 66.360 ;
        RECT 43.170 66.340 43.570 66.360 ;
        RECT 43.180 66.330 43.570 66.340 ;
        RECT -88.050 65.160 -26.950 65.170 ;
        RECT -88.050 63.280 -25.860 65.160 ;
        RECT -88.050 63.090 -26.950 63.280 ;
        RECT -92.890 -171.000 -90.060 -167.220 ;
        RECT -92.400 -171.560 -90.320 -171.000 ;
        RECT -88.050 -195.800 -85.970 63.090 ;
        RECT -83.890 60.410 -26.950 60.470 ;
        RECT -83.890 58.530 -25.790 60.410 ;
        RECT 76.880 59.980 77.200 60.300 ;
        RECT 77.820 59.980 78.140 60.300 ;
        RECT -83.890 58.390 -26.950 58.530 ;
        RECT -88.400 -199.520 -85.750 -195.800 ;
        RECT -88.050 -199.530 -85.970 -199.520 ;
        RECT -83.890 -224.500 -81.810 58.390 ;
        RECT -84.080 -228.030 -81.410 -224.500 ;
        RECT -22.350 -233.860 -19.010 58.530 ;
        RECT 172.300 -51.510 174.390 79.920 ;
        RECT 176.540 -25.040 178.630 85.430 ;
        RECT 180.670 3.440 182.760 90.470 ;
        RECT 184.760 32.210 186.850 95.670 ;
        RECT 188.840 60.710 190.930 100.550 ;
        RECT 192.980 89.270 195.070 105.950 ;
        RECT 192.780 85.730 195.210 89.270 ;
        RECT 192.980 85.060 195.070 85.730 ;
        RECT 188.600 57.140 191.110 60.710 ;
        RECT 184.560 28.500 187.080 32.210 ;
        RECT 184.760 28.470 186.850 28.500 ;
        RECT 180.400 0.020 182.760 3.440 ;
        RECT 180.670 -0.690 182.760 0.020 ;
        RECT 176.370 -28.750 178.800 -25.040 ;
        RECT 172.310 -53.410 174.390 -51.510 ;
        RECT 172.310 -53.530 174.400 -53.410 ;
        RECT 172.200 -53.590 174.400 -53.530 ;
        RECT 171.940 -57.270 174.470 -53.590 ;
        RECT 172.200 -57.290 174.290 -57.270 ;
      LAYER via2 ;
        RECT 49.580 113.550 49.900 113.870 ;
        RECT 50.610 113.540 50.930 113.860 ;
        RECT 50.690 110.060 51.030 110.400 ;
        RECT 49.620 106.580 49.950 106.930 ;
        RECT 50.710 104.010 51.050 104.370 ;
      LAYER met3 ;
        RECT 49.510 113.180 49.960 113.930 ;
        RECT 49.510 107.020 49.880 113.180 ;
        RECT 50.550 113.170 51.000 113.920 ;
        RECT 50.630 110.530 51.000 113.170 ;
        RECT 50.630 109.930 51.070 110.530 ;
        RECT 49.510 106.690 50.000 107.020 ;
        RECT 49.560 106.530 50.000 106.690 ;
        RECT 50.630 104.820 51.000 109.930 ;
        RECT 50.620 103.950 51.090 104.820 ;
  END
END sky130_hilas_TopProtectStructure

MACRO sky130_hilas_capacitorSize01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_capacitorSize01 ;
  ORIGIN -14.140 0.480 ;
  SIZE 10.420 BY 5.830 ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 23.740 2.130 24.400 2.790 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 14.250 2.720 14.910 2.780 ;
        RECT 15.300 2.720 16.310 2.730 ;
        RECT 14.250 2.220 17.940 2.720 ;
        RECT 14.250 2.210 15.660 2.220 ;
        RECT 14.250 2.120 14.910 2.210 ;
        RECT 17.300 1.100 17.930 2.220 ;
        RECT 17.300 1.090 19.450 1.100 ;
        RECT 16.490 0.620 19.530 1.090 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 14.140 4.800 24.560 4.980 ;
        RECT 14.140 4.370 24.560 4.550 ;
        RECT 14.170 3.370 24.560 3.550 ;
        RECT 22.650 3.120 24.560 3.130 ;
        RECT 14.170 2.940 24.560 3.120 ;
        RECT 14.380 2.600 14.750 2.660 ;
        RECT 14.160 2.320 14.750 2.600 ;
        RECT 14.380 2.260 14.750 2.320 ;
        RECT 23.870 2.610 24.240 2.670 ;
        RECT 23.870 2.330 24.560 2.610 ;
        RECT 23.870 2.270 24.240 2.330 ;
        RECT 14.170 1.790 24.560 1.960 ;
        RECT 14.170 1.370 24.560 1.540 ;
        RECT 14.170 0.390 24.560 0.560 ;
        RECT 14.170 -0.050 24.560 0.120 ;
      LAYER via2 ;
        RECT 14.430 2.320 14.710 2.600 ;
        RECT 23.920 2.330 24.200 2.610 ;
      LAYER met3 ;
        RECT 15.600 5.320 18.420 5.350 ;
        RECT 15.600 2.820 22.800 5.320 ;
        RECT 14.160 2.060 14.950 2.810 ;
        RECT 15.600 2.070 24.440 2.820 ;
        RECT 15.600 -0.460 22.800 2.070 ;
        RECT 18.390 -0.480 22.800 -0.460 ;
      LAYER via3 ;
        RECT 14.350 2.210 14.780 2.690 ;
        RECT 23.840 2.220 24.270 2.700 ;
  END
END sky130_hilas_capacitorSize01

MACRO sky130_hilas_TA2SignalBiasCell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TA2SignalBiasCell ;
  ORIGIN 5.690 -1.400 ;
  SIZE 8.880 BY 6.050 ;
  PIN VOUT_AMP2
    USE ANALOG ;
    ANTENNADIFFAREA 0.308800 ;
    PORT
      LAYER met2 ;
        RECT 0.270 4.970 0.580 5.030 ;
        RECT 2.570 4.970 2.880 4.990 ;
        RECT 0.270 4.740 3.190 4.970 ;
        RECT 0.270 4.700 0.580 4.740 ;
        RECT 2.570 4.660 2.880 4.740 ;
    END
  END VOUT_AMP2
  PIN VOUT_AMP1
    USE ANALOG ;
    ANTENNADIFFAREA 0.308800 ;
    PORT
      LAYER met2 ;
        RECT 0.270 4.140 0.580 4.190 ;
        RECT 2.560 4.140 2.870 4.270 ;
        RECT 0.270 3.920 3.190 4.140 ;
        RECT 0.270 3.860 0.580 3.920 ;
    END
  END VOUT_AMP1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 1.230 1.400 1.570 7.450 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -5.690 7.440 -1.650 7.450 ;
        RECT -5.690 1.410 -0.090 7.440 ;
        RECT -1.950 1.400 -0.090 1.410 ;
        RECT 1.910 1.400 3.190 7.450 ;
      LAYER met2 ;
        RECT -4.900 7.270 -4.660 7.450 ;
        RECT -4.940 6.980 -4.630 7.270 ;
        RECT -5.420 6.940 -4.630 6.980 ;
        RECT -5.420 6.630 -4.660 6.940 ;
        RECT -5.420 6.400 -0.880 6.630 ;
        RECT -5.420 6.160 -4.660 6.400 ;
        RECT -5.420 6.150 -4.970 6.160 ;
        RECT -1.110 6.040 -0.880 6.400 ;
        RECT 1.910 6.040 2.240 6.190 ;
        RECT -1.110 5.840 2.240 6.040 ;
        RECT -0.850 5.830 2.240 5.840 ;
        RECT 1.910 5.260 2.240 5.830 ;
        RECT -4.980 2.780 -4.670 3.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.900 6.190 2.170 7.450 ;
        RECT 1.900 5.260 2.250 6.190 ;
        RECT 1.900 3.280 2.170 5.260 ;
        RECT 1.900 2.990 2.180 3.280 ;
        RECT 1.900 1.400 2.170 2.990 ;
      LAYER via ;
        RECT 1.940 5.290 2.200 6.150 ;
    END
  END VPWR
  PIN VIN22
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -1.300 7.430 -1.050 7.440 ;
        RECT -0.700 7.430 -0.390 7.440 ;
        RECT -1.300 7.180 -0.390 7.430 ;
        RECT -0.700 7.110 -0.390 7.180 ;
    END
  END VIN22
  PIN VIN21
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -0.940 4.750 -0.630 4.790 ;
        RECT -1.030 4.740 -0.600 4.750 ;
        RECT -1.260 4.510 -0.160 4.740 ;
        RECT -0.940 4.460 -0.630 4.510 ;
    END
  END VIN21
  PIN VIN11
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -2.500 4.340 -2.190 4.390 ;
        RECT -2.820 4.110 -1.720 4.340 ;
        RECT -2.820 4.100 -2.160 4.110 ;
        RECT -2.500 4.060 -2.190 4.100 ;
    END
  END VIN11
  PIN VIN12
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -2.260 1.670 -1.950 1.740 ;
        RECT -2.860 1.420 -1.950 1.670 ;
        RECT -2.260 1.410 -1.950 1.420 ;
    END
  END VIN12
  PIN VBIAS2
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -4.010 1.670 -3.700 1.740 ;
        RECT -4.580 1.660 -3.700 1.670 ;
        RECT -5.640 1.430 -3.700 1.660 ;
        RECT -4.580 1.420 -3.700 1.430 ;
        RECT -4.010 1.410 -3.700 1.420 ;
    END
  END VBIAS2
  PIN VBIAS1
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -4.250 4.340 -3.940 4.390 ;
        RECT -5.680 4.110 -3.470 4.340 ;
        RECT -5.680 4.100 -3.910 4.110 ;
        RECT -5.680 4.090 -5.040 4.100 ;
        RECT -4.250 4.060 -3.940 4.100 ;
    END
  END VBIAS1
  OBS
      LAYER li1 ;
        RECT -0.960 7.400 -0.790 7.450 ;
        RECT -4.930 7.190 -4.610 7.230 ;
        RECT -4.930 7.000 -4.600 7.190 ;
        RECT -0.960 7.140 -0.400 7.400 ;
        RECT 0.510 7.150 0.710 7.190 ;
        RECT -0.960 7.120 -0.790 7.140 ;
        RECT -4.930 6.980 -4.610 7.000 ;
        RECT -5.020 6.970 -4.610 6.980 ;
        RECT -5.270 6.780 -4.670 6.970 ;
        RECT -5.440 6.240 -4.670 6.780 ;
        RECT -5.440 4.910 -5.270 6.240 ;
        RECT -5.430 1.970 -5.260 3.750 ;
        RECT -4.850 3.070 -4.670 6.240 ;
        RECT -4.040 5.950 -3.870 6.970 ;
        RECT -4.090 5.910 -3.770 5.950 ;
        RECT -4.090 5.720 -3.760 5.910 ;
        RECT -4.090 5.690 -3.770 5.720 ;
        RECT -4.040 5.190 -3.870 5.690 ;
        RECT -4.120 5.130 -3.580 5.190 ;
        RECT -4.120 5.020 -3.570 5.130 ;
        RECT -3.760 4.900 -3.570 5.020 ;
        RECT -4.290 4.600 -4.120 4.760 ;
        RECT -4.290 4.430 -4.070 4.600 ;
        RECT -4.240 4.350 -4.070 4.430 ;
        RECT -4.240 4.310 -3.920 4.350 ;
        RECT -4.240 4.120 -3.910 4.310 ;
        RECT -4.240 4.090 -3.920 4.120 ;
        RECT -4.970 3.030 -4.650 3.070 ;
        RECT -4.970 2.840 -4.640 3.030 ;
        RECT -4.970 2.810 -4.650 2.840 ;
        RECT -4.850 1.880 -4.670 2.810 ;
        RECT -4.040 2.540 -3.870 3.920 ;
        RECT -3.100 3.070 -2.920 6.980 ;
        RECT -2.290 5.190 -2.120 6.970 ;
        RECT -1.540 6.040 -1.360 6.970 ;
        RECT 0.280 6.890 0.710 7.150 ;
        RECT -0.810 6.710 -0.480 6.880 ;
        RECT 0.510 6.860 0.710 6.890 ;
        RECT -0.730 6.570 -0.480 6.710 ;
        RECT -0.730 6.310 -0.250 6.570 ;
        RECT 0.100 6.500 0.270 6.540 ;
        RECT 0.510 6.500 0.710 6.530 ;
        RECT -1.660 6.010 -1.340 6.040 ;
        RECT -1.660 5.820 -1.330 6.010 ;
        RECT -1.660 5.780 -1.340 5.820 ;
        RECT -2.370 5.130 -1.830 5.190 ;
        RECT -2.370 5.020 -1.820 5.130 ;
        RECT -2.010 4.900 -1.820 5.020 ;
        RECT -2.540 4.600 -2.370 4.760 ;
        RECT -2.540 4.430 -2.320 4.600 ;
        RECT -2.490 4.350 -2.320 4.430 ;
        RECT -2.490 4.310 -2.170 4.350 ;
        RECT -2.490 4.120 -2.160 4.310 ;
        RECT -2.490 4.090 -2.170 4.120 ;
        RECT -3.220 3.030 -2.900 3.070 ;
        RECT -3.220 2.840 -2.890 3.030 ;
        RECT -3.220 2.810 -2.900 2.840 ;
        RECT -4.040 2.280 -3.560 2.540 ;
        RECT -4.040 2.140 -3.790 2.280 ;
        RECT -4.120 1.970 -3.790 2.140 ;
        RECT -3.100 1.880 -2.920 2.810 ;
        RECT -2.290 2.540 -2.120 3.920 ;
        RECT -2.290 2.280 -1.810 2.540 ;
        RECT -2.290 2.140 -2.040 2.280 ;
        RECT -2.370 1.970 -2.040 2.140 ;
        RECT -1.540 1.870 -1.360 5.780 ;
        RECT -0.730 4.930 -0.560 6.310 ;
        RECT 0.100 6.240 0.710 6.500 ;
        RECT 0.100 6.210 0.270 6.240 ;
        RECT 0.510 6.200 0.710 6.240 ;
        RECT 1.100 6.200 1.650 7.190 ;
        RECT 2.470 7.040 3.100 7.210 ;
        RECT 2.470 6.940 2.860 7.040 ;
        RECT 2.470 6.910 2.850 6.940 ;
        RECT 2.470 6.760 2.830 6.910 ;
        RECT 2.120 6.590 2.830 6.760 ;
        RECT 0.100 5.650 0.270 5.680 ;
        RECT 0.510 5.650 0.710 5.690 ;
        RECT 0.100 5.390 0.710 5.650 ;
        RECT 0.100 5.350 0.270 5.390 ;
        RECT 0.510 5.360 0.710 5.390 ;
        RECT 0.510 5.000 0.710 5.030 ;
        RECT -0.930 4.730 -0.610 4.760 ;
        RECT 0.280 4.740 0.710 5.000 ;
        RECT -0.930 4.540 -0.600 4.730 ;
        RECT 0.510 4.700 0.710 4.740 ;
        RECT 1.100 4.700 1.650 5.690 ;
        RECT 1.960 5.270 2.820 6.150 ;
        RECT 1.960 5.260 2.170 5.270 ;
        RECT 2.580 4.910 2.900 4.950 ;
        RECT 2.580 4.850 2.910 4.910 ;
        RECT 2.110 4.720 2.910 4.850 ;
        RECT 2.110 4.690 2.900 4.720 ;
        RECT 2.110 4.670 2.810 4.690 ;
        RECT -0.930 4.500 -0.610 4.540 ;
        RECT -0.930 4.420 -0.760 4.500 ;
        RECT -0.980 4.250 -0.760 4.420 ;
        RECT -0.980 4.090 -0.810 4.250 ;
        RECT 2.570 4.190 2.890 4.230 ;
        RECT 0.510 4.150 0.710 4.190 ;
        RECT -0.450 3.830 -0.260 3.950 ;
        RECT 0.280 3.890 0.710 4.150 ;
        RECT 0.510 3.860 0.710 3.890 ;
        RECT -0.810 3.720 -0.260 3.830 ;
        RECT -0.810 3.660 -0.270 3.720 ;
        RECT -0.730 1.880 -0.560 3.660 ;
        RECT 0.100 3.500 0.270 3.540 ;
        RECT 0.510 3.500 0.710 3.530 ;
        RECT 0.100 3.240 0.710 3.500 ;
        RECT 0.100 3.210 0.270 3.240 ;
        RECT 0.510 3.200 0.710 3.240 ;
        RECT 1.100 3.200 1.650 4.190 ;
        RECT 2.110 4.010 2.900 4.190 ;
        RECT 2.570 4.000 2.900 4.010 ;
        RECT 2.570 3.970 2.890 4.000 ;
        RECT 2.120 3.250 2.820 3.590 ;
        RECT 1.970 3.020 2.820 3.250 ;
        RECT 2.120 2.710 2.820 3.020 ;
        RECT 0.100 2.650 0.270 2.680 ;
        RECT 0.510 2.650 0.710 2.690 ;
        RECT 0.100 2.390 0.710 2.650 ;
        RECT 0.100 2.350 0.270 2.390 ;
        RECT 0.510 2.360 0.710 2.390 ;
        RECT 0.510 2.000 0.710 2.030 ;
        RECT 0.280 1.740 0.710 2.000 ;
        RECT -4.270 1.710 -4.100 1.730 ;
        RECT -2.520 1.710 -2.350 1.730 ;
        RECT -4.270 1.450 -3.710 1.710 ;
        RECT -2.520 1.450 -1.960 1.710 ;
        RECT 0.510 1.700 0.710 1.740 ;
        RECT 1.100 1.700 1.650 2.690 ;
        RECT 2.120 2.100 2.830 2.270 ;
        RECT 2.470 1.820 2.830 2.100 ;
        RECT 2.470 1.650 3.100 1.820 ;
        RECT -4.270 1.400 -4.100 1.450 ;
        RECT -2.520 1.400 -2.350 1.450 ;
      LAYER mcon ;
        RECT -4.870 7.010 -4.700 7.180 ;
        RECT -0.630 7.180 -0.460 7.350 ;
        RECT -5.440 6.610 -5.270 6.780 ;
        RECT -4.850 6.560 -4.680 6.730 ;
        RECT -5.440 6.270 -5.270 6.440 ;
        RECT -5.440 5.930 -5.270 6.100 ;
        RECT -5.440 5.590 -5.270 5.760 ;
        RECT -5.440 5.250 -5.270 5.420 ;
        RECT -4.850 6.220 -4.680 6.390 ;
        RECT -5.430 3.580 -5.260 3.750 ;
        RECT -5.430 3.240 -5.260 3.410 ;
        RECT -4.030 5.730 -3.860 5.900 ;
        RECT -3.750 4.930 -3.580 5.100 ;
        RECT -4.180 4.130 -4.010 4.300 ;
        RECT -5.430 2.900 -5.260 3.070 ;
        RECT -4.910 2.850 -4.740 3.020 ;
        RECT -5.430 2.560 -5.260 2.730 ;
        RECT -5.430 2.220 -5.260 2.390 ;
        RECT 0.340 6.930 0.510 7.100 ;
        RECT 1.320 6.610 1.490 6.780 ;
        RECT 2.590 6.950 2.760 7.120 ;
        RECT -0.480 6.350 -0.310 6.520 ;
        RECT -1.600 5.830 -1.430 6.000 ;
        RECT -2.000 4.930 -1.830 5.100 ;
        RECT -2.430 4.130 -2.260 4.300 ;
        RECT -3.160 2.850 -2.990 3.020 ;
        RECT -3.790 2.330 -3.620 2.500 ;
        RECT -2.040 2.330 -1.870 2.500 ;
        RECT 0.290 6.280 0.460 6.450 ;
        RECT 1.980 5.980 2.150 6.150 ;
        RECT 0.290 5.440 0.460 5.610 ;
        RECT 1.320 5.110 1.490 5.280 ;
        RECT 1.980 5.640 2.150 5.810 ;
        RECT 1.980 5.280 2.150 5.450 ;
        RECT 0.340 4.790 0.510 4.960 ;
        RECT -0.870 4.550 -0.700 4.720 ;
        RECT 2.640 4.730 2.810 4.900 ;
        RECT -0.440 3.750 -0.270 3.920 ;
        RECT 0.340 3.930 0.510 4.100 ;
        RECT 2.630 4.010 2.800 4.180 ;
        RECT 1.320 3.610 1.490 3.780 ;
        RECT 0.290 3.280 0.460 3.450 ;
        RECT 1.980 3.050 2.150 3.220 ;
        RECT 0.290 2.440 0.460 2.610 ;
        RECT 1.320 2.110 1.490 2.280 ;
        RECT 0.340 1.790 0.510 1.960 ;
        RECT -3.940 1.500 -3.770 1.670 ;
        RECT 2.550 1.760 2.720 1.930 ;
        RECT -2.190 1.500 -2.020 1.670 ;
      LAYER met1 ;
        RECT -4.940 6.990 -4.620 7.260 ;
        RECT -0.710 7.110 -0.390 7.430 ;
        RECT -5.470 6.940 -4.620 6.990 ;
        RECT -5.470 6.670 -4.650 6.940 ;
        RECT 0.270 6.860 0.590 7.180 ;
        RECT 2.520 6.880 2.840 7.200 ;
        RECT -5.470 6.380 -4.620 6.670 ;
        RECT -5.470 6.130 -4.650 6.380 ;
        RECT -0.560 6.280 -0.240 6.600 ;
        RECT 0.220 6.210 0.540 6.530 ;
        RECT -5.470 3.100 -4.830 6.130 ;
        RECT -4.100 5.660 -3.780 5.980 ;
        RECT -1.670 5.750 -1.350 6.070 ;
        RECT -0.450 5.590 -0.240 5.700 ;
        RECT -0.470 5.270 -0.210 5.590 ;
        RECT 0.220 5.360 0.540 5.680 ;
        RECT -3.780 4.870 -3.550 5.160 ;
        RECT -2.030 4.870 -1.800 5.160 ;
        RECT -4.250 4.060 -3.930 4.380 ;
        RECT -3.760 3.580 -3.550 4.870 ;
        RECT -2.500 4.060 -2.180 4.380 ;
        RECT -2.010 3.580 -1.800 4.870 ;
        RECT -0.940 4.470 -0.620 4.790 ;
        RECT -0.450 3.980 -0.240 5.270 ;
        RECT 0.270 4.710 0.590 5.030 ;
        RECT 2.570 4.660 2.890 4.980 ;
        RECT -0.470 3.690 -0.240 3.980 ;
        RECT 0.270 3.860 0.590 4.180 ;
        RECT 2.560 3.940 2.880 4.260 ;
        RECT -3.780 3.260 -3.520 3.580 ;
        RECT -2.030 3.260 -1.770 3.580 ;
        RECT -3.760 3.150 -3.550 3.260 ;
        RECT -2.010 3.150 -1.800 3.260 ;
        RECT 0.220 3.210 0.540 3.530 ;
        RECT -5.470 2.780 -4.660 3.100 ;
        RECT -3.230 2.780 -2.910 3.100 ;
        RECT -5.470 1.950 -4.830 2.780 ;
        RECT -3.870 2.250 -3.550 2.570 ;
        RECT -2.120 2.250 -1.800 2.570 ;
        RECT 0.220 2.360 0.540 2.680 ;
        RECT -5.250 1.940 -4.830 1.950 ;
        RECT -4.020 1.420 -3.700 1.740 ;
        RECT -2.270 1.420 -1.950 1.740 ;
        RECT 0.270 1.710 0.590 2.030 ;
        RECT 2.480 1.690 2.800 2.010 ;
      LAYER via ;
        RECT -4.910 6.970 -4.650 7.230 ;
        RECT -0.680 7.140 -0.420 7.400 ;
        RECT -5.350 6.190 -4.760 6.910 ;
        RECT 0.300 6.890 0.560 7.150 ;
        RECT 2.550 6.910 2.810 7.170 ;
        RECT -0.530 6.310 -0.270 6.570 ;
        RECT 0.250 6.240 0.510 6.500 ;
        RECT -4.070 5.690 -3.810 5.950 ;
        RECT -1.640 5.780 -1.380 6.040 ;
        RECT -0.470 5.300 -0.210 5.560 ;
        RECT 0.250 5.390 0.510 5.650 ;
        RECT -4.220 4.090 -3.960 4.350 ;
        RECT -2.470 4.090 -2.210 4.350 ;
        RECT -0.910 4.500 -0.650 4.760 ;
        RECT 0.300 4.740 0.560 5.000 ;
        RECT 2.600 4.690 2.860 4.950 ;
        RECT 0.300 3.890 0.560 4.150 ;
        RECT 2.590 3.970 2.850 4.230 ;
        RECT -3.780 3.290 -3.520 3.550 ;
        RECT -2.030 3.290 -1.770 3.550 ;
        RECT 0.250 3.240 0.510 3.500 ;
        RECT -4.950 2.810 -4.690 3.070 ;
        RECT -3.200 2.810 -2.940 3.070 ;
        RECT -3.840 2.280 -3.580 2.540 ;
        RECT -2.090 2.280 -1.830 2.540 ;
        RECT 0.250 2.390 0.510 2.650 ;
        RECT 0.300 1.740 0.560 2.000 ;
        RECT -3.990 1.450 -3.730 1.710 ;
        RECT 2.510 1.720 2.770 1.980 ;
        RECT -2.240 1.450 -1.980 1.710 ;
      LAYER met2 ;
        RECT 0.270 7.110 0.580 7.190 ;
        RECT 2.520 7.110 2.830 7.210 ;
        RECT 0.270 6.880 2.830 7.110 ;
        RECT 0.270 6.860 0.580 6.880 ;
        RECT -0.550 6.570 -0.240 6.610 ;
        RECT -0.730 6.460 0.010 6.570 ;
        RECT 0.220 6.460 0.530 6.540 ;
        RECT -0.730 6.320 0.530 6.460 ;
        RECT -0.550 6.280 0.530 6.320 ;
        RECT -0.240 6.250 0.530 6.280 ;
        RECT -0.240 6.200 0.010 6.250 ;
        RECT 0.220 6.210 0.530 6.250 ;
        RECT -4.100 5.930 -3.790 5.990 ;
        RECT -1.670 5.930 -1.360 6.070 ;
        RECT -4.100 5.740 -1.360 5.930 ;
        RECT -4.100 5.710 -1.620 5.740 ;
        RECT -4.100 5.660 -3.790 5.710 ;
        RECT 0.220 5.640 0.530 5.680 ;
        RECT -0.210 5.560 0.530 5.640 ;
        RECT -0.500 5.540 0.530 5.560 ;
        RECT -0.550 5.430 0.530 5.540 ;
        RECT -0.550 5.350 0.000 5.430 ;
        RECT 0.220 5.350 0.530 5.430 ;
        RECT -0.550 5.290 -0.080 5.350 ;
        RECT -3.860 3.310 -3.390 3.560 ;
        RECT -2.110 3.470 -1.640 3.560 ;
        RECT -2.110 3.460 0.000 3.470 ;
        RECT 0.220 3.460 0.530 3.540 ;
        RECT -2.110 3.310 0.530 3.460 ;
        RECT -3.810 3.290 -3.490 3.310 ;
        RECT -2.060 3.290 0.530 3.310 ;
        RECT -1.770 3.270 0.530 3.290 ;
        RECT -0.080 3.250 0.530 3.270 ;
        RECT 0.220 3.210 0.530 3.250 ;
        RECT -3.230 3.100 -2.920 3.110 ;
        RECT -3.340 2.920 -2.920 3.100 ;
        RECT -3.360 2.910 -2.920 2.920 ;
        RECT -3.580 2.780 -2.920 2.910 ;
        RECT -3.580 2.570 -3.220 2.780 ;
        RECT -2.060 2.640 0.000 2.670 ;
        RECT 0.220 2.640 0.530 2.680 ;
        RECT -2.060 2.570 0.530 2.640 ;
        RECT -3.860 2.530 -3.220 2.570 ;
        RECT -2.110 2.530 0.530 2.570 ;
        RECT -4.040 2.290 -3.220 2.530 ;
        RECT -2.290 2.460 0.530 2.530 ;
        RECT -4.040 2.280 -3.490 2.290 ;
        RECT -2.290 2.280 -1.740 2.460 ;
        RECT -0.080 2.430 0.530 2.460 ;
        RECT 0.220 2.350 0.530 2.430 ;
        RECT -3.860 2.240 -3.550 2.280 ;
        RECT -2.110 2.240 -1.800 2.280 ;
        RECT 0.270 1.980 0.580 2.030 ;
        RECT 2.480 1.980 2.790 2.020 ;
        RECT 0.270 1.750 2.980 1.980 ;
        RECT 0.270 1.700 0.580 1.750 ;
        RECT 2.480 1.690 2.790 1.750 ;
  END
END sky130_hilas_TA2SignalBiasCell

MACRO sky130_hilas_StepUpDigital
  CLASS BLOCK ;
  FOREIGN sky130_hilas_StepUpDigital ;
  ORIGIN -0.190 0.440 ;
  SIZE 8.700 BY 1.750 ;
  OBS
      LAYER nwell ;
        RECT 0.190 -0.440 2.690 1.310 ;
        RECT 6.560 -0.440 8.330 1.310 ;
      LAYER li1 ;
        RECT 1.470 0.800 1.920 0.950 ;
        RECT 0.530 0.620 0.860 0.790 ;
        RECT 1.320 0.630 1.920 0.800 ;
        RECT 0.600 0.160 0.780 0.620 ;
        RECT 2.120 0.190 2.290 0.950 ;
        RECT 2.620 0.860 2.910 0.880 ;
        RECT 2.620 0.820 3.080 0.860 ;
        RECT 2.620 0.800 4.060 0.820 ;
        RECT 2.620 0.640 4.100 0.800 ;
        RECT 2.910 0.630 4.100 0.640 ;
        RECT 4.550 0.770 5.010 0.800 ;
        RECT 6.320 0.770 6.670 0.870 ;
        RECT 4.550 0.630 5.660 0.770 ;
        RECT 4.840 0.600 5.660 0.630 ;
        RECT 5.900 0.600 7.070 0.770 ;
        RECT 7.320 0.600 8.080 0.770 ;
        RECT 4.840 0.460 5.100 0.600 ;
        RECT 3.920 0.290 5.100 0.460 ;
        RECT 7.850 0.590 8.080 0.600 ;
        RECT 2.120 0.180 2.500 0.190 ;
        RECT 0.600 -0.010 1.560 0.160 ;
        RECT 2.030 0.120 2.500 0.180 ;
        RECT 2.030 0.010 3.370 0.120 ;
        RECT 2.110 -0.050 3.370 0.010 ;
        RECT 2.110 -0.100 2.500 -0.050 ;
        RECT 3.920 -0.150 4.100 0.290 ;
        RECT 4.840 0.150 5.100 0.290 ;
        RECT 6.310 0.150 6.640 0.410 ;
        RECT 7.850 0.150 8.120 0.590 ;
        RECT 4.340 -0.210 4.550 0.120 ;
        RECT 4.840 -0.020 5.170 0.150 ;
        RECT 5.410 -0.020 7.570 0.150 ;
        RECT 4.840 -0.070 5.010 -0.020 ;
        RECT 7.820 -0.030 8.150 0.150 ;
        RECT 8.500 0.010 8.670 0.070 ;
        RECT 8.480 -0.210 8.700 0.010 ;
        RECT 8.500 -0.260 8.670 -0.210 ;
      LAYER mcon ;
        RECT 1.640 0.700 1.810 0.870 ;
        RECT 0.600 0.360 0.770 0.530 ;
        RECT 2.680 0.660 2.850 0.830 ;
        RECT 6.380 0.640 6.590 0.850 ;
        RECT 0.600 0.000 0.770 0.170 ;
        RECT 7.890 0.270 8.060 0.440 ;
      LAYER met1 ;
        RECT 0.530 -0.440 0.820 1.310 ;
        RECT 1.570 0.650 1.890 0.950 ;
        RECT 2.620 0.880 2.930 0.890 ;
        RECT 2.610 0.610 2.930 0.880 ;
        RECT 2.620 0.600 2.910 0.610 ;
        RECT 4.310 -0.150 4.590 0.180 ;
        RECT 4.840 -0.440 5.150 1.310 ;
        RECT 6.320 0.600 6.670 0.890 ;
        RECT 6.470 0.580 6.670 0.600 ;
        RECT 7.850 -0.440 8.090 1.310 ;
        RECT 8.420 -0.260 8.830 0.070 ;
      LAYER via ;
        RECT 1.600 0.660 1.860 0.920 ;
        RECT 2.640 0.620 2.900 0.880 ;
        RECT 4.320 -0.110 4.580 0.150 ;
        RECT 6.360 0.610 6.620 0.870 ;
        RECT 8.460 -0.230 8.720 0.030 ;
      LAYER met2 ;
        RECT 1.570 0.870 1.890 0.920 ;
        RECT 2.600 0.880 2.920 0.890 ;
        RECT 2.600 0.870 2.930 0.880 ;
        RECT 0.260 0.670 2.930 0.870 ;
        RECT 1.570 0.660 1.890 0.670 ;
        RECT 2.600 0.620 2.930 0.670 ;
        RECT 2.600 0.600 2.920 0.620 ;
        RECT 4.280 0.100 4.620 0.160 ;
        RECT 6.360 0.100 6.620 0.900 ;
        RECT 4.280 -0.120 6.720 0.100 ;
        RECT 8.430 -0.260 8.890 0.060 ;
  END
END sky130_hilas_StepUpDigital

MACRO sky130_hilas_Tgate4Double01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_Tgate4Double01 ;
  ORIGIN 0.360 1.410 ;
  SIZE 7.080 BY 6.050 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER nwell ;
        RECT -0.240 -1.410 3.230 4.640 ;
      LAYER met1 ;
        RECT 0.380 3.770 0.580 4.640 ;
        RECT 0.370 3.480 0.600 3.770 ;
        RECT 0.380 2.770 0.580 3.480 ;
        RECT 0.370 2.480 0.600 2.770 ;
        RECT 0.380 0.750 0.580 2.480 ;
        RECT 0.370 0.460 0.600 0.750 ;
        RECT 0.380 -0.250 0.580 0.460 ;
        RECT 0.370 -0.540 0.600 -0.250 ;
        RECT 0.380 -1.410 0.580 -0.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.210 3.770 6.400 4.640 ;
        RECT 6.190 3.480 6.420 3.770 ;
        RECT 6.210 2.770 6.400 3.480 ;
        RECT 6.190 2.480 6.420 2.770 ;
        RECT 6.210 0.750 6.400 2.480 ;
        RECT 6.190 0.460 6.420 0.750 ;
        RECT 6.210 -0.250 6.400 0.460 ;
        RECT 6.190 -0.540 6.420 -0.250 ;
        RECT 6.210 -1.410 6.400 -0.540 ;
    END
  END VGND
  PIN INPUT1_1
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.090 4.530 2.400 4.540 ;
        RECT -0.360 4.330 5.480 4.530 ;
        RECT 2.090 4.210 2.400 4.330 ;
        RECT 5.170 4.200 5.480 4.330 ;
    END
  END INPUT1_1
  PIN SELECT1
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER met2 ;
        RECT -0.360 3.350 0.250 3.550 ;
        RECT -0.070 3.260 0.250 3.350 ;
    END
  END SELECT1
  PIN SELECT2
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER met2 ;
        RECT -0.070 2.900 0.250 2.990 ;
        RECT -0.360 2.700 0.250 2.900 ;
    END
  END SELECT2
  PIN INPUT2_2
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 0.740 2.400 1.050 2.410 ;
        RECT 3.660 2.400 3.970 2.410 ;
        RECT -0.360 2.200 4.010 2.400 ;
        RECT 0.740 2.080 1.050 2.200 ;
        RECT 3.660 2.080 3.970 2.200 ;
    END
  END INPUT2_2
  PIN INPUT1_2
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.090 1.920 2.400 2.040 ;
        RECT 5.170 1.920 5.480 2.050 ;
        RECT -0.360 1.720 5.480 1.920 ;
        RECT 2.090 1.710 2.400 1.720 ;
    END
  END INPUT1_2
  PIN SELECT3
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER met2 ;
        RECT -0.360 0.330 0.250 0.530 ;
        RECT -0.070 0.240 0.250 0.330 ;
    END
  END SELECT3
  PIN INPUT2_3
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 0.740 1.030 1.050 1.150 ;
        RECT 3.660 1.030 3.970 1.150 ;
        RECT -0.360 0.830 4.010 1.030 ;
        RECT 0.740 0.820 1.050 0.830 ;
        RECT 3.660 0.820 3.970 0.830 ;
    END
  END INPUT2_3
  PIN SELECT4
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER met2 ;
        RECT -0.070 -0.120 0.250 -0.030 ;
        RECT -0.360 -0.320 0.250 -0.120 ;
    END
  END SELECT4
  PIN INPUT2_4
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 0.740 -0.620 1.050 -0.610 ;
        RECT 3.660 -0.620 3.970 -0.610 ;
        RECT -0.360 -0.820 4.010 -0.620 ;
        RECT 0.740 -0.940 1.050 -0.820 ;
        RECT 3.660 -0.940 3.970 -0.820 ;
    END
  END INPUT2_4
  PIN INPUT1_4
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.090 -1.100 2.400 -0.980 ;
        RECT 5.170 -1.100 5.480 -0.970 ;
        RECT -0.360 -1.300 5.480 -1.100 ;
        RECT 2.090 -1.310 2.400 -1.300 ;
    END
  END INPUT1_4
  PIN OUTPUT4
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER met2 ;
        RECT 1.320 -0.120 1.640 -0.110 ;
        RECT 2.740 -0.120 3.060 -0.100 ;
        RECT 4.490 -0.120 4.810 -0.080 ;
        RECT 5.530 -0.120 5.850 -0.090 ;
        RECT 1.320 -0.320 6.720 -0.120 ;
        RECT 1.320 -0.370 1.640 -0.320 ;
        RECT 2.740 -0.360 3.060 -0.320 ;
        RECT 4.490 -0.340 4.810 -0.320 ;
        RECT 5.530 -0.350 5.850 -0.320 ;
    END
  END OUTPUT4
  PIN OUTPUT3
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER met2 ;
        RECT 1.320 0.530 1.640 0.580 ;
        RECT 2.740 0.530 3.060 0.570 ;
        RECT 4.490 0.530 4.810 0.550 ;
        RECT 5.530 0.530 5.850 0.560 ;
        RECT 1.320 0.330 6.720 0.530 ;
        RECT 1.320 0.320 1.640 0.330 ;
        RECT 2.740 0.310 3.060 0.330 ;
        RECT 4.490 0.290 4.810 0.330 ;
        RECT 5.530 0.300 5.850 0.330 ;
    END
  END OUTPUT3
  PIN OUTPUT2
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER met2 ;
        RECT 1.320 2.900 1.640 2.910 ;
        RECT 2.740 2.900 3.060 2.920 ;
        RECT 4.490 2.900 4.810 2.940 ;
        RECT 5.530 2.900 5.850 2.930 ;
        RECT 1.320 2.700 6.720 2.900 ;
        RECT 1.320 2.650 1.640 2.700 ;
        RECT 2.740 2.660 3.060 2.700 ;
        RECT 4.490 2.680 4.810 2.700 ;
        RECT 5.530 2.670 5.850 2.700 ;
    END
  END OUTPUT2
  PIN OUTPUT1
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER met2 ;
        RECT 1.320 3.550 1.640 3.600 ;
        RECT 2.740 3.550 3.060 3.590 ;
        RECT 4.490 3.550 4.810 3.570 ;
        RECT 5.530 3.550 5.850 3.580 ;
        RECT 1.320 3.350 6.720 3.550 ;
        RECT 1.320 3.340 1.640 3.350 ;
        RECT 2.740 3.330 3.060 3.350 ;
        RECT 4.490 3.310 4.810 3.350 ;
        RECT 5.530 3.320 5.850 3.350 ;
    END
  END OUTPUT1
  PIN INPUT2_1
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 0.740 4.050 1.050 4.170 ;
        RECT 3.660 4.050 3.970 4.170 ;
        RECT -0.360 3.850 4.010 4.050 ;
        RECT 0.740 3.840 1.050 3.850 ;
        RECT 3.660 3.840 3.970 3.850 ;
    END
  END INPUT2_1
  PIN INPUT1_3
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.090 1.510 2.400 1.520 ;
        RECT -0.360 1.310 5.480 1.510 ;
        RECT 2.090 1.190 2.400 1.310 ;
        RECT 5.170 1.180 5.480 1.310 ;
    END
  END INPUT1_3
  OBS
      LAYER li1 ;
        RECT 2.100 4.480 2.420 4.510 ;
        RECT 0.070 4.130 0.240 4.410 ;
        RECT 0.580 4.170 0.930 4.340 ;
        RECT 0.750 4.140 0.930 4.170 ;
        RECT 1.350 4.150 1.520 4.420 ;
        RECT 2.100 4.290 2.430 4.480 ;
        RECT 5.180 4.470 5.500 4.500 ;
        RECT 2.100 4.250 2.420 4.290 ;
        RECT 0.070 4.090 0.280 4.130 ;
        RECT 0.750 4.110 1.070 4.140 ;
        RECT 0.070 4.070 0.300 4.090 ;
        RECT 0.070 4.050 0.330 4.070 ;
        RECT 0.070 4.000 0.410 4.050 ;
        RECT 0.070 3.940 0.560 4.000 ;
        RECT 0.070 3.910 0.580 3.940 ;
        RECT 0.110 3.880 0.580 3.910 ;
        RECT 0.750 3.920 1.080 4.110 ;
        RECT 1.350 3.930 1.550 4.150 ;
        RECT 2.130 4.080 2.300 4.250 ;
        RECT 2.820 4.130 2.990 4.420 ;
        RECT 3.780 4.140 3.950 4.420 ;
        RECT 4.520 4.140 4.690 4.430 ;
        RECT 5.180 4.280 5.510 4.470 ;
        RECT 5.750 4.330 5.940 4.360 ;
        RECT 5.180 4.240 5.500 4.280 ;
        RECT 1.360 3.920 1.550 3.930 ;
        RECT 0.750 3.880 1.070 3.920 ;
        RECT 2.810 3.900 3.000 4.130 ;
        RECT 3.670 4.110 3.990 4.140 ;
        RECT 3.670 3.920 4.000 4.110 ;
        RECT 3.670 3.880 3.990 3.920 ;
        RECT 4.520 3.910 4.710 4.140 ;
        RECT 5.240 4.080 5.410 4.240 ;
        RECT 5.750 4.160 6.190 4.330 ;
        RECT 5.750 4.130 5.940 4.160 ;
        RECT 0.240 3.830 0.580 3.880 ;
        RECT 0.360 3.820 0.580 3.830 ;
        RECT 0.370 3.790 0.580 3.820 ;
        RECT 0.390 3.710 0.580 3.790 ;
        RECT 1.750 3.710 2.080 3.830 ;
        RECT 6.470 3.740 6.640 4.420 ;
        RECT -0.100 3.660 0.070 3.680 ;
        RECT -0.120 3.230 0.090 3.660 ;
        RECT 0.390 3.540 0.910 3.710 ;
        RECT 0.390 3.510 0.580 3.540 ;
        RECT 1.260 3.530 5.480 3.710 ;
        RECT 6.210 3.700 6.640 3.740 ;
        RECT 5.860 3.540 6.640 3.700 ;
        RECT 5.860 3.530 6.400 3.540 ;
        RECT 6.210 3.510 6.400 3.530 ;
        RECT -0.120 2.590 0.090 3.020 ;
        RECT 0.390 2.710 0.580 2.740 ;
        RECT 6.210 2.720 6.400 2.740 ;
        RECT -0.100 2.570 0.070 2.590 ;
        RECT 0.390 2.540 0.910 2.710 ;
        RECT 1.260 2.540 5.480 2.720 ;
        RECT 5.860 2.710 6.400 2.720 ;
        RECT 5.860 2.550 6.640 2.710 ;
        RECT 0.390 2.460 0.580 2.540 ;
        RECT 0.370 2.430 0.580 2.460 ;
        RECT 0.360 2.420 0.580 2.430 ;
        RECT 1.750 2.420 2.080 2.540 ;
        RECT 6.210 2.510 6.640 2.550 ;
        RECT 0.240 2.370 0.580 2.420 ;
        RECT 0.110 2.340 0.580 2.370 ;
        RECT 0.070 2.310 0.580 2.340 ;
        RECT 0.750 2.330 1.070 2.370 ;
        RECT 0.070 2.250 0.560 2.310 ;
        RECT 0.070 2.200 0.410 2.250 ;
        RECT 0.070 2.180 0.330 2.200 ;
        RECT 0.070 2.160 0.300 2.180 ;
        RECT 0.070 2.120 0.280 2.160 ;
        RECT 0.750 2.140 1.080 2.330 ;
        RECT 1.360 2.320 1.550 2.330 ;
        RECT 0.070 1.840 0.240 2.120 ;
        RECT 0.750 2.110 1.070 2.140 ;
        RECT 0.750 2.080 0.930 2.110 ;
        RECT 0.580 1.910 0.930 2.080 ;
        RECT 1.350 2.100 1.550 2.320 ;
        RECT 1.350 1.830 1.520 2.100 ;
        RECT 2.130 2.000 2.300 2.170 ;
        RECT 2.810 2.120 3.000 2.350 ;
        RECT 3.670 2.330 3.990 2.370 ;
        RECT 3.670 2.140 4.000 2.330 ;
        RECT 2.100 1.960 2.420 2.000 ;
        RECT 2.100 1.770 2.430 1.960 ;
        RECT 2.820 1.830 2.990 2.120 ;
        RECT 3.670 2.110 3.990 2.140 ;
        RECT 4.520 2.110 4.710 2.340 ;
        RECT 3.780 1.830 3.950 2.110 ;
        RECT 4.520 1.820 4.690 2.110 ;
        RECT 5.240 2.010 5.410 2.170 ;
        RECT 5.750 2.090 5.940 2.120 ;
        RECT 5.180 1.970 5.500 2.010 ;
        RECT 5.180 1.780 5.510 1.970 ;
        RECT 5.750 1.920 6.190 2.090 ;
        RECT 5.750 1.890 5.940 1.920 ;
        RECT 6.470 1.830 6.640 2.510 ;
        RECT 2.100 1.740 2.420 1.770 ;
        RECT 5.180 1.750 5.500 1.780 ;
        RECT 2.100 1.460 2.420 1.490 ;
        RECT 0.070 1.110 0.240 1.390 ;
        RECT 0.580 1.150 0.930 1.320 ;
        RECT 0.750 1.120 0.930 1.150 ;
        RECT 1.350 1.130 1.520 1.400 ;
        RECT 2.100 1.270 2.430 1.460 ;
        RECT 5.180 1.450 5.500 1.480 ;
        RECT 2.100 1.230 2.420 1.270 ;
        RECT 0.070 1.070 0.280 1.110 ;
        RECT 0.750 1.090 1.070 1.120 ;
        RECT 0.070 1.050 0.300 1.070 ;
        RECT 0.070 1.030 0.330 1.050 ;
        RECT 0.070 0.980 0.410 1.030 ;
        RECT 0.070 0.920 0.560 0.980 ;
        RECT 0.070 0.890 0.580 0.920 ;
        RECT 0.110 0.860 0.580 0.890 ;
        RECT 0.750 0.900 1.080 1.090 ;
        RECT 1.350 0.910 1.550 1.130 ;
        RECT 2.130 1.060 2.300 1.230 ;
        RECT 2.820 1.110 2.990 1.400 ;
        RECT 3.780 1.120 3.950 1.400 ;
        RECT 4.520 1.120 4.690 1.410 ;
        RECT 5.180 1.260 5.510 1.450 ;
        RECT 5.750 1.310 5.940 1.340 ;
        RECT 5.180 1.220 5.500 1.260 ;
        RECT 1.360 0.900 1.550 0.910 ;
        RECT 0.750 0.860 1.070 0.900 ;
        RECT 2.810 0.880 3.000 1.110 ;
        RECT 3.670 1.090 3.990 1.120 ;
        RECT 3.670 0.900 4.000 1.090 ;
        RECT 3.670 0.860 3.990 0.900 ;
        RECT 4.520 0.890 4.710 1.120 ;
        RECT 5.240 1.060 5.410 1.220 ;
        RECT 5.750 1.140 6.190 1.310 ;
        RECT 5.750 1.110 5.940 1.140 ;
        RECT 0.240 0.810 0.580 0.860 ;
        RECT 0.360 0.800 0.580 0.810 ;
        RECT 0.370 0.770 0.580 0.800 ;
        RECT 0.390 0.690 0.580 0.770 ;
        RECT 1.750 0.690 2.080 0.810 ;
        RECT 6.470 0.720 6.640 1.400 ;
        RECT -0.100 0.640 0.070 0.660 ;
        RECT -0.120 0.210 0.090 0.640 ;
        RECT 0.390 0.520 0.910 0.690 ;
        RECT 0.390 0.490 0.580 0.520 ;
        RECT 1.260 0.510 5.480 0.690 ;
        RECT 6.210 0.680 6.640 0.720 ;
        RECT 5.860 0.520 6.640 0.680 ;
        RECT 5.860 0.510 6.400 0.520 ;
        RECT 6.210 0.490 6.400 0.510 ;
        RECT -0.120 -0.430 0.090 0.000 ;
        RECT 0.390 -0.310 0.580 -0.280 ;
        RECT 6.210 -0.300 6.400 -0.280 ;
        RECT -0.100 -0.450 0.070 -0.430 ;
        RECT 0.390 -0.480 0.910 -0.310 ;
        RECT 1.260 -0.480 5.480 -0.300 ;
        RECT 5.860 -0.310 6.400 -0.300 ;
        RECT 5.860 -0.470 6.640 -0.310 ;
        RECT 0.390 -0.560 0.580 -0.480 ;
        RECT 0.370 -0.590 0.580 -0.560 ;
        RECT 0.360 -0.600 0.580 -0.590 ;
        RECT 1.750 -0.600 2.080 -0.480 ;
        RECT 6.210 -0.510 6.640 -0.470 ;
        RECT 0.240 -0.650 0.580 -0.600 ;
        RECT 0.110 -0.680 0.580 -0.650 ;
        RECT 0.070 -0.710 0.580 -0.680 ;
        RECT 0.750 -0.690 1.070 -0.650 ;
        RECT 0.070 -0.770 0.560 -0.710 ;
        RECT 0.070 -0.820 0.410 -0.770 ;
        RECT 0.070 -0.840 0.330 -0.820 ;
        RECT 0.070 -0.860 0.300 -0.840 ;
        RECT 0.070 -0.900 0.280 -0.860 ;
        RECT 0.750 -0.880 1.080 -0.690 ;
        RECT 1.360 -0.700 1.550 -0.690 ;
        RECT 0.070 -1.180 0.240 -0.900 ;
        RECT 0.750 -0.910 1.070 -0.880 ;
        RECT 0.750 -0.940 0.930 -0.910 ;
        RECT 0.580 -1.110 0.930 -0.940 ;
        RECT 1.350 -0.920 1.550 -0.700 ;
        RECT 1.350 -1.190 1.520 -0.920 ;
        RECT 2.130 -1.020 2.300 -0.850 ;
        RECT 2.810 -0.900 3.000 -0.670 ;
        RECT 3.670 -0.690 3.990 -0.650 ;
        RECT 3.670 -0.880 4.000 -0.690 ;
        RECT 2.100 -1.060 2.420 -1.020 ;
        RECT 2.100 -1.250 2.430 -1.060 ;
        RECT 2.820 -1.190 2.990 -0.900 ;
        RECT 3.670 -0.910 3.990 -0.880 ;
        RECT 4.520 -0.910 4.710 -0.680 ;
        RECT 3.780 -1.190 3.950 -0.910 ;
        RECT 4.520 -1.200 4.690 -0.910 ;
        RECT 5.240 -1.010 5.410 -0.850 ;
        RECT 5.750 -0.930 5.940 -0.900 ;
        RECT 5.180 -1.050 5.500 -1.010 ;
        RECT 5.180 -1.240 5.510 -1.050 ;
        RECT 5.750 -1.100 6.190 -0.930 ;
        RECT 5.750 -1.130 5.940 -1.100 ;
        RECT 6.470 -1.190 6.640 -0.510 ;
        RECT 2.100 -1.280 2.420 -1.250 ;
        RECT 5.180 -1.270 5.500 -1.240 ;
      LAYER mcon ;
        RECT 2.160 4.300 2.330 4.470 ;
        RECT 0.810 3.930 0.980 4.100 ;
        RECT 1.370 3.950 1.540 4.120 ;
        RECT 5.240 4.290 5.410 4.460 ;
        RECT 2.820 3.930 2.990 4.100 ;
        RECT 3.730 3.930 3.900 4.100 ;
        RECT 4.530 3.940 4.700 4.110 ;
        RECT 5.760 4.160 5.930 4.330 ;
        RECT -0.100 3.510 0.070 3.680 ;
        RECT 0.400 3.540 0.570 3.710 ;
        RECT 6.220 3.540 6.390 3.710 ;
        RECT 0.400 2.540 0.570 2.710 ;
        RECT 6.220 2.540 6.390 2.710 ;
        RECT 0.810 2.150 0.980 2.320 ;
        RECT 1.370 2.130 1.540 2.300 ;
        RECT 2.820 2.150 2.990 2.320 ;
        RECT 3.730 2.150 3.900 2.320 ;
        RECT 4.530 2.140 4.700 2.310 ;
        RECT 2.160 1.780 2.330 1.950 ;
        RECT 5.240 1.790 5.410 1.960 ;
        RECT 5.760 1.920 5.930 2.090 ;
        RECT 2.160 1.280 2.330 1.450 ;
        RECT 0.810 0.910 0.980 1.080 ;
        RECT 1.370 0.930 1.540 1.100 ;
        RECT 5.240 1.270 5.410 1.440 ;
        RECT 2.820 0.910 2.990 1.080 ;
        RECT 3.730 0.910 3.900 1.080 ;
        RECT 4.530 0.920 4.700 1.090 ;
        RECT 5.760 1.140 5.930 1.310 ;
        RECT -0.100 0.490 0.070 0.660 ;
        RECT 0.400 0.520 0.570 0.690 ;
        RECT 6.220 0.520 6.390 0.690 ;
        RECT 0.400 -0.480 0.570 -0.310 ;
        RECT 6.220 -0.480 6.390 -0.310 ;
        RECT 0.810 -0.870 0.980 -0.700 ;
        RECT 1.370 -0.890 1.540 -0.720 ;
        RECT 2.820 -0.870 2.990 -0.700 ;
        RECT 3.730 -0.870 3.900 -0.700 ;
        RECT 4.530 -0.880 4.700 -0.710 ;
        RECT 2.160 -1.240 2.330 -1.070 ;
        RECT 5.240 -1.230 5.410 -1.060 ;
        RECT 5.760 -1.100 5.930 -0.930 ;
      LAYER met1 ;
        RECT 2.090 4.220 2.410 4.540 ;
        RECT 5.170 4.210 5.490 4.530 ;
        RECT 0.740 3.850 1.060 4.170 ;
        RECT 1.340 3.890 1.570 4.180 ;
        RECT -0.130 3.550 0.100 3.740 ;
        RECT 1.360 3.630 1.530 3.890 ;
        RECT 2.790 3.870 3.020 4.160 ;
        RECT -0.130 3.450 0.220 3.550 ;
        RECT -0.120 3.230 0.220 3.450 ;
        RECT 1.350 3.310 1.610 3.630 ;
        RECT 2.810 3.620 2.980 3.870 ;
        RECT 3.660 3.850 3.980 4.170 ;
        RECT 4.500 3.880 4.730 4.170 ;
        RECT 5.730 4.100 5.960 4.390 ;
        RECT 2.770 3.300 3.030 3.620 ;
        RECT 4.530 3.600 4.700 3.880 ;
        RECT 5.730 3.610 5.920 4.100 ;
        RECT 4.520 3.280 4.780 3.600 ;
        RECT 5.560 3.360 5.920 3.610 ;
        RECT 5.560 3.290 5.820 3.360 ;
        RECT -0.120 2.800 0.220 3.020 ;
        RECT -0.130 2.700 0.220 2.800 ;
        RECT -0.130 2.510 0.100 2.700 ;
        RECT 1.350 2.620 1.610 2.940 ;
        RECT 2.770 2.630 3.030 2.950 ;
        RECT 4.520 2.650 4.780 2.970 ;
        RECT 5.560 2.890 5.820 2.960 ;
        RECT 0.740 2.080 1.060 2.400 ;
        RECT 1.360 2.360 1.530 2.620 ;
        RECT 2.810 2.380 2.980 2.630 ;
        RECT 1.340 2.070 1.570 2.360 ;
        RECT 2.790 2.090 3.020 2.380 ;
        RECT 3.660 2.080 3.980 2.400 ;
        RECT 4.530 2.370 4.700 2.650 ;
        RECT 5.560 2.640 5.920 2.890 ;
        RECT 4.500 2.080 4.730 2.370 ;
        RECT 5.730 2.150 5.920 2.640 ;
        RECT 2.090 1.710 2.410 2.030 ;
        RECT 5.170 1.720 5.490 2.040 ;
        RECT 5.730 1.860 5.960 2.150 ;
        RECT 2.090 1.200 2.410 1.520 ;
        RECT 5.170 1.190 5.490 1.510 ;
        RECT 0.740 0.830 1.060 1.150 ;
        RECT 1.340 0.870 1.570 1.160 ;
        RECT -0.130 0.530 0.100 0.720 ;
        RECT 1.360 0.610 1.530 0.870 ;
        RECT 2.790 0.850 3.020 1.140 ;
        RECT -0.130 0.430 0.220 0.530 ;
        RECT -0.120 0.210 0.220 0.430 ;
        RECT 1.350 0.290 1.610 0.610 ;
        RECT 2.810 0.600 2.980 0.850 ;
        RECT 3.660 0.830 3.980 1.150 ;
        RECT 4.500 0.860 4.730 1.150 ;
        RECT 5.730 1.080 5.960 1.370 ;
        RECT 2.770 0.280 3.030 0.600 ;
        RECT 4.530 0.580 4.700 0.860 ;
        RECT 5.730 0.590 5.920 1.080 ;
        RECT 4.520 0.260 4.780 0.580 ;
        RECT 5.560 0.340 5.920 0.590 ;
        RECT 5.560 0.270 5.820 0.340 ;
        RECT -0.120 -0.220 0.220 0.000 ;
        RECT -0.130 -0.320 0.220 -0.220 ;
        RECT -0.130 -0.510 0.100 -0.320 ;
        RECT 1.350 -0.400 1.610 -0.080 ;
        RECT 2.770 -0.390 3.030 -0.070 ;
        RECT 4.520 -0.370 4.780 -0.050 ;
        RECT 5.560 -0.130 5.820 -0.060 ;
        RECT 0.740 -0.940 1.060 -0.620 ;
        RECT 1.360 -0.660 1.530 -0.400 ;
        RECT 2.810 -0.640 2.980 -0.390 ;
        RECT 1.340 -0.950 1.570 -0.660 ;
        RECT 2.790 -0.930 3.020 -0.640 ;
        RECT 3.660 -0.940 3.980 -0.620 ;
        RECT 4.530 -0.650 4.700 -0.370 ;
        RECT 5.560 -0.380 5.920 -0.130 ;
        RECT 4.500 -0.940 4.730 -0.650 ;
        RECT 5.730 -0.870 5.920 -0.380 ;
        RECT 2.090 -1.310 2.410 -0.990 ;
        RECT 5.170 -1.300 5.490 -0.980 ;
        RECT 5.730 -1.160 5.960 -0.870 ;
      LAYER via ;
        RECT 2.120 4.250 2.380 4.510 ;
        RECT 5.200 4.240 5.460 4.500 ;
        RECT 0.770 3.880 1.030 4.140 ;
        RECT 3.690 3.880 3.950 4.140 ;
        RECT -0.040 3.260 0.220 3.520 ;
        RECT 1.350 3.340 1.610 3.600 ;
        RECT 2.770 3.330 3.030 3.590 ;
        RECT 4.520 3.310 4.780 3.570 ;
        RECT 5.560 3.320 5.820 3.580 ;
        RECT -0.040 2.730 0.220 2.990 ;
        RECT 1.350 2.650 1.610 2.910 ;
        RECT 2.770 2.660 3.030 2.920 ;
        RECT 4.520 2.680 4.780 2.940 ;
        RECT 5.560 2.670 5.820 2.930 ;
        RECT 0.770 2.110 1.030 2.370 ;
        RECT 3.690 2.110 3.950 2.370 ;
        RECT 2.120 1.740 2.380 2.000 ;
        RECT 5.200 1.750 5.460 2.010 ;
        RECT 2.120 1.230 2.380 1.490 ;
        RECT 5.200 1.220 5.460 1.480 ;
        RECT 0.770 0.860 1.030 1.120 ;
        RECT 3.690 0.860 3.950 1.120 ;
        RECT -0.040 0.240 0.220 0.500 ;
        RECT 1.350 0.320 1.610 0.580 ;
        RECT 2.770 0.310 3.030 0.570 ;
        RECT 4.520 0.290 4.780 0.550 ;
        RECT 5.560 0.300 5.820 0.560 ;
        RECT -0.040 -0.290 0.220 -0.030 ;
        RECT 1.350 -0.370 1.610 -0.110 ;
        RECT 2.770 -0.360 3.030 -0.100 ;
        RECT 4.520 -0.340 4.780 -0.080 ;
        RECT 5.560 -0.350 5.820 -0.090 ;
        RECT 0.770 -0.910 1.030 -0.650 ;
        RECT 3.690 -0.910 3.950 -0.650 ;
        RECT 2.120 -1.280 2.380 -1.020 ;
        RECT 5.200 -1.270 5.460 -1.010 ;
  END
END sky130_hilas_Tgate4Double01

END LIBRARY