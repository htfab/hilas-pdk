* Qucs 0.0.22 /home/ubuntu/.qucs/Hilas_prj/Trans2med.sch
* Qucs 0.0.22  /home/ubuntu/.qucs/Hilas_prj/Trans2med.sch
M1 _net0  Gate2p  Drain2p  Well MOSP
M4 Drain2n  Gate2n  Source2n  0 MOSN
M5 Drain1n  Gate1n  Source1n  0 MOSN
M6 _net1  Gate1p  Drain1p  Well MOSP
.control
echo "" > spice4qucs.cir.noise
echo "" > spice4qucs.cir.pz
exit
.endc
.END
