magic
tech sky130A
magscale 1 2
timestamp 1632256349
<< checkpaint >>
rect -990 -1124 1954 2002
<< error_s >>
rect 354 1198 368 1232
rect 382 1214 396 1260
rect 568 1200 576 1250
rect 602 1222 610 1274
rect 14 1096 42 1150
rect 410 1108 474 1110
rect 410 1098 476 1108
rect 384 1080 446 1082
rect 384 1074 448 1080
rect 450 1074 476 1098
rect 390 1070 476 1074
rect 420 1062 476 1070
rect 602 1076 622 1082
rect 602 1066 624 1076
rect 14 1014 46 1048
rect 356 1000 370 1034
rect 384 1016 398 1062
rect 420 1052 486 1062
rect 574 1060 594 1066
rect 422 1050 448 1052
rect 450 1050 476 1052
rect 422 1016 514 1050
rect 426 988 514 1016
rect 570 1008 594 1060
rect 602 1032 626 1066
rect 602 1024 624 1032
rect 602 1018 622 1024
rect 570 1002 578 1008
rect 14 912 42 946
rect 14 830 48 864
rect 70 848 76 892
rect 356 802 370 836
rect 384 818 398 864
rect 422 818 448 882
rect 450 798 476 910
rect 570 804 578 854
rect 604 826 612 878
rect 410 786 588 798
rect 14 756 42 762
rect 14 728 56 756
rect 434 754 526 756
rect 334 726 376 752
rect 410 740 526 754
rect 410 730 458 740
rect 382 724 428 726
rect 382 718 430 724
rect 66 700 84 716
rect 368 702 430 718
rect 14 646 46 680
rect 66 650 74 700
rect 366 692 410 702
rect 366 674 372 692
rect 338 636 344 674
rect 366 666 402 674
rect 366 660 372 666
rect 398 636 402 666
rect 422 660 430 702
rect 434 676 436 698
rect 450 632 458 730
rect 594 626 600 676
rect 628 646 634 698
rect 420 612 471 617
rect 420 604 476 612
rect 14 524 42 562
rect 422 554 448 584
rect 338 532 448 554
rect 338 530 384 532
rect 390 526 448 532
rect 366 520 384 526
rect 422 520 448 526
rect 366 512 432 520
rect 366 500 434 512
rect 366 498 436 500
rect 14 440 42 478
rect 366 476 372 498
rect 338 438 344 476
rect 366 468 402 476
rect 366 462 372 468
rect 398 438 402 468
rect 422 462 430 498
rect 434 478 436 498
rect 450 492 476 604
rect 450 434 458 492
rect 594 428 600 478
rect 628 448 634 500
rect 420 414 471 419
rect 420 406 476 414
rect 14 392 42 394
rect 0 366 42 392
rect 422 380 448 386
rect 14 332 42 366
rect 270 322 448 380
rect 0 282 42 310
rect 14 248 42 282
rect 270 302 434 322
rect 270 280 436 302
rect 450 294 476 406
rect 270 264 434 280
rect 450 264 458 294
rect 270 240 506 264
rect 270 210 514 240
rect 270 208 476 210
rect 14 194 42 196
rect 0 168 42 194
rect 270 188 434 208
rect 270 168 448 188
rect 14 140 448 168
rect 28 126 448 140
rect 28 94 398 126
rect 422 124 448 126
rect 450 96 476 208
rect 502 194 514 210
rect 530 166 542 268
rect 594 230 600 280
rect 628 250 634 302
rect 542 126 602 136
rect 14 56 398 94
rect 28 36 398 56
rect 542 36 566 126
<< nwell >>
rect 434 264 542 618
rect 422 210 542 264
rect 434 126 542 210
rect 398 36 542 126
rect 28 0 542 36
<< psubdiff >>
rect 426 1036 514 1050
rect 426 1002 456 1036
rect 490 1002 514 1036
rect 426 988 514 1002
<< nsubdiff >>
rect 422 254 506 264
rect 422 220 446 254
rect 480 220 506 254
rect 422 210 506 220
<< psubdiffcont >>
rect 456 1002 490 1036
<< nsubdiffcont >>
rect 446 220 480 254
<< locali >>
rect 80 1024 122 1074
rect 454 1052 488 1062
rect 452 1046 488 1052
rect 452 1036 538 1046
rect 452 1002 456 1036
rect 490 1002 538 1036
rect 452 996 538 1002
rect 452 990 490 996
rect 454 984 490 990
rect 430 220 446 254
rect 480 220 496 254
<< metal1 >>
rect 450 254 494 1176
rect 446 220 494 254
rect 450 0 494 220
rect 530 0 574 1176
<< metal2 >>
rect 14 1142 28 1150
rect 14 1096 42 1142
rect 410 1098 574 1132
rect 14 1014 46 1048
rect 14 912 42 946
rect 410 914 574 948
rect 14 830 48 864
rect 14 756 42 762
rect 14 728 56 756
rect 410 730 574 764
rect 14 646 46 680
rect 14 524 42 562
rect 414 510 574 550
rect 14 440 42 478
rect 14 366 42 370
rect 14 332 28 366
rect 414 318 574 358
rect 14 282 42 286
rect 14 248 28 282
rect 14 168 42 178
rect 14 140 28 168
rect 412 126 574 166
rect 14 90 42 94
rect 14 56 44 90
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1632251332
transform 0 1 456 -1 0 240
box 0 0 46 58
use sky130_hilas_pFETdevice01e  sky130_hilas_pFETdevice01e_2
timestamp 1632256325
transform 1 0 270 0 1 136
box 0 0 424 210
use sky130_hilas_pFETdevice01e  sky130_hilas_pFETdevice01e_1
timestamp 1632256325
transform 1 0 270 0 1 334
box 0 0 424 210
use sky130_hilas_pFETdevice01e  sky130_hilas_pFETdevice01e_0
timestamp 1632256325
transform 1 0 270 0 1 532
box 0 0 424 210
use sky130_hilas_nFET03a  sky130_hilas_nFET03a_0
timestamp 1632255311
transform 1 0 250 0 1 716
box 0 0 420 180
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1632251356
transform 1 0 66 0 1 650
box 0 0 68 66
use sky130_hilas_nFET03a  sky130_hilas_nFET03a_1
timestamp 1632255311
transform 1 0 250 0 1 914
box 0 0 420 180
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1632251356
transform 1 0 70 0 1 848
box 0 0 68 66
use sky130_hilas_nFET03a  sky130_hilas_nFET03a_3
timestamp 1632255311
transform 1 0 248 0 1 1112
box 0 0 420 180
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1632251332
transform 1 0 548 0 1 1008
box 0 0 46 58
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1632251356
transform 1 0 74 0 1 1032
box 0 0 68 66
<< labels >>
rlabel metal1 450 0 494 18 0 WELL
port 13 nsew power default
rlabel metal1 530 0 574 18 0 VGND
port 14 nsew ground default
rlabel metal1 450 1158 494 1176 0 WELL
port 13 nsew ground default
rlabel metal1 530 1158 574 1176 0 VGND
port 14 nsew power default
rlabel metal2 14 1096 28 1130 0 NFET_SOURCE1
port 1 nsew analog default
rlabel metal2 14 1014 28 1048 0 NFET_GATE1
port 2 nsew analog default
rlabel metal2 14 912 28 946 0 NFET_SOURCE2
port 3 nsew analog default
rlabel metal2 14 830 28 864 0 NFET_GATE2
port 4 nsew analog default
rlabel metal2 14 728 28 762 0 NFET_SOURCE3
port 5 nsew analog default
rlabel metal2 14 646 28 680 0 NFET_GATE3
port 6 nsew analog default
rlabel metal2 14 440 28 478 0 PFET_GATE1
port 8 nsew analog default
rlabel metal2 14 524 28 562 0 PFET_SOURCE1
port 7 nsew analog default
rlabel metal2 14 332 28 370 0 PFET_SOURCE2
port 9 nsew analog default
rlabel metal2 14 248 28 286 0 PFET_GATE2
port 10 nsew analog default
rlabel metal2 14 140 28 178 0 PFET_SOURCE3
port 11 nsew analog default
rlabel metal2 14 56 28 94 0 PFET_GATE3
port 12 nsew analog default
rlabel metal2 562 510 574 550 0 PFET_DRAIN1
port 17 nsew analog default
rlabel metal2 562 318 574 358 0 PFET_DRAIN2
port 16 nsew analog default
rlabel metal2 562 126 574 166 0 PFET_DRAIN3
port 15 nsew analog default
rlabel metal2 564 1098 574 1132 0 NFET_DRAIN1
port 20 nsew analog default
rlabel metal2 564 914 574 948 0 NFET_DRAIN2
port 19 nsew analog default
rlabel metal2 564 730 574 764 0 NFET_DRAIN3
port 18 nsew analog default
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
