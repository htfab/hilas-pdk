magic
tech sky130A
timestamp 1629137210
<< checkpaint >>
rect -630 681 663 816
rect -630 -495 821 681
rect -472 -630 821 -495
<< error_s >>
rect 67 148 106 151
rect 67 106 106 109
<< nwell >>
rect 6 50 167 171
<< pmos >>
rect 67 109 106 148
<< pdiff >>
rect 40 137 67 148
rect 40 120 44 137
rect 61 120 67 137
rect 40 109 67 120
rect 106 137 133 148
rect 106 120 112 137
rect 129 120 133 137
rect 106 109 133 120
<< pdiffc >>
rect 44 120 61 137
rect 112 120 129 137
<< poly >>
rect 67 148 106 161
rect 67 101 106 109
rect 67 86 157 101
rect 141 69 157 86
rect 141 58 158 69
rect 141 54 157 58
rect 143 52 157 54
rect 143 44 149 52
<< locali >>
rect 44 137 61 145
rect 44 112 61 120
rect 112 137 129 145
rect 112 112 129 120
use sky130_hilas_poly2m1  sky130_hilas_poly2m1_2
timestamp 1629137133
transform 1 0 158 0 -1 51
box 0 0 33 51
use sky130_hilas_poly2m1  sky130_hilas_poly2m1_0
timestamp 1629137133
transform 1 0 0 0 1 135
box 0 0 33 51
<< end >>
