magic
tech sky130A
timestamp 1627250433
<< error_s >>
rect -539 538 -533 544
rect -434 538 -428 544
rect 432 538 438 544
rect 537 538 543 544
rect -113 528 -107 534
rect -60 528 -54 534
rect 58 528 64 534
rect 111 528 117 534
rect -545 474 -539 480
rect -428 474 -422 480
rect -119 478 -113 484
rect -54 478 -48 484
rect 52 478 58 484
rect 117 478 123 484
rect 426 474 432 480
rect 543 474 549 480
rect -539 421 -533 427
rect -434 421 -428 427
rect -113 419 -107 425
rect -60 419 -54 425
rect 58 419 64 425
rect 111 419 117 425
rect 432 421 438 427
rect 537 421 543 427
rect -119 369 -113 375
rect -54 369 -48 375
rect 52 369 58 375
rect 117 369 123 375
rect -545 357 -539 363
rect -428 357 -422 363
rect 426 357 432 363
rect 543 357 549 363
rect -539 236 -533 242
rect -434 236 -428 242
rect 432 236 438 242
rect 537 236 543 242
rect -113 230 -107 236
rect -60 230 -54 236
rect 58 230 64 236
rect 111 230 117 236
rect -119 180 -113 186
rect -54 180 -48 186
rect 52 180 58 186
rect 117 180 123 186
rect -545 172 -539 178
rect -428 172 -422 178
rect 426 172 432 178
rect 543 172 549 178
rect -539 120 -533 126
rect -434 120 -428 126
rect 432 120 438 126
rect 537 120 543 126
rect -113 113 -107 119
rect -60 113 -54 119
rect 58 113 64 119
rect 111 113 117 119
rect -119 63 -113 69
rect -54 63 -48 69
rect 52 63 58 69
rect 117 63 123 69
rect -545 56 -539 62
rect -428 56 -422 62
rect 426 56 432 62
rect 543 56 549 62
<< metal1 >>
rect -968 597 -952 601
rect -984 595 -952 597
rect -927 596 -908 601
rect -887 596 -871 601
rect -984 569 -981 595
rect -955 569 -952 595
rect -693 592 -669 601
rect -475 591 -437 601
rect -300 595 -276 601
rect -72 588 -32 601
rect 36 591 76 601
rect 280 596 304 601
rect 441 591 479 601
rect 673 594 697 601
rect 875 596 891 601
rect 912 596 931 601
rect 956 597 972 601
rect 956 595 988 597
rect -984 567 -952 569
rect -32 565 36 587
rect 956 569 959 595
rect 985 569 988 595
rect 956 567 988 569
rect -968 -4 -952 2
rect -927 -3 -908 3
rect -887 -3 -871 3
rect -693 -4 -669 4
rect -475 -4 -437 5
rect -300 -4 -276 3
rect -72 -4 -32 8
rect 36 -4 76 8
rect 280 -4 304 3
rect 441 -4 479 11
rect 673 -4 697 2
rect 875 -3 891 3
rect 912 -3 931 3
rect 956 -3 972 3
<< via1 >>
rect -981 569 -955 595
rect 959 569 985 595
<< metal2 >>
rect -984 595 -699 597
rect -984 569 -981 595
rect -955 587 -699 595
rect 705 595 988 597
rect 705 587 959 595
rect -955 579 959 587
rect -955 569 -942 579
rect -743 569 725 579
rect 956 569 959 579
rect 985 569 988 595
rect -984 567 -942 569
rect 956 567 988 569
rect -1004 533 -990 552
rect 999 533 1008 551
rect -1004 490 -990 509
rect 999 490 1008 508
rect -1004 390 -989 409
rect 996 390 1009 408
rect -1004 347 -991 365
rect 995 347 1009 365
rect -1004 232 -997 250
rect 1000 232 1009 250
rect -1004 189 -997 207
rect 1000 189 1009 207
rect -334 134 342 152
rect -1004 90 -997 108
rect 1000 90 1009 108
rect -1004 47 -997 65
rect 1000 47 1009 65
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_0
timestamp 1627219133
transform 1 0 264 0 1 378
box -264 -382 744 223
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_1
timestamp 1627219133
transform -1 0 -260 0 1 378
box -264 -382 744 223
<< labels >>
rlabel metal1 441 591 479 601 0 GATE2
port 1 nsew analog default
rlabel metal1 -72 -4 -32 8 0 VTUN
port 2 nsew power default
rlabel metal1 36 -4 76 8 0 VTUN
port 2 nsew power default
rlabel metal1 36 591 76 601 0 VTUN
port 2 nsew power default
rlabel metal1 -72 588 -32 601 0 VTUN
port 2 nsew power default
rlabel metal1 -475 591 -437 601 0 GATE1
port 3 nsew analog default
rlabel metal1 -475 -4 -437 5 0 GATE1
port 3 nsew analog default
rlabel metal1 956 -3 972 3 0 VINJ
port 4 nsew power default
rlabel metal1 441 -4 479 11 0 GATE2
port 1 nsew analog default
rlabel metal1 912 596 931 601 0 SelectGate2
rlabel metal1 956 596 972 601 0 VINJ
port 6 nsew power default
rlabel metal1 -968 596 -952 601 0 VINJ
port 6 nsew power default
rlabel metal1 -927 596 -908 601 0 GATESELECT1
port 10 nsew analog default
rlabel metal1 -968 -4 -952 2 0 VINJ
port 6 nsew power default
rlabel metal1 -927 -3 -908 3 0 GATESELECT1
port 10 nsew analog default
rlabel metal1 -887 596 -871 601 0 COL1
port 12 nsew analog default
rlabel metal1 -887 -3 -871 3 0 COL1
port 12 nsew analog default
rlabel metal1 912 -3 931 3 0 GATESELECT2
port 11 nsew analog default
rlabel metal1 875 -3 891 3 0 COL2
port 13 nsew analog default
rlabel metal1 875 596 891 601 0 COL2
port 13 nsew analog default
rlabel metal2 -1004 490 -997 509 0 ROW1
port 14 nsew analog default
rlabel metal2 -1004 390 -997 409 0 ROW2
port 15 nsew analog default
rlabel metal2 -1004 533 -997 552 0 DRAIN1
port 16 nsew analog default
rlabel metal2 -1004 347 -997 365 0 DRAIN2
port 17 nsew analog default
rlabel metal2 -1004 232 -997 250 0 DRAIN3
port 18 nsew analog default
rlabel metal2 -1004 189 -997 207 0 ROW3
port 19 nsew analog default
rlabel metal2 -1004 90 -997 108 0 ROW4
port 20 nsew analog default
rlabel metal2 -1004 47 -997 65 0 DRAIN4
port 21 nsew analog default
rlabel metal2 999 533 1008 551 0 DRAIN1
port 16 nsew analog default
rlabel metal2 999 490 1008 508 0 ROW1
port 14 nsew analog default
rlabel metal2 1000 390 1009 408 0 ROW2
port 15 nsew
rlabel metal2 1000 347 1009 365 0 DRAIN2
port 17 nsew analog default
rlabel metal2 1000 232 1009 250 0 DRAIN3
port 18 nsew analog default
rlabel metal2 1000 189 1009 207 0 ROW3
port 19 nsew analog default
rlabel metal2 1000 90 1009 108 0 ROW4
port 20 nsew analog default
rlabel metal2 1000 47 1009 65 0 DRAIN4
port 21 nsew
rlabel metal1 -693 595 -669 601 0 VGND
port 22 nsew
rlabel metal1 -693 -4 -669 4 0 VGND
port 22 nsew
rlabel metal1 -300 -4 -276 3 0 VGND
port 22 nsew
rlabel metal1 -300 595 -276 601 0 VGND
port 22 nsew
rlabel metal1 280 -4 304 3 0 VGND
port 22 nsew
rlabel metal1 673 -4 697 2 0 VGND
port 22 nsew
rlabel metal1 280 596 304 601 0 VGND
port 22 nsew
rlabel metal1 673 594 697 601 0 VGND
port 22 nsew
<< end >>
