magic
tech sky130A
timestamp 1627400024
<< error_s >>
rect 58 532 64 538
rect 111 532 117 538
rect 52 482 58 488
rect 117 482 123 488
rect 481 473 487 479
rect 586 473 592 479
rect 475 423 481 429
rect 592 423 598 429
rect 481 172 487 178
rect 586 172 592 178
rect 58 118 64 124
rect 111 118 117 124
rect 475 122 481 128
rect 592 122 598 128
rect 52 68 58 74
rect 117 68 123 74
<< nwell >>
rect 1665 587 1792 605
rect 1145 431 1311 453
rect 1191 270 1219 294
rect 1664 0 1792 19
<< locali >>
rect 283 339 329 348
rect 283 322 286 339
rect 303 322 329 339
rect 283 270 329 322
rect 283 253 286 270
rect 303 253 329 270
rect 283 247 329 253
<< viali >>
rect 286 322 303 339
rect 286 253 303 270
<< metal1 >>
rect 35 598 77 605
rect 405 597 428 605
rect 1057 597 1076 605
rect 1101 597 1129 605
rect 1596 591 1630 605
rect 1663 590 1690 605
rect 279 344 317 348
rect 279 251 283 344
rect 312 251 317 344
rect 279 247 317 251
rect 1596 0 1630 19
rect 1663 0 1690 21
<< via1 >>
rect 1600 439 1626 465
rect 283 339 312 344
rect 283 322 286 339
rect 286 322 303 339
rect 303 322 312 339
rect 283 270 312 322
rect 283 253 286 270
rect 286 253 303 270
rect 303 253 312 270
rect 283 251 312 253
<< metal2 >>
rect 1343 578 1368 604
rect 0 537 7 555
rect 1449 480 1474 517
rect 1596 465 1630 469
rect 1596 460 1600 465
rect 1145 431 1311 453
rect 1361 441 1600 460
rect 1361 384 1380 441
rect 1596 439 1600 441
rect 1626 439 1630 465
rect 1596 436 1630 439
rect 1452 395 1473 424
rect 282 365 1380 384
rect 282 347 301 365
rect 280 344 315 347
rect 280 251 283 344
rect 312 251 315 344
rect 1777 334 1792 356
rect 1347 311 1372 334
rect 1191 270 1219 294
rect 1777 252 1792 274
rect 280 248 315 251
rect 1296 187 1473 207
rect 1139 138 1155 178
rect 1267 106 1473 127
rect 0 52 8 67
rect 1187 2 1213 27
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1608069483
transform 1 0 1637 0 1 41
box -172 -22 155 550
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1608384750
transform 1 0 1145 0 -1 165
box 133 -440 320 165
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_0
timestamp 1608384750
transform 1 0 989 0 1 440
box 133 -440 320 165
use sky130_hilas_FGBias2x1cell  sky130_hilas_FGBias2x1cell_0
timestamp 1625491133
transform 1 0 396 0 1 382
box -396 -382 757 223
<< labels >>
rlabel metal1 1596 0 1630 6 0 VGND
port 7 nsew ground default
rlabel metal1 1663 0 1690 6 0 VPWR
port 8 nsew power default
rlabel metal1 1596 600 1630 605 0 VGND
port 7 nsew ground default
rlabel metal1 1663 600 1690 605 0 VPWR
port 8 nsew power default
rlabel metal2 1347 311 1372 334 0 VIN21
port 3 nsew
rlabel metal2 1187 2 1210 27 0 VIN12
port 2 nsew analog default
rlabel metal2 1343 578 1368 604 0 VIN22
port 4 nsew
rlabel metal2 1777 252 1792 274 0 OUTPUT1
port 5 nsew
rlabel metal2 1777 334 1792 356 0 OUTPUT2
port 6 nsew
rlabel metal1 1057 597 1076 605 0 COLSEL1
port 1 nsew
rlabel metal2 0 537 7 555 0 DRAIN1
port 9 nsew
rlabel metal2 0 52 8 67 0 DRAIN2
port 10 nsew
rlabel metal1 35 598 77 605 0 VTUN
port 11 nsew
rlabel metal1 405 597 428 605 0 GATE1
port 12 nsew
rlabel metal1 1101 597 1129 605 0 VINJ
port 13 nsew
rlabel metal2 1191 270 1214 294 0 VIN11
port 14 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
