magic
tech sky130A
timestamp 1628616987
<< checkpaint >>
rect -658 7833 3642 8386
rect -658 7129 4554 7833
rect 7307 7129 13890 7929
rect -658 5968 13890 7129
rect -658 5709 3642 5968
rect 1438 4660 3220 5709
rect 1629 4510 3220 4660
rect 3716 4337 13890 5968
rect 1393 3972 3006 4115
rect 3716 3995 13286 4337
rect 1393 3497 3473 3972
rect 1151 2119 3473 3497
rect 3712 3734 13286 3995
rect 3712 3280 13257 3734
rect 3712 3103 12297 3280
rect 3712 2750 10585 3103
rect 3712 2205 12216 2750
rect 1151 2117 3330 2119
rect 1151 2095 3183 2117
rect 1151 1634 3041 2095
rect 3712 1948 8395 2205
rect 1179 883 3041 1634
rect 4455 1009 8395 1948
rect 4455 1007 6909 1009
rect 1184 863 3041 883
rect 1184 464 2908 863
rect 9611 -248 12216 2205
rect 9611 -630 11691 -248
<< error_s >>
rect 2694 7164 2723 7180
rect 2773 7164 2802 7180
rect 2852 7164 2881 7180
rect 2931 7164 2960 7180
rect 2694 7130 2695 7131
rect 2722 7130 2723 7131
rect 2773 7130 2774 7131
rect 2801 7130 2802 7131
rect 2852 7130 2853 7131
rect 2880 7130 2881 7131
rect 2931 7130 2932 7131
rect 2959 7130 2960 7131
rect 2644 7101 2661 7130
rect 2693 7129 2724 7130
rect 2772 7129 2803 7130
rect 2851 7129 2882 7130
rect 2930 7129 2961 7130
rect 2694 7122 2723 7129
rect 2773 7122 2802 7129
rect 2852 7122 2881 7129
rect 2931 7122 2960 7129
rect 2694 7108 2703 7122
rect 2950 7108 2960 7122
rect 2694 7102 2723 7108
rect 2773 7102 2802 7108
rect 2852 7102 2881 7108
rect 2931 7102 2960 7108
rect 2693 7101 2724 7102
rect 2772 7101 2803 7102
rect 2851 7101 2882 7102
rect 2930 7101 2961 7102
rect 2992 7101 3010 7130
rect 2694 7100 2695 7101
rect 2722 7100 2723 7101
rect 2773 7100 2774 7101
rect 2801 7100 2802 7101
rect 2852 7100 2853 7101
rect 2880 7100 2881 7101
rect 2931 7100 2932 7101
rect 2959 7100 2960 7101
rect 2694 7051 2723 7066
rect 2773 7051 2802 7066
rect 2852 7051 2881 7066
rect 2931 7051 2960 7066
rect 2694 6884 2723 6900
rect 2773 6884 2802 6900
rect 2852 6884 2881 6900
rect 2931 6884 2960 6900
rect 2694 6850 2695 6851
rect 2722 6850 2723 6851
rect 2773 6850 2774 6851
rect 2801 6850 2802 6851
rect 2852 6850 2853 6851
rect 2880 6850 2881 6851
rect 2931 6850 2932 6851
rect 2959 6850 2960 6851
rect 2644 6821 2661 6850
rect 2693 6849 2724 6850
rect 2772 6849 2803 6850
rect 2851 6849 2882 6850
rect 2930 6849 2961 6850
rect 2694 6842 2723 6849
rect 2773 6842 2802 6849
rect 2852 6842 2881 6849
rect 2931 6842 2960 6849
rect 2694 6828 2703 6842
rect 2950 6828 2960 6842
rect 2694 6822 2723 6828
rect 2773 6822 2802 6828
rect 2852 6822 2881 6828
rect 2931 6822 2960 6828
rect 2693 6821 2724 6822
rect 2772 6821 2803 6822
rect 2851 6821 2882 6822
rect 2930 6821 2961 6822
rect 2992 6821 3010 6850
rect 2694 6820 2695 6821
rect 2722 6820 2723 6821
rect 2773 6820 2774 6821
rect 2801 6820 2802 6821
rect 2852 6820 2853 6821
rect 2880 6820 2881 6821
rect 2931 6820 2932 6821
rect 2959 6820 2960 6821
rect 3790 6802 3819 6820
rect 2694 6771 2723 6786
rect 2773 6771 2802 6786
rect 2852 6771 2881 6786
rect 2931 6771 2960 6786
rect 3790 6770 3791 6771
rect 3818 6770 3819 6771
rect 2694 6729 2723 6745
rect 2773 6729 2802 6745
rect 2852 6729 2881 6745
rect 2931 6729 2960 6745
rect 3740 6741 3758 6770
rect 3789 6769 3820 6770
rect 3790 6760 3819 6769
rect 3790 6751 3800 6760
rect 3809 6751 3819 6760
rect 3790 6742 3819 6751
rect 3789 6741 3820 6742
rect 3851 6741 3869 6770
rect 3790 6740 3791 6741
rect 3818 6740 3819 6741
rect 2694 6695 2695 6696
rect 2722 6695 2723 6696
rect 2773 6695 2774 6696
rect 2801 6695 2802 6696
rect 2852 6695 2853 6696
rect 2880 6695 2881 6696
rect 2931 6695 2932 6696
rect 2959 6695 2960 6696
rect 2644 6666 2661 6695
rect 2693 6694 2724 6695
rect 2772 6694 2803 6695
rect 2851 6694 2882 6695
rect 2930 6694 2961 6695
rect 2694 6687 2723 6694
rect 2773 6687 2802 6694
rect 2852 6687 2881 6694
rect 2931 6687 2960 6694
rect 2694 6673 2703 6687
rect 2950 6673 2960 6687
rect 2694 6667 2723 6673
rect 2773 6667 2802 6673
rect 2852 6667 2881 6673
rect 2931 6667 2960 6673
rect 2693 6666 2724 6667
rect 2772 6666 2803 6667
rect 2851 6666 2882 6667
rect 2930 6666 2961 6667
rect 2992 6666 3010 6695
rect 3790 6691 3819 6709
rect 2694 6665 2695 6666
rect 2722 6665 2723 6666
rect 2773 6665 2774 6666
rect 2801 6665 2802 6666
rect 2852 6665 2853 6666
rect 2880 6665 2881 6666
rect 2931 6665 2932 6666
rect 2959 6665 2960 6666
rect 2694 6616 2723 6631
rect 2773 6616 2802 6631
rect 2852 6616 2881 6631
rect 2931 6616 2960 6631
rect 4572 6062 4600 6068
rect 4714 6061 4742 6068
rect 4849 6062 4899 6068
rect 5172 6061 5222 6067
rect 4572 6020 4600 6026
rect 4714 6019 4742 6026
rect 4849 6020 4899 6026
rect 5172 6019 5222 6025
rect 4523 5990 4551 5996
rect 4763 5990 4791 5996
rect 4920 5990 4971 5996
rect 5101 5995 5151 6001
rect 4523 5948 4551 5954
rect 4763 5948 4791 5954
rect 4920 5948 4971 5954
rect 5101 5953 5151 5959
rect 4572 5887 4600 5893
rect 4714 5886 4742 5893
rect 4849 5887 4899 5893
rect 5172 5886 5222 5892
rect 4572 5845 4600 5851
rect 4714 5844 4742 5851
rect 4849 5845 4899 5851
rect 5172 5844 5222 5850
rect 4523 5815 4551 5821
rect 4763 5815 4791 5821
rect 4920 5815 4971 5821
rect 5101 5820 5151 5826
rect 4523 5773 4551 5779
rect 4763 5773 4791 5779
rect 4920 5773 4971 5779
rect 5101 5778 5151 5784
rect 4572 5712 4600 5718
rect 4714 5711 4742 5718
rect 4849 5712 4899 5718
rect 5172 5711 5222 5717
rect 6016 5684 6066 5690
rect 6088 5684 6138 5690
rect 8057 5684 8107 5690
rect 8129 5684 8179 5690
rect 8517 5688 8544 5694
rect 4572 5670 4600 5676
rect 4714 5669 4742 5676
rect 4849 5670 4899 5676
rect 5172 5669 5222 5675
rect 4523 5640 4551 5646
rect 4763 5640 4791 5646
rect 4920 5640 4971 5646
rect 5101 5645 5151 5651
rect 6016 5642 6066 5648
rect 6088 5642 6138 5648
rect 8057 5642 8107 5648
rect 8129 5642 8179 5648
rect 8517 5646 8544 5652
rect 8517 5621 8544 5627
rect 4523 5598 4551 5604
rect 4763 5598 4791 5604
rect 4920 5598 4971 5604
rect 5101 5603 5151 5609
rect 4572 5537 4600 5543
rect 4714 5536 4742 5543
rect 4849 5537 4899 5543
rect 5172 5536 5222 5542
rect 6201 5540 6204 5590
rect 6243 5540 6246 5590
rect 6337 5540 6339 5590
rect 6379 5540 6381 5590
rect 8517 5579 8544 5585
rect 8517 5538 8544 5544
rect 4572 5495 4600 5501
rect 4714 5494 4742 5501
rect 4849 5495 4899 5501
rect 5172 5494 5222 5500
rect 4523 5465 4551 5471
rect 4763 5465 4791 5471
rect 4920 5465 4971 5471
rect 5101 5470 5151 5476
rect 6201 5461 6204 5511
rect 6243 5461 6246 5511
rect 6337 5461 6339 5511
rect 6379 5461 6381 5511
rect 8517 5496 8544 5502
rect 8517 5471 8544 5477
rect 4523 5423 4551 5429
rect 4763 5423 4791 5429
rect 4920 5423 4971 5429
rect 5101 5428 5151 5434
rect 8517 5429 8544 5435
rect 11275 5431 11315 5437
rect 11425 5431 11465 5437
rect 8517 5388 8544 5394
rect 11275 5389 11315 5395
rect 11425 5389 11465 5395
rect 5426 5371 5476 5376
rect 5606 5371 5656 5377
rect 5746 5371 5796 5376
rect 4523 5362 4551 5368
rect 4763 5362 4791 5368
rect 4920 5362 4971 5368
rect 11199 5365 11239 5370
rect 11425 5363 11465 5370
rect 5101 5357 5151 5363
rect 5426 5329 5476 5334
rect 5606 5329 5656 5335
rect 5746 5329 5796 5334
rect 4523 5320 4551 5326
rect 4763 5320 4791 5326
rect 4920 5320 4971 5326
rect 5101 5315 5151 5321
rect 5426 5304 5476 5310
rect 5746 5304 5796 5310
rect 6201 5308 6204 5358
rect 6243 5308 6246 5358
rect 6337 5308 6339 5358
rect 6379 5308 6381 5358
rect 8517 5346 8544 5352
rect 8517 5321 8544 5327
rect 11199 5323 11239 5328
rect 11425 5321 11465 5328
rect 4572 5290 4600 5296
rect 4714 5290 4742 5297
rect 4849 5290 4899 5296
rect 5172 5291 5222 5297
rect 8517 5279 8544 5285
rect 5426 5262 5476 5268
rect 5746 5262 5796 5268
rect 4572 5248 4600 5254
rect 4714 5248 4742 5255
rect 4849 5248 4899 5254
rect 5172 5249 5222 5255
rect 6201 5229 6204 5279
rect 6243 5229 6246 5279
rect 6337 5229 6339 5279
rect 6379 5229 6381 5279
rect 11199 5261 11239 5266
rect 11425 5261 11465 5268
rect 8517 5238 8544 5244
rect 11199 5219 11239 5224
rect 11425 5219 11465 5226
rect 5426 5201 5476 5207
rect 5746 5201 5796 5207
rect 8517 5196 8544 5202
rect 11275 5194 11315 5200
rect 11425 5194 11465 5200
rect 4523 5187 4551 5193
rect 4763 5187 4791 5193
rect 4920 5187 4971 5193
rect 5101 5182 5151 5188
rect 6016 5171 6066 5177
rect 6088 5171 6138 5177
rect 8057 5171 8107 5177
rect 8129 5171 8179 5177
rect 8517 5171 8544 5177
rect 5426 5159 5476 5165
rect 5746 5159 5796 5165
rect 11275 5152 11315 5158
rect 11425 5152 11465 5158
rect 4523 5145 4551 5151
rect 4763 5145 4791 5151
rect 4920 5145 4971 5151
rect 5101 5140 5151 5146
rect 5426 5135 5476 5140
rect 5606 5134 5656 5140
rect 5746 5135 5796 5140
rect 6016 5129 6066 5135
rect 6088 5129 6138 5135
rect 8057 5129 8107 5135
rect 8129 5129 8179 5135
rect 8517 5129 8544 5135
rect 4572 5115 4600 5121
rect 4714 5115 4742 5122
rect 4849 5115 4899 5121
rect 5172 5116 5222 5122
rect 11275 5111 11315 5117
rect 11425 5111 11465 5117
rect 5426 5093 5476 5098
rect 5606 5092 5656 5098
rect 5746 5093 5796 5098
rect 6017 5081 6067 5087
rect 6089 5081 6139 5087
rect 8057 5081 8107 5087
rect 8129 5081 8179 5087
rect 8517 5085 8544 5091
rect 4572 5073 4600 5079
rect 4714 5073 4742 5080
rect 4849 5073 4899 5079
rect 5172 5074 5222 5080
rect 11275 5069 11315 5075
rect 11425 5069 11465 5075
rect 5426 5051 5476 5056
rect 5606 5051 5656 5057
rect 5746 5051 5796 5056
rect 6017 5039 6067 5045
rect 6089 5039 6139 5045
rect 8057 5039 8107 5045
rect 8129 5039 8179 5045
rect 8517 5043 8544 5049
rect 11199 5045 11239 5050
rect 11425 5043 11465 5050
rect 8517 5018 8544 5024
rect 4523 5012 4551 5018
rect 4763 5012 4791 5018
rect 4920 5012 4971 5018
rect 5101 5007 5151 5013
rect 5426 5009 5476 5014
rect 5606 5009 5656 5015
rect 5746 5009 5796 5014
rect 11199 5003 11239 5008
rect 11425 5001 11465 5008
rect 5426 4984 5476 4990
rect 5746 4984 5796 4990
rect 8517 4976 8544 4982
rect 4523 4970 4551 4976
rect 4763 4970 4791 4976
rect 4920 4970 4971 4976
rect 5101 4965 5151 4971
rect 4572 4940 4600 4946
rect 4714 4940 4742 4947
rect 4849 4940 4899 4946
rect 5172 4941 5222 4947
rect 5426 4942 5476 4948
rect 5746 4942 5796 4948
rect 11199 4941 11239 4946
rect 11425 4941 11465 4948
rect 8517 4935 8544 4941
rect 4572 4898 4600 4904
rect 4714 4898 4742 4905
rect 4849 4898 4899 4904
rect 5172 4899 5222 4905
rect 11199 4899 11239 4904
rect 11425 4899 11465 4906
rect 8517 4893 8544 4899
rect 5426 4881 5476 4887
rect 5746 4881 5796 4887
rect 11275 4874 11315 4880
rect 11425 4874 11465 4880
rect 8517 4868 8544 4874
rect 4523 4837 4551 4843
rect 4763 4837 4791 4843
rect 4920 4837 4971 4843
rect 5426 4839 5476 4845
rect 5746 4839 5796 4845
rect 5101 4832 5151 4838
rect 11275 4832 11315 4838
rect 11425 4832 11465 4838
rect 8517 4826 8544 4832
rect 5426 4815 5476 4820
rect 5606 4814 5656 4820
rect 5746 4815 5796 4820
rect 4523 4795 4551 4801
rect 4763 4795 4791 4801
rect 4920 4795 4971 4801
rect 5101 4790 5151 4796
rect 8517 4785 8544 4791
rect 5426 4773 5476 4778
rect 5606 4772 5656 4778
rect 5746 4773 5796 4778
rect 4572 4765 4600 4771
rect 4714 4765 4742 4772
rect 4849 4765 4899 4771
rect 5172 4766 5222 4772
rect 8517 4743 8544 4749
rect 4572 4723 4600 4729
rect 4714 4723 4742 4730
rect 4849 4723 4899 4729
rect 5172 4724 5222 4730
rect 8517 4718 8544 4724
rect 8517 4676 8544 4682
rect 8517 4635 8544 4641
rect 8517 4593 8544 4599
rect 6017 4568 6067 4574
rect 6089 4568 6139 4574
rect 8057 4568 8107 4574
rect 8129 4568 8179 4574
rect 8517 4568 8544 4574
rect 6017 4526 6067 4532
rect 6089 4526 6139 4532
rect 8057 4526 8107 4532
rect 8129 4526 8179 4532
rect 8517 4526 8544 4532
rect 4523 4349 4551 4355
rect 4763 4349 4791 4355
rect 4920 4349 4971 4355
rect 5101 4344 5151 4350
rect 5424 4324 5474 4329
rect 5604 4324 5654 4330
rect 5744 4324 5794 4329
rect 6158 4323 6208 4329
rect 6230 4323 6280 4329
rect 7914 4323 7964 4329
rect 7986 4323 8036 4329
rect 4523 4307 4551 4313
rect 4763 4307 4791 4313
rect 4920 4307 4971 4313
rect 5101 4302 5151 4308
rect 4572 4277 4600 4283
rect 4714 4277 4742 4284
rect 4849 4277 4899 4283
rect 5172 4278 5222 4284
rect 5424 4282 5474 4287
rect 5604 4282 5654 4288
rect 5744 4282 5794 4287
rect 6158 4281 6208 4287
rect 6230 4281 6280 4287
rect 7914 4281 7964 4287
rect 7986 4281 8036 4287
rect 5424 4257 5474 4263
rect 5744 4257 5794 4263
rect 6230 4254 6280 4260
rect 7914 4254 7964 4260
rect 4572 4235 4600 4241
rect 4714 4235 4742 4242
rect 4849 4235 4899 4241
rect 5172 4236 5222 4242
rect 5424 4215 5474 4221
rect 5744 4215 5794 4221
rect 6230 4212 6280 4218
rect 7914 4212 7964 4218
rect 4523 4174 4551 4180
rect 4763 4174 4791 4180
rect 4920 4174 4971 4180
rect 5101 4169 5151 4175
rect 6230 4169 6280 4175
rect 7914 4169 7964 4175
rect 5424 4154 5474 4160
rect 5744 4154 5794 4160
rect 4523 4132 4551 4138
rect 4763 4132 4791 4138
rect 4920 4132 4971 4138
rect 5101 4127 5151 4133
rect 6230 4127 6280 4133
rect 7914 4127 7964 4133
rect 5424 4112 5474 4118
rect 5744 4112 5794 4118
rect 4572 4102 4600 4108
rect 4714 4102 4742 4109
rect 4849 4102 4899 4108
rect 5172 4103 5222 4109
rect 6158 4100 6208 4106
rect 6230 4100 6280 4106
rect 7914 4100 7964 4106
rect 7986 4100 8036 4106
rect 5424 4088 5474 4093
rect 5604 4087 5654 4093
rect 5744 4088 5794 4093
rect 4572 4060 4600 4066
rect 4714 4060 4742 4067
rect 4849 4060 4899 4066
rect 5172 4061 5222 4067
rect 6158 4058 6208 4064
rect 6230 4058 6280 4064
rect 7914 4058 7964 4064
rect 7986 4058 8036 4064
rect 5424 4046 5474 4051
rect 5604 4045 5654 4051
rect 5744 4046 5794 4051
rect 4523 3999 4551 4005
rect 4763 3999 4791 4005
rect 4920 3999 4971 4005
rect 5424 4004 5474 4009
rect 5604 4004 5654 4010
rect 5744 4004 5794 4009
rect 5101 3994 5151 4000
rect 6158 3999 6208 4005
rect 6230 3999 6280 4005
rect 7914 3999 7964 4005
rect 7986 3999 8036 4005
rect 4523 3957 4551 3963
rect 4763 3957 4791 3963
rect 4920 3957 4971 3963
rect 5424 3962 5474 3967
rect 5604 3962 5654 3968
rect 5744 3962 5794 3967
rect 5101 3952 5151 3958
rect 6158 3957 6208 3963
rect 6230 3957 6280 3963
rect 7914 3957 7964 3963
rect 7986 3957 8036 3963
rect 5424 3937 5474 3943
rect 5744 3937 5794 3943
rect 4572 3927 4600 3933
rect 4714 3927 4742 3934
rect 4849 3927 4899 3933
rect 5172 3928 5222 3934
rect 6230 3930 6280 3936
rect 7914 3930 7964 3936
rect 5424 3895 5474 3901
rect 5744 3895 5794 3901
rect 4572 3885 4600 3891
rect 4714 3885 4742 3892
rect 4849 3885 4899 3891
rect 5172 3886 5222 3892
rect 6230 3888 6280 3894
rect 7914 3888 7964 3894
rect 6230 3846 6280 3852
rect 7914 3846 7964 3852
rect 5424 3834 5474 3840
rect 5744 3834 5794 3840
rect 4523 3824 4551 3830
rect 4763 3824 4791 3830
rect 4920 3824 4971 3830
rect 5101 3819 5151 3825
rect 6230 3804 6280 3810
rect 7914 3804 7964 3810
rect 5424 3792 5474 3798
rect 5744 3792 5794 3798
rect 4523 3782 4551 3788
rect 4763 3782 4791 3788
rect 4920 3782 4971 3788
rect 5101 3777 5151 3783
rect 6158 3777 6208 3783
rect 6230 3777 6280 3783
rect 7914 3777 7964 3783
rect 7986 3777 8036 3783
rect 5424 3768 5474 3773
rect 5604 3767 5654 3773
rect 5744 3768 5794 3773
rect 4572 3752 4600 3758
rect 4714 3752 4742 3759
rect 4849 3752 4899 3758
rect 5172 3753 5222 3759
rect 6158 3735 6208 3741
rect 6230 3735 6280 3741
rect 7914 3735 7964 3741
rect 7986 3735 8036 3741
rect 5424 3726 5474 3731
rect 5604 3725 5654 3731
rect 5744 3726 5794 3731
rect 4572 3710 4600 3716
rect 4714 3710 4742 3717
rect 4849 3710 4899 3716
rect 5172 3711 5222 3717
rect 4519 3443 4547 3449
rect 4759 3443 4787 3449
rect 4916 3443 4967 3449
rect 5097 3438 5147 3444
rect 4519 3401 4547 3407
rect 4759 3401 4787 3407
rect 4916 3401 4967 3407
rect 5097 3396 5147 3402
rect 5427 3397 5477 3402
rect 5607 3397 5657 3403
rect 5747 3397 5797 3402
rect 6161 3390 6211 3396
rect 6233 3390 6283 3396
rect 4568 3371 4596 3377
rect 4710 3371 4738 3378
rect 4845 3371 4895 3377
rect 5168 3372 5218 3378
rect 5427 3355 5477 3360
rect 5607 3355 5657 3361
rect 5747 3355 5797 3360
rect 6161 3348 6211 3354
rect 6233 3348 6283 3354
rect 4568 3329 4596 3335
rect 4710 3329 4738 3336
rect 4845 3329 4895 3335
rect 5168 3330 5218 3336
rect 5427 3330 5477 3336
rect 5747 3330 5797 3336
rect 6233 3321 6283 3327
rect 5427 3288 5477 3294
rect 5747 3288 5797 3294
rect 6233 3279 6283 3285
rect 4519 3268 4547 3274
rect 4759 3268 4787 3274
rect 4916 3268 4967 3274
rect 5097 3263 5147 3269
rect 6233 3238 6283 3244
rect 4519 3226 4547 3232
rect 4759 3226 4787 3232
rect 4916 3226 4967 3232
rect 5427 3227 5477 3233
rect 5747 3227 5797 3233
rect 5097 3221 5147 3227
rect 4568 3196 4596 3202
rect 4710 3196 4738 3203
rect 4845 3196 4895 3202
rect 5168 3197 5218 3203
rect 6233 3196 6283 3202
rect 5427 3185 5477 3191
rect 5747 3185 5797 3191
rect 6161 3169 6211 3175
rect 6233 3169 6283 3175
rect 5427 3161 5477 3166
rect 4568 3154 4596 3160
rect 4710 3154 4738 3161
rect 4845 3154 4895 3160
rect 5168 3155 5218 3161
rect 5607 3160 5657 3166
rect 5747 3161 5797 3166
rect 6161 3127 6211 3133
rect 6233 3127 6283 3133
rect 5427 3119 5477 3124
rect 5607 3118 5657 3124
rect 5747 3119 5797 3124
rect 4519 3093 4547 3099
rect 4759 3093 4787 3099
rect 4916 3093 4967 3099
rect 5097 3088 5147 3094
rect 5427 3077 5477 3082
rect 5607 3077 5657 3083
rect 5747 3077 5797 3082
rect 6161 3066 6211 3072
rect 6233 3066 6283 3072
rect 4519 3051 4547 3057
rect 4759 3051 4787 3057
rect 4916 3051 4967 3057
rect 5097 3046 5147 3052
rect 5427 3035 5477 3040
rect 5607 3035 5657 3041
rect 5747 3035 5797 3040
rect 4568 3021 4596 3027
rect 4710 3021 4738 3028
rect 4845 3021 4895 3027
rect 5168 3022 5218 3028
rect 6161 3024 6211 3030
rect 6233 3024 6283 3030
rect 5427 3010 5477 3016
rect 5747 3010 5797 3016
rect 6233 2997 6283 3003
rect 4568 2979 4596 2985
rect 4710 2979 4738 2986
rect 4845 2979 4895 2985
rect 5168 2980 5218 2986
rect 5427 2968 5477 2974
rect 5747 2968 5797 2974
rect 6233 2955 6283 2961
rect 4519 2918 4547 2924
rect 4759 2918 4787 2924
rect 4916 2918 4967 2924
rect 5097 2913 5147 2919
rect 6233 2913 6283 2919
rect 5427 2907 5477 2913
rect 5747 2907 5797 2913
rect 4519 2876 4547 2882
rect 4759 2876 4787 2882
rect 4916 2876 4967 2882
rect 5097 2871 5147 2877
rect 6233 2871 6283 2877
rect 5427 2865 5477 2871
rect 5747 2865 5797 2871
rect 4568 2846 4596 2852
rect 4710 2846 4738 2853
rect 4845 2846 4895 2852
rect 5168 2847 5218 2853
rect 5427 2841 5477 2846
rect 5607 2840 5657 2846
rect 5747 2841 5797 2846
rect 6161 2844 6211 2850
rect 6233 2844 6283 2850
rect 4568 2804 4596 2810
rect 4710 2804 4738 2811
rect 4845 2804 4895 2810
rect 5168 2805 5218 2811
rect 5427 2799 5477 2804
rect 5607 2798 5657 2804
rect 5747 2799 5797 2804
rect 6161 2802 6211 2808
rect 6233 2802 6283 2808
rect 10789 1930 10792 1969
rect 10831 1930 10834 1969
rect 10885 1930 10888 1969
rect 10927 1930 10930 1969
rect 10981 1930 10984 1969
rect 11023 1930 11026 1969
rect 11077 1930 11080 1969
rect 11119 1930 11122 1969
rect 11173 1930 11176 1969
rect 11215 1930 11218 1969
rect 11269 1930 11272 1969
rect 11311 1930 11314 1969
rect 10789 1769 10792 1808
rect 10831 1769 10834 1808
rect 10885 1768 10888 1807
rect 10927 1768 10930 1807
rect 10981 1768 10984 1807
rect 11023 1768 11026 1807
rect 11077 1768 11080 1807
rect 11119 1768 11122 1807
rect 11173 1768 11176 1807
rect 11215 1768 11218 1807
rect 11269 1769 11272 1808
rect 11311 1769 11314 1808
rect 10789 1608 10792 1647
rect 10831 1608 10834 1647
rect 10885 1607 10888 1646
rect 10927 1607 10930 1646
rect 10981 1607 10984 1646
rect 11023 1607 11026 1646
rect 11077 1607 11080 1646
rect 11119 1607 11122 1646
rect 11173 1607 11176 1646
rect 11215 1607 11218 1646
rect 11269 1608 11272 1647
rect 11311 1608 11314 1647
rect 10789 1447 10792 1486
rect 10831 1447 10834 1486
rect 10885 1446 10888 1485
rect 10927 1446 10930 1485
rect 10981 1446 10984 1485
rect 11023 1446 11026 1485
rect 11077 1446 11080 1485
rect 11119 1446 11122 1485
rect 11173 1446 11176 1485
rect 11215 1446 11218 1485
rect 11269 1447 11272 1486
rect 11311 1447 11314 1486
rect 10789 1286 10792 1325
rect 10831 1286 10834 1325
rect 10885 1285 10888 1324
rect 10927 1285 10930 1324
rect 10981 1285 10984 1324
rect 11023 1285 11026 1324
rect 11077 1285 11080 1324
rect 11119 1285 11122 1324
rect 11173 1285 11176 1324
rect 11215 1285 11218 1324
rect 11269 1286 11272 1325
rect 11311 1286 11314 1325
rect 11057 1235 11061 1236
rect 10789 1125 10792 1164
rect 10831 1125 10834 1164
rect 10885 1124 10888 1163
rect 10927 1124 10930 1163
rect 10981 1124 10984 1163
rect 11023 1124 11026 1163
rect 11077 1124 11080 1163
rect 11119 1124 11122 1163
rect 11173 1124 11176 1163
rect 11215 1124 11218 1163
rect 11269 1125 11272 1164
rect 11311 1125 11314 1164
rect 10789 964 10792 1003
rect 10831 964 10834 1003
rect 10885 963 10888 1002
rect 10927 963 10930 1002
rect 10981 963 10984 1002
rect 11023 963 11026 1002
rect 11077 963 11080 1002
rect 11119 963 11122 1002
rect 11173 963 11176 1002
rect 11215 963 11218 1002
rect 11269 964 11272 1003
rect 11311 964 11314 1003
rect 10789 803 10792 842
rect 10831 803 10834 842
rect 10885 802 10888 841
rect 10927 802 10930 841
rect 10981 802 10984 841
rect 11023 802 11026 841
rect 11077 802 11080 841
rect 11119 802 11122 841
rect 11173 802 11176 841
rect 11215 802 11218 841
rect 11269 803 11272 842
rect 11311 803 11314 842
rect 10789 642 10792 681
rect 10831 642 10834 681
rect 10885 641 10888 680
rect 10927 641 10930 680
rect 10981 641 10984 680
rect 11023 641 11026 680
rect 11077 641 11080 680
rect 11119 641 11122 680
rect 11173 641 11176 680
rect 11215 641 11218 680
rect 11269 642 11272 681
rect 11311 642 11314 681
rect 10789 481 10792 520
rect 10831 481 10834 520
rect 10885 481 10888 520
rect 10927 481 10930 520
rect 10981 481 10984 520
rect 11023 481 11026 520
rect 11077 481 11080 520
rect 11119 481 11122 520
rect 11173 481 11176 520
rect 11215 481 11218 520
rect 11269 481 11272 520
rect 11311 481 11314 520
<< nwell >>
rect 5949 5404 5952 5405
rect 4473 5390 4650 5401
rect 5037 5390 5287 5401
rect 5881 5374 5952 5404
rect 5881 5370 5949 5374
rect 5880 4765 5950 5370
rect 6927 5161 6928 5280
rect 6927 5156 6932 5161
rect 6927 5146 6933 5156
rect 6928 5034 6933 5146
rect 8270 5055 8326 5109
rect 5881 4745 5950 4765
rect 5880 2793 6055 3390
rect 5880 2790 6182 2793
rect 6094 2774 6182 2790
rect 6070 2077 6272 2646
rect 11334 465 11469 2012
rect 11333 418 11469 465
<< psubdiff >>
rect 1216 6247 3018 6260
rect 1216 6176 2588 6247
rect 2677 6176 3018 6247
rect 1216 6169 3018 6176
rect 2927 2439 3018 6169
rect 7322 5942 8933 5947
rect 7322 5860 7335 5942
rect 7361 5941 8933 5942
rect 7361 5863 8668 5941
rect 8757 5863 8933 5941
rect 7361 5860 8933 5863
rect 7322 5856 8933 5860
rect 8842 4037 8933 5856
rect 2927 2405 2938 2439
rect 2955 2422 2972 2439
rect 2989 2422 3018 2439
rect 3006 2405 3018 2422
rect 2927 2387 3018 2405
rect 2927 2326 2941 2387
rect 2994 2326 3018 2387
rect 2361 1560 2612 1569
rect 2361 1518 2389 1560
rect 2362 1208 2389 1518
rect 2406 1208 2425 1560
rect 2442 1208 2460 1560
rect 2477 1208 2495 1560
rect 2512 1208 2531 1560
rect 2548 1208 2566 1560
rect 2583 1208 2612 1560
rect 2362 1195 2612 1208
rect 2927 1276 3018 2326
rect 8593 3946 8933 4037
rect 8593 1276 8684 3946
rect 2362 1194 2397 1195
rect 2927 1185 10085 1276
rect 2927 788 3018 1185
<< nsubdiff >>
rect 11375 1981 11432 1989
rect 11375 1587 11388 1981
rect 11379 1527 11388 1587
rect 11375 1426 11388 1527
rect 11379 1366 11388 1426
rect 11375 1265 11388 1366
rect 11378 1205 11388 1265
rect 11375 1103 11388 1205
rect 11379 1043 11388 1103
rect 11375 942 11388 1043
rect 11378 882 11388 942
rect 11375 695 11388 882
rect 11378 486 11388 695
rect 11405 486 11432 1981
rect 11378 474 11432 486
<< psubdiffcont >>
rect 2588 6176 2677 6247
rect 7335 5860 7361 5942
rect 8668 5863 8757 5941
rect 2938 2422 2955 2439
rect 2972 2422 2989 2439
rect 2938 2405 3006 2422
rect 2941 2326 2994 2387
rect 2389 1208 2406 1560
rect 2425 1208 2442 1560
rect 2460 1208 2477 1560
rect 2495 1208 2512 1560
rect 2531 1208 2548 1560
rect 2566 1208 2583 1560
<< nsubdiffcont >>
rect 11388 486 11405 1981
<< locali >>
rect 2530 6252 2682 6253
rect 2530 6250 2685 6252
rect 2530 6176 2537 6250
rect 2580 6247 2685 6250
rect 2580 6176 2588 6247
rect 2677 6176 2685 6247
rect 2530 6173 2685 6176
rect 7327 5942 7394 5944
rect 7327 5860 7335 5942
rect 7361 5860 7366 5942
rect 7392 5860 7394 5942
rect 7327 5857 7394 5860
rect 8555 5942 8765 5944
rect 8555 5863 8561 5942
rect 8593 5941 8765 5942
rect 8593 5863 8668 5941
rect 8757 5863 8765 5941
rect 8555 5859 8765 5863
rect 2930 2405 2938 2439
rect 2969 2422 2972 2439
rect 2930 2397 3006 2405
rect 2932 2387 3006 2397
rect 2932 2326 2941 2387
rect 2994 2326 3006 2387
rect 2932 2318 3006 2326
rect 11388 1982 11425 1989
rect 11388 1981 11408 1982
rect 2365 1560 2604 1565
rect 2365 1528 2371 1560
rect 2370 1208 2371 1528
rect 2388 1208 2389 1560
rect 2406 1208 2407 1560
rect 2424 1208 2425 1560
rect 2442 1208 2443 1560
rect 2477 1208 2495 1560
rect 2529 1208 2531 1560
rect 2565 1208 2566 1560
rect 2583 1208 2584 1560
rect 2601 1208 2604 1560
rect 2370 1202 2604 1208
rect 2370 1201 2603 1202
rect 11405 487 11408 1981
rect 11425 487 11426 502
rect 11405 486 11426 487
rect 11388 477 11426 486
<< viali >>
rect 2537 6176 2580 6250
rect 7366 5860 7392 5942
rect 8561 5863 8593 5942
rect 2952 2422 2955 2439
rect 2955 2422 2969 2439
rect 2989 2422 3006 2439
rect 2952 2405 2969 2422
rect 2989 2405 3006 2422
rect 2371 1208 2388 1560
rect 2407 1208 2424 1560
rect 2443 1208 2460 1560
rect 2512 1208 2529 1560
rect 2548 1208 2565 1560
rect 2584 1208 2601 1560
rect 11408 487 11425 1982
<< metal1 >>
rect 8563 7642 8597 7656
rect 9351 7642 9423 7816
rect 8563 7570 9423 7642
rect 3356 7325 3490 7370
rect 746 7285 796 7289
rect 746 7246 751 7285
rect 790 7246 796 7285
rect 3356 7283 4708 7325
rect 4887 7316 5206 7428
rect 3356 7269 3490 7283
rect 746 7241 796 7246
rect 756 6945 795 7241
rect 2815 7209 3092 7233
rect 2815 7168 2839 7209
rect 756 6940 803 6945
rect 756 6901 759 6940
rect 798 6901 803 6940
rect 756 6896 803 6901
rect 756 6895 801 6896
rect 756 1084 795 6895
rect 897 6810 923 6813
rect 897 6781 923 6784
rect 898 6559 922 6781
rect 889 6556 931 6559
rect 889 6511 931 6514
rect 1478 6435 1507 6627
rect 1476 6432 1517 6435
rect 1476 6374 1484 6432
rect 1513 6374 1517 6432
rect 1476 6368 1517 6374
rect 2814 6299 2838 6622
rect 2809 6294 2843 6299
rect 2809 6268 2813 6294
rect 2839 6268 2843 6294
rect 2809 6265 2843 6268
rect 2534 6255 2583 6256
rect 2533 6250 2584 6255
rect 2533 6176 2537 6250
rect 2580 6176 2584 6250
rect 2141 5386 2164 5734
rect 2208 5672 2230 5734
rect 2477 5706 2499 6161
rect 2533 6140 2584 6176
rect 3068 6162 3092 7209
rect 3399 7176 3702 7203
rect 3870 7177 3896 7283
rect 3396 6259 3427 6629
rect 3388 6256 3427 6259
rect 3388 6225 3392 6256
rect 3423 6225 3427 6256
rect 3388 6222 3427 6225
rect 3675 6208 3702 7176
rect 4666 6958 4708 7283
rect 5047 7034 5089 7316
rect 5047 7031 5094 7034
rect 5047 6989 5050 7031
rect 5092 6989 5094 7031
rect 5047 6986 5094 6989
rect 4662 6955 4710 6958
rect 4662 6913 4665 6955
rect 4707 6913 4710 6955
rect 4662 6910 4710 6913
rect 5217 6796 5261 6799
rect 5217 6749 5261 6752
rect 5789 6796 5833 6799
rect 5789 6749 5833 6752
rect 5968 6793 6041 7432
rect 6483 7417 6581 7432
rect 5968 6749 5971 6793
rect 6015 6749 6041 6793
rect 4775 6694 4819 6697
rect 4775 6647 4819 6650
rect 3792 6308 3817 6623
rect 4496 6374 4528 6378
rect 4496 6373 4499 6374
rect 4487 6348 4499 6373
rect 4525 6348 4528 6374
rect 4487 6344 4528 6348
rect 3788 6305 3821 6308
rect 3788 6279 3792 6305
rect 3818 6279 3821 6305
rect 3788 6272 3821 6279
rect 3671 6206 3705 6208
rect 3671 6180 3675 6206
rect 3702 6180 3705 6206
rect 3671 6177 3705 6180
rect 2528 6137 2584 6140
rect 2528 6130 2542 6137
rect 2517 6102 2542 6130
rect 2577 6102 2584 6137
rect 3063 6159 3097 6162
rect 3063 6133 3067 6159
rect 3093 6133 3097 6159
rect 3063 6130 3097 6133
rect 2517 6090 2584 6102
rect 2517 6087 2583 6090
rect 2517 5706 2539 6087
rect 4487 5994 4511 6344
rect 4781 5987 4812 6647
rect 5224 5989 5253 6749
rect 5343 6650 5346 6694
rect 5390 6650 5393 6694
rect 2639 5917 2674 5921
rect 2639 5878 2644 5917
rect 2670 5878 2674 5917
rect 2639 5875 2674 5878
rect 4282 5905 4319 5908
rect 4282 5879 4284 5905
rect 4317 5879 4319 5905
rect 4282 5877 4319 5879
rect 2579 5839 2604 5851
rect 2576 5836 2608 5839
rect 2576 5796 2580 5836
rect 2606 5796 2608 5836
rect 2576 5793 2608 5796
rect 2579 5714 2604 5793
rect 2579 5711 2608 5714
rect 2579 5685 2582 5711
rect 2579 5682 2608 5685
rect 2205 5669 2231 5672
rect 2205 5640 2231 5643
rect 2208 5580 2230 5640
rect 2202 5577 2230 5580
rect 2228 5551 2230 5577
rect 2202 5548 2230 5551
rect 2208 5488 2230 5548
rect 2203 5485 2230 5488
rect 2229 5459 2230 5485
rect 2203 5456 2230 5459
rect 2138 5383 2164 5386
rect 2138 5354 2164 5357
rect 2141 5290 2164 5354
rect 2134 5287 2164 5290
rect 2160 5261 2164 5287
rect 2134 5258 2164 5261
rect 2141 5194 2164 5258
rect 2138 5191 2164 5194
rect 2138 5162 2164 5165
rect 2141 3687 2164 5162
rect 2208 3687 2230 5456
rect 2579 5622 2604 5682
rect 2579 5619 2608 5622
rect 2579 5593 2582 5619
rect 2579 5590 2608 5593
rect 2579 5530 2604 5590
rect 2579 5527 2605 5530
rect 2579 5498 2605 5501
rect 2130 3684 2164 3687
rect 2130 3637 2134 3684
rect 2160 3637 2164 3684
rect 2130 3634 2164 3637
rect 2196 3684 2230 3687
rect 2196 3637 2198 3684
rect 2224 3637 2230 3684
rect 2196 3634 2230 3637
rect 1999 3560 2022 3567
rect 1995 3534 1998 3560
rect 2024 3534 2027 3560
rect 1950 3523 1973 3527
rect 1946 3520 1973 3523
rect 1972 3494 1973 3520
rect 1946 3491 1973 3494
rect 1015 3435 1087 3437
rect 1015 3369 1018 3435
rect 1084 3369 1087 3435
rect 1015 3367 1087 3369
rect 1016 2852 1082 3367
rect 1950 3139 1973 3491
rect 1999 3287 2022 3534
rect 2141 3525 2164 3634
rect 2208 3561 2230 3634
rect 2384 3563 2411 3567
rect 2206 3558 2232 3561
rect 2206 3529 2232 3532
rect 2382 3560 2411 3563
rect 2409 3533 2411 3560
rect 2382 3530 2411 3533
rect 2140 3522 2166 3525
rect 2140 3493 2166 3496
rect 2329 3376 2358 3379
rect 1999 3250 2072 3287
rect 1950 3132 1976 3139
rect 1948 3131 1976 3132
rect 1945 3129 1977 3131
rect 1945 3103 1948 3129
rect 1974 3103 1977 3129
rect 1945 3100 1977 3103
rect 1535 2954 1578 2957
rect 1535 2917 1539 2954
rect 1576 2917 1578 2954
rect 1535 2914 1578 2917
rect 1016 2849 1090 2852
rect 1016 2783 1022 2849
rect 1088 2783 1090 2849
rect 1016 2780 1090 2783
rect 1540 2333 1577 2914
rect 1999 2500 2022 3250
rect 2384 3233 2411 3530
rect 2372 3208 2411 3233
rect 2432 3523 2456 3527
rect 2432 3520 2458 3523
rect 2432 3491 2458 3494
rect 2432 3177 2456 3491
rect 2372 3154 2456 3177
rect 1999 2477 2244 2500
rect 2212 2444 2244 2477
rect 1536 2330 1579 2333
rect 1536 2293 1538 2330
rect 1575 2293 1579 2330
rect 1536 2290 1579 2293
rect 2288 2287 2321 2290
rect 2274 2279 2292 2287
rect 2250 2255 2292 2279
rect 2288 2251 2292 2255
rect 2318 2251 2321 2287
rect 2288 2248 2321 2251
rect 1837 1756 1866 1759
rect 1837 1724 1866 1727
rect 1838 1667 1864 1724
rect 2432 1688 2456 3154
rect 2477 3087 2499 5162
rect 2517 3348 2539 5162
rect 2579 3463 2604 5498
rect 2641 5421 2667 5875
rect 4218 5740 4257 5742
rect 4218 5707 4221 5740
rect 4254 5707 4257 5740
rect 4218 5705 4257 5707
rect 4160 5592 4199 5595
rect 4160 5559 4164 5592
rect 4197 5559 4199 5592
rect 4160 5556 4199 5559
rect 4096 5432 4135 5435
rect 2641 5418 2669 5421
rect 2641 5392 2643 5418
rect 4096 5399 4100 5432
rect 4133 5399 4135 5432
rect 4096 5397 4135 5399
rect 2641 5389 2669 5392
rect 4099 5396 4133 5397
rect 2641 5325 2667 5389
rect 4035 5377 4069 5378
rect 4034 5375 4070 5377
rect 4034 5342 4036 5375
rect 4069 5342 4070 5375
rect 4034 5338 4070 5342
rect 2641 5322 2670 5325
rect 2641 5296 2644 5322
rect 2641 5293 2670 5296
rect 2641 5229 2667 5293
rect 2641 5226 2669 5229
rect 2641 5200 2643 5226
rect 2641 5197 2669 5200
rect 3973 5218 4009 5221
rect 2579 3461 2605 3463
rect 2578 3460 2606 3461
rect 2578 3434 2579 3460
rect 2605 3434 2606 3460
rect 2578 3433 2606 3434
rect 2579 3431 2605 3433
rect 2513 3345 2545 3348
rect 2513 3319 2517 3345
rect 2543 3319 2545 3345
rect 2513 3316 2545 3319
rect 2473 3084 2501 3087
rect 2473 3058 2475 3084
rect 2473 3055 2501 3058
rect 2477 1758 2499 3055
rect 2517 2534 2539 3316
rect 2517 2531 2546 2534
rect 2517 2489 2519 2531
rect 2545 2489 2546 2531
rect 2517 2486 2546 2489
rect 2517 2290 2539 2486
rect 2515 2287 2541 2290
rect 2515 2248 2541 2251
rect 2517 1786 2539 2248
rect 2579 1924 2604 3431
rect 2641 3030 2667 5197
rect 3973 5185 3975 5218
rect 4008 5185 4009 5218
rect 3973 5182 4009 5185
rect 3908 5065 3949 5068
rect 3908 5032 3912 5065
rect 3945 5032 3949 5065
rect 3908 5028 3949 5032
rect 3855 4908 3891 4911
rect 3855 4875 3856 4908
rect 3889 4875 3891 4908
rect 3855 4872 3891 4875
rect 3797 4366 3830 4368
rect 3791 4361 3830 4366
rect 3791 4328 3794 4361
rect 3827 4328 3830 4361
rect 3791 4324 3830 4328
rect 3734 4205 3767 4207
rect 3729 4202 3768 4205
rect 3729 4169 3731 4202
rect 3764 4169 3768 4202
rect 3729 4166 3768 4169
rect 3672 4050 3705 4051
rect 3669 4047 3705 4050
rect 3702 4014 3705 4047
rect 3669 4011 3705 4014
rect 3607 3899 3646 3903
rect 3607 3866 3609 3899
rect 3642 3866 3646 3899
rect 3607 3863 3646 3866
rect 3540 3382 3583 3386
rect 3540 3349 3545 3382
rect 3578 3349 3583 3382
rect 3540 3346 3583 3349
rect 3474 3225 3515 3229
rect 3474 3192 3478 3225
rect 3511 3192 3515 3225
rect 3474 3189 3515 3192
rect 3413 3061 3452 3065
rect 2640 3027 2671 3030
rect 2640 3001 2643 3027
rect 2669 3001 2671 3027
rect 3413 3028 3416 3061
rect 3449 3028 3452 3061
rect 3413 3025 3452 3028
rect 2640 2998 2671 3001
rect 2575 1921 2605 1924
rect 2575 1888 2577 1921
rect 2603 1888 2605 1921
rect 2575 1884 2605 1888
rect 2517 1772 2541 1786
rect 2473 1755 2504 1758
rect 2473 1726 2474 1755
rect 2503 1726 2504 1755
rect 2473 1723 2504 1726
rect 2518 1709 2541 1772
rect 2353 1685 2456 1688
rect 2353 1625 2358 1685
rect 2418 1632 2456 1685
rect 2517 1706 2541 1709
rect 2418 1625 2432 1632
rect 2353 1621 2432 1625
rect 2517 1567 2539 1706
rect 2364 1560 2606 1567
rect 2364 1208 2371 1560
rect 2388 1208 2407 1560
rect 2424 1208 2443 1560
rect 2460 1208 2512 1560
rect 2529 1208 2548 1560
rect 2565 1208 2584 1560
rect 2601 1208 2606 1560
rect 2364 1199 2606 1208
rect 2641 1170 2667 2998
rect 3344 2917 3385 2920
rect 3344 2884 3348 2917
rect 3381 2884 3385 2917
rect 3344 2881 3385 2884
rect 2923 2519 3016 2531
rect 2923 2448 2944 2519
rect 3002 2448 3016 2519
rect 2923 2439 3016 2448
rect 2923 2405 2952 2439
rect 2969 2405 2989 2439
rect 3006 2405 3016 2439
rect 2923 2366 3016 2405
rect 2932 2318 3006 2366
rect 2632 1166 2667 1170
rect 2632 1132 2636 1166
rect 2662 1132 2667 1166
rect 2632 1129 2667 1132
rect 739 1077 795 1084
rect 739 1038 745 1077
rect 784 1038 795 1077
rect 739 1032 795 1038
rect 3350 547 3383 2881
rect 3345 546 3388 547
rect 3342 544 3391 546
rect 3342 501 3345 544
rect 3388 501 3391 544
rect 3342 500 3391 501
rect 3345 498 3388 500
rect 3415 468 3448 3025
rect 3406 465 3455 468
rect 3406 422 3410 465
rect 3453 422 3455 465
rect 3406 419 3455 422
rect 3480 397 3513 3189
rect 3477 394 3517 397
rect 3477 351 3517 354
rect 3456 311 3514 313
rect 3456 260 3460 311
rect 3511 302 3514 311
rect 3547 302 3580 3346
rect 3611 760 3644 3863
rect 3611 314 3643 760
rect 3672 375 3705 4011
rect 3734 436 3767 4166
rect 3797 503 3830 4324
rect 3857 569 3890 4872
rect 3915 626 3948 5028
rect 3976 693 4009 5182
rect 4035 754 4068 5338
rect 4099 821 4132 5396
rect 4161 886 4194 5556
rect 4221 949 4254 5705
rect 4284 1010 4317 5877
rect 4497 5390 4521 5401
rect 4791 5390 4822 5401
rect 5224 5386 5253 5402
rect 5370 5350 5389 6650
rect 5798 5346 5823 6749
rect 5968 6745 6041 6749
rect 5984 5706 6001 6745
rect 6484 6692 6581 7417
rect 7746 7315 8065 7427
rect 7023 6955 7170 6961
rect 7023 6913 7027 6955
rect 7162 6913 7170 6955
rect 7023 6908 7170 6913
rect 6786 6694 6830 6697
rect 6482 6690 6583 6692
rect 6482 6649 6485 6690
rect 6580 6649 6583 6690
rect 6482 6645 6583 6649
rect 6786 6647 6830 6650
rect 6206 6298 6240 6301
rect 6206 6272 6211 6298
rect 6237 6272 6240 6298
rect 6211 6269 6237 6272
rect 6023 5945 6049 5948
rect 6023 5916 6049 5919
rect 6026 5693 6045 5916
rect 6213 5691 6234 6269
rect 6570 6209 6596 6210
rect 6568 6207 6598 6209
rect 6568 6181 6570 6207
rect 6596 6181 6598 6207
rect 6568 6179 6598 6181
rect 6570 6178 6596 6179
rect 6253 6105 6287 6108
rect 6253 6079 6257 6105
rect 6283 6079 6287 6105
rect 6253 6076 6287 6079
rect 6260 5693 6279 6076
rect 6297 5896 6326 5899
rect 6297 5870 6299 5896
rect 6325 5870 6326 5896
rect 6297 5867 6326 5870
rect 6301 5691 6322 5867
rect 6401 5848 6435 5851
rect 6401 5822 6405 5848
rect 6431 5822 6435 5848
rect 6401 5819 6435 5822
rect 6409 5694 6427 5819
rect 6573 5155 6593 6178
rect 6796 5689 6819 6647
rect 6886 6299 6914 6302
rect 6886 6273 6887 6299
rect 6913 6273 6914 6299
rect 6886 6270 6914 6273
rect 6842 6208 6870 6211
rect 6842 6182 6843 6208
rect 6869 6182 6870 6208
rect 6842 6179 6870 6182
rect 6571 5142 6593 5155
rect 6566 5139 6599 5142
rect 6566 5112 6569 5139
rect 6596 5112 6599 5139
rect 6566 5109 6599 5112
rect 6819 5098 6820 5114
rect 6845 5025 6867 6179
rect 6844 5018 6867 5025
rect 6843 4958 6863 5018
rect 6888 4973 6911 6270
rect 7025 5670 7067 6908
rect 7128 5670 7170 6908
rect 7366 6690 7410 6693
rect 7366 6643 7410 6646
rect 7376 5945 7399 6643
rect 7818 6118 7946 7315
rect 8194 6796 8222 6808
rect 8194 6793 8227 6796
rect 8194 6749 8199 6793
rect 8194 6746 8227 6749
rect 7818 6110 7948 6118
rect 7817 6109 7948 6110
rect 7817 6083 7821 6109
rect 7943 6083 7948 6109
rect 7817 6080 7948 6083
rect 7495 6044 7525 6047
rect 7495 6018 7497 6044
rect 7523 6018 7525 6044
rect 7495 6015 7525 6018
rect 7363 5944 7399 5945
rect 7360 5942 7399 5944
rect 7360 5860 7366 5942
rect 7392 5860 7399 5942
rect 7360 5855 7399 5860
rect 7376 5689 7399 5855
rect 7498 5689 7521 6015
rect 8126 5990 8169 5994
rect 8126 5964 8130 5990
rect 8156 5964 8169 5990
rect 8126 5960 8169 5964
rect 8150 5693 8169 5960
rect 8194 5684 8222 6746
rect 8364 6299 8390 6302
rect 8364 6270 8390 6273
rect 8275 6212 8301 6215
rect 8275 6183 8301 6186
rect 8278 5811 8297 6183
rect 8366 5811 8388 6270
rect 8563 5948 8597 7570
rect 10603 7318 10922 7430
rect 9013 7224 9050 7225
rect 9008 7220 9058 7224
rect 9008 7183 9016 7220
rect 9053 7183 9058 7220
rect 9008 7179 9058 7183
rect 8628 6371 8660 6375
rect 8628 6344 8631 6371
rect 8657 6344 8660 6371
rect 8628 6338 8660 6344
rect 8558 5942 8597 5948
rect 8558 5940 8561 5942
rect 8557 5863 8561 5940
rect 8593 5863 8597 5942
rect 8558 5856 8597 5863
rect 8261 5791 8329 5811
rect 8261 5765 8275 5791
rect 8301 5765 8329 5791
rect 8261 5742 8329 5765
rect 8365 5792 8433 5811
rect 8365 5766 8377 5792
rect 8403 5766 8433 5792
rect 8365 5742 8433 5766
rect 8563 5678 8597 5856
rect 8630 5800 8657 6338
rect 8630 5797 8698 5800
rect 8630 5754 8652 5797
rect 8695 5754 8698 5797
rect 8630 5750 8698 5754
rect 8630 5685 8657 5750
rect 6844 4955 6867 4958
rect 4487 4349 4511 4786
rect 4781 4342 4812 4793
rect 5224 4344 5253 4791
rect 5370 4395 5389 4785
rect 5501 4405 5524 4789
rect 5798 4406 5823 4791
rect 6845 4635 6867 4955
rect 6845 4626 6880 4635
rect 6845 4604 6896 4626
rect 5368 4345 5389 4395
rect 5499 4364 5524 4405
rect 5796 4364 5823 4406
rect 5974 4421 6002 4532
rect 6027 4463 6046 4523
rect 6227 4479 6266 4481
rect 6226 4476 6266 4479
rect 6226 4470 6233 4476
rect 6211 4469 6233 4470
rect 6027 4444 6187 4463
rect 5974 4393 6146 4421
rect 6126 4370 6146 4393
rect 5368 4332 5387 4345
rect 5499 4321 5522 4364
rect 5796 4327 5821 4364
rect 6127 4340 6143 4370
rect 6168 4332 6187 4444
rect 6208 4448 6233 4469
rect 6261 4448 6266 4476
rect 6208 4445 6266 4448
rect 6208 4443 6265 4445
rect 6208 4442 6227 4443
rect 6208 4358 6225 4442
rect 6675 4436 6698 4527
rect 6797 4439 6820 4527
rect 6623 4429 6698 4436
rect 6620 4413 6698 4429
rect 6795 4433 6820 4439
rect 7128 4446 7170 4546
rect 6620 4368 6661 4413
rect 6208 4331 6224 4358
rect 6620 4319 6658 4368
rect 6795 4333 6819 4433
rect 7128 4428 7171 4446
rect 7128 4389 7172 4428
rect 7376 4407 7399 4527
rect 7131 4368 7172 4389
rect 7131 4317 7171 4368
rect 7375 4333 7399 4407
rect 7498 4438 7521 4527
rect 7498 4400 7574 4438
rect 8150 4425 8169 4523
rect 7536 4354 7574 4400
rect 7967 4417 7995 4420
rect 7967 4391 7968 4417
rect 7994 4391 7995 4417
rect 7967 4388 7995 4391
rect 8010 4406 8169 4425
rect 7970 4340 7986 4388
rect 8010 4373 8029 4406
rect 8194 4387 8222 4532
rect 9013 4488 9050 7179
rect 9092 6874 9138 6877
rect 9092 6837 9098 6874
rect 9135 6837 9138 6874
rect 9092 6834 9138 6837
rect 9010 4483 9055 4488
rect 9010 4446 9017 4483
rect 9054 4446 9055 4483
rect 9010 4442 9055 4446
rect 9013 4438 9050 4442
rect 9094 4429 9131 6834
rect 9169 6403 9214 6406
rect 9169 6366 9175 6403
rect 9212 6366 9214 6403
rect 9169 6363 9214 6366
rect 8055 4386 8222 4387
rect 8007 4362 8029 4373
rect 8007 4332 8026 4362
rect 8051 4359 8222 4386
rect 9091 4424 9135 4429
rect 9091 4387 9094 4424
rect 9131 4387 9135 4424
rect 9091 4383 9135 4387
rect 9094 4378 9131 4383
rect 8051 4340 8067 4359
rect 9171 4194 9208 6363
rect 9826 6311 9884 6314
rect 9826 6261 9830 6311
rect 9880 6261 9884 6311
rect 9826 6258 9884 6261
rect 9708 6251 9764 6255
rect 9600 6204 9656 6208
rect 9505 6155 9561 6166
rect 9505 6105 9508 6155
rect 9558 6105 9561 6155
rect 9505 6101 9561 6105
rect 9600 6154 9603 6204
rect 9653 6154 9656 6204
rect 9708 6201 9711 6251
rect 9761 6201 9764 6251
rect 9708 6196 9764 6201
rect 9600 6150 9656 6154
rect 9258 5896 9301 5899
rect 9258 5859 9263 5896
rect 9300 5859 9301 5896
rect 9258 5855 9301 5859
rect 9168 4193 9208 4194
rect 9167 4191 9209 4193
rect 9167 4154 9168 4191
rect 9205 4154 9209 4191
rect 9167 4151 9209 4154
rect 9171 4150 9208 4151
rect 4487 3687 4511 3773
rect 4781 3687 4812 3780
rect 4487 3396 4521 3687
rect 4781 3396 4822 3687
rect 5224 3396 5253 3778
rect 4497 3372 4521 3396
rect 4791 3369 4822 3396
rect 5370 3369 5389 3778
rect 5501 3674 5524 3782
rect 5492 3670 5525 3674
rect 5492 3629 5496 3670
rect 5522 3629 5525 3670
rect 5492 3626 5525 3629
rect 5501 3365 5524 3626
rect 5798 3386 5823 3784
rect 6130 3380 6146 3785
rect 6405 3421 6429 3793
rect 6403 3396 6442 3421
rect 6417 3371 6442 3396
rect 6623 3358 6661 3807
rect 6798 3419 6822 3793
rect 6798 3392 6845 3419
rect 6818 3369 6845 3392
rect 7026 3356 7066 3809
rect 7378 3542 7402 3793
rect 9259 3676 9296 5855
rect 9255 3670 9304 3676
rect 9255 3629 9261 3670
rect 9298 3629 9304 3670
rect 9255 3625 9304 3629
rect 9259 3622 9296 3625
rect 7378 3518 7436 3542
rect 7412 3384 7436 3518
rect 5933 3283 5965 3287
rect 5933 3257 5936 3283
rect 5962 3257 5965 3283
rect 7924 3281 7950 3284
rect 5933 3253 5965 3257
rect 7923 3255 7924 3278
rect 4487 1533 4511 2796
rect 4781 2688 4812 2803
rect 5224 2739 5253 2801
rect 5274 2770 5308 2773
rect 5274 2744 5278 2770
rect 5304 2744 5308 2770
rect 5274 2741 5308 2744
rect 5221 2736 5256 2739
rect 5221 2707 5224 2736
rect 5253 2707 5256 2736
rect 5221 2704 5256 2707
rect 4777 2687 4814 2688
rect 4777 2656 4780 2687
rect 4811 2656 4814 2687
rect 5224 2658 5253 2704
rect 5274 2680 5299 2741
rect 5370 2682 5389 2802
rect 5798 2735 5823 2808
rect 5941 2777 5962 3253
rect 7923 3252 7950 3255
rect 7872 3188 7898 3191
rect 7872 3159 7898 3162
rect 6067 3084 6106 3109
rect 5995 3005 6029 3008
rect 5995 2979 5999 3005
rect 6025 2979 6029 3005
rect 5995 2974 6029 2979
rect 5999 2972 6021 2974
rect 5938 2774 5966 2777
rect 5938 2748 5939 2774
rect 5965 2748 5966 2774
rect 5938 2745 5966 2748
rect 5999 2744 6019 2972
rect 6045 2790 6064 2826
rect 6041 2773 6069 2790
rect 6041 2747 6042 2773
rect 6068 2747 6069 2773
rect 5995 2741 6023 2744
rect 6041 2743 6069 2747
rect 5795 2733 5829 2735
rect 5795 2707 5799 2733
rect 5825 2707 5829 2733
rect 5995 2715 5996 2741
rect 6022 2715 6023 2741
rect 5995 2712 6023 2715
rect 5795 2706 5829 2707
rect 4777 2655 4814 2656
rect 4781 2534 4812 2655
rect 5167 2630 5253 2658
rect 5159 2629 5253 2630
rect 5269 2669 5299 2680
rect 5364 2679 5396 2682
rect 5159 2627 5205 2629
rect 5159 2585 5161 2627
rect 5203 2585 5205 2627
rect 5159 2582 5205 2585
rect 4776 2531 4818 2534
rect 5269 2518 5288 2669
rect 5364 2653 5367 2679
rect 5393 2653 5396 2679
rect 5364 2650 5396 2653
rect 5632 2629 5707 2648
rect 5657 2545 5707 2629
rect 6088 2621 6106 3084
rect 7825 3004 7851 3007
rect 7825 2975 7851 2978
rect 7775 2911 7801 2914
rect 7775 2882 7801 2885
rect 6220 2737 6246 2740
rect 6218 2735 6248 2737
rect 6218 2709 6220 2735
rect 6246 2709 6248 2735
rect 6218 2707 6248 2709
rect 6220 2706 6246 2707
rect 6088 2617 6136 2621
rect 6088 2591 6100 2617
rect 6096 2584 6100 2591
rect 6133 2584 6136 2617
rect 6221 2614 6243 2706
rect 6417 2693 6442 2816
rect 6818 2695 6845 2818
rect 7100 2775 7143 2778
rect 7100 2740 7104 2775
rect 7139 2740 7143 2775
rect 7100 2738 7143 2740
rect 6416 2667 6419 2693
rect 6445 2667 6448 2693
rect 6818 2691 6853 2695
rect 6818 2664 6823 2691
rect 6850 2664 6853 2691
rect 6096 2580 6136 2584
rect 6215 2611 6249 2614
rect 6215 2574 6249 2577
rect 6221 2566 6243 2574
rect 6616 2547 6710 2640
rect 7104 2595 7139 2738
rect 7286 2682 7308 2814
rect 7412 2742 7435 2814
rect 7412 2719 7733 2742
rect 7412 2718 7435 2719
rect 7104 2563 7108 2595
rect 7134 2563 7139 2595
rect 7104 2559 7139 2563
rect 7257 2658 7308 2682
rect 4776 2486 4818 2489
rect 5225 2512 5288 2518
rect 5608 2513 5632 2545
rect 5732 2513 5756 2545
rect 6589 2515 6613 2547
rect 6713 2515 6737 2547
rect 7257 2533 7280 2658
rect 7710 2622 7733 2719
rect 7705 2619 7736 2622
rect 7705 2585 7707 2619
rect 7733 2585 7736 2619
rect 7705 2582 7736 2585
rect 7246 2530 7292 2533
rect 5225 2480 5229 2512
rect 5261 2486 5288 2512
rect 7246 2492 7250 2530
rect 7288 2492 7292 2530
rect 7246 2489 7292 2492
rect 5261 2480 5269 2486
rect 5225 2476 5269 2480
rect 5608 2379 5632 2411
rect 5732 2378 5756 2410
rect 6589 2381 6613 2413
rect 6713 2380 6737 2412
rect 7710 2265 7733 2582
rect 7697 2243 7733 2265
rect 7677 2220 7733 2243
rect 7677 2219 7731 2220
rect 5246 1958 5278 2133
rect 5608 2102 5632 2134
rect 5732 2101 5756 2133
rect 5632 2036 5658 2082
rect 5706 2038 5732 2082
rect 5631 2033 5659 2036
rect 5631 2002 5659 2005
rect 5705 2035 5733 2038
rect 5705 2004 5733 2007
rect 5234 1948 5288 1958
rect 5234 1902 5239 1948
rect 5285 1902 5288 1948
rect 5234 1898 5288 1902
rect 5632 1861 5658 2002
rect 5706 1861 5732 2004
rect 4447 1516 4512 1533
rect 5632 1518 5732 1861
rect 6083 1856 6117 2135
rect 6077 1853 6123 1856
rect 6077 1804 6123 1807
rect 6226 1767 6260 2134
rect 6589 2104 6613 2136
rect 6713 2104 6737 2136
rect 6613 2036 6639 2085
rect 6612 2033 6640 2036
rect 6612 2002 6640 2005
rect 6613 1884 6639 2002
rect 6687 1884 6713 2085
rect 6217 1764 6269 1767
rect 6217 1718 6220 1764
rect 6266 1718 6269 1764
rect 6217 1715 6269 1718
rect 6613 1524 6713 1884
rect 7068 1679 7095 2138
rect 7775 2098 7800 2882
rect 7825 2188 7850 2975
rect 7873 2279 7898 3159
rect 7923 2368 7948 3252
rect 9507 2518 9557 6101
rect 9600 3046 9650 6150
rect 9713 3569 9763 6196
rect 9826 4086 9876 6258
rect 10712 6098 10840 7318
rect 10711 6095 10840 6098
rect 10839 5967 10840 6095
rect 10711 5964 10840 5967
rect 10712 5915 10840 5964
rect 11148 5797 11168 5800
rect 11139 5794 11170 5797
rect 11139 5751 11143 5794
rect 11169 5751 11170 5794
rect 11139 5747 11170 5751
rect 10757 5665 10792 5668
rect 10757 5623 10760 5665
rect 10786 5623 10792 5665
rect 10757 5620 10792 5623
rect 10358 5343 10405 5349
rect 10358 5303 10360 5343
rect 10400 5303 10405 5343
rect 10358 5300 10405 5303
rect 9821 4083 9876 4086
rect 9871 4033 9876 4083
rect 9821 4030 9876 4033
rect 9712 3561 9764 3569
rect 9712 3514 9713 3561
rect 9763 3514 9764 3561
rect 9712 3513 9764 3514
rect 9599 3045 9651 3046
rect 9599 2995 9600 3045
rect 9650 2995 9651 3045
rect 9599 2994 9651 2995
rect 9491 2515 9557 2518
rect 9491 2465 9495 2515
rect 9545 2465 9557 2515
rect 9491 2461 9557 2465
rect 7918 2364 7955 2368
rect 7918 2314 7922 2364
rect 7948 2314 7955 2364
rect 7918 2310 7955 2314
rect 7865 2274 7902 2279
rect 7865 2224 7868 2274
rect 7894 2224 7902 2274
rect 7865 2221 7902 2224
rect 7816 2184 7853 2188
rect 7816 2134 7821 2184
rect 7847 2134 7853 2184
rect 7816 2130 7853 2134
rect 7769 2094 7804 2098
rect 7057 1673 7106 1679
rect 7057 1627 7059 1673
rect 7105 1627 7106 1673
rect 7057 1623 7106 1627
rect 6613 1520 6815 1524
rect 4447 1404 4452 1516
rect 4478 1404 4512 1516
rect 5584 1514 5777 1518
rect 4447 1401 4512 1404
rect 5530 1512 5777 1514
rect 5530 1510 5663 1512
rect 5530 1398 5589 1510
rect 5775 1400 5777 1512
rect 5701 1398 5777 1400
rect 5530 1395 5777 1398
rect 6565 1514 6815 1520
rect 6565 1395 6570 1514
rect 6756 1395 6815 1514
rect 4282 1008 4319 1010
rect 4282 975 4284 1008
rect 4317 975 4319 1008
rect 4282 972 4319 975
rect 4217 946 4256 949
rect 4217 913 4222 946
rect 4255 913 4256 946
rect 4217 910 4256 913
rect 4157 883 4195 886
rect 4157 850 4159 883
rect 4192 850 4195 883
rect 4157 847 4195 850
rect 4098 820 4133 821
rect 4098 787 4099 820
rect 4132 787 4133 820
rect 4098 784 4133 787
rect 4034 752 4070 754
rect 4034 719 4035 752
rect 4068 719 4070 752
rect 4034 716 4070 719
rect 3975 692 4009 693
rect 3973 690 4011 692
rect 3973 657 3975 690
rect 4008 657 4011 690
rect 3973 655 4011 657
rect 3975 654 4008 655
rect 3915 590 3948 593
rect 3857 533 3890 536
rect 3797 500 3832 503
rect 3797 470 3799 500
rect 3799 464 3832 467
rect 3734 400 3767 403
rect 3670 372 3705 375
rect 3703 342 3705 372
rect 3670 335 3703 338
rect 3511 269 3580 302
rect 3609 311 3653 314
rect 3609 274 3612 311
rect 3649 274 3653 311
rect 3609 272 3653 274
rect 3511 260 3514 269
rect 3456 258 3514 260
rect 5530 246 5624 1395
rect 6565 1392 6815 1395
rect 6726 392 6815 1392
rect 7642 1077 7675 2076
rect 7769 2044 7773 2094
rect 7799 2044 7804 2094
rect 7769 2041 7804 2044
rect 9507 1679 9557 2461
rect 9600 1770 9650 2994
rect 9713 1857 9763 3513
rect 9826 1959 9876 4030
rect 10115 2767 10173 2771
rect 10115 2717 10119 2767
rect 10169 2717 10173 2767
rect 10115 2715 10173 2717
rect 10118 2714 10169 2715
rect 9826 1956 9882 1959
rect 9826 1906 9832 1956
rect 9826 1903 9882 1906
rect 9826 1890 9876 1903
rect 9713 1808 9763 1811
rect 9600 1721 9650 1724
rect 9507 1630 9557 1633
rect 10118 1527 10168 2714
rect 10055 1516 10168 1527
rect 10055 1404 10061 1516
rect 10155 1404 10168 1516
rect 10055 1399 10168 1404
rect 7636 1074 7679 1077
rect 7636 1041 7640 1074
rect 7673 1041 7679 1074
rect 7636 1038 7679 1041
rect 10363 965 10403 5300
rect 10455 5239 10458 5275
rect 10494 5239 10497 5275
rect 10362 962 10409 965
rect 10362 922 10366 962
rect 10406 922 10409 962
rect 10362 919 10409 922
rect 10456 885 10495 5239
rect 10547 5041 10592 5043
rect 10547 5002 10550 5041
rect 10589 5002 10592 5041
rect 10547 5000 10592 5002
rect 10453 881 10499 885
rect 10453 842 10457 881
rect 10496 842 10499 881
rect 10453 838 10499 842
rect 10549 803 10588 5000
rect 10633 4974 10671 4975
rect 10631 4972 10673 4974
rect 10631 4946 10633 4972
rect 10671 4946 10673 4972
rect 10631 4944 10673 4946
rect 10547 799 10594 803
rect 10547 760 10550 799
rect 10589 760 10594 799
rect 10547 757 10594 760
rect 10633 723 10671 4944
rect 10767 2621 10790 5620
rect 11148 5422 11168 5747
rect 11499 5423 11518 7450
rect 11833 6571 11915 6574
rect 11833 6565 11838 6571
rect 11827 6500 11838 6565
rect 11909 6500 11915 6571
rect 11827 6496 11915 6500
rect 11827 4596 11898 6496
rect 11814 4592 11898 4596
rect 11814 4521 11819 4592
rect 11890 4521 11898 4592
rect 11814 4517 11898 4521
rect 11386 2767 11458 2770
rect 11386 2716 11399 2767
rect 11450 2716 11458 2767
rect 11386 2713 11458 2716
rect 10767 2598 10791 2621
rect 10767 2017 10790 2598
rect 11392 2012 11443 2713
rect 11378 2007 11443 2012
rect 11377 1989 11443 2007
rect 11374 1988 11443 1989
rect 11374 1982 11434 1988
rect 11374 1764 11408 1982
rect 11339 1665 11408 1764
rect 11374 1587 11408 1665
rect 11379 1527 11408 1587
rect 11375 1526 11408 1527
rect 11374 1426 11408 1526
rect 11379 1366 11408 1426
rect 11374 1265 11408 1366
rect 11378 1205 11408 1265
rect 11374 1103 11408 1205
rect 11379 1043 11408 1103
rect 11374 942 11408 1043
rect 11378 882 11408 942
rect 10630 719 10674 723
rect 10630 681 10632 719
rect 10670 681 10674 719
rect 11374 695 11408 882
rect 10630 677 10674 681
rect 11378 487 11408 695
rect 11425 1951 11434 1982
rect 11425 487 11432 1951
rect 11378 474 11432 487
rect 6726 319 6818 392
rect 6723 246 6815 319
<< via1 >>
rect 751 7246 790 7285
rect 759 6901 798 6940
rect 897 6784 923 6810
rect 889 6514 931 6556
rect 1484 6374 1513 6432
rect 2813 6268 2839 6294
rect 3392 6225 3423 6256
rect 5050 6989 5092 7031
rect 4665 6913 4707 6955
rect 5217 6752 5261 6796
rect 5789 6752 5833 6796
rect 5971 6749 6015 6793
rect 4775 6650 4819 6694
rect 4499 6348 4525 6374
rect 3792 6279 3818 6305
rect 3675 6180 3702 6206
rect 2542 6102 2577 6137
rect 3067 6133 3093 6159
rect 5346 6650 5390 6694
rect 2644 5878 2670 5917
rect 4284 5879 4317 5905
rect 2580 5796 2606 5836
rect 2582 5685 2608 5711
rect 2205 5643 2231 5669
rect 2202 5551 2228 5577
rect 2203 5459 2229 5485
rect 2138 5357 2164 5383
rect 2134 5261 2160 5287
rect 2138 5165 2164 5191
rect 2582 5593 2608 5619
rect 2579 5501 2605 5527
rect 2134 3637 2160 3684
rect 2198 3637 2224 3684
rect 1998 3534 2024 3560
rect 1946 3494 1972 3520
rect 1018 3369 1084 3435
rect 2206 3532 2232 3558
rect 2382 3533 2409 3560
rect 2140 3496 2166 3522
rect 1948 3103 1974 3129
rect 1539 2917 1576 2954
rect 1022 2783 1088 2849
rect 2432 3494 2458 3520
rect 1538 2293 1575 2330
rect 2292 2251 2318 2287
rect 1837 1727 1866 1756
rect 4221 5707 4254 5740
rect 4164 5559 4197 5592
rect 2643 5392 2669 5418
rect 4100 5399 4133 5432
rect 4036 5342 4069 5375
rect 2644 5296 2670 5322
rect 2643 5200 2669 5226
rect 2579 3434 2605 3460
rect 2517 3319 2543 3345
rect 2475 3058 2501 3084
rect 2519 2489 2545 2531
rect 2515 2251 2541 2287
rect 3975 5185 4008 5218
rect 3912 5032 3945 5065
rect 3856 4875 3889 4908
rect 3794 4328 3827 4361
rect 3731 4169 3764 4202
rect 3669 4014 3702 4047
rect 3609 3866 3642 3899
rect 3545 3349 3578 3382
rect 3478 3192 3511 3225
rect 2643 3001 2669 3027
rect 3416 3028 3449 3061
rect 2577 1888 2603 1921
rect 2474 1726 2503 1755
rect 2358 1625 2418 1685
rect 3348 2884 3381 2917
rect 2944 2448 3002 2519
rect 2636 1132 2662 1166
rect 745 1038 784 1077
rect 3345 501 3388 544
rect 3410 422 3453 465
rect 3477 354 3517 394
rect 3460 260 3511 311
rect 7027 6913 7162 6955
rect 6485 6649 6580 6690
rect 6786 6650 6830 6694
rect 6211 6272 6237 6298
rect 6023 5919 6049 5945
rect 6570 6181 6596 6207
rect 6257 6079 6283 6105
rect 6299 5870 6325 5896
rect 6405 5822 6431 5848
rect 6887 6273 6913 6299
rect 6843 6182 6869 6208
rect 6569 5112 6596 5139
rect 7366 6646 7410 6690
rect 8199 6749 8227 6793
rect 7821 6083 7943 6109
rect 7497 6018 7523 6044
rect 8130 5964 8156 5990
rect 8364 6273 8390 6299
rect 8275 6186 8301 6212
rect 9016 7183 9053 7220
rect 8631 6344 8657 6371
rect 8275 5765 8301 5791
rect 8377 5766 8403 5792
rect 8652 5754 8695 5797
rect 6233 4448 6261 4476
rect 7968 4391 7994 4417
rect 9098 6837 9135 6874
rect 9017 4446 9054 4483
rect 9175 6366 9212 6403
rect 9094 4387 9131 4424
rect 9830 6261 9880 6311
rect 9508 6105 9558 6155
rect 9603 6154 9653 6204
rect 9711 6201 9761 6251
rect 9263 5859 9300 5896
rect 9168 4154 9205 4191
rect 5496 3629 5522 3670
rect 9261 3629 9298 3670
rect 5936 3257 5962 3283
rect 7924 3255 7950 3281
rect 5278 2744 5304 2770
rect 5224 2707 5253 2736
rect 4780 2656 4811 2687
rect 7872 3162 7898 3188
rect 5999 2979 6025 3005
rect 5939 2748 5965 2774
rect 6042 2747 6068 2773
rect 5799 2707 5825 2733
rect 5996 2715 6022 2741
rect 5161 2585 5203 2627
rect 4776 2489 4818 2531
rect 5367 2653 5393 2679
rect 7825 2978 7851 3004
rect 7775 2885 7801 2911
rect 6220 2709 6246 2735
rect 6100 2584 6133 2617
rect 7104 2740 7139 2775
rect 6419 2667 6445 2693
rect 6823 2664 6850 2691
rect 6215 2577 6249 2611
rect 7108 2563 7134 2595
rect 7707 2585 7733 2619
rect 5229 2480 5261 2512
rect 7250 2492 7288 2530
rect 5631 2005 5659 2033
rect 5705 2007 5733 2035
rect 5239 1902 5285 1948
rect 6077 1807 6123 1853
rect 6612 2005 6640 2033
rect 6220 1718 6266 1764
rect 10711 5967 10839 6095
rect 11143 5751 11169 5794
rect 10760 5623 10786 5665
rect 10360 5303 10400 5343
rect 9821 4033 9871 4083
rect 9713 3514 9763 3561
rect 9600 2995 9650 3045
rect 9495 2465 9545 2515
rect 7922 2314 7948 2364
rect 7868 2224 7894 2274
rect 7821 2134 7847 2184
rect 7059 1627 7105 1673
rect 4452 1404 4478 1516
rect 5663 1510 5775 1512
rect 5589 1400 5775 1510
rect 5589 1398 5701 1400
rect 6570 1395 6756 1514
rect 4284 975 4317 1008
rect 4222 913 4255 946
rect 4159 850 4192 883
rect 4099 787 4132 820
rect 4035 719 4068 752
rect 3975 657 4008 690
rect 3915 593 3948 626
rect 3857 536 3890 569
rect 3799 467 3832 500
rect 3734 403 3767 436
rect 3670 338 3703 372
rect 3612 274 3649 311
rect 7773 2044 7799 2094
rect 10119 2717 10169 2767
rect 9832 1906 9882 1956
rect 9713 1811 9763 1857
rect 9600 1724 9650 1770
rect 9507 1633 9557 1679
rect 10061 1404 10155 1516
rect 7640 1041 7673 1074
rect 10458 5239 10494 5275
rect 10366 922 10406 962
rect 10550 5002 10589 5041
rect 10457 842 10496 881
rect 10633 4946 10671 4972
rect 10550 760 10589 799
rect 11838 6500 11909 6571
rect 11819 4521 11890 4592
rect 11399 2716 11450 2767
rect 10632 681 10670 719
<< metal2 >>
rect 625 7277 693 7399
rect 748 7285 793 7287
rect 748 7277 751 7285
rect 625 7254 751 7277
rect 625 7167 693 7254
rect 748 7246 751 7254
rect 790 7246 793 7285
rect 748 7244 793 7246
rect 9010 7220 9056 7222
rect 12097 7220 12183 7355
rect 9010 7183 9016 7220
rect 9053 7183 12183 7220
rect 9010 7181 9056 7183
rect 12097 7145 12183 7183
rect 610 7057 858 7058
rect 610 7018 1005 7057
rect 837 6981 1005 7018
rect 2603 7048 2678 7049
rect 2603 7018 2765 7048
rect 5048 7031 5093 7033
rect 5047 7025 5050 7031
rect 2603 7001 2627 7018
rect 2735 6996 2765 7018
rect 2808 6995 5050 7025
rect 5047 6989 5050 6995
rect 5092 6989 5095 7031
rect 5048 6987 5093 6989
rect 4663 6955 4708 6957
rect 7024 6955 7166 6958
rect 625 6858 693 6946
rect 758 6940 801 6944
rect 758 6901 759 6940
rect 798 6901 801 6940
rect 4662 6913 4665 6955
rect 4707 6954 4710 6955
rect 7024 6954 7027 6955
rect 4707 6914 7027 6954
rect 4707 6913 4710 6914
rect 7024 6913 7027 6914
rect 7162 6954 7166 6955
rect 7162 6914 7171 6954
rect 7162 6913 7166 6914
rect 4663 6911 4708 6913
rect 7024 6910 7166 6913
rect 758 6897 801 6901
rect 758 6896 952 6897
rect 767 6874 952 6896
rect 9093 6874 9137 6876
rect 12097 6874 12183 6942
rect 625 6826 961 6858
rect 9093 6837 9098 6874
rect 9135 6837 12183 6874
rect 9093 6835 9137 6837
rect 625 6714 693 6826
rect 894 6784 897 6810
rect 923 6787 952 6810
rect 923 6784 926 6787
rect 5214 6752 5217 6796
rect 5261 6793 5264 6796
rect 5786 6793 5789 6796
rect 5261 6752 5789 6793
rect 5833 6793 5836 6796
rect 5833 6752 5971 6793
rect 5229 6749 5971 6752
rect 6015 6749 8199 6793
rect 8227 6749 8230 6793
rect 12097 6732 12183 6837
rect 5346 6694 5390 6697
rect 825 6677 978 6693
rect 644 6644 978 6677
rect 4772 6650 4775 6694
rect 4819 6692 4822 6694
rect 4819 6650 5346 6692
rect 6783 6692 6786 6694
rect 5390 6690 6786 6692
rect 5390 6650 6485 6690
rect 4787 6649 6485 6650
rect 6580 6650 6786 6690
rect 6830 6692 6833 6694
rect 6830 6690 7423 6692
rect 6830 6650 7366 6690
rect 6580 6649 7366 6650
rect 4787 6648 7366 6649
rect 5346 6647 5390 6648
rect 7363 6646 7366 6648
rect 7410 6648 7423 6690
rect 7410 6646 7413 6648
rect 644 6637 871 6644
rect 644 6617 684 6637
rect 609 6577 684 6617
rect 11835 6556 11838 6571
rect 886 6514 889 6556
rect 931 6514 11838 6556
rect 11835 6500 11838 6514
rect 11909 6500 11912 6571
rect 580 6432 648 6499
rect 1472 6432 1519 6434
rect 580 6374 1484 6432
rect 1513 6374 1519 6432
rect 9171 6403 9213 6405
rect 12094 6403 12180 6533
rect 580 6350 652 6374
rect 1472 6372 1519 6374
rect 4497 6374 4527 6377
rect 580 6267 648 6350
rect 4497 6348 4499 6374
rect 4525 6371 4527 6374
rect 8629 6371 8659 6374
rect 4525 6348 8631 6371
rect 4497 6345 4527 6348
rect 8629 6344 8631 6348
rect 8657 6348 8666 6371
rect 9171 6366 9175 6403
rect 9212 6366 12180 6403
rect 9171 6364 9213 6366
rect 8657 6344 8659 6348
rect 8629 6340 8659 6344
rect 12094 6323 12180 6366
rect 3789 6305 3820 6307
rect 2810 6297 2842 6298
rect 3789 6297 3792 6305
rect 2810 6294 3792 6297
rect 2810 6268 2813 6294
rect 2839 6279 3792 6294
rect 3818 6297 3821 6305
rect 6207 6298 6239 6300
rect 6884 6299 6916 6300
rect 6207 6297 6211 6298
rect 3818 6279 6211 6297
rect 2839 6274 6211 6279
rect 2839 6268 2842 6274
rect 3789 6273 3820 6274
rect 6207 6272 6211 6274
rect 6237 6297 6240 6298
rect 6884 6297 6887 6299
rect 6237 6274 6887 6297
rect 6237 6272 6240 6274
rect 6884 6273 6887 6274
rect 6913 6297 6916 6299
rect 8361 6297 8364 6299
rect 6913 6274 8364 6297
rect 6913 6273 6916 6274
rect 8361 6273 8364 6274
rect 8390 6297 8393 6299
rect 9827 6297 9830 6311
rect 8390 6274 9830 6297
rect 8390 6273 8393 6274
rect 6884 6272 6916 6273
rect 2810 6266 2842 6268
rect 9827 6261 9830 6274
rect 9880 6261 9883 6311
rect 9827 6260 9883 6261
rect 3389 6256 3426 6258
rect 580 6217 631 6229
rect 3389 6225 3392 6256
rect 3423 6252 3426 6256
rect 9709 6252 9763 6254
rect 3423 6251 9763 6252
rect 3423 6229 9711 6251
rect 3423 6225 3426 6229
rect 3389 6223 3426 6225
rect 580 6188 890 6217
rect 6840 6208 6872 6209
rect 6569 6207 6597 6208
rect 631 6187 890 6188
rect 3672 6206 3703 6207
rect 6567 6206 6570 6207
rect 3672 6180 3675 6206
rect 3702 6183 6570 6206
rect 3702 6180 3705 6183
rect 6567 6181 6570 6183
rect 6596 6206 6599 6207
rect 6840 6206 6843 6208
rect 6596 6183 6843 6206
rect 6596 6181 6599 6183
rect 6840 6182 6843 6183
rect 6869 6206 6872 6208
rect 8272 6206 8275 6212
rect 6869 6186 8275 6206
rect 8301 6206 8304 6212
rect 9601 6206 9655 6207
rect 8301 6204 9655 6206
rect 8301 6186 9603 6204
rect 6869 6183 9603 6186
rect 6869 6182 6872 6183
rect 6840 6181 6872 6182
rect 6569 6180 6597 6181
rect 3672 6178 3703 6180
rect 3064 6160 3096 6161
rect 9507 6160 9560 6163
rect 3064 6159 9560 6160
rect 576 6137 627 6139
rect 2540 6137 2580 6138
rect 576 6102 2542 6137
rect 2577 6102 2580 6137
rect 3064 6133 3067 6159
rect 3093 6155 9560 6159
rect 3093 6137 9508 6155
rect 3093 6133 3096 6137
rect 3064 6131 3096 6133
rect 7819 6109 7947 6112
rect 576 6098 627 6102
rect 2540 6099 2580 6102
rect 6254 6105 6286 6106
rect 6254 6079 6257 6105
rect 6283 6102 6286 6105
rect 7819 6102 7821 6109
rect 6283 6083 7821 6102
rect 7943 6083 7947 6109
rect 9507 6105 9508 6137
rect 9558 6105 9560 6155
rect 9601 6154 9603 6183
rect 9653 6154 9655 6204
rect 9709 6201 9711 6229
rect 9761 6201 9763 6251
rect 9709 6198 9763 6201
rect 9601 6151 9655 6154
rect 9507 6102 9560 6105
rect 6283 6081 7947 6083
rect 6283 6079 6286 6081
rect 6254 6078 6286 6079
rect 548 5917 675 6063
rect 5260 6037 5545 6057
rect 7496 6044 7524 6046
rect 5525 5987 5545 6037
rect 7494 6018 7497 6044
rect 7523 6041 7526 6044
rect 10708 6041 10711 6095
rect 7523 6020 10711 6041
rect 7523 6018 7526 6020
rect 7496 6016 7524 6018
rect 8127 5990 8158 5993
rect 8127 5987 8130 5990
rect 4378 5952 4434 5969
rect 5525 5967 8130 5987
rect 8127 5964 8130 5967
rect 8156 5964 8158 5990
rect 10708 5967 10711 6020
rect 10839 5967 10842 6095
rect 8127 5961 8158 5964
rect 1683 5917 1713 5918
rect 2642 5917 2671 5919
rect 548 5878 2644 5917
rect 2670 5878 2674 5917
rect 4281 5879 4284 5905
rect 4317 5896 4320 5905
rect 4378 5896 4395 5952
rect 6020 5940 6023 5945
rect 5520 5920 6023 5940
rect 4317 5879 4396 5896
rect 5520 5882 5540 5920
rect 6020 5919 6023 5920
rect 6049 5940 6052 5945
rect 6049 5920 6057 5940
rect 6049 5919 6052 5920
rect 6296 5896 6327 5897
rect 9259 5896 9302 5898
rect 12094 5896 12180 6094
rect 6296 5893 6299 5896
rect 548 5875 675 5878
rect 2642 5876 2671 5878
rect 5260 5862 5540 5882
rect 5571 5873 6299 5893
rect 2578 5836 2607 5838
rect 1333 5796 2580 5836
rect 2606 5796 2609 5836
rect 577 5527 704 5614
rect 1333 5527 1373 5796
rect 2578 5795 2607 5796
rect 4378 5769 4434 5786
rect 4221 5742 4254 5743
rect 4219 5740 4256 5742
rect 1713 5728 1750 5729
rect 1534 5705 1750 5728
rect 2579 5706 2582 5711
rect 1534 5692 2276 5705
rect 1534 5622 1596 5692
rect 1713 5688 2276 5692
rect 2522 5689 2582 5706
rect 2579 5685 2582 5689
rect 2608 5706 2611 5711
rect 4219 5707 4221 5740
rect 4254 5732 4256 5740
rect 4378 5732 4395 5769
rect 4254 5715 4395 5732
rect 4254 5707 4256 5715
rect 4378 5714 4395 5715
rect 5571 5707 5591 5873
rect 6296 5870 6299 5873
rect 6325 5870 6328 5896
rect 6296 5869 6327 5870
rect 9259 5859 9263 5896
rect 9300 5884 12180 5896
rect 9300 5859 12169 5884
rect 9259 5856 9300 5859
rect 6402 5848 6434 5849
rect 6402 5845 6405 5848
rect 2608 5689 2617 5706
rect 4219 5704 4256 5707
rect 2608 5685 2611 5689
rect 5260 5687 5591 5707
rect 5626 5825 6405 5845
rect 2202 5643 2205 5669
rect 2231 5664 2234 5669
rect 2231 5647 2276 5664
rect 2231 5643 2234 5647
rect 1713 5622 1750 5626
rect 577 5487 1373 5527
rect 1481 5613 1750 5622
rect 2579 5614 2582 5619
rect 1481 5596 2276 5613
rect 2522 5597 2582 5614
rect 1481 5585 1750 5596
rect 2579 5593 2582 5597
rect 2608 5614 2611 5619
rect 2608 5597 2617 5614
rect 2608 5593 2611 5597
rect 4374 5596 4434 5613
rect 4161 5592 4200 5594
rect 1481 5574 1596 5585
rect 1481 5529 1592 5574
rect 2199 5551 2202 5577
rect 2228 5572 2231 5577
rect 2228 5555 2276 5572
rect 4161 5559 4164 5592
rect 4197 5584 4200 5592
rect 4374 5584 4391 5596
rect 4197 5567 4391 5584
rect 4197 5559 4200 5567
rect 4161 5557 4200 5559
rect 2228 5551 2231 5555
rect 1713 5529 1750 5533
rect 5626 5532 5646 5825
rect 6402 5822 6405 5825
rect 6431 5845 6434 5848
rect 6431 5825 6442 5845
rect 6431 5822 6434 5825
rect 6402 5821 6434 5822
rect 8266 5794 8324 5809
rect 8266 5791 8278 5794
rect 8266 5765 8275 5791
rect 8310 5765 8324 5794
rect 8368 5793 8426 5808
rect 8368 5792 8381 5793
rect 8368 5766 8377 5792
rect 8266 5762 8278 5765
rect 8310 5762 8330 5765
rect 8266 5746 8330 5762
rect 8306 5685 8330 5746
rect 8368 5761 8381 5766
rect 8413 5761 8426 5793
rect 8368 5745 8426 5761
rect 8650 5797 8697 5800
rect 8650 5754 8652 5797
rect 8695 5794 8697 5797
rect 11140 5795 11169 5796
rect 11140 5794 11170 5795
rect 12193 5794 12238 5796
rect 8695 5754 11143 5794
rect 8650 5751 11143 5754
rect 11169 5751 12239 5794
rect 11140 5750 11170 5751
rect 11140 5748 11169 5750
rect 12143 5683 12179 5684
rect 10758 5665 10788 5667
rect 12087 5665 12179 5683
rect 1481 5521 1750 5529
rect 2576 5522 2579 5527
rect 1481 5504 2276 5521
rect 2522 5505 2579 5522
rect 1481 5492 1750 5504
rect 2576 5501 2579 5505
rect 2605 5522 2608 5527
rect 2605 5505 2617 5522
rect 5256 5512 5646 5532
rect 5941 5645 5970 5663
rect 2605 5501 2608 5505
rect 1481 5488 1571 5492
rect 577 5426 704 5487
rect 620 5033 747 5121
rect 1481 5033 1518 5488
rect 2200 5459 2203 5485
rect 2229 5480 2232 5485
rect 2229 5463 2276 5480
rect 2229 5459 2232 5463
rect 4097 5432 4136 5433
rect 1629 5419 2278 5421
rect 620 4996 1518 5033
rect 1600 5402 2278 5419
rect 2640 5415 2643 5418
rect 1600 5384 1750 5402
rect 2519 5395 2643 5415
rect 2640 5392 2643 5395
rect 2669 5415 2672 5418
rect 2669 5395 2682 5415
rect 4097 5399 4100 5432
rect 4133 5424 4136 5432
rect 4391 5424 4434 5441
rect 4133 5407 4454 5424
rect 4133 5399 4136 5407
rect 4391 5405 4408 5407
rect 4097 5398 4136 5399
rect 2669 5392 2672 5395
rect 1600 5325 1666 5384
rect 1713 5380 1750 5384
rect 2135 5357 2138 5383
rect 2164 5379 2167 5383
rect 2164 5360 2278 5379
rect 4033 5375 4072 5378
rect 2164 5357 2167 5360
rect 4033 5342 4036 5375
rect 4069 5367 4072 5375
rect 4069 5350 4454 5367
rect 5941 5361 5959 5645
rect 10757 5623 10760 5665
rect 10786 5655 12179 5665
rect 10786 5623 12183 5655
rect 10758 5621 10788 5623
rect 12087 5589 12183 5623
rect 8376 5447 8436 5458
rect 8376 5413 8389 5447
rect 8423 5413 8436 5447
rect 8736 5441 9259 5464
rect 9296 5441 10211 5464
rect 12093 5446 12183 5589
rect 8376 5402 8436 5413
rect 10182 5431 10211 5441
rect 10980 5431 11094 5439
rect 10182 5419 11094 5431
rect 10182 5411 11015 5419
rect 10182 5410 10211 5411
rect 4069 5342 4072 5350
rect 5864 5344 5959 5361
rect 8737 5359 9259 5381
rect 9296 5359 10117 5381
rect 4033 5340 4072 5342
rect 1600 5306 2278 5325
rect 2641 5319 2644 5322
rect 1600 5288 1750 5306
rect 2519 5299 2644 5319
rect 2641 5296 2644 5299
rect 2670 5319 2673 5322
rect 2670 5299 2682 5319
rect 5298 5301 5318 5313
rect 2670 5296 2673 5299
rect 1600 5287 1667 5288
rect 1600 5283 1666 5287
rect 1713 5284 1750 5288
rect 620 4933 747 4996
rect 614 4557 741 4646
rect 1600 4557 1637 5283
rect 2131 5261 2134 5287
rect 2160 5283 2163 5287
rect 2160 5264 2278 5283
rect 5298 5281 5333 5301
rect 5298 5279 5318 5281
rect 2160 5261 2163 5264
rect 5260 5259 5318 5279
rect 614 4520 1637 4557
rect 1713 5210 2278 5229
rect 2640 5223 2643 5226
rect 614 4458 741 4520
rect 620 4073 747 4164
rect 1713 4073 1750 5210
rect 2519 5203 2643 5223
rect 2640 5200 2643 5203
rect 2669 5223 2672 5226
rect 2669 5203 2682 5223
rect 3972 5218 4011 5220
rect 2669 5200 2672 5203
rect 2135 5165 2138 5191
rect 2164 5187 2167 5191
rect 2164 5168 2278 5187
rect 3972 5185 3975 5218
rect 4008 5210 4011 5218
rect 4008 5193 4454 5210
rect 4008 5185 4011 5193
rect 3972 5183 4011 5185
rect 4399 5177 4434 5193
rect 2164 5165 2167 5168
rect 5293 5159 5330 5179
rect 5293 5104 5313 5159
rect 5897 5156 5970 5174
rect 10095 5171 10117 5359
rect 10357 5343 10403 5346
rect 10357 5303 10360 5343
rect 10400 5333 10403 5343
rect 10988 5333 11094 5341
rect 10400 5321 11094 5333
rect 11530 5321 11702 5341
rect 10400 5313 11015 5321
rect 11530 5313 11701 5321
rect 10400 5303 10403 5313
rect 10357 5301 10403 5303
rect 10458 5275 10494 5278
rect 11681 5268 11701 5313
rect 10494 5248 11094 5268
rect 11530 5248 11701 5268
rect 10458 5236 10494 5239
rect 10095 5170 10255 5171
rect 5897 5135 5915 5156
rect 10095 5150 11094 5170
rect 10095 5149 10255 5150
rect 11681 5143 11701 5248
rect 12090 5143 12180 5210
rect 6567 5140 6598 5141
rect 5858 5117 5915 5135
rect 6566 5139 6599 5140
rect 6566 5134 6569 5139
rect 6531 5129 6569 5134
rect 6208 5112 6569 5129
rect 6596 5112 6599 5139
rect 8814 5113 9259 5129
rect 6208 5107 6598 5112
rect 8811 5109 9259 5113
rect 9296 5119 11015 5129
rect 9296 5109 11094 5119
rect 5260 5084 5313 5104
rect 8270 5100 8326 5109
rect 3909 5065 3951 5066
rect 3909 5032 3912 5065
rect 3945 5057 3951 5065
rect 8270 5065 8282 5100
rect 8315 5065 8326 5100
rect 3945 5040 4399 5057
rect 3945 5032 3951 5040
rect 3909 5031 3951 5032
rect 4382 5022 4399 5040
rect 5907 5041 5962 5059
rect 8270 5055 8326 5065
rect 5907 5039 5925 5041
rect 5865 5023 5925 5039
rect 4382 5005 4434 5022
rect 5296 4948 5328 4992
rect 5296 4929 5316 4948
rect 5260 4909 5316 4929
rect 3853 4908 3892 4909
rect 3853 4875 3856 4908
rect 3889 4900 3892 4908
rect 3889 4883 4390 4900
rect 3889 4875 3892 4883
rect 3853 4874 3892 4875
rect 4374 4872 4390 4883
rect 4374 4842 4391 4872
rect 8811 4861 8834 5109
rect 10985 5099 11094 5109
rect 11681 5100 12180 5143
rect 10550 5042 10589 5044
rect 10549 5041 10590 5042
rect 10549 5002 10550 5041
rect 10589 5031 10590 5041
rect 11681 5031 11701 5100
rect 10589 5021 11015 5031
rect 10589 5011 11094 5021
rect 10589 5002 10590 5011
rect 10549 5001 10590 5002
rect 10992 5001 11094 5011
rect 11530 5001 11701 5031
rect 12090 5001 12180 5100
rect 10550 4999 10589 5001
rect 10632 4972 10672 4973
rect 10630 4946 10633 4972
rect 10671 4966 10674 4972
rect 11681 4966 11701 5001
rect 10671 4948 11015 4966
rect 11530 4948 11701 4966
rect 10671 4946 11094 4948
rect 10632 4945 10672 4946
rect 10980 4928 11094 4946
rect 11524 4934 11701 4948
rect 11524 4928 11700 4934
rect 4374 4825 4434 4842
rect 5289 4836 5327 4854
rect 8374 4844 8436 4853
rect 5289 4754 5307 4836
rect 5863 4791 5935 4809
rect 8374 4808 8391 4844
rect 8425 4808 8436 4844
rect 8736 4838 8834 4861
rect 8895 4848 9259 4868
rect 9296 4850 11015 4868
rect 9296 4848 11094 4850
rect 8374 4800 8436 4808
rect 5260 4734 5308 4754
rect 5917 4572 5935 4791
rect 8895 4778 8915 4848
rect 10989 4830 11094 4848
rect 8737 4763 8915 4778
rect 8737 4756 8912 4763
rect 11816 4592 11894 4595
rect 5917 4554 5971 4572
rect 11816 4521 11819 4592
rect 11890 4580 11894 4592
rect 12090 4580 12180 4672
rect 11890 4533 12180 4580
rect 11890 4521 11894 4533
rect 11816 4518 11894 4521
rect 9012 4483 9058 4485
rect 6231 4478 6263 4479
rect 9012 4478 9017 4483
rect 6231 4476 9017 4478
rect 6231 4448 6233 4476
rect 6261 4450 9017 4476
rect 6261 4448 6263 4450
rect 6231 4445 6263 4448
rect 9012 4446 9017 4450
rect 9054 4446 9058 4483
rect 12090 4463 12180 4533
rect 9012 4444 9058 4446
rect 9091 4424 9134 4426
rect 9091 4418 9094 4424
rect 7965 4417 9094 4418
rect 7965 4391 7968 4417
rect 7994 4392 9094 4417
rect 7994 4391 7997 4392
rect 9091 4387 9094 4392
rect 9131 4387 9134 4424
rect 9091 4385 9134 4387
rect 3792 4361 3829 4365
rect 3792 4328 3794 4361
rect 3827 4353 3829 4361
rect 3827 4336 4424 4353
rect 3827 4328 3829 4336
rect 3792 4325 3829 4328
rect 5909 4312 5927 4313
rect 5875 4301 5927 4312
rect 5875 4294 6110 4301
rect 5909 4283 6110 4294
rect 5267 4246 5327 4266
rect 3728 4202 3767 4203
rect 3728 4169 3731 4202
rect 3764 4194 3767 4202
rect 3764 4182 4424 4194
rect 9165 4191 9209 4193
rect 3764 4177 4434 4182
rect 9165 4181 9168 4191
rect 3764 4169 3767 4177
rect 3728 4168 3767 4169
rect 4395 4165 4434 4177
rect 9152 4163 9168 4181
rect 9164 4154 9168 4163
rect 9205 4154 9209 4191
rect 9164 4153 9209 4154
rect 9164 4147 9204 4153
rect 8081 4129 9204 4147
rect 5287 4126 5325 4127
rect 5285 4109 5325 4126
rect 5285 4091 5305 4109
rect 620 4036 1750 4073
rect 5260 4071 5305 4091
rect 5883 4088 6116 4104
rect 5861 4086 6116 4088
rect 5861 4070 5901 4086
rect 9818 4083 9878 4087
rect 620 3976 747 4036
rect 3666 4014 3669 4047
rect 3702 4039 3705 4047
rect 3702 4022 4384 4039
rect 9818 4033 9821 4083
rect 9871 4081 9878 4083
rect 12090 4081 12180 4184
rect 9871 4034 12180 4081
rect 9871 4033 9878 4034
rect 9818 4029 9878 4033
rect 3702 4014 3705 4022
rect 4369 4015 4384 4022
rect 4369 4004 4386 4015
rect 4369 3987 4434 4004
rect 5863 3991 5903 3992
rect 5863 3977 5904 3991
rect 5863 3976 6114 3977
rect 5886 3959 6114 3976
rect 12090 3975 12180 4034
rect 5280 3931 5325 3944
rect 5280 3916 5329 3931
rect 5260 3911 5329 3916
rect 3605 3899 3647 3900
rect 3605 3866 3609 3899
rect 3642 3891 3647 3899
rect 5260 3896 5315 3911
rect 3642 3874 4386 3891
rect 3642 3866 3647 3874
rect 3605 3864 3647 3866
rect 4369 3825 4386 3874
rect 4369 3808 4434 3825
rect 5284 3789 5327 3812
rect 614 3658 741 3742
rect 5284 3741 5304 3789
rect 5882 3763 6112 3781
rect 5882 3762 5902 3763
rect 5861 3744 5902 3762
rect 5260 3721 5304 3741
rect 2131 3684 2162 3686
rect 2197 3684 2228 3686
rect 614 3621 1584 3658
rect 2131 3637 2134 3684
rect 2160 3637 2198 3684
rect 2224 3637 2863 3684
rect 2131 3635 2162 3637
rect 2197 3635 2228 3637
rect 614 3554 741 3621
rect 1547 3486 1584 3621
rect 2816 3569 2863 3637
rect 5493 3670 5524 3672
rect 9257 3670 9302 3673
rect 5493 3629 5496 3670
rect 5522 3629 9261 3670
rect 9298 3629 9302 3670
rect 5493 3627 5524 3629
rect 9257 3627 9302 3629
rect 12093 3569 12183 3666
rect 1998 3560 2024 3563
rect 2816 3561 12183 3569
rect 2203 3556 2206 3558
rect 2024 3537 2206 3556
rect 1998 3531 2024 3534
rect 2203 3532 2206 3537
rect 2232 3556 2235 3558
rect 2379 3556 2382 3560
rect 2232 3537 2382 3556
rect 2232 3532 2235 3537
rect 2379 3533 2382 3537
rect 2409 3533 2412 3560
rect 2816 3522 9713 3561
rect 1943 3494 1946 3520
rect 1972 3516 1975 3520
rect 2137 3516 2140 3522
rect 1972 3497 2140 3516
rect 1972 3494 1975 3497
rect 2137 3496 2140 3497
rect 2166 3516 2169 3522
rect 2429 3516 2432 3520
rect 2166 3497 2432 3516
rect 2166 3496 2169 3497
rect 2429 3494 2432 3497
rect 2458 3494 2461 3520
rect 9709 3514 9713 3522
rect 9763 3522 12183 3561
rect 9763 3514 9766 3522
rect 9709 3510 9766 3514
rect 1547 3485 1750 3486
rect 1547 3467 1772 3485
rect 1547 3461 1912 3467
rect 1547 3449 2045 3461
rect 2577 3460 2607 3462
rect 2576 3458 2579 3460
rect 1713 3445 2045 3449
rect 1750 3439 2045 3445
rect 1013 3435 1090 3439
rect 1013 3369 1018 3435
rect 1084 3420 1090 3435
rect 2354 3436 2579 3458
rect 1713 3420 1752 3422
rect 1084 3416 1752 3420
rect 1084 3395 2044 3416
rect 1084 3383 1751 3395
rect 2354 3392 2376 3436
rect 2576 3434 2579 3436
rect 2605 3434 2608 3460
rect 12093 3457 12183 3522
rect 2577 3432 2607 3434
rect 4388 3428 4430 3445
rect 4388 3418 4426 3428
rect 4388 3396 4416 3418
rect 1084 3369 1090 3383
rect 1713 3381 1750 3383
rect 3541 3382 3582 3384
rect 1013 3365 1090 3369
rect 3541 3349 3545 3382
rect 3578 3374 3582 3382
rect 4388 3374 4415 3396
rect 3578 3357 4415 3374
rect 5864 3368 5895 3386
rect 3578 3349 3582 3357
rect 4388 3356 4405 3357
rect 3541 3348 3582 3349
rect 2515 3345 2544 3347
rect 2514 3341 2517 3345
rect 620 3255 747 3332
rect 2357 3322 2517 3341
rect 2514 3319 2517 3322
rect 2543 3319 2546 3345
rect 5256 3340 5317 3360
rect 5877 3350 6112 3368
rect 5297 3336 5317 3340
rect 2515 3317 2544 3319
rect 5297 3316 5339 3336
rect 5941 3287 6058 3302
rect 5935 3283 5963 3287
rect 620 3218 1219 3255
rect 4382 3252 4430 3269
rect 5935 3257 5936 3283
rect 5962 3257 5963 3283
rect 7921 3276 7924 3281
rect 7443 3260 7924 3276
rect 5935 3254 5963 3257
rect 7921 3255 7924 3260
rect 7950 3255 7953 3281
rect 620 3144 747 3218
rect 1182 3052 1219 3218
rect 3475 3225 3514 3228
rect 3475 3192 3478 3225
rect 3511 3217 3514 3225
rect 4382 3223 4399 3252
rect 4382 3217 4398 3223
rect 3511 3201 4398 3217
rect 3511 3200 4363 3201
rect 3511 3192 3514 3200
rect 3475 3190 3514 3192
rect 5296 3185 5328 3201
rect 5256 3165 5328 3185
rect 7869 3183 7872 3188
rect 5875 3160 6054 3173
rect 7443 3167 7872 3183
rect 7869 3162 7872 3167
rect 7898 3162 7901 3188
rect 5861 3155 6054 3160
rect 5861 3140 5893 3155
rect 5861 3132 5879 3140
rect 1946 3129 1975 3130
rect 1945 3103 1948 3129
rect 1974 3127 1977 3129
rect 1974 3105 2045 3127
rect 1974 3103 1977 3105
rect 1946 3101 1975 3103
rect 2472 3084 2504 3086
rect 2472 3081 2475 3084
rect 2355 3060 2475 3081
rect 2472 3058 2475 3060
rect 2501 3058 2504 3084
rect 4374 3071 4430 3088
rect 4374 3067 4391 3071
rect 2472 3056 2504 3058
rect 3414 3063 3451 3064
rect 4374 3063 4390 3067
rect 3414 3061 4390 3063
rect 1182 3034 1777 3052
rect 1182 3027 1784 3034
rect 1923 3027 2045 3028
rect 2641 3027 2670 3029
rect 3414 3028 3416 3061
rect 3449 3046 4390 3061
rect 5866 3049 5886 3065
rect 3449 3028 3451 3046
rect 1182 3015 2045 3027
rect 2640 3024 2643 3027
rect 1713 3011 2045 3015
rect 1749 3006 2045 3011
rect 2355 3003 2643 3024
rect 1536 2954 1577 2956
rect 1713 2954 1912 2956
rect 620 2841 747 2923
rect 1536 2917 1539 2954
rect 1576 2950 1912 2954
rect 1576 2928 2045 2950
rect 1576 2917 1751 2928
rect 2355 2921 2376 3003
rect 2640 3001 2643 3003
rect 2669 3001 2672 3027
rect 3414 3025 3451 3028
rect 5868 3044 5886 3049
rect 9597 3045 9652 3046
rect 5868 3026 6057 3044
rect 5256 3008 5325 3010
rect 2641 2999 2670 3001
rect 5256 2990 5333 3008
rect 5304 2981 5333 2990
rect 5996 3005 6028 3007
rect 5996 2979 5999 3005
rect 6025 3003 6028 3005
rect 6025 2982 6057 3003
rect 7822 2999 7825 3004
rect 7443 2983 7825 2999
rect 6025 2979 6042 2982
rect 5996 2975 6042 2979
rect 7822 2978 7825 2983
rect 7851 2978 7854 3004
rect 9597 2995 9600 3045
rect 9650 3043 9653 3045
rect 12090 3043 12180 3158
rect 9650 2996 12180 3043
rect 9650 2995 9653 2996
rect 9597 2993 9652 2995
rect 12090 2949 12180 2996
rect 3345 2917 3384 2919
rect 1536 2915 1577 2917
rect 1713 2915 1750 2917
rect 3345 2884 3348 2917
rect 3381 2909 3384 2917
rect 4365 2909 4430 2916
rect 3381 2899 4430 2909
rect 7772 2906 7775 2911
rect 3381 2892 4394 2899
rect 5302 2893 5332 2897
rect 3381 2884 3384 2892
rect 4377 2890 4394 2892
rect 3345 2882 3384 2884
rect 5301 2869 5332 2893
rect 7443 2890 7775 2906
rect 7772 2885 7775 2890
rect 7801 2885 7804 2911
rect 1013 2849 1093 2855
rect 1013 2841 1022 2849
rect 620 2791 1022 2841
rect 620 2735 747 2791
rect 1013 2783 1022 2791
rect 1088 2783 1093 2849
rect 5301 2835 5321 2869
rect 5892 2835 6055 2848
rect 5256 2815 5321 2835
rect 5861 2830 6055 2835
rect 5861 2817 5910 2830
rect 1013 2778 1093 2783
rect 5936 2774 5968 2775
rect 5275 2744 5278 2770
rect 5304 2765 5307 2770
rect 5936 2765 5939 2774
rect 5304 2749 5939 2765
rect 5304 2744 5307 2749
rect 5936 2748 5939 2749
rect 5965 2748 5968 2774
rect 5936 2747 5968 2748
rect 6039 2773 6071 2794
rect 6039 2747 6042 2773
rect 6068 2763 6071 2773
rect 7101 2775 7142 2776
rect 7101 2765 7104 2775
rect 6404 2763 7104 2765
rect 6068 2749 7104 2763
rect 6068 2747 6071 2749
rect 6039 2746 6071 2747
rect 6396 2742 7104 2749
rect 5995 2741 6023 2742
rect 5222 2736 5255 2738
rect 5221 2707 5224 2736
rect 5253 2728 5256 2736
rect 5796 2733 5828 2734
rect 5796 2728 5799 2733
rect 5253 2712 5799 2728
rect 5253 2707 5256 2712
rect 5796 2707 5799 2712
rect 5825 2707 5828 2733
rect 5993 2732 5996 2741
rect 5990 2716 5996 2732
rect 5993 2715 5996 2716
rect 6022 2732 6025 2741
rect 7101 2740 7104 2742
rect 7139 2740 7142 2775
rect 7101 2739 7142 2740
rect 10116 2767 10172 2769
rect 6217 2732 6220 2735
rect 6022 2716 6220 2732
rect 6022 2715 6025 2716
rect 5995 2714 6023 2715
rect 6217 2709 6220 2716
rect 6246 2709 6249 2735
rect 10116 2717 10119 2767
rect 10169 2762 10172 2767
rect 11388 2767 11456 2768
rect 11388 2762 11399 2767
rect 10169 2721 11399 2762
rect 10169 2717 10172 2721
rect 10116 2716 10172 2717
rect 11388 2716 11399 2721
rect 11450 2762 11456 2767
rect 12141 2762 12207 2826
rect 11450 2721 12207 2762
rect 11450 2716 11456 2721
rect 11388 2715 11456 2716
rect 12141 2711 12207 2721
rect 6219 2708 6247 2709
rect 5221 2705 5256 2707
rect 6418 2693 6446 2696
rect 4779 2687 4812 2690
rect 4779 2656 4780 2687
rect 4811 2666 4812 2687
rect 5365 2679 5395 2680
rect 5364 2666 5367 2679
rect 4811 2656 5367 2666
rect 4779 2653 5367 2656
rect 5393 2666 5396 2679
rect 6418 2667 6419 2693
rect 6445 2667 6446 2693
rect 6418 2666 6446 2667
rect 6821 2691 6851 2694
rect 6821 2666 6823 2691
rect 5393 2664 6823 2666
rect 6850 2664 6851 2691
rect 5393 2661 6850 2664
rect 5393 2653 6844 2661
rect 4779 2650 6844 2653
rect 5160 2628 5204 2629
rect 628 2627 5204 2628
rect 628 2586 5161 2627
rect 4475 2585 4523 2586
rect 5158 2585 5161 2586
rect 5203 2585 5206 2627
rect 6097 2617 6135 2620
rect 7705 2619 7735 2621
rect 5160 2584 5204 2585
rect 6097 2584 6100 2617
rect 6133 2584 6135 2617
rect 6097 2581 6135 2584
rect 6212 2577 6215 2611
rect 6249 2577 6252 2611
rect 7071 2595 7137 2597
rect 7071 2563 7108 2595
rect 7134 2563 7137 2595
rect 7634 2585 7707 2619
rect 7733 2585 7736 2619
rect 7705 2583 7736 2585
rect 7071 2561 7137 2563
rect 626 2489 2519 2531
rect 2545 2519 4776 2531
rect 2545 2489 2944 2519
rect 2931 2448 2944 2489
rect 3002 2489 4776 2519
rect 4818 2489 4824 2531
rect 7246 2530 7291 2532
rect 5227 2512 5265 2515
rect 3002 2448 3014 2489
rect 5227 2480 5229 2512
rect 5261 2480 5265 2512
rect 7246 2492 7250 2530
rect 7288 2492 7291 2530
rect 7246 2489 7291 2492
rect 9492 2515 9552 2518
rect 5227 2477 5265 2480
rect 9492 2465 9495 2515
rect 9545 2513 9552 2515
rect 12133 2513 12343 2607
rect 9545 2466 12343 2513
rect 9545 2465 9552 2466
rect 9492 2462 9552 2465
rect 2931 2439 3014 2448
rect 614 2330 741 2408
rect 12133 2399 12343 2466
rect 12135 2398 12212 2399
rect 1537 2330 1578 2332
rect 614 2293 1538 2330
rect 1575 2293 1578 2330
rect 7919 2314 7922 2364
rect 7948 2314 13573 2364
rect 614 2220 741 2293
rect 1537 2291 1578 2293
rect 2290 2287 2319 2289
rect 2513 2287 2544 2289
rect 2289 2251 2292 2287
rect 2318 2251 2515 2287
rect 2541 2251 2544 2287
rect 12963 2274 13164 2276
rect 2290 2249 2319 2251
rect 2513 2249 2544 2251
rect 7865 2224 7868 2274
rect 7894 2224 13164 2274
rect 7818 2134 7821 2184
rect 7847 2182 12745 2184
rect 7847 2134 12756 2182
rect 7770 2044 7773 2094
rect 7799 2093 12349 2094
rect 7799 2044 12370 2093
rect 5629 2035 6719 2036
rect 5629 2033 5705 2035
rect 5628 2005 5631 2033
rect 5659 2008 5705 2033
rect 5659 2005 5662 2008
rect 5702 2007 5705 2008
rect 5733 2033 6719 2035
rect 5733 2008 6612 2033
rect 5733 2007 5736 2008
rect 6609 2005 6612 2008
rect 6640 2008 6719 2033
rect 6640 2005 6643 2008
rect 1709 1991 1746 1992
rect 620 1909 747 1979
rect 1577 1953 1838 1991
rect 5236 1954 5286 1955
rect 9829 1954 9832 1956
rect 1577 1909 1615 1953
rect 1709 1951 1746 1953
rect 5236 1948 9832 1954
rect 2576 1921 2604 1922
rect 620 1871 1615 1909
rect 2217 1888 2577 1921
rect 2603 1888 2606 1921
rect 5236 1902 5239 1948
rect 5285 1908 9832 1948
rect 5285 1902 5288 1908
rect 9829 1906 9832 1908
rect 9882 1906 9885 1956
rect 5236 1900 5286 1902
rect 2576 1886 2604 1888
rect 620 1791 747 1871
rect 6067 1857 9775 1863
rect 6067 1853 9713 1857
rect 6067 1817 6077 1853
rect 6074 1807 6077 1817
rect 6123 1817 9713 1853
rect 6123 1807 6126 1817
rect 9710 1811 9713 1817
rect 9763 1817 9775 1857
rect 9763 1811 9766 1817
rect 6211 1770 9666 1772
rect 6211 1765 9600 1770
rect 6210 1764 9600 1765
rect 1834 1727 1837 1756
rect 1866 1753 1869 1756
rect 2472 1755 2505 1759
rect 2471 1753 2474 1755
rect 1866 1727 2474 1753
rect 1838 1726 2474 1727
rect 2503 1753 2506 1755
rect 2503 1726 2837 1753
rect 1838 1724 2837 1726
rect 2472 1722 2505 1724
rect 2218 1685 2452 1690
rect 2218 1630 2358 1685
rect 2355 1625 2358 1630
rect 2418 1656 2452 1685
rect 2418 1632 2456 1656
rect 2418 1630 2452 1632
rect 2418 1625 2421 1630
rect 2355 1623 2421 1625
rect 2358 1622 2418 1623
rect 2807 1516 2836 1724
rect 6210 1718 6220 1764
rect 6266 1726 9600 1764
rect 6266 1718 6275 1726
rect 9597 1724 9600 1726
rect 9650 1726 9666 1770
rect 9650 1724 9653 1726
rect 6210 1713 6275 1718
rect 7055 1678 7107 1680
rect 9504 1678 9507 1679
rect 7055 1673 9507 1678
rect 7055 1627 7059 1673
rect 7105 1633 9507 1673
rect 9557 1678 9560 1679
rect 9557 1633 9569 1678
rect 7105 1632 9569 1633
rect 7105 1627 7108 1632
rect 7055 1622 7107 1627
rect 4449 1516 4481 1518
rect 10049 1516 10165 1519
rect 620 1386 747 1477
rect 2788 1404 4452 1516
rect 4478 1514 10061 1516
rect 4478 1512 6570 1514
rect 4478 1510 5663 1512
rect 4478 1404 5589 1510
rect 4449 1402 4481 1404
rect 5586 1398 5589 1404
rect 5775 1404 6570 1512
rect 5775 1400 5778 1404
rect 5701 1398 5778 1400
rect 5586 1396 5778 1398
rect 6567 1395 6570 1404
rect 6756 1404 10061 1514
rect 10155 1404 10165 1516
rect 6756 1395 6760 1404
rect 10049 1401 10165 1404
rect 6567 1393 6760 1395
rect 620 1348 1617 1386
rect 620 1289 747 1348
rect 1579 1263 1617 1348
rect 1709 1263 1746 1264
rect 1579 1225 1851 1263
rect 1709 1223 1746 1225
rect 2634 1166 2665 1168
rect 2211 1132 2636 1166
rect 2662 1132 2665 1166
rect 2634 1130 2665 1132
rect 741 1077 791 1082
rect 741 1038 745 1077
rect 784 1071 791 1077
rect 7638 1074 7677 1075
rect 7637 1071 7640 1074
rect 784 1043 7640 1071
rect 784 1038 791 1043
rect 7637 1041 7640 1043
rect 7673 1041 7677 1074
rect 7638 1040 7677 1041
rect 741 1035 791 1038
rect 4279 1008 4321 1009
rect 4279 975 4284 1008
rect 4317 983 8306 1008
rect 4317 975 8307 983
rect 4279 974 4321 975
rect 7703 973 8307 975
rect 4219 946 4257 947
rect 607 735 734 923
rect 4219 913 4222 946
rect 4255 913 7899 946
rect 4219 912 4257 913
rect 7292 912 7899 913
rect 4155 883 4197 884
rect 4155 850 4159 883
rect 4192 850 7491 883
rect 4155 849 4197 850
rect 4096 820 4136 821
rect 4096 787 4099 820
rect 4132 819 4136 820
rect 4132 787 7090 819
rect 4096 786 7090 787
rect 4096 785 4136 786
rect 4030 752 4071 753
rect 4029 719 4035 752
rect 4068 719 6681 752
rect 4030 717 4071 719
rect 3972 690 4013 691
rect 3972 657 3975 690
rect 4008 688 6279 690
rect 4008 657 6280 688
rect 3972 656 4013 657
rect 3912 593 3915 626
rect 3948 625 3951 626
rect 3948 593 5881 625
rect 3922 592 5881 593
rect 3340 544 3394 547
rect 3340 543 3345 544
rect 2057 539 3345 543
rect 2052 501 3345 539
rect 3388 501 3394 544
rect 3854 536 3857 569
rect 3890 564 3893 569
rect 3890 536 5490 564
rect 3880 531 5490 536
rect 2052 500 3394 501
rect 614 260 741 448
rect 2052 312 2253 500
rect 3340 497 3394 500
rect 3796 467 3799 500
rect 3832 467 5070 500
rect 3405 465 3459 466
rect 3405 459 3410 465
rect 2462 422 3410 459
rect 3453 422 3459 465
rect 4457 437 4659 439
rect 3741 436 4662 437
rect 2462 416 3459 422
rect 2462 315 2660 416
rect 3731 403 3734 436
rect 3767 404 4662 436
rect 3767 403 3770 404
rect 3473 394 3522 398
rect 3473 378 3477 394
rect 2912 376 3477 378
rect 2855 354 3477 376
rect 3517 354 3522 394
rect 2855 348 3522 354
rect 2855 338 3513 348
rect 3667 338 3670 372
rect 3703 338 4265 372
rect 2855 315 3053 338
rect 3456 315 3521 316
rect 2050 246 2253 312
rect 2457 249 2660 315
rect 2853 249 3056 315
rect 3253 311 3521 315
rect 3253 260 3460 311
rect 3511 260 3521 311
rect 3606 313 3661 315
rect 3606 311 3861 313
rect 4062 312 4266 338
rect 3606 274 3612 311
rect 3649 274 3861 311
rect 3606 270 3861 274
rect 3253 252 3521 260
rect 3253 249 3456 252
rect 3658 247 3861 270
rect 4061 246 4266 312
rect 4454 249 4662 404
rect 4865 337 5068 467
rect 4865 308 5069 337
rect 4866 247 5069 308
rect 5283 249 5486 531
rect 5682 321 5881 592
rect 5681 246 5884 321
rect 6080 319 6280 657
rect 6077 249 6280 319
rect 6490 312 6681 719
rect 6894 314 7089 786
rect 7292 314 7491 850
rect 7703 880 7899 912
rect 8113 923 8307 973
rect 10365 962 10408 964
rect 8515 959 8711 962
rect 10363 959 10366 962
rect 8515 924 10366 959
rect 7703 314 7898 880
rect 8113 316 8306 923
rect 6482 247 6685 312
rect 6889 249 7092 314
rect 7292 249 7495 314
rect 7697 249 7900 314
rect 8104 238 8307 316
rect 8515 314 8711 924
rect 10363 922 10366 924
rect 10406 922 10409 962
rect 10365 921 10408 922
rect 10455 881 10498 883
rect 10454 880 10457 881
rect 8908 842 10457 880
rect 10496 842 10499 881
rect 8512 249 8715 314
rect 8908 312 9104 842
rect 10455 840 10498 842
rect 10547 798 10550 799
rect 9323 760 10550 798
rect 10589 760 10592 799
rect 9323 314 9521 760
rect 10631 719 10673 722
rect 9734 681 10632 719
rect 10670 681 10673 719
rect 8907 247 9110 312
rect 9319 249 9522 314
rect 9734 311 9932 681
rect 10631 678 10673 681
rect 10241 382 10865 402
rect 10241 314 10261 382
rect 10957 361 10977 402
rect 10734 341 10977 361
rect 10734 314 10754 341
rect 11054 314 11075 403
rect 9733 246 9936 311
rect 10132 249 10335 314
rect 10534 284 10754 314
rect 10534 249 10737 284
rect 10942 249 11145 314
rect 11247 305 11268 403
rect 11344 384 11363 401
rect 11344 365 11844 384
rect 11825 319 11844 365
rect 11360 305 11563 314
rect 11825 312 11928 319
rect 12169 314 12370 2044
rect 11247 284 11563 305
rect 11360 249 11563 284
rect 11758 247 11961 312
rect 12163 262 12370 314
rect 12555 314 12756 2134
rect 12163 249 12366 262
rect 12555 249 12762 314
rect 12963 312 13164 2224
rect 13372 314 13573 2314
rect 12555 245 12756 249
rect 12963 247 13167 312
rect 13369 256 13573 314
rect 13369 249 13572 256
rect 12963 239 13164 247
<< via2 >>
rect 8278 5791 8310 5794
rect 8278 5765 8301 5791
rect 8301 5765 8310 5791
rect 8381 5792 8413 5793
rect 8381 5766 8403 5792
rect 8403 5766 8413 5792
rect 8278 5762 8310 5765
rect 8381 5761 8413 5766
rect 8389 5413 8423 5447
rect 8282 5065 8315 5100
rect 8391 4808 8425 4844
<< metal3 >>
rect 8271 5794 8316 5800
rect 8271 5762 8278 5794
rect 8310 5762 8316 5794
rect 8271 5725 8316 5762
rect 8375 5793 8420 5799
rect 8375 5761 8381 5793
rect 8413 5761 8420 5793
rect 8271 5109 8308 5725
rect 8375 5724 8420 5761
rect 8383 5460 8420 5724
rect 8383 5447 8427 5460
rect 8383 5413 8389 5447
rect 8423 5413 8427 5447
rect 8383 5400 8427 5413
rect 8271 5100 8320 5109
rect 8271 5076 8282 5100
rect 8276 5065 8282 5076
rect 8315 5065 8320 5100
rect 8276 5060 8320 5065
rect 8383 4889 8420 5400
rect 8382 4844 8429 4889
rect 8382 4808 8391 4844
rect 8425 4808 8429 4844
rect 8382 4802 8429 4808
use sky130_hilas_nFETLarge  sky130_hilas_nFETLarge_0
timestamp 1628616966
transform -1 0 2338 0 -1 2867
box 0 0 557 603
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_0
timestamp 1628616754
transform -1 0 2342 0 -1 2112
box 0 0 464 599
use sky130_hilas_nFETLarge  sky130_hilas_nFETLarge_1
timestamp 1628616966
transform -1 0 7765 0 1 1639
box 0 0 557 603
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_1
timestamp 1628616754
transform 1 0 5154 0 1 1637
box 0 0 464 599
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_2
timestamp 1628616754
transform -1 0 6210 0 1 1637
box 0 0 464 599
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_3
timestamp 1628616754
transform 1 0 6135 0 1 1640
box 0 0 464 599
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_4
timestamp 1628616754
transform -1 0 7191 0 1 1640
box 0 0 464 599
use sky130_hilas_DAC5bit01  sky130_hilas_DAC5bit01_0
timestamp 1628616972
transform 0 1 10242 1 0 0
box 0 0 1658 799
use sky130_hilas_Trans2med  sky130_hilas_Trans2med_0
timestamp 1628616970
transform 1 0 2403 0 -1 3342
box 0 0 440 593
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_2
timestamp 1628616740
transform -1 0 5257 0 -1 4271
box 0 0 889 787
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_3
timestamp 1628616740
transform -1 0 5253 0 -1 3365
box 0 0 889 787
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_1
timestamp 1628616740
transform -1 0 5257 0 -1 5284
box 0 0 889 787
use sky130_hilas_WTA4Stage01  sky130_hilas_WTA4Stage01_0
timestamp 1628616963
transform 1 0 7155 0 1 2835
box 0 0 2692 1487
use sky130_hilas_swc4x2cell  sky130_hilas_swc4x2cell_0
timestamp 1628616697
transform 1 0 7095 0 1 3733
box 0 0 4572 1472
use sky130_hilas_TA2Cell_1FG  sky130_hilas_TA2Cell_1FG_0
timestamp 1628616976
transform 1 0 8566 0 1 4364
box 0 0 4090 2332
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_3
timestamp 1628616972
transform -1 0 6932 0 -1 3402
box 0 0 800 611
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_2
timestamp 1628616972
transform -1 0 6929 0 -1 4329
box 0 0 800 611
use sky130_hilas_Trans4small  sky130_hilas_Trans4small_0
timestamp 1628616972
transform 1 0 2068 0 1 5290
box 0 0 340 646
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_0
timestamp 1628616740
transform -1 0 5257 0 1 5507
box 0 0 889 787
use sky130_hilas_FGcharacterization01  sky130_hilas_FGcharacterization01_0
timestamp 1628616982
transform -1 0 3012 0 1 6339
box 0 0 3012 1417
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_1
timestamp 1628616972
transform -1 0 6931 0 -1 5376
box 0 0 800 611
use sky130_hilas_TA2Cell_1FG_Strong  sky130_hilas_TA2Cell_1FG_Strong_0
timestamp 1628616985
transform 1 0 8566 0 1 4967
box 0 0 4694 2332
use sky130_hilas_Tgate4Single01  sky130_hilas_Tgate4Single01_0
timestamp 1628616972
transform 1 0 11110 0 1 4978
box 0 0 739 1047
<< labels >>
rlabel metal2 13369 249 13572 314 1 DIG24 
port 1 n
rlabel metal2 12964 247 13167 312 0 DIG23
port 2 nsew
rlabel metal2 12559 249 12762 314 0 DIG22
port 3 nsew
rlabel metal2 12163 249 12366 314 0 DIG21
port 4 nsew
rlabel metal2 11758 247 11961 312 0 DIG29
port 5 nsew
rlabel metal2 11360 249 11563 314 0 DIG28
port 6 nsew
rlabel metal2 10942 249 11145 314 0 DIG27
port 7 nsew
rlabel metal2 10534 249 10737 314 0 DIG26
port 8 nsew
rlabel metal2 10132 249 10335 314 0 DIG25
port 9 nsew
rlabel metal2 9733 246 9936 311 0 DIG20
port 10 nsew
rlabel metal2 9319 249 9522 314 0 DIG19
port 11 nsew
rlabel metal2 8907 247 9110 312 0 DIG18
port 12 nsew
rlabel metal2 8512 249 8715 314 0 DIG17
port 13 nsew
rlabel metal2 8104 251 8307 316 0 DIG16
port 14 nsew
rlabel metal2 7697 249 7900 314 0 DIG15
port 15 nsew
rlabel metal2 7292 249 7495 314 0 DIG14
port 16 nsew
rlabel metal2 6889 249 7092 314 0 DIG13
port 17 nsew
rlabel metal2 6482 247 6685 312 0 DIG12
port 18 nsew
rlabel metal2 6077 253 6280 319 0 DIG11
port 19 nsew
rlabel metal2 5681 255 5884 321 0 DIG10
port 20 nsew
rlabel metal2 5283 249 5486 315 0 DIG09
port 21 nsew
rlabel metal2 4866 247 5069 313 0 DIG08
port 22 nsew
rlabel metal2 4457 249 4660 315 0 DIG07
port 23 nsew
rlabel metal2 4061 246 4264 312 0 DIG06
port 24 nsew
rlabel metal2 3658 247 3861 313 0 DIG05
port 25 nsew
rlabel metal2 3253 249 3456 315 0 DIG04
port 26 nsew
rlabel metal2 2853 249 3056 315 0 DIG03
port 27 nsew
rlabel metal2 2457 249 2660 315 0 DIG02
port 28 nsew
rlabel metal2 2050 246 2253 312 0 DIG01
port 29 nsew
rlabel metal2 12135 2398 12212 2607 0 CAP2    
port 30 nsew
rlabel metal2 12090 2949 12180 3158 0 GENERALGATE01   
port 31 nsew
rlabel metal2 12093 3457 12183 3666 0 GATEANDCAP1    
port 32 nsew
rlabel metal2 12090 3975 12180 4184 0 GENERALGATE02
port 33 nsew
rlabel metal2 12090 4463 12180 4672 0 OUTPUTTA1    
port 34 nsew
rlabel metal2 12090 5001 12180 5210 0 GATENFET1   
port 35 nsew
rlabel metal2 12093 5446 12183 5655 0 DACOUTPUT  
port 36 nsew
rlabel metal2 12094 5884 12180 6094 0 DRAINOUT
port 37 nsew
rlabel metal2 12094 6323 12180 6533 0 ROWTERM2
port 38 nsew
rlabel metal2 12097 6732 12183 6942 0 COLUMN2
port 39 nsew
rlabel metal2 12097 7145 12183 7355 0 COLUMN1
port 40 nsew
rlabel metal1 10603 7318 10922 7430 0 GATE2
port 41 nsew
rlabel metal1 7746 7315 8065 7427 0 GATE1
port 61 nsew
rlabel metal1 4887 7316 5206 7428 0 DRAININJECT
port 42 nsew
rlabel metal1 3356 7269 3490 7370 0 VTUN
port 43 nsew
rlabel metal2 625 7167 693 7399 0 VREFCHAR
port 44 nsew
rlabel metal2 625 6714 693 6946 0 CHAROUTPUT
port 45 nsew
rlabel metal2 580 6267 648 6499 0 LARGECAPACITOR
port 46 nsew
rlabel metal2 1709 1951 1746 1992 0 DRAIN6N
port 47 nsew
rlabel metal2 1709 1223 1746 1264 0 DRAIN6P
port 48 nsew
rlabel metal2 1713 2915 1750 2956 0 DRAIN5P
port 49 nsew
rlabel metal2 1713 3011 1750 3052 0 DARIN4P
port 50 nsew
rlabel metal2 1713 3381 1750 3422 0 DRAIN5N
port 51 nsew
rlabel metal2 1713 3445 1750 3486 0 DRAIN4N
port 52 nsew
rlabel metal2 1713 5188 1750 5229 0 DRAIN3P
port 53 nsew
rlabel metal2 1713 5284 1750 5325 0 DRAIN2P
port 54 nsew
rlabel metal2 1713 5380 1750 5421 0 DRAIN1P
port 55 nsew
rlabel metal2 1713 5492 1750 5533 0 DRAIN3N
port 56 nsew
rlabel metal2 1713 5585 1750 5626 0 DRAIN2N
port 57 nsew
rlabel metal2 1713 5688 1750 5729 0 DRAIN1N
port 58 nsew
rlabel metal2 1683 5796 1713 5836 0 SOURCEN
port 59 nsew
rlabel metal2 1683 5878 1713 5918 0 SOURCEP
port 60 nsew
rlabel metal2 609 6577 654 6617 0 VGND
port 63 nsew
rlabel metal2 613 7018 658 7058 0 VINJ
port 62 nsew
rlabel metal2 580 6188 631 6229 0 VINJ
port 62 nsew
rlabel metal2 576 6098 627 6139 0 VGND
port 63 nsew
rlabel metal2 628 2586 691 2628 0 VINJ
port 62 nsew
rlabel metal2 626 2489 689 2531 0 VGND
port 63 nsew
rlabel metal2 12193 5751 12238 5796 0 VPWR
port 64 nsew
rlabel metal1 5968 7402 6041 7432 0 VINJ
port 62 nsew
rlabel metal1 6484 7411 6581 7432 0 VGND
port 63 nsew
rlabel metal2 12141 2711 12207 2826 0 VPWR
port 64 nsew
rlabel metal1 5530 246 5622 319 0 VPWR
port 64 nsew
rlabel metal1 6723 246 6815 319 0 VPWR
port 64 nsew
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
