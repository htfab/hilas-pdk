magic
tech sky130A
timestamp 1629472382
<< checkpaint >>
rect -630 -248 5202 2102
rect 33 -252 4539 -248
rect 102 -257 4470 -252
rect 650 -652 3922 -257
<< error_s >>
rect 1347 594 1397 600
rect 1419 594 1469 600
rect 3103 594 3153 600
rect 3175 594 3225 600
rect 1347 552 1397 558
rect 1419 552 1469 558
rect 3103 552 3153 558
rect 3175 552 3225 558
rect 1419 525 1469 531
rect 3103 525 3153 531
rect 1419 483 1469 489
rect 3103 483 3153 489
rect 1419 440 1469 446
rect 3103 440 3153 446
rect 1419 398 1469 404
rect 3103 398 3153 404
rect 1347 371 1397 377
rect 1419 371 1469 377
rect 3103 371 3153 377
rect 3175 371 3225 377
rect 1347 329 1397 335
rect 1419 329 1469 335
rect 3103 329 3153 335
rect 3175 329 3225 335
rect 1347 270 1397 276
rect 1419 270 1469 276
rect 3103 270 3153 276
rect 3175 270 3225 276
rect 1347 228 1397 234
rect 1419 228 1469 234
rect 3103 228 3153 234
rect 3175 228 3225 234
rect 1419 201 1469 207
rect 3103 201 3153 207
rect 1419 159 1469 165
rect 3103 159 3153 165
rect 1419 117 1469 123
rect 3103 117 3153 123
rect 1419 75 1469 81
rect 3103 75 3153 81
rect 1347 48 1397 54
rect 1419 48 1469 54
rect 3103 48 3153 54
rect 3175 48 3225 54
rect 1347 6 1397 12
rect 1419 6 1469 12
rect 3103 6 3153 12
rect 3175 6 3225 12
<< nwell >>
rect 3264 587 3273 617
rect 1280 369 1293 375
rect 1280 357 1287 369
<< metal1 >>
rect 3241 615 3273 616
rect 1301 614 1332 615
rect 1301 601 1304 614
rect 1300 588 1304 601
rect 1330 588 1332 614
rect 3241 605 3244 615
rect 1357 600 1376 605
rect 1397 600 1413 605
rect 1591 596 1615 605
rect 1809 595 1847 605
rect 1984 599 2008 605
rect 2212 592 2252 605
rect 2320 595 2360 605
rect 2564 600 2588 605
rect 2725 595 2763 605
rect 2957 598 2981 605
rect 3159 600 3175 605
rect 3196 600 3215 605
rect 1300 586 1332 588
rect 1316 571 1332 586
rect 2252 569 2320 591
rect 3240 589 3244 605
rect 3270 589 3273 615
rect 3240 588 3273 589
rect 3240 571 3256 588
rect 1316 0 1332 6
rect 1357 1 1376 7
rect 1397 1 1413 7
rect 1591 0 1615 8
rect 1809 0 1847 9
rect 1984 0 2008 7
rect 2212 0 2252 12
rect 2320 0 2360 12
rect 2564 0 2588 7
rect 2725 0 2763 15
rect 2957 0 2981 6
rect 3159 1 3175 7
rect 3196 1 3215 7
rect 3240 1 3256 7
<< via1 >>
rect 1304 588 1330 614
rect 3244 589 3270 615
<< metal2 >>
rect 1300 615 3274 618
rect 1300 614 3244 615
rect 1300 588 1304 614
rect 1330 600 3244 614
rect 1330 588 1342 600
rect 1300 586 1342 588
rect 3240 589 3244 600
rect 3270 589 3274 615
rect 3240 587 3274 589
rect 1280 554 1286 572
rect 3283 554 3292 572
rect 1280 511 1287 529
rect 3283 511 3292 529
rect 1280 400 1286 418
rect 3286 400 3292 418
rect 1280 357 1293 375
rect 3286 357 3292 375
rect 1280 230 1287 248
rect 3283 230 3292 248
rect 1280 187 1287 205
rect 3283 187 3292 205
rect 1950 138 2626 156
rect 1280 77 1287 95
rect 3283 77 3292 95
rect 1280 34 1287 52
rect 3283 34 3292 52
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_0
timestamp 1629137274
transform 1 0 2548 0 1 382
box 0 0 2024 1090
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_1
timestamp 1629137274
transform -1 0 2024 0 1 382
box 0 0 2024 1090
<< labels >>
rlabel metal1 2725 595 2763 605 0 GATE2
port 1 nsew analog default
rlabel metal1 2212 0 2252 12 0 VTUN
port 2 nsew power default
rlabel metal1 2320 0 2360 12 0 VTUN
port 2 nsew power default
rlabel metal1 2320 595 2360 605 0 VTUN
port 2 nsew power default
rlabel metal1 2212 592 2252 605 0 VTUN
port 2 nsew power default
rlabel metal1 1809 595 1847 605 0 GATE1
port 3 nsew analog default
rlabel metal1 1809 0 1847 9 0 GATE1
port 3 nsew analog default
rlabel metal1 3240 1 3256 7 0 VINJ
port 4 nsew power default
rlabel metal1 2725 0 2763 15 0 GATE2
port 1 nsew analog default
rlabel metal1 3196 600 3215 605 0 SelectGate2
rlabel metal1 3240 600 3256 605 0 VINJ
port 6 nsew power default
rlabel metal1 1316 600 1332 605 0 VINJ
port 6 nsew power default
rlabel metal1 1357 600 1376 605 0 GATESELECT1
port 10 nsew analog default
rlabel metal1 1316 0 1332 6 0 VINJ
port 6 nsew power default
rlabel metal1 1357 1 1376 7 0 GATESELECT1
port 10 nsew analog default
rlabel metal1 1397 600 1413 605 0 COL1
port 12 nsew analog default
rlabel metal1 1397 1 1413 7 0 COL1
port 12 nsew analog default
rlabel metal1 3196 1 3215 7 0 GATESELECT2
port 11 nsew analog default
rlabel metal1 3159 1 3175 7 0 COL2
port 13 nsew analog default
rlabel metal1 3159 600 3175 605 0 COL2
port 13 nsew analog default
rlabel metal1 1591 599 1615 605 0 VGND
port 22 nsew
rlabel metal1 1591 0 1615 8 0 VGND
port 22 nsew
rlabel metal1 1984 0 2008 7 0 VGND
port 22 nsew
rlabel metal1 1984 599 2008 605 0 VGND
port 22 nsew
rlabel metal1 2564 0 2588 7 0 VGND
port 22 nsew
rlabel metal1 2957 0 2981 6 0 VGND
port 22 nsew
rlabel metal1 2564 600 2588 605 0 VGND
port 22 nsew
rlabel metal1 2957 598 2981 605 0 VGND
port 22 nsew
rlabel metal2 1280 34 1287 52 0 DRAIN4
port 21 nsew
rlabel metal2 1280 77 1287 95 0 ROW4
port 20 nsew
rlabel metal2 1280 187 1287 205 0 ROW3
port 19 nsew
rlabel metal2 1280 230 1287 248 0 DRAIN3
port 18 nsew
rlabel metal2 1280 357 1287 375 0 DRAIN2
port 17 nsew
rlabel metal2 1280 400 1286 418 0 ROW2
port 15 nsew
rlabel metal2 1280 511 1287 529 0 ROW1
port 14 nsew
rlabel metal2 1280 554 1286 572 0 DRAIN1
port 16 nsew
rlabel metal2 3283 511 3292 529 0 ROW1
port 14 nsew
rlabel metal2 3286 400 3292 418 0 ROW2
port 15 nsew
rlabel metal2 3286 357 3292 375 0 DRAIN2
port 17 nsew
rlabel metal2 3283 230 3292 248 0 DRAIN3
port 18 nsew
rlabel metal2 3283 187 3292 205 0 ROW3
port 19 nsew
rlabel metal2 3283 77 3292 95 0 ROW4
port 20 nsew
rlabel metal2 3283 34 3292 52 0 DRAIN4
port 21 nsew
rlabel metal2 3283 554 3292 572 0 DRAIN1
port 16 nsew
<< end >>
