VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_overlapcap01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_overlapcap01 ;
  ORIGIN 2.870 0.710 ;
  SIZE 2.870 BY 2.080 ;
  OBS
      LAYER nwell ;
        RECT -2.810 -0.650 -0.090 1.310 ;
      LAYER li1 ;
        RECT -2.410 -0.260 -0.460 0.910 ;
      LAYER mcon ;
        RECT -1.930 0.570 -1.760 0.740 ;
        RECT -1.930 0.230 -1.760 0.400 ;
        RECT -1.930 -0.110 -1.760 0.060 ;
      LAYER met1 ;
        RECT -1.970 0.320 -1.710 0.800 ;
        RECT -1.980 -0.200 -1.710 0.320 ;
        RECT -1.980 -0.650 -1.720 -0.200 ;
  END
END sky130_hilas_overlapcap01
END LIBRARY

