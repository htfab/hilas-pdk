VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_hilas_TA2Cell_1FG_Strong
  CLASS CORE ;
  FOREIGN sky130_hilas_TA2Cell_1FG_Strong ;
  ORIGIN 0.000 0.000 ;
  SIZE 46.940 BY 23.320 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 25.760 14.880 26.180 15.030 ;
        RECT 26.790 14.880 27.210 15.030 ;
        RECT 25.760 14.740 27.210 14.880 ;
    END
  END VTUN
  PIN PROG
    PORT
      LAYER met1 ;
        RECT 18.520 14.970 18.730 15.030 ;
    END
  END PROG
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT 30.490 14.950 30.720 15.030 ;
    END
  END GATE1
  PIN VIN11
    PORT
      LAYER met1 ;
        RECT 17.640 14.920 17.850 15.030 ;
    END
  END VIN11
  PIN VINJ
    PORT
      LAYER met2 ;
        RECT 15.200 14.890 15.520 15.010 ;
        RECT 37.470 14.890 37.790 15.010 ;
        RECT 15.200 14.710 37.790 14.890 ;
    END
    PORT
      LAYER met1 ;
        RECT 37.450 15.010 37.730 15.030 ;
        RECT 37.450 14.950 37.790 15.010 ;
        RECT 37.470 14.710 37.790 14.950 ;
      LAYER via ;
        RECT 37.500 14.730 37.760 14.990 ;
    END
    PORT
      LAYER met1 ;
        RECT 37.450 8.980 37.730 9.030 ;
    END
  END VINJ
  PIN VIN22
    PORT
      LAYER met2 ;
        RECT 38.570 14.760 38.880 15.000 ;
    END
  END VIN22
  PIN VIN21
    PORT
      LAYER met2 ;
        RECT 38.650 12.090 38.970 12.330 ;
    END
  END VIN21
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 41.800 14.880 42.080 15.030 ;
    END
    PORT
      LAYER met1 ;
        RECT 41.810 8.980 42.080 9.190 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 41.570 16.460 41.890 16.540 ;
        RECT 40.580 16.280 41.890 16.460 ;
        RECT 40.580 16.110 41.760 16.280 ;
        RECT 40.630 15.960 40.950 16.110 ;
    END
    PORT
      LAYER met2 ;
        RECT 39.610 9.330 39.930 9.480 ;
        RECT 23.420 9.180 39.930 9.330 ;
        RECT 23.420 9.030 23.740 9.180 ;
        RECT 29.220 9.030 29.540 9.180 ;
    END
  END VGND
  PIN OUTPUT2
    PORT
      LAYER met2 ;
        RECT 42.990 11.500 43.100 11.720 ;
    END
  END OUTPUT2
  PIN OUTPUT1
    PORT
      LAYER met2 ;
        RECT 42.990 12.320 43.100 12.550 ;
    END
  END OUTPUT1
  PIN GATESEL1
    PORT
      LAYER met1 ;
        RECT 15.520 15.030 15.940 19.320 ;
        RECT 15.360 15.010 15.960 15.030 ;
        RECT 15.200 14.970 15.960 15.010 ;
        RECT 15.200 14.710 15.940 14.970 ;
        RECT 15.520 13.270 15.940 14.710 ;
      LAYER via ;
        RECT 15.230 14.730 15.490 14.990 ;
    END
  END GATESEL1
  PIN GATESEL2
    PORT
      LAYER met1 ;
        RECT 37.010 8.980 37.200 9.030 ;
    END
    PORT
      LAYER met1 ;
        RECT 37.010 14.950 37.200 15.030 ;
    END
  END GATESEL2
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 15.000 14.350 15.080 14.530 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 15.000 9.480 15.080 9.660 ;
    END
  END DRAIN2
  PIN VIN12
    PORT
      LAYER met1 ;
        RECT 17.650 8.990 17.880 9.110 ;
    END
  END VIN12
  PIN GATE2
    PORT
      LAYER met1 ;
        RECT 18.110 14.950 18.300 15.030 ;
    END
  END GATE2
  PIN RUN
    PORT
      LAYER met1 ;
        RECT 19.600 14.960 19.780 15.030 ;
    END
  END RUN
  OBS
      LAYER nwell ;
        RECT 0.040 22.980 1.770 23.320 ;
        RECT 44.920 22.980 46.650 23.320 ;
        RECT 0.040 21.420 1.790 22.980 ;
        RECT 0.060 19.790 1.790 21.420 ;
        RECT 44.900 21.420 46.650 22.980 ;
        RECT 44.900 19.790 46.630 21.420 ;
        RECT 0.000 16.620 3.310 19.790 ;
        RECT 43.380 19.400 46.690 19.790 ;
        RECT 19.850 19.360 22.560 19.400 ;
        RECT 43.380 19.360 46.930 19.400 ;
        RECT 19.850 17.710 22.570 19.360 ;
        RECT 38.620 19.310 41.930 19.320 ;
        RECT 40.970 19.280 41.160 19.310 ;
        RECT 43.380 17.710 46.940 19.360 ;
        RECT 0.000 12.800 3.310 15.970 ;
        RECT 15.140 15.030 15.700 17.090 ;
        RECT 15.000 15.020 18.310 15.030 ;
        RECT 15.140 14.670 15.700 15.020 ;
        RECT 15.520 13.280 15.940 13.350 ;
        RECT 19.850 13.130 22.570 14.780 ;
        RECT 30.990 14.670 31.550 17.090 ;
        RECT 43.380 16.620 46.690 17.710 ;
        RECT 43.800 15.970 45.080 16.620 ;
        RECT 37.970 15.020 39.310 15.030 ;
        RECT 37.470 14.710 37.790 15.010 ;
        RECT 41.820 14.850 43.100 15.030 ;
        RECT 43.380 14.780 46.690 15.970 ;
        RECT 43.380 13.130 46.940 14.780 ;
        RECT 19.850 13.090 22.560 13.130 ;
        RECT 43.380 13.090 46.930 13.130 ;
        RECT 43.380 12.800 46.690 13.090 ;
        RECT 43.800 9.470 45.080 12.310 ;
        RECT 41.820 8.980 43.100 9.170 ;
        RECT 37.970 7.550 38.420 7.780 ;
        RECT 36.630 7.420 38.490 7.490 ;
        RECT 40.260 3.050 42.120 6.040 ;
        RECT 40.260 0.000 42.120 2.990 ;
      LAYER li1 ;
        RECT 0.820 21.590 1.370 22.020 ;
        RECT 45.320 21.590 45.870 22.020 ;
        RECT 0.820 19.860 1.370 20.290 ;
        RECT 45.320 19.860 45.870 20.290 ;
        RECT 0.400 19.060 0.600 19.410 ;
        RECT 1.880 19.160 2.410 19.330 ;
        RECT 44.280 19.160 44.810 19.330 ;
        RECT 0.390 19.030 0.600 19.060 ;
        RECT 46.090 19.060 46.290 19.410 ;
        RECT 46.090 19.030 46.300 19.060 ;
        RECT 0.390 18.450 0.610 19.030 ;
        RECT 0.390 18.440 0.600 18.450 ;
        RECT 0.770 18.270 0.960 18.280 ;
        RECT 0.760 17.980 0.960 18.270 ;
        RECT 0.700 17.650 0.970 17.980 ;
        RECT 1.160 17.170 1.330 18.780 ;
        RECT 7.310 18.770 7.500 19.000 ;
        RECT 1.150 16.980 1.330 17.170 ;
        RECT 1.990 17.080 2.160 18.770 ;
        RECT 2.580 18.580 2.910 18.750 ;
        RECT 3.930 18.580 4.280 18.750 ;
        RECT 7.590 18.720 8.470 18.890 ;
        RECT 7.780 18.330 7.970 18.440 ;
        RECT 7.670 18.210 7.970 18.330 ;
        RECT 8.300 18.330 8.470 18.720 ;
        RECT 7.670 18.160 7.890 18.210 ;
        RECT 8.300 18.160 8.690 18.330 ;
        RECT 20.150 18.230 20.380 18.920 ;
        RECT 44.520 18.230 44.750 18.920 ;
        RECT 2.580 17.790 2.910 17.960 ;
        RECT 3.930 17.790 4.280 17.960 ;
        RECT 39.750 17.940 40.070 17.980 ;
        RECT 39.750 17.750 40.080 17.940 ;
        RECT 39.750 17.720 40.070 17.750 ;
        RECT 6.380 17.370 6.700 17.410 ;
        RECT 7.630 17.370 8.710 17.540 ;
        RECT 9.040 17.370 10.120 17.540 ;
        RECT 6.370 17.180 6.700 17.370 ;
        RECT 2.580 17.000 2.910 17.170 ;
        RECT 3.930 17.000 4.270 17.170 ;
        RECT 6.380 17.150 6.700 17.180 ;
        RECT 44.530 17.080 44.700 18.230 ;
        RECT 45.360 17.170 45.530 18.780 ;
        RECT 46.080 18.450 46.300 19.030 ;
        RECT 46.090 18.440 46.300 18.450 ;
        RECT 45.730 18.270 45.920 18.280 ;
        RECT 45.730 17.980 45.930 18.270 ;
        RECT 45.720 17.650 46.010 17.980 ;
        RECT 7.310 16.780 7.500 17.010 ;
        RECT 45.360 16.980 45.540 17.170 ;
        RECT 7.610 16.580 7.690 16.750 ;
        RECT 8.170 16.430 8.380 16.860 ;
        RECT 8.190 16.410 8.360 16.430 ;
        RECT 6.370 15.680 6.690 15.720 ;
        RECT 7.320 15.710 7.510 15.940 ;
        RECT 7.640 15.840 7.690 16.010 ;
        RECT 7.780 15.890 7.970 16.120 ;
        RECT 8.780 16.010 8.950 16.580 ;
        RECT 13.060 16.430 13.250 16.750 ;
        RECT 33.440 16.430 33.630 16.750 ;
        RECT 13.060 16.340 13.340 16.430 ;
        RECT 9.700 16.200 13.340 16.340 ;
        RECT 33.350 16.340 33.630 16.430 ;
        RECT 44.360 16.540 44.690 16.710 ;
        RECT 44.800 16.630 45.130 16.800 ;
        RECT 33.350 16.200 36.990 16.340 ;
        RECT 44.360 16.260 44.720 16.540 ;
        RECT 9.700 16.160 13.250 16.200 ;
        RECT 8.060 15.980 8.110 15.990 ;
        RECT 8.690 15.980 8.770 15.990 ;
        RECT 8.060 15.940 8.770 15.980 ;
        RECT 8.060 15.900 8.790 15.940 ;
        RECT 8.020 15.780 8.860 15.900 ;
        RECT 13.060 15.740 13.250 16.160 ;
        RECT 33.440 16.160 36.990 16.200 ;
        RECT 33.440 15.740 33.630 16.160 ;
        RECT 42.290 16.010 42.610 16.050 ;
        RECT 42.290 15.820 42.620 16.010 ;
        RECT 42.290 15.790 42.610 15.820 ;
        RECT 42.690 15.800 42.890 16.130 ;
        RECT 43.280 15.940 43.480 16.130 ;
        RECT 44.010 16.090 44.720 16.260 ;
        RECT 43.950 15.970 44.270 16.010 ;
        RECT 1.150 15.420 1.330 15.610 ;
        RECT 0.700 14.610 0.970 14.940 ;
        RECT 0.760 14.320 0.960 14.610 ;
        RECT 0.770 14.310 0.960 14.320 ;
        RECT 0.390 14.140 0.600 14.150 ;
        RECT 0.390 13.560 0.610 14.140 ;
        RECT 1.160 13.810 1.330 15.420 ;
        RECT 1.990 13.820 2.160 15.510 ;
        RECT 2.580 15.420 2.910 15.590 ;
        RECT 3.930 15.420 4.270 15.590 ;
        RECT 6.360 15.490 6.690 15.680 ;
        RECT 6.370 15.460 6.690 15.490 ;
        RECT 42.970 15.610 43.160 15.620 ;
        RECT 43.170 15.610 43.520 15.940 ;
        RECT 43.950 15.780 44.280 15.970 ;
        RECT 43.950 15.750 44.270 15.780 ;
        RECT 7.630 15.050 8.710 15.220 ;
        RECT 9.030 15.050 10.270 15.220 ;
        RECT 39.750 15.180 40.070 15.220 ;
        RECT 34.470 15.120 34.700 15.160 ;
        RECT 39.750 14.990 40.080 15.180 ;
        RECT 42.060 15.100 42.230 15.430 ;
        RECT 42.240 15.360 42.560 15.400 ;
        RECT 42.240 15.170 42.570 15.360 ;
        RECT 42.240 15.140 42.560 15.170 ;
        RECT 42.690 15.140 42.890 15.470 ;
        RECT 42.970 15.280 43.520 15.610 ;
        RECT 39.750 14.960 40.070 14.990 ;
        RECT 43.170 14.950 43.520 15.280 ;
        RECT 2.580 14.630 2.910 14.800 ;
        RECT 3.930 14.630 4.280 14.800 ;
        RECT 9.360 14.730 9.530 14.790 ;
        RECT 44.010 14.770 44.710 15.650 ;
        RECT 45.360 15.420 45.540 15.610 ;
        RECT 7.770 14.430 7.960 14.540 ;
        RECT 9.340 14.520 9.550 14.730 ;
        RECT 9.360 14.450 9.530 14.520 ;
        RECT 7.670 14.310 7.960 14.430 ;
        RECT 8.230 14.420 8.690 14.430 ;
        RECT 7.670 14.260 7.880 14.310 ;
        RECT 8.230 14.270 8.700 14.420 ;
        RECT 43.350 14.380 43.540 14.610 ;
        RECT 44.530 14.350 44.700 14.770 ;
        RECT 8.230 14.260 8.690 14.270 ;
        RECT 2.580 13.840 2.910 14.010 ;
        RECT 3.930 13.840 4.280 14.010 ;
        RECT 7.340 13.920 7.530 14.030 ;
        RECT 8.230 13.920 8.420 14.260 ;
        RECT 7.340 13.800 8.420 13.920 ;
        RECT 7.460 13.740 8.420 13.800 ;
        RECT 20.150 13.570 20.380 14.260 ;
        RECT 42.060 13.840 42.230 14.170 ;
        RECT 42.240 14.100 42.560 14.130 ;
        RECT 42.240 13.910 42.570 14.100 ;
        RECT 42.240 13.870 42.560 13.910 ;
        RECT 42.690 13.800 42.890 14.130 ;
        RECT 43.170 13.990 43.520 14.320 ;
        RECT 44.000 14.260 44.700 14.350 ;
        RECT 44.000 14.170 44.750 14.260 ;
        RECT 42.970 13.660 43.520 13.990 ;
        RECT 42.970 13.650 43.160 13.660 ;
        RECT 0.390 13.530 0.600 13.560 ;
        RECT 0.400 13.180 0.600 13.530 ;
        RECT 42.290 13.450 42.610 13.480 ;
        RECT 1.880 13.260 2.410 13.430 ;
        RECT 42.290 13.260 42.620 13.450 ;
        RECT 42.290 13.220 42.610 13.260 ;
        RECT 42.690 13.140 42.890 13.470 ;
        RECT 43.170 13.330 43.520 13.660 ;
        RECT 44.000 13.750 44.320 13.790 ;
        RECT 44.000 13.560 44.330 13.750 ;
        RECT 44.520 13.570 44.750 14.170 ;
        RECT 45.360 13.810 45.530 15.420 ;
        RECT 45.720 14.610 46.010 14.940 ;
        RECT 45.730 14.320 45.930 14.610 ;
        RECT 45.730 14.310 45.920 14.320 ;
        RECT 46.090 14.140 46.300 14.150 ;
        RECT 46.080 13.560 46.300 14.140 ;
        RECT 44.000 13.530 44.320 13.560 ;
        RECT 46.090 13.530 46.300 13.560 ;
        RECT 43.280 13.140 43.480 13.330 ;
        RECT 44.280 13.260 44.810 13.430 ;
        RECT 46.090 13.180 46.290 13.530 ;
        RECT 42.290 13.010 42.610 13.050 ;
        RECT 42.290 12.820 42.620 13.010 ;
        RECT 42.290 12.790 42.610 12.820 ;
        RECT 42.690 12.800 42.890 13.130 ;
        RECT 43.280 12.940 43.480 13.130 ;
        RECT 43.990 13.030 44.310 13.070 ;
        RECT 42.970 12.610 43.160 12.620 ;
        RECT 43.170 12.610 43.520 12.940 ;
        RECT 43.990 12.840 44.320 13.030 ;
        RECT 43.990 12.810 44.310 12.840 ;
        RECT 42.060 12.100 42.230 12.430 ;
        RECT 42.240 12.360 42.560 12.400 ;
        RECT 42.240 12.170 42.570 12.360 ;
        RECT 42.240 12.140 42.560 12.170 ;
        RECT 42.690 12.140 42.890 12.470 ;
        RECT 42.970 12.280 43.520 12.610 ;
        RECT 43.170 12.020 43.520 12.280 ;
        RECT 43.170 11.950 43.540 12.020 ;
        RECT 43.350 11.790 43.540 11.950 ;
        RECT 44.000 11.890 44.700 12.070 ;
        RECT 42.060 10.840 42.230 11.170 ;
        RECT 42.240 11.100 42.560 11.130 ;
        RECT 42.240 10.910 42.570 11.100 ;
        RECT 42.240 10.870 42.560 10.910 ;
        RECT 42.690 10.800 42.890 11.130 ;
        RECT 43.170 10.990 43.520 11.320 ;
        RECT 42.970 10.660 43.520 10.990 ;
        RECT 44.010 10.820 44.710 11.470 ;
        RECT 42.970 10.650 43.160 10.660 ;
        RECT 37.720 10.550 38.040 10.590 ;
        RECT 37.710 10.360 38.040 10.550 ;
        RECT 37.720 10.350 38.040 10.360 ;
        RECT 37.710 10.330 38.040 10.350 ;
        RECT 42.290 10.450 42.610 10.480 ;
        RECT 37.710 10.020 37.880 10.330 ;
        RECT 42.290 10.260 42.620 10.450 ;
        RECT 42.290 10.220 42.610 10.260 ;
        RECT 42.690 10.140 42.890 10.470 ;
        RECT 43.170 10.330 43.520 10.660 ;
        RECT 43.910 10.590 44.710 10.820 ;
        RECT 43.910 10.560 44.230 10.590 ;
        RECT 43.280 10.140 43.480 10.330 ;
        RECT 44.010 9.980 44.720 10.150 ;
        RECT 37.870 9.720 38.190 9.760 ;
        RECT 37.860 9.530 38.190 9.720 ;
        RECT 44.360 9.700 44.720 9.980 ;
        RECT 44.360 9.530 44.690 9.700 ;
        RECT 37.870 9.500 38.190 9.530 ;
        RECT 44.800 9.440 45.130 9.610 ;
        RECT 37.060 8.900 37.380 8.930 ;
        RECT 37.060 8.710 37.390 8.900 ;
        RECT 37.060 8.670 37.380 8.710 ;
        RECT 37.040 6.950 37.220 8.010 ;
        RECT 37.790 7.620 38.110 7.650 ;
        RECT 37.790 7.550 38.120 7.620 ;
        RECT 37.650 7.430 38.120 7.550 ;
        RECT 37.650 7.420 38.110 7.430 ;
        RECT 37.770 7.390 38.110 7.420 ;
        RECT 37.770 7.320 37.820 7.390 ;
        RECT 37.690 6.990 37.860 7.320 ;
        RECT 38.090 6.790 38.170 6.870 ;
        RECT 38.230 6.790 38.420 6.910 ;
        RECT 38.090 6.700 38.420 6.790 ;
        RECT 38.230 6.680 38.420 6.700 ;
        RECT 40.670 3.520 40.850 5.570 ;
        RECT 41.400 5.310 41.730 5.480 ;
        RECT 41.480 3.530 41.650 5.310 ;
        RECT 40.670 0.470 40.850 2.520 ;
        RECT 41.400 2.260 41.730 2.430 ;
        RECT 41.480 0.480 41.650 2.260 ;
      LAYER mcon ;
        RECT 1.100 21.670 1.370 21.940 ;
        RECT 45.320 21.670 45.590 21.940 ;
        RECT 1.100 19.940 1.370 20.210 ;
        RECT 45.320 19.940 45.590 20.210 ;
        RECT 2.230 19.160 2.410 19.330 ;
        RECT 0.420 18.860 0.590 19.030 ;
        RECT 7.320 18.800 7.490 18.970 ;
        RECT 0.770 18.020 0.950 18.210 ;
        RECT 7.790 18.240 7.960 18.410 ;
        RECT 20.180 18.710 20.350 18.880 ;
        RECT 20.180 18.260 20.350 18.430 ;
        RECT 44.550 18.710 44.720 18.880 ;
        RECT 46.100 18.860 46.270 19.030 ;
        RECT 44.550 18.260 44.720 18.430 ;
        RECT 39.810 17.760 39.980 17.930 ;
        RECT 6.470 17.190 6.640 17.360 ;
        RECT 45.740 18.020 45.920 18.210 ;
        RECT 7.320 16.810 7.490 16.980 ;
        RECT 7.330 15.740 7.500 15.910 ;
        RECT 7.790 15.920 7.960 16.090 ;
        RECT 13.160 16.230 13.330 16.400 ;
        RECT 33.360 16.230 33.530 16.400 ;
        RECT 42.350 15.830 42.520 16.000 ;
        RECT 0.770 14.380 0.950 14.570 ;
        RECT 6.460 15.500 6.630 15.670 ;
        RECT 44.010 15.790 44.180 15.960 ;
        RECT 39.810 15.000 39.980 15.170 ;
        RECT 42.300 15.180 42.470 15.350 ;
        RECT 43.290 15.440 43.460 15.610 ;
        RECT 7.780 14.340 7.950 14.510 ;
        RECT 43.360 14.410 43.530 14.580 ;
        RECT 7.350 13.830 7.520 14.000 ;
        RECT 20.180 14.060 20.350 14.230 ;
        RECT 42.300 13.920 42.470 14.090 ;
        RECT 0.420 13.560 0.590 13.730 ;
        RECT 20.180 13.610 20.350 13.780 ;
        RECT 43.290 13.660 43.460 13.830 ;
        RECT 44.550 14.060 44.720 14.230 ;
        RECT 2.230 13.260 2.410 13.430 ;
        RECT 42.350 13.270 42.520 13.440 ;
        RECT 45.740 14.380 45.920 14.570 ;
        RECT 44.060 13.570 44.230 13.740 ;
        RECT 44.550 13.610 44.720 13.780 ;
        RECT 46.100 13.560 46.270 13.730 ;
        RECT 42.350 12.830 42.520 13.000 ;
        RECT 44.050 12.850 44.220 13.020 ;
        RECT 42.300 12.180 42.470 12.350 ;
        RECT 43.290 12.440 43.460 12.610 ;
        RECT 43.360 11.820 43.530 11.990 ;
        RECT 42.300 10.920 42.470 11.090 ;
        RECT 43.290 10.660 43.460 10.830 ;
        RECT 37.810 10.370 37.980 10.540 ;
        RECT 42.350 10.270 42.520 10.440 ;
        RECT 43.970 10.600 44.140 10.770 ;
        RECT 37.960 9.540 38.130 9.710 ;
        RECT 37.120 8.720 37.290 8.890 ;
        RECT 37.850 7.440 38.020 7.610 ;
        RECT 38.240 6.710 38.410 6.880 ;
      LAYER met1 ;
        RECT 0.360 19.090 0.520 19.730 ;
        RECT 0.360 18.540 0.630 19.090 ;
        RECT 0.350 18.490 0.630 18.540 ;
        RECT 0.350 18.400 0.520 18.490 ;
        RECT 0.360 16.710 0.520 18.400 ;
        RECT 0.770 18.280 0.960 19.730 ;
        RECT 1.040 19.400 1.430 22.990 ;
        RECT 45.260 19.400 45.650 22.990 ;
        RECT 2.170 18.920 2.480 19.360 ;
        RECT 5.120 19.270 5.280 19.320 ;
        RECT 5.530 19.260 5.720 19.320 ;
        RECT 7.400 19.030 7.610 19.320 ;
        RECT 7.290 18.740 7.610 19.030 ;
        RECT 0.740 18.250 0.960 18.280 ;
        RECT 0.730 17.980 0.980 18.250 ;
        RECT 0.730 17.970 0.970 17.980 ;
        RECT 0.740 17.730 0.970 17.970 ;
        RECT 0.770 16.710 0.930 17.730 ;
        RECT 1.120 16.920 1.360 17.300 ;
        RECT 6.390 17.120 6.710 17.440 ;
        RECT 7.400 17.040 7.610 18.740 ;
        RECT 7.870 18.470 8.060 19.320 ;
        RECT 7.760 18.180 8.060 18.470 ;
        RECT 7.290 16.750 7.610 17.040 ;
        RECT 5.760 16.500 6.020 16.560 ;
        RECT 7.400 16.530 7.610 16.750 ;
        RECT 5.760 16.240 6.120 16.500 ;
        RECT 5.880 16.080 6.120 16.240 ;
        RECT 7.870 16.150 8.060 18.180 ;
        RECT 8.280 16.860 8.490 19.320 ;
        RECT 8.160 16.350 8.490 16.860 ;
        RECT 7.420 15.970 7.610 16.020 ;
        RECT 0.360 14.190 0.520 15.880 ;
        RECT 0.770 14.860 0.930 15.880 ;
        RECT 1.120 15.290 1.360 15.670 ;
        RECT 6.380 15.430 6.700 15.750 ;
        RECT 7.300 15.680 7.610 15.970 ;
        RECT 7.760 15.860 8.060 16.150 ;
        RECT 0.740 14.620 0.970 14.860 ;
        RECT 0.730 14.610 0.970 14.620 ;
        RECT 0.730 14.340 0.980 14.610 ;
        RECT 0.740 14.310 0.960 14.340 ;
        RECT 0.350 14.100 0.520 14.190 ;
        RECT 0.350 14.050 0.630 14.100 ;
        RECT 0.360 13.500 0.630 14.050 ;
        RECT 0.360 12.860 0.520 13.500 ;
        RECT 0.770 12.860 0.960 14.310 ;
        RECT 7.420 14.060 7.610 15.680 ;
        RECT 7.870 14.570 8.060 15.860 ;
        RECT 7.750 14.280 8.060 14.570 ;
        RECT 7.100 13.770 7.110 13.780 ;
        RECT 7.320 13.770 7.610 14.060 ;
        RECT 2.170 13.230 2.480 13.670 ;
        RECT 5.120 13.270 5.280 13.320 ;
        RECT 5.530 13.270 5.720 13.320 ;
        RECT 7.410 13.270 7.640 13.770 ;
        RECT 7.870 13.270 8.060 14.280 ;
        RECT 8.280 13.270 8.490 16.350 ;
        RECT 9.360 14.790 9.540 19.320 ;
        RECT 13.230 16.460 13.460 19.320 ;
        RECT 20.130 18.180 20.390 18.970 ;
        RECT 13.130 16.170 13.460 16.460 ;
        RECT 9.300 14.450 9.590 14.790 ;
        RECT 9.360 13.270 9.540 14.450 ;
        RECT 13.230 13.270 13.460 16.170 ;
        RECT 20.130 13.520 20.390 14.310 ;
        RECT 30.750 13.270 31.170 19.320 ;
        RECT 33.230 16.460 33.460 19.320 ;
        RECT 33.230 16.170 33.560 16.460 ;
        RECT 33.230 13.270 33.460 16.170 ;
        RECT 34.450 13.270 34.680 19.320 ;
        RECT 40.970 19.280 41.160 19.320 ;
        RECT 39.740 17.690 40.060 18.010 ;
        RECT 40.660 16.530 40.920 16.850 ;
        RECT 41.410 16.570 41.690 19.320 ;
        RECT 44.210 18.970 44.520 19.360 ;
        RECT 44.210 18.920 44.760 18.970 ;
        RECT 44.500 18.180 44.760 18.920 ;
        RECT 45.730 18.280 45.920 19.730 ;
        RECT 46.170 19.090 46.330 19.730 ;
        RECT 46.060 18.540 46.330 19.090 ;
        RECT 46.060 18.490 46.340 18.540 ;
        RECT 46.170 18.400 46.340 18.490 ;
        RECT 45.730 18.250 45.950 18.280 ;
        RECT 45.710 17.980 45.960 18.250 ;
        RECT 45.720 17.970 45.960 17.980 ;
        RECT 45.720 17.730 45.950 17.970 ;
        RECT 45.330 16.920 45.570 17.300 ;
        RECT 45.760 16.710 45.920 17.730 ;
        RECT 46.170 16.710 46.330 18.400 ;
        RECT 41.410 16.250 41.860 16.570 ;
        RECT 40.660 15.930 40.920 16.250 ;
        RECT 39.740 14.930 40.060 15.250 ;
        RECT 41.410 15.030 41.690 16.250 ;
        RECT 42.280 16.000 42.600 16.080 ;
        RECT 42.280 15.760 42.850 16.000 ;
        RECT 42.510 15.430 42.850 15.760 ;
        RECT 42.230 15.110 42.850 15.430 ;
        RECT 41.140 14.890 41.690 15.030 ;
        RECT 40.970 13.270 41.160 13.320 ;
        RECT 41.410 13.270 41.690 14.890 ;
        RECT 42.510 14.160 42.850 15.110 ;
        RECT 42.230 13.840 42.850 14.160 ;
        RECT 42.510 13.510 42.850 13.840 ;
        RECT 42.280 13.190 42.850 13.510 ;
        RECT 42.510 13.080 42.850 13.190 ;
        RECT 42.280 12.760 42.850 13.080 ;
        RECT 42.510 12.430 42.850 12.760 ;
        RECT 42.230 12.110 42.850 12.430 ;
        RECT 42.510 11.160 42.850 12.110 ;
        RECT 42.230 10.840 42.850 11.160 ;
        RECT 37.730 10.300 38.050 10.620 ;
        RECT 42.510 10.510 42.850 10.840 ;
        RECT 42.280 10.280 42.850 10.510 ;
        RECT 43.180 15.670 43.450 15.990 ;
        RECT 43.940 15.720 44.260 16.040 ;
        RECT 43.180 15.380 43.490 15.670 ;
        RECT 43.180 14.640 43.450 15.380 ;
        RECT 45.330 15.290 45.570 15.670 ;
        RECT 45.760 14.860 45.920 15.880 ;
        RECT 43.180 14.350 43.560 14.640 ;
        RECT 45.720 14.620 45.950 14.860 ;
        RECT 45.720 14.610 45.960 14.620 ;
        RECT 43.180 13.890 43.450 14.350 ;
        RECT 45.710 14.340 45.960 14.610 ;
        RECT 45.730 14.310 45.950 14.340 ;
        RECT 43.180 13.600 43.490 13.890 ;
        RECT 43.990 13.670 44.310 13.820 ;
        RECT 44.500 13.670 44.760 14.310 ;
        RECT 43.180 12.670 43.450 13.600 ;
        RECT 43.990 13.520 44.760 13.670 ;
        RECT 43.990 13.500 44.520 13.520 ;
        RECT 44.210 13.230 44.520 13.500 ;
        RECT 43.980 12.780 44.300 13.100 ;
        RECT 45.730 12.860 45.920 14.310 ;
        RECT 46.170 14.190 46.330 15.880 ;
        RECT 46.170 14.100 46.340 14.190 ;
        RECT 46.060 14.050 46.340 14.100 ;
        RECT 46.060 13.500 46.330 14.050 ;
        RECT 46.170 12.860 46.330 13.500 ;
        RECT 43.180 12.380 43.490 12.670 ;
        RECT 43.180 12.050 43.450 12.380 ;
        RECT 43.180 11.760 43.560 12.050 ;
        RECT 43.180 10.890 43.450 11.760 ;
        RECT 43.180 10.600 43.490 10.890 ;
        RECT 43.180 10.290 43.450 10.600 ;
        RECT 43.900 10.530 44.220 10.850 ;
        RECT 42.280 10.190 42.600 10.280 ;
        RECT 37.880 9.470 38.200 9.790 ;
        RECT 23.420 9.030 23.740 9.330 ;
        RECT 29.220 9.030 29.540 9.330 ;
        RECT 39.610 9.180 39.930 9.480 ;
        RECT 39.610 9.150 40.040 9.180 ;
        RECT 40.640 9.170 41.150 9.180 ;
        RECT 40.640 9.150 41.480 9.170 ;
        RECT 39.610 9.120 41.480 9.150 ;
        RECT 39.760 9.070 41.480 9.120 ;
        RECT 39.790 9.040 41.480 9.070 ;
        RECT 39.820 9.020 41.480 9.040 ;
        RECT 39.890 9.010 40.850 9.020 ;
        RECT 41.140 8.980 41.480 9.020 ;
        RECT 37.050 8.640 37.370 8.960 ;
        RECT 38.130 8.530 38.340 8.740 ;
        RECT 38.130 8.210 38.460 8.530 ;
        RECT 37.780 7.360 38.100 7.680 ;
        RECT 38.130 6.970 38.340 8.210 ;
        RECT 38.210 6.650 38.440 6.940 ;
      LAYER via ;
        RECT 2.190 18.950 2.450 19.210 ;
        RECT 6.420 17.150 6.680 17.410 ;
        RECT 5.760 16.270 6.020 16.530 ;
        RECT 6.410 15.460 6.670 15.720 ;
        RECT 2.190 13.380 2.450 13.640 ;
        RECT 39.770 17.720 40.030 17.980 ;
        RECT 40.660 16.560 40.920 16.820 ;
        RECT 44.240 18.950 44.500 19.210 ;
        RECT 41.600 16.280 41.860 16.540 ;
        RECT 40.660 15.960 40.920 16.220 ;
        RECT 39.770 14.960 40.030 15.220 ;
        RECT 42.310 15.790 42.570 16.050 ;
        RECT 42.260 15.140 42.520 15.400 ;
        RECT 42.260 13.870 42.520 14.130 ;
        RECT 42.310 13.220 42.570 13.480 ;
        RECT 42.310 12.790 42.570 13.050 ;
        RECT 42.260 12.140 42.520 12.400 ;
        RECT 42.260 10.870 42.520 11.130 ;
        RECT 37.760 10.330 38.020 10.590 ;
        RECT 42.310 10.220 42.570 10.480 ;
        RECT 43.970 15.750 44.230 16.010 ;
        RECT 44.020 13.640 44.280 13.790 ;
        RECT 44.020 13.530 44.500 13.640 ;
        RECT 44.240 13.380 44.500 13.530 ;
        RECT 44.010 12.810 44.270 13.070 ;
        RECT 43.930 10.560 44.190 10.820 ;
        RECT 37.910 9.500 38.170 9.760 ;
        RECT 23.450 9.050 23.710 9.310 ;
        RECT 29.250 9.050 29.510 9.310 ;
        RECT 39.640 9.200 39.900 9.460 ;
        RECT 37.080 8.670 37.340 8.930 ;
        RECT 38.200 8.240 38.460 8.500 ;
        RECT 37.810 7.390 38.070 7.650 ;
      LAYER met2 ;
        RECT 2.170 19.240 2.480 19.250 ;
        RECT 0.000 19.060 2.480 19.240 ;
        RECT 2.170 18.920 2.480 19.060 ;
        RECT 44.210 19.240 44.520 19.250 ;
        RECT 44.210 19.060 46.690 19.240 ;
        RECT 44.210 18.920 44.520 19.060 ;
        RECT 7.170 18.820 7.490 18.840 ;
        RECT 4.760 18.640 4.840 18.820 ;
        RECT 7.170 18.640 16.280 18.820 ;
        RECT 30.400 18.640 39.520 18.820 ;
        RECT 39.740 17.800 40.050 18.020 ;
        RECT 39.740 17.690 41.930 17.800 ;
        RECT 39.900 17.580 41.930 17.690 ;
        RECT 6.400 17.280 6.710 17.450 ;
        RECT 6.400 17.120 16.280 17.280 ;
        RECT 6.570 17.090 16.280 17.120 ;
        RECT 40.630 16.560 40.950 16.820 ;
        RECT 5.730 16.270 6.050 16.530 ;
        RECT 6.120 16.360 16.280 16.400 ;
        RECT 6.110 16.170 16.280 16.360 ;
        RECT 42.280 15.800 42.590 16.090 ;
        RECT 43.940 15.800 44.250 16.050 ;
        RECT 6.390 15.430 6.700 15.760 ;
        RECT 41.560 15.720 44.250 15.800 ;
        RECT 41.560 15.570 44.100 15.720 ;
        RECT 6.560 15.230 16.280 15.420 ;
        RECT 39.740 15.040 40.050 15.260 ;
        RECT 41.790 15.040 42.120 15.210 ;
        RECT 42.230 15.110 42.540 15.440 ;
        RECT 39.740 15.000 42.120 15.040 ;
        RECT 39.740 14.930 41.930 15.000 ;
        RECT 39.890 14.830 41.930 14.930 ;
        RECT 39.680 14.130 39.900 14.150 ;
        RECT 4.760 13.770 4.840 13.950 ;
        RECT 7.070 13.940 7.230 13.960 ;
        RECT 39.460 13.940 39.620 13.960 ;
        RECT 7.070 13.890 16.280 13.940 ;
        RECT 7.190 13.790 16.280 13.890 ;
        RECT 30.400 13.890 39.620 13.940 ;
        RECT 30.400 13.790 39.500 13.890 ;
        RECT 39.630 13.790 39.900 14.130 ;
        RECT 41.790 14.060 42.120 14.270 ;
        RECT 42.230 13.830 42.540 14.160 ;
        RECT 43.990 13.670 44.300 13.830 ;
        RECT 2.170 13.530 2.480 13.670 ;
        RECT 43.990 13.660 44.520 13.670 ;
        RECT 0.000 13.350 2.480 13.530 ;
        RECT 41.820 13.530 44.520 13.660 ;
        RECT 2.170 13.340 2.480 13.350 ;
        RECT 37.890 13.290 38.240 13.510 ;
        RECT 41.820 13.430 46.690 13.530 ;
        RECT 39.700 13.220 39.900 13.230 ;
        RECT 26.510 12.800 34.500 13.000 ;
        RECT 39.700 12.890 39.920 13.220 ;
        RECT 42.280 13.180 42.590 13.430 ;
        RECT 44.210 13.350 46.690 13.430 ;
        RECT 44.210 13.340 44.520 13.350 ;
        RECT 39.720 12.880 39.920 12.890 ;
        RECT 42.280 12.830 42.590 13.090 ;
        RECT 43.980 12.830 44.290 13.110 ;
        RECT 33.100 12.120 33.320 12.130 ;
        RECT 26.520 11.870 33.350 12.120 ;
        RECT 34.280 12.080 34.500 12.800 ;
        RECT 41.560 12.610 44.470 12.830 ;
        RECT 26.520 10.950 30.030 11.140 ;
        RECT 29.800 10.350 30.030 10.950 ;
        RECT 33.060 10.700 33.350 11.870 ;
        RECT 34.250 12.040 34.500 12.080 ;
        RECT 34.250 11.400 34.510 12.040 ;
        RECT 41.790 12.000 42.120 12.210 ;
        RECT 42.230 12.110 42.540 12.440 ;
        RECT 34.250 11.190 38.380 11.400 ;
        RECT 38.170 11.050 38.380 11.190 ;
        RECT 41.790 11.060 42.120 11.270 ;
        RECT 38.170 10.840 40.180 11.050 ;
        RECT 42.230 10.830 42.540 11.160 ;
        RECT 33.060 10.480 35.950 10.700 ;
        RECT 43.900 10.670 44.210 10.860 ;
        RECT 33.060 10.470 33.350 10.480 ;
        RECT 37.740 10.470 38.050 10.630 ;
        RECT 29.800 10.200 30.020 10.350 ;
        RECT 37.310 10.250 38.190 10.470 ;
        RECT 41.550 10.440 44.260 10.670 ;
        RECT 34.170 10.200 40.170 10.250 ;
        RECT 29.800 10.050 40.170 10.200 ;
        RECT 42.280 10.180 42.590 10.440 ;
        RECT 29.800 10.040 40.040 10.050 ;
        RECT 29.800 9.980 34.560 10.040 ;
        RECT 37.890 9.610 38.200 9.800 ;
        RECT 37.850 9.360 38.400 9.610 ;
        RECT 37.050 8.630 37.360 8.960 ;
        RECT 38.030 8.330 38.500 8.580 ;
        RECT 38.170 8.240 38.490 8.330 ;
        RECT 37.550 7.780 37.980 7.790 ;
        RECT 37.550 7.550 38.420 7.780 ;
        RECT 37.780 7.350 38.090 7.550 ;
  END
END sky130_hilas_TA2Cell_1FG_Strong

MACRO sky130_hilas_TA2Cell_NoFG
  CLASS CORE ;
  FOREIGN sky130_hilas_TA2Cell_NoFG ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.500 BY 24.010 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN COLSEL1
    PORT
      LAYER met1 ;
        RECT 10.570 14.950 10.760 15.030 ;
    END
  END COLSEL1
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 11.870 9.000 12.130 9.250 ;
    END
  END VIN12
  PIN VIN21
    PORT
      LAYER met2 ;
        RECT 13.470 12.090 13.720 12.320 ;
    END
  END VIN21
  PIN VIN22
    PORT
      LAYER met2 ;
        RECT 13.300 15.040 13.610 15.260 ;
        RECT 13.300 14.930 15.490 15.040 ;
        RECT 13.430 14.830 15.490 14.930 ;
        RECT 13.430 14.760 13.680 14.830 ;
    END
  END VIN22
  PIN OUTPUT1
    PORT
      LAYER met2 ;
        RECT 17.770 11.500 17.920 11.720 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    PORT
      LAYER met2 ;
        RECT 17.770 12.320 17.920 12.540 ;
    END
  END OUTPUT2
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 15.960 8.980 16.300 9.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.960 14.890 16.300 15.030 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 16.630 8.980 16.900 9.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 16.630 14.880 16.900 15.030 ;
    END
  END VPWR
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 0.000 14.350 0.070 14.530 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 0.000 9.500 0.080 9.650 ;
    END
  END DRAIN2
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 0.350 14.960 0.770 15.030 ;
    END
  END VTUN
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT 4.050 14.950 4.280 15.030 ;
    END
  END GATE1
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 11.010 14.950 11.290 15.030 ;
    END
  END VINJ
  PIN VIN11
    PORT
      LAYER met2 ;
        RECT 11.910 11.680 12.190 11.920 ;
    END
  END VIN11
  OBS
      LAYER nwell ;
        RECT 13.520 21.020 15.380 24.010 ;
        RECT 18.480 22.980 20.210 23.320 ;
        RECT 18.460 21.420 20.210 22.980 ;
        RECT 13.520 19.320 15.380 20.960 ;
        RECT 18.460 19.790 20.190 21.420 ;
        RECT 16.940 19.400 20.250 19.790 ;
        RECT 16.940 19.360 20.490 19.400 ;
        RECT 12.180 19.310 15.490 19.320 ;
        RECT 13.520 17.970 15.380 19.310 ;
        RECT 16.940 17.710 20.500 19.360 ;
        RECT 4.550 14.670 5.110 17.090 ;
        RECT 16.940 16.620 20.250 17.710 ;
        RECT 9.890 16.520 11.750 16.590 ;
        RECT 11.230 16.230 11.680 16.460 ;
        RECT 18.620 15.970 19.900 16.620 ;
        RECT 16.940 15.030 20.250 15.970 ;
        RECT 16.650 14.850 20.250 15.030 ;
        RECT 16.940 14.780 20.250 14.850 ;
        RECT 11.450 13.290 13.110 13.510 ;
        RECT 16.940 13.130 20.500 14.780 ;
        RECT 16.940 13.090 20.490 13.130 ;
        RECT 16.940 12.800 20.250 13.090 ;
        RECT 11.910 11.680 12.190 11.920 ;
        RECT 18.620 9.470 19.900 12.310 ;
        RECT 16.640 8.980 17.920 9.170 ;
        RECT 12.790 7.550 13.240 7.780 ;
        RECT 11.450 7.420 13.310 7.490 ;
        RECT 15.080 3.050 16.940 6.040 ;
        RECT 15.080 0.000 16.940 2.990 ;
      LAYER li1 ;
        RECT 13.930 21.490 14.110 23.540 ;
        RECT 14.740 21.750 14.910 23.530 ;
        RECT 14.660 21.580 14.990 21.750 ;
        RECT 18.880 21.590 19.430 22.020 ;
        RECT 13.930 18.440 14.110 20.490 ;
        RECT 14.740 18.700 14.910 20.480 ;
        RECT 18.880 19.860 19.430 20.290 ;
        RECT 17.840 19.160 18.370 19.330 ;
        RECT 19.650 19.060 19.850 19.410 ;
        RECT 19.650 19.030 19.860 19.060 ;
        RECT 14.660 18.530 14.990 18.700 ;
        RECT 18.080 18.230 18.310 18.920 ;
        RECT 13.310 17.940 13.630 17.980 ;
        RECT 13.310 17.750 13.640 17.940 ;
        RECT 13.310 17.720 13.630 17.750 ;
        RECT 11.490 17.310 11.680 17.330 ;
        RECT 11.350 17.220 11.680 17.310 ;
        RECT 11.350 17.140 11.430 17.220 ;
        RECT 11.490 17.100 11.680 17.220 ;
        RECT 18.090 17.080 18.260 18.230 ;
        RECT 18.920 17.170 19.090 18.780 ;
        RECT 19.640 18.450 19.860 19.030 ;
        RECT 19.650 18.440 19.860 18.450 ;
        RECT 19.290 18.270 19.480 18.280 ;
        RECT 19.290 17.980 19.490 18.270 ;
        RECT 19.280 17.650 19.570 17.980 ;
        RECT 7.000 16.430 7.190 16.750 ;
        RECT 6.910 16.340 7.190 16.430 ;
        RECT 10.300 16.340 10.480 17.060 ;
        RECT 10.950 16.690 11.120 17.020 ;
        RECT 18.920 16.980 19.100 17.170 ;
        RECT 11.030 16.620 11.080 16.690 ;
        RECT 11.030 16.590 11.370 16.620 ;
        RECT 10.910 16.580 11.370 16.590 ;
        RECT 10.910 16.460 11.380 16.580 ;
        RECT 11.050 16.390 11.380 16.460 ;
        RECT 19.180 16.540 19.510 16.710 ;
        RECT 19.620 16.630 19.950 16.800 ;
        RECT 11.050 16.360 11.370 16.390 ;
        RECT 6.910 16.200 10.550 16.340 ;
        RECT 19.180 16.260 19.540 16.540 ;
        RECT 7.000 16.160 10.550 16.200 ;
        RECT 7.000 15.740 7.190 16.160 ;
        RECT 10.300 16.000 10.480 16.160 ;
        RECT 17.110 16.010 17.430 16.050 ;
        RECT 17.110 15.820 17.440 16.010 ;
        RECT 17.110 15.790 17.430 15.820 ;
        RECT 17.510 15.800 17.710 16.130 ;
        RECT 18.100 15.940 18.300 16.130 ;
        RECT 18.830 16.090 19.540 16.260 ;
        RECT 18.770 15.970 19.090 16.010 ;
        RECT 17.790 15.610 17.980 15.620 ;
        RECT 17.990 15.610 18.340 15.940 ;
        RECT 18.770 15.780 19.100 15.970 ;
        RECT 18.770 15.750 19.090 15.780 ;
        RECT 10.320 15.300 10.640 15.340 ;
        RECT 8.030 15.120 8.260 15.160 ;
        RECT 10.320 15.110 10.650 15.300 ;
        RECT 13.310 15.180 13.630 15.220 ;
        RECT 10.320 15.080 10.640 15.110 ;
        RECT 13.310 14.990 13.640 15.180 ;
        RECT 16.880 15.100 17.050 15.430 ;
        RECT 17.060 15.360 17.380 15.400 ;
        RECT 17.060 15.170 17.390 15.360 ;
        RECT 17.060 15.140 17.380 15.170 ;
        RECT 17.510 15.140 17.710 15.470 ;
        RECT 17.790 15.280 18.340 15.610 ;
        RECT 13.310 14.960 13.630 14.990 ;
        RECT 17.990 14.950 18.340 15.280 ;
        RECT 18.090 14.610 18.260 14.950 ;
        RECT 18.830 14.940 19.530 15.650 ;
        RECT 18.830 14.770 19.570 14.940 ;
        RECT 11.130 14.480 11.450 14.510 ;
        RECT 11.120 14.290 11.450 14.480 ;
        RECT 18.090 14.380 18.360 14.610 ;
        RECT 18.090 14.320 18.260 14.380 ;
        RECT 18.920 14.350 19.090 14.770 ;
        RECT 19.280 14.610 19.570 14.770 ;
        RECT 19.290 14.350 19.490 14.610 ;
        RECT 11.130 14.250 11.450 14.290 ;
        RECT 10.970 13.680 11.140 13.990 ;
        RECT 16.880 13.840 17.050 14.170 ;
        RECT 17.060 14.100 17.380 14.130 ;
        RECT 17.060 13.910 17.390 14.100 ;
        RECT 17.060 13.870 17.380 13.910 ;
        RECT 17.510 13.800 17.710 14.130 ;
        RECT 17.990 13.990 18.340 14.320 ;
        RECT 18.820 14.170 19.520 14.350 ;
        RECT 10.970 13.660 11.300 13.680 ;
        RECT 10.980 13.650 11.300 13.660 ;
        RECT 17.790 13.660 18.340 13.990 ;
        RECT 18.920 13.810 19.090 14.170 ;
        RECT 19.650 14.140 19.860 14.150 ;
        RECT 17.790 13.650 17.980 13.660 ;
        RECT 10.970 13.460 11.300 13.650 ;
        RECT 10.980 13.420 11.300 13.460 ;
        RECT 17.110 13.450 17.430 13.480 ;
        RECT 17.110 13.260 17.440 13.450 ;
        RECT 17.110 13.220 17.430 13.260 ;
        RECT 17.510 13.140 17.710 13.470 ;
        RECT 17.990 13.430 18.340 13.660 ;
        RECT 18.820 13.750 19.140 13.790 ;
        RECT 18.820 13.560 19.150 13.750 ;
        RECT 19.640 13.560 19.860 14.140 ;
        RECT 18.820 13.530 19.140 13.560 ;
        RECT 19.650 13.530 19.860 13.560 ;
        RECT 17.840 13.260 18.370 13.430 ;
        RECT 18.100 13.140 18.300 13.260 ;
        RECT 19.650 13.180 19.850 13.530 ;
        RECT 17.110 13.010 17.430 13.050 ;
        RECT 17.110 12.820 17.440 13.010 ;
        RECT 17.110 12.790 17.430 12.820 ;
        RECT 17.510 12.800 17.710 13.130 ;
        RECT 18.100 12.940 18.300 13.130 ;
        RECT 18.810 13.030 19.130 13.070 ;
        RECT 17.790 12.610 17.980 12.620 ;
        RECT 17.990 12.610 18.340 12.940 ;
        RECT 18.810 12.840 19.140 13.030 ;
        RECT 18.810 12.810 19.130 12.840 ;
        RECT 2.830 11.450 3.290 12.460 ;
        RECT 16.880 12.100 17.050 12.430 ;
        RECT 17.060 12.360 17.380 12.400 ;
        RECT 17.060 12.170 17.390 12.360 ;
        RECT 17.060 12.140 17.380 12.170 ;
        RECT 17.510 12.140 17.710 12.470 ;
        RECT 17.790 12.280 18.340 12.610 ;
        RECT 17.990 12.020 18.340 12.280 ;
        RECT 17.990 11.950 18.360 12.020 ;
        RECT 18.170 11.790 18.360 11.950 ;
        RECT 18.820 11.890 19.520 12.070 ;
        RECT 16.880 10.840 17.050 11.170 ;
        RECT 17.060 11.100 17.380 11.130 ;
        RECT 17.060 10.910 17.390 11.100 ;
        RECT 17.060 10.870 17.380 10.910 ;
        RECT 17.510 10.800 17.710 11.130 ;
        RECT 17.990 10.990 18.340 11.320 ;
        RECT 17.790 10.660 18.340 10.990 ;
        RECT 18.830 10.820 19.530 11.470 ;
        RECT 17.790 10.650 17.980 10.660 ;
        RECT 12.540 10.550 12.860 10.590 ;
        RECT 12.530 10.360 12.860 10.550 ;
        RECT 12.540 10.350 12.860 10.360 ;
        RECT 12.530 10.330 12.860 10.350 ;
        RECT 17.110 10.450 17.430 10.480 ;
        RECT 12.530 10.020 12.700 10.330 ;
        RECT 17.110 10.260 17.440 10.450 ;
        RECT 17.110 10.220 17.430 10.260 ;
        RECT 17.510 10.140 17.710 10.470 ;
        RECT 17.990 10.330 18.340 10.660 ;
        RECT 18.730 10.590 19.530 10.820 ;
        RECT 18.730 10.560 19.050 10.590 ;
        RECT 18.100 10.140 18.300 10.330 ;
        RECT 18.830 9.980 19.540 10.150 ;
        RECT 12.690 9.720 13.010 9.760 ;
        RECT 12.680 9.530 13.010 9.720 ;
        RECT 19.180 9.700 19.540 9.980 ;
        RECT 19.180 9.530 19.510 9.700 ;
        RECT 12.690 9.500 13.010 9.530 ;
        RECT 19.620 9.440 19.950 9.610 ;
        RECT 11.880 8.900 12.200 8.930 ;
        RECT 11.880 8.710 12.210 8.900 ;
        RECT 11.880 8.670 12.200 8.710 ;
        RECT 11.860 6.950 12.040 8.010 ;
        RECT 12.610 7.620 12.930 7.650 ;
        RECT 12.610 7.550 12.940 7.620 ;
        RECT 12.470 7.430 12.940 7.550 ;
        RECT 12.470 7.420 12.930 7.430 ;
        RECT 12.590 7.390 12.930 7.420 ;
        RECT 12.590 7.320 12.640 7.390 ;
        RECT 12.510 6.990 12.680 7.320 ;
        RECT 12.910 6.790 12.990 6.870 ;
        RECT 13.050 6.790 13.240 6.910 ;
        RECT 12.910 6.700 13.240 6.790 ;
        RECT 13.050 6.680 13.240 6.700 ;
        RECT 15.490 3.520 15.670 5.570 ;
        RECT 16.220 5.310 16.550 5.480 ;
        RECT 16.300 3.530 16.470 5.310 ;
        RECT 15.490 0.470 15.670 2.520 ;
        RECT 16.220 2.260 16.550 2.430 ;
        RECT 16.300 0.480 16.470 2.260 ;
      LAYER mcon ;
        RECT 18.880 21.670 19.150 21.940 ;
        RECT 18.880 19.940 19.150 20.210 ;
        RECT 18.110 18.710 18.280 18.880 ;
        RECT 19.660 18.860 19.830 19.030 ;
        RECT 18.110 18.260 18.280 18.430 ;
        RECT 13.370 17.760 13.540 17.930 ;
        RECT 11.500 17.130 11.670 17.300 ;
        RECT 19.300 18.020 19.480 18.210 ;
        RECT 6.920 16.230 7.090 16.400 ;
        RECT 11.110 16.400 11.280 16.570 ;
        RECT 17.170 15.830 17.340 16.000 ;
        RECT 18.830 15.790 19.000 15.960 ;
        RECT 10.380 15.120 10.550 15.290 ;
        RECT 13.370 15.000 13.540 15.170 ;
        RECT 17.120 15.180 17.290 15.350 ;
        RECT 18.110 15.440 18.280 15.610 ;
        RECT 18.920 15.420 19.100 15.610 ;
        RECT 11.220 14.300 11.390 14.470 ;
        RECT 18.180 14.410 18.350 14.580 ;
        RECT 19.300 14.380 19.480 14.570 ;
        RECT 17.120 13.920 17.290 14.090 ;
        RECT 18.110 14.060 18.280 14.230 ;
        RECT 11.070 13.470 11.240 13.640 ;
        RECT 18.110 13.610 18.280 13.830 ;
        RECT 17.170 13.270 17.340 13.440 ;
        RECT 18.880 13.570 19.050 13.740 ;
        RECT 19.660 13.560 19.830 13.730 ;
        RECT 17.170 12.830 17.340 13.000 ;
        RECT 18.870 12.850 19.040 13.020 ;
        RECT 2.860 12.200 3.030 12.370 ;
        RECT 17.120 12.180 17.290 12.350 ;
        RECT 18.110 12.440 18.280 12.610 ;
        RECT 18.180 11.820 18.350 11.990 ;
        RECT 2.860 11.510 3.030 11.680 ;
        RECT 17.120 10.920 17.290 11.090 ;
        RECT 18.110 10.660 18.280 10.830 ;
        RECT 12.630 10.370 12.800 10.540 ;
        RECT 17.170 10.270 17.340 10.440 ;
        RECT 18.790 10.600 18.960 10.770 ;
        RECT 12.780 9.540 12.950 9.710 ;
        RECT 11.940 8.720 12.110 8.890 ;
        RECT 12.670 7.440 12.840 7.610 ;
        RECT 13.060 6.710 13.230 6.880 ;
      LAYER met1 ;
        RECT 18.820 19.400 19.210 22.990 ;
        RECT 4.310 13.270 4.730 19.320 ;
        RECT 6.790 16.460 7.020 19.320 ;
        RECT 6.790 16.170 7.120 16.460 ;
        RECT 6.790 13.270 7.020 16.170 ;
        RECT 8.010 13.270 8.240 19.320 ;
        RECT 14.530 19.280 14.720 19.320 ;
        RECT 13.300 17.690 13.620 18.010 ;
        RECT 11.470 17.070 11.700 17.360 ;
        RECT 11.040 16.330 11.360 16.650 ;
        RECT 11.390 15.800 11.600 17.040 ;
        RECT 14.220 16.530 14.480 16.850 ;
        RECT 14.970 16.570 15.250 19.320 ;
        RECT 17.770 18.970 18.080 19.360 ;
        RECT 17.770 18.920 18.320 18.970 ;
        RECT 18.060 18.180 18.320 18.920 ;
        RECT 19.290 18.280 19.480 19.730 ;
        RECT 19.730 19.090 19.890 19.730 ;
        RECT 19.620 18.540 19.890 19.090 ;
        RECT 19.620 18.490 19.900 18.540 ;
        RECT 19.730 18.400 19.900 18.490 ;
        RECT 19.290 18.250 19.510 18.280 ;
        RECT 19.270 17.980 19.520 18.250 ;
        RECT 19.280 17.970 19.520 17.980 ;
        RECT 19.280 17.730 19.510 17.970 ;
        RECT 18.890 16.920 19.130 17.300 ;
        RECT 19.320 16.710 19.480 17.730 ;
        RECT 19.730 16.710 19.890 18.400 ;
        RECT 14.970 16.250 15.420 16.570 ;
        RECT 14.220 15.930 14.480 16.250 ;
        RECT 11.390 15.480 11.720 15.800 ;
        RECT 10.310 15.050 10.630 15.370 ;
        RECT 11.390 15.270 11.600 15.480 ;
        RECT 13.300 14.930 13.620 15.250 ;
        RECT 11.140 14.220 11.460 14.540 ;
        RECT 10.990 13.390 11.310 13.710 ;
        RECT 14.530 13.270 14.720 13.320 ;
        RECT 14.970 13.270 15.250 16.250 ;
        RECT 17.100 16.000 17.420 16.080 ;
        RECT 17.100 15.760 17.670 16.000 ;
        RECT 17.330 15.430 17.670 15.760 ;
        RECT 17.050 15.110 17.670 15.430 ;
        RECT 17.330 14.160 17.670 15.110 ;
        RECT 17.050 13.840 17.670 14.160 ;
        RECT 16.000 13.370 16.260 13.630 ;
        RECT 17.330 13.510 17.670 13.840 ;
        RECT 18.000 15.670 18.270 15.990 ;
        RECT 18.760 15.720 19.080 16.040 ;
        RECT 18.000 15.380 18.310 15.670 ;
        RECT 18.000 14.640 18.270 15.380 ;
        RECT 18.890 15.290 19.130 15.670 ;
        RECT 19.320 14.860 19.480 15.880 ;
        RECT 18.000 14.350 18.380 14.640 ;
        RECT 19.280 14.620 19.510 14.860 ;
        RECT 19.280 14.610 19.520 14.620 ;
        RECT 18.000 14.310 18.270 14.350 ;
        RECT 19.270 14.340 19.520 14.610 ;
        RECT 19.290 14.310 19.510 14.340 ;
        RECT 18.000 13.670 18.320 14.310 ;
        RECT 17.100 13.190 17.670 13.510 ;
        RECT 17.770 13.520 18.320 13.670 ;
        RECT 17.770 13.230 18.270 13.520 ;
        RECT 18.810 13.500 19.130 13.820 ;
        RECT 17.330 13.080 17.670 13.190 ;
        RECT 17.100 12.760 17.670 13.080 ;
        RECT 2.790 11.450 3.170 12.460 ;
        RECT 17.330 12.430 17.670 12.760 ;
        RECT 17.050 12.110 17.670 12.430 ;
        RECT 17.330 11.160 17.670 12.110 ;
        RECT 17.050 10.840 17.670 11.160 ;
        RECT 12.550 10.300 12.870 10.620 ;
        RECT 17.330 10.510 17.670 10.840 ;
        RECT 17.100 10.280 17.670 10.510 ;
        RECT 18.000 12.670 18.270 13.230 ;
        RECT 18.800 12.780 19.120 13.100 ;
        RECT 19.290 12.860 19.480 14.310 ;
        RECT 19.730 14.190 19.890 15.880 ;
        RECT 19.730 14.100 19.900 14.190 ;
        RECT 19.620 14.050 19.900 14.100 ;
        RECT 19.620 13.500 19.890 14.050 ;
        RECT 19.730 12.860 19.890 13.500 ;
        RECT 18.000 12.380 18.310 12.670 ;
        RECT 18.000 12.050 18.270 12.380 ;
        RECT 18.000 11.760 18.380 12.050 ;
        RECT 18.000 10.890 18.270 11.760 ;
        RECT 18.000 10.600 18.310 10.890 ;
        RECT 18.000 10.290 18.270 10.600 ;
        RECT 18.720 10.530 19.040 10.850 ;
        RECT 17.100 10.190 17.420 10.280 ;
        RECT 12.700 9.470 13.020 9.790 ;
        RECT 11.870 8.640 12.190 8.960 ;
        RECT 12.950 8.530 13.160 8.740 ;
        RECT 12.950 8.210 13.280 8.530 ;
        RECT 12.600 7.360 12.920 7.680 ;
        RECT 12.950 6.970 13.160 8.210 ;
        RECT 13.030 6.650 13.260 6.940 ;
      LAYER via ;
        RECT 13.330 17.720 13.590 17.980 ;
        RECT 11.070 16.360 11.330 16.620 ;
        RECT 14.220 16.560 14.480 16.820 ;
        RECT 17.800 18.950 18.060 19.210 ;
        RECT 15.160 16.280 15.420 16.540 ;
        RECT 14.220 15.960 14.480 16.220 ;
        RECT 11.460 15.510 11.720 15.770 ;
        RECT 10.340 15.080 10.600 15.340 ;
        RECT 13.330 14.960 13.590 15.220 ;
        RECT 11.170 14.250 11.430 14.510 ;
        RECT 11.020 13.420 11.280 13.680 ;
        RECT 17.130 15.790 17.390 16.050 ;
        RECT 17.080 15.140 17.340 15.400 ;
        RECT 17.080 13.870 17.340 14.130 ;
        RECT 18.790 15.750 19.050 16.010 ;
        RECT 17.130 13.220 17.390 13.480 ;
        RECT 17.800 13.380 18.060 13.640 ;
        RECT 18.840 13.530 19.100 13.790 ;
        RECT 17.130 12.790 17.390 13.050 ;
        RECT 2.830 11.490 3.120 12.420 ;
        RECT 17.080 12.140 17.340 12.400 ;
        RECT 17.080 10.870 17.340 11.130 ;
        RECT 12.580 10.330 12.840 10.590 ;
        RECT 17.130 10.220 17.390 10.480 ;
        RECT 18.830 12.810 19.090 13.070 ;
        RECT 18.750 10.560 19.010 10.820 ;
        RECT 12.730 9.500 12.990 9.760 ;
        RECT 11.900 8.670 12.160 8.930 ;
        RECT 13.020 8.240 13.280 8.500 ;
        RECT 12.630 7.390 12.890 7.650 ;
      LAYER met2 ;
        RECT 17.770 19.240 18.080 19.250 ;
        RECT 17.770 19.060 20.250 19.240 ;
        RECT 17.770 18.920 18.080 19.060 ;
        RECT 3.960 18.640 13.080 18.820 ;
        RECT 13.300 17.800 13.610 18.020 ;
        RECT 13.300 17.690 15.490 17.800 ;
        RECT 13.460 17.580 15.490 17.690 ;
        RECT 11.040 16.460 11.350 16.660 ;
        RECT 14.190 16.560 14.510 16.820 ;
        RECT 15.130 16.460 15.450 16.540 ;
        RECT 10.810 16.230 11.680 16.460 ;
        RECT 14.140 16.280 15.450 16.460 ;
        RECT 10.810 16.220 11.240 16.230 ;
        RECT 14.140 16.110 15.320 16.280 ;
        RECT 14.190 15.960 14.510 16.110 ;
        RECT 17.100 15.800 17.410 16.090 ;
        RECT 18.760 15.800 19.070 16.050 ;
        RECT 11.430 15.680 11.750 15.770 ;
        RECT 16.380 15.720 19.070 15.800 ;
        RECT 11.290 15.430 11.760 15.680 ;
        RECT 16.380 15.570 18.920 15.720 ;
        RECT 10.310 15.050 10.620 15.380 ;
        RECT 16.610 15.000 16.940 15.210 ;
        RECT 17.050 15.110 17.360 15.440 ;
        RECT 11.110 14.400 11.660 14.650 ;
        RECT 11.150 14.210 11.460 14.400 ;
        RECT 13.020 13.940 13.180 13.960 ;
        RECT 3.960 13.890 13.180 13.940 ;
        RECT 3.960 13.790 13.060 13.890 ;
        RECT 10.570 13.540 11.450 13.790 ;
        RECT 14.490 13.780 14.740 14.150 ;
        RECT 16.610 14.060 16.940 14.270 ;
        RECT 17.050 13.830 17.360 14.160 ;
        RECT 15.960 13.580 16.300 13.670 ;
        RECT 17.770 13.660 18.080 13.670 ;
        RECT 18.810 13.660 19.120 13.830 ;
        RECT 11.000 13.380 11.310 13.540 ;
        RECT 11.450 13.290 13.110 13.510 ;
        RECT 13.610 13.390 16.300 13.580 ;
        RECT 16.640 13.530 19.290 13.660 ;
        RECT 16.640 13.430 20.250 13.530 ;
        RECT 13.610 12.820 13.800 13.390 ;
        RECT 15.960 13.340 16.300 13.390 ;
        RECT 14.520 12.930 14.730 13.220 ;
        RECT 17.100 13.180 17.410 13.430 ;
        RECT 17.770 13.350 20.250 13.430 ;
        RECT 17.770 13.340 18.080 13.350 ;
        RECT 17.100 12.830 17.410 13.090 ;
        RECT 18.800 12.830 19.110 13.110 ;
        RECT 2.820 12.630 13.800 12.820 ;
        RECT 2.820 12.450 3.010 12.630 ;
        RECT 16.380 12.610 19.290 12.830 ;
        RECT 2.800 11.460 3.150 12.450 ;
        RECT 16.610 12.000 16.940 12.210 ;
        RECT 17.050 12.110 17.360 12.440 ;
        RECT 16.610 11.060 16.940 11.270 ;
        RECT 12.960 10.850 14.730 11.050 ;
        RECT 17.050 10.830 17.360 11.160 ;
        RECT 11.390 10.360 11.550 10.760 ;
        RECT 18.720 10.670 19.030 10.860 ;
        RECT 12.560 10.470 12.870 10.630 ;
        RECT 12.130 10.250 13.010 10.470 ;
        RECT 16.370 10.440 19.080 10.670 ;
        RECT 12.130 10.220 14.730 10.250 ;
        RECT 12.670 10.040 14.730 10.220 ;
        RECT 17.100 10.180 17.410 10.440 ;
        RECT 12.710 9.610 13.020 9.800 ;
        RECT 12.670 9.360 13.220 9.610 ;
        RECT 11.870 8.630 12.180 8.960 ;
        RECT 12.850 8.330 13.320 8.580 ;
        RECT 12.990 8.240 13.310 8.330 ;
        RECT 12.370 7.780 12.800 7.790 ;
        RECT 12.370 7.550 13.240 7.780 ;
        RECT 12.600 7.350 12.910 7.550 ;
  END
END sky130_hilas_TA2Cell_NoFG

MACRO sky130_hilas_TopLevelTextStructure
  CLASS CORE ;
  FOREIGN sky130_hilas_TopLevelTextStructure ;
  ORIGIN 0.000 0.000 ;
  SIZE 135.730 BY 78.160 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DIG24 
    ANTENNADIFFAREA 0.272000 ;
    PORT
      LAYER nwell ;
        RECT 78.830 32.310 81.390 34.220 ;
      LAYER met2 ;
        RECT 79.210 32.760 79.530 32.810 ;
        RECT 74.430 32.600 79.530 32.760 ;
        RECT 79.210 32.550 79.530 32.600 ;
        RECT 79.190 23.140 135.730 23.640 ;
        RECT 133.720 3.140 135.730 23.140 ;
        RECT 133.690 2.560 135.730 3.140 ;
        RECT 133.690 2.490 135.720 2.560 ;
    END
  END DIG24 
  PIN DIG23
    PORT
      LAYER met2 ;
        RECT 78.690 31.830 79.010 31.880 ;
        RECT 74.430 31.670 79.010 31.830 ;
        RECT 78.690 31.620 79.010 31.670 ;
        RECT 129.630 22.740 131.640 22.760 ;
        RECT 78.650 22.240 131.640 22.740 ;
        RECT 129.630 3.120 131.640 22.240 ;
        RECT 129.630 2.470 131.670 3.120 ;
        RECT 129.630 2.390 131.640 2.470 ;
    END
  END DIG23
  PIN DIG22
    PORT
      LAYER met2 ;
        RECT 78.220 29.990 78.540 30.040 ;
        RECT 74.430 29.830 78.540 29.990 ;
        RECT 78.220 29.780 78.540 29.830 ;
        RECT 78.180 21.820 127.450 21.840 ;
        RECT 78.180 21.340 127.560 21.820 ;
        RECT 125.550 3.140 127.560 21.340 ;
        RECT 125.550 2.490 127.620 3.140 ;
        RECT 125.550 2.450 127.560 2.490 ;
    END
  END DIG22
  PIN DIG21
    PORT
      LAYER met2 ;
        RECT 77.720 29.060 78.040 29.110 ;
        RECT 74.430 28.900 78.040 29.060 ;
        RECT 77.720 28.850 78.040 28.900 ;
        RECT 77.700 20.930 123.490 20.940 ;
        RECT 77.700 20.440 123.700 20.930 ;
        RECT 121.690 3.140 123.700 20.440 ;
        RECT 121.630 2.620 123.700 3.140 ;
        RECT 121.630 2.490 123.660 2.620 ;
    END
  END DIG21
  PIN DIG29
    PORT
      LAYER met2 ;
        RECT 113.440 3.840 113.630 4.010 ;
        RECT 113.440 3.650 118.440 3.840 ;
        RECT 118.250 3.190 118.440 3.650 ;
        RECT 118.250 3.120 119.280 3.190 ;
        RECT 117.580 2.470 119.610 3.120 ;
    END
  END DIG29
  PIN DIG28
    PORT
      LAYER met2 ;
        RECT 112.470 3.050 112.680 4.030 ;
        RECT 113.600 3.050 115.630 3.140 ;
        RECT 112.470 2.840 115.630 3.050 ;
        RECT 113.600 2.490 115.630 2.840 ;
    END
  END DIG28
  PIN DIG27
    PORT
      LAYER met2 ;
        RECT 110.540 3.140 110.750 4.030 ;
        RECT 109.420 2.490 111.450 3.140 ;
    END
  END DIG27
  PIN DIG26
    ANTENNAGATEAREA 53.084400 ;
    ANTENNADIFFAREA 276.667206 ;
    PORT
      LAYER nwell ;
        RECT 85.700 72.650 87.430 72.990 ;
        RECT 85.700 71.090 87.450 72.650 ;
        RECT 85.720 69.460 87.450 71.090 ;
        RECT 85.660 66.290 88.970 69.460 ;
        RECT 124.540 66.620 126.270 66.960 ;
        RECT 85.950 65.640 87.700 66.290 ;
        RECT 85.660 63.430 88.970 65.640 ;
        RECT 124.520 65.060 126.270 66.620 ;
        RECT 124.520 64.700 126.250 65.060 ;
        RECT 123.630 64.690 126.250 64.700 ;
        RECT 124.520 63.430 126.250 64.690 ;
        RECT 85.660 61.350 89.220 63.430 ;
        RECT 85.910 60.260 89.220 61.350 ;
        RECT 123.000 63.040 126.310 63.430 ;
        RECT 123.000 63.000 126.550 63.040 ;
        RECT 123.000 61.350 126.560 63.000 ;
        RECT 123.000 60.260 126.310 61.350 ;
        RECT 123.420 59.610 124.700 60.260 ;
        RECT 85.910 58.420 89.220 59.610 ;
        RECT 85.660 56.770 89.220 58.420 ;
        RECT 113.850 57.710 116.610 58.480 ;
        RECT 123.000 58.420 126.310 59.610 ;
        RECT 113.850 57.540 115.840 57.710 ;
        RECT 113.850 56.920 115.830 57.540 ;
        RECT 123.000 57.160 126.560 58.420 ;
        RECT 122.290 57.090 126.560 57.160 ;
        RECT 116.140 56.920 117.280 56.960 ;
        RECT 113.850 56.870 117.280 56.920 ;
        RECT 85.670 56.730 89.220 56.770 ;
        RECT 21.960 53.640 23.990 56.610 ;
        RECT 85.910 56.440 89.220 56.730 ;
        RECT 116.140 56.370 117.280 56.870 ;
        RECT 123.000 56.770 126.560 57.090 ;
        RECT 123.000 56.730 126.550 56.770 ;
        RECT 123.000 56.440 126.310 56.730 ;
        RECT 115.650 56.360 117.280 56.370 ;
        RECT 113.850 55.530 117.280 56.360 ;
        RECT 113.850 55.520 115.840 55.530 ;
        RECT 113.850 54.510 116.610 55.520 ;
        RECT 113.850 54.500 115.840 54.510 ;
        RECT 113.850 53.670 117.280 54.500 ;
        RECT 115.650 53.660 117.280 53.670 ;
        RECT 22.780 53.530 23.320 53.640 ;
        RECT 22.600 53.080 23.320 53.530 ;
        RECT 116.140 53.160 117.280 53.660 ;
        RECT 20.750 52.900 23.320 53.080 ;
        RECT 113.850 53.110 117.280 53.160 ;
        RECT 123.420 53.110 124.700 55.950 ;
        RECT 113.850 52.490 115.830 53.110 ;
        RECT 116.140 53.070 117.280 53.110 ;
        RECT 113.850 52.320 115.840 52.490 ;
        RECT 113.850 51.550 116.610 52.320 ;
        RECT 49.810 27.890 52.310 33.210 ;
        RECT 49.810 27.690 52.340 27.890 ;
        RECT 49.810 26.210 52.310 27.690 ;
        RECT 113.340 4.650 114.690 20.120 ;
        RECT 113.330 4.180 114.690 4.650 ;
      LAYER met3 ;
        RECT 82.710 57.250 83.160 58.000 ;
        RECT 82.710 51.090 83.080 57.250 ;
        RECT 83.750 57.240 84.200 57.990 ;
        RECT 83.830 54.600 84.200 57.240 ;
        RECT 83.830 54.000 84.270 54.600 ;
        RECT 82.710 50.760 83.200 51.090 ;
        RECT 82.760 50.600 83.200 50.760 ;
        RECT 83.830 48.890 84.200 54.000 ;
        RECT 83.820 48.020 84.290 48.890 ;
    END
  END DIG26
  PIN DIG25
    ANTENNAGATEAREA 53.084400 ;
    ANTENNADIFFAREA 253.798294 ;
    PORT
      LAYER met2 ;
        RECT 6.250 72.770 6.930 73.990 ;
        RECT 7.480 72.770 7.930 72.870 ;
        RECT 6.250 72.540 7.930 72.770 ;
        RECT 6.250 71.670 6.930 72.540 ;
        RECT 7.480 72.440 7.930 72.540 ;
        RECT 7.580 68.970 8.010 69.440 ;
        RECT 7.580 68.960 9.520 68.970 ;
        RECT 7.670 68.740 9.520 68.960 ;
        RECT 44.970 63.710 45.270 63.770 ;
        RECT 86.290 63.710 86.590 63.740 ;
        RECT 44.970 63.480 86.660 63.710 ;
        RECT 44.970 63.450 45.270 63.480 ;
        RECT 86.290 63.400 86.590 63.480 ;
        RECT 87.830 63.200 88.140 63.340 ;
        RECT 37.890 63.050 38.200 63.070 ;
        RECT 28.100 62.970 28.420 62.980 ;
        RECT 37.890 62.970 38.210 63.050 ;
        RECT 85.660 63.020 88.140 63.200 ;
        RECT 87.830 63.010 88.140 63.020 ;
        RECT 62.070 62.980 62.390 63.000 ;
        RECT 62.070 62.970 62.400 62.980 ;
        RECT 68.840 62.970 69.160 63.000 ;
        RECT 83.610 62.970 83.930 62.990 ;
        RECT 98.270 62.970 98.830 63.110 ;
        RECT 28.100 62.740 98.830 62.970 ;
        RECT 28.100 62.660 28.420 62.740 ;
        RECT 37.890 62.730 38.200 62.740 ;
        RECT 62.070 62.720 62.400 62.740 ;
        RECT 68.840 62.720 69.160 62.740 ;
        RECT 83.610 62.730 83.930 62.740 ;
        RECT 85.910 62.700 88.390 62.740 ;
        RECT 33.890 62.520 34.260 62.580 ;
        RECT 48.700 62.520 48.960 62.590 ;
        RECT 88.080 62.560 88.390 62.700 ;
        RECT 98.270 62.600 98.830 62.740 ;
        RECT 97.090 62.520 97.630 62.540 ;
        RECT 33.890 62.460 97.630 62.520 ;
        RECT 112.170 62.470 120.160 62.670 ;
        RECT 33.890 62.290 102.200 62.460 ;
        RECT 33.890 62.230 34.260 62.290 ;
        RECT 36.720 62.060 37.030 62.070 ;
        RECT 48.700 62.060 48.960 62.290 ;
        RECT 93.080 62.280 102.200 62.290 ;
        RECT 49.620 62.080 49.940 62.090 ;
        RECT 49.610 62.070 49.940 62.080 ;
        RECT 50.650 62.070 50.970 62.120 ;
        RECT 65.690 62.070 65.970 62.080 ;
        RECT 49.610 62.060 52.280 62.070 ;
        RECT 65.670 62.060 65.990 62.070 ;
        RECT 68.400 62.060 68.720 62.090 ;
        RECT 82.720 62.060 83.040 62.120 ;
        RECT 96.010 62.060 96.550 62.070 ;
        RECT 36.720 61.830 96.550 62.060 ;
        RECT 97.090 61.980 97.630 62.280 ;
        RECT 36.720 61.800 37.050 61.830 ;
        RECT 36.720 61.780 37.030 61.800 ;
        RECT 48.700 61.790 48.960 61.830 ;
        RECT 49.610 61.820 49.940 61.830 ;
        RECT 49.620 61.800 49.940 61.820 ;
        RECT 50.700 61.790 51.040 61.830 ;
        RECT 65.670 61.810 65.990 61.830 ;
        RECT 68.400 61.810 68.720 61.830 ;
        RECT 65.690 61.800 65.970 61.810 ;
        RECT 30.640 61.600 30.960 61.610 ;
        RECT 46.430 61.600 46.890 61.750 ;
        RECT 48.600 61.600 51.040 61.790 ;
        RECT 52.220 61.600 52.380 61.630 ;
        RECT 92.550 61.600 92.860 61.660 ;
        RECT 95.070 61.600 95.600 61.630 ;
        RECT 30.640 61.430 95.600 61.600 ;
        RECT 96.010 61.510 96.550 61.830 ;
        RECT 118.760 61.790 118.980 61.800 ;
        RECT 112.180 61.540 119.010 61.790 ;
        RECT 119.940 61.750 120.160 62.470 ;
        RECT 119.910 61.710 120.160 61.750 ;
        RECT 5.760 61.370 6.270 61.390 ;
        RECT 25.400 61.370 25.800 61.380 ;
        RECT 5.760 61.020 25.800 61.370 ;
        RECT 30.640 61.370 102.200 61.430 ;
        RECT 30.640 61.310 30.960 61.370 ;
        RECT 90.670 61.220 102.200 61.370 ;
        RECT 91.980 61.210 102.200 61.220 ;
        RECT 95.070 61.020 95.600 61.210 ;
        RECT 5.760 60.980 6.270 61.020 ;
        RECT 25.400 60.990 25.800 61.020 ;
        RECT 48.700 60.040 48.960 60.840 ;
        RECT 112.180 60.620 115.690 60.810 ;
        RECT 49.620 60.330 49.940 60.340 ;
        RECT 49.610 60.320 49.940 60.330 ;
        RECT 50.650 60.320 50.970 60.370 ;
        RECT 49.610 60.120 52.280 60.320 ;
        RECT 49.610 60.070 49.940 60.120 ;
        RECT 50.650 60.110 50.970 60.120 ;
        RECT 49.620 60.050 49.940 60.070 ;
        RECT 50.700 60.040 51.040 60.100 ;
        RECT 46.430 59.680 46.890 60.000 ;
        RECT 48.600 59.820 51.040 60.040 ;
        RECT 114.820 60.020 115.140 60.150 ;
        RECT 115.460 60.020 115.690 60.620 ;
        RECT 118.720 60.370 119.010 61.540 ;
        RECT 119.360 61.440 119.670 61.660 ;
        RECT 119.910 61.440 120.170 61.710 ;
        RECT 119.360 61.330 121.550 61.440 ;
        RECT 119.520 61.220 121.550 61.330 ;
        RECT 119.910 61.070 120.170 61.220 ;
        RECT 119.910 60.860 124.040 61.070 ;
        RECT 120.250 60.370 120.570 60.460 ;
        RECT 120.940 60.370 121.800 60.860 ;
        RECT 123.830 60.720 124.040 60.860 ;
        RECT 123.830 60.510 125.840 60.720 ;
        RECT 118.720 60.150 121.800 60.370 ;
        RECT 118.720 60.140 119.010 60.150 ;
        RECT 117.050 60.020 117.370 60.140 ;
        RECT 120.940 60.100 121.800 60.150 ;
        RECT 123.400 60.140 123.710 60.300 ;
        RECT 114.040 59.870 115.920 60.020 ;
        RECT 116.910 59.880 117.370 60.020 ;
        RECT 120.200 59.920 121.800 60.100 ;
        RECT 122.970 59.920 123.850 60.140 ;
        RECT 116.910 59.870 117.280 59.880 ;
        RECT 119.830 59.870 125.830 59.920 ;
        RECT 114.040 59.820 125.830 59.870 ;
        RECT 115.460 59.720 125.830 59.820 ;
        RECT 115.460 59.710 125.700 59.720 ;
        RECT 115.460 59.650 120.220 59.710 ;
        RECT 120.250 59.600 120.570 59.710 ;
        RECT 120.940 59.440 121.800 59.710 ;
        RECT 121.900 59.440 122.210 59.710 ;
        RECT 123.560 59.470 123.870 59.690 ;
        RECT 123.550 59.440 123.870 59.470 ;
        RECT 120.940 59.360 123.870 59.440 ;
        RECT 20.980 58.360 21.290 58.390 ;
        RECT 25.780 58.360 26.070 58.380 ;
        RECT 13.330 57.960 26.090 58.360 ;
        RECT 48.700 58.290 48.960 59.090 ;
        RECT 114.510 59.040 114.820 59.320 ;
        RECT 114.040 59.000 114.820 59.040 ;
        RECT 115.650 59.040 115.870 59.050 ;
        RECT 116.180 59.040 116.490 59.320 ;
        RECT 120.940 59.280 123.860 59.360 ;
        RECT 120.940 59.210 124.060 59.280 ;
        RECT 115.650 59.000 117.280 59.040 ;
        RECT 120.940 59.000 121.800 59.210 ;
        RECT 121.850 59.000 122.160 59.080 ;
        RECT 123.510 59.030 124.060 59.210 ;
        RECT 125.270 59.000 125.590 59.150 ;
        RECT 92.590 58.960 93.020 58.980 ;
        RECT 109.080 58.960 125.590 59.000 ;
        RECT 92.590 58.900 125.590 58.960 ;
        RECT 92.550 58.850 125.590 58.900 ;
        RECT 92.550 58.840 121.800 58.850 ;
        RECT 92.550 58.680 121.740 58.840 ;
        RECT 121.850 58.750 122.160 58.850 ;
        RECT 90.670 58.640 121.740 58.680 ;
        RECT 49.620 58.580 49.940 58.590 ;
        RECT 49.610 58.570 49.940 58.580 ;
        RECT 50.650 58.570 50.970 58.620 ;
        RECT 90.670 58.590 121.690 58.640 ;
        RECT 49.610 58.370 52.280 58.570 ;
        RECT 90.670 58.500 102.200 58.590 ;
        RECT 117.070 58.500 117.390 58.590 ;
        RECT 90.670 58.470 117.390 58.500 ;
        RECT 91.980 58.460 117.390 58.470 ;
        RECT 49.610 58.320 49.940 58.370 ;
        RECT 50.650 58.360 50.970 58.370 ;
        RECT 49.620 58.300 49.940 58.320 ;
        RECT 50.700 58.290 51.040 58.350 ;
        RECT 94.870 58.320 117.390 58.460 ;
        RECT 118.190 58.400 118.500 58.590 ;
        RECT 119.360 58.570 121.550 58.590 ;
        RECT 119.510 58.470 121.550 58.570 ;
        RECT 5.770 55.270 7.040 56.140 ;
        RECT 13.330 55.270 13.730 57.960 ;
        RECT 21.860 57.900 22.460 57.960 ;
        RECT 23.720 57.910 23.940 57.960 ;
        RECT 25.780 57.950 26.070 57.960 ;
        RECT 46.430 57.930 46.890 58.250 ;
        RECT 48.600 58.070 51.040 58.290 ;
        RECT 82.660 57.650 83.240 58.090 ;
        RECT 82.660 57.460 83.300 57.650 ;
        RECT 25.790 57.060 26.110 57.110 ;
        RECT 25.220 56.890 26.170 57.060 ;
        RECT 25.790 56.850 26.110 56.890 ;
        RECT 22.020 56.640 22.340 56.690 ;
        RECT 22.660 56.640 23.480 56.720 ;
        RECT 22.020 56.550 23.480 56.640 ;
        RECT 22.020 56.470 22.760 56.550 ;
        RECT 48.700 56.540 48.960 57.340 ;
        RECT 49.620 56.830 49.940 56.840 ;
        RECT 49.610 56.820 49.940 56.830 ;
        RECT 50.650 56.820 50.970 56.870 ;
        RECT 83.060 56.850 83.300 57.460 ;
        RECT 83.680 57.450 84.260 58.080 ;
        RECT 99.840 58.050 100.150 58.320 ;
        RECT 114.110 58.210 114.430 58.320 ;
        RECT 86.500 57.940 86.970 58.000 ;
        RECT 100.250 57.940 102.200 58.150 ;
        RECT 113.730 58.140 114.430 58.210 ;
        RECT 111.100 57.940 111.150 58.060 ;
        RECT 113.730 58.010 114.340 58.140 ;
        RECT 123.690 58.000 124.160 58.250 ;
        RECT 111.400 57.950 111.690 57.960 ;
        RECT 111.400 57.940 111.700 57.950 ;
        RECT 121.930 57.940 122.380 57.960 ;
        RECT 86.500 57.510 122.390 57.940 ;
        RECT 123.830 57.910 124.150 58.000 ;
        RECT 93.100 57.430 102.200 57.510 ;
        RECT 103.530 57.390 104.370 57.510 ;
        RECT 110.020 57.430 119.120 57.510 ;
        RECT 119.250 57.430 119.520 57.510 ;
        RECT 121.850 57.470 122.160 57.510 ;
        RECT 123.610 57.460 123.920 57.470 ;
        RECT 123.210 57.450 123.920 57.460 ;
        RECT 123.210 57.310 124.080 57.450 ;
        RECT 123.210 57.300 124.140 57.310 ;
        RECT 114.600 57.230 115.720 57.240 ;
        RECT 113.730 57.140 115.720 57.230 ;
        RECT 103.980 57.030 115.720 57.140 ;
        RECT 121.440 57.170 124.140 57.300 ;
        RECT 121.440 57.070 126.310 57.170 ;
        RECT 103.980 56.920 114.120 57.030 ;
        RECT 114.600 57.020 115.720 57.030 ;
        RECT 111.100 56.880 111.160 56.920 ;
        RECT 113.900 56.820 114.120 56.920 ;
        RECT 114.820 56.820 115.140 56.950 ;
        RECT 117.050 56.820 117.370 56.940 ;
        RECT 49.610 56.620 52.280 56.820 ;
        RECT 107.580 56.650 107.880 56.670 ;
        RECT 113.900 56.650 115.920 56.820 ;
        RECT 116.910 56.680 117.370 56.820 ;
        RECT 119.320 56.860 119.520 56.870 ;
        RECT 116.910 56.650 117.280 56.680 ;
        RECT 119.320 56.650 119.540 56.860 ;
        RECT 121.430 56.830 121.790 56.840 ;
        RECT 120.870 56.650 121.790 56.830 ;
        RECT 121.900 56.820 122.210 57.070 ;
        RECT 123.440 57.020 123.750 57.070 ;
        RECT 123.830 56.990 126.310 57.070 ;
        RECT 123.830 56.980 124.140 56.990 ;
        RECT 49.610 56.570 49.940 56.620 ;
        RECT 50.650 56.610 50.970 56.620 ;
        RECT 49.620 56.550 49.940 56.570 ;
        RECT 50.700 56.540 51.040 56.600 ;
        RECT 22.020 56.430 22.340 56.470 ;
        RECT 22.440 56.260 22.750 56.470 ;
        RECT 25.790 56.140 26.110 56.190 ;
        RECT 46.430 56.180 46.890 56.500 ;
        RECT 48.600 56.320 51.040 56.540 ;
        RECT 107.570 56.550 121.790 56.650 ;
        RECT 107.570 56.470 121.830 56.550 ;
        RECT 121.900 56.470 122.210 56.730 ;
        RECT 123.600 56.470 123.910 56.750 ;
        RECT 107.570 56.250 124.090 56.470 ;
        RECT 107.570 56.230 121.830 56.250 ;
        RECT 107.580 56.210 107.880 56.230 ;
        RECT 111.100 56.170 111.160 56.230 ;
        RECT 113.900 56.200 114.120 56.230 ;
        RECT 114.600 56.200 115.720 56.210 ;
        RECT 25.220 55.970 26.170 56.140 ;
        RECT 25.790 55.930 26.110 55.970 ;
        RECT 103.930 55.950 112.940 56.170 ;
        RECT 113.730 56.000 115.720 56.200 ;
        RECT 115.790 56.150 115.860 56.230 ;
        RECT 21.960 55.720 22.340 55.910 ;
        RECT 22.530 55.720 22.850 55.880 ;
        RECT 21.990 55.650 22.850 55.720 ;
        RECT 21.990 55.550 23.480 55.650 ;
        RECT 21.990 55.510 22.310 55.550 ;
        RECT 22.440 55.450 23.480 55.550 ;
        RECT 22.440 55.270 22.750 55.450 ;
        RECT 5.770 54.870 13.730 55.270 ;
        RECT 25.760 55.220 26.080 55.270 ;
        RECT 25.220 55.050 26.170 55.220 ;
        RECT 25.760 55.010 26.080 55.050 ;
        RECT 5.770 54.260 7.040 54.870 ;
        RECT 21.960 54.800 22.340 54.920 ;
        RECT 22.530 54.800 22.850 54.890 ;
        RECT 21.960 54.730 22.850 54.800 ;
        RECT 22.000 54.690 22.850 54.730 ;
        RECT 22.000 54.630 23.480 54.690 ;
        RECT 22.000 54.590 22.320 54.630 ;
        RECT 22.530 54.610 23.480 54.630 ;
        RECT 22.440 54.490 23.480 54.610 ;
        RECT 22.440 54.280 22.750 54.490 ;
        RECT 92.960 54.410 102.110 54.640 ;
        RECT 101.820 54.310 102.110 54.410 ;
        RECT 103.980 54.310 109.640 54.390 ;
        RECT 109.800 54.310 110.940 54.390 ;
        RECT 101.820 54.190 110.940 54.310 ;
        RECT 112.720 54.340 112.940 55.950 ;
        RECT 113.900 55.840 114.120 56.000 ;
        RECT 114.510 55.990 115.720 56.000 ;
        RECT 114.510 55.840 114.820 55.990 ;
        RECT 120.870 55.890 121.830 56.230 ;
        RECT 113.900 55.790 114.820 55.840 ;
        RECT 113.900 55.720 114.610 55.790 ;
        RECT 113.870 55.640 114.610 55.720 ;
        RECT 113.870 55.220 114.130 55.640 ;
        RECT 113.730 55.200 114.340 55.220 ;
        RECT 113.730 55.040 114.430 55.200 ;
        RECT 113.730 55.020 118.000 55.040 ;
        RECT 113.870 55.010 118.000 55.020 ;
        RECT 113.730 54.830 118.000 55.010 ;
        RECT 113.730 54.810 114.340 54.830 ;
        RECT 117.790 54.690 118.000 54.830 ;
        RECT 117.790 54.480 119.810 54.690 ;
        RECT 120.930 54.460 121.830 55.890 ;
        RECT 121.850 55.750 122.160 56.080 ;
        RECT 121.850 54.470 122.160 54.800 ;
        RECT 114.040 54.340 114.610 54.390 ;
        RECT 101.820 54.110 110.150 54.190 ;
        RECT 112.720 54.120 115.570 54.340 ;
        RECT 123.520 54.310 123.830 54.500 ;
        RECT 101.820 54.100 102.110 54.110 ;
        RECT 21.350 53.790 21.670 53.830 ;
        RECT 21.960 53.790 22.340 53.930 ;
        RECT 22.530 53.790 22.850 53.900 ;
        RECT 21.350 53.730 22.850 53.790 ;
        RECT 109.420 53.840 109.640 54.110 ;
        RECT 114.510 54.040 114.820 54.120 ;
        RECT 117.360 54.110 117.670 54.270 ;
        RECT 114.510 54.030 115.720 54.040 ;
        RECT 113.730 53.890 115.720 54.030 ;
        RECT 116.930 53.890 117.810 54.110 ;
        RECT 121.170 54.080 123.880 54.310 ;
        RECT 111.100 53.840 111.160 53.880 ;
        RECT 113.730 53.840 119.810 53.890 ;
        RECT 21.350 53.600 23.480 53.730 ;
        RECT 109.420 53.680 119.810 53.840 ;
        RECT 121.900 53.820 122.210 54.080 ;
        RECT 109.420 53.620 114.180 53.680 ;
        RECT 21.350 53.570 21.670 53.600 ;
        RECT 22.530 53.580 23.480 53.600 ;
        RECT 22.670 53.530 23.480 53.580 ;
        RECT 114.040 53.350 117.280 53.410 ;
        RECT 114.040 53.210 117.370 53.350 ;
        RECT 108.810 52.970 109.130 52.980 ;
        RECT 111.100 52.970 111.160 53.150 ;
        RECT 114.820 53.080 115.140 53.210 ;
        RECT 115.300 53.130 117.010 53.210 ;
        RECT 114.600 53.000 115.720 53.010 ;
        RECT 113.730 52.970 115.720 53.000 ;
        RECT 115.790 52.970 115.860 53.130 ;
        RECT 116.810 52.970 117.010 53.130 ;
        RECT 117.050 53.090 117.370 53.210 ;
        RECT 119.250 52.970 119.580 53.110 ;
        RECT 21.310 52.830 21.630 52.870 ;
        RECT 21.310 52.640 22.780 52.830 ;
        RECT 108.810 52.810 119.580 52.970 ;
        RECT 108.810 52.800 109.500 52.810 ;
        RECT 113.730 52.800 115.720 52.810 ;
        RECT 104.580 52.680 104.940 52.780 ;
        RECT 108.810 52.680 109.130 52.800 ;
        RECT 114.600 52.790 115.720 52.800 ;
        RECT 116.810 52.680 117.010 52.810 ;
        RECT 21.310 52.610 21.630 52.640 ;
        RECT 104.580 52.480 110.940 52.680 ;
        RECT 115.300 52.480 117.010 52.680 ;
        RECT 104.580 52.360 104.940 52.480 ;
        RECT 116.670 52.270 117.010 52.480 ;
        RECT 21.350 51.870 21.670 51.910 ;
        RECT 21.350 51.680 22.780 51.870 ;
        RECT 21.350 51.650 21.670 51.680 ;
        RECT 116.810 51.430 117.010 52.270 ;
        RECT 120.900 51.430 121.800 52.100 ;
        RECT 65.670 51.400 65.980 51.410 ;
        RECT 65.660 51.340 65.990 51.400 ;
        RECT 65.310 51.290 65.990 51.340 ;
        RECT 62.080 51.120 65.990 51.290 ;
        RECT 115.650 51.190 115.870 51.200 ;
        RECT 116.810 51.190 121.800 51.430 ;
        RECT 62.080 51.070 65.980 51.120 ;
        RECT 115.650 51.000 121.800 51.190 ;
        RECT 115.650 50.990 117.280 51.000 ;
        RECT 117.400 50.990 117.710 51.000 ;
        RECT 115.650 50.980 115.870 50.990 ;
        RECT 116.180 50.710 116.490 50.990 ;
        RECT 105.500 50.420 105.890 50.440 ;
        RECT 105.490 50.310 105.900 50.420 ;
        RECT 116.810 50.310 117.010 50.990 ;
        RECT 105.490 50.210 110.150 50.310 ;
        RECT 115.300 50.210 117.010 50.310 ;
        RECT 105.490 50.110 110.940 50.210 ;
        RECT 105.490 50.010 105.900 50.110 ;
        RECT 109.920 50.010 110.940 50.110 ;
        RECT 114.040 50.150 117.280 50.210 ;
        RECT 114.040 50.010 117.370 50.150 ;
        RECT 120.900 50.010 121.800 51.000 ;
        RECT 105.500 49.990 105.890 50.010 ;
        RECT 114.820 49.880 115.140 50.010 ;
        RECT 106.320 49.720 106.720 49.730 ;
        RECT 106.300 49.660 106.740 49.720 ;
        RECT 116.810 49.660 117.010 50.010 ;
        RECT 117.050 49.890 117.370 50.010 ;
        RECT 106.300 49.480 110.150 49.660 ;
        RECT 115.300 49.480 117.010 49.660 ;
        RECT 106.300 49.460 110.940 49.480 ;
        RECT 106.320 49.450 106.720 49.460 ;
        RECT 109.800 49.280 110.940 49.460 ;
        RECT 115.240 49.340 117.010 49.480 ;
        RECT 115.240 49.280 117.000 49.340 ;
        RECT 46.430 41.280 46.890 41.600 ;
        RECT 48.600 41.240 51.040 41.460 ;
        RECT 48.700 40.440 48.960 41.240 ;
        RECT 49.620 41.210 49.940 41.230 ;
        RECT 49.610 41.160 49.940 41.210 ;
        RECT 50.700 41.180 51.040 41.240 ;
        RECT 50.650 41.160 50.970 41.170 ;
        RECT 49.610 40.960 52.280 41.160 ;
        RECT 49.610 40.950 49.940 40.960 ;
        RECT 49.620 40.940 49.940 40.950 ;
        RECT 50.650 40.910 50.970 40.960 ;
        RECT 98.180 40.810 98.780 40.870 ;
        RECT 120.900 40.810 121.800 41.840 ;
        RECT 98.180 40.340 121.800 40.810 ;
        RECT 98.180 40.290 98.780 40.340 ;
        RECT 46.430 39.530 46.890 39.850 ;
        RECT 120.900 39.750 121.800 40.340 ;
        RECT 48.600 39.490 51.040 39.710 ;
        RECT 48.700 38.690 48.960 39.490 ;
        RECT 49.620 39.460 49.940 39.480 ;
        RECT 49.610 39.410 49.940 39.460 ;
        RECT 50.700 39.430 51.040 39.490 ;
        RECT 50.650 39.410 50.970 39.420 ;
        RECT 49.610 39.210 52.280 39.410 ;
        RECT 49.610 39.200 49.940 39.210 ;
        RECT 49.620 39.190 49.940 39.200 ;
        RECT 50.650 39.160 50.970 39.210 ;
        RECT 46.430 37.780 46.890 38.100 ;
        RECT 48.600 37.740 51.040 37.960 ;
        RECT 48.700 36.940 48.960 37.740 ;
        RECT 49.620 37.710 49.940 37.730 ;
        RECT 49.610 37.660 49.940 37.710 ;
        RECT 50.700 37.680 51.040 37.740 ;
        RECT 50.650 37.660 50.970 37.670 ;
        RECT 49.610 37.460 52.280 37.660 ;
        RECT 49.610 37.450 49.940 37.460 ;
        RECT 49.620 37.440 49.940 37.450 ;
        RECT 50.650 37.410 50.970 37.460 ;
        RECT 21.310 36.840 21.620 36.860 ;
        RECT 21.970 36.840 22.280 36.860 ;
        RECT 21.310 36.370 28.630 36.840 ;
        RECT 21.310 36.350 21.620 36.370 ;
        RECT 21.970 36.350 22.280 36.370 ;
        RECT 28.160 35.690 28.630 36.370 ;
        RECT 54.930 36.700 55.240 36.720 ;
        RECT 78.830 36.710 81.000 36.730 ;
        RECT 78.830 36.700 81.160 36.710 ;
        RECT 81.300 36.700 81.390 36.730 ;
        RECT 81.720 36.700 81.810 36.710 ;
        RECT 92.570 36.700 93.020 36.730 ;
        RECT 46.430 36.030 46.890 36.350 ;
        RECT 54.930 36.290 93.020 36.700 ;
        RECT 54.930 36.270 55.240 36.290 ;
        RECT 48.600 35.990 51.040 36.210 ;
        RECT 78.830 36.160 81.010 36.290 ;
        RECT 92.570 36.270 93.020 36.290 ;
        RECT 78.830 36.120 81.160 36.160 ;
        RECT 48.700 35.690 48.960 35.990 ;
        RECT 49.620 35.960 49.940 35.980 ;
        RECT 49.610 35.910 49.940 35.960 ;
        RECT 50.700 35.930 51.040 35.990 ;
        RECT 50.650 35.910 50.970 35.920 ;
        RECT 49.610 35.710 52.280 35.910 ;
        RECT 80.850 35.830 81.160 36.120 ;
        RECT 78.830 35.790 81.160 35.830 ;
        RECT 49.610 35.700 49.940 35.710 ;
        RECT 49.620 35.690 49.940 35.700 ;
        RECT 50.650 35.690 50.970 35.710 ;
        RECT 78.830 35.690 81.010 35.790 ;
        RECT 120.930 35.690 121.830 36.660 ;
        RECT 19.980 35.560 20.240 35.630 ;
        RECT 22.030 35.560 22.350 35.580 ;
        RECT 23.790 35.560 24.120 35.600 ;
        RECT 19.980 35.370 24.120 35.560 ;
        RECT 19.980 35.310 20.240 35.370 ;
        RECT 22.030 35.320 22.350 35.370 ;
        RECT 23.790 35.330 24.120 35.370 ;
        RECT 28.160 35.220 121.830 35.690 ;
        RECT 19.430 35.160 19.750 35.200 ;
        RECT 21.370 35.160 21.690 35.220 ;
        RECT 24.290 35.160 24.610 35.200 ;
        RECT 48.700 35.190 48.960 35.220 ;
        RECT 19.430 34.970 24.610 35.160 ;
        RECT 97.090 35.100 97.660 35.220 ;
        RECT 19.430 34.940 19.750 34.970 ;
        RECT 21.370 34.960 21.690 34.970 ;
        RECT 24.290 34.940 24.610 34.970 ;
        RECT 25.770 34.600 26.070 34.620 ;
        RECT 25.760 34.580 26.080 34.600 ;
        RECT 23.540 34.360 26.080 34.580 ;
        RECT 120.930 34.570 121.830 35.220 ;
        RECT 23.540 33.920 23.760 34.360 ;
        RECT 25.760 34.340 26.080 34.360 ;
        RECT 25.770 34.320 26.070 34.340 ;
        RECT 25.150 33.450 25.440 33.470 ;
        RECT 25.140 33.420 25.460 33.450 ;
        RECT 24.900 33.410 26.890 33.420 ;
        RECT 23.570 33.220 26.890 33.410 ;
        RECT 27.740 33.310 28.430 33.390 ;
        RECT 24.900 33.200 26.890 33.220 ;
        RECT 25.140 33.190 25.460 33.200 ;
        RECT 25.150 33.170 25.440 33.190 ;
        RECT 27.580 33.180 28.430 33.310 ;
        RECT 27.580 32.980 27.890 33.180 ;
        RECT 96.030 33.160 96.340 33.420 ;
        RECT 95.880 33.000 98.470 33.160 ;
        RECT 25.710 32.540 26.020 32.870 ;
        RECT 95.880 32.830 96.190 33.000 ;
        RECT 95.880 32.570 96.190 32.740 ;
        RECT 46.390 32.220 46.850 32.540 ;
        RECT 95.880 32.410 98.470 32.570 ;
        RECT 48.560 32.180 51.000 32.400 ;
        RECT 19.460 31.290 19.750 31.300 ;
        RECT 19.450 31.270 19.770 31.290 ;
        RECT 25.210 31.280 25.530 31.540 ;
        RECT 48.660 31.380 48.920 32.180 ;
        RECT 49.580 32.150 49.900 32.170 ;
        RECT 49.570 32.100 49.900 32.150 ;
        RECT 50.660 32.120 51.000 32.180 ;
        RECT 96.030 32.150 96.340 32.410 ;
        RECT 96.670 32.250 97.930 32.410 ;
        RECT 50.610 32.100 50.930 32.110 ;
        RECT 49.570 31.900 52.240 32.100 ;
        RECT 49.570 31.890 49.900 31.900 ;
        RECT 49.580 31.880 49.900 31.890 ;
        RECT 50.610 31.850 50.930 31.900 ;
        RECT 19.450 31.050 20.450 31.270 ;
        RECT 19.450 31.030 19.770 31.050 ;
        RECT 27.610 31.040 27.930 31.070 ;
        RECT 19.460 31.010 19.750 31.030 ;
        RECT 24.900 30.860 27.930 31.040 ;
        RECT 24.720 30.830 27.930 30.860 ;
        RECT 24.720 30.810 25.040 30.830 ;
        RECT 23.550 30.640 25.040 30.810 ;
        RECT 27.610 30.750 27.930 30.830 ;
        RECT 23.550 30.600 27.880 30.640 ;
        RECT 24.720 30.560 27.880 30.600 ;
        RECT 24.900 30.530 27.880 30.560 ;
        RECT 24.900 30.430 27.940 30.530 ;
        RECT 46.390 30.470 46.850 30.790 ;
        RECT 48.560 30.430 51.000 30.650 ;
        RECT 96.030 30.460 96.340 30.650 ;
        RECT 27.620 30.210 27.940 30.430 ;
        RECT 25.210 29.730 25.530 29.990 ;
        RECT 48.660 29.630 48.920 30.430 ;
        RECT 49.580 30.400 49.900 30.420 ;
        RECT 49.570 30.350 49.900 30.400 ;
        RECT 50.660 30.370 51.000 30.430 ;
        RECT 95.970 30.450 96.520 30.460 ;
        RECT 95.970 30.430 96.530 30.450 ;
        RECT 96.670 30.430 97.930 30.570 ;
        RECT 120.900 30.430 121.800 31.580 ;
        RECT 95.970 30.390 121.800 30.430 ;
        RECT 50.610 30.350 50.930 30.360 ;
        RECT 49.570 30.150 52.240 30.350 ;
        RECT 49.570 30.140 49.900 30.150 ;
        RECT 49.580 30.130 49.900 30.140 ;
        RECT 50.610 30.100 50.930 30.150 ;
        RECT 95.880 30.080 121.800 30.390 ;
        RECT 91.130 29.960 121.800 30.080 ;
        RECT 91.130 29.910 97.810 29.960 ;
        RECT 95.880 29.800 96.190 29.910 ;
        RECT 97.480 29.880 97.810 29.910 ;
        RECT 95.880 29.640 98.470 29.800 ;
        RECT 96.030 29.380 96.340 29.640 ;
        RECT 96.690 29.480 97.930 29.640 ;
        RECT 120.900 29.490 121.800 29.960 ;
        RECT 25.740 28.660 26.050 28.990 ;
        RECT 46.390 28.720 46.850 29.040 ;
        RECT 48.560 28.680 51.000 28.900 ;
        RECT 19.240 28.220 21.950 28.230 ;
        RECT 19.010 27.900 21.950 28.220 ;
        RECT 19.010 27.750 19.630 27.900 ;
        RECT 20.420 27.760 20.730 27.900 ;
        RECT 21.510 27.760 21.820 27.900 ;
        RECT 48.660 27.880 48.920 28.680 ;
        RECT 49.580 28.650 49.900 28.670 ;
        RECT 49.570 28.600 49.900 28.650 ;
        RECT 50.660 28.620 51.000 28.680 ;
        RECT 50.610 28.600 50.930 28.610 ;
        RECT 49.570 28.400 52.240 28.600 ;
        RECT 49.570 28.390 49.900 28.400 ;
        RECT 49.580 28.380 49.900 28.390 ;
        RECT 50.610 28.350 50.930 28.400 ;
        RECT 19.010 26.280 19.360 27.750 ;
        RECT 101.160 27.620 101.720 27.690 ;
        RECT 113.880 27.620 114.560 27.680 ;
        RECT 121.410 27.620 122.070 28.260 ;
        RECT 19.980 27.410 23.140 27.550 ;
        RECT 19.870 27.230 23.140 27.410 ;
        RECT 52.220 27.360 52.550 27.380 ;
        RECT 52.210 27.290 52.560 27.360 ;
        RECT 19.870 27.080 20.180 27.230 ;
        RECT 20.970 27.080 21.280 27.230 ;
        RECT 22.070 27.080 22.380 27.230 ;
        RECT 22.820 26.280 23.140 27.230 ;
        RECT 46.390 26.970 46.850 27.290 ;
        RECT 52.180 27.280 52.560 27.290 ;
        RECT 57.960 27.280 58.280 27.340 ;
        RECT 48.560 26.930 51.000 27.150 ;
        RECT 52.180 27.120 58.280 27.280 ;
        RECT 101.160 27.210 122.070 27.620 ;
        RECT 101.160 27.160 101.720 27.210 ;
        RECT 113.880 27.150 114.560 27.210 ;
        RECT 52.180 27.090 52.560 27.120 ;
        RECT 52.210 27.050 52.560 27.090 ;
        RECT 57.960 27.070 58.280 27.120 ;
        RECT 121.410 27.110 122.070 27.210 ;
        RECT 47.790 26.660 48.120 26.900 ;
        RECT 48.660 26.660 48.920 26.930 ;
        RECT 49.580 26.900 49.900 26.920 ;
        RECT 49.570 26.850 49.900 26.900 ;
        RECT 50.660 26.870 51.000 26.930 ;
        RECT 50.610 26.850 50.930 26.860 ;
        RECT 49.570 26.660 52.240 26.850 ;
        RECT 53.650 26.790 53.950 26.800 ;
        RECT 53.640 26.660 53.960 26.790 ;
        RECT 64.180 26.660 64.460 26.960 ;
        RECT 68.210 26.660 68.510 26.940 ;
        RECT 47.790 26.640 68.510 26.660 ;
        RECT 47.790 26.610 68.500 26.640 ;
        RECT 47.790 26.500 68.440 26.610 ;
        RECT 48.660 26.280 48.920 26.500 ;
        RECT 51.600 26.280 52.040 26.290 ;
        RECT 6.280 26.270 52.040 26.280 ;
        RECT 6.280 25.860 52.060 26.270 ;
        RECT 19.010 25.460 19.360 25.860 ;
        RECT 19.870 25.710 20.180 25.860 ;
        RECT 20.970 25.710 21.280 25.860 ;
        RECT 22.070 25.710 22.380 25.860 ;
        RECT 19.010 25.310 21.960 25.460 ;
        RECT 22.820 25.310 23.140 25.860 ;
        RECT 44.750 25.850 45.230 25.860 ;
        RECT 51.580 25.850 52.060 25.860 ;
        RECT 51.600 25.840 52.040 25.850 ;
        RECT 6.260 24.890 48.240 25.310 ;
        RECT 94.920 25.130 95.520 25.180 ;
        RECT 121.330 25.130 123.430 26.070 ;
        RECT 19.010 24.260 19.360 24.890 ;
        RECT 19.010 24.130 19.390 24.260 ;
        RECT 19.010 24.090 19.760 24.130 ;
        RECT 19.010 23.790 21.950 24.090 ;
        RECT 19.310 23.640 19.620 23.790 ;
        RECT 20.420 23.630 20.730 23.790 ;
        RECT 21.510 23.610 21.820 23.790 ;
        RECT 22.820 23.410 23.140 24.890 ;
        RECT 29.310 24.390 30.140 24.890 ;
        RECT 94.920 24.660 123.430 25.130 ;
        RECT 94.920 24.620 95.520 24.660 ;
        RECT 121.330 23.990 123.430 24.660 ;
        RECT 121.350 23.980 122.120 23.990 ;
        RECT 19.990 23.270 23.140 23.410 ;
        RECT 19.870 23.080 23.140 23.270 ;
        RECT 19.870 23.070 23.050 23.080 ;
        RECT 19.870 22.940 20.180 23.070 ;
        RECT 20.970 22.930 21.280 23.070 ;
        RECT 22.060 22.930 22.370 23.070 ;
        RECT 22.900 22.870 23.190 22.890 ;
        RECT 25.130 22.870 25.440 22.890 ;
        RECT 22.890 22.510 25.440 22.870 ;
        RECT 22.900 22.490 23.190 22.510 ;
        RECT 25.130 22.490 25.440 22.510 ;
        RECT 52.550 21.980 52.860 22.120 ;
        RECT 53.640 21.980 53.950 22.120 ;
        RECT 54.740 21.980 55.050 22.110 ;
        RECT 51.870 21.970 55.050 21.980 ;
        RECT 51.780 21.780 55.050 21.970 ;
        RECT 58.590 21.980 58.900 22.110 ;
        RECT 59.690 21.980 60.000 22.120 ;
        RECT 60.780 21.980 61.090 22.120 ;
        RECT 62.360 22.010 62.670 22.150 ;
        RECT 63.450 22.010 63.760 22.150 ;
        RECT 64.550 22.010 64.860 22.140 ;
        RECT 61.680 22.000 64.860 22.010 ;
        RECT 61.590 21.980 64.860 22.000 ;
        RECT 58.590 21.810 64.860 21.980 ;
        RECT 68.400 22.010 68.710 22.140 ;
        RECT 69.500 22.010 69.810 22.150 ;
        RECT 70.590 22.010 70.900 22.150 ;
        RECT 68.400 22.000 71.580 22.010 ;
        RECT 68.400 21.810 71.670 22.000 ;
        RECT 58.590 21.780 64.740 21.810 ;
        RECT 51.780 21.640 54.930 21.780 ;
        RECT 58.710 21.670 64.740 21.780 ;
        RECT 68.520 21.670 71.670 21.810 ;
        RECT 74.140 21.990 74.450 22.120 ;
        RECT 75.240 21.990 75.550 22.130 ;
        RECT 76.330 21.990 76.640 22.130 ;
        RECT 74.140 21.980 77.320 21.990 ;
        RECT 74.140 21.790 77.410 21.980 ;
        RECT 58.710 21.640 61.910 21.670 ;
        RECT 19.280 20.660 21.990 20.670 ;
        RECT 19.050 20.340 21.990 20.660 ;
        RECT 19.050 20.190 19.670 20.340 ;
        RECT 20.460 20.200 20.770 20.340 ;
        RECT 21.550 20.200 21.860 20.340 ;
        RECT 19.050 17.900 19.400 20.190 ;
        RECT 20.020 19.850 23.180 19.990 ;
        RECT 19.910 19.670 23.180 19.850 ;
        RECT 19.910 19.520 20.220 19.670 ;
        RECT 21.010 19.520 21.320 19.670 ;
        RECT 22.110 19.520 22.420 19.670 ;
        RECT 22.860 19.210 23.180 19.670 ;
        RECT 25.760 19.210 26.040 19.220 ;
        RECT 22.170 18.880 26.060 19.210 ;
        RECT 51.780 19.190 52.100 21.640 ;
        RECT 53.100 21.260 53.410 21.440 ;
        RECT 54.190 21.260 54.500 21.420 ;
        RECT 55.300 21.260 55.610 21.410 ;
        RECT 58.030 21.260 58.340 21.410 ;
        RECT 59.140 21.260 59.450 21.420 ;
        RECT 60.230 21.260 60.540 21.440 ;
        RECT 52.970 20.960 55.910 21.260 ;
        RECT 55.160 20.920 55.910 20.960 ;
        RECT 55.530 20.790 55.910 20.920 ;
        RECT 55.560 20.070 55.910 20.790 ;
        RECT 57.730 20.960 60.670 21.260 ;
        RECT 57.730 20.920 58.480 20.960 ;
        RECT 57.730 20.790 58.110 20.920 ;
        RECT 57.730 20.360 58.080 20.790 ;
        RECT 61.540 20.360 61.910 21.640 ;
        RECT 62.910 21.290 63.220 21.470 ;
        RECT 64.000 21.290 64.310 21.450 ;
        RECT 65.110 21.290 65.420 21.440 ;
        RECT 67.840 21.290 68.150 21.440 ;
        RECT 68.950 21.290 69.260 21.450 ;
        RECT 70.040 21.290 70.350 21.470 ;
        RECT 62.780 20.990 65.720 21.290 ;
        RECT 64.970 20.950 65.720 20.990 ;
        RECT 65.340 20.820 65.720 20.950 ;
        RECT 65.370 20.360 65.720 20.820 ;
        RECT 67.540 20.990 70.480 21.290 ;
        RECT 67.540 20.950 68.290 20.990 ;
        RECT 67.540 20.820 67.920 20.950 ;
        RECT 56.290 20.330 67.190 20.360 ;
        RECT 53.100 19.920 53.410 20.070 ;
        RECT 54.190 19.920 54.500 20.070 ;
        RECT 55.290 19.920 55.910 20.070 ;
        RECT 56.280 20.080 67.190 20.330 ;
        RECT 67.540 20.100 67.890 20.820 ;
        RECT 56.280 20.050 56.620 20.080 ;
        RECT 57.020 20.070 57.360 20.080 ;
        RECT 57.730 20.070 58.080 20.080 ;
        RECT 52.960 19.590 55.910 19.920 ;
        RECT 52.360 19.540 52.860 19.550 ;
        RECT 55.560 19.540 55.910 19.590 ;
        RECT 57.730 19.920 58.350 20.070 ;
        RECT 59.140 19.920 59.450 20.070 ;
        RECT 60.230 19.920 60.540 20.070 ;
        RECT 57.730 19.590 60.680 19.920 ;
        RECT 57.730 19.540 58.080 19.590 ;
        RECT 61.540 19.540 61.910 20.080 ;
        RECT 62.910 19.950 63.220 20.080 ;
        RECT 64.000 19.950 64.310 20.080 ;
        RECT 65.100 19.950 65.720 20.080 ;
        RECT 66.090 20.050 66.430 20.080 ;
        RECT 62.770 19.620 65.720 19.950 ;
        RECT 65.370 19.540 65.720 19.620 ;
        RECT 67.540 19.950 68.160 20.100 ;
        RECT 68.950 19.950 69.260 20.100 ;
        RECT 70.040 19.950 70.350 20.100 ;
        RECT 67.540 19.620 70.490 19.950 ;
        RECT 67.540 19.540 67.890 19.620 ;
        RECT 71.350 19.540 71.670 21.670 ;
        RECT 74.260 21.650 77.410 21.790 ;
        RECT 73.580 21.270 73.890 21.420 ;
        RECT 74.690 21.270 75.000 21.430 ;
        RECT 75.780 21.270 76.090 21.450 ;
        RECT 73.280 20.970 76.220 21.270 ;
        RECT 73.280 20.930 74.030 20.970 ;
        RECT 73.280 20.800 73.660 20.930 ;
        RECT 73.280 20.080 73.630 20.800 ;
        RECT 73.280 19.930 73.900 20.080 ;
        RECT 74.690 19.930 75.000 20.080 ;
        RECT 75.780 19.930 76.090 20.080 ;
        RECT 73.280 19.600 76.230 19.930 ;
        RECT 73.280 19.540 73.630 19.600 ;
        RECT 77.090 19.540 77.410 21.650 ;
        RECT 98.290 19.540 98.850 19.560 ;
        RECT 52.360 19.190 98.850 19.540 ;
        RECT 51.780 19.080 98.850 19.190 ;
        RECT 51.780 19.010 55.050 19.080 ;
        RECT 22.860 18.630 23.180 18.880 ;
        RECT 25.760 18.860 26.040 18.880 ;
        RECT 51.780 18.860 54.940 19.010 ;
        RECT 20.020 18.480 23.180 18.630 ;
        RECT 19.910 18.300 23.180 18.480 ;
        RECT 19.910 18.150 20.220 18.300 ;
        RECT 21.010 18.150 21.320 18.300 ;
        RECT 22.110 18.150 22.420 18.300 ;
        RECT 19.050 17.570 22.000 17.900 ;
        RECT 18.340 17.530 18.690 17.560 ;
        RECT 19.050 17.530 19.670 17.570 ;
        RECT 20.460 17.530 20.770 17.570 ;
        RECT 21.550 17.530 21.860 17.570 ;
        RECT 22.860 17.530 23.180 18.300 ;
        RECT 51.780 17.820 52.100 18.860 ;
        RECT 52.540 17.820 52.850 17.970 ;
        RECT 53.640 17.820 53.950 17.970 ;
        RECT 54.740 17.820 55.050 17.970 ;
        RECT 51.780 17.640 55.050 17.820 ;
        RECT 24.720 17.550 25.050 17.590 ;
        RECT 24.710 17.530 25.060 17.550 ;
        RECT 18.340 17.270 28.370 17.530 ;
        RECT 51.780 17.500 54.940 17.640 ;
        RECT 55.560 17.300 55.910 19.080 ;
        RECT 18.380 17.240 28.370 17.270 ;
        RECT 19.050 16.700 19.400 17.240 ;
        RECT 22.860 16.900 23.180 17.240 ;
        RECT 24.720 17.220 25.050 17.240 ;
        RECT 19.050 16.570 19.430 16.700 ;
        RECT 19.050 16.530 19.800 16.570 ;
        RECT 22.180 16.560 24.520 16.900 ;
        RECT 19.050 16.230 21.990 16.530 ;
        RECT 22.180 16.320 24.560 16.560 ;
        RECT 22.180 16.300 24.520 16.320 ;
        RECT 19.350 16.080 19.660 16.230 ;
        RECT 20.460 16.070 20.770 16.230 ;
        RECT 21.550 16.050 21.860 16.230 ;
        RECT 22.860 15.850 23.180 16.300 ;
        RECT 23.550 16.230 24.210 16.300 ;
        RECT 23.580 16.220 24.180 16.230 ;
        RECT 20.030 15.710 23.180 15.850 ;
        RECT 19.910 15.520 23.180 15.710 ;
        RECT 19.910 15.510 23.090 15.520 ;
        RECT 19.910 15.380 20.220 15.510 ;
        RECT 21.010 15.370 21.320 15.510 ;
        RECT 22.100 15.370 22.410 15.510 ;
        RECT 28.070 15.160 28.360 17.240 ;
        RECT 53.100 17.150 53.410 17.290 ;
        RECT 54.190 17.150 54.500 17.290 ;
        RECT 55.290 17.150 55.910 17.300 ;
        RECT 52.970 16.830 55.910 17.150 ;
        RECT 57.730 17.300 58.080 19.080 ;
        RECT 58.590 19.040 64.860 19.080 ;
        RECT 58.590 19.010 64.750 19.040 ;
        RECT 58.700 18.890 64.750 19.010 ;
        RECT 58.700 18.860 61.910 18.890 ;
        RECT 61.540 18.630 61.910 18.860 ;
        RECT 65.370 18.630 65.720 19.080 ;
        RECT 67.540 18.630 67.890 19.080 ;
        RECT 68.400 19.040 71.670 19.080 ;
        RECT 68.510 18.890 71.670 19.040 ;
        RECT 71.350 18.630 71.670 18.890 ;
        RECT 73.280 18.630 73.630 19.080 ;
        RECT 74.140 19.020 77.410 19.080 ;
        RECT 98.290 19.060 98.850 19.080 ;
        RECT 74.250 18.870 77.410 19.020 ;
        RECT 77.090 18.630 77.410 18.870 ;
        RECT 60.670 18.170 97.750 18.630 ;
        RECT 60.740 18.070 61.260 18.170 ;
        RECT 58.590 17.820 58.900 17.970 ;
        RECT 59.690 17.820 60.000 17.970 ;
        RECT 60.790 17.820 61.100 17.970 ;
        RECT 61.540 17.850 61.910 18.170 ;
        RECT 62.350 17.850 62.660 18.000 ;
        RECT 63.450 17.850 63.760 18.000 ;
        RECT 64.550 17.850 64.860 18.000 ;
        RECT 61.540 17.820 64.860 17.850 ;
        RECT 58.590 17.720 64.860 17.820 ;
        RECT 65.370 17.720 65.720 18.170 ;
        RECT 67.540 17.720 67.890 18.170 ;
        RECT 68.400 17.850 68.710 18.000 ;
        RECT 69.500 17.850 69.810 18.000 ;
        RECT 70.600 17.850 70.910 18.000 ;
        RECT 71.350 17.850 71.670 18.170 ;
        RECT 68.400 17.720 71.670 17.850 ;
        RECT 73.280 17.720 73.630 18.170 ;
        RECT 74.140 17.830 74.450 17.980 ;
        RECT 75.240 17.830 75.550 17.980 ;
        RECT 76.340 17.830 76.650 17.980 ;
        RECT 77.090 17.830 77.410 18.170 ;
        RECT 97.100 18.110 97.660 18.170 ;
        RECT 74.140 17.720 77.410 17.830 ;
        RECT 58.590 17.640 96.660 17.720 ;
        RECT 58.700 17.530 96.660 17.640 ;
        RECT 58.700 17.500 61.860 17.530 ;
        RECT 57.730 17.150 58.350 17.300 ;
        RECT 59.140 17.150 59.450 17.290 ;
        RECT 60.230 17.150 60.540 17.290 ;
        RECT 61.360 17.230 61.670 17.330 ;
        RECT 61.780 17.230 62.090 17.360 ;
        RECT 61.350 17.200 62.090 17.230 ;
        RECT 62.100 17.260 96.660 17.530 ;
        RECT 62.100 17.200 62.750 17.260 ;
        RECT 57.730 16.830 60.670 17.150 ;
        RECT 52.970 16.820 55.680 16.830 ;
        RECT 57.960 16.820 60.670 16.830 ;
        RECT 61.350 17.130 62.750 17.200 ;
        RECT 62.910 17.180 63.220 17.260 ;
        RECT 64.000 17.180 64.310 17.260 ;
        RECT 65.100 17.180 65.720 17.260 ;
        RECT 61.350 16.410 62.100 17.130 ;
        RECT 62.780 16.860 65.720 17.180 ;
        RECT 67.540 17.180 68.160 17.260 ;
        RECT 68.950 17.180 69.260 17.260 ;
        RECT 70.040 17.180 70.350 17.260 ;
        RECT 71.170 17.230 71.480 17.260 ;
        RECT 67.540 16.860 70.480 17.180 ;
        RECT 71.170 17.030 71.910 17.230 ;
        RECT 71.310 16.890 71.910 17.030 ;
        RECT 62.780 16.850 65.490 16.860 ;
        RECT 67.770 16.850 70.480 16.860 ;
        RECT 61.500 16.380 62.100 16.410 ;
        RECT 70.550 16.780 71.070 16.800 ;
        RECT 71.160 16.780 71.910 16.890 ;
        RECT 73.280 17.160 73.900 17.260 ;
        RECT 74.690 17.160 75.000 17.260 ;
        RECT 75.780 17.160 76.090 17.260 ;
        RECT 76.910 17.210 77.220 17.260 ;
        RECT 95.970 17.240 96.530 17.260 ;
        RECT 73.280 16.840 76.220 17.160 ;
        RECT 76.910 17.010 77.650 17.210 ;
        RECT 77.050 16.870 77.650 17.010 ;
        RECT 73.510 16.830 76.220 16.840 ;
        RECT 76.900 16.780 77.650 16.870 ;
        RECT 95.040 16.780 95.600 16.790 ;
        RECT 70.550 16.320 95.690 16.780 ;
        RECT 70.550 16.270 71.080 16.320 ;
        RECT 70.550 16.220 71.070 16.270 ;
        RECT 44.490 15.160 44.810 15.180 ;
        RECT 100.490 15.160 101.650 15.190 ;
        RECT 27.880 14.040 101.650 15.160 ;
        RECT 44.490 14.020 44.810 14.040 ;
        RECT 55.860 13.960 57.780 14.040 ;
        RECT 65.670 13.930 67.600 14.040 ;
        RECT 100.490 14.010 101.650 14.040 ;
        RECT 104.320 11.860 104.520 11.870 ;
        RECT 104.320 11.710 108.260 11.860 ;
        RECT 7.410 10.710 7.910 10.820 ;
        RECT 76.380 10.740 76.770 10.750 ;
        RECT 76.370 10.710 76.770 10.740 ;
        RECT 7.410 10.430 76.770 10.710 ;
        RECT 7.410 10.350 7.910 10.430 ;
        RECT 76.370 10.410 76.770 10.430 ;
        RECT 76.380 10.400 76.770 10.410 ;
        RECT 104.320 8.800 104.520 11.710 ;
        RECT 108.340 11.680 108.660 12.000 ;
        RECT 105.290 10.110 108.100 10.310 ;
        RECT 104.550 8.810 104.980 8.830 ;
        RECT 104.540 8.800 104.990 8.810 ;
        RECT 89.080 8.420 104.990 8.800 ;
        RECT 89.080 3.120 91.040 8.420 ;
        RECT 103.200 8.350 103.530 8.420 ;
        RECT 103.200 7.980 103.400 8.350 ;
        RECT 104.320 7.980 104.520 8.420 ;
        RECT 104.550 8.400 104.980 8.420 ;
        RECT 105.290 7.990 105.500 10.110 ;
        RECT 108.340 10.070 108.660 10.390 ;
        RECT 107.070 8.650 107.380 8.680 ;
        RECT 107.070 8.400 108.140 8.650 ;
        RECT 108.330 8.460 108.650 8.780 ;
        RECT 105.290 7.980 105.920 7.990 ;
        RECT 93.230 7.600 105.920 7.980 ;
        RECT 93.230 3.140 95.210 7.600 ;
        RECT 103.200 7.190 103.400 7.600 ;
        RECT 104.320 7.190 104.520 7.600 ;
        RECT 105.290 7.190 105.500 7.600 ;
        RECT 106.310 7.190 106.730 7.220 ;
        RECT 97.340 6.810 106.730 7.190 ;
        RECT 89.070 2.470 91.100 3.120 ;
        RECT 93.190 2.490 95.220 3.140 ;
        RECT 97.340 3.110 99.320 6.810 ;
        RECT 103.200 4.020 103.400 6.810 ;
        RECT 104.320 4.020 104.520 6.810 ;
        RECT 105.290 4.020 105.500 6.810 ;
        RECT 106.310 6.780 106.730 6.810 ;
        RECT 107.070 4.020 107.370 8.400 ;
        RECT 108.340 7.050 108.660 7.160 ;
        RECT 108.190 6.840 108.660 7.050 ;
        RECT 108.190 5.550 108.380 6.840 ;
        RECT 108.190 5.230 108.650 5.550 ;
        RECT 107.570 4.020 107.890 4.070 ;
        RECT 108.190 4.020 108.380 5.230 ;
        RECT 102.410 3.820 108.650 4.020 ;
        RECT 102.410 3.140 102.610 3.820 ;
        RECT 103.200 3.140 103.400 3.820 ;
        RECT 97.330 2.460 99.360 3.110 ;
        RECT 101.320 2.490 103.400 3.140 ;
        RECT 103.200 0.000 103.400 2.490 ;
        RECT 104.320 0.140 104.520 3.820 ;
        RECT 105.290 3.140 105.500 3.820 ;
        RECT 107.070 3.700 107.370 3.820 ;
        RECT 107.570 3.750 107.890 3.820 ;
        RECT 107.070 3.610 107.830 3.700 ;
        RECT 108.190 3.610 108.380 3.820 ;
        RECT 109.570 3.610 109.770 4.020 ;
        RECT 107.070 3.410 109.770 3.610 ;
        RECT 107.070 3.140 107.540 3.410 ;
        RECT 105.290 2.840 107.540 3.140 ;
        RECT 105.290 2.490 107.370 2.840 ;
        RECT 105.290 0.640 105.500 2.490 ;
        RECT 107.070 2.060 107.370 2.490 ;
        RECT 108.190 2.350 108.380 3.410 ;
        RECT 107.070 1.900 107.430 2.060 ;
        RECT 105.090 0.320 105.500 0.640 ;
        RECT 107.220 0.620 107.430 1.900 ;
        RECT 104.310 0.000 104.520 0.140 ;
        RECT 105.290 0.000 105.500 0.320 ;
        RECT 106.980 0.260 107.430 0.620 ;
        RECT 108.190 2.030 108.650 2.350 ;
        RECT 108.190 0.640 108.380 2.030 ;
        RECT 108.190 0.320 108.610 0.640 ;
        RECT 108.190 0.290 108.380 0.320 ;
        RECT 107.220 0.000 107.430 0.260 ;
        RECT 108.170 0.000 108.380 0.290 ;
      LAYER via2 ;
        RECT 82.780 57.620 83.100 57.940 ;
        RECT 83.810 57.610 84.130 57.930 ;
    END
  END DIG25
  PIN DIG17
    ANTENNADIFFAREA 2.024600 ;
    PORT
      LAYER met2 ;
        RECT 103.570 53.330 104.030 53.460 ;
        RECT 109.880 53.330 110.940 53.410 ;
        RECT 103.570 53.210 110.940 53.330 ;
        RECT 103.570 53.130 110.150 53.210 ;
        RECT 103.570 53.010 104.030 53.130 ;
        RECT 83.950 43.330 103.690 43.510 ;
        RECT 83.950 43.190 88.440 43.330 ;
        RECT 84.190 43.160 88.440 43.190 ;
        RECT 84.190 43.110 84.510 43.160 ;
        RECT 88.120 43.090 88.440 43.160 ;
        RECT 99.180 43.200 103.690 43.330 ;
        RECT 99.180 43.160 103.430 43.200 ;
        RECT 99.180 43.090 99.500 43.160 ;
        RECT 103.110 43.110 103.430 43.160 ;
        RECT 103.650 9.620 104.080 9.640 ;
        RECT 85.150 9.590 87.110 9.620 ;
        RECT 103.630 9.590 104.090 9.620 ;
        RECT 85.150 9.240 104.090 9.590 ;
        RECT 85.150 3.140 87.110 9.240 ;
        RECT 103.630 9.220 104.090 9.240 ;
        RECT 103.650 9.210 104.080 9.220 ;
        RECT 85.120 2.490 87.150 3.140 ;
    END
  END DIG17
  PIN DIG16
    PORT
      LAYER met2 ;
        RECT 43.780 59.520 44.340 59.690 ;
        RECT 43.780 59.070 43.950 59.520 ;
        RECT 42.810 58.960 43.200 59.050 ;
        RECT 43.680 58.960 43.950 59.070 ;
        RECT 42.810 58.790 43.960 58.960 ;
        RECT 43.680 58.750 43.780 58.790 ;
        RECT 42.790 10.080 43.210 10.090 ;
        RECT 42.790 9.830 83.060 10.080 ;
        RECT 42.790 9.750 83.070 9.830 ;
        RECT 42.790 9.740 43.210 9.750 ;
        RECT 77.030 9.730 83.070 9.750 ;
        RECT 81.130 9.230 83.070 9.730 ;
        RECT 81.130 3.160 83.060 9.230 ;
        RECT 81.040 2.380 83.070 3.160 ;
    END
  END DIG16
  PIN DIG15
    PORT
      LAYER met2 ;
        RECT 43.780 57.690 44.340 57.860 ;
        RECT 42.210 57.420 42.540 57.430 ;
        RECT 42.190 57.320 42.560 57.420 ;
        RECT 43.780 57.320 43.950 57.690 ;
        RECT 42.190 57.150 43.950 57.320 ;
        RECT 42.190 57.040 42.560 57.150 ;
        RECT 43.680 57.140 43.950 57.150 ;
        RECT 43.680 57.000 43.780 57.140 ;
        RECT 42.190 9.460 42.570 9.470 ;
        RECT 42.190 9.130 78.990 9.460 ;
        RECT 42.190 9.120 42.570 9.130 ;
        RECT 72.920 9.120 78.990 9.130 ;
        RECT 77.030 8.800 78.990 9.120 ;
        RECT 77.030 3.140 78.980 8.800 ;
        RECT 76.970 2.490 79.000 3.140 ;
    END
  END DIG15
  PIN DIG14
    PORT
      LAYER met2 ;
        RECT 43.740 55.960 44.340 56.130 ;
        RECT 41.610 55.840 42.000 55.940 ;
        RECT 43.740 55.840 43.910 55.960 ;
        RECT 41.610 55.670 43.910 55.840 ;
        RECT 41.610 55.570 42.000 55.670 ;
        RECT 41.550 8.830 41.970 8.840 ;
        RECT 41.550 8.500 74.910 8.830 ;
        RECT 41.550 8.490 41.970 8.500 ;
        RECT 72.920 3.140 74.910 8.500 ;
        RECT 72.920 2.490 74.950 3.140 ;
    END
  END DIG14
  PIN DIG13
    PORT
      LAYER met2 ;
        RECT 40.970 54.240 41.360 54.330 ;
        RECT 43.910 54.240 44.340 54.410 ;
        RECT 40.970 54.070 44.540 54.240 ;
        RECT 40.970 53.980 41.360 54.070 ;
        RECT 43.910 54.050 44.080 54.070 ;
        RECT 40.960 8.190 41.360 8.210 ;
        RECT 40.960 7.860 70.900 8.190 ;
        RECT 40.960 7.850 41.360 7.860 ;
        RECT 68.940 3.140 70.890 7.860 ;
        RECT 68.890 2.490 70.920 3.140 ;
    END
  END DIG13
  PIN DIG12
    PORT
      LAYER met2 ;
        RECT 40.330 53.670 40.720 53.780 ;
        RECT 40.330 53.500 44.540 53.670 ;
        RECT 40.330 53.400 40.720 53.500 ;
        RECT 40.300 7.520 40.710 7.530 ;
        RECT 40.290 7.190 66.810 7.520 ;
        RECT 40.300 7.170 40.710 7.190 ;
        RECT 64.900 3.120 66.810 7.190 ;
        RECT 64.820 2.470 66.850 3.120 ;
    END
  END DIG12
  PIN DIG11
    PORT
      LAYER met2 ;
        RECT 39.720 52.100 40.110 52.200 ;
        RECT 39.720 51.930 44.540 52.100 ;
        RECT 39.720 51.830 40.110 51.930 ;
        RECT 43.990 51.770 44.340 51.930 ;
        RECT 39.720 6.900 40.130 6.910 ;
        RECT 39.720 6.880 62.790 6.900 ;
        RECT 39.720 6.570 62.800 6.880 ;
        RECT 39.720 6.560 40.130 6.570 ;
        RECT 60.800 3.190 62.800 6.570 ;
        RECT 60.770 2.490 62.800 3.190 ;
    END
  END DIG11
  PIN DIG10
    PORT
      LAYER met2 ;
        RECT 39.090 50.570 39.510 50.660 ;
        RECT 39.090 50.400 43.990 50.570 ;
        RECT 39.090 50.310 39.510 50.400 ;
        RECT 43.820 50.220 43.990 50.400 ;
        RECT 43.820 50.050 44.340 50.220 ;
        RECT 39.120 6.250 39.510 6.260 ;
        RECT 39.120 5.930 58.810 6.250 ;
        RECT 39.220 5.920 58.810 5.930 ;
        RECT 56.820 3.210 58.810 5.920 ;
        RECT 56.810 2.460 58.840 3.210 ;
    END
  END DIG10
  PIN DIG09
    PORT
      LAYER met2 ;
        RECT 38.530 49.000 38.920 49.090 ;
        RECT 43.680 49.000 43.780 49.160 ;
        RECT 38.530 48.830 43.900 49.000 ;
        RECT 38.530 48.740 38.920 48.830 ;
        RECT 43.740 48.720 43.900 48.830 ;
        RECT 43.740 48.420 43.910 48.720 ;
        RECT 43.740 48.250 44.340 48.420 ;
        RECT 38.540 5.640 38.930 5.690 ;
        RECT 38.540 5.360 54.900 5.640 ;
        RECT 38.800 5.310 54.900 5.360 ;
        RECT 52.830 2.490 54.860 5.310 ;
    END
  END DIG09
  PIN DIG08
    PORT
      LAYER met2 ;
        RECT 37.920 43.530 38.290 43.650 ;
        RECT 37.920 43.360 44.240 43.530 ;
        RECT 37.920 43.250 38.290 43.360 ;
        RECT 37.960 4.670 50.700 5.000 ;
        RECT 48.650 3.370 50.680 4.670 ;
        RECT 48.650 3.080 50.690 3.370 ;
        RECT 48.660 2.470 50.690 3.080 ;
    END
  END DIG08
  PIN DIG07
    PORT
      LAYER met2 ;
        RECT 37.280 41.940 37.670 42.030 ;
        RECT 37.280 41.820 44.240 41.940 ;
        RECT 37.280 41.770 44.340 41.820 ;
        RECT 37.280 41.680 37.670 41.770 ;
        RECT 43.950 41.650 44.340 41.770 ;
        RECT 44.570 4.370 46.590 4.390 ;
        RECT 37.410 4.360 46.620 4.370 ;
        RECT 37.310 4.040 46.620 4.360 ;
        RECT 37.310 4.030 37.700 4.040 ;
        RECT 44.540 2.490 46.620 4.040 ;
    END
  END DIG07
  PIN DIG06
    PORT
      LAYER met2 ;
        RECT 36.660 40.390 37.050 40.470 ;
        RECT 36.660 40.220 43.840 40.390 ;
        RECT 36.660 40.140 37.050 40.220 ;
        RECT 43.690 40.150 43.840 40.220 ;
        RECT 43.690 40.040 43.860 40.150 ;
        RECT 43.690 39.870 44.340 40.040 ;
        RECT 36.670 3.380 42.650 3.720 ;
        RECT 40.620 3.120 42.660 3.380 ;
        RECT 40.610 2.460 42.660 3.120 ;
    END
  END DIG06
  PIN DIG05
    PORT
      LAYER met2 ;
        RECT 36.050 38.910 36.470 39.000 ;
        RECT 43.680 38.910 43.780 39.030 ;
        RECT 36.050 38.740 43.860 38.910 ;
        RECT 36.050 38.640 36.470 38.740 ;
        RECT 43.680 38.710 43.860 38.740 ;
        RECT 43.690 38.250 43.860 38.710 ;
        RECT 43.690 38.080 44.340 38.250 ;
        RECT 36.060 3.130 36.610 3.150 ;
        RECT 36.060 2.700 38.610 3.130 ;
        RECT 36.580 2.470 38.610 2.700 ;
    END
  END DIG05
  PIN DIG04
    PORT
      LAYER met2 ;
        RECT 43.880 34.280 44.300 34.450 ;
        RECT 43.880 34.180 44.260 34.280 ;
        RECT 43.880 33.960 44.160 34.180 ;
        RECT 35.410 33.740 35.820 33.840 ;
        RECT 43.880 33.740 44.150 33.960 ;
        RECT 35.410 33.570 44.150 33.740 ;
        RECT 35.410 33.480 35.820 33.570 ;
        RECT 43.880 33.560 44.050 33.570 ;
        RECT 34.560 3.150 35.210 3.160 ;
        RECT 32.530 2.520 35.210 3.150 ;
        RECT 32.530 2.490 34.560 2.520 ;
    END
  END DIG04
  PIN DIG03
    PORT
      LAYER met2 ;
        RECT 43.820 32.520 44.300 32.690 ;
        RECT 34.750 32.170 35.140 32.280 ;
        RECT 43.820 32.230 43.990 32.520 ;
        RECT 43.820 32.170 43.980 32.230 ;
        RECT 34.750 32.010 43.980 32.170 ;
        RECT 34.750 32.000 43.630 32.010 ;
        RECT 34.750 31.900 35.140 32.000 ;
        RECT 34.730 3.780 35.220 3.980 ;
        RECT 29.120 3.760 35.220 3.780 ;
        RECT 28.550 3.480 35.220 3.760 ;
        RECT 28.550 3.380 35.130 3.480 ;
        RECT 28.550 3.150 30.530 3.380 ;
        RECT 28.530 2.490 30.560 3.150 ;
    END
  END DIG03
  PIN DIG02
    PORT
      LAYER met2 ;
        RECT 43.740 30.710 44.300 30.880 ;
        RECT 43.740 30.670 43.910 30.710 ;
        RECT 34.140 30.630 34.510 30.640 ;
        RECT 43.740 30.630 43.900 30.670 ;
        RECT 34.140 30.460 43.900 30.630 ;
        RECT 34.140 30.250 34.510 30.460 ;
        RECT 34.050 4.590 34.590 4.660 ;
        RECT 24.620 4.160 34.590 4.590 ;
        RECT 24.620 3.150 26.600 4.160 ;
        RECT 24.570 2.490 26.600 3.150 ;
    END
  END DIG02
  PIN DIG01
    PORT
      LAYER met2 ;
        RECT 33.450 29.090 33.840 29.190 ;
        RECT 43.650 29.090 44.300 29.160 ;
        RECT 33.450 28.990 44.300 29.090 ;
        RECT 33.450 28.920 43.940 28.990 ;
        RECT 33.450 28.820 33.840 28.920 ;
        RECT 43.770 28.900 43.940 28.920 ;
        RECT 33.400 5.430 33.940 5.470 ;
        RECT 20.570 5.390 33.940 5.430 ;
        RECT 20.520 5.000 33.940 5.390 ;
        RECT 20.520 3.120 22.530 5.000 ;
        RECT 33.400 4.970 33.940 5.000 ;
        RECT 20.500 2.460 22.530 3.120 ;
    END
  END DIG01
  PIN OUTPUTTA1    
    ANTENNAGATEAREA 0.335600 ;
    ANTENNADIFFAREA 3.191500 ;
    PORT
      LAYER nwell ;
        RECT 0.550 65.890 3.290 69.390 ;
      LAYER met2 ;
        RECT 6.250 68.580 6.930 69.460 ;
        RECT 0.960 68.020 1.280 68.280 ;
        RECT 1.640 68.010 1.950 68.340 ;
        RECT 2.370 68.030 2.690 68.290 ;
        RECT 6.250 68.260 9.610 68.580 ;
        RECT 6.250 68.110 6.930 68.260 ;
        RECT 3.120 67.980 17.770 68.110 ;
        RECT 0.450 67.900 17.770 67.980 ;
        RECT 0.450 67.730 3.260 67.900 ;
        RECT 0.450 67.220 3.120 67.730 ;
        RECT 3.520 67.690 3.840 67.900 ;
        RECT 0.960 67.150 1.280 67.220 ;
        RECT 1.640 67.170 1.950 67.220 ;
        RECT 2.390 67.170 2.710 67.220 ;
        RECT 6.250 67.140 6.930 67.900 ;
        RECT 8.940 67.870 9.520 67.900 ;
        RECT 8.940 67.840 9.260 67.870 ;
        RECT 17.190 67.600 17.430 67.900 ;
        RECT 17.030 67.270 17.430 67.600 ;
        RECT 17.190 67.230 17.430 67.270 ;
        RECT 118.350 65.560 119.120 65.710 ;
        RECT 8.860 65.140 119.120 65.560 ;
        RECT 92.050 65.100 92.360 65.140 ;
        RECT 118.350 65.000 119.120 65.140 ;
        RECT 118.160 45.800 118.940 45.950 ;
        RECT 120.900 45.800 121.800 46.720 ;
        RECT 118.160 45.330 121.800 45.800 ;
        RECT 118.160 45.180 118.940 45.330 ;
        RECT 120.900 44.630 121.800 45.330 ;
    END
  END OUTPUTTA1    
  PIN DRAINOUT
    PORT
      LAYER met1 ;
        RECT 121.030 60.210 121.310 62.960 ;
        RECT 121.030 59.890 121.480 60.210 ;
        RECT 121.030 58.670 121.310 59.890 ;
        RECT 120.760 58.530 121.310 58.670 ;
        RECT 121.030 56.910 121.310 58.530 ;
      LAYER via ;
        RECT 121.220 59.920 121.480 60.180 ;
    END
  END DRAINOUT
  PIN ROWTERM2
    PORT
      LAYER met2 ;
        RECT 100.860 64.560 101.180 64.680 ;
        RECT 120.940 64.560 121.800 65.330 ;
        RECT 123.130 64.560 123.450 64.680 ;
        RECT 100.860 64.380 123.450 64.560 ;
        RECT 91.710 64.030 92.130 64.050 ;
        RECT 100.660 64.030 100.740 64.200 ;
        RECT 120.940 64.030 121.800 64.380 ;
        RECT 91.710 63.660 121.800 64.030 ;
        RECT 91.710 63.640 92.130 63.660 ;
        RECT 120.940 63.610 121.800 63.660 ;
        RECT 125.120 63.610 125.280 63.630 ;
        RECT 116.060 63.560 125.280 63.610 ;
        RECT 116.060 63.460 125.160 63.560 ;
        RECT 120.940 63.230 121.800 63.460 ;
        RECT 74.960 60.440 75.240 60.460 ;
        RECT 74.940 60.410 75.260 60.440 ;
        RECT 91.650 60.410 102.200 60.460 ;
        RECT 107.080 60.410 108.420 60.950 ;
        RECT 74.940 60.200 108.420 60.410 ;
        RECT 74.940 60.180 75.260 60.200 ;
        RECT 74.960 60.160 75.240 60.180 ;
        RECT 91.760 59.860 92.020 60.100 ;
        RECT 91.650 59.750 92.020 59.860 ;
        RECT 91.650 59.600 91.970 59.750 ;
        RECT 107.080 59.670 108.420 60.200 ;
        RECT 91.650 41.810 92.090 41.930 ;
        RECT 91.520 41.630 92.090 41.810 ;
        RECT 91.640 41.530 92.090 41.630 ;
        RECT 83.750 41.470 83.810 41.510 ;
        RECT 91.640 41.470 92.040 41.530 ;
        RECT 80.810 41.290 92.040 41.470 ;
    END
  END ROWTERM2
  PIN COLUMN2
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 90.930 68.740 91.370 68.760 ;
        RECT 120.970 68.740 121.830 69.420 ;
        RECT 90.930 68.490 121.830 68.740 ;
        RECT 90.930 68.370 125.180 68.490 ;
        RECT 90.930 68.350 91.370 68.370 ;
        RECT 92.830 68.310 101.940 68.370 ;
        RECT 116.060 68.310 125.180 68.370 ;
        RECT 120.970 67.320 121.830 68.310 ;
        RECT 80.250 44.240 80.560 44.410 ;
        RECT 78.230 44.180 80.560 44.240 ;
        RECT 80.700 44.180 80.790 44.240 ;
        RECT 83.570 44.180 91.340 44.260 ;
        RECT 78.230 44.060 91.340 44.180 ;
        RECT 79.650 43.920 91.340 44.060 ;
        RECT 79.650 43.910 79.970 43.920 ;
        RECT 90.910 43.850 91.340 43.920 ;
    END
  END COLUMN2
  PIN COLUMN1
    ANTENNADIFFAREA 0.176000 ;
    PORT
      LAYER met2 ;
        RECT 90.100 72.200 90.560 72.220 ;
        RECT 120.970 72.200 121.830 73.550 ;
        RECT 90.100 71.830 121.830 72.200 ;
        RECT 90.100 71.810 90.560 71.830 ;
        RECT 120.970 71.450 121.830 71.830 ;
        RECT 78.230 44.980 80.410 45.120 ;
        RECT 78.230 44.940 80.560 44.980 ;
        RECT 62.310 44.780 62.630 44.790 ;
        RECT 80.250 44.780 80.560 44.940 ;
        RECT 90.120 44.780 90.580 44.850 ;
        RECT 62.310 44.500 90.580 44.780 ;
        RECT 62.310 44.450 62.630 44.500 ;
        RECT 78.230 44.490 80.410 44.500 ;
        RECT 90.120 44.440 90.580 44.500 ;
    END
  END COLUMN1
  PIN GATE2
    PORT
      LAYER met1 ;
        RECT 106.030 73.180 109.220 74.300 ;
        RECT 107.120 60.980 108.400 73.180 ;
        RECT 107.110 59.640 108.400 60.980 ;
        RECT 107.120 59.150 108.400 59.640 ;
      LAYER via ;
        RECT 107.110 59.670 108.390 60.950 ;
    END
  END GATE2
  PIN DRAININJECT
    PORT
      LAYER met2 ;
        RECT 50.480 70.310 50.930 70.330 ;
        RECT 50.470 70.250 50.950 70.310 ;
        RECT 28.080 69.950 50.950 70.250 ;
        RECT 50.470 69.890 50.950 69.950 ;
        RECT 50.480 69.870 50.930 69.890 ;
    END
  END DRAININJECT
  PIN VTUN
    PORT
      LAYER met2 ;
        RECT 46.630 69.550 47.080 69.570 ;
        RECT 46.620 69.540 47.100 69.550 ;
        RECT 70.240 69.540 71.660 69.580 ;
        RECT 46.620 69.140 71.710 69.540 ;
        RECT 46.620 69.130 47.100 69.140 ;
        RECT 46.630 69.110 47.080 69.130 ;
        RECT 70.240 69.100 71.660 69.140 ;
    END
  END VTUN
  PIN LARGECAPACITOR
    ANTENNADIFFAREA 4.612400 ;
    PORT
      LAYER met2 ;
        RECT 0.450 64.010 4.330 64.340 ;
        RECT 5.800 64.320 6.480 64.990 ;
        RECT 14.720 64.320 15.190 64.340 ;
        RECT 0.450 63.920 4.340 64.010 ;
        RECT 0.450 63.850 4.330 63.920 ;
        RECT 0.830 63.790 1.140 63.850 ;
        RECT 1.760 63.790 2.070 63.850 ;
        RECT 2.460 63.790 2.770 63.850 ;
        RECT 3.200 63.790 3.510 63.850 ;
        RECT 3.650 63.780 4.220 63.850 ;
        RECT 3.650 63.670 4.090 63.780 ;
        RECT 5.800 63.740 15.190 64.320 ;
        RECT 5.800 63.670 6.520 63.740 ;
        RECT 14.720 63.720 15.190 63.740 ;
        RECT 16.310 63.670 16.620 63.940 ;
        RECT 26.170 63.670 26.480 63.960 ;
        RECT 3.360 63.460 26.590 63.670 ;
        RECT 5.800 62.670 6.480 63.460 ;
    END
  END LARGECAPACITOR
  PIN DRAIN6N
    PORT
      LAYER met2 ;
        RECT 17.090 19.910 17.460 19.920 ;
        RECT 6.200 19.090 7.470 19.790 ;
        RECT 15.770 19.530 18.380 19.910 ;
        RECT 15.770 19.090 16.150 19.530 ;
        RECT 17.090 19.510 17.460 19.530 ;
        RECT 6.200 18.710 16.150 19.090 ;
        RECT 6.200 17.910 7.470 18.710 ;
    END
  END DRAIN6N
  PIN DRAIN6P
    PORT
      LAYER met2 ;
        RECT 6.200 13.860 7.470 14.770 ;
        RECT 6.200 13.480 16.170 13.860 ;
        RECT 6.200 12.890 7.470 13.480 ;
        RECT 15.790 12.630 16.170 13.480 ;
        RECT 17.090 12.630 17.460 12.640 ;
        RECT 15.790 12.250 18.510 12.630 ;
        RECT 17.090 12.230 17.460 12.250 ;
    END
  END DRAIN6P
  PIN DRAIN5P
    PORT
      LAYER met2 ;
        RECT 15.360 29.540 15.770 29.560 ;
        RECT 17.130 29.540 19.120 29.560 ;
        RECT 15.360 29.500 19.120 29.540 ;
        RECT 15.360 29.280 20.450 29.500 ;
        RECT 15.360 29.170 17.510 29.280 ;
        RECT 15.360 29.150 15.770 29.170 ;
        RECT 17.130 29.150 17.500 29.170 ;
        RECT 6.140 23.300 7.410 24.080 ;
        RECT 15.370 23.300 15.780 23.320 ;
        RECT 6.140 22.930 15.780 23.300 ;
        RECT 6.140 22.200 7.410 22.930 ;
        RECT 15.370 22.910 15.780 22.930 ;
    END
  END DRAIN5P
  PIN DARIN4P
    PORT
      LAYER met2 ;
        RECT 6.200 32.550 7.470 33.320 ;
        RECT 6.200 32.180 12.190 32.550 ;
        RECT 6.200 31.440 7.470 32.180 ;
        RECT 11.820 30.520 12.190 32.180 ;
        RECT 11.820 30.340 17.770 30.520 ;
        RECT 11.820 30.270 17.840 30.340 ;
        RECT 19.230 30.270 20.450 30.280 ;
        RECT 11.820 30.150 20.450 30.270 ;
        RECT 17.130 30.110 20.450 30.150 ;
        RECT 17.490 30.060 20.450 30.110 ;
    END
  END DARIN4P
  PIN DRAIN5N
    PORT
      LAYER met2 ;
        RECT 10.130 34.200 10.900 34.390 ;
        RECT 17.130 34.200 17.520 34.220 ;
        RECT 10.130 34.160 17.520 34.200 ;
        RECT 10.130 33.950 20.440 34.160 ;
        RECT 10.130 33.830 17.510 33.950 ;
        RECT 10.130 33.650 10.900 33.830 ;
        RECT 17.130 33.810 17.500 33.830 ;
        RECT 6.200 28.410 7.470 29.230 ;
        RECT 10.130 28.410 10.930 28.550 ;
        RECT 6.200 27.910 10.930 28.410 ;
        RECT 6.200 27.350 7.470 27.910 ;
        RECT 10.130 27.780 10.930 27.910 ;
    END
  END DRAIN5N
  PIN DRAIN4N
    PORT
      LAYER met2 ;
        RECT 6.140 36.580 7.410 37.420 ;
        RECT 6.140 36.210 15.840 36.580 ;
        RECT 6.140 35.540 7.410 36.210 ;
        RECT 15.470 34.860 15.840 36.210 ;
        RECT 15.470 34.850 17.500 34.860 ;
        RECT 15.470 34.670 17.720 34.850 ;
        RECT 15.470 34.610 19.120 34.670 ;
        RECT 15.470 34.490 20.450 34.610 ;
        RECT 17.130 34.450 20.450 34.490 ;
        RECT 17.500 34.390 20.450 34.450 ;
    END
  END DRAIN4N
  PIN DRAIN3P
    PORT
      LAYER met2 ;
        RECT 17.130 52.100 22.780 52.290 ;
        RECT 6.200 40.730 7.470 41.640 ;
        RECT 17.130 40.730 17.500 52.100 ;
        RECT 6.200 40.360 17.500 40.730 ;
        RECT 6.200 39.760 7.470 40.360 ;
    END
  END DRAIN3P
  PIN DRAIN2P
    PORT
      LAYER met2 ;
        RECT 20.680 54.310 20.820 54.330 ;
        RECT 20.680 54.210 20.750 54.310 ;
        RECT 21.960 54.210 22.330 54.350 ;
        RECT 16.290 54.190 22.780 54.210 ;
        RECT 16.000 54.020 22.780 54.190 ;
        RECT 16.000 53.840 17.500 54.020 ;
        RECT 16.000 53.250 16.660 53.840 ;
        RECT 17.130 53.800 17.500 53.840 ;
        RECT 20.680 53.350 20.820 53.370 ;
        RECT 20.680 53.250 20.830 53.350 ;
        RECT 16.000 53.060 22.780 53.250 ;
        RECT 16.000 52.880 17.500 53.060 ;
        RECT 16.000 52.870 16.670 52.880 ;
        RECT 16.000 52.830 16.660 52.870 ;
        RECT 17.130 52.840 17.500 52.880 ;
        RECT 6.140 45.570 7.410 46.460 ;
        RECT 16.000 45.570 16.370 52.830 ;
        RECT 6.140 45.200 16.370 45.570 ;
        RECT 6.140 44.580 7.410 45.200 ;
    END
  END DRAIN2P
  PIN DRAIN3N
    ANTENNADIFFAREA 0.130200 ;
    PORT
      LAYER met2 ;
        RECT 17.130 57.280 17.500 57.290 ;
        RECT 15.340 57.050 17.500 57.280 ;
        RECT 20.680 57.050 20.850 57.220 ;
        RECT 21.860 57.050 22.460 57.080 ;
        RECT 22.530 57.050 22.840 57.320 ;
        RECT 15.340 56.990 22.840 57.050 ;
        RECT 15.340 56.920 22.760 56.990 ;
        RECT 15.340 56.220 15.960 56.920 ;
        RECT 17.130 56.880 22.760 56.920 ;
        RECT 17.130 56.220 17.500 56.260 ;
        RECT 14.810 56.130 17.500 56.220 ;
        RECT 20.680 56.130 20.840 56.300 ;
        RECT 14.810 55.960 22.760 56.130 ;
        RECT 14.810 55.850 17.500 55.960 ;
        RECT 14.810 55.740 15.960 55.850 ;
        RECT 14.810 55.290 15.920 55.740 ;
        RECT 17.130 55.290 17.500 55.330 ;
        RECT 14.810 55.210 17.500 55.290 ;
        RECT 20.680 55.210 20.820 55.290 ;
        RECT 21.960 55.210 22.330 55.340 ;
        RECT 14.810 55.040 22.760 55.210 ;
        RECT 14.810 54.920 17.500 55.040 ;
        RECT 14.810 54.880 15.710 54.920 ;
        RECT 6.200 50.330 7.470 51.210 ;
        RECT 14.810 50.330 15.180 54.880 ;
        RECT 6.200 49.960 15.180 50.330 ;
        RECT 6.200 49.330 7.470 49.960 ;
    END
  END DRAIN3N
  PIN SOURCEP
    ANTENNADIFFAREA 0.819000 ;
    PORT
      LAYER met2 ;
        RECT 5.480 59.170 6.750 60.630 ;
        RECT 16.830 59.170 17.130 59.180 ;
        RECT 22.520 59.170 22.830 59.300 ;
        RECT 23.610 59.170 23.920 59.310 ;
        RECT 26.420 59.170 26.710 59.190 ;
        RECT 5.480 58.780 26.740 59.170 ;
        RECT 5.480 58.750 6.750 58.780 ;
        RECT 26.420 58.760 26.710 58.780 ;
        RECT 26.400 54.150 26.720 54.180 ;
        RECT 25.190 53.950 26.820 54.150 ;
        RECT 26.400 53.920 26.720 53.950 ;
        RECT 26.410 53.190 26.730 53.220 ;
        RECT 25.190 52.990 26.820 53.190 ;
        RECT 26.410 52.960 26.730 52.990 ;
        RECT 26.400 52.230 26.720 52.260 ;
        RECT 25.190 52.030 26.820 52.230 ;
        RECT 26.400 52.000 26.720 52.030 ;
        RECT 26.560 32.870 28.430 32.950 ;
        RECT 26.410 32.730 28.430 32.870 ;
        RECT 26.410 32.540 26.720 32.730 ;
        RECT 26.410 30.270 26.700 30.290 ;
        RECT 26.400 30.240 26.720 30.270 ;
        RECT 23.550 30.030 26.720 30.240 ;
        RECT 23.550 29.210 23.760 30.030 ;
        RECT 24.900 29.860 25.150 30.030 ;
        RECT 26.400 30.010 26.720 30.030 ;
        RECT 26.410 29.990 26.700 30.010 ;
        RECT 26.600 28.980 28.430 29.060 ;
        RECT 26.430 28.850 28.430 28.980 ;
        RECT 26.430 28.650 26.740 28.850 ;
        RECT 26.340 11.660 26.650 11.680 ;
        RECT 22.110 11.320 26.650 11.660 ;
        RECT 26.340 11.300 26.650 11.320 ;
    END
  END SOURCEP
  PIN GATE1
    PORT
      LAYER met2 ;
        RECT 62.540 61.020 62.860 61.060 ;
        RECT 78.190 61.020 79.470 61.120 ;
        RECT 62.540 60.810 79.470 61.020 ;
        RECT 62.540 60.780 62.860 60.810 ;
    END
  END GATE1
  PIN VINJ
    PORT
      LAYER met2 ;
        RECT 6.100 70.570 8.580 70.580 ;
        RECT 6.100 70.180 10.050 70.570 ;
        RECT 8.370 69.810 10.050 70.180 ;
    END
    PORT
      LAYER met2 ;
        RECT 5.800 62.170 6.310 62.290 ;
        RECT 5.800 61.880 8.900 62.170 ;
        RECT 6.310 61.870 8.900 61.880 ;
    END
    PORT
      LAYER met2 ;
        RECT 52.140 67.930 52.640 67.960 ;
        RECT 57.860 67.930 58.360 67.960 ;
        RECT 52.140 67.520 82.300 67.930 ;
        RECT 52.290 67.490 82.300 67.520 ;
    END
  END VINJ
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 8.250 66.770 9.780 66.930 ;
        RECT 6.440 66.440 9.780 66.770 ;
        RECT 6.440 66.370 8.710 66.440 ;
        RECT 6.440 66.170 6.840 66.370 ;
        RECT 6.090 65.770 6.840 66.170 ;
    END
    PORT
      LAYER met2 ;
        RECT 47.720 66.920 48.220 66.940 ;
        RECT 53.460 66.920 53.900 66.970 ;
        RECT 67.830 66.920 68.330 66.940 ;
        RECT 47.720 66.500 74.230 66.920 ;
        RECT 47.870 66.480 74.230 66.500 ;
        RECT 53.460 66.470 53.900 66.480 ;
        RECT 73.630 66.460 74.130 66.480 ;
        RECT 88.080 57.170 88.390 57.310 ;
        RECT 85.910 56.990 88.390 57.170 ;
        RECT 88.080 56.980 88.390 56.990 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 121.900 59.640 122.220 59.720 ;
        RECT 121.900 59.400 122.470 59.640 ;
        RECT 122.130 59.070 122.470 59.400 ;
        RECT 121.850 58.750 122.470 59.070 ;
        RECT 122.130 57.800 122.470 58.750 ;
        RECT 121.850 57.480 122.470 57.800 ;
        RECT 122.130 57.150 122.470 57.480 ;
        RECT 121.900 56.830 122.470 57.150 ;
        RECT 122.130 56.720 122.470 56.830 ;
        RECT 121.900 56.400 122.470 56.720 ;
        RECT 122.130 56.070 122.470 56.400 ;
        RECT 121.850 55.750 122.470 56.070 ;
        RECT 122.130 54.800 122.470 55.750 ;
        RECT 121.850 54.480 122.470 54.800 ;
        RECT 122.130 54.150 122.470 54.480 ;
        RECT 121.900 53.920 122.470 54.150 ;
        RECT 121.900 53.830 122.220 53.920 ;
      LAYER via ;
        RECT 121.930 59.430 122.190 59.690 ;
        RECT 121.880 58.780 122.140 59.040 ;
        RECT 121.880 57.510 122.140 57.770 ;
        RECT 121.930 56.860 122.190 57.120 ;
        RECT 121.930 56.430 122.190 56.690 ;
        RECT 121.880 55.780 122.140 56.040 ;
        RECT 121.880 54.510 122.140 54.770 ;
        RECT 121.930 53.860 122.190 54.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.320 20.360 56.580 20.820 ;
        RECT 57.060 20.380 57.320 20.820 ;
        RECT 56.310 20.020 56.590 20.360 ;
        RECT 57.050 20.040 57.330 20.380 ;
        RECT 56.320 18.610 56.580 20.020 ;
        RECT 57.060 18.610 57.320 20.040 ;
        RECT 56.320 15.180 57.320 18.610 ;
        RECT 55.840 15.140 57.770 15.180 ;
        RECT 55.300 13.950 57.770 15.140 ;
        RECT 55.300 2.460 56.240 13.950 ;
      LAYER via ;
        RECT 56.310 20.050 56.590 20.330 ;
        RECT 57.050 20.070 57.330 20.350 ;
        RECT 56.630 15.100 57.750 15.120 ;
        RECT 55.890 14.000 57.750 15.100 ;
        RECT 55.890 13.980 57.010 14.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 66.130 20.360 66.390 20.850 ;
        RECT 66.120 20.020 66.400 20.360 ;
        RECT 66.130 18.840 66.390 20.020 ;
        RECT 66.870 18.840 67.130 20.850 ;
        RECT 66.130 15.240 67.130 18.840 ;
        RECT 66.130 15.200 68.150 15.240 ;
        RECT 65.650 13.920 68.150 15.200 ;
        RECT 67.260 3.920 68.150 13.920 ;
        RECT 67.260 3.190 68.180 3.920 ;
        RECT 67.230 2.460 68.150 3.190 ;
      LAYER via ;
        RECT 66.120 20.050 66.400 20.330 ;
        RECT 65.700 13.950 67.560 15.140 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 0.600 72.960 10.290 77.560 ;
        RECT 12.940 73.180 15.650 73.220 ;
        RECT 0.000 71.570 10.290 72.960 ;
        RECT 12.930 71.530 15.650 73.180 ;
        RECT 18.130 71.480 20.350 73.170 ;
        RECT 130.580 72.650 132.310 72.990 ;
        RECT 130.560 71.090 132.310 72.650 ;
        RECT 12.940 70.190 15.650 70.230 ;
        RECT 12.930 69.920 15.650 70.190 ;
        RECT 12.220 68.280 16.220 69.920 ;
        RECT 130.560 69.460 132.290 71.090 ;
        RECT 129.040 69.070 132.350 69.460 ;
        RECT 105.510 69.030 108.220 69.070 ;
        RECT 129.040 69.030 132.590 69.070 ;
        RECT 12.930 67.530 15.650 68.280 ;
        RECT 17.430 67.770 19.040 68.560 ;
        RECT 19.540 67.770 20.050 67.940 ;
        RECT 20.090 67.770 21.240 67.940 ;
        RECT 12.220 63.930 16.220 67.120 ;
        RECT 17.430 66.590 21.430 67.770 ;
        RECT 105.510 67.380 108.230 69.030 ;
        RECT 124.280 68.980 127.590 68.990 ;
        RECT 126.630 68.950 126.820 68.980 ;
        RECT 129.040 67.380 132.600 69.030 ;
        RECT 17.430 66.580 18.220 66.590 ;
        RECT 19.540 66.580 21.430 66.590 ;
        RECT 18.220 66.390 18.490 66.570 ;
        RECT 19.540 66.380 20.050 66.580 ;
        RECT 20.090 66.390 21.240 66.580 ;
        RECT 25.150 65.070 25.370 65.180 ;
        RECT 100.800 64.700 101.360 66.760 ;
        RECT 100.660 64.690 103.970 64.700 ;
        RECT 100.800 64.340 101.360 64.690 ;
        RECT 101.180 62.950 101.600 63.020 ;
        RECT 44.210 62.440 45.980 62.510 ;
        RECT 46.990 61.340 48.760 62.930 ;
        RECT 105.510 62.800 108.230 64.450 ;
        RECT 116.650 64.340 117.210 66.760 ;
        RECT 129.040 66.290 132.350 67.380 ;
        RECT 129.460 65.640 130.740 66.290 ;
        RECT 123.130 64.380 123.450 64.680 ;
        RECT 127.480 64.520 128.760 64.700 ;
        RECT 129.040 64.450 132.350 65.640 ;
        RECT 118.240 62.950 121.550 62.960 ;
        RECT 120.590 62.920 120.780 62.950 ;
        RECT 129.040 62.800 132.600 64.450 ;
        RECT 105.510 62.760 108.220 62.800 ;
        RECT 129.040 62.760 132.590 62.800 ;
        RECT 44.210 60.690 45.980 60.850 ;
        RECT 46.990 59.590 48.760 61.180 ;
        RECT 49.850 61.030 52.350 62.510 ;
        RECT 129.040 62.470 132.350 62.760 ;
        RECT 49.850 60.830 52.380 61.030 ;
        RECT 44.210 58.940 45.980 59.100 ;
        RECT 46.990 57.840 48.760 59.430 ;
        RECT 44.210 57.190 45.980 57.350 ;
        RECT 46.990 56.090 48.760 57.680 ;
        RECT 44.210 55.510 45.980 55.600 ;
        RECT 49.850 55.510 52.350 60.830 ;
        RECT 94.630 58.660 96.610 58.670 ;
        RECT 101.050 58.310 101.610 60.730 ;
        RECT 110.610 58.310 111.170 60.730 ;
        RECT 116.140 59.570 117.280 60.160 ;
        RECT 115.650 58.730 117.280 59.570 ;
        RECT 129.460 59.140 130.740 61.980 ;
        RECT 117.590 58.660 119.060 58.670 ;
        RECT 121.440 58.490 122.720 58.670 ;
        RECT 127.480 58.650 128.760 58.840 ;
        RECT 94.630 57.990 94.700 58.170 ;
        RECT 111.220 57.300 111.230 57.680 ;
        RECT 59.490 54.040 59.520 54.050 ;
        RECT 44.730 53.900 46.500 54.010 ;
        RECT 50.370 53.900 52.870 54.010 ;
        RECT 58.810 53.740 59.520 54.040 ;
        RECT 58.810 53.700 59.490 53.740 ;
        RECT 44.210 52.310 45.980 52.400 ;
        RECT 44.210 50.560 45.980 50.720 ;
        RECT 46.990 50.230 48.760 51.820 ;
        RECT 44.210 48.810 45.980 48.970 ;
        RECT 46.990 48.480 48.760 50.070 ;
        RECT 44.210 47.060 45.980 47.220 ;
        RECT 46.990 46.730 48.760 48.320 ;
        RECT 49.850 47.080 52.350 52.400 ;
        RECT 58.800 47.650 59.500 53.700 ;
        RECT 63.570 52.350 66.990 53.580 ;
        RECT 94.630 53.120 94.710 53.300 ;
        RECT 69.270 52.350 69.280 52.800 ;
        RECT 121.440 52.620 122.720 52.810 ;
        RECT 125.920 52.720 127.780 55.710 ;
        RECT 63.570 52.330 69.310 52.350 ;
        RECT 63.570 51.090 66.990 52.330 ;
        RECT 69.270 51.610 69.280 52.330 ;
        RECT 74.950 52.000 76.680 52.050 ;
        RECT 110.940 52.000 112.670 52.050 ;
        RECT 69.270 51.560 69.320 51.610 ;
        RECT 69.270 51.460 69.330 51.560 ;
        RECT 63.570 49.140 66.990 50.380 ;
        RECT 69.280 50.340 69.330 51.460 ;
        RECT 63.570 49.130 69.310 49.140 ;
        RECT 63.570 47.890 66.990 49.130 ;
        RECT 70.950 48.470 72.680 50.310 ;
        RECT 58.810 47.450 59.500 47.650 ;
        RECT 49.850 46.880 52.380 47.080 ;
        RECT 44.210 45.400 45.980 45.470 ;
        RECT 46.990 44.980 48.760 46.570 ;
        RECT 49.850 45.400 52.350 46.880 ;
        RECT 74.950 45.560 77.870 52.000 ;
        RECT 82.700 50.550 83.260 51.090 ;
        RECT 78.230 46.560 80.790 48.470 ;
        RECT 91.120 46.720 91.190 46.900 ;
        RECT 96.430 46.720 96.500 46.900 ;
        RECT 106.830 46.560 109.390 48.470 ;
        RECT 85.770 46.310 86.880 46.540 ;
        RECT 90.030 46.370 90.620 46.480 ;
        RECT 97.000 46.370 97.590 46.480 ;
        RECT 100.740 46.310 101.850 46.540 ;
        RECT 75.640 45.510 77.870 45.560 ;
        RECT 78.230 43.320 80.790 46.290 ;
        RECT 81.890 44.880 82.240 44.890 ;
        RECT 81.890 44.720 81.900 44.880 ;
        RECT 82.070 44.720 82.240 44.880 ;
        RECT 105.380 44.880 105.730 44.890 ;
        RECT 105.380 44.720 105.550 44.880 ;
        RECT 105.720 44.720 105.730 44.880 ;
        RECT 75.550 43.160 77.280 43.220 ;
        RECT 44.210 42.180 45.980 42.270 ;
        RECT 44.210 40.430 45.980 40.590 ;
        RECT 46.990 40.100 48.760 41.690 ;
        RECT 44.210 38.680 45.980 38.840 ;
        RECT 46.990 38.350 48.760 39.940 ;
        RECT 44.210 36.930 45.980 37.090 ;
        RECT 46.990 36.600 48.760 38.190 ;
        RECT 49.850 36.950 52.350 42.270 ;
        RECT 63.550 41.880 66.970 43.110 ;
        RECT 75.550 43.060 78.470 43.160 ;
        RECT 85.770 43.070 86.880 43.340 ;
        RECT 90.030 43.090 90.620 43.280 ;
        RECT 97.000 43.090 97.590 43.280 ;
        RECT 100.740 43.070 101.850 43.340 ;
        RECT 103.590 43.200 103.680 43.500 ;
        RECT 106.830 43.320 109.390 46.290 ;
        RECT 109.750 45.560 112.670 52.000 ;
        RECT 115.650 51.130 117.280 51.300 ;
        RECT 117.590 51.190 118.040 51.420 ;
        RECT 115.650 51.060 118.110 51.130 ;
        RECT 115.650 50.460 117.280 51.060 ;
        RECT 116.140 50.310 117.280 50.460 ;
        RECT 114.940 49.870 117.280 50.310 ;
        RECT 114.940 48.470 116.670 49.870 ;
        RECT 119.880 46.690 121.740 49.680 ;
        RECT 125.920 49.670 127.780 52.660 ;
        RECT 109.750 45.510 111.980 45.560 ;
        RECT 119.880 43.640 121.740 46.630 ;
        RECT 63.550 41.860 69.290 41.880 ;
        RECT 63.550 40.620 66.970 41.860 ;
        RECT 63.550 38.670 66.970 39.910 ;
        RECT 71.550 39.590 73.280 41.430 ;
        RECT 75.550 41.150 80.790 43.060 ;
        RECT 106.830 41.150 109.390 43.060 ;
        RECT 63.550 38.660 69.290 38.670 ;
        RECT 63.550 37.420 66.970 38.660 ;
        RECT 49.850 36.750 52.380 36.950 ;
        RECT 44.210 35.270 45.980 35.340 ;
        RECT 46.990 34.850 48.760 36.440 ;
        RECT 49.850 35.270 52.350 36.750 ;
        RECT 75.550 36.720 78.470 41.150 ;
        RECT 83.750 41.020 83.880 41.080 ;
        RECT 83.750 40.900 83.820 41.020 ;
        RECT 78.830 37.720 81.390 39.630 ;
        RECT 76.240 36.670 78.470 36.720 ;
        RECT 78.830 34.480 81.390 37.470 ;
        RECT 86.370 37.430 87.480 37.700 ;
        RECT 90.630 37.490 91.220 37.650 ;
        RECT 84.190 36.510 84.280 36.590 ;
        RECT 82.670 36.010 82.840 36.070 ;
        RECT 82.490 36.000 82.840 36.010 ;
        RECT 82.490 35.900 82.500 36.000 ;
        RECT 82.670 35.900 82.840 36.000 ;
        RECT 83.960 34.530 86.920 34.540 ;
        RECT 83.960 34.380 84.370 34.530 ;
        RECT 89.650 34.440 90.030 34.540 ;
        RECT 83.960 34.370 84.550 34.380 ;
        RECT 44.170 33.120 45.940 33.210 ;
        RECT 44.170 31.370 45.940 31.530 ;
        RECT 46.950 31.040 48.720 32.630 ;
        RECT 24.030 27.490 26.400 30.360 ;
        RECT 27.870 28.410 28.430 30.380 ;
        RECT 44.170 29.620 45.940 29.780 ;
        RECT 46.950 29.290 48.720 30.880 ;
        RECT 44.170 27.870 45.940 28.030 ;
        RECT 46.950 27.540 48.720 29.130 ;
        RECT 58.800 27.930 60.550 33.900 ;
        RECT 63.580 32.610 67.000 33.840 ;
        RECT 83.960 32.610 84.370 34.370 ;
        RECT 86.370 34.230 87.480 34.420 ;
        RECT 93.680 34.400 94.080 34.540 ;
        RECT 90.630 34.250 91.220 34.400 ;
        RECT 63.580 32.590 69.320 32.610 ;
        RECT 63.580 31.350 67.000 32.590 ;
        RECT 83.850 32.190 84.370 32.610 ;
        RECT 83.850 31.990 84.360 32.190 ;
        RECT 83.850 31.460 84.370 31.990 ;
        RECT 63.580 29.400 67.000 30.640 ;
        RECT 63.580 29.390 69.320 29.400 ;
        RECT 63.580 28.150 67.000 29.390 ;
        RECT 83.960 28.500 84.370 31.460 ;
        RECT 58.800 27.900 61.820 27.930 ;
        RECT 60.940 27.740 61.820 27.900 ;
        RECT 44.170 26.210 45.940 26.280 ;
        RECT 46.950 25.790 48.720 27.380 ;
        RECT 60.700 22.370 62.720 26.460 ;
        RECT 60.700 22.340 65.520 22.370 ;
        RECT 52.320 22.250 55.710 22.340 ;
        RECT 57.930 22.280 65.520 22.340 ;
        RECT 67.740 22.280 71.130 22.370 ;
        RECT 57.930 22.250 65.990 22.280 ;
        RECT 18.780 20.850 19.400 20.940 ;
        RECT 18.780 15.240 22.640 20.850 ;
        RECT 52.320 16.640 56.180 22.250 ;
        RECT 55.560 16.550 56.180 16.640 ;
        RECT 57.460 20.770 65.990 22.250 ;
        RECT 57.460 16.640 61.320 20.770 ;
        RECT 62.130 16.670 65.990 20.770 ;
        RECT 57.460 16.550 58.080 16.640 ;
        RECT 65.370 16.580 65.990 16.670 ;
        RECT 67.270 16.670 71.130 22.280 ;
        RECT 67.270 16.580 67.890 16.670 ;
        RECT 19.250 15.150 22.640 15.240 ;
        RECT 104.400 1.890 105.250 16.370 ;
        RECT 105.360 8.320 110.410 16.370 ;
        RECT 105.360 6.710 107.530 8.320 ;
        RECT 107.780 6.770 110.410 8.320 ;
        RECT 108.240 6.710 110.410 6.770 ;
        RECT 105.360 1.890 110.410 6.710 ;
        RECT 105.360 1.880 109.450 1.890 ;
        RECT 104.400 0.270 105.250 1.880 ;
        RECT 105.360 0.270 110.410 1.880 ;
      LAYER li1 ;
        RECT 0.460 71.870 0.630 72.540 ;
        RECT 15.120 72.050 15.350 72.740 ;
        RECT 19.820 72.000 20.050 72.690 ;
        RECT 86.480 71.260 87.030 71.690 ;
        RECT 130.980 71.260 131.530 71.690 ;
        RECT 15.120 69.590 15.350 69.750 ;
        RECT 0.420 69.080 0.590 69.410 ;
        RECT 0.660 68.970 0.750 69.110 ;
        RECT 1.820 69.080 1.990 69.410 ;
        RECT 0.550 68.790 1.550 68.970 ;
        RECT 2.040 68.960 2.120 69.110 ;
        RECT 3.750 69.000 4.420 69.170 ;
        RECT 1.950 68.790 2.960 68.960 ;
        RECT 12.560 68.610 15.870 69.590 ;
        RECT 86.480 69.530 87.030 69.960 ;
        RECT 130.980 69.530 131.530 69.960 ;
        RECT 86.060 68.730 86.260 69.080 ;
        RECT 87.540 68.830 88.070 69.000 ;
        RECT 129.940 68.830 130.470 69.000 ;
        RECT 86.050 68.700 86.260 68.730 ;
        RECT 131.750 68.730 131.950 69.080 ;
        RECT 131.750 68.700 131.960 68.730 ;
        RECT 1.620 68.260 1.940 68.300 ;
        RECT 1.610 68.110 1.940 68.260 ;
        RECT 0.880 67.940 2.960 68.110 ;
        RECT 3.490 68.080 4.160 68.250 ;
        RECT 15.120 68.050 15.350 68.610 ;
        RECT 17.810 67.970 17.980 68.300 ;
        RECT 18.490 67.970 18.660 68.300 ;
        RECT 86.050 68.120 86.270 68.700 ;
        RECT 86.050 68.110 86.260 68.120 ;
        RECT 1.060 67.530 2.880 67.700 ;
        RECT 3.580 67.540 3.790 67.970 ;
        RECT 86.430 67.940 86.620 67.950 ;
        RECT 3.600 67.520 3.770 67.540 ;
        RECT 17.010 67.520 17.330 67.560 ;
        RECT 1.620 67.420 1.940 67.460 ;
        RECT 1.610 67.290 1.940 67.420 ;
        RECT 17.000 67.330 17.330 67.520 ;
        RECT 17.880 67.410 18.050 67.760 ;
        RECT 86.420 67.650 86.620 67.940 ;
        RECT 18.370 67.600 18.690 67.640 ;
        RECT 18.360 67.410 18.690 67.600 ;
        RECT 19.060 67.590 19.380 67.630 ;
        RECT 17.010 67.300 17.330 67.330 ;
        RECT 0.880 67.120 2.960 67.290 ;
        RECT 17.450 67.150 18.050 67.410 ;
        RECT 18.370 67.380 18.690 67.410 ;
        RECT 19.050 67.400 19.380 67.590 ;
        RECT 19.060 67.370 19.380 67.400 ;
        RECT 86.360 67.320 86.630 67.650 ;
        RECT 26.380 67.170 26.550 67.190 ;
        RECT 3.490 66.650 4.160 66.820 ;
        RECT 0.880 66.280 1.550 66.450 ;
        RECT 2.280 66.280 2.960 66.450 ;
        RECT 3.160 66.160 3.350 66.300 ;
        RECT 3.160 66.070 4.430 66.160 ;
        RECT 3.290 65.990 4.430 66.070 ;
        RECT 12.560 65.810 15.870 66.790 ;
        RECT 3.280 65.560 3.450 65.600 ;
        RECT 3.280 65.530 3.660 65.560 ;
        RECT 0.880 65.160 1.550 65.330 ;
        RECT 1.850 65.200 2.020 65.530 ;
        RECT 3.280 65.340 3.670 65.530 ;
        RECT 3.760 65.380 4.430 65.550 ;
        RECT 2.080 65.160 2.960 65.330 ;
        RECT 3.280 65.300 3.660 65.340 ;
        RECT 3.280 65.270 3.450 65.300 ;
        RECT 1.600 64.620 1.920 64.660 ;
        RECT 3.030 64.640 3.350 64.680 ;
        RECT 1.590 64.490 1.920 64.620 ;
        RECT 3.020 64.490 3.350 64.640 ;
        RECT 0.870 64.320 4.450 64.490 ;
        RECT 12.560 64.260 15.870 65.240 ;
        RECT 16.510 64.290 16.680 66.940 ;
        RECT 17.880 66.750 18.050 67.150 ;
        RECT 23.490 67.000 26.550 67.170 ;
        RECT 26.380 66.350 26.550 67.000 ;
        RECT 86.820 66.840 86.990 68.450 ;
        RECT 92.970 68.440 93.160 68.670 ;
        RECT 86.810 66.650 86.990 66.840 ;
        RECT 87.650 66.750 87.820 68.440 ;
        RECT 88.240 68.250 88.570 68.420 ;
        RECT 89.590 68.250 89.940 68.420 ;
        RECT 93.250 68.390 94.130 68.560 ;
        RECT 93.440 68.000 93.630 68.110 ;
        RECT 93.330 67.880 93.630 68.000 ;
        RECT 93.960 68.000 94.130 68.390 ;
        RECT 93.330 67.830 93.550 67.880 ;
        RECT 93.960 67.830 94.350 68.000 ;
        RECT 105.810 67.900 106.040 68.590 ;
        RECT 130.180 67.900 130.410 68.590 ;
        RECT 88.240 67.460 88.570 67.630 ;
        RECT 89.590 67.460 89.940 67.630 ;
        RECT 125.410 67.610 125.730 67.650 ;
        RECT 125.410 67.420 125.740 67.610 ;
        RECT 125.410 67.390 125.730 67.420 ;
        RECT 92.040 67.040 92.360 67.080 ;
        RECT 93.290 67.040 94.370 67.210 ;
        RECT 94.700 67.040 95.780 67.210 ;
        RECT 92.030 66.850 92.360 67.040 ;
        RECT 88.240 66.670 88.570 66.840 ;
        RECT 89.590 66.670 89.930 66.840 ;
        RECT 92.040 66.820 92.360 66.850 ;
        RECT 130.190 66.750 130.360 67.900 ;
        RECT 131.020 66.840 131.190 68.450 ;
        RECT 131.740 68.120 131.960 68.700 ;
        RECT 131.750 68.110 131.960 68.120 ;
        RECT 131.390 67.940 131.580 67.950 ;
        RECT 131.390 67.650 131.590 67.940 ;
        RECT 131.380 67.320 131.670 67.650 ;
        RECT 92.970 66.450 93.160 66.680 ;
        RECT 131.020 66.650 131.200 66.840 ;
        RECT 26.380 66.180 27.650 66.350 ;
        RECT 93.270 66.250 93.350 66.420 ;
        RECT 0.810 64.040 1.130 64.080 ;
        RECT 1.740 64.040 2.060 64.080 ;
        RECT 2.440 64.040 2.760 64.080 ;
        RECT 3.180 64.040 3.500 64.080 ;
        RECT 0.800 63.850 1.130 64.040 ;
        RECT 1.730 63.850 2.060 64.040 ;
        RECT 2.430 63.850 2.760 64.040 ;
        RECT 3.170 63.870 3.500 64.040 ;
        RECT 3.890 64.030 4.210 64.070 ;
        RECT 3.880 63.870 4.210 64.030 ;
        RECT 16.510 63.900 16.690 64.290 ;
        RECT 26.380 63.920 26.550 66.180 ;
        RECT 93.830 66.100 94.040 66.530 ;
        RECT 93.850 66.080 94.020 66.100 ;
        RECT 28.500 64.960 28.670 65.850 ;
        RECT 86.730 65.230 87.280 65.660 ;
        RECT 92.030 65.350 92.350 65.390 ;
        RECT 92.980 65.380 93.170 65.610 ;
        RECT 93.300 65.510 93.350 65.680 ;
        RECT 93.440 65.560 93.630 65.790 ;
        RECT 94.440 65.680 94.610 66.250 ;
        RECT 98.720 66.100 98.910 66.420 ;
        RECT 119.100 66.100 119.290 66.420 ;
        RECT 98.720 66.010 99.000 66.100 ;
        RECT 95.360 65.870 99.000 66.010 ;
        RECT 119.010 66.010 119.290 66.100 ;
        RECT 130.020 66.210 130.350 66.380 ;
        RECT 130.460 66.300 130.790 66.470 ;
        RECT 119.010 65.870 122.650 66.010 ;
        RECT 130.020 65.930 130.380 66.210 ;
        RECT 95.360 65.830 98.910 65.870 ;
        RECT 93.720 65.650 93.770 65.660 ;
        RECT 94.350 65.650 94.430 65.660 ;
        RECT 93.720 65.610 94.430 65.650 ;
        RECT 93.720 65.570 94.450 65.610 ;
        RECT 93.680 65.450 94.520 65.570 ;
        RECT 98.720 65.410 98.910 65.830 ;
        RECT 119.100 65.830 122.650 65.870 ;
        RECT 119.100 65.410 119.290 65.830 ;
        RECT 127.950 65.680 128.270 65.720 ;
        RECT 86.810 65.090 86.990 65.230 ;
        RECT 86.360 64.280 86.630 64.610 ;
        RECT 86.420 63.990 86.620 64.280 ;
        RECT 86.430 63.980 86.620 63.990 ;
        RECT 86.820 63.930 86.990 65.090 ;
        RECT 3.170 63.850 4.210 63.870 ;
        RECT 16.290 63.860 16.690 63.900 ;
        RECT 26.150 63.880 26.550 63.920 ;
        RECT 0.810 63.820 1.130 63.850 ;
        RECT 1.740 63.820 2.060 63.850 ;
        RECT 2.440 63.820 2.760 63.850 ;
        RECT 3.180 63.820 4.210 63.850 ;
        RECT 0.920 63.810 4.210 63.820 ;
        RECT 0.920 63.650 4.350 63.810 ;
        RECT 16.280 63.670 16.690 63.860 ;
        RECT 26.140 63.770 26.550 63.880 ;
        RECT 86.050 63.810 86.260 63.820 ;
        RECT 26.140 63.690 26.470 63.770 ;
        RECT 3.500 63.640 4.350 63.650 ;
        RECT 16.290 63.640 16.690 63.670 ;
        RECT 26.150 63.660 26.470 63.690 ;
        RECT 16.510 63.560 16.690 63.640 ;
        RECT 86.050 63.230 86.270 63.810 ;
        RECT 86.730 63.500 87.280 63.930 ;
        RECT 86.820 63.480 86.990 63.500 ;
        RECT 87.650 63.490 87.820 65.180 ;
        RECT 88.240 65.090 88.570 65.260 ;
        RECT 89.590 65.090 89.930 65.260 ;
        RECT 92.020 65.160 92.350 65.350 ;
        RECT 124.940 65.230 125.490 65.660 ;
        RECT 127.950 65.490 128.280 65.680 ;
        RECT 127.950 65.460 128.270 65.490 ;
        RECT 128.350 65.470 128.550 65.800 ;
        RECT 128.940 65.610 129.140 65.800 ;
        RECT 129.670 65.760 130.380 65.930 ;
        RECT 129.610 65.640 129.930 65.680 ;
        RECT 128.630 65.280 128.820 65.290 ;
        RECT 128.830 65.280 129.180 65.610 ;
        RECT 129.610 65.450 129.940 65.640 ;
        RECT 129.610 65.420 129.930 65.450 ;
        RECT 92.030 65.130 92.350 65.160 ;
        RECT 93.290 64.720 94.370 64.890 ;
        RECT 94.690 64.720 95.930 64.890 ;
        RECT 125.410 64.850 125.730 64.890 ;
        RECT 120.130 64.790 120.360 64.830 ;
        RECT 125.410 64.660 125.740 64.850 ;
        RECT 127.720 64.770 127.890 65.100 ;
        RECT 127.900 65.030 128.220 65.070 ;
        RECT 127.900 64.840 128.230 65.030 ;
        RECT 127.900 64.810 128.220 64.840 ;
        RECT 128.350 64.810 128.550 65.140 ;
        RECT 128.630 64.950 129.180 65.280 ;
        RECT 125.410 64.630 125.730 64.660 ;
        RECT 128.830 64.620 129.180 64.950 ;
        RECT 88.240 64.300 88.570 64.470 ;
        RECT 89.590 64.300 89.940 64.470 ;
        RECT 95.020 64.400 95.190 64.460 ;
        RECT 129.670 64.440 130.370 65.320 ;
        RECT 131.020 65.090 131.200 65.280 ;
        RECT 93.430 64.100 93.620 64.210 ;
        RECT 95.000 64.190 95.210 64.400 ;
        RECT 95.020 64.120 95.190 64.190 ;
        RECT 93.330 63.980 93.620 64.100 ;
        RECT 93.890 64.090 94.350 64.100 ;
        RECT 93.330 63.930 93.540 63.980 ;
        RECT 93.890 63.940 94.360 64.090 ;
        RECT 129.010 64.050 129.200 64.280 ;
        RECT 130.190 64.020 130.360 64.440 ;
        RECT 93.890 63.930 94.350 63.940 ;
        RECT 88.240 63.510 88.570 63.680 ;
        RECT 89.590 63.510 89.940 63.680 ;
        RECT 93.000 63.590 93.190 63.700 ;
        RECT 93.890 63.590 94.080 63.930 ;
        RECT 93.000 63.470 94.080 63.590 ;
        RECT 93.120 63.410 94.080 63.470 ;
        RECT 105.810 63.240 106.040 63.930 ;
        RECT 124.940 63.500 125.490 63.930 ;
        RECT 127.720 63.510 127.890 63.840 ;
        RECT 127.900 63.770 128.220 63.800 ;
        RECT 127.900 63.580 128.230 63.770 ;
        RECT 127.900 63.540 128.220 63.580 ;
        RECT 128.350 63.470 128.550 63.800 ;
        RECT 128.830 63.660 129.180 63.990 ;
        RECT 129.660 63.930 130.360 64.020 ;
        RECT 129.660 63.840 130.410 63.930 ;
        RECT 128.630 63.330 129.180 63.660 ;
        RECT 128.630 63.320 128.820 63.330 ;
        RECT 86.050 63.200 86.260 63.230 ;
        RECT 86.060 62.850 86.260 63.200 ;
        RECT 127.950 63.120 128.270 63.150 ;
        RECT 86.310 62.700 86.510 63.050 ;
        RECT 87.540 62.970 88.070 63.100 ;
        RECT 87.540 62.930 88.320 62.970 ;
        RECT 87.790 62.800 88.320 62.930 ;
        RECT 123.900 62.800 124.430 62.970 ;
        RECT 86.300 62.670 86.510 62.700 ;
        RECT 25.300 62.520 26.820 62.530 ;
        RECT 25.300 61.730 26.850 62.520 ;
        RECT 48.650 62.460 49.000 62.560 ;
        RECT 52.240 62.510 52.410 62.550 ;
        RECT 51.260 62.490 52.410 62.510 ;
        RECT 50.310 62.460 50.770 62.490 ;
        RECT 47.240 62.290 48.000 62.460 ;
        RECT 48.250 62.290 49.420 62.460 ;
        RECT 49.660 62.320 50.770 62.460 ;
        RECT 51.220 62.320 52.410 62.490 ;
        RECT 49.660 62.290 50.480 62.320 ;
        RECT 47.240 62.280 47.470 62.290 ;
        RECT 47.200 61.840 47.470 62.280 ;
        RECT 50.220 62.150 50.480 62.290 ;
        RECT 48.680 61.840 49.010 62.100 ;
        RECT 49.630 62.050 49.920 62.080 ;
        RECT 49.590 61.880 49.920 62.050 ;
        RECT 49.630 61.840 49.920 61.880 ;
        RECT 50.220 61.980 51.400 62.150 ;
        RECT 86.300 62.090 86.520 62.670 ;
        RECT 86.300 62.080 86.510 62.090 ;
        RECT 50.220 61.840 50.480 61.980 ;
        RECT 46.650 61.700 46.820 61.760 ;
        RECT 46.620 61.480 46.840 61.700 ;
        RECT 47.170 61.660 47.500 61.840 ;
        RECT 47.750 61.670 49.910 61.840 ;
        RECT 50.150 61.670 50.480 61.840 ;
        RECT 50.620 61.830 51.400 61.980 ;
        RECT 50.250 61.620 50.480 61.670 ;
        RECT 46.650 61.430 46.820 61.480 ;
        RECT 50.250 61.390 50.420 61.620 ;
        RECT 50.770 61.480 50.980 61.810 ;
        RECT 51.220 61.540 51.400 61.830 ;
        RECT 51.680 61.820 52.010 61.990 ;
        RECT 86.680 61.910 86.870 61.920 ;
        RECT 50.040 61.380 50.420 61.390 ;
        RECT 50.040 61.320 50.510 61.380 ;
        RECT 51.760 61.360 51.940 61.820 ;
        RECT 51.950 61.640 52.570 61.810 ;
        RECT 86.670 61.620 86.870 61.910 ;
        RECT 49.700 61.270 50.510 61.320 ;
        RECT 49.690 61.210 50.510 61.270 ;
        RECT 49.690 61.150 50.430 61.210 ;
        RECT 50.980 61.190 51.940 61.360 ;
        RECT 86.590 61.290 86.880 61.620 ;
        RECT 50.040 61.100 50.430 61.150 ;
        RECT 87.070 60.810 87.240 62.420 ;
        RECT 87.850 61.870 88.080 62.560 ;
        RECT 95.270 61.950 100.330 62.780 ;
        RECT 125.710 62.700 125.910 63.050 ;
        RECT 127.950 62.930 128.280 63.120 ;
        RECT 127.950 62.890 128.270 62.930 ;
        RECT 128.350 62.810 128.550 63.140 ;
        RECT 128.830 63.000 129.180 63.330 ;
        RECT 129.660 63.420 129.980 63.460 ;
        RECT 129.660 63.230 129.990 63.420 ;
        RECT 130.180 63.240 130.410 63.840 ;
        RECT 131.020 63.480 131.190 65.090 ;
        RECT 131.380 64.280 131.670 64.610 ;
        RECT 131.390 63.990 131.590 64.280 ;
        RECT 131.390 63.980 131.580 63.990 ;
        RECT 131.750 63.810 131.960 63.820 ;
        RECT 131.740 63.230 131.960 63.810 ;
        RECT 129.660 63.200 129.980 63.230 ;
        RECT 131.750 63.200 131.960 63.230 ;
        RECT 128.940 62.810 129.140 63.000 ;
        RECT 129.940 62.930 130.470 63.100 ;
        RECT 131.750 62.850 131.950 63.200 ;
        RECT 125.710 62.670 125.920 62.700 ;
        RECT 99.780 61.870 100.260 61.950 ;
        RECT 124.140 61.870 124.370 62.560 ;
        RECT 48.650 60.710 49.000 60.810 ;
        RECT 52.240 60.760 52.410 60.800 ;
        RECT 51.260 60.740 52.410 60.760 ;
        RECT 50.310 60.710 50.770 60.740 ;
        RECT 47.240 60.540 48.000 60.710 ;
        RECT 48.250 60.540 49.420 60.710 ;
        RECT 49.660 60.570 50.770 60.710 ;
        RECT 51.220 60.570 52.410 60.740 ;
        RECT 87.060 60.620 87.240 60.810 ;
        RECT 87.900 60.720 88.070 61.870 ;
        RECT 99.780 61.770 100.110 61.870 ;
        RECT 99.780 61.620 99.930 61.770 ;
        RECT 92.530 61.580 92.850 61.620 ;
        RECT 92.520 61.390 92.850 61.580 ;
        RECT 92.530 61.360 92.850 61.390 ;
        RECT 119.370 61.580 119.690 61.620 ;
        RECT 119.370 61.390 119.700 61.580 ;
        RECT 119.370 61.360 119.690 61.390 ;
        RECT 124.150 60.720 124.320 61.870 ;
        RECT 124.980 60.810 125.150 62.420 ;
        RECT 125.700 62.090 125.920 62.670 ;
        RECT 127.950 62.680 128.270 62.720 ;
        RECT 127.950 62.490 128.280 62.680 ;
        RECT 127.950 62.460 128.270 62.490 ;
        RECT 128.350 62.470 128.550 62.800 ;
        RECT 128.940 62.610 129.140 62.800 ;
        RECT 129.650 62.700 129.970 62.740 ;
        RECT 128.630 62.280 128.820 62.290 ;
        RECT 128.830 62.280 129.180 62.610 ;
        RECT 129.650 62.510 129.980 62.700 ;
        RECT 129.650 62.480 129.970 62.510 ;
        RECT 125.710 62.080 125.920 62.090 ;
        RECT 125.350 61.910 125.540 61.920 ;
        RECT 125.350 61.620 125.550 61.910 ;
        RECT 127.720 61.770 127.890 62.100 ;
        RECT 127.900 62.030 128.220 62.070 ;
        RECT 127.900 61.840 128.230 62.030 ;
        RECT 127.900 61.810 128.220 61.840 ;
        RECT 128.350 61.810 128.550 62.140 ;
        RECT 128.630 61.950 129.180 62.280 ;
        RECT 128.830 61.690 129.180 61.950 ;
        RECT 128.830 61.620 129.200 61.690 ;
        RECT 125.340 61.290 125.630 61.620 ;
        RECT 129.010 61.460 129.200 61.620 ;
        RECT 129.660 61.560 130.360 61.740 ;
        RECT 124.980 60.620 125.160 60.810 ;
        RECT 49.660 60.540 50.480 60.570 ;
        RECT 47.240 60.530 47.470 60.540 ;
        RECT 47.200 60.090 47.470 60.530 ;
        RECT 50.220 60.400 50.480 60.540 ;
        RECT 127.720 60.510 127.890 60.840 ;
        RECT 127.900 60.770 128.220 60.800 ;
        RECT 127.900 60.580 128.230 60.770 ;
        RECT 127.900 60.540 128.220 60.580 ;
        RECT 128.350 60.470 128.550 60.800 ;
        RECT 128.830 60.660 129.180 60.990 ;
        RECT 48.680 60.090 49.010 60.350 ;
        RECT 49.630 60.300 49.920 60.330 ;
        RECT 49.590 60.130 49.920 60.300 ;
        RECT 49.630 60.090 49.920 60.130 ;
        RECT 50.220 60.230 51.400 60.400 ;
        RECT 50.220 60.090 50.480 60.230 ;
        RECT 46.650 59.950 46.820 60.010 ;
        RECT 46.620 59.730 46.840 59.950 ;
        RECT 47.170 59.910 47.500 60.090 ;
        RECT 47.750 59.920 49.910 60.090 ;
        RECT 50.150 59.920 50.480 60.090 ;
        RECT 50.620 60.080 51.400 60.230 ;
        RECT 50.250 59.870 50.480 59.920 ;
        RECT 46.650 59.680 46.820 59.730 ;
        RECT 50.250 59.640 50.420 59.870 ;
        RECT 50.770 59.730 50.980 60.060 ;
        RECT 51.220 59.790 51.400 60.080 ;
        RECT 51.680 60.070 52.010 60.240 ;
        RECT 98.970 60.070 99.160 60.390 ;
        RECT 113.060 60.070 113.250 60.390 ;
        RECT 123.380 60.220 123.700 60.260 ;
        RECT 50.040 59.630 50.420 59.640 ;
        RECT 50.040 59.570 50.510 59.630 ;
        RECT 51.760 59.610 51.940 60.070 ;
        RECT 51.950 59.890 52.570 60.060 ;
        RECT 98.970 59.980 99.250 60.070 ;
        RECT 95.610 59.840 99.250 59.980 ;
        RECT 112.970 59.980 113.250 60.070 ;
        RECT 123.370 60.030 123.700 60.220 ;
        RECT 123.380 60.020 123.700 60.030 ;
        RECT 123.370 60.000 123.700 60.020 ;
        RECT 123.980 60.180 124.310 60.350 ;
        RECT 124.420 60.270 124.750 60.440 ;
        RECT 128.630 60.330 129.180 60.660 ;
        RECT 129.670 60.490 130.370 61.140 ;
        RECT 128.630 60.320 128.820 60.330 ;
        RECT 112.970 59.840 116.610 59.980 ;
        RECT 95.610 59.800 99.160 59.840 ;
        RECT 49.700 59.520 50.510 59.570 ;
        RECT 49.690 59.460 50.510 59.520 ;
        RECT 49.690 59.400 50.430 59.460 ;
        RECT 50.980 59.440 51.940 59.610 ;
        RECT 50.040 59.350 50.430 59.400 ;
        RECT 22.530 59.220 22.850 59.260 ;
        RECT 23.620 59.230 23.940 59.270 ;
        RECT 22.530 59.150 22.860 59.220 ;
        RECT 22.530 59.000 22.900 59.150 ;
        RECT 22.700 58.820 22.900 59.000 ;
        RECT 23.290 58.820 23.490 59.150 ;
        RECT 23.620 59.040 23.950 59.230 ;
        RECT 23.620 59.010 23.940 59.040 ;
        RECT 48.650 58.960 49.000 59.060 ;
        RECT 52.240 59.010 52.410 59.050 ;
        RECT 51.260 58.990 52.410 59.010 ;
        RECT 50.310 58.960 50.770 58.990 ;
        RECT 47.240 58.790 48.000 58.960 ;
        RECT 48.250 58.790 49.420 58.960 ;
        RECT 49.660 58.820 50.770 58.960 ;
        RECT 51.220 58.820 52.410 58.990 ;
        RECT 49.660 58.790 50.480 58.820 ;
        RECT 47.240 58.780 47.470 58.790 ;
        RECT 22.150 58.510 22.480 58.680 ;
        RECT 20.990 58.310 21.310 58.350 ;
        RECT 47.200 58.340 47.470 58.780 ;
        RECT 50.220 58.650 50.480 58.790 ;
        RECT 48.680 58.340 49.010 58.600 ;
        RECT 49.630 58.550 49.920 58.580 ;
        RECT 49.590 58.380 49.920 58.550 ;
        RECT 49.630 58.340 49.920 58.380 ;
        RECT 50.220 58.480 51.400 58.650 ;
        RECT 73.270 58.570 73.940 59.440 ;
        RECT 85.550 58.590 87.650 59.440 ;
        RECT 98.970 59.380 99.160 59.800 ;
        RECT 113.060 59.800 117.280 59.840 ;
        RECT 113.060 59.380 113.250 59.800 ;
        RECT 114.040 59.660 114.680 59.800 ;
        RECT 115.060 59.670 115.410 59.800 ;
        RECT 115.510 59.710 115.840 59.800 ;
        RECT 115.590 59.630 115.840 59.710 ;
        RECT 116.140 59.660 117.280 59.800 ;
        RECT 114.440 59.280 114.610 59.290 ;
        RECT 114.440 59.240 114.840 59.280 ;
        RECT 50.220 58.340 50.480 58.480 ;
        RECT 20.990 58.120 21.320 58.310 ;
        RECT 22.540 58.230 22.860 58.270 ;
        RECT 23.630 58.240 23.950 58.280 ;
        RECT 22.540 58.160 22.870 58.230 ;
        RECT 22.880 58.160 23.050 58.210 ;
        RECT 23.370 58.160 23.560 58.200 ;
        RECT 22.540 58.130 23.050 58.160 ;
        RECT 23.300 58.130 23.560 58.160 ;
        RECT 20.990 58.090 21.310 58.120 ;
        RECT 21.010 58.020 21.220 58.090 ;
        RECT 22.540 58.010 23.560 58.130 ;
        RECT 23.630 58.050 23.960 58.240 ;
        RECT 46.650 58.200 46.820 58.260 ;
        RECT 23.630 58.020 23.950 58.050 ;
        RECT 22.710 57.970 23.560 58.010 ;
        RECT 46.620 57.980 46.840 58.200 ;
        RECT 47.170 58.160 47.500 58.340 ;
        RECT 47.750 58.170 49.910 58.340 ;
        RECT 50.150 58.170 50.480 58.340 ;
        RECT 50.620 58.330 51.400 58.480 ;
        RECT 50.250 58.120 50.480 58.170 ;
        RECT 22.710 57.880 23.500 57.970 ;
        RECT 46.650 57.930 46.820 57.980 ;
        RECT 50.250 57.890 50.420 58.120 ;
        RECT 50.770 57.980 50.980 58.310 ;
        RECT 51.220 58.040 51.400 58.330 ;
        RECT 51.680 58.320 52.010 58.490 ;
        RECT 22.710 57.830 23.060 57.880 ;
        RECT 23.300 57.830 23.500 57.880 ;
        RECT 50.040 57.880 50.420 57.890 ;
        RECT 22.880 57.820 23.060 57.830 ;
        RECT 50.040 57.820 50.510 57.880 ;
        RECT 51.760 57.860 51.940 58.320 ;
        RECT 51.950 58.140 52.570 58.310 ;
        RECT 86.590 58.250 86.880 58.580 ;
        RECT 86.670 57.960 86.870 58.250 ;
        RECT 86.680 57.950 86.870 57.960 ;
        RECT 49.700 57.770 50.510 57.820 ;
        RECT 49.690 57.710 50.510 57.770 ;
        RECT 22.160 57.520 22.490 57.690 ;
        RECT 49.690 57.650 50.430 57.710 ;
        RECT 50.980 57.690 51.940 57.860 ;
        RECT 86.300 57.780 86.510 57.790 ;
        RECT 50.040 57.600 50.430 57.650 ;
        RECT 20.970 57.390 21.290 57.430 ;
        RECT 20.970 57.200 21.300 57.390 ;
        RECT 22.540 57.240 22.860 57.280 ;
        RECT 23.630 57.250 23.950 57.290 ;
        RECT 20.970 57.170 21.290 57.200 ;
        RECT 22.540 57.170 22.870 57.240 ;
        RECT 22.540 57.020 22.910 57.170 ;
        RECT 22.710 56.840 22.910 57.020 ;
        RECT 23.300 56.840 23.500 57.170 ;
        RECT 23.630 57.060 23.960 57.250 ;
        RECT 48.650 57.210 49.000 57.310 ;
        RECT 52.240 57.260 52.410 57.300 ;
        RECT 51.260 57.240 52.410 57.260 ;
        RECT 50.310 57.210 50.770 57.240 ;
        RECT 23.630 57.030 23.950 57.060 ;
        RECT 47.240 57.040 48.000 57.210 ;
        RECT 48.250 57.040 49.420 57.210 ;
        RECT 49.660 57.070 50.770 57.210 ;
        RECT 51.220 57.070 52.410 57.240 ;
        RECT 86.300 57.200 86.520 57.780 ;
        RECT 87.070 57.450 87.240 58.590 ;
        RECT 87.900 57.900 88.070 59.150 ;
        RECT 114.440 59.050 114.850 59.240 ;
        RECT 115.050 59.210 115.240 59.320 ;
        RECT 115.050 59.090 115.390 59.210 ;
        RECT 114.440 59.020 114.840 59.050 ;
        RECT 115.100 59.040 115.390 59.090 ;
        RECT 114.440 58.990 114.610 59.020 ;
        RECT 115.670 58.950 115.840 59.630 ;
        RECT 121.910 59.650 122.230 59.690 ;
        RECT 121.910 59.460 122.240 59.650 ;
        RECT 121.910 59.430 122.230 59.460 ;
        RECT 122.310 59.440 122.510 59.770 ;
        RECT 122.900 59.580 123.100 59.770 ;
        RECT 123.370 59.690 123.540 60.000 ;
        RECT 123.980 59.900 124.340 60.180 ;
        RECT 123.630 59.730 124.340 59.900 ;
        RECT 127.950 60.120 128.270 60.150 ;
        RECT 127.950 59.930 128.280 60.120 ;
        RECT 127.950 59.890 128.270 59.930 ;
        RECT 128.350 59.810 128.550 60.140 ;
        RECT 128.830 60.000 129.180 60.330 ;
        RECT 129.570 60.260 130.370 60.490 ;
        RECT 129.570 60.230 129.890 60.260 ;
        RECT 128.940 59.810 129.140 60.000 ;
        RECT 129.670 59.650 130.380 59.820 ;
        RECT 123.570 59.610 123.890 59.650 ;
        RECT 116.180 59.280 116.350 59.290 ;
        RECT 116.180 59.240 116.510 59.280 ;
        RECT 116.180 59.050 116.520 59.240 ;
        RECT 117.160 59.220 117.350 59.330 ;
        RECT 117.040 59.210 117.350 59.220 ;
        RECT 116.790 59.100 117.350 59.210 ;
        RECT 122.590 59.250 122.780 59.260 ;
        RECT 122.790 59.250 123.140 59.580 ;
        RECT 123.570 59.430 123.900 59.610 ;
        RECT 123.530 59.420 123.900 59.430 ;
        RECT 123.530 59.390 123.890 59.420 ;
        RECT 116.180 59.020 116.510 59.050 ;
        RECT 116.790 59.040 117.170 59.100 ;
        RECT 116.180 58.990 116.350 59.020 ;
        RECT 92.530 58.820 92.850 58.860 ;
        RECT 92.520 58.630 92.850 58.820 ;
        RECT 119.370 58.820 119.690 58.860 ;
        RECT 97.900 58.760 98.130 58.800 ;
        RECT 114.090 58.760 114.320 58.800 ;
        RECT 92.530 58.600 92.850 58.630 ;
        RECT 119.370 58.630 119.700 58.820 ;
        RECT 121.680 58.740 121.850 59.070 ;
        RECT 121.860 59.000 122.180 59.040 ;
        RECT 121.860 58.810 122.190 59.000 ;
        RECT 121.860 58.780 122.180 58.810 ;
        RECT 122.310 58.780 122.510 59.110 ;
        RECT 122.590 58.920 123.140 59.250 ;
        RECT 123.520 59.290 123.850 59.390 ;
        RECT 130.020 59.370 130.380 59.650 ;
        RECT 123.520 59.200 124.330 59.290 ;
        RECT 123.530 59.170 124.330 59.200 ;
        RECT 119.370 58.600 119.690 58.630 ;
        RECT 122.790 58.600 123.140 58.920 ;
        RECT 122.720 58.590 123.140 58.600 ;
        RECT 99.820 58.300 100.140 58.340 ;
        RECT 99.810 58.110 100.140 58.300 ;
        RECT 114.060 58.160 114.270 58.590 ;
        RECT 122.720 58.570 123.040 58.590 ;
        RECT 122.720 58.380 123.050 58.570 ;
        RECT 123.630 58.410 124.330 59.170 ;
        RECT 124.980 59.060 125.160 59.250 ;
        RECT 130.020 59.200 130.350 59.370 ;
        RECT 130.460 59.110 130.790 59.280 ;
        RECT 122.720 58.340 123.040 58.380 ;
        RECT 114.080 58.140 114.250 58.160 ;
        RECT 99.820 58.080 100.140 58.110 ;
        RECT 99.940 57.940 99.960 58.080 ;
        RECT 114.580 58.020 114.770 58.130 ;
        RECT 87.850 57.210 88.080 57.900 ;
        RECT 99.940 57.860 100.290 57.940 ;
        RECT 114.580 57.900 115.000 58.020 ;
        RECT 86.300 57.170 86.510 57.200 ;
        RECT 49.660 57.040 50.480 57.070 ;
        RECT 47.240 57.030 47.470 57.040 ;
        RECT 22.160 56.550 22.490 56.700 ;
        RECT 47.200 56.590 47.470 57.030 ;
        RECT 50.220 56.900 50.480 57.040 ;
        RECT 48.680 56.590 49.010 56.850 ;
        RECT 49.630 56.800 49.920 56.830 ;
        RECT 49.590 56.630 49.920 56.800 ;
        RECT 49.630 56.590 49.920 56.630 ;
        RECT 50.220 56.730 51.400 56.900 ;
        RECT 86.310 56.820 86.510 57.170 ;
        RECT 87.790 56.900 88.320 57.070 ;
        RECT 95.240 57.010 100.290 57.860 ;
        RECT 114.480 57.850 115.000 57.900 ;
        RECT 115.350 57.850 116.610 58.030 ;
        RECT 122.970 58.020 123.160 58.250 ;
        RECT 124.150 57.990 124.320 58.410 ;
        RECT 114.480 57.770 114.670 57.850 ;
        RECT 114.460 57.740 114.670 57.770 ;
        RECT 114.450 57.730 114.670 57.740 ;
        RECT 115.840 57.730 116.170 57.850 ;
        RECT 114.330 57.680 114.670 57.730 ;
        RECT 114.200 57.650 114.670 57.680 ;
        RECT 114.160 57.620 114.670 57.650 ;
        RECT 114.160 57.560 114.650 57.620 ;
        RECT 114.160 57.510 114.500 57.560 ;
        RECT 114.160 57.490 114.420 57.510 ;
        RECT 114.160 57.470 114.390 57.490 ;
        RECT 121.680 57.480 121.850 57.810 ;
        RECT 121.860 57.740 122.180 57.770 ;
        RECT 121.860 57.550 122.190 57.740 ;
        RECT 121.860 57.510 122.180 57.550 ;
        RECT 114.160 57.430 114.370 57.470 ;
        RECT 122.310 57.440 122.510 57.770 ;
        RECT 122.790 57.680 123.140 57.960 ;
        RECT 123.620 57.900 124.320 57.990 ;
        RECT 123.620 57.810 124.370 57.900 ;
        RECT 122.700 57.630 123.140 57.680 ;
        RECT 114.160 57.150 114.330 57.430 ;
        RECT 122.590 57.290 123.140 57.630 ;
        RECT 123.620 57.390 123.940 57.430 ;
        RECT 123.620 57.320 123.950 57.390 ;
        RECT 121.910 57.090 122.230 57.120 ;
        RECT 121.910 56.900 122.240 57.090 ;
        RECT 121.910 56.860 122.230 56.900 ;
        RECT 122.310 56.780 122.510 57.110 ;
        RECT 122.700 56.970 123.140 57.290 ;
        RECT 123.450 57.220 123.950 57.320 ;
        RECT 123.310 57.200 123.950 57.220 ;
        RECT 124.140 57.210 124.370 57.810 ;
        RECT 124.980 57.450 125.150 59.060 ;
        RECT 125.340 58.250 125.630 58.580 ;
        RECT 125.350 57.960 125.550 58.250 ;
        RECT 125.350 57.950 125.540 57.960 ;
        RECT 125.710 57.780 125.920 57.790 ;
        RECT 125.700 57.200 125.920 57.780 ;
        RECT 123.310 57.170 123.940 57.200 ;
        RECT 125.710 57.170 125.920 57.200 ;
        RECT 123.310 57.100 123.780 57.170 ;
        RECT 123.310 57.090 123.770 57.100 ;
        RECT 123.430 57.060 123.770 57.090 ;
        RECT 123.430 56.990 123.480 57.060 ;
        RECT 50.220 56.590 50.480 56.730 ;
        RECT 22.160 56.530 22.770 56.550 ;
        RECT 22.450 56.510 22.770 56.530 ;
        RECT 20.950 56.400 21.270 56.440 ;
        RECT 20.950 56.210 21.280 56.400 ;
        RECT 22.450 56.340 22.780 56.510 ;
        RECT 46.650 56.450 46.820 56.510 ;
        RECT 23.750 56.410 24.070 56.450 ;
        RECT 22.450 56.290 22.930 56.340 ;
        RECT 20.950 56.180 21.270 56.210 ;
        RECT 22.620 56.160 22.930 56.290 ;
        RECT 22.600 56.140 22.930 56.160 ;
        RECT 22.760 56.010 22.930 56.140 ;
        RECT 23.440 56.010 23.610 56.340 ;
        RECT 23.750 56.220 24.080 56.410 ;
        RECT 46.620 56.230 46.840 56.450 ;
        RECT 47.170 56.410 47.500 56.590 ;
        RECT 47.750 56.420 49.910 56.590 ;
        RECT 50.150 56.420 50.480 56.590 ;
        RECT 50.620 56.580 51.400 56.730 ;
        RECT 50.250 56.370 50.480 56.420 ;
        RECT 23.750 56.190 24.070 56.220 ;
        RECT 46.650 56.180 46.820 56.230 ;
        RECT 50.250 56.140 50.420 56.370 ;
        RECT 50.770 56.230 50.980 56.560 ;
        RECT 51.220 56.290 51.400 56.580 ;
        RECT 51.680 56.570 52.010 56.740 ;
        RECT 50.040 56.130 50.420 56.140 ;
        RECT 50.040 56.070 50.510 56.130 ;
        RECT 51.760 56.110 51.940 56.570 ;
        RECT 51.950 56.390 52.570 56.560 ;
        RECT 114.040 56.460 114.680 56.640 ;
        RECT 115.060 56.470 115.410 56.640 ;
        RECT 115.510 56.630 115.700 56.740 ;
        RECT 121.910 56.650 122.230 56.690 ;
        RECT 115.510 56.510 115.840 56.630 ;
        RECT 115.590 56.430 115.840 56.510 ;
        RECT 116.140 56.460 117.280 56.640 ;
        RECT 121.910 56.460 122.240 56.650 ;
        RECT 121.910 56.430 122.230 56.460 ;
        RECT 122.310 56.440 122.510 56.770 ;
        RECT 122.700 56.620 122.880 56.970 ;
        RECT 122.900 56.780 123.100 56.970 ;
        RECT 122.900 56.580 123.100 56.770 ;
        RECT 123.350 56.660 123.520 56.990 ;
        RECT 123.900 56.900 124.430 57.070 ;
        RECT 125.710 56.820 125.910 57.170 ;
        RECT 123.610 56.670 123.930 56.710 ;
        RECT 123.610 56.580 123.940 56.670 ;
        RECT 49.700 56.020 50.510 56.070 ;
        RECT 49.690 55.960 50.510 56.020 ;
        RECT 49.690 55.900 50.430 55.960 ;
        RECT 50.980 55.940 51.940 56.110 ;
        RECT 50.040 55.850 50.430 55.900 ;
        RECT 22.380 55.810 22.810 55.830 ;
        RECT 22.360 55.640 22.810 55.810 ;
        RECT 22.380 55.620 22.810 55.640 ;
        RECT 22.450 55.520 22.770 55.560 ;
        RECT 22.450 55.350 22.780 55.520 ;
        RECT 23.750 55.420 24.070 55.460 ;
        RECT 22.450 55.300 22.930 55.350 ;
        RECT 22.620 55.170 22.930 55.300 ;
        RECT 22.600 55.150 22.930 55.170 ;
        RECT 22.760 55.020 22.930 55.150 ;
        RECT 23.440 55.020 23.610 55.350 ;
        RECT 23.750 55.230 24.080 55.420 ;
        RECT 23.750 55.200 24.070 55.230 ;
        RECT 103.120 55.090 103.320 56.100 ;
        RECT 108.870 55.090 109.160 56.100 ;
        RECT 114.440 56.080 114.610 56.090 ;
        RECT 114.160 55.800 114.330 56.080 ;
        RECT 114.440 56.040 114.840 56.080 ;
        RECT 114.440 55.850 114.850 56.040 ;
        RECT 115.050 56.010 115.240 56.120 ;
        RECT 115.050 55.890 115.390 56.010 ;
        RECT 114.440 55.820 114.840 55.850 ;
        RECT 115.100 55.840 115.390 55.890 ;
        RECT 114.160 55.760 114.370 55.800 ;
        RECT 114.440 55.790 114.610 55.820 ;
        RECT 114.160 55.740 114.390 55.760 ;
        RECT 115.670 55.750 115.840 56.430 ;
        RECT 122.590 56.250 122.780 56.260 ;
        RECT 122.790 56.250 123.140 56.580 ;
        RECT 123.610 56.450 124.080 56.580 ;
        RECT 123.750 56.370 124.080 56.450 ;
        RECT 123.890 56.350 124.080 56.370 ;
        RECT 116.180 56.080 116.350 56.090 ;
        RECT 116.180 56.040 116.510 56.080 ;
        RECT 116.180 55.850 116.520 56.040 ;
        RECT 117.160 56.020 117.350 56.130 ;
        RECT 117.040 56.010 117.350 56.020 ;
        RECT 116.790 55.900 117.350 56.010 ;
        RECT 116.180 55.820 116.510 55.850 ;
        RECT 116.790 55.840 117.170 55.900 ;
        RECT 116.180 55.790 116.350 55.820 ;
        RECT 121.680 55.740 121.850 56.070 ;
        RECT 121.860 56.000 122.180 56.040 ;
        RECT 121.860 55.810 122.190 56.000 ;
        RECT 121.860 55.780 122.180 55.810 ;
        RECT 122.310 55.780 122.510 56.110 ;
        RECT 122.590 55.920 123.140 56.250 ;
        RECT 114.160 55.720 114.420 55.740 ;
        RECT 114.160 55.670 114.500 55.720 ;
        RECT 114.160 55.610 114.650 55.670 ;
        RECT 122.790 55.660 123.140 55.920 ;
        RECT 114.160 55.580 114.670 55.610 ;
        RECT 122.790 55.590 123.160 55.660 ;
        RECT 114.200 55.550 114.670 55.580 ;
        RECT 114.330 55.500 114.670 55.550 ;
        RECT 114.450 55.490 114.670 55.500 ;
        RECT 114.460 55.460 114.670 55.490 ;
        RECT 22.380 54.820 22.810 54.840 ;
        RECT 22.360 54.650 22.810 54.820 ;
        RECT 22.380 54.630 22.810 54.650 ;
        RECT 114.060 54.640 114.270 55.390 ;
        RECT 114.480 55.380 114.670 55.460 ;
        RECT 115.840 55.380 116.170 55.500 ;
        RECT 122.970 55.430 123.160 55.590 ;
        RECT 123.620 55.530 124.320 55.710 ;
        RECT 114.480 55.330 115.000 55.380 ;
        RECT 114.580 55.210 115.000 55.330 ;
        RECT 114.580 55.100 114.770 55.210 ;
        RECT 115.350 55.200 116.610 55.380 ;
        RECT 114.580 54.820 114.770 54.930 ;
        RECT 114.580 54.700 115.000 54.820 ;
        RECT 114.480 54.650 115.000 54.700 ;
        RECT 115.350 54.650 116.610 54.830 ;
        RECT 114.480 54.570 114.670 54.650 ;
        RECT 22.450 54.530 22.770 54.570 ;
        RECT 114.460 54.540 114.670 54.570 ;
        RECT 114.450 54.530 114.670 54.540 ;
        RECT 115.840 54.530 116.170 54.650 ;
        RECT 22.450 54.360 22.780 54.530 ;
        RECT 114.330 54.480 114.670 54.530 ;
        RECT 121.680 54.480 121.850 54.810 ;
        RECT 121.860 54.740 122.180 54.770 ;
        RECT 121.860 54.550 122.190 54.740 ;
        RECT 121.860 54.510 122.180 54.550 ;
        RECT 23.750 54.430 24.070 54.470 ;
        RECT 114.200 54.450 114.670 54.480 ;
        RECT 22.450 54.310 22.930 54.360 ;
        RECT 22.620 54.180 22.930 54.310 ;
        RECT 22.600 54.170 22.930 54.180 ;
        RECT 22.600 54.160 23.090 54.170 ;
        RECT 22.760 54.080 23.090 54.160 ;
        RECT 22.760 54.000 23.150 54.080 ;
        RECT 23.440 54.030 23.610 54.360 ;
        RECT 23.750 54.240 24.080 54.430 ;
        RECT 114.160 54.420 114.670 54.450 ;
        RECT 122.310 54.440 122.510 54.770 ;
        RECT 122.790 54.630 123.140 54.960 ;
        RECT 114.160 54.360 114.650 54.420 ;
        RECT 114.160 54.310 114.500 54.360 ;
        RECT 114.160 54.290 114.420 54.310 ;
        RECT 122.590 54.300 123.140 54.630 ;
        RECT 123.630 54.460 124.330 55.110 ;
        RECT 122.590 54.290 122.780 54.300 ;
        RECT 114.160 54.270 114.390 54.290 ;
        RECT 23.750 54.210 24.070 54.240 ;
        RECT 114.160 54.230 114.370 54.270 ;
        RECT 22.920 53.890 23.150 54.000 ;
        RECT 114.160 53.950 114.330 54.230 ;
        RECT 114.440 54.210 114.610 54.240 ;
        RECT 114.440 54.180 114.840 54.210 ;
        RECT 114.440 53.990 114.850 54.180 ;
        RECT 115.100 54.140 115.390 54.190 ;
        RECT 115.050 54.020 115.390 54.140 ;
        RECT 114.440 53.950 114.840 53.990 ;
        RECT 114.440 53.940 114.610 53.950 ;
        RECT 115.050 53.910 115.240 54.020 ;
        RECT 22.380 53.830 22.810 53.850 ;
        RECT 22.360 53.660 22.810 53.830 ;
        RECT 22.380 53.640 22.810 53.660 ;
        RECT 115.670 53.600 115.840 54.280 ;
        RECT 116.180 54.210 116.350 54.240 ;
        RECT 116.180 54.180 116.510 54.210 ;
        RECT 117.340 54.190 117.660 54.230 ;
        RECT 116.180 53.990 116.520 54.180 ;
        RECT 116.790 54.130 117.170 54.190 ;
        RECT 117.330 54.130 117.660 54.190 ;
        RECT 116.790 54.020 117.660 54.130 ;
        RECT 117.040 54.010 117.660 54.020 ;
        RECT 116.180 53.950 116.510 53.990 ;
        RECT 117.160 53.970 117.660 54.010 ;
        RECT 121.910 54.090 122.230 54.120 ;
        RECT 116.180 53.940 116.350 53.950 ;
        RECT 117.160 53.900 117.500 53.970 ;
        RECT 117.330 53.660 117.500 53.900 ;
        RECT 121.910 53.900 122.240 54.090 ;
        RECT 121.910 53.860 122.230 53.900 ;
        RECT 122.310 53.780 122.510 54.110 ;
        RECT 122.790 53.970 123.140 54.300 ;
        RECT 123.530 54.230 124.330 54.460 ;
        RECT 123.530 54.200 123.850 54.230 ;
        RECT 122.900 53.780 123.100 53.970 ;
        RECT 123.630 53.620 124.340 53.790 ;
        RECT 114.040 53.390 114.680 53.570 ;
        RECT 115.060 53.390 115.410 53.560 ;
        RECT 115.590 53.520 115.840 53.600 ;
        RECT 115.510 53.400 115.840 53.520 ;
        RECT 115.510 53.290 115.700 53.400 ;
        RECT 116.140 53.390 117.280 53.570 ;
        RECT 117.490 53.360 117.810 53.400 ;
        RECT 61.630 52.830 61.800 53.250 ;
        RECT 62.440 53.130 62.680 53.160 ;
        RECT 62.110 52.960 62.680 53.130 ;
        RECT 62.920 52.960 64.260 53.130 ;
        RECT 64.710 52.960 65.670 53.130 ;
        RECT 62.440 52.920 62.680 52.960 ;
        RECT 65.220 52.950 65.390 52.960 ;
        RECT 61.560 52.610 61.730 52.650 ;
        RECT 61.500 52.440 61.730 52.610 ;
        RECT 64.850 52.510 65.190 52.690 ;
        RECT 61.560 52.230 61.730 52.440 ;
        RECT 61.500 52.060 61.730 52.230 ;
        RECT 61.800 52.220 61.990 52.450 ;
        RECT 62.090 52.340 62.460 52.510 ;
        RECT 62.920 52.340 65.670 52.510 ;
        RECT 62.090 52.160 62.460 52.330 ;
        RECT 62.920 52.160 65.670 52.330 ;
        RECT 50.040 52.010 50.430 52.060 ;
        RECT 61.560 52.020 61.730 52.060 ;
        RECT 49.690 51.950 50.430 52.010 ;
        RECT 64.850 51.980 65.190 52.160 ;
        RECT 49.690 51.890 50.510 51.950 ;
        RECT 49.700 51.840 50.510 51.890 ;
        RECT 50.040 51.780 50.510 51.840 ;
        RECT 50.980 51.800 51.940 51.970 ;
        RECT 50.040 51.770 50.420 51.780 ;
        RECT 46.650 51.680 46.820 51.730 ;
        RECT 46.620 51.460 46.840 51.680 ;
        RECT 50.250 51.540 50.420 51.770 ;
        RECT 46.650 51.400 46.820 51.460 ;
        RECT 47.170 51.320 47.500 51.500 ;
        RECT 50.250 51.490 50.480 51.540 ;
        RECT 47.750 51.320 49.910 51.490 ;
        RECT 50.150 51.320 50.480 51.490 ;
        RECT 50.770 51.350 50.980 51.680 ;
        RECT 51.220 51.330 51.400 51.620 ;
        RECT 51.760 51.340 51.940 51.800 ;
        RECT 51.950 51.350 52.570 51.520 ;
        RECT 61.630 51.420 61.800 51.840 ;
        RECT 62.440 51.710 62.680 51.750 ;
        RECT 65.220 51.710 65.390 51.720 ;
        RECT 62.110 51.540 62.680 51.710 ;
        RECT 62.920 51.540 64.260 51.710 ;
        RECT 64.710 51.540 65.670 51.710 ;
        RECT 62.440 51.510 62.680 51.540 ;
        RECT 66.200 51.470 66.370 53.200 ;
        RECT 66.600 52.360 66.770 53.250 ;
        RECT 117.480 53.170 117.810 53.360 ;
        RECT 123.980 53.340 124.340 53.620 ;
        RECT 123.980 53.170 124.310 53.340 ;
        RECT 117.490 53.140 117.810 53.170 ;
        RECT 124.420 53.080 124.750 53.250 ;
        RECT 126.330 53.190 126.510 55.240 ;
        RECT 127.060 54.980 127.390 55.150 ;
        RECT 127.140 53.200 127.310 54.980 ;
        RECT 114.160 52.600 114.330 52.880 ;
        RECT 114.160 52.560 114.370 52.600 ;
        RECT 114.160 52.540 114.390 52.560 ;
        RECT 116.680 52.540 117.000 52.570 ;
        RECT 114.160 52.520 114.420 52.540 ;
        RECT 114.160 52.470 114.500 52.520 ;
        RECT 114.160 52.410 114.650 52.470 ;
        RECT 114.160 52.380 114.670 52.410 ;
        RECT 114.200 52.350 114.670 52.380 ;
        RECT 66.600 51.420 66.770 52.310 ;
        RECT 114.330 52.300 114.670 52.350 ;
        RECT 116.680 52.350 117.010 52.540 ;
        RECT 116.680 52.310 117.000 52.350 ;
        RECT 114.450 52.290 114.670 52.300 ;
        RECT 114.460 52.260 114.670 52.290 ;
        RECT 114.480 52.180 114.670 52.260 ;
        RECT 115.840 52.180 116.170 52.300 ;
        RECT 114.480 52.130 115.000 52.180 ;
        RECT 114.580 52.010 115.000 52.130 ;
        RECT 114.580 51.900 114.770 52.010 ;
        RECT 115.350 52.000 116.610 52.180 ;
        RECT 114.080 51.870 114.250 51.890 ;
        RECT 114.060 51.440 114.270 51.870 ;
        RECT 47.200 50.880 47.470 51.320 ;
        RECT 48.680 51.060 49.010 51.320 ;
        RECT 49.630 51.280 49.920 51.320 ;
        RECT 49.590 51.110 49.920 51.280 ;
        RECT 49.630 51.080 49.920 51.110 ;
        RECT 50.220 51.180 50.480 51.320 ;
        RECT 50.620 51.180 51.400 51.330 ;
        RECT 47.240 50.870 47.470 50.880 ;
        RECT 50.220 51.010 51.400 51.180 ;
        RECT 51.680 51.170 52.010 51.340 ;
        RECT 114.440 51.010 114.610 51.040 ;
        RECT 50.220 50.870 50.480 51.010 ;
        RECT 47.240 50.700 48.000 50.870 ;
        RECT 48.250 50.700 49.420 50.870 ;
        RECT 49.660 50.840 50.480 50.870 ;
        RECT 114.440 50.980 114.840 51.010 ;
        RECT 49.660 50.700 50.770 50.840 ;
        RECT 48.650 50.600 49.000 50.700 ;
        RECT 50.310 50.670 50.770 50.700 ;
        RECT 51.220 50.670 52.410 50.840 ;
        RECT 114.440 50.790 114.850 50.980 ;
        RECT 115.100 50.940 115.390 50.990 ;
        RECT 115.050 50.820 115.390 50.940 ;
        RECT 114.440 50.750 114.840 50.790 ;
        RECT 114.440 50.740 114.610 50.750 ;
        RECT 115.050 50.710 115.240 50.820 ;
        RECT 51.260 50.650 52.410 50.670 ;
        RECT 52.240 50.610 52.410 50.650 ;
        RECT 115.670 50.400 115.840 51.080 ;
        RECT 116.180 51.010 116.350 51.040 ;
        RECT 116.180 50.980 116.510 51.010 ;
        RECT 116.660 50.990 116.840 51.650 ;
        RECT 117.410 51.260 117.730 51.290 ;
        RECT 117.410 51.190 117.740 51.260 ;
        RECT 117.270 51.070 117.740 51.190 ;
        RECT 117.270 51.060 117.730 51.070 ;
        RECT 117.390 51.030 117.730 51.060 ;
        RECT 116.180 50.790 116.520 50.980 ;
        RECT 116.660 50.930 117.170 50.990 ;
        RECT 117.390 50.960 117.440 51.030 ;
        RECT 117.310 50.930 117.480 50.960 ;
        RECT 116.660 50.820 117.480 50.930 ;
        RECT 116.180 50.750 116.510 50.790 ;
        RECT 116.180 50.740 116.350 50.750 ;
        RECT 116.660 50.590 116.840 50.820 ;
        RECT 117.040 50.810 117.480 50.820 ;
        RECT 117.160 50.700 117.480 50.810 ;
        RECT 117.310 50.630 117.480 50.700 ;
        RECT 50.040 50.260 50.430 50.310 ;
        RECT 49.690 50.200 50.430 50.260 ;
        RECT 49.690 50.140 50.510 50.200 ;
        RECT 49.700 50.090 50.510 50.140 ;
        RECT 50.040 50.030 50.510 50.090 ;
        RECT 50.980 50.050 51.940 50.220 ;
        RECT 114.040 50.190 114.680 50.370 ;
        RECT 115.060 50.190 115.410 50.360 ;
        RECT 115.590 50.320 115.840 50.400 ;
        RECT 117.710 50.430 117.790 50.510 ;
        RECT 117.850 50.430 118.040 50.550 ;
        RECT 115.510 50.200 115.840 50.320 ;
        RECT 115.510 50.090 115.700 50.200 ;
        RECT 116.140 50.190 117.280 50.370 ;
        RECT 117.710 50.340 118.040 50.430 ;
        RECT 117.850 50.320 118.040 50.340 ;
        RECT 126.330 50.140 126.510 52.190 ;
        RECT 127.060 51.930 127.390 52.100 ;
        RECT 127.140 50.150 127.310 51.930 ;
        RECT 50.040 50.020 50.420 50.030 ;
        RECT 46.650 49.930 46.820 49.980 ;
        RECT 46.620 49.710 46.840 49.930 ;
        RECT 50.250 49.790 50.420 50.020 ;
        RECT 46.650 49.650 46.820 49.710 ;
        RECT 47.170 49.570 47.500 49.750 ;
        RECT 50.250 49.740 50.480 49.790 ;
        RECT 47.750 49.570 49.910 49.740 ;
        RECT 50.150 49.570 50.480 49.740 ;
        RECT 50.770 49.600 50.980 49.930 ;
        RECT 51.220 49.580 51.400 49.870 ;
        RECT 51.760 49.590 51.940 50.050 ;
        RECT 51.950 49.600 52.570 49.770 ;
        RECT 61.630 49.630 61.800 50.050 ;
        RECT 62.440 49.930 62.680 49.960 ;
        RECT 62.110 49.760 62.680 49.930 ;
        RECT 62.920 49.760 64.260 49.930 ;
        RECT 64.710 49.760 65.670 49.930 ;
        RECT 62.440 49.720 62.680 49.760 ;
        RECT 65.220 49.750 65.390 49.760 ;
        RECT 47.200 49.130 47.470 49.570 ;
        RECT 48.680 49.310 49.010 49.570 ;
        RECT 49.630 49.530 49.920 49.570 ;
        RECT 49.590 49.360 49.920 49.530 ;
        RECT 49.630 49.330 49.920 49.360 ;
        RECT 50.220 49.430 50.480 49.570 ;
        RECT 50.620 49.430 51.400 49.580 ;
        RECT 47.240 49.120 47.470 49.130 ;
        RECT 50.220 49.260 51.400 49.430 ;
        RECT 51.680 49.420 52.010 49.590 ;
        RECT 61.560 49.410 61.730 49.450 ;
        RECT 50.220 49.120 50.480 49.260 ;
        RECT 61.500 49.240 61.730 49.410 ;
        RECT 64.850 49.310 65.190 49.490 ;
        RECT 47.240 48.950 48.000 49.120 ;
        RECT 48.250 48.950 49.420 49.120 ;
        RECT 49.660 49.090 50.480 49.120 ;
        RECT 49.660 48.950 50.770 49.090 ;
        RECT 48.650 48.850 49.000 48.950 ;
        RECT 50.310 48.920 50.770 48.950 ;
        RECT 51.220 48.920 52.410 49.090 ;
        RECT 61.560 49.030 61.730 49.240 ;
        RECT 51.260 48.900 52.410 48.920 ;
        RECT 52.240 48.860 52.410 48.900 ;
        RECT 61.500 48.860 61.730 49.030 ;
        RECT 61.800 49.020 61.990 49.250 ;
        RECT 62.090 49.140 62.460 49.310 ;
        RECT 62.920 49.140 65.670 49.310 ;
        RECT 62.090 48.960 62.460 49.130 ;
        RECT 62.920 48.960 65.670 49.130 ;
        RECT 61.560 48.820 61.730 48.860 ;
        RECT 64.850 48.780 65.190 48.960 ;
        RECT 50.040 48.510 50.430 48.560 ;
        RECT 49.690 48.450 50.430 48.510 ;
        RECT 49.690 48.390 50.510 48.450 ;
        RECT 49.700 48.340 50.510 48.390 ;
        RECT 50.040 48.280 50.510 48.340 ;
        RECT 50.980 48.300 51.940 48.470 ;
        RECT 50.040 48.270 50.420 48.280 ;
        RECT 46.650 48.180 46.820 48.230 ;
        RECT 46.620 47.960 46.840 48.180 ;
        RECT 50.250 48.040 50.420 48.270 ;
        RECT 46.650 47.900 46.820 47.960 ;
        RECT 47.170 47.820 47.500 48.000 ;
        RECT 50.250 47.990 50.480 48.040 ;
        RECT 47.750 47.820 49.910 47.990 ;
        RECT 50.150 47.820 50.480 47.990 ;
        RECT 50.770 47.850 50.980 48.180 ;
        RECT 51.220 47.830 51.400 48.120 ;
        RECT 51.760 47.840 51.940 48.300 ;
        RECT 61.630 48.220 61.800 48.640 ;
        RECT 62.440 48.510 62.680 48.550 ;
        RECT 65.220 48.510 65.390 48.520 ;
        RECT 62.110 48.340 62.680 48.510 ;
        RECT 62.920 48.340 64.260 48.510 ;
        RECT 64.710 48.340 65.670 48.510 ;
        RECT 62.440 48.310 62.680 48.340 ;
        RECT 66.200 48.270 66.370 50.000 ;
        RECT 66.600 49.160 66.770 50.050 ;
        RECT 66.600 48.220 66.770 49.110 ;
        RECT 71.710 48.920 72.260 49.350 ;
        RECT 75.740 48.990 76.290 49.420 ;
        RECT 111.330 48.990 111.880 49.420 ;
        RECT 115.360 48.920 115.910 49.350 ;
        RECT 80.230 48.120 80.550 48.160 ;
        RECT 51.950 47.850 52.570 48.020 ;
        RECT 47.200 47.380 47.470 47.820 ;
        RECT 48.680 47.560 49.010 47.820 ;
        RECT 49.630 47.780 49.920 47.820 ;
        RECT 49.590 47.610 49.920 47.780 ;
        RECT 49.630 47.580 49.920 47.610 ;
        RECT 50.220 47.680 50.480 47.820 ;
        RECT 50.620 47.680 51.400 47.830 ;
        RECT 47.240 47.370 47.470 47.380 ;
        RECT 50.220 47.510 51.400 47.680 ;
        RECT 51.680 47.670 52.010 47.840 ;
        RECT 78.630 47.730 78.830 48.080 ;
        RECT 80.220 48.000 80.550 48.120 ;
        RECT 80.110 47.900 80.550 48.000 ;
        RECT 107.070 48.120 107.390 48.160 ;
        RECT 107.070 48.000 107.400 48.120 ;
        RECT 107.070 47.900 107.510 48.000 ;
        RECT 80.110 47.830 80.450 47.900 ;
        RECT 107.170 47.830 107.510 47.900 ;
        RECT 78.620 47.700 78.830 47.730 ;
        RECT 108.790 47.730 108.990 48.080 ;
        RECT 50.220 47.370 50.480 47.510 ;
        RECT 47.240 47.200 48.000 47.370 ;
        RECT 48.250 47.200 49.420 47.370 ;
        RECT 49.660 47.340 50.480 47.370 ;
        RECT 49.660 47.200 50.770 47.340 ;
        RECT 48.650 47.100 49.000 47.200 ;
        RECT 50.310 47.170 50.770 47.200 ;
        RECT 51.220 47.170 52.410 47.340 ;
        RECT 51.260 47.150 52.410 47.170 ;
        RECT 52.240 47.110 52.410 47.150 ;
        RECT 78.620 47.110 78.840 47.700 ;
        RECT 79.360 47.110 79.560 47.710 ;
        RECT 80.230 47.570 80.550 47.610 ;
        RECT 80.220 47.380 80.550 47.570 ;
        RECT 80.110 47.350 80.550 47.380 ;
        RECT 107.070 47.570 107.390 47.610 ;
        RECT 107.070 47.380 107.400 47.570 ;
        RECT 107.070 47.350 107.510 47.380 ;
        RECT 80.110 47.210 80.450 47.350 ;
        RECT 107.170 47.210 107.510 47.350 ;
        RECT 108.060 47.110 108.260 47.710 ;
        RECT 108.790 47.700 109.000 47.730 ;
        RECT 108.780 47.110 109.000 47.700 ;
        RECT 120.290 47.160 120.470 49.210 ;
        RECT 121.020 48.950 121.350 49.120 ;
        RECT 121.100 47.170 121.270 48.950 ;
        RECT 50.040 46.760 50.430 46.810 ;
        RECT 49.690 46.700 50.430 46.760 ;
        RECT 49.690 46.640 50.510 46.700 ;
        RECT 49.700 46.590 50.510 46.640 ;
        RECT 50.040 46.530 50.510 46.590 ;
        RECT 50.980 46.550 51.940 46.720 ;
        RECT 50.040 46.520 50.420 46.530 ;
        RECT 46.650 46.430 46.820 46.480 ;
        RECT 46.620 46.210 46.840 46.430 ;
        RECT 50.250 46.290 50.420 46.520 ;
        RECT 46.650 46.150 46.820 46.210 ;
        RECT 47.170 46.070 47.500 46.250 ;
        RECT 50.250 46.240 50.480 46.290 ;
        RECT 47.750 46.070 49.910 46.240 ;
        RECT 50.150 46.070 50.480 46.240 ;
        RECT 50.770 46.100 50.980 46.430 ;
        RECT 51.220 46.080 51.400 46.370 ;
        RECT 51.760 46.090 51.940 46.550 ;
        RECT 51.950 46.100 52.570 46.270 ;
        RECT 47.200 45.630 47.470 46.070 ;
        RECT 48.680 45.810 49.010 46.070 ;
        RECT 49.630 46.030 49.920 46.070 ;
        RECT 49.590 45.860 49.920 46.030 ;
        RECT 49.630 45.830 49.920 45.860 ;
        RECT 50.220 45.930 50.480 46.070 ;
        RECT 50.620 45.930 51.400 46.080 ;
        RECT 47.240 45.620 47.470 45.630 ;
        RECT 50.220 45.760 51.400 45.930 ;
        RECT 51.680 45.920 52.010 46.090 ;
        RECT 84.260 46.070 84.430 46.600 ;
        RECT 88.200 46.080 88.370 46.610 ;
        RECT 99.250 46.080 99.420 46.610 ;
        RECT 103.190 46.070 103.360 46.600 ;
        RECT 50.220 45.620 50.480 45.760 ;
        RECT 47.240 45.450 48.000 45.620 ;
        RECT 48.250 45.450 49.420 45.620 ;
        RECT 49.660 45.590 50.480 45.620 ;
        RECT 49.660 45.450 50.770 45.590 ;
        RECT 48.650 45.350 49.000 45.450 ;
        RECT 50.310 45.420 50.770 45.450 ;
        RECT 51.220 45.420 52.410 45.590 ;
        RECT 51.260 45.400 52.410 45.420 ;
        RECT 52.240 45.360 52.410 45.400 ;
        RECT 78.620 45.150 78.840 45.740 ;
        RECT 78.620 45.120 78.830 45.150 ;
        RECT 79.360 45.140 79.560 45.740 ;
        RECT 80.110 45.500 80.450 45.640 ;
        RECT 107.170 45.500 107.510 45.640 ;
        RECT 80.110 45.470 80.550 45.500 ;
        RECT 80.220 45.280 80.550 45.470 ;
        RECT 107.070 45.470 107.510 45.500 ;
        RECT 80.230 45.240 80.550 45.280 ;
        RECT 78.630 44.490 78.830 45.120 ;
        RECT 80.110 44.950 80.450 45.020 ;
        RECT 80.110 44.850 80.550 44.950 ;
        RECT 80.220 44.760 80.550 44.850 ;
        RECT 80.110 44.660 80.550 44.760 ;
        RECT 81.890 44.720 82.330 44.890 ;
        RECT 80.110 44.590 80.450 44.660 ;
        RECT 78.620 44.460 78.830 44.490 ;
        RECT 78.620 43.870 78.840 44.460 ;
        RECT 79.360 43.870 79.560 44.470 ;
        RECT 80.230 44.330 80.550 44.370 ;
        RECT 80.220 44.140 80.550 44.330 ;
        RECT 84.260 44.230 84.430 45.240 ;
        RECT 88.190 44.370 88.360 45.380 ;
        RECT 99.260 44.370 99.430 45.380 ;
        RECT 107.070 45.280 107.400 45.470 ;
        RECT 107.070 45.240 107.390 45.280 ;
        RECT 103.190 44.230 103.360 45.240 ;
        RECT 108.060 45.140 108.260 45.740 ;
        RECT 108.780 45.150 109.000 45.740 ;
        RECT 108.790 45.120 109.000 45.150 ;
        RECT 107.170 44.950 107.510 45.020 ;
        RECT 105.290 44.720 105.730 44.890 ;
        RECT 107.070 44.850 107.510 44.950 ;
        RECT 107.070 44.760 107.400 44.850 ;
        RECT 107.070 44.660 107.510 44.760 ;
        RECT 107.170 44.590 107.510 44.660 ;
        RECT 108.790 44.490 108.990 45.120 ;
        RECT 107.070 44.330 107.390 44.370 ;
        RECT 80.110 44.110 80.550 44.140 ;
        RECT 107.070 44.140 107.400 44.330 ;
        RECT 107.070 44.110 107.510 44.140 ;
        RECT 80.110 43.970 80.450 44.110 ;
        RECT 107.170 43.970 107.510 44.110 ;
        RECT 108.060 43.870 108.260 44.470 ;
        RECT 108.790 44.460 109.000 44.490 ;
        RECT 108.780 43.870 109.000 44.460 ;
        RECT 120.290 44.110 120.470 46.160 ;
        RECT 121.020 45.900 121.350 46.070 ;
        RECT 121.100 44.120 121.270 45.900 ;
        RECT 61.610 42.360 61.780 42.780 ;
        RECT 62.420 42.660 62.660 42.690 ;
        RECT 62.090 42.490 62.660 42.660 ;
        RECT 62.900 42.490 64.240 42.660 ;
        RECT 64.690 42.490 65.650 42.660 ;
        RECT 62.420 42.450 62.660 42.490 ;
        RECT 65.200 42.480 65.370 42.490 ;
        RECT 61.540 42.140 61.710 42.180 ;
        RECT 61.480 41.970 61.710 42.140 ;
        RECT 64.830 42.040 65.170 42.220 ;
        RECT 50.040 41.880 50.430 41.930 ;
        RECT 49.690 41.820 50.430 41.880 ;
        RECT 49.690 41.760 50.510 41.820 ;
        RECT 49.700 41.710 50.510 41.760 ;
        RECT 50.040 41.650 50.510 41.710 ;
        RECT 50.980 41.670 51.940 41.840 ;
        RECT 61.540 41.760 61.710 41.970 ;
        RECT 50.040 41.640 50.420 41.650 ;
        RECT 46.650 41.550 46.820 41.600 ;
        RECT 46.620 41.330 46.840 41.550 ;
        RECT 50.250 41.410 50.420 41.640 ;
        RECT 46.650 41.270 46.820 41.330 ;
        RECT 47.170 41.190 47.500 41.370 ;
        RECT 50.250 41.360 50.480 41.410 ;
        RECT 47.750 41.190 49.910 41.360 ;
        RECT 50.150 41.190 50.480 41.360 ;
        RECT 50.770 41.220 50.980 41.550 ;
        RECT 51.220 41.200 51.400 41.490 ;
        RECT 51.760 41.210 51.940 41.670 ;
        RECT 61.480 41.590 61.710 41.760 ;
        RECT 61.780 41.750 61.970 41.980 ;
        RECT 62.070 41.870 62.440 42.040 ;
        RECT 62.900 41.870 65.650 42.040 ;
        RECT 62.070 41.690 62.440 41.860 ;
        RECT 62.900 41.690 65.650 41.860 ;
        RECT 61.540 41.550 61.710 41.590 ;
        RECT 64.830 41.510 65.170 41.690 ;
        RECT 51.950 41.220 52.570 41.390 ;
        RECT 47.200 40.750 47.470 41.190 ;
        RECT 48.680 40.930 49.010 41.190 ;
        RECT 49.630 41.150 49.920 41.190 ;
        RECT 49.590 40.980 49.920 41.150 ;
        RECT 49.630 40.950 49.920 40.980 ;
        RECT 50.220 41.050 50.480 41.190 ;
        RECT 50.620 41.050 51.400 41.200 ;
        RECT 47.240 40.740 47.470 40.750 ;
        RECT 50.220 40.880 51.400 41.050 ;
        RECT 51.680 41.040 52.010 41.210 ;
        RECT 61.610 40.950 61.780 41.370 ;
        RECT 62.420 41.240 62.660 41.280 ;
        RECT 65.200 41.240 65.370 41.250 ;
        RECT 62.090 41.070 62.660 41.240 ;
        RECT 62.900 41.070 64.240 41.240 ;
        RECT 64.690 41.070 65.650 41.240 ;
        RECT 62.420 41.040 62.660 41.070 ;
        RECT 66.180 41.000 66.350 42.730 ;
        RECT 66.580 41.890 66.750 42.780 ;
        RECT 78.620 41.920 78.840 42.510 ;
        RECT 78.620 41.890 78.830 41.920 ;
        RECT 79.360 41.910 79.560 42.510 ;
        RECT 80.110 42.270 80.450 42.410 ;
        RECT 107.170 42.270 107.510 42.410 ;
        RECT 80.110 42.240 80.550 42.270 ;
        RECT 80.220 42.050 80.550 42.240 ;
        RECT 80.230 42.010 80.550 42.050 ;
        RECT 107.070 42.240 107.510 42.270 ;
        RECT 107.070 42.050 107.400 42.240 ;
        RECT 107.070 42.010 107.390 42.050 ;
        RECT 108.060 41.910 108.260 42.510 ;
        RECT 108.780 41.920 109.000 42.510 ;
        RECT 66.580 40.950 66.750 41.840 ;
        RECT 78.630 41.540 78.830 41.890 ;
        RECT 108.790 41.890 109.000 41.920 ;
        RECT 80.110 41.720 80.450 41.790 ;
        RECT 107.170 41.720 107.510 41.790 ;
        RECT 80.110 41.620 80.550 41.720 ;
        RECT 80.220 41.500 80.550 41.620 ;
        RECT 80.230 41.460 80.550 41.500 ;
        RECT 107.070 41.620 107.510 41.720 ;
        RECT 107.070 41.500 107.400 41.620 ;
        RECT 108.790 41.540 108.990 41.890 ;
        RECT 107.070 41.460 107.390 41.500 ;
        RECT 50.220 40.740 50.480 40.880 ;
        RECT 47.240 40.570 48.000 40.740 ;
        RECT 48.250 40.570 49.420 40.740 ;
        RECT 49.660 40.710 50.480 40.740 ;
        RECT 49.660 40.570 50.770 40.710 ;
        RECT 48.650 40.470 49.000 40.570 ;
        RECT 50.310 40.540 50.770 40.570 ;
        RECT 51.220 40.540 52.410 40.710 ;
        RECT 51.260 40.520 52.410 40.540 ;
        RECT 52.240 40.480 52.410 40.520 ;
        RECT 50.040 40.130 50.430 40.180 ;
        RECT 49.690 40.070 50.430 40.130 ;
        RECT 49.690 40.010 50.510 40.070 ;
        RECT 49.700 39.960 50.510 40.010 ;
        RECT 50.040 39.900 50.510 39.960 ;
        RECT 50.980 39.920 51.940 40.090 ;
        RECT 72.310 40.040 72.860 40.470 ;
        RECT 76.340 40.110 76.890 40.540 ;
        RECT 50.040 39.890 50.420 39.900 ;
        RECT 46.650 39.800 46.820 39.850 ;
        RECT 46.620 39.580 46.840 39.800 ;
        RECT 50.250 39.660 50.420 39.890 ;
        RECT 46.650 39.520 46.820 39.580 ;
        RECT 47.170 39.440 47.500 39.620 ;
        RECT 50.250 39.610 50.480 39.660 ;
        RECT 47.750 39.440 49.910 39.610 ;
        RECT 50.150 39.440 50.480 39.610 ;
        RECT 50.770 39.470 50.980 39.800 ;
        RECT 51.220 39.450 51.400 39.740 ;
        RECT 51.760 39.460 51.940 39.920 ;
        RECT 51.950 39.470 52.570 39.640 ;
        RECT 47.200 39.000 47.470 39.440 ;
        RECT 48.680 39.180 49.010 39.440 ;
        RECT 49.630 39.400 49.920 39.440 ;
        RECT 49.590 39.230 49.920 39.400 ;
        RECT 49.630 39.200 49.920 39.230 ;
        RECT 50.220 39.300 50.480 39.440 ;
        RECT 50.620 39.300 51.400 39.450 ;
        RECT 47.240 38.990 47.470 39.000 ;
        RECT 50.220 39.130 51.400 39.300 ;
        RECT 51.680 39.290 52.010 39.460 ;
        RECT 61.610 39.160 61.780 39.580 ;
        RECT 62.420 39.460 62.660 39.490 ;
        RECT 62.090 39.290 62.660 39.460 ;
        RECT 62.900 39.290 64.240 39.460 ;
        RECT 64.690 39.290 65.650 39.460 ;
        RECT 62.420 39.250 62.660 39.290 ;
        RECT 65.200 39.280 65.370 39.290 ;
        RECT 50.220 38.990 50.480 39.130 ;
        RECT 47.240 38.820 48.000 38.990 ;
        RECT 48.250 38.820 49.420 38.990 ;
        RECT 49.660 38.960 50.480 38.990 ;
        RECT 49.660 38.820 50.770 38.960 ;
        RECT 48.650 38.720 49.000 38.820 ;
        RECT 50.310 38.790 50.770 38.820 ;
        RECT 51.220 38.790 52.410 38.960 ;
        RECT 61.540 38.940 61.710 38.980 ;
        RECT 51.260 38.770 52.410 38.790 ;
        RECT 61.480 38.770 61.710 38.940 ;
        RECT 64.830 38.840 65.170 39.020 ;
        RECT 52.240 38.730 52.410 38.770 ;
        RECT 61.540 38.560 61.710 38.770 ;
        RECT 50.040 38.380 50.430 38.430 ;
        RECT 61.480 38.390 61.710 38.560 ;
        RECT 61.780 38.550 61.970 38.780 ;
        RECT 62.070 38.670 62.440 38.840 ;
        RECT 62.900 38.670 65.650 38.840 ;
        RECT 62.070 38.490 62.440 38.660 ;
        RECT 62.900 38.490 65.650 38.660 ;
        RECT 49.690 38.320 50.430 38.380 ;
        RECT 61.540 38.350 61.710 38.390 ;
        RECT 49.690 38.260 50.510 38.320 ;
        RECT 49.700 38.210 50.510 38.260 ;
        RECT 50.040 38.150 50.510 38.210 ;
        RECT 50.980 38.170 51.940 38.340 ;
        RECT 64.830 38.310 65.170 38.490 ;
        RECT 50.040 38.140 50.420 38.150 ;
        RECT 46.650 38.050 46.820 38.100 ;
        RECT 46.620 37.830 46.840 38.050 ;
        RECT 50.250 37.910 50.420 38.140 ;
        RECT 46.650 37.770 46.820 37.830 ;
        RECT 47.170 37.690 47.500 37.870 ;
        RECT 50.250 37.860 50.480 37.910 ;
        RECT 47.750 37.690 49.910 37.860 ;
        RECT 50.150 37.690 50.480 37.860 ;
        RECT 50.770 37.720 50.980 38.050 ;
        RECT 51.220 37.700 51.400 37.990 ;
        RECT 51.760 37.710 51.940 38.170 ;
        RECT 51.950 37.720 52.570 37.890 ;
        RECT 61.610 37.750 61.780 38.170 ;
        RECT 62.420 38.040 62.660 38.080 ;
        RECT 65.200 38.040 65.370 38.050 ;
        RECT 62.090 37.870 62.660 38.040 ;
        RECT 62.900 37.870 64.240 38.040 ;
        RECT 64.690 37.870 65.650 38.040 ;
        RECT 62.420 37.840 62.660 37.870 ;
        RECT 66.180 37.800 66.350 39.530 ;
        RECT 66.580 38.690 66.750 39.580 ;
        RECT 80.830 39.280 81.150 39.320 ;
        RECT 79.230 38.890 79.430 39.240 ;
        RECT 80.820 39.160 81.150 39.280 ;
        RECT 80.710 39.060 81.150 39.160 ;
        RECT 80.710 38.990 81.050 39.060 ;
        RECT 79.220 38.860 79.430 38.890 ;
        RECT 66.580 37.750 66.750 38.640 ;
        RECT 79.220 38.270 79.440 38.860 ;
        RECT 79.960 38.270 80.160 38.870 ;
        RECT 80.830 38.730 81.150 38.770 ;
        RECT 80.820 38.540 81.150 38.730 ;
        RECT 80.710 38.510 81.150 38.540 ;
        RECT 80.710 38.370 81.050 38.510 ;
        RECT 47.200 37.250 47.470 37.690 ;
        RECT 48.680 37.430 49.010 37.690 ;
        RECT 49.630 37.650 49.920 37.690 ;
        RECT 49.590 37.480 49.920 37.650 ;
        RECT 49.630 37.450 49.920 37.480 ;
        RECT 50.220 37.550 50.480 37.690 ;
        RECT 50.620 37.550 51.400 37.700 ;
        RECT 47.240 37.240 47.470 37.250 ;
        RECT 50.220 37.380 51.400 37.550 ;
        RECT 51.680 37.540 52.010 37.710 ;
        RECT 50.220 37.240 50.480 37.380 ;
        RECT 47.240 37.070 48.000 37.240 ;
        RECT 48.250 37.070 49.420 37.240 ;
        RECT 49.660 37.210 50.480 37.240 ;
        RECT 49.660 37.070 50.770 37.210 ;
        RECT 48.650 36.970 49.000 37.070 ;
        RECT 50.310 37.040 50.770 37.070 ;
        RECT 51.220 37.040 52.410 37.210 ;
        RECT 84.990 37.170 85.160 37.700 ;
        RECT 89.010 37.200 89.180 37.730 ;
        RECT 51.260 37.020 52.410 37.040 ;
        RECT 52.240 36.980 52.410 37.020 ;
        RECT 50.040 36.630 50.430 36.680 ;
        RECT 49.690 36.570 50.430 36.630 ;
        RECT 49.690 36.510 50.510 36.570 ;
        RECT 49.700 36.460 50.510 36.510 ;
        RECT 50.040 36.400 50.510 36.460 ;
        RECT 50.980 36.420 51.940 36.590 ;
        RECT 50.040 36.390 50.420 36.400 ;
        RECT 46.650 36.300 46.820 36.350 ;
        RECT 46.620 36.080 46.840 36.300 ;
        RECT 50.250 36.160 50.420 36.390 ;
        RECT 46.650 36.020 46.820 36.080 ;
        RECT 47.170 35.940 47.500 36.120 ;
        RECT 50.250 36.110 50.480 36.160 ;
        RECT 47.750 35.940 49.910 36.110 ;
        RECT 50.150 35.940 50.480 36.110 ;
        RECT 50.770 35.970 50.980 36.300 ;
        RECT 51.220 35.950 51.400 36.240 ;
        RECT 51.760 35.960 51.940 36.420 ;
        RECT 79.220 36.330 79.440 36.920 ;
        RECT 79.220 36.300 79.430 36.330 ;
        RECT 79.960 36.320 80.160 36.920 ;
        RECT 80.710 36.680 81.050 36.820 ;
        RECT 80.710 36.650 81.150 36.680 ;
        RECT 80.820 36.460 81.150 36.650 ;
        RECT 80.830 36.420 81.150 36.460 ;
        RECT 51.950 35.970 52.570 36.140 ;
        RECT 47.200 35.500 47.470 35.940 ;
        RECT 48.680 35.680 49.010 35.940 ;
        RECT 49.630 35.900 49.920 35.940 ;
        RECT 49.590 35.730 49.920 35.900 ;
        RECT 49.630 35.700 49.920 35.730 ;
        RECT 50.220 35.800 50.480 35.940 ;
        RECT 50.620 35.800 51.400 35.950 ;
        RECT 47.240 35.490 47.470 35.500 ;
        RECT 50.220 35.630 51.400 35.800 ;
        RECT 51.680 35.790 52.010 35.960 ;
        RECT 79.230 35.650 79.430 36.300 ;
        RECT 80.710 36.130 81.050 36.200 ;
        RECT 80.710 36.030 81.150 36.130 ;
        RECT 80.820 35.920 81.150 36.030 ;
        RECT 80.710 35.820 81.150 35.920 ;
        RECT 82.490 35.900 82.930 36.070 ;
        RECT 80.710 35.750 81.050 35.820 ;
        RECT 50.220 35.490 50.480 35.630 ;
        RECT 47.240 35.320 48.000 35.490 ;
        RECT 48.250 35.320 49.420 35.490 ;
        RECT 49.660 35.460 50.480 35.490 ;
        RECT 79.220 35.620 79.430 35.650 ;
        RECT 49.660 35.320 50.770 35.460 ;
        RECT 48.650 35.220 49.000 35.320 ;
        RECT 50.310 35.290 50.770 35.320 ;
        RECT 51.220 35.290 52.410 35.460 ;
        RECT 51.260 35.270 52.410 35.290 ;
        RECT 52.240 35.230 52.410 35.270 ;
        RECT 79.220 35.030 79.440 35.620 ;
        RECT 79.960 35.030 80.160 35.630 ;
        RECT 80.830 35.490 81.150 35.530 ;
        RECT 80.820 35.300 81.150 35.490 ;
        RECT 84.980 35.310 85.150 36.500 ;
        RECT 80.710 35.270 81.150 35.300 ;
        RECT 89.000 35.270 89.170 36.440 ;
        RECT 80.710 35.130 81.050 35.270 ;
        RECT 26.940 33.250 27.260 33.280 ;
        RECT 27.590 33.250 27.910 33.280 ;
        RECT 26.940 33.060 27.270 33.250 ;
        RECT 27.590 33.060 27.920 33.250 ;
        RECT 61.640 33.090 61.810 33.510 ;
        RECT 62.450 33.390 62.690 33.420 ;
        RECT 62.120 33.220 62.690 33.390 ;
        RECT 62.930 33.220 64.270 33.390 ;
        RECT 64.720 33.220 65.680 33.390 ;
        RECT 62.450 33.180 62.690 33.220 ;
        RECT 65.230 33.210 65.400 33.220 ;
        RECT 25.850 32.840 26.020 33.040 ;
        RECT 26.400 32.840 26.570 33.040 ;
        RECT 26.940 33.020 27.260 33.060 ;
        RECT 27.590 33.020 27.910 33.060 ;
        RECT 25.720 32.810 26.040 32.840 ;
        RECT 26.400 32.810 26.740 32.840 ;
        RECT 25.720 32.620 26.050 32.810 ;
        RECT 26.400 32.620 26.750 32.810 ;
        RECT 25.720 32.580 26.040 32.620 ;
        RECT 26.400 32.580 26.740 32.620 ;
        RECT 25.100 31.010 25.270 31.030 ;
        RECT 25.080 30.890 25.290 31.010 ;
        RECT 25.080 30.580 25.480 30.890 ;
        RECT 25.850 30.640 26.020 32.580 ;
        RECT 26.400 30.640 26.570 32.580 ;
        RECT 27.040 30.640 27.210 33.020 ;
        RECT 27.590 31.020 27.760 33.020 ;
        RECT 61.570 32.870 61.740 32.910 ;
        RECT 50.000 32.820 50.390 32.870 ;
        RECT 49.650 32.760 50.390 32.820 ;
        RECT 49.650 32.700 50.470 32.760 ;
        RECT 49.660 32.650 50.470 32.700 ;
        RECT 50.000 32.590 50.470 32.650 ;
        RECT 50.940 32.610 51.900 32.780 ;
        RECT 61.510 32.700 61.740 32.870 ;
        RECT 64.860 32.770 65.200 32.950 ;
        RECT 50.000 32.580 50.380 32.590 ;
        RECT 28.020 31.720 28.190 32.570 ;
        RECT 46.610 32.490 46.780 32.540 ;
        RECT 46.580 32.270 46.800 32.490 ;
        RECT 50.210 32.350 50.380 32.580 ;
        RECT 46.610 32.210 46.780 32.270 ;
        RECT 47.130 32.130 47.460 32.310 ;
        RECT 50.210 32.300 50.440 32.350 ;
        RECT 47.710 32.130 49.870 32.300 ;
        RECT 50.110 32.130 50.440 32.300 ;
        RECT 50.730 32.160 50.940 32.490 ;
        RECT 51.180 32.140 51.360 32.430 ;
        RECT 51.720 32.150 51.900 32.610 ;
        RECT 61.570 32.490 61.740 32.700 ;
        RECT 51.910 32.160 52.530 32.330 ;
        RECT 61.510 32.320 61.740 32.490 ;
        RECT 61.810 32.480 62.000 32.710 ;
        RECT 62.100 32.600 62.470 32.770 ;
        RECT 62.930 32.600 65.680 32.770 ;
        RECT 62.100 32.420 62.470 32.590 ;
        RECT 62.930 32.420 65.680 32.590 ;
        RECT 61.570 32.280 61.740 32.320 ;
        RECT 64.860 32.240 65.200 32.420 ;
        RECT 47.160 31.690 47.430 32.130 ;
        RECT 48.640 31.870 48.970 32.130 ;
        RECT 49.590 32.090 49.880 32.130 ;
        RECT 49.550 31.920 49.880 32.090 ;
        RECT 49.590 31.890 49.880 31.920 ;
        RECT 50.180 31.990 50.440 32.130 ;
        RECT 50.580 31.990 51.360 32.140 ;
        RECT 47.200 31.680 47.430 31.690 ;
        RECT 50.180 31.820 51.360 31.990 ;
        RECT 51.640 31.980 51.970 32.150 ;
        RECT 50.180 31.680 50.440 31.820 ;
        RECT 61.640 31.680 61.810 32.100 ;
        RECT 62.450 31.970 62.690 32.010 ;
        RECT 65.230 31.970 65.400 31.980 ;
        RECT 62.120 31.800 62.690 31.970 ;
        RECT 62.930 31.800 64.270 31.970 ;
        RECT 64.720 31.800 65.680 31.970 ;
        RECT 62.450 31.770 62.690 31.800 ;
        RECT 66.210 31.730 66.380 33.460 ;
        RECT 66.610 32.620 66.780 33.510 ;
        RECT 79.220 33.080 79.440 33.670 ;
        RECT 79.220 33.050 79.430 33.080 ;
        RECT 79.960 33.070 80.160 33.670 ;
        RECT 96.830 33.630 97.040 33.650 ;
        RECT 80.710 33.430 81.050 33.570 ;
        RECT 96.810 33.460 97.480 33.630 ;
        RECT 80.710 33.400 81.150 33.430 ;
        RECT 80.820 33.210 81.150 33.400 ;
        RECT 80.830 33.170 81.150 33.210 ;
        RECT 96.040 33.340 96.360 33.380 ;
        RECT 96.040 33.250 96.370 33.340 ;
        RECT 96.810 33.250 97.060 33.460 ;
        RECT 96.040 33.230 97.540 33.250 ;
        RECT 96.040 33.130 97.620 33.230 ;
        RECT 95.890 33.080 97.620 33.130 ;
        RECT 79.230 32.700 79.430 33.050 ;
        RECT 80.710 32.880 81.050 32.950 ;
        RECT 95.890 32.910 96.560 33.080 ;
        RECT 96.730 33.060 97.060 33.080 ;
        RECT 97.280 33.060 97.620 33.080 ;
        RECT 80.710 32.780 81.150 32.880 ;
        RECT 95.890 32.870 96.210 32.910 ;
        RECT 80.820 32.660 81.150 32.780 ;
        RECT 80.830 32.620 81.150 32.660 ;
        RECT 95.890 32.660 96.210 32.700 ;
        RECT 96.220 32.660 96.560 32.910 ;
        RECT 96.810 32.890 96.980 33.060 ;
        RECT 97.370 32.890 97.540 33.060 ;
        RECT 96.730 32.680 97.060 32.890 ;
        RECT 97.280 32.680 97.620 32.890 ;
        RECT 66.610 31.680 66.780 32.570 ;
        RECT 95.890 32.490 96.560 32.660 ;
        RECT 96.810 32.510 96.980 32.680 ;
        RECT 97.370 32.510 97.540 32.680 ;
        RECT 96.730 32.490 97.060 32.510 ;
        RECT 97.280 32.490 97.620 32.510 ;
        RECT 95.890 32.440 97.620 32.490 ;
        RECT 96.040 32.340 97.620 32.440 ;
        RECT 96.040 32.320 97.540 32.340 ;
        RECT 96.040 32.230 96.370 32.320 ;
        RECT 96.040 32.190 96.360 32.230 ;
        RECT 96.810 32.110 97.060 32.320 ;
        RECT 97.940 32.260 98.450 33.310 ;
        RECT 96.810 31.940 97.480 32.110 ;
        RECT 96.830 31.920 97.040 31.940 ;
        RECT 47.200 31.510 47.960 31.680 ;
        RECT 48.210 31.510 49.380 31.680 ;
        RECT 49.620 31.650 50.440 31.680 ;
        RECT 49.620 31.510 50.730 31.650 ;
        RECT 48.610 31.410 48.960 31.510 ;
        RECT 50.270 31.480 50.730 31.510 ;
        RECT 51.180 31.480 52.370 31.650 ;
        RECT 51.220 31.460 52.370 31.480 ;
        RECT 52.200 31.420 52.370 31.460 ;
        RECT 50.000 31.070 50.390 31.120 ;
        RECT 27.590 31.000 28.080 31.020 ;
        RECT 49.650 31.010 50.390 31.070 ;
        RECT 27.590 30.830 28.100 31.000 ;
        RECT 49.650 30.950 50.470 31.010 ;
        RECT 49.660 30.900 50.470 30.950 ;
        RECT 50.000 30.840 50.470 30.900 ;
        RECT 50.940 30.860 51.900 31.030 ;
        RECT 96.830 30.860 97.040 30.880 ;
        RECT 50.000 30.830 50.380 30.840 ;
        RECT 27.590 30.810 28.080 30.830 ;
        RECT 27.590 30.640 27.760 30.810 ;
        RECT 46.610 30.740 46.780 30.790 ;
        RECT 25.270 30.460 25.480 30.580 ;
        RECT 46.580 30.520 46.800 30.740 ;
        RECT 50.210 30.600 50.380 30.830 ;
        RECT 27.660 30.460 28.090 30.480 ;
        RECT 46.610 30.460 46.780 30.520 ;
        RECT 25.290 30.440 25.460 30.460 ;
        RECT 27.660 30.290 28.110 30.460 ;
        RECT 47.130 30.380 47.460 30.560 ;
        RECT 50.210 30.550 50.440 30.600 ;
        RECT 47.710 30.380 49.870 30.550 ;
        RECT 50.110 30.380 50.440 30.550 ;
        RECT 50.730 30.410 50.940 30.740 ;
        RECT 51.180 30.390 51.360 30.680 ;
        RECT 51.720 30.400 51.900 30.860 ;
        RECT 96.810 30.690 97.480 30.860 ;
        RECT 51.910 30.410 52.530 30.580 ;
        RECT 96.040 30.570 96.360 30.610 ;
        RECT 96.040 30.480 96.370 30.570 ;
        RECT 96.810 30.480 97.060 30.690 ;
        RECT 96.040 30.460 97.540 30.480 ;
        RECT 27.660 30.270 28.090 30.290 ;
        RECT 22.670 28.490 23.180 28.670 ;
        RECT 22.610 28.460 23.180 28.490 ;
        RECT 22.600 28.270 23.180 28.460 ;
        RECT 22.610 28.230 23.180 28.270 ;
        RECT 19.300 28.020 19.620 28.050 ;
        RECT 20.400 28.030 20.720 28.060 ;
        RECT 21.490 28.030 21.810 28.060 ;
        RECT 19.290 27.960 19.620 28.020 ;
        RECT 20.390 27.960 20.720 28.030 ;
        RECT 17.860 25.560 18.030 27.960 ;
        RECT 18.410 25.560 18.580 27.960 ;
        RECT 18.960 25.560 19.130 27.960 ;
        RECT 19.290 27.830 19.680 27.960 ;
        RECT 19.300 27.790 19.680 27.830 ;
        RECT 19.510 25.490 19.680 27.790 ;
        RECT 20.060 27.380 20.230 27.960 ;
        RECT 20.390 27.840 20.780 27.960 ;
        RECT 21.480 27.840 21.810 28.030 ;
        RECT 22.670 28.020 23.180 28.230 ;
        RECT 22.620 27.990 23.180 28.020 ;
        RECT 20.400 27.800 20.780 27.840 ;
        RECT 21.490 27.800 21.810 27.840 ;
        RECT 22.610 27.800 23.190 27.990 ;
        RECT 19.850 27.350 20.230 27.380 ;
        RECT 19.840 27.160 20.230 27.350 ;
        RECT 19.850 27.120 20.230 27.160 ;
        RECT 20.060 26.010 20.230 27.120 ;
        RECT 19.850 25.980 20.230 26.010 ;
        RECT 19.840 25.790 20.230 25.980 ;
        RECT 19.850 25.750 20.230 25.790 ;
        RECT 20.060 25.490 20.230 25.750 ;
        RECT 20.610 25.490 20.780 27.800 ;
        RECT 22.620 27.760 23.190 27.800 ;
        RECT 22.680 27.660 23.190 27.760 ;
        RECT 24.270 27.720 24.440 30.210 ;
        RECT 24.820 27.720 24.990 30.220 ;
        RECT 25.450 27.720 25.620 30.210 ;
        RECT 26.000 28.960 26.170 30.220 ;
        RECT 47.160 29.940 47.430 30.380 ;
        RECT 48.640 30.120 48.970 30.380 ;
        RECT 49.590 30.340 49.880 30.380 ;
        RECT 49.550 30.170 49.880 30.340 ;
        RECT 49.590 30.140 49.880 30.170 ;
        RECT 50.180 30.240 50.440 30.380 ;
        RECT 50.580 30.240 51.360 30.390 ;
        RECT 47.200 29.930 47.430 29.940 ;
        RECT 50.180 30.070 51.360 30.240 ;
        RECT 51.640 30.230 51.970 30.400 ;
        RECT 96.040 30.360 97.620 30.460 ;
        RECT 95.890 30.310 97.620 30.360 ;
        RECT 50.180 29.930 50.440 30.070 ;
        RECT 28.010 29.170 28.180 29.840 ;
        RECT 47.200 29.760 47.960 29.930 ;
        RECT 48.210 29.760 49.380 29.930 ;
        RECT 49.620 29.900 50.440 29.930 ;
        RECT 49.620 29.760 50.730 29.900 ;
        RECT 48.610 29.660 48.960 29.760 ;
        RECT 50.270 29.730 50.730 29.760 ;
        RECT 51.180 29.730 52.370 29.900 ;
        RECT 61.640 29.890 61.810 30.310 ;
        RECT 62.450 30.190 62.690 30.220 ;
        RECT 62.120 30.020 62.690 30.190 ;
        RECT 62.930 30.020 64.270 30.190 ;
        RECT 64.720 30.020 65.680 30.190 ;
        RECT 62.450 29.980 62.690 30.020 ;
        RECT 65.230 30.010 65.400 30.020 ;
        RECT 51.220 29.710 52.370 29.730 ;
        RECT 52.200 29.670 52.370 29.710 ;
        RECT 61.570 29.670 61.740 29.710 ;
        RECT 61.510 29.500 61.740 29.670 ;
        RECT 64.860 29.570 65.200 29.750 ;
        RECT 50.000 29.320 50.390 29.370 ;
        RECT 49.650 29.260 50.390 29.320 ;
        RECT 61.570 29.290 61.740 29.500 ;
        RECT 49.650 29.200 50.470 29.260 ;
        RECT 49.660 29.150 50.470 29.200 ;
        RECT 50.000 29.090 50.470 29.150 ;
        RECT 50.940 29.110 51.900 29.280 ;
        RECT 61.510 29.120 61.740 29.290 ;
        RECT 61.810 29.280 62.000 29.510 ;
        RECT 62.100 29.400 62.470 29.570 ;
        RECT 62.930 29.400 65.680 29.570 ;
        RECT 62.100 29.220 62.470 29.390 ;
        RECT 62.930 29.220 65.680 29.390 ;
        RECT 50.000 29.080 50.380 29.090 ;
        RECT 46.610 28.990 46.780 29.040 ;
        RECT 25.750 28.700 26.170 28.960 ;
        RECT 26.000 27.720 26.170 28.700 ;
        RECT 26.440 28.920 26.760 28.950 ;
        RECT 26.440 28.730 26.770 28.920 ;
        RECT 46.580 28.770 46.800 28.990 ;
        RECT 50.210 28.850 50.380 29.080 ;
        RECT 26.440 28.690 26.760 28.730 ;
        RECT 46.610 28.710 46.780 28.770 ;
        RECT 47.130 28.630 47.460 28.810 ;
        RECT 50.210 28.800 50.440 28.850 ;
        RECT 47.710 28.630 49.870 28.800 ;
        RECT 50.110 28.630 50.440 28.800 ;
        RECT 50.730 28.660 50.940 28.990 ;
        RECT 51.180 28.640 51.360 28.930 ;
        RECT 51.720 28.650 51.900 29.110 ;
        RECT 61.570 29.080 61.740 29.120 ;
        RECT 64.860 29.040 65.200 29.220 ;
        RECT 51.910 28.660 52.530 28.830 ;
        RECT 47.160 28.190 47.430 28.630 ;
        RECT 48.640 28.370 48.970 28.630 ;
        RECT 49.590 28.590 49.880 28.630 ;
        RECT 49.550 28.420 49.880 28.590 ;
        RECT 49.590 28.390 49.880 28.420 ;
        RECT 50.180 28.490 50.440 28.630 ;
        RECT 50.580 28.490 51.360 28.640 ;
        RECT 47.200 28.180 47.430 28.190 ;
        RECT 50.180 28.320 51.360 28.490 ;
        RECT 51.640 28.480 51.970 28.650 ;
        RECT 61.640 28.480 61.810 28.900 ;
        RECT 62.450 28.770 62.690 28.810 ;
        RECT 65.230 28.770 65.400 28.780 ;
        RECT 62.120 28.600 62.690 28.770 ;
        RECT 62.930 28.600 64.270 28.770 ;
        RECT 64.720 28.600 65.680 28.770 ;
        RECT 62.450 28.570 62.690 28.600 ;
        RECT 66.210 28.530 66.380 30.260 ;
        RECT 66.610 29.420 66.780 30.310 ;
        RECT 95.890 30.140 96.560 30.310 ;
        RECT 96.730 30.290 97.060 30.310 ;
        RECT 97.280 30.290 97.620 30.310 ;
        RECT 95.890 30.100 96.210 30.140 ;
        RECT 95.890 29.890 96.210 29.930 ;
        RECT 96.220 29.890 96.560 30.140 ;
        RECT 96.810 30.120 96.980 30.290 ;
        RECT 97.370 30.120 97.540 30.290 ;
        RECT 96.730 29.910 97.060 30.120 ;
        RECT 97.280 29.910 97.620 30.120 ;
        RECT 83.910 29.760 84.230 29.800 ;
        RECT 83.910 29.590 84.240 29.760 ;
        RECT 95.890 29.720 96.560 29.890 ;
        RECT 96.810 29.740 96.980 29.910 ;
        RECT 97.370 29.740 97.540 29.910 ;
        RECT 96.730 29.720 97.060 29.740 ;
        RECT 97.280 29.720 97.620 29.740 ;
        RECT 95.890 29.670 97.620 29.720 ;
        RECT 83.820 29.570 84.240 29.590 ;
        RECT 96.040 29.570 97.620 29.670 ;
        RECT 83.820 29.540 84.230 29.570 ;
        RECT 96.040 29.550 97.540 29.570 ;
        RECT 66.610 28.480 66.780 29.370 ;
        RECT 83.820 28.840 84.000 29.540 ;
        RECT 96.040 29.460 96.370 29.550 ;
        RECT 96.040 29.420 96.360 29.460 ;
        RECT 96.810 29.340 97.060 29.550 ;
        RECT 97.940 29.490 98.450 30.540 ;
        RECT 96.810 29.170 97.480 29.340 ;
        RECT 96.830 29.150 97.040 29.170 ;
        RECT 83.820 28.800 84.280 28.840 ;
        RECT 83.820 28.670 84.290 28.800 ;
        RECT 83.960 28.610 84.290 28.670 ;
        RECT 83.960 28.580 84.280 28.610 ;
        RECT 50.180 28.180 50.440 28.320 ;
        RECT 26.920 28.150 27.240 28.180 ;
        RECT 26.920 27.960 27.250 28.150 ;
        RECT 27.630 28.090 27.950 28.120 ;
        RECT 26.920 27.920 27.240 27.960 ;
        RECT 27.630 27.900 27.960 28.090 ;
        RECT 47.200 28.010 47.960 28.180 ;
        RECT 48.210 28.010 49.380 28.180 ;
        RECT 49.620 28.150 50.440 28.180 ;
        RECT 49.620 28.010 50.730 28.150 ;
        RECT 48.610 27.910 48.960 28.010 ;
        RECT 50.270 27.980 50.730 28.010 ;
        RECT 51.180 27.980 52.370 28.150 ;
        RECT 51.220 27.960 52.370 27.980 ;
        RECT 52.200 27.920 52.370 27.960 ;
        RECT 27.630 27.860 27.950 27.900 ;
        RECT 50.000 27.570 50.390 27.620 ;
        RECT 49.650 27.510 50.390 27.570 ;
        RECT 20.950 27.350 21.270 27.380 ;
        RECT 22.050 27.350 22.370 27.380 ;
        RECT 20.940 27.160 21.270 27.350 ;
        RECT 22.040 27.160 22.370 27.350 ;
        RECT 20.950 27.120 21.270 27.160 ;
        RECT 22.050 27.120 22.370 27.160 ;
        RECT 22.970 26.250 23.140 27.470 ;
        RECT 49.650 27.450 50.470 27.510 ;
        RECT 49.660 27.400 50.470 27.450 ;
        RECT 50.000 27.340 50.470 27.400 ;
        RECT 50.940 27.360 51.900 27.530 ;
        RECT 50.000 27.330 50.380 27.340 ;
        RECT 46.610 27.240 46.780 27.290 ;
        RECT 46.580 27.020 46.800 27.240 ;
        RECT 50.210 27.100 50.380 27.330 ;
        RECT 46.610 26.960 46.780 27.020 ;
        RECT 47.130 26.880 47.460 27.060 ;
        RECT 50.210 27.050 50.440 27.100 ;
        RECT 47.710 26.880 49.870 27.050 ;
        RECT 50.110 26.880 50.440 27.050 ;
        RECT 50.730 26.910 50.940 27.240 ;
        RECT 51.180 26.890 51.360 27.180 ;
        RECT 51.720 26.900 51.900 27.360 ;
        RECT 51.910 26.910 52.530 27.080 ;
        RECT 47.160 26.440 47.430 26.880 ;
        RECT 48.640 26.620 48.970 26.880 ;
        RECT 49.590 26.840 49.880 26.880 ;
        RECT 49.550 26.670 49.880 26.840 ;
        RECT 49.590 26.640 49.880 26.670 ;
        RECT 50.180 26.740 50.440 26.880 ;
        RECT 50.580 26.740 51.360 26.890 ;
        RECT 47.200 26.430 47.430 26.440 ;
        RECT 50.180 26.570 51.360 26.740 ;
        RECT 51.640 26.730 51.970 26.900 ;
        RECT 50.180 26.430 50.440 26.570 ;
        RECT 47.200 26.260 47.960 26.430 ;
        RECT 48.210 26.260 49.380 26.430 ;
        RECT 49.620 26.400 50.440 26.430 ;
        RECT 49.620 26.260 50.730 26.400 ;
        RECT 48.610 26.160 48.960 26.260 ;
        RECT 50.270 26.230 50.730 26.260 ;
        RECT 51.180 26.230 52.370 26.400 ;
        RECT 51.220 26.210 52.370 26.230 ;
        RECT 52.200 26.170 52.370 26.210 ;
        RECT 20.950 25.980 21.270 26.010 ;
        RECT 22.050 25.980 22.370 26.010 ;
        RECT 20.940 25.870 21.270 25.980 ;
        RECT 22.040 25.870 22.370 25.980 ;
        RECT 20.940 25.790 21.330 25.870 ;
        RECT 20.950 25.750 21.330 25.790 ;
        RECT 21.160 25.490 21.330 25.750 ;
        RECT 21.710 25.490 21.880 25.870 ;
        RECT 22.040 25.790 22.430 25.870 ;
        RECT 22.050 25.750 22.430 25.790 ;
        RECT 22.260 25.490 22.430 25.750 ;
        RECT 19.300 25.250 19.620 25.280 ;
        RECT 20.400 25.250 20.720 25.280 ;
        RECT 21.490 25.250 21.810 25.280 ;
        RECT 19.290 25.180 19.620 25.250 ;
        RECT 20.390 25.180 20.720 25.250 ;
        RECT 17.860 22.780 18.030 25.180 ;
        RECT 18.410 22.780 18.580 25.180 ;
        RECT 18.960 22.780 19.130 25.180 ;
        RECT 19.290 25.060 19.680 25.180 ;
        RECT 19.300 25.020 19.680 25.060 ;
        RECT 19.510 23.940 19.680 25.020 ;
        RECT 19.290 23.910 19.680 23.940 ;
        RECT 19.280 23.720 19.680 23.910 ;
        RECT 19.290 23.680 19.680 23.720 ;
        RECT 19.510 22.780 19.680 23.680 ;
        RECT 20.060 23.240 20.230 25.180 ;
        RECT 20.390 25.060 20.780 25.180 ;
        RECT 21.480 25.060 21.810 25.250 ;
        RECT 20.400 25.020 20.780 25.060 ;
        RECT 21.490 25.020 21.810 25.060 ;
        RECT 20.610 23.930 20.780 25.020 ;
        RECT 29.300 23.970 30.060 24.390 ;
        RECT 20.400 23.900 20.780 23.930 ;
        RECT 20.390 23.710 20.780 23.900 ;
        RECT 21.490 23.880 21.810 23.910 ;
        RECT 20.400 23.670 20.780 23.710 ;
        RECT 21.480 23.690 21.810 23.880 ;
        RECT 19.850 23.210 20.230 23.240 ;
        RECT 19.840 23.020 20.230 23.210 ;
        RECT 19.850 22.980 20.230 23.020 ;
        RECT 20.060 22.780 20.230 22.980 ;
        RECT 20.610 22.780 20.780 23.670 ;
        RECT 21.490 23.650 21.810 23.690 ;
        RECT 20.950 23.200 21.270 23.230 ;
        RECT 22.040 23.200 22.360 23.230 ;
        RECT 20.940 23.010 21.270 23.200 ;
        RECT 22.030 23.010 22.360 23.200 ;
        RECT 29.320 23.180 30.060 23.970 ;
        RECT 20.950 22.970 21.270 23.010 ;
        RECT 22.040 22.970 22.360 23.010 ;
        RECT 62.370 22.110 62.540 22.140 ;
        RECT 52.560 22.080 52.730 22.110 ;
        RECT 52.560 22.040 52.880 22.080 ;
        RECT 52.560 21.850 52.890 22.040 ;
        RECT 52.560 21.820 52.880 21.850 ;
        RECT 22.710 20.930 23.220 21.110 ;
        RECT 22.650 20.900 23.220 20.930 ;
        RECT 22.640 20.710 23.220 20.900 ;
        RECT 19.480 20.490 19.650 20.710 ;
        RECT 19.340 20.460 19.660 20.490 ;
        RECT 19.330 20.270 19.660 20.460 ;
        RECT 19.340 20.230 19.660 20.270 ;
        RECT 19.480 18.310 19.650 20.230 ;
        RECT 20.030 19.820 20.200 20.710 ;
        RECT 20.580 20.500 20.750 20.710 ;
        RECT 20.440 20.470 20.760 20.500 ;
        RECT 20.430 20.280 20.760 20.470 ;
        RECT 20.440 20.240 20.760 20.280 ;
        RECT 19.890 19.790 20.210 19.820 ;
        RECT 19.880 19.600 20.210 19.790 ;
        RECT 19.890 19.560 20.210 19.600 ;
        RECT 20.030 18.450 20.200 19.560 ;
        RECT 19.890 18.420 20.210 18.450 ;
        RECT 19.880 18.310 20.210 18.420 ;
        RECT 20.580 18.310 20.750 20.240 ;
        RECT 21.130 19.820 21.300 20.710 ;
        RECT 21.680 20.500 21.850 20.710 ;
        RECT 21.530 20.470 21.850 20.500 ;
        RECT 21.520 20.280 21.850 20.470 ;
        RECT 21.530 20.240 21.850 20.280 ;
        RECT 20.990 19.790 21.310 19.820 ;
        RECT 20.980 19.600 21.310 19.790 ;
        RECT 20.990 19.560 21.310 19.600 ;
        RECT 21.130 18.450 21.300 19.560 ;
        RECT 20.990 18.420 21.310 18.450 ;
        RECT 20.980 18.310 21.310 18.420 ;
        RECT 21.680 18.310 21.850 20.240 ;
        RECT 22.230 19.820 22.400 20.700 ;
        RECT 22.650 20.670 23.220 20.710 ;
        RECT 22.710 20.460 23.220 20.670 ;
        RECT 22.660 20.430 23.220 20.460 ;
        RECT 22.650 20.240 23.230 20.430 ;
        RECT 22.660 20.200 23.230 20.240 ;
        RECT 22.710 20.180 23.230 20.200 ;
        RECT 22.720 20.100 23.230 20.180 ;
        RECT 22.090 19.790 22.410 19.820 ;
        RECT 22.080 19.600 22.410 19.790 ;
        RECT 52.560 19.620 52.730 21.820 ;
        RECT 53.110 21.400 53.280 22.110 ;
        RECT 53.660 22.080 53.830 22.110 ;
        RECT 53.650 22.040 53.970 22.080 ;
        RECT 53.650 21.850 53.980 22.040 ;
        RECT 53.650 21.820 53.970 21.850 ;
        RECT 53.110 21.360 53.430 21.400 ;
        RECT 53.110 21.170 53.440 21.360 ;
        RECT 53.110 21.140 53.430 21.170 ;
        RECT 53.110 20.030 53.280 21.140 ;
        RECT 53.110 19.990 53.430 20.030 ;
        RECT 53.110 19.800 53.440 19.990 ;
        RECT 53.110 19.770 53.430 19.800 ;
        RECT 53.110 19.610 53.280 19.770 ;
        RECT 53.660 19.610 53.830 21.820 ;
        RECT 54.210 21.380 54.380 22.110 ;
        RECT 54.760 22.070 54.930 22.110 ;
        RECT 54.750 22.030 55.070 22.070 ;
        RECT 54.750 21.840 55.080 22.030 ;
        RECT 54.750 21.810 55.070 21.840 ;
        RECT 54.200 21.340 54.520 21.380 ;
        RECT 54.200 21.150 54.530 21.340 ;
        RECT 54.200 21.120 54.520 21.150 ;
        RECT 54.210 20.030 54.380 21.120 ;
        RECT 54.200 19.990 54.520 20.030 ;
        RECT 54.200 19.800 54.530 19.990 ;
        RECT 54.200 19.770 54.520 19.800 ;
        RECT 54.210 19.610 54.380 19.770 ;
        RECT 54.760 19.610 54.930 21.810 ;
        RECT 55.310 21.370 55.480 22.110 ;
        RECT 55.310 21.330 55.630 21.370 ;
        RECT 55.310 21.140 55.640 21.330 ;
        RECT 55.790 21.290 55.960 22.050 ;
        RECT 57.680 21.290 57.850 22.050 ;
        RECT 58.160 21.370 58.330 22.110 ;
        RECT 58.710 22.070 58.880 22.110 ;
        RECT 58.570 22.030 58.890 22.070 ;
        RECT 58.560 21.840 58.890 22.030 ;
        RECT 58.570 21.810 58.890 21.840 ;
        RECT 58.010 21.330 58.330 21.370 ;
        RECT 58.000 21.140 58.330 21.330 ;
        RECT 55.310 21.110 55.630 21.140 ;
        RECT 58.010 21.110 58.330 21.140 ;
        RECT 55.310 20.030 55.480 21.110 ;
        RECT 58.160 20.030 58.330 21.110 ;
        RECT 55.300 19.990 55.620 20.030 ;
        RECT 58.020 19.990 58.340 20.030 ;
        RECT 55.300 19.800 55.630 19.990 ;
        RECT 58.010 19.800 58.340 19.990 ;
        RECT 55.300 19.770 55.620 19.800 ;
        RECT 58.020 19.770 58.340 19.800 ;
        RECT 55.310 19.610 55.480 19.770 ;
        RECT 58.160 19.610 58.330 19.770 ;
        RECT 58.710 19.610 58.880 21.810 ;
        RECT 59.260 21.380 59.430 22.110 ;
        RECT 59.810 22.080 59.980 22.110 ;
        RECT 59.670 22.040 59.990 22.080 ;
        RECT 59.660 21.850 59.990 22.040 ;
        RECT 59.670 21.820 59.990 21.850 ;
        RECT 59.120 21.340 59.440 21.380 ;
        RECT 59.110 21.150 59.440 21.340 ;
        RECT 59.120 21.120 59.440 21.150 ;
        RECT 59.260 20.030 59.430 21.120 ;
        RECT 59.120 19.990 59.440 20.030 ;
        RECT 59.110 19.800 59.440 19.990 ;
        RECT 59.120 19.770 59.440 19.800 ;
        RECT 59.260 19.610 59.430 19.770 ;
        RECT 59.810 19.610 59.980 21.820 ;
        RECT 60.360 21.400 60.530 22.110 ;
        RECT 60.910 22.080 61.080 22.110 ;
        RECT 60.760 22.040 61.080 22.080 ;
        RECT 60.750 21.850 61.080 22.040 ;
        RECT 60.760 21.820 61.080 21.850 ;
        RECT 60.210 21.360 60.530 21.400 ;
        RECT 60.200 21.170 60.530 21.360 ;
        RECT 60.210 21.140 60.530 21.170 ;
        RECT 60.360 20.030 60.530 21.140 ;
        RECT 60.210 19.990 60.530 20.030 ;
        RECT 60.200 19.800 60.530 19.990 ;
        RECT 60.210 19.770 60.530 19.800 ;
        RECT 60.360 19.610 60.530 19.770 ;
        RECT 60.910 19.620 61.080 21.820 ;
        RECT 62.370 22.070 62.690 22.110 ;
        RECT 62.370 21.880 62.700 22.070 ;
        RECT 62.370 21.850 62.690 21.880 ;
        RECT 62.370 19.650 62.540 21.850 ;
        RECT 62.920 21.430 63.090 22.140 ;
        RECT 63.470 22.110 63.640 22.140 ;
        RECT 63.460 22.070 63.780 22.110 ;
        RECT 63.460 21.880 63.790 22.070 ;
        RECT 63.460 21.850 63.780 21.880 ;
        RECT 62.920 21.390 63.240 21.430 ;
        RECT 62.920 21.200 63.250 21.390 ;
        RECT 62.920 21.170 63.240 21.200 ;
        RECT 62.920 20.060 63.090 21.170 ;
        RECT 62.920 20.020 63.240 20.060 ;
        RECT 62.920 19.830 63.250 20.020 ;
        RECT 62.920 19.800 63.240 19.830 ;
        RECT 62.920 19.640 63.090 19.800 ;
        RECT 63.470 19.640 63.640 21.850 ;
        RECT 64.020 21.410 64.190 22.140 ;
        RECT 64.570 22.100 64.740 22.140 ;
        RECT 64.560 22.060 64.880 22.100 ;
        RECT 64.560 21.870 64.890 22.060 ;
        RECT 64.560 21.840 64.880 21.870 ;
        RECT 64.010 21.370 64.330 21.410 ;
        RECT 64.010 21.180 64.340 21.370 ;
        RECT 64.010 21.150 64.330 21.180 ;
        RECT 64.020 20.060 64.190 21.150 ;
        RECT 64.010 20.020 64.330 20.060 ;
        RECT 64.010 19.830 64.340 20.020 ;
        RECT 64.010 19.800 64.330 19.830 ;
        RECT 64.020 19.640 64.190 19.800 ;
        RECT 64.570 19.640 64.740 21.840 ;
        RECT 65.120 21.400 65.290 22.140 ;
        RECT 65.120 21.360 65.440 21.400 ;
        RECT 65.120 21.170 65.450 21.360 ;
        RECT 65.600 21.320 65.770 22.080 ;
        RECT 67.490 21.320 67.660 22.080 ;
        RECT 67.970 21.400 68.140 22.140 ;
        RECT 68.520 22.100 68.690 22.140 ;
        RECT 68.380 22.060 68.700 22.100 ;
        RECT 68.370 21.870 68.700 22.060 ;
        RECT 68.380 21.840 68.700 21.870 ;
        RECT 67.820 21.360 68.140 21.400 ;
        RECT 67.810 21.170 68.140 21.360 ;
        RECT 65.120 21.140 65.440 21.170 ;
        RECT 67.820 21.140 68.140 21.170 ;
        RECT 65.120 20.060 65.290 21.140 ;
        RECT 67.970 20.060 68.140 21.140 ;
        RECT 65.110 20.020 65.430 20.060 ;
        RECT 67.830 20.020 68.150 20.060 ;
        RECT 65.110 19.830 65.440 20.020 ;
        RECT 67.820 19.830 68.150 20.020 ;
        RECT 65.110 19.800 65.430 19.830 ;
        RECT 67.830 19.800 68.150 19.830 ;
        RECT 65.120 19.640 65.290 19.800 ;
        RECT 67.970 19.640 68.140 19.800 ;
        RECT 68.520 19.640 68.690 21.840 ;
        RECT 69.070 21.410 69.240 22.140 ;
        RECT 69.620 22.110 69.790 22.140 ;
        RECT 69.480 22.070 69.800 22.110 ;
        RECT 69.470 21.880 69.800 22.070 ;
        RECT 69.480 21.850 69.800 21.880 ;
        RECT 68.930 21.370 69.250 21.410 ;
        RECT 68.920 21.180 69.250 21.370 ;
        RECT 68.930 21.150 69.250 21.180 ;
        RECT 69.070 20.060 69.240 21.150 ;
        RECT 68.930 20.020 69.250 20.060 ;
        RECT 68.920 19.830 69.250 20.020 ;
        RECT 68.930 19.800 69.250 19.830 ;
        RECT 69.070 19.640 69.240 19.800 ;
        RECT 69.620 19.640 69.790 21.850 ;
        RECT 70.170 21.430 70.340 22.140 ;
        RECT 70.720 22.110 70.890 22.140 ;
        RECT 70.570 22.070 70.890 22.110 ;
        RECT 70.560 21.880 70.890 22.070 ;
        RECT 70.570 21.850 70.890 21.880 ;
        RECT 70.020 21.390 70.340 21.430 ;
        RECT 70.010 21.200 70.340 21.390 ;
        RECT 70.020 21.170 70.340 21.200 ;
        RECT 70.170 20.060 70.340 21.170 ;
        RECT 70.020 20.020 70.340 20.060 ;
        RECT 70.010 19.830 70.340 20.020 ;
        RECT 70.020 19.800 70.340 19.830 ;
        RECT 70.170 19.640 70.340 19.800 ;
        RECT 70.720 19.650 70.890 21.850 ;
        RECT 72.130 19.880 72.300 22.280 ;
        RECT 72.680 19.880 72.850 22.280 ;
        RECT 73.230 19.880 73.400 22.280 ;
        RECT 73.780 21.380 73.950 22.280 ;
        RECT 74.330 22.080 74.500 22.280 ;
        RECT 74.120 22.040 74.500 22.080 ;
        RECT 74.110 21.850 74.500 22.040 ;
        RECT 74.120 21.820 74.500 21.850 ;
        RECT 73.560 21.340 73.950 21.380 ;
        RECT 73.550 21.150 73.950 21.340 ;
        RECT 73.560 21.120 73.950 21.150 ;
        RECT 73.780 20.040 73.950 21.120 ;
        RECT 73.570 20.000 73.950 20.040 ;
        RECT 73.560 19.880 73.950 20.000 ;
        RECT 74.330 19.880 74.500 21.820 ;
        RECT 74.880 21.390 75.050 22.280 ;
        RECT 75.220 22.050 75.540 22.090 ;
        RECT 76.310 22.050 76.630 22.090 ;
        RECT 75.210 21.860 75.540 22.050 ;
        RECT 76.300 21.860 76.630 22.050 ;
        RECT 75.220 21.830 75.540 21.860 ;
        RECT 76.310 21.830 76.630 21.860 ;
        RECT 74.670 21.350 75.050 21.390 ;
        RECT 75.760 21.370 76.080 21.410 ;
        RECT 74.660 21.160 75.050 21.350 ;
        RECT 75.750 21.180 76.080 21.370 ;
        RECT 74.670 21.130 75.050 21.160 ;
        RECT 75.760 21.150 76.080 21.180 ;
        RECT 74.880 20.040 75.050 21.130 ;
        RECT 74.670 20.000 75.050 20.040 ;
        RECT 75.760 20.000 76.080 20.040 ;
        RECT 74.660 19.880 75.050 20.000 ;
        RECT 73.560 19.810 73.890 19.880 ;
        RECT 74.660 19.810 74.990 19.880 ;
        RECT 75.750 19.810 76.080 20.000 ;
        RECT 73.570 19.780 73.890 19.810 ;
        RECT 74.670 19.780 74.990 19.810 ;
        RECT 75.760 19.780 76.080 19.810 ;
        RECT 22.090 19.560 22.410 19.600 ;
        RECT 22.230 18.450 22.400 19.560 ;
        RECT 52.500 19.530 52.660 19.560 ;
        RECT 52.500 19.300 52.670 19.530 ;
        RECT 53.050 19.520 53.210 19.560 ;
        RECT 52.500 19.260 52.870 19.300 ;
        RECT 53.050 19.280 53.220 19.520 ;
        RECT 53.600 19.300 53.770 19.590 ;
        RECT 54.150 19.520 54.310 19.560 ;
        RECT 54.700 19.520 54.860 19.560 ;
        RECT 55.250 19.540 55.410 19.560 ;
        RECT 58.230 19.540 58.390 19.560 ;
        RECT 52.500 19.180 52.880 19.260 ;
        RECT 53.050 19.180 53.280 19.280 ;
        RECT 53.600 19.260 53.970 19.300 ;
        RECT 54.150 19.280 54.320 19.520 ;
        RECT 54.700 19.300 54.870 19.520 ;
        RECT 53.600 19.180 53.980 19.260 ;
        RECT 54.150 19.180 54.380 19.280 ;
        RECT 54.700 19.260 55.070 19.300 ;
        RECT 55.250 19.280 55.420 19.540 ;
        RECT 58.220 19.280 58.390 19.540 ;
        RECT 58.780 19.520 58.940 19.560 ;
        RECT 59.330 19.520 59.490 19.560 ;
        RECT 58.770 19.300 58.940 19.520 ;
        RECT 54.700 19.180 55.080 19.260 ;
        RECT 55.250 19.180 55.480 19.280 ;
        RECT 52.550 19.070 52.880 19.180 ;
        RECT 52.550 19.040 52.870 19.070 ;
        RECT 22.090 18.420 22.410 18.450 ;
        RECT 22.080 18.310 22.410 18.420 ;
        RECT 19.480 18.210 19.710 18.310 ;
        RECT 19.880 18.230 20.260 18.310 ;
        RECT 19.540 17.950 19.710 18.210 ;
        RECT 19.890 18.190 20.260 18.230 ;
        RECT 20.580 18.210 20.810 18.310 ;
        RECT 20.980 18.230 21.360 18.310 ;
        RECT 20.090 17.970 20.260 18.190 ;
        RECT 20.640 17.970 20.810 18.210 ;
        RECT 20.990 18.190 21.360 18.230 ;
        RECT 21.680 18.210 21.910 18.310 ;
        RECT 22.080 18.230 22.460 18.310 ;
        RECT 19.550 17.930 19.710 17.950 ;
        RECT 20.100 17.930 20.260 17.970 ;
        RECT 20.650 17.930 20.810 17.970 ;
        RECT 21.190 17.900 21.360 18.190 ;
        RECT 21.740 17.970 21.910 18.210 ;
        RECT 22.090 18.190 22.460 18.230 ;
        RECT 21.750 17.930 21.910 17.970 ;
        RECT 22.290 17.960 22.460 18.190 ;
        RECT 22.300 17.930 22.460 17.960 ;
        RECT 52.560 17.930 52.730 19.040 ;
        RECT 52.550 17.890 52.870 17.930 ;
        RECT 19.480 17.720 19.650 17.880 ;
        RECT 19.340 17.690 19.660 17.720 ;
        RECT 19.330 17.500 19.660 17.690 ;
        RECT 19.340 17.460 19.660 17.500 ;
        RECT 19.480 16.380 19.650 17.460 ;
        RECT 19.330 16.350 19.650 16.380 ;
        RECT 19.000 15.440 19.170 16.200 ;
        RECT 19.320 16.160 19.650 16.350 ;
        RECT 19.330 16.120 19.650 16.160 ;
        RECT 19.480 15.380 19.650 16.120 ;
        RECT 20.030 15.680 20.200 17.880 ;
        RECT 20.580 17.720 20.750 17.880 ;
        RECT 20.440 17.690 20.760 17.720 ;
        RECT 20.430 17.500 20.760 17.690 ;
        RECT 20.440 17.460 20.760 17.500 ;
        RECT 20.580 16.370 20.750 17.460 ;
        RECT 20.440 16.340 20.760 16.370 ;
        RECT 20.430 16.150 20.760 16.340 ;
        RECT 20.440 16.110 20.760 16.150 ;
        RECT 19.890 15.650 20.210 15.680 ;
        RECT 19.880 15.460 20.210 15.650 ;
        RECT 19.890 15.420 20.210 15.460 ;
        RECT 20.030 15.380 20.200 15.420 ;
        RECT 20.580 15.380 20.750 16.110 ;
        RECT 21.130 15.670 21.300 17.880 ;
        RECT 21.680 17.720 21.850 17.880 ;
        RECT 21.530 17.690 21.850 17.720 ;
        RECT 21.520 17.500 21.850 17.690 ;
        RECT 21.530 17.460 21.850 17.500 ;
        RECT 21.680 16.350 21.850 17.460 ;
        RECT 21.530 16.320 21.850 16.350 ;
        RECT 21.520 16.130 21.850 16.320 ;
        RECT 21.530 16.090 21.850 16.130 ;
        RECT 20.990 15.640 21.310 15.670 ;
        RECT 20.980 15.450 21.310 15.640 ;
        RECT 20.990 15.410 21.310 15.450 ;
        RECT 21.130 15.380 21.300 15.410 ;
        RECT 21.680 15.380 21.850 16.090 ;
        RECT 22.230 15.670 22.400 17.870 ;
        RECT 52.550 17.700 52.880 17.890 ;
        RECT 52.550 17.670 52.870 17.700 ;
        RECT 51.730 17.310 52.240 17.390 ;
        RECT 51.730 17.290 52.250 17.310 ;
        RECT 51.730 17.250 52.300 17.290 ;
        RECT 51.730 17.060 52.310 17.250 ;
        RECT 51.740 17.030 52.300 17.060 ;
        RECT 51.740 16.820 52.250 17.030 ;
        RECT 51.740 16.780 52.310 16.820 ;
        RECT 52.560 16.790 52.730 17.670 ;
        RECT 53.110 17.250 53.280 19.180 ;
        RECT 53.650 19.070 53.980 19.180 ;
        RECT 53.650 19.040 53.970 19.070 ;
        RECT 53.660 17.930 53.830 19.040 ;
        RECT 53.650 17.890 53.970 17.930 ;
        RECT 53.650 17.700 53.980 17.890 ;
        RECT 53.650 17.670 53.970 17.700 ;
        RECT 53.110 17.210 53.430 17.250 ;
        RECT 53.110 17.020 53.440 17.210 ;
        RECT 53.110 16.990 53.430 17.020 ;
        RECT 53.110 16.780 53.280 16.990 ;
        RECT 53.660 16.780 53.830 17.670 ;
        RECT 54.210 17.250 54.380 19.180 ;
        RECT 54.750 19.070 55.080 19.180 ;
        RECT 54.750 19.040 55.070 19.070 ;
        RECT 54.760 17.930 54.930 19.040 ;
        RECT 54.750 17.890 55.070 17.930 ;
        RECT 54.750 17.700 55.080 17.890 ;
        RECT 54.750 17.670 55.070 17.700 ;
        RECT 54.200 17.210 54.520 17.250 ;
        RECT 54.200 17.020 54.530 17.210 ;
        RECT 54.200 16.990 54.520 17.020 ;
        RECT 54.210 16.780 54.380 16.990 ;
        RECT 54.760 16.780 54.930 17.670 ;
        RECT 55.310 17.260 55.480 19.180 ;
        RECT 58.160 19.180 58.390 19.280 ;
        RECT 58.570 19.260 58.940 19.300 ;
        RECT 59.320 19.280 59.490 19.520 ;
        RECT 59.870 19.300 60.040 19.590 ;
        RECT 62.310 19.560 62.470 19.590 ;
        RECT 60.430 19.520 60.590 19.560 ;
        RECT 60.980 19.530 61.140 19.560 ;
        RECT 58.560 19.180 58.940 19.260 ;
        RECT 59.260 19.180 59.490 19.280 ;
        RECT 59.670 19.260 60.040 19.300 ;
        RECT 60.420 19.280 60.590 19.520 ;
        RECT 60.970 19.300 61.140 19.530 ;
        RECT 59.660 19.180 60.040 19.260 ;
        RECT 60.360 19.180 60.590 19.280 ;
        RECT 60.770 19.260 61.140 19.300 ;
        RECT 60.760 19.180 61.140 19.260 ;
        RECT 62.310 19.330 62.480 19.560 ;
        RECT 62.860 19.550 63.020 19.590 ;
        RECT 62.310 19.290 62.680 19.330 ;
        RECT 62.860 19.310 63.030 19.550 ;
        RECT 63.410 19.330 63.580 19.620 ;
        RECT 63.960 19.550 64.120 19.590 ;
        RECT 64.510 19.550 64.670 19.590 ;
        RECT 65.060 19.570 65.220 19.590 ;
        RECT 68.040 19.570 68.200 19.590 ;
        RECT 62.310 19.210 62.690 19.290 ;
        RECT 62.860 19.210 63.090 19.310 ;
        RECT 63.410 19.290 63.780 19.330 ;
        RECT 63.960 19.310 64.130 19.550 ;
        RECT 64.510 19.330 64.680 19.550 ;
        RECT 63.410 19.210 63.790 19.290 ;
        RECT 63.960 19.210 64.190 19.310 ;
        RECT 64.510 19.290 64.880 19.330 ;
        RECT 65.060 19.310 65.230 19.570 ;
        RECT 68.030 19.310 68.200 19.570 ;
        RECT 68.590 19.550 68.750 19.590 ;
        RECT 69.140 19.550 69.300 19.590 ;
        RECT 68.580 19.330 68.750 19.550 ;
        RECT 64.510 19.210 64.890 19.290 ;
        RECT 65.060 19.210 65.290 19.310 ;
        RECT 58.160 17.260 58.330 19.180 ;
        RECT 58.560 19.070 58.890 19.180 ;
        RECT 58.570 19.040 58.890 19.070 ;
        RECT 58.710 17.930 58.880 19.040 ;
        RECT 58.570 17.890 58.890 17.930 ;
        RECT 58.560 17.700 58.890 17.890 ;
        RECT 58.570 17.670 58.890 17.700 ;
        RECT 55.300 17.220 55.620 17.260 ;
        RECT 58.020 17.220 58.340 17.260 ;
        RECT 55.300 17.030 55.630 17.220 ;
        RECT 58.010 17.030 58.340 17.220 ;
        RECT 55.300 17.000 55.620 17.030 ;
        RECT 58.020 17.000 58.340 17.030 ;
        RECT 55.310 16.780 55.480 17.000 ;
        RECT 58.160 16.780 58.330 17.000 ;
        RECT 58.710 16.780 58.880 17.670 ;
        RECT 59.260 17.250 59.430 19.180 ;
        RECT 59.660 19.070 59.990 19.180 ;
        RECT 59.670 19.040 59.990 19.070 ;
        RECT 59.810 17.930 59.980 19.040 ;
        RECT 59.670 17.890 59.990 17.930 ;
        RECT 59.660 17.700 59.990 17.890 ;
        RECT 59.670 17.670 59.990 17.700 ;
        RECT 59.120 17.210 59.440 17.250 ;
        RECT 59.110 17.020 59.440 17.210 ;
        RECT 59.120 16.990 59.440 17.020 ;
        RECT 59.260 16.780 59.430 16.990 ;
        RECT 59.810 16.780 59.980 17.670 ;
        RECT 60.360 17.250 60.530 19.180 ;
        RECT 60.760 19.070 61.090 19.180 ;
        RECT 62.360 19.100 62.690 19.210 ;
        RECT 62.360 19.070 62.680 19.100 ;
        RECT 60.770 19.040 61.090 19.070 ;
        RECT 60.910 17.930 61.080 19.040 ;
        RECT 62.370 17.960 62.540 19.070 ;
        RECT 60.770 17.890 61.090 17.930 ;
        RECT 60.760 17.700 61.090 17.890 ;
        RECT 62.360 17.920 62.680 17.960 ;
        RECT 62.360 17.730 62.690 17.920 ;
        RECT 62.360 17.700 62.680 17.730 ;
        RECT 60.770 17.670 61.090 17.700 ;
        RECT 60.210 17.210 60.530 17.250 ;
        RECT 60.200 17.020 60.530 17.210 ;
        RECT 60.210 16.990 60.530 17.020 ;
        RECT 60.360 16.780 60.530 16.990 ;
        RECT 60.910 16.790 61.080 17.670 ;
        RECT 61.540 17.390 62.050 17.420 ;
        RECT 61.400 17.340 62.050 17.390 ;
        RECT 61.400 17.320 62.060 17.340 ;
        RECT 61.400 17.310 62.110 17.320 ;
        RECT 61.390 17.290 62.110 17.310 ;
        RECT 61.340 17.280 62.110 17.290 ;
        RECT 61.340 17.250 62.120 17.280 ;
        RECT 61.330 17.090 62.120 17.250 ;
        RECT 61.330 17.060 62.110 17.090 ;
        RECT 61.340 17.030 62.060 17.060 ;
        RECT 61.390 16.850 62.060 17.030 ;
        RECT 61.390 16.820 62.120 16.850 ;
        RECT 62.370 16.820 62.540 17.700 ;
        RECT 62.920 17.280 63.090 19.210 ;
        RECT 63.460 19.100 63.790 19.210 ;
        RECT 63.460 19.070 63.780 19.100 ;
        RECT 63.470 17.960 63.640 19.070 ;
        RECT 63.460 17.920 63.780 17.960 ;
        RECT 63.460 17.730 63.790 17.920 ;
        RECT 63.460 17.700 63.780 17.730 ;
        RECT 62.920 17.240 63.240 17.280 ;
        RECT 62.920 17.050 63.250 17.240 ;
        RECT 62.920 17.020 63.240 17.050 ;
        RECT 61.330 16.810 62.120 16.820 ;
        RECT 62.920 16.810 63.090 17.020 ;
        RECT 63.470 16.810 63.640 17.700 ;
        RECT 64.020 17.280 64.190 19.210 ;
        RECT 64.560 19.100 64.890 19.210 ;
        RECT 64.560 19.070 64.880 19.100 ;
        RECT 64.570 17.960 64.740 19.070 ;
        RECT 64.560 17.920 64.880 17.960 ;
        RECT 64.560 17.730 64.890 17.920 ;
        RECT 64.560 17.700 64.880 17.730 ;
        RECT 64.010 17.240 64.330 17.280 ;
        RECT 64.010 17.050 64.340 17.240 ;
        RECT 64.010 17.020 64.330 17.050 ;
        RECT 64.020 16.810 64.190 17.020 ;
        RECT 64.570 16.810 64.740 17.700 ;
        RECT 65.120 17.290 65.290 19.210 ;
        RECT 67.970 19.210 68.200 19.310 ;
        RECT 68.380 19.290 68.750 19.330 ;
        RECT 69.130 19.310 69.300 19.550 ;
        RECT 69.680 19.330 69.850 19.620 ;
        RECT 70.240 19.550 70.400 19.590 ;
        RECT 70.790 19.560 70.950 19.590 ;
        RECT 68.370 19.210 68.750 19.290 ;
        RECT 69.070 19.210 69.300 19.310 ;
        RECT 69.480 19.290 69.850 19.330 ;
        RECT 70.230 19.310 70.400 19.550 ;
        RECT 70.780 19.330 70.950 19.560 ;
        RECT 69.470 19.210 69.850 19.290 ;
        RECT 70.170 19.210 70.400 19.310 ;
        RECT 70.580 19.290 70.950 19.330 ;
        RECT 70.570 19.210 70.950 19.290 ;
        RECT 67.970 17.290 68.140 19.210 ;
        RECT 68.370 19.100 68.700 19.210 ;
        RECT 68.380 19.070 68.700 19.100 ;
        RECT 68.520 17.960 68.690 19.070 ;
        RECT 68.380 17.920 68.700 17.960 ;
        RECT 68.370 17.730 68.700 17.920 ;
        RECT 68.380 17.700 68.700 17.730 ;
        RECT 65.110 17.250 65.430 17.290 ;
        RECT 67.830 17.250 68.150 17.290 ;
        RECT 65.110 17.060 65.440 17.250 ;
        RECT 67.820 17.060 68.150 17.250 ;
        RECT 65.110 17.030 65.430 17.060 ;
        RECT 67.830 17.030 68.150 17.060 ;
        RECT 65.120 16.810 65.290 17.030 ;
        RECT 67.970 16.810 68.140 17.030 ;
        RECT 68.520 16.810 68.690 17.700 ;
        RECT 69.070 17.280 69.240 19.210 ;
        RECT 69.470 19.100 69.800 19.210 ;
        RECT 69.480 19.070 69.800 19.100 ;
        RECT 69.620 17.960 69.790 19.070 ;
        RECT 69.480 17.920 69.800 17.960 ;
        RECT 69.470 17.730 69.800 17.920 ;
        RECT 69.480 17.700 69.800 17.730 ;
        RECT 68.930 17.240 69.250 17.280 ;
        RECT 68.920 17.050 69.250 17.240 ;
        RECT 68.930 17.020 69.250 17.050 ;
        RECT 69.070 16.810 69.240 17.020 ;
        RECT 69.620 16.810 69.790 17.700 ;
        RECT 70.170 17.280 70.340 19.210 ;
        RECT 70.570 19.100 70.900 19.210 ;
        RECT 70.580 19.070 70.900 19.100 ;
        RECT 70.720 17.960 70.890 19.070 ;
        RECT 70.580 17.920 70.900 17.960 ;
        RECT 70.570 17.730 70.900 17.920 ;
        RECT 70.580 17.700 70.900 17.730 ;
        RECT 70.020 17.240 70.340 17.280 ;
        RECT 70.010 17.050 70.340 17.240 ;
        RECT 70.020 17.020 70.340 17.050 ;
        RECT 70.170 16.810 70.340 17.020 ;
        RECT 70.720 16.820 70.890 17.700 ;
        RECT 71.210 17.340 71.720 17.420 ;
        RECT 71.200 17.320 71.720 17.340 ;
        RECT 71.150 17.280 71.720 17.320 ;
        RECT 71.140 17.090 71.720 17.280 ;
        RECT 72.130 17.100 72.300 19.500 ;
        RECT 72.680 17.100 72.850 19.500 ;
        RECT 73.230 17.100 73.400 19.500 ;
        RECT 73.780 17.270 73.950 19.570 ;
        RECT 74.330 19.310 74.500 19.570 ;
        RECT 74.120 19.270 74.500 19.310 ;
        RECT 74.110 19.080 74.500 19.270 ;
        RECT 74.120 19.050 74.500 19.080 ;
        RECT 74.330 17.940 74.500 19.050 ;
        RECT 74.120 17.900 74.500 17.940 ;
        RECT 74.110 17.710 74.500 17.900 ;
        RECT 74.120 17.680 74.500 17.710 ;
        RECT 73.570 17.230 73.950 17.270 ;
        RECT 73.560 17.100 73.950 17.230 ;
        RECT 74.330 17.100 74.500 17.680 ;
        RECT 74.880 17.260 75.050 19.570 ;
        RECT 75.430 19.310 75.600 19.570 ;
        RECT 75.220 19.270 75.600 19.310 ;
        RECT 75.210 19.190 75.600 19.270 ;
        RECT 75.980 19.190 76.150 19.570 ;
        RECT 76.530 19.310 76.700 19.570 ;
        RECT 76.320 19.270 76.700 19.310 ;
        RECT 76.310 19.190 76.700 19.270 ;
        RECT 75.210 19.080 75.540 19.190 ;
        RECT 76.310 19.080 76.640 19.190 ;
        RECT 75.220 19.050 75.540 19.080 ;
        RECT 76.320 19.050 76.640 19.080 ;
        RECT 75.220 17.900 75.540 17.940 ;
        RECT 76.320 17.900 76.640 17.940 ;
        RECT 75.210 17.710 75.540 17.900 ;
        RECT 76.310 17.710 76.640 17.900 ;
        RECT 75.220 17.680 75.540 17.710 ;
        RECT 76.320 17.680 76.640 17.710 ;
        RECT 77.240 17.590 77.410 18.810 ;
        RECT 76.950 17.300 77.460 17.400 ;
        RECT 76.890 17.260 77.460 17.300 ;
        RECT 74.670 17.220 75.050 17.260 ;
        RECT 75.760 17.220 76.080 17.260 ;
        RECT 74.660 17.100 75.050 17.220 ;
        RECT 71.150 17.060 71.710 17.090 ;
        RECT 71.200 16.850 71.710 17.060 ;
        RECT 73.560 17.040 73.890 17.100 ;
        RECT 73.570 17.010 73.890 17.040 ;
        RECT 74.660 17.030 74.990 17.100 ;
        RECT 75.750 17.030 76.080 17.220 ;
        RECT 76.880 17.070 77.460 17.260 ;
        RECT 76.890 17.040 77.450 17.070 ;
        RECT 74.670 17.000 74.990 17.030 ;
        RECT 75.760 17.000 76.080 17.030 ;
        RECT 71.140 16.810 71.710 16.850 ;
        RECT 76.940 16.830 77.450 17.040 ;
        RECT 61.330 16.780 62.130 16.810 ;
        RECT 51.740 16.590 52.320 16.780 ;
        RECT 61.320 16.620 62.130 16.780 ;
        RECT 71.130 16.620 71.710 16.810 ;
        RECT 76.880 16.790 77.450 16.830 ;
        RECT 61.320 16.590 62.120 16.620 ;
        RECT 71.140 16.590 71.710 16.620 ;
        RECT 76.870 16.600 77.450 16.790 ;
        RECT 51.740 16.560 52.310 16.590 ;
        RECT 61.330 16.560 62.060 16.590 ;
        RECT 51.740 16.380 52.250 16.560 ;
        RECT 61.390 16.410 62.060 16.560 ;
        RECT 71.200 16.410 71.710 16.590 ;
        RECT 76.880 16.570 77.450 16.600 ;
        RECT 61.390 16.380 61.900 16.410 ;
        RECT 76.940 16.390 77.450 16.570 ;
        RECT 22.080 15.640 22.400 15.670 ;
        RECT 22.070 15.450 22.400 15.640 ;
        RECT 22.080 15.410 22.400 15.450 ;
        RECT 22.230 15.380 22.400 15.410 ;
        RECT 23.650 15.280 26.040 15.650 ;
        RECT 23.700 12.020 26.040 15.280 ;
        RECT 102.520 14.480 102.750 14.590 ;
        RECT 102.420 14.380 107.080 14.480 ;
        RECT 102.420 14.310 107.270 14.380 ;
        RECT 105.980 14.210 106.310 14.310 ;
        RECT 106.940 14.210 107.270 14.310 ;
        RECT 107.900 14.210 108.230 14.380 ;
        RECT 108.860 14.210 109.190 14.380 ;
        RECT 108.130 13.970 108.320 13.980 ;
        RECT 103.640 13.790 107.440 13.800 ;
        RECT 108.100 13.790 108.360 13.970 ;
        RECT 103.640 13.650 108.360 13.790 ;
        RECT 103.640 13.630 108.230 13.650 ;
        RECT 105.980 13.530 106.310 13.630 ;
        RECT 106.940 13.620 108.230 13.630 ;
        RECT 106.940 13.530 107.440 13.620 ;
        RECT 107.900 13.530 108.230 13.620 ;
        RECT 108.860 13.530 109.190 13.700 ;
        RECT 107.210 13.160 107.440 13.530 ;
        RECT 108.130 13.300 108.320 13.310 ;
        RECT 108.100 13.160 108.360 13.300 ;
        RECT 107.210 12.980 108.360 13.160 ;
        RECT 102.520 12.870 102.750 12.980 ;
        RECT 107.210 12.950 108.220 12.980 ;
        RECT 102.420 12.700 106.900 12.870 ;
        RECT 107.210 12.770 107.440 12.950 ;
        RECT 105.980 12.600 106.310 12.700 ;
        RECT 106.940 12.600 107.440 12.770 ;
        RECT 107.900 12.600 108.230 12.770 ;
        RECT 108.860 12.600 109.190 12.770 ;
        RECT 107.210 12.190 107.440 12.600 ;
        RECT 103.670 12.020 107.440 12.190 ;
        RECT 23.700 12.010 26.030 12.020 ;
        RECT 105.980 11.920 106.310 12.020 ;
        RECT 106.940 11.920 107.440 12.020 ;
        RECT 107.900 11.940 108.230 12.090 ;
        RECT 107.900 11.920 108.620 11.940 ;
        RECT 108.860 11.920 109.190 12.090 ;
        RECT 102.520 11.270 102.750 11.380 ;
        RECT 102.420 11.100 106.920 11.270 ;
        RECT 107.210 11.160 107.440 11.920 ;
        RECT 108.170 11.750 108.620 11.920 ;
        RECT 108.190 11.730 108.620 11.750 ;
        RECT 105.980 10.990 106.310 11.100 ;
        RECT 106.940 10.990 107.440 11.160 ;
        RECT 107.900 10.990 108.230 11.160 ;
        RECT 108.860 10.990 109.190 11.160 ;
        RECT 107.210 10.580 107.440 10.990 ;
        RECT 103.680 10.410 107.440 10.580 ;
        RECT 105.980 10.310 106.310 10.410 ;
        RECT 106.940 10.310 107.440 10.410 ;
        RECT 107.900 10.330 108.230 10.480 ;
        RECT 107.900 10.310 108.620 10.330 ;
        RECT 108.860 10.310 109.190 10.480 ;
        RECT 106.420 10.120 106.850 10.140 ;
        RECT 106.400 9.950 106.850 10.120 ;
        RECT 106.420 9.930 106.850 9.950 ;
        RECT 102.520 9.650 102.750 9.760 ;
        RECT 102.420 9.480 106.920 9.650 ;
        RECT 105.980 9.380 106.310 9.480 ;
        RECT 107.210 8.980 107.440 10.310 ;
        RECT 108.170 10.140 108.620 10.310 ;
        RECT 108.190 10.120 108.620 10.140 ;
        RECT 107.900 9.380 108.230 9.550 ;
        RECT 108.860 9.380 109.190 9.550 ;
        RECT 103.670 8.810 107.440 8.980 ;
        RECT 105.980 8.700 106.310 8.810 ;
        RECT 107.210 8.560 107.440 8.810 ;
        RECT 107.900 8.720 108.230 8.870 ;
        RECT 107.900 8.700 108.610 8.720 ;
        RECT 108.860 8.700 109.190 8.870 ;
        RECT 107.210 8.540 107.710 8.560 ;
        RECT 107.210 8.370 107.730 8.540 ;
        RECT 108.160 8.530 108.610 8.700 ;
        RECT 108.180 8.510 108.610 8.530 ;
        RECT 107.210 8.350 107.710 8.370 ;
        RECT 102.520 8.050 102.750 8.160 ;
        RECT 102.420 7.880 106.870 8.050 ;
        RECT 107.210 7.940 107.440 8.350 ;
        RECT 105.980 7.770 106.310 7.880 ;
        RECT 106.940 7.770 107.440 7.940 ;
        RECT 108.400 7.830 108.730 8.000 ;
        RECT 108.860 7.770 109.190 7.940 ;
        RECT 107.210 7.360 107.440 7.770 ;
        RECT 103.650 7.190 107.440 7.360 ;
        RECT 105.980 7.090 106.310 7.190 ;
        RECT 106.940 7.090 107.440 7.190 ;
        RECT 108.400 7.150 108.730 7.320 ;
        RECT 102.520 6.430 102.750 6.540 ;
        RECT 102.420 6.260 106.920 6.430 ;
        RECT 107.210 6.330 107.440 7.090 ;
        RECT 108.190 7.080 108.620 7.100 ;
        RECT 108.860 7.090 109.190 7.260 ;
        RECT 108.170 6.910 108.620 7.080 ;
        RECT 108.710 6.960 109.140 6.980 ;
        RECT 108.190 6.890 108.620 6.910 ;
        RECT 108.690 6.790 109.140 6.960 ;
        RECT 108.710 6.770 109.140 6.790 ;
        RECT 105.980 6.160 106.310 6.260 ;
        RECT 106.940 6.160 107.440 6.330 ;
        RECT 107.900 6.160 108.230 6.330 ;
        RECT 108.860 6.160 109.190 6.330 ;
        RECT 107.210 5.740 107.440 6.160 ;
        RECT 103.650 5.570 107.440 5.740 ;
        RECT 105.980 5.480 106.310 5.570 ;
        RECT 106.940 5.480 107.440 5.570 ;
        RECT 107.900 5.490 108.230 5.650 ;
        RECT 107.900 5.480 108.610 5.490 ;
        RECT 108.860 5.480 109.190 5.650 ;
        RECT 102.520 4.830 102.750 4.940 ;
        RECT 102.420 4.660 106.840 4.830 ;
        RECT 107.210 4.720 107.440 5.480 ;
        RECT 108.180 5.470 108.610 5.480 ;
        RECT 108.160 5.300 108.610 5.470 ;
        RECT 108.180 5.280 108.610 5.300 ;
        RECT 113.880 5.020 114.250 19.890 ;
        RECT 113.880 4.770 114.260 5.020 ;
        RECT 105.980 4.550 106.310 4.660 ;
        RECT 106.940 4.550 107.440 4.720 ;
        RECT 107.900 4.550 108.230 4.720 ;
        RECT 108.860 4.550 109.190 4.720 ;
        RECT 107.210 4.150 107.440 4.550 ;
        RECT 103.650 3.980 107.450 4.150 ;
        RECT 105.980 3.870 106.310 3.980 ;
        RECT 106.940 3.870 107.440 3.980 ;
        RECT 102.520 3.200 102.750 3.320 ;
        RECT 102.420 3.030 106.880 3.200 ;
        RECT 107.210 3.110 107.440 3.870 ;
        RECT 107.630 3.600 107.840 4.030 ;
        RECT 107.900 3.870 108.230 4.040 ;
        RECT 108.860 3.870 109.190 4.040 ;
        RECT 107.650 3.580 107.820 3.600 ;
        RECT 105.980 2.940 106.310 3.030 ;
        RECT 106.940 2.940 107.440 3.110 ;
        RECT 107.900 2.940 108.230 3.110 ;
        RECT 108.860 2.940 109.190 3.110 ;
        RECT 107.210 2.540 107.440 2.940 ;
        RECT 103.650 2.370 107.440 2.540 ;
        RECT 105.980 2.260 106.310 2.370 ;
        RECT 106.940 2.260 107.270 2.370 ;
        RECT 107.900 2.290 108.230 2.430 ;
        RECT 107.900 2.260 108.610 2.290 ;
        RECT 108.860 2.260 109.190 2.430 ;
        RECT 108.160 2.100 108.610 2.260 ;
        RECT 108.180 2.080 108.610 2.100 ;
        RECT 104.940 0.560 105.370 0.580 ;
        RECT 105.880 0.560 106.310 0.580 ;
        RECT 108.140 0.560 108.570 0.580 ;
        RECT 104.920 0.390 105.370 0.560 ;
        RECT 105.860 0.390 106.310 0.560 ;
        RECT 106.830 0.540 107.260 0.560 ;
        RECT 104.940 0.370 105.370 0.390 ;
        RECT 105.880 0.370 106.310 0.390 ;
        RECT 106.810 0.370 107.260 0.540 ;
        RECT 108.120 0.390 108.570 0.560 ;
        RECT 108.140 0.370 108.570 0.390 ;
        RECT 106.830 0.350 107.260 0.370 ;
      LAYER mcon ;
        RECT 0.460 72.120 0.630 72.290 ;
        RECT 15.150 72.530 15.320 72.700 ;
        RECT 15.150 72.080 15.320 72.250 ;
        RECT 19.850 72.480 20.020 72.650 ;
        RECT 19.850 72.030 20.020 72.200 ;
        RECT 86.760 71.340 87.030 71.610 ;
        RECT 130.980 71.340 131.250 71.610 ;
        RECT 15.150 69.540 15.320 69.710 ;
        RECT 86.760 69.610 87.030 69.880 ;
        RECT 130.980 69.610 131.250 69.880 ;
        RECT 14.130 69.360 14.300 69.530 ;
        RECT 4.000 69.000 4.170 69.170 ;
        RECT 15.150 69.090 15.320 69.260 ;
        RECT 1.130 68.790 1.300 68.960 ;
        RECT 2.540 68.790 2.710 68.960 ;
        RECT 14.130 68.670 14.300 68.840 ;
        RECT 87.890 68.830 88.070 69.000 ;
        RECT 15.150 68.530 15.320 68.700 ;
        RECT 86.080 68.530 86.250 68.700 ;
        RECT 1.130 67.940 1.300 68.110 ;
        RECT 1.710 68.080 1.880 68.250 ;
        RECT 2.540 67.940 2.710 68.110 ;
        RECT 3.740 68.080 3.910 68.250 ;
        RECT 15.150 68.080 15.320 68.250 ;
        RECT 92.980 68.470 93.150 68.640 ;
        RECT 1.310 67.530 1.480 67.700 ;
        RECT 2.370 67.530 2.540 67.700 ;
        RECT 1.130 67.120 1.300 67.290 ;
        RECT 1.710 67.240 1.880 67.410 ;
        RECT 17.100 67.340 17.270 67.510 ;
        RECT 86.430 67.690 86.610 67.880 ;
        RECT 18.460 67.420 18.630 67.590 ;
        RECT 2.540 67.120 2.710 67.290 ;
        RECT 19.150 67.410 19.320 67.580 ;
        RECT 3.740 66.650 3.910 66.820 ;
        RECT 14.130 66.560 14.300 66.730 ;
        RECT 1.130 66.280 1.300 66.450 ;
        RECT 2.540 66.280 2.710 66.450 ;
        RECT 3.170 66.100 3.340 66.270 ;
        RECT 14.130 65.870 14.300 66.040 ;
        RECT 1.130 65.160 1.300 65.330 ;
        RECT 3.400 65.350 3.570 65.520 ;
        RECT 4.010 65.380 4.180 65.550 ;
        RECT 2.540 65.160 2.710 65.330 ;
        RECT 14.130 65.010 14.300 65.180 ;
        RECT 1.690 64.440 1.860 64.610 ;
        RECT 3.120 64.460 3.290 64.630 ;
        RECT 14.130 64.320 14.300 64.490 ;
        RECT 93.450 67.910 93.620 68.080 ;
        RECT 105.840 68.380 106.010 68.550 ;
        RECT 105.840 67.930 106.010 68.100 ;
        RECT 130.210 68.380 130.380 68.550 ;
        RECT 131.760 68.530 131.930 68.700 ;
        RECT 130.210 67.930 130.380 68.100 ;
        RECT 125.470 67.430 125.640 67.600 ;
        RECT 92.130 66.860 92.300 67.030 ;
        RECT 131.400 67.690 131.580 67.880 ;
        RECT 92.980 66.480 93.150 66.650 ;
        RECT 0.900 63.860 1.070 64.030 ;
        RECT 1.830 63.860 2.000 64.030 ;
        RECT 2.530 63.860 2.700 64.030 ;
        RECT 3.270 63.860 3.440 64.030 ;
        RECT 3.980 63.850 4.150 64.020 ;
        RECT 28.500 65.650 28.670 65.820 ;
        RECT 87.010 65.310 87.280 65.580 ;
        RECT 92.990 65.410 93.160 65.580 ;
        RECT 93.450 65.590 93.620 65.760 ;
        RECT 98.820 65.900 98.990 66.070 ;
        RECT 119.020 65.900 119.190 66.070 ;
        RECT 86.430 64.050 86.610 64.240 ;
        RECT 16.380 63.680 16.550 63.850 ;
        RECT 26.240 63.700 26.410 63.870 ;
        RECT 87.010 63.580 87.280 63.850 ;
        RECT 92.120 65.170 92.290 65.340 ;
        RECT 124.940 65.310 125.210 65.580 ;
        RECT 128.010 65.500 128.180 65.670 ;
        RECT 129.670 65.460 129.840 65.630 ;
        RECT 125.470 64.670 125.640 64.840 ;
        RECT 127.960 64.850 128.130 65.020 ;
        RECT 128.950 65.110 129.120 65.280 ;
        RECT 93.440 64.010 93.610 64.180 ;
        RECT 129.020 64.080 129.190 64.250 ;
        RECT 93.010 63.500 93.180 63.670 ;
        RECT 105.840 63.730 106.010 63.900 ;
        RECT 124.940 63.580 125.210 63.850 ;
        RECT 127.960 63.590 128.130 63.760 ;
        RECT 86.080 63.230 86.250 63.400 ;
        RECT 105.840 63.280 106.010 63.450 ;
        RECT 128.950 63.330 129.120 63.500 ;
        RECT 130.210 63.730 130.380 63.900 ;
        RECT 87.890 62.930 88.070 63.100 ;
        RECT 88.140 62.800 88.320 62.970 ;
        RECT 25.370 61.760 25.800 62.500 ;
        RECT 48.730 62.330 48.940 62.540 ;
        RECT 86.330 62.500 86.500 62.670 ;
        RECT 47.260 61.960 47.430 62.130 ;
        RECT 49.690 61.860 49.860 62.030 ;
        RECT 50.730 61.900 50.900 62.070 ;
        RECT 51.770 61.560 51.940 61.730 ;
        RECT 86.680 61.660 86.860 61.850 ;
        RECT 51.770 61.200 51.940 61.370 ;
        RECT 87.880 62.350 88.050 62.520 ;
        RECT 87.880 61.900 88.050 62.070 ;
        RECT 128.010 62.940 128.180 63.110 ;
        RECT 131.400 64.050 131.580 64.240 ;
        RECT 129.720 63.240 129.890 63.410 ;
        RECT 130.210 63.280 130.380 63.450 ;
        RECT 131.760 63.230 131.930 63.400 ;
        RECT 48.730 60.580 48.940 60.790 ;
        RECT 99.880 61.810 100.050 61.980 ;
        RECT 124.170 62.350 124.340 62.520 ;
        RECT 125.720 62.500 125.890 62.670 ;
        RECT 124.170 61.900 124.340 62.070 ;
        RECT 92.620 61.400 92.790 61.570 ;
        RECT 119.430 61.400 119.600 61.570 ;
        RECT 128.010 62.500 128.180 62.670 ;
        RECT 129.710 62.520 129.880 62.690 ;
        RECT 125.360 61.660 125.540 61.850 ;
        RECT 127.960 61.850 128.130 62.020 ;
        RECT 128.950 62.110 129.120 62.280 ;
        RECT 129.020 61.490 129.190 61.660 ;
        RECT 47.260 60.210 47.430 60.380 ;
        RECT 127.960 60.590 128.130 60.760 ;
        RECT 49.690 60.110 49.860 60.280 ;
        RECT 50.730 60.150 50.900 60.320 ;
        RECT 51.770 59.810 51.940 59.980 ;
        RECT 99.070 59.870 99.240 60.040 ;
        RECT 112.980 59.870 113.150 60.040 ;
        RECT 123.470 60.040 123.640 60.210 ;
        RECT 128.950 60.330 129.120 60.500 ;
        RECT 51.770 59.450 51.940 59.620 ;
        RECT 22.590 59.040 22.760 59.210 ;
        RECT 23.680 59.050 23.850 59.220 ;
        RECT 48.730 58.830 48.940 59.040 ;
        RECT 47.260 58.460 47.430 58.630 ;
        RECT 49.690 58.360 49.860 58.530 ;
        RECT 73.660 58.600 73.920 59.420 ;
        RECT 85.610 58.630 85.930 59.420 ;
        RECT 115.520 59.740 115.690 59.910 ;
        RECT 87.060 59.060 87.240 59.250 ;
        RECT 21.050 58.130 21.220 58.300 ;
        RECT 22.600 58.050 22.770 58.220 ;
        RECT 23.380 58.000 23.550 58.170 ;
        RECT 23.690 58.060 23.860 58.230 ;
        RECT 50.730 58.400 50.900 58.570 ;
        RECT 51.770 58.060 51.940 58.230 ;
        RECT 86.680 58.020 86.860 58.210 ;
        RECT 51.770 57.700 51.940 57.870 ;
        RECT 21.030 57.210 21.200 57.380 ;
        RECT 114.580 59.060 114.750 59.230 ;
        RECT 115.060 59.120 115.230 59.290 ;
        RECT 121.970 59.470 122.140 59.640 ;
        RECT 128.010 59.940 128.180 60.110 ;
        RECT 129.630 60.270 129.800 60.440 ;
        RECT 116.250 59.060 116.420 59.230 ;
        RECT 117.170 59.130 117.340 59.300 ;
        RECT 123.630 59.430 123.800 59.600 ;
        RECT 92.620 58.640 92.790 58.810 ;
        RECT 119.430 58.640 119.600 58.810 ;
        RECT 121.920 58.820 122.090 58.990 ;
        RECT 122.910 59.080 123.080 59.250 ;
        RECT 123.620 59.210 123.790 59.380 ;
        RECT 99.910 58.120 100.080 58.290 ;
        RECT 122.780 58.390 122.950 58.560 ;
        RECT 87.880 57.700 88.050 57.870 ;
        RECT 114.590 57.930 114.760 58.100 ;
        RECT 122.980 58.050 123.150 58.220 ;
        RECT 22.600 57.060 22.770 57.230 ;
        RECT 23.690 57.070 23.860 57.240 ;
        RECT 48.730 57.080 48.940 57.290 ;
        RECT 86.330 57.200 86.500 57.370 ;
        RECT 87.880 57.250 88.050 57.420 ;
        RECT 47.260 56.710 47.430 56.880 ;
        RECT 49.690 56.610 49.860 56.780 ;
        RECT 88.140 56.900 88.320 57.070 ;
        RECT 121.920 57.560 122.090 57.730 ;
        RECT 122.910 57.300 123.080 57.470 ;
        RECT 124.170 57.700 124.340 57.870 ;
        RECT 125.360 58.020 125.540 58.210 ;
        RECT 121.970 56.910 122.140 57.080 ;
        RECT 21.010 56.220 21.180 56.390 ;
        RECT 22.510 56.330 22.680 56.500 ;
        RECT 23.810 56.230 23.980 56.400 ;
        RECT 50.730 56.650 50.900 56.820 ;
        RECT 123.680 57.280 123.850 57.380 ;
        RECT 123.510 57.210 123.850 57.280 ;
        RECT 124.170 57.250 124.340 57.420 ;
        RECT 123.510 57.110 123.680 57.210 ;
        RECT 125.720 57.200 125.890 57.370 ;
        RECT 51.770 56.310 51.940 56.480 ;
        RECT 115.520 56.540 115.690 56.710 ;
        RECT 121.970 56.470 122.140 56.640 ;
        RECT 51.770 55.950 51.940 56.120 ;
        RECT 103.130 55.860 103.300 56.030 ;
        RECT 22.510 55.340 22.680 55.510 ;
        RECT 23.810 55.240 23.980 55.410 ;
        RECT 103.140 55.140 103.310 55.310 ;
        RECT 108.920 55.860 109.090 56.030 ;
        RECT 114.580 55.860 114.750 56.030 ;
        RECT 115.060 55.920 115.230 56.090 ;
        RECT 123.670 56.490 123.840 56.660 ;
        RECT 123.900 56.380 124.070 56.550 ;
        RECT 116.250 55.860 116.420 56.030 ;
        RECT 117.170 55.930 117.340 56.100 ;
        RECT 121.920 55.820 122.090 55.990 ;
        RECT 122.910 56.080 123.080 56.250 ;
        RECT 108.920 55.140 109.090 55.310 ;
        RECT 122.980 55.460 123.150 55.630 ;
        RECT 114.080 54.920 114.250 55.110 ;
        RECT 114.590 55.130 114.760 55.300 ;
        RECT 114.590 54.730 114.760 54.900 ;
        RECT 22.510 54.350 22.680 54.520 ;
        RECT 121.920 54.560 122.090 54.730 ;
        RECT 22.950 53.900 23.120 54.070 ;
        RECT 23.810 54.250 23.980 54.420 ;
        RECT 122.910 54.300 123.080 54.470 ;
        RECT 114.580 54.000 114.750 54.170 ;
        RECT 115.060 53.940 115.230 54.110 ;
        RECT 116.250 54.000 116.420 54.170 ;
        RECT 117.170 53.930 117.340 54.100 ;
        RECT 117.430 54.010 117.600 54.180 ;
        RECT 121.970 53.910 122.140 54.080 ;
        RECT 123.590 54.240 123.760 54.410 ;
        RECT 115.520 53.320 115.690 53.490 ;
        RECT 61.630 53.080 61.800 53.250 ;
        RECT 62.470 52.960 62.640 53.130 ;
        RECT 63.220 52.960 63.390 53.130 ;
        RECT 61.500 52.440 61.670 52.610 ;
        RECT 66.200 52.630 66.370 52.800 ;
        RECT 61.810 52.250 61.980 52.420 ;
        RECT 66.600 53.080 66.770 53.250 ;
        RECT 117.580 53.180 117.750 53.350 ;
        RECT 66.600 52.720 66.770 52.890 ;
        RECT 51.770 51.790 51.940 51.960 ;
        RECT 66.200 51.870 66.370 52.040 ;
        RECT 51.770 51.430 51.940 51.600 ;
        RECT 62.470 51.540 62.640 51.710 ;
        RECT 63.220 51.540 63.390 51.710 ;
        RECT 65.220 51.550 65.390 51.720 ;
        RECT 66.600 52.140 66.770 52.310 ;
        RECT 116.740 52.360 116.910 52.530 ;
        RECT 66.600 51.780 66.770 51.950 ;
        RECT 114.590 51.930 114.760 52.100 ;
        RECT 114.080 51.720 114.250 51.890 ;
        RECT 47.260 51.030 47.430 51.200 ;
        RECT 49.690 51.130 49.860 51.300 ;
        RECT 50.730 51.090 50.900 51.260 ;
        RECT 48.730 50.620 48.940 50.830 ;
        RECT 114.580 50.800 114.750 50.970 ;
        RECT 115.060 50.740 115.230 50.910 ;
        RECT 117.470 51.080 117.640 51.250 ;
        RECT 116.250 50.800 116.420 50.970 ;
        RECT 117.170 50.730 117.340 50.900 ;
        RECT 51.770 50.040 51.940 50.210 ;
        RECT 115.520 50.120 115.690 50.290 ;
        RECT 117.860 50.350 118.030 50.520 ;
        RECT 51.770 49.680 51.940 49.850 ;
        RECT 61.630 49.880 61.800 50.050 ;
        RECT 62.470 49.760 62.640 49.930 ;
        RECT 63.220 49.760 63.390 49.930 ;
        RECT 47.260 49.280 47.430 49.450 ;
        RECT 49.690 49.380 49.860 49.550 ;
        RECT 50.730 49.340 50.900 49.510 ;
        RECT 61.500 49.240 61.670 49.410 ;
        RECT 66.200 49.430 66.370 49.600 ;
        RECT 48.730 48.870 48.940 49.080 ;
        RECT 61.810 49.050 61.980 49.220 ;
        RECT 66.600 49.880 66.770 50.050 ;
        RECT 66.600 49.520 66.770 49.690 ;
        RECT 66.200 48.670 66.370 48.840 ;
        RECT 51.770 48.290 51.940 48.460 ;
        RECT 62.470 48.340 62.640 48.510 ;
        RECT 63.220 48.340 63.390 48.510 ;
        RECT 65.220 48.350 65.390 48.520 ;
        RECT 66.600 48.940 66.770 49.110 ;
        RECT 71.990 49.000 72.260 49.270 ;
        RECT 76.020 49.070 76.290 49.340 ;
        RECT 111.330 49.070 111.600 49.340 ;
        RECT 115.360 49.000 115.630 49.270 ;
        RECT 66.600 48.580 66.770 48.750 ;
        RECT 51.770 47.930 51.940 48.100 ;
        RECT 47.260 47.530 47.430 47.700 ;
        RECT 49.690 47.630 49.860 47.800 ;
        RECT 50.730 47.590 50.900 47.760 ;
        RECT 80.320 47.940 80.490 48.110 ;
        RECT 107.130 47.940 107.300 48.110 ;
        RECT 78.650 47.530 78.820 47.700 ;
        RECT 48.730 47.120 48.940 47.330 ;
        RECT 79.380 47.500 79.550 47.670 ;
        RECT 80.320 47.390 80.490 47.560 ;
        RECT 107.130 47.390 107.300 47.560 ;
        RECT 108.070 47.500 108.240 47.670 ;
        RECT 108.800 47.530 108.970 47.700 ;
        RECT 51.770 46.540 51.940 46.710 ;
        RECT 51.770 46.180 51.940 46.350 ;
        RECT 84.260 46.430 84.430 46.600 ;
        RECT 47.260 45.780 47.430 45.950 ;
        RECT 49.690 45.880 49.860 46.050 ;
        RECT 50.730 45.840 50.900 46.010 ;
        RECT 88.200 46.440 88.370 46.610 ;
        RECT 99.250 46.440 99.420 46.610 ;
        RECT 103.190 46.430 103.360 46.600 ;
        RECT 48.730 45.370 48.940 45.580 ;
        RECT 78.650 45.150 78.820 45.320 ;
        RECT 79.380 45.180 79.550 45.350 ;
        RECT 80.320 45.290 80.490 45.460 ;
        RECT 80.320 44.700 80.490 44.910 ;
        RECT 84.260 44.840 84.430 45.010 ;
        RECT 84.260 44.480 84.430 44.650 ;
        RECT 78.650 44.290 78.820 44.460 ;
        RECT 79.380 44.260 79.550 44.430 ;
        RECT 80.320 44.150 80.490 44.320 ;
        RECT 88.190 44.980 88.360 45.150 ;
        RECT 88.190 44.620 88.360 44.790 ;
        RECT 107.130 45.290 107.300 45.460 ;
        RECT 99.260 44.980 99.430 45.150 ;
        RECT 99.260 44.620 99.430 44.790 ;
        RECT 108.070 45.180 108.240 45.350 ;
        RECT 108.800 45.150 108.970 45.320 ;
        RECT 103.190 44.840 103.360 45.010 ;
        RECT 105.550 44.720 105.730 44.890 ;
        RECT 107.130 44.700 107.300 44.910 ;
        RECT 103.190 44.480 103.360 44.650 ;
        RECT 107.130 44.150 107.300 44.320 ;
        RECT 108.070 44.260 108.240 44.430 ;
        RECT 108.800 44.290 108.970 44.460 ;
        RECT 61.610 42.610 61.780 42.780 ;
        RECT 62.450 42.490 62.620 42.660 ;
        RECT 63.200 42.490 63.370 42.660 ;
        RECT 61.480 41.970 61.650 42.140 ;
        RECT 66.180 42.160 66.350 42.330 ;
        RECT 51.770 41.660 51.940 41.830 ;
        RECT 61.790 41.780 61.960 41.950 ;
        RECT 66.580 42.610 66.750 42.780 ;
        RECT 66.580 42.250 66.750 42.420 ;
        RECT 78.650 41.920 78.820 42.090 ;
        RECT 79.380 41.950 79.550 42.120 ;
        RECT 80.320 42.060 80.490 42.230 ;
        RECT 107.130 42.060 107.300 42.230 ;
        RECT 108.070 41.950 108.240 42.120 ;
        RECT 108.800 41.920 108.970 42.090 ;
        RECT 51.770 41.300 51.940 41.470 ;
        RECT 66.180 41.400 66.350 41.570 ;
        RECT 47.260 40.900 47.430 41.070 ;
        RECT 49.690 41.000 49.860 41.170 ;
        RECT 50.730 40.960 50.900 41.130 ;
        RECT 62.450 41.070 62.620 41.240 ;
        RECT 63.200 41.070 63.370 41.240 ;
        RECT 65.200 41.080 65.370 41.250 ;
        RECT 66.580 41.670 66.750 41.840 ;
        RECT 80.320 41.510 80.490 41.680 ;
        RECT 66.580 41.310 66.750 41.480 ;
        RECT 107.130 41.510 107.300 41.680 ;
        RECT 48.730 40.490 48.940 40.700 ;
        RECT 72.590 40.120 72.860 40.390 ;
        RECT 51.770 39.910 51.940 40.080 ;
        RECT 76.620 40.190 76.890 40.460 ;
        RECT 51.770 39.550 51.940 39.720 ;
        RECT 47.260 39.150 47.430 39.320 ;
        RECT 49.690 39.250 49.860 39.420 ;
        RECT 50.730 39.210 50.900 39.380 ;
        RECT 61.610 39.410 61.780 39.580 ;
        RECT 62.450 39.290 62.620 39.460 ;
        RECT 63.200 39.290 63.370 39.460 ;
        RECT 48.730 38.740 48.940 38.950 ;
        RECT 61.480 38.770 61.650 38.940 ;
        RECT 66.180 38.960 66.350 39.130 ;
        RECT 61.790 38.580 61.960 38.750 ;
        RECT 51.770 38.160 51.940 38.330 ;
        RECT 66.580 39.410 66.750 39.580 ;
        RECT 66.580 39.050 66.750 39.220 ;
        RECT 80.920 39.100 81.090 39.270 ;
        RECT 79.250 38.690 79.420 38.860 ;
        RECT 66.180 38.200 66.350 38.370 ;
        RECT 51.770 37.800 51.940 37.970 ;
        RECT 62.450 37.870 62.620 38.040 ;
        RECT 63.200 37.870 63.370 38.040 ;
        RECT 65.200 37.880 65.370 38.050 ;
        RECT 66.580 38.470 66.750 38.640 ;
        RECT 66.580 38.110 66.750 38.280 ;
        RECT 79.980 38.660 80.150 38.830 ;
        RECT 80.920 38.550 81.090 38.720 ;
        RECT 47.260 37.400 47.430 37.570 ;
        RECT 49.690 37.500 49.860 37.670 ;
        RECT 50.730 37.460 50.900 37.630 ;
        RECT 84.990 37.530 85.160 37.700 ;
        RECT 48.730 36.990 48.940 37.200 ;
        RECT 89.010 37.560 89.180 37.730 ;
        RECT 51.770 36.410 51.940 36.580 ;
        RECT 79.250 36.330 79.420 36.500 ;
        RECT 79.980 36.360 80.150 36.530 ;
        RECT 80.920 36.470 81.090 36.640 ;
        RECT 84.980 36.330 85.150 36.500 ;
        RECT 51.770 36.050 51.940 36.220 ;
        RECT 47.260 35.650 47.430 35.820 ;
        RECT 49.690 35.750 49.860 35.920 ;
        RECT 50.730 35.710 50.900 35.880 ;
        RECT 80.920 35.860 81.090 36.090 ;
        RECT 48.730 35.240 48.940 35.450 ;
        RECT 84.980 35.670 85.150 35.840 ;
        RECT 79.250 35.450 79.420 35.620 ;
        RECT 79.980 35.420 80.150 35.590 ;
        RECT 80.920 35.310 81.090 35.480 ;
        RECT 89.000 36.270 89.170 36.440 ;
        RECT 89.000 35.630 89.170 35.800 ;
        RECT 61.640 33.340 61.810 33.510 ;
        RECT 27.000 33.070 27.170 33.240 ;
        RECT 27.650 33.070 27.820 33.240 ;
        RECT 62.480 33.220 62.650 33.390 ;
        RECT 63.230 33.220 63.400 33.390 ;
        RECT 25.780 32.630 25.950 32.800 ;
        RECT 26.480 32.630 26.650 32.800 ;
        RECT 25.100 30.860 25.270 31.030 ;
        RECT 51.730 32.600 51.900 32.770 ;
        RECT 61.510 32.700 61.680 32.870 ;
        RECT 66.210 32.890 66.380 33.060 ;
        RECT 28.020 32.400 28.190 32.570 ;
        RECT 51.730 32.240 51.900 32.410 ;
        RECT 61.820 32.510 61.990 32.680 ;
        RECT 66.610 33.340 66.780 33.510 ;
        RECT 66.610 32.980 66.780 33.150 ;
        RECT 79.250 33.080 79.420 33.250 ;
        RECT 96.850 33.460 97.020 33.630 ;
        RECT 79.980 33.110 80.150 33.280 ;
        RECT 80.920 33.220 81.090 33.390 ;
        RECT 96.100 33.160 96.270 33.330 ;
        RECT 95.950 32.920 96.120 33.090 ;
        RECT 80.920 32.670 81.090 32.840 ;
        RECT 98.110 32.890 98.280 33.060 ;
        RECT 47.220 31.840 47.390 32.010 ;
        RECT 49.650 31.940 49.820 32.110 ;
        RECT 50.690 31.900 50.860 32.070 ;
        RECT 66.210 32.130 66.380 32.300 ;
        RECT 62.480 31.800 62.650 31.970 ;
        RECT 63.230 31.800 63.400 31.970 ;
        RECT 65.230 31.810 65.400 31.980 ;
        RECT 66.610 32.400 66.780 32.570 ;
        RECT 95.950 32.480 96.120 32.650 ;
        RECT 98.110 32.510 98.280 32.680 ;
        RECT 66.610 32.040 66.780 32.210 ;
        RECT 96.100 32.240 96.270 32.410 ;
        RECT 96.850 31.940 97.020 32.110 ;
        RECT 48.690 31.430 48.900 31.640 ;
        RECT 27.930 30.830 28.100 31.000 ;
        RECT 51.730 30.850 51.900 31.020 ;
        RECT 27.940 30.290 28.110 30.460 ;
        RECT 51.730 30.490 51.900 30.660 ;
        RECT 96.850 30.690 97.020 30.860 ;
        RECT 22.700 28.280 22.870 28.450 ;
        RECT 19.390 27.840 19.560 28.010 ;
        RECT 20.490 27.850 20.660 28.020 ;
        RECT 21.580 27.850 21.750 28.020 ;
        RECT 22.710 27.810 22.880 27.980 ;
        RECT 19.940 27.170 20.110 27.340 ;
        RECT 19.940 25.800 20.110 25.970 ;
        RECT 47.220 30.090 47.390 30.260 ;
        RECT 49.650 30.190 49.820 30.360 ;
        RECT 50.690 30.150 50.860 30.320 ;
        RECT 96.100 30.390 96.270 30.560 ;
        RECT 61.640 30.140 61.810 30.310 ;
        RECT 48.690 29.680 48.900 29.890 ;
        RECT 62.480 30.020 62.650 30.190 ;
        RECT 63.230 30.020 63.400 30.190 ;
        RECT 28.010 29.420 28.180 29.590 ;
        RECT 61.510 29.500 61.680 29.670 ;
        RECT 66.210 29.690 66.380 29.860 ;
        RECT 51.730 29.100 51.900 29.270 ;
        RECT 61.820 29.310 61.990 29.480 ;
        RECT 25.810 28.750 25.980 28.920 ;
        RECT 26.500 28.740 26.670 28.910 ;
        RECT 66.610 30.140 66.780 30.310 ;
        RECT 95.950 30.150 96.120 30.320 ;
        RECT 66.610 29.780 66.780 29.950 ;
        RECT 98.110 30.120 98.280 30.290 ;
        RECT 83.970 29.580 84.140 29.750 ;
        RECT 95.950 29.710 96.120 29.880 ;
        RECT 98.110 29.740 98.280 29.910 ;
        RECT 51.730 28.740 51.900 28.910 ;
        RECT 66.210 28.930 66.380 29.100 ;
        RECT 47.220 28.340 47.390 28.510 ;
        RECT 49.650 28.440 49.820 28.610 ;
        RECT 50.690 28.400 50.860 28.570 ;
        RECT 62.480 28.600 62.650 28.770 ;
        RECT 63.230 28.600 63.400 28.770 ;
        RECT 65.230 28.610 65.400 28.780 ;
        RECT 66.610 29.200 66.780 29.370 ;
        RECT 66.610 28.840 66.780 29.010 ;
        RECT 96.100 29.470 96.270 29.640 ;
        RECT 96.850 29.170 97.020 29.340 ;
        RECT 84.020 28.620 84.190 28.790 ;
        RECT 26.980 27.970 27.150 28.140 ;
        RECT 27.690 27.910 27.860 28.080 ;
        RECT 48.690 27.930 48.900 28.140 ;
        RECT 21.040 27.170 21.210 27.340 ;
        RECT 22.140 27.170 22.310 27.340 ;
        RECT 22.970 27.300 23.140 27.470 ;
        RECT 51.730 27.350 51.900 27.520 ;
        RECT 51.730 26.990 51.900 27.160 ;
        RECT 22.970 26.610 23.140 26.780 ;
        RECT 47.220 26.590 47.390 26.760 ;
        RECT 49.650 26.690 49.820 26.860 ;
        RECT 50.690 26.650 50.860 26.820 ;
        RECT 48.690 26.180 48.900 26.390 ;
        RECT 21.040 25.800 21.210 25.970 ;
        RECT 22.140 25.800 22.310 25.970 ;
        RECT 19.390 25.070 19.560 25.240 ;
        RECT 19.380 23.730 19.550 23.900 ;
        RECT 20.490 25.070 20.660 25.240 ;
        RECT 21.580 25.070 21.750 25.240 ;
        RECT 29.520 24.050 29.690 24.390 ;
        RECT 29.890 24.050 30.060 24.390 ;
        RECT 20.490 23.720 20.660 23.890 ;
        RECT 21.580 23.700 21.750 23.870 ;
        RECT 19.940 23.030 20.110 23.200 ;
        RECT 21.040 23.020 21.210 23.190 ;
        RECT 22.130 23.020 22.300 23.190 ;
        RECT 52.620 21.860 52.790 22.030 ;
        RECT 22.740 20.720 22.910 20.890 ;
        RECT 19.430 20.280 19.600 20.450 ;
        RECT 20.530 20.290 20.700 20.460 ;
        RECT 19.980 19.610 20.150 19.780 ;
        RECT 19.980 18.240 20.150 18.410 ;
        RECT 21.620 20.290 21.790 20.460 ;
        RECT 21.080 19.610 21.250 19.780 ;
        RECT 21.080 18.240 21.250 18.410 ;
        RECT 22.750 20.250 22.920 20.420 ;
        RECT 22.180 19.610 22.350 19.780 ;
        RECT 53.710 21.860 53.880 22.030 ;
        RECT 53.170 21.180 53.340 21.350 ;
        RECT 53.170 19.810 53.340 19.980 ;
        RECT 54.810 21.850 54.980 22.020 ;
        RECT 54.260 21.160 54.430 21.330 ;
        RECT 54.260 19.810 54.430 19.980 ;
        RECT 55.790 21.880 55.960 22.050 ;
        RECT 55.790 21.520 55.960 21.690 ;
        RECT 55.370 21.150 55.540 21.320 ;
        RECT 57.680 21.880 57.850 22.050 ;
        RECT 57.680 21.520 57.850 21.690 ;
        RECT 58.660 21.850 58.830 22.020 ;
        RECT 58.100 21.150 58.270 21.320 ;
        RECT 55.360 19.810 55.530 19.980 ;
        RECT 58.110 19.810 58.280 19.980 ;
        RECT 59.760 21.860 59.930 22.030 ;
        RECT 59.210 21.160 59.380 21.330 ;
        RECT 59.210 19.810 59.380 19.980 ;
        RECT 60.850 21.860 61.020 22.030 ;
        RECT 60.300 21.180 60.470 21.350 ;
        RECT 60.300 19.810 60.470 19.980 ;
        RECT 62.430 21.890 62.600 22.060 ;
        RECT 63.520 21.890 63.690 22.060 ;
        RECT 62.980 21.210 63.150 21.380 ;
        RECT 62.980 19.840 63.150 20.010 ;
        RECT 64.620 21.880 64.790 22.050 ;
        RECT 64.070 21.190 64.240 21.360 ;
        RECT 64.070 19.840 64.240 20.010 ;
        RECT 65.600 21.910 65.770 22.080 ;
        RECT 65.600 21.550 65.770 21.720 ;
        RECT 65.180 21.180 65.350 21.350 ;
        RECT 67.490 21.910 67.660 22.080 ;
        RECT 67.490 21.550 67.660 21.720 ;
        RECT 68.470 21.880 68.640 22.050 ;
        RECT 67.910 21.180 68.080 21.350 ;
        RECT 65.170 19.840 65.340 20.010 ;
        RECT 67.920 19.840 68.090 20.010 ;
        RECT 69.570 21.890 69.740 22.060 ;
        RECT 69.020 21.190 69.190 21.360 ;
        RECT 69.020 19.840 69.190 20.010 ;
        RECT 70.660 21.890 70.830 22.060 ;
        RECT 70.110 21.210 70.280 21.380 ;
        RECT 70.110 19.840 70.280 20.010 ;
        RECT 74.210 21.860 74.380 22.030 ;
        RECT 73.650 21.160 73.820 21.330 ;
        RECT 73.660 19.820 73.830 19.990 ;
        RECT 75.310 21.870 75.480 22.040 ;
        RECT 76.400 21.870 76.570 22.040 ;
        RECT 74.760 21.170 74.930 21.340 ;
        RECT 75.850 21.190 76.020 21.360 ;
        RECT 74.760 19.820 74.930 19.990 ;
        RECT 75.850 19.820 76.020 19.990 ;
        RECT 52.610 19.080 52.780 19.250 ;
        RECT 22.180 18.240 22.350 18.410 ;
        RECT 19.430 17.510 19.600 17.680 ;
        RECT 19.420 16.170 19.590 16.340 ;
        RECT 19.000 15.800 19.170 15.970 ;
        RECT 20.530 17.510 20.700 17.680 ;
        RECT 20.530 16.160 20.700 16.330 ;
        RECT 19.980 15.470 20.150 15.640 ;
        RECT 21.620 17.510 21.790 17.680 ;
        RECT 21.620 16.140 21.790 16.310 ;
        RECT 21.080 15.460 21.250 15.630 ;
        RECT 52.610 17.710 52.780 17.880 ;
        RECT 52.040 17.070 52.210 17.240 ;
        RECT 53.710 19.080 53.880 19.250 ;
        RECT 53.710 17.710 53.880 17.880 ;
        RECT 53.170 17.030 53.340 17.200 ;
        RECT 54.810 19.080 54.980 19.250 ;
        RECT 54.810 17.710 54.980 17.880 ;
        RECT 54.260 17.030 54.430 17.200 ;
        RECT 58.660 19.080 58.830 19.250 ;
        RECT 58.660 17.710 58.830 17.880 ;
        RECT 55.360 17.040 55.530 17.210 ;
        RECT 58.110 17.040 58.280 17.210 ;
        RECT 59.760 19.080 59.930 19.250 ;
        RECT 59.760 17.710 59.930 17.880 ;
        RECT 59.210 17.030 59.380 17.200 ;
        RECT 60.860 19.080 61.030 19.250 ;
        RECT 62.420 19.110 62.590 19.280 ;
        RECT 60.860 17.710 61.030 17.880 ;
        RECT 62.420 17.740 62.590 17.910 ;
        RECT 60.300 17.030 60.470 17.200 ;
        RECT 61.430 17.070 61.600 17.240 ;
        RECT 61.850 17.100 62.020 17.270 ;
        RECT 63.520 19.110 63.690 19.280 ;
        RECT 63.520 17.740 63.690 17.910 ;
        RECT 62.980 17.060 63.150 17.230 ;
        RECT 64.620 19.110 64.790 19.280 ;
        RECT 64.620 17.740 64.790 17.910 ;
        RECT 64.070 17.060 64.240 17.230 ;
        RECT 68.470 19.110 68.640 19.280 ;
        RECT 68.470 17.740 68.640 17.910 ;
        RECT 65.170 17.070 65.340 17.240 ;
        RECT 67.920 17.070 68.090 17.240 ;
        RECT 69.570 19.110 69.740 19.280 ;
        RECT 69.570 17.740 69.740 17.910 ;
        RECT 69.020 17.060 69.190 17.230 ;
        RECT 70.670 19.110 70.840 19.280 ;
        RECT 70.670 17.740 70.840 17.910 ;
        RECT 70.110 17.060 70.280 17.230 ;
        RECT 71.240 17.100 71.410 17.270 ;
        RECT 74.210 19.090 74.380 19.260 ;
        RECT 74.210 17.720 74.380 17.890 ;
        RECT 73.660 17.050 73.830 17.220 ;
        RECT 75.310 19.090 75.480 19.260 ;
        RECT 76.410 19.090 76.580 19.260 ;
        RECT 77.240 18.640 77.410 18.810 ;
        RECT 77.240 18.280 77.410 18.450 ;
        RECT 75.310 17.720 75.480 17.890 ;
        RECT 76.410 17.720 76.580 17.890 ;
        RECT 74.760 17.040 74.930 17.210 ;
        RECT 75.850 17.040 76.020 17.210 ;
        RECT 76.980 17.080 77.150 17.250 ;
        RECT 52.050 16.600 52.220 16.770 ;
        RECT 61.420 16.600 61.590 16.770 ;
        RECT 61.860 16.630 62.030 16.800 ;
        RECT 71.230 16.630 71.400 16.800 ;
        RECT 76.970 16.610 77.140 16.780 ;
        RECT 22.170 15.460 22.340 15.630 ;
        RECT 23.710 12.080 23.880 15.600 ;
        RECT 24.070 12.080 24.240 15.600 ;
        RECT 24.430 12.080 24.600 15.600 ;
        RECT 25.120 12.080 25.290 15.600 ;
        RECT 25.480 12.080 25.650 15.600 ;
        RECT 25.840 12.080 26.010 15.600 ;
        RECT 102.550 14.410 102.720 14.580 ;
        RECT 108.140 13.710 108.310 13.880 ;
        RECT 108.140 13.040 108.310 13.210 ;
        RECT 102.550 12.800 102.720 12.970 ;
        RECT 102.550 11.200 102.720 11.370 ;
        RECT 102.550 9.580 102.720 9.750 ;
        RECT 107.560 8.370 107.730 8.540 ;
        RECT 102.550 7.980 102.720 8.150 ;
        RECT 102.550 6.360 102.720 6.530 ;
        RECT 102.550 4.760 102.720 4.930 ;
        RECT 114.080 4.870 114.250 19.820 ;
        RECT 102.550 3.140 102.720 3.310 ;
      LAYER met1 ;
        RECT 85.630 76.420 85.970 76.560 ;
        RECT 93.510 76.420 94.230 78.160 ;
        RECT 85.630 75.700 94.230 76.420 ;
        RECT 33.560 73.250 34.900 73.700 ;
        RECT 7.460 72.410 7.960 72.890 ;
        RECT 33.560 72.830 47.080 73.250 ;
        RECT 48.870 73.160 52.060 74.280 ;
        RECT 0.420 72.030 0.660 72.390 ;
        RECT 7.560 69.450 7.950 72.410 ;
        RECT 15.110 72.000 15.370 72.790 ;
        RECT 19.810 71.950 20.070 72.740 ;
        RECT 33.560 72.690 34.900 72.830 ;
        RECT 28.150 72.090 30.920 72.330 ;
        RECT 28.150 71.680 28.390 72.090 ;
        RECT 1.000 69.040 1.260 69.340 ;
        RECT 3.860 69.200 4.120 69.390 ;
        RECT 3.860 69.070 4.230 69.200 ;
        RECT 1.000 69.020 1.410 69.040 ;
        RECT 1.030 68.730 1.410 69.020 ;
        RECT 2.440 68.730 3.470 69.040 ;
        RECT 3.940 68.970 4.230 69.070 ;
        RECT 0.990 68.170 1.250 68.310 ;
        RECT 0.990 67.990 1.340 68.170 ;
        RECT 1.630 68.010 1.950 68.330 ;
        RECT 2.400 68.170 2.660 68.320 ;
        RECT 2.400 68.000 2.740 68.170 ;
        RECT 1.100 67.940 1.340 67.990 ;
        RECT 2.510 67.940 2.740 68.000 ;
        RECT 1.040 67.860 2.790 67.940 ;
        RECT 0.990 67.540 2.790 67.860 ;
        RECT 1.040 67.440 2.790 67.540 ;
        RECT 0.990 67.280 2.790 67.440 ;
        RECT 0.990 67.120 1.340 67.280 ;
        RECT 1.630 67.170 1.950 67.280 ;
        RECT 2.420 67.140 2.740 67.280 ;
        RECT 1.100 67.060 1.340 67.120 ;
        RECT 2.510 67.060 2.740 67.140 ;
        RECT 1.100 66.090 1.330 66.510 ;
        RECT 0.990 65.770 1.330 66.090 ;
        RECT 1.100 65.100 1.330 65.770 ;
        RECT 2.510 65.100 2.740 66.510 ;
        RECT 3.230 66.330 3.470 68.730 ;
        RECT 7.560 68.960 8.030 69.450 ;
        RECT 7.560 68.950 8.010 68.960 ;
        RECT 14.100 68.950 14.340 69.590 ;
        RECT 15.110 69.010 15.370 69.800 ;
        RECT 19.310 69.030 19.550 69.440 ;
        RECT 3.950 68.280 4.220 68.410 ;
        RECT 3.630 68.050 4.310 68.280 ;
        RECT 3.520 67.690 3.840 68.010 ;
        RECT 3.890 67.990 4.310 68.050 ;
        RECT 3.570 67.460 3.800 67.690 ;
        RECT 4.080 67.050 4.310 67.990 ;
        RECT 3.950 66.870 4.310 67.050 ;
        RECT 3.950 66.850 4.220 66.870 ;
        RECT 3.630 66.620 4.220 66.850 ;
        RECT 3.140 66.040 3.470 66.330 ;
        RECT 3.230 65.960 3.470 66.040 ;
        RECT 3.330 65.270 3.650 65.590 ;
        RECT 3.950 65.580 4.220 66.620 ;
        RECT 3.950 65.350 4.280 65.580 ;
        RECT 1.610 64.370 1.930 64.690 ;
        RECT 3.040 64.390 3.360 64.710 ;
        RECT 0.820 63.790 1.140 64.110 ;
        RECT 1.750 63.790 2.070 64.110 ;
        RECT 2.450 63.790 2.770 64.110 ;
        RECT 3.190 63.790 3.510 64.110 ;
        RECT 3.900 63.780 4.220 64.100 ;
        RECT 5.940 63.390 6.230 64.450 ;
        RECT 7.560 10.840 7.950 68.950 ;
        RECT 14.100 68.690 14.330 68.950 ;
        RECT 14.090 68.470 14.330 68.690 ;
        RECT 8.970 67.810 9.230 68.130 ;
        RECT 15.110 68.000 15.370 68.790 ;
        RECT 25.150 68.190 25.420 69.440 ;
        RECT 29.860 68.550 30.120 69.440 ;
        RECT 8.980 65.590 9.220 67.810 ;
        RECT 17.020 67.270 17.340 67.590 ;
        RECT 18.380 67.350 18.700 67.670 ;
        RECT 19.070 67.340 19.390 67.660 ;
        RECT 14.100 66.150 14.340 66.790 ;
        RECT 14.100 65.890 14.330 66.150 ;
        RECT 14.090 65.670 14.330 65.890 ;
        RECT 8.890 65.110 9.310 65.590 ;
        RECT 14.100 64.600 14.340 65.240 ;
        RECT 14.100 64.340 14.330 64.600 ;
        RECT 14.780 64.350 15.070 66.270 ;
        RECT 14.090 64.120 14.330 64.340 ;
        RECT 14.760 63.680 15.170 64.350 ;
        RECT 16.300 63.610 16.620 63.930 ;
        RECT 19.300 63.390 19.540 65.270 ;
        RECT 25.120 63.390 25.430 65.980 ;
        RECT 26.160 63.630 26.480 63.950 ;
        RECT 28.140 62.990 28.380 66.220 ;
        RECT 28.470 64.750 28.700 66.040 ;
        RECT 29.080 63.570 29.330 65.440 ;
        RECT 29.080 63.390 29.340 63.570 ;
        RECT 28.090 62.650 28.430 62.990 ;
        RECT 25.340 62.550 25.830 62.560 ;
        RECT 22.520 58.970 22.840 59.290 ;
        RECT 23.610 58.980 23.930 59.300 ;
        RECT 20.980 58.060 21.300 58.380 ;
        RECT 22.530 57.980 22.850 58.300 ;
        RECT 20.960 57.140 21.280 57.460 ;
        RECT 20.940 56.150 21.260 56.470 ;
        RECT 21.410 53.860 21.640 57.340 ;
        RECT 22.080 56.720 22.300 57.340 ;
        RECT 22.530 56.990 22.850 57.310 ;
        RECT 22.050 56.400 22.310 56.720 ;
        RECT 22.080 55.840 22.300 56.400 ;
        RECT 22.440 56.260 22.760 56.580 ;
        RECT 22.530 55.840 22.850 55.880 ;
        RECT 22.080 55.800 22.850 55.840 ;
        RECT 22.020 55.610 22.850 55.800 ;
        RECT 22.020 55.480 22.300 55.610 ;
        RECT 22.530 55.590 22.850 55.610 ;
        RECT 22.080 54.880 22.300 55.480 ;
        RECT 22.440 55.560 22.850 55.590 ;
        RECT 22.440 55.270 22.760 55.560 ;
        RECT 22.030 54.850 22.300 54.880 ;
        RECT 22.530 54.850 22.850 54.890 ;
        RECT 22.030 54.620 22.850 54.850 ;
        RECT 22.030 54.560 22.300 54.620 ;
        RECT 22.530 54.600 22.850 54.620 ;
        RECT 21.380 53.540 21.640 53.860 ;
        RECT 21.410 52.900 21.640 53.540 ;
        RECT 21.340 52.580 21.640 52.900 ;
        RECT 21.410 51.940 21.640 52.580 ;
        RECT 21.380 51.620 21.640 51.940 ;
        RECT 21.410 36.870 21.640 51.620 ;
        RECT 22.080 53.860 22.300 54.560 ;
        RECT 22.440 54.570 22.850 54.600 ;
        RECT 22.440 54.280 22.760 54.570 ;
        RECT 22.860 54.170 23.080 58.780 ;
        RECT 22.840 54.100 23.080 54.170 ;
        RECT 23.260 58.230 23.480 58.780 ;
        RECT 23.260 57.940 23.580 58.230 ;
        RECT 23.620 57.990 23.940 58.310 ;
        RECT 22.840 54.000 23.180 54.100 ;
        RECT 22.530 53.860 22.850 53.900 ;
        RECT 22.080 53.630 22.850 53.860 ;
        RECT 22.080 36.870 22.300 53.630 ;
        RECT 22.530 53.580 22.850 53.630 ;
        RECT 22.860 53.870 23.180 54.000 ;
        RECT 22.860 52.900 23.080 53.870 ;
        RECT 23.260 52.900 23.480 57.940 ;
        RECT 23.620 57.000 23.940 57.320 ;
        RECT 24.770 57.060 24.990 61.610 ;
        RECT 25.330 61.400 25.840 62.550 ;
        RECT 30.680 61.620 30.920 72.090 ;
        RECT 33.990 71.760 37.020 72.030 ;
        RECT 38.700 71.770 38.960 72.830 ;
        RECT 33.960 62.590 34.270 66.290 ;
        RECT 33.880 62.220 34.270 62.590 ;
        RECT 36.750 62.080 37.020 71.760 ;
        RECT 46.660 69.580 47.080 72.830 ;
        RECT 50.470 70.340 50.890 73.160 ;
        RECT 50.470 69.860 50.940 70.340 ;
        RECT 46.620 69.100 47.100 69.580 ;
        RECT 52.170 67.490 52.610 67.990 ;
        RECT 57.890 67.490 58.330 67.990 ;
        RECT 47.750 66.470 48.190 66.970 ;
        RECT 37.920 63.080 38.170 66.230 ;
        RECT 44.960 63.730 45.280 63.780 ;
        RECT 44.870 63.440 45.280 63.730 ;
        RECT 37.880 62.720 38.210 63.080 ;
        RECT 44.450 62.440 44.690 62.510 ;
        RECT 36.710 61.770 37.050 62.080 ;
        RECT 44.480 62.020 44.720 62.070 ;
        RECT 25.280 61.300 25.840 61.400 ;
        RECT 30.630 61.300 30.970 61.620 ;
        RECT 25.170 60.900 25.840 61.300 ;
        RECT 25.170 60.870 25.830 60.900 ;
        RECT 25.170 57.060 25.390 60.870 ;
        RECT 44.450 60.690 44.690 60.760 ;
        RECT 44.870 59.940 45.110 63.440 ;
        RECT 47.230 62.510 47.470 62.930 ;
        RECT 47.230 62.450 47.700 62.510 ;
        RECT 47.230 62.070 47.470 62.450 ;
        RECT 47.230 62.010 47.730 62.070 ;
        RECT 46.490 61.430 46.900 61.760 ;
        RECT 47.230 61.250 47.470 62.010 ;
        RECT 47.230 60.760 47.470 61.180 ;
        RECT 47.230 60.700 47.700 60.760 ;
        RECT 46.490 59.680 46.900 60.010 ;
        RECT 47.230 59.500 47.470 60.700 ;
        RECT 47.810 59.870 48.120 66.470 ;
        RECT 48.650 62.290 49.000 62.580 ;
        RECT 48.650 62.270 48.850 62.290 ;
        RECT 49.610 62.080 49.920 62.090 ;
        RECT 49.610 61.810 49.930 62.080 ;
        RECT 49.630 61.800 49.920 61.810 ;
        RECT 50.170 61.250 50.480 62.940 ;
        RECT 50.650 61.870 50.970 62.150 ;
        RECT 51.720 62.070 52.010 62.510 ;
        RECT 51.720 61.980 52.040 62.070 ;
        RECT 50.650 61.850 51.010 61.870 ;
        RECT 50.730 61.540 51.010 61.850 ;
        RECT 48.650 60.540 49.000 60.830 ;
        RECT 48.650 60.520 48.850 60.540 ;
        RECT 49.610 60.330 49.920 60.340 ;
        RECT 49.610 60.060 49.930 60.330 ;
        RECT 49.630 60.050 49.920 60.060 ;
        RECT 50.170 59.500 50.480 61.190 ;
        RECT 50.650 60.120 50.970 60.400 ;
        RECT 50.650 60.100 51.010 60.120 ;
        RECT 50.730 59.790 51.010 60.100 ;
        RECT 26.390 58.750 26.740 59.210 ;
        RECT 42.820 58.770 43.190 59.080 ;
        RECT 47.230 59.010 47.470 59.430 ;
        RECT 44.450 58.940 44.690 59.010 ;
        RECT 47.230 58.950 47.700 59.010 ;
        RECT 25.790 58.390 26.040 58.510 ;
        RECT 25.760 57.930 26.080 58.390 ;
        RECT 25.790 57.140 26.040 57.930 ;
        RECT 25.790 56.820 26.080 57.140 ;
        RECT 23.740 56.160 24.060 56.480 ;
        RECT 25.790 56.220 26.040 56.820 ;
        RECT 25.790 55.900 26.080 56.220 ;
        RECT 23.740 55.170 24.060 55.490 ;
        RECT 25.790 55.300 26.040 55.900 ;
        RECT 25.790 54.980 26.050 55.300 ;
        RECT 23.740 54.180 24.060 54.500 ;
        RECT 21.300 36.340 21.640 36.870 ;
        RECT 21.960 36.340 22.300 36.870 ;
        RECT 19.990 35.600 20.220 35.670 ;
        RECT 19.950 35.340 20.270 35.600 ;
        RECT 19.500 35.230 19.730 35.270 ;
        RECT 19.460 34.910 19.730 35.230 ;
        RECT 10.150 33.670 10.870 34.370 ;
        RECT 10.160 28.520 10.820 33.670 ;
        RECT 19.500 31.390 19.730 34.910 ;
        RECT 19.990 32.870 20.220 35.340 ;
        RECT 21.410 35.250 21.640 36.340 ;
        RECT 22.080 35.610 22.300 36.340 ;
        RECT 23.840 35.630 24.110 35.670 ;
        RECT 22.060 35.290 22.320 35.610 ;
        RECT 23.820 35.300 24.110 35.630 ;
        RECT 21.400 34.930 21.660 35.250 ;
        RECT 23.290 33.760 23.580 33.790 ;
        RECT 19.990 32.500 20.720 32.870 ;
        RECT 19.500 31.320 19.760 31.390 ;
        RECT 19.480 31.310 19.760 31.320 ;
        RECT 19.450 31.000 19.770 31.310 ;
        RECT 15.350 29.140 15.780 29.570 ;
        RECT 10.160 27.800 10.900 28.520 ;
        RECT 15.400 23.330 15.770 29.140 ;
        RECT 19.310 27.760 19.630 28.080 ;
        RECT 19.990 27.410 20.220 32.500 ;
        RECT 23.840 32.330 24.110 35.300 ;
        RECT 23.720 32.080 24.110 32.330 ;
        RECT 24.320 35.230 24.560 35.270 ;
        RECT 24.320 34.910 24.580 35.230 ;
        RECT 24.320 31.770 24.560 34.910 ;
        RECT 23.720 31.540 24.560 31.770 ;
        RECT 22.620 28.200 22.940 28.520 ;
        RECT 20.410 27.770 20.730 28.090 ;
        RECT 21.500 27.770 21.820 28.090 ;
        RECT 22.630 27.730 22.950 28.050 ;
        RECT 19.860 27.090 20.220 27.410 ;
        RECT 20.960 27.090 21.280 27.410 ;
        RECT 22.060 27.090 22.380 27.410 ;
        RECT 19.990 26.040 20.220 27.090 ;
        RECT 22.910 27.070 23.200 27.500 ;
        RECT 22.910 27.050 23.380 27.070 ;
        RECT 22.920 26.750 23.380 27.050 ;
        RECT 22.920 26.220 23.200 26.750 ;
        RECT 22.930 26.190 23.200 26.220 ;
        RECT 19.860 25.720 20.220 26.040 ;
        RECT 20.960 25.720 21.280 26.040 ;
        RECT 22.060 25.720 22.380 26.040 ;
        RECT 19.310 24.990 19.630 25.310 ;
        RECT 19.990 25.000 20.220 25.720 ;
        RECT 20.410 25.000 20.730 25.310 ;
        RECT 21.500 25.000 21.820 25.310 ;
        RECT 19.990 24.770 22.440 25.000 ;
        RECT 22.120 24.440 22.440 24.770 ;
        RECT 19.300 23.650 19.620 23.970 ;
        RECT 20.410 23.640 20.730 23.960 ;
        RECT 21.500 23.620 21.820 23.940 ;
        RECT 15.360 22.900 15.790 23.330 ;
        RECT 19.860 22.950 20.180 23.270 ;
        RECT 20.960 22.940 21.280 23.260 ;
        RECT 22.050 22.940 22.370 23.260 ;
        RECT 22.880 22.870 23.210 22.900 ;
        RECT 22.740 22.790 23.210 22.870 ;
        RECT 22.500 22.550 23.210 22.790 ;
        RECT 22.880 22.480 23.210 22.550 ;
        RECT 18.370 17.240 18.660 17.590 ;
        RECT 18.380 16.670 18.640 17.240 ;
        RECT 19.020 16.140 19.280 21.120 ;
        RECT 22.660 20.640 22.980 20.960 ;
        RECT 19.350 20.200 19.670 20.520 ;
        RECT 20.450 20.210 20.770 20.530 ;
        RECT 21.540 20.210 21.860 20.530 ;
        RECT 22.670 20.170 22.990 20.490 ;
        RECT 19.900 19.530 20.220 19.850 ;
        RECT 21.000 19.530 21.320 19.850 ;
        RECT 22.100 19.530 22.420 19.850 ;
        RECT 19.900 18.160 20.220 18.480 ;
        RECT 21.000 18.160 21.320 18.480 ;
        RECT 22.100 18.160 22.420 18.480 ;
        RECT 19.350 17.430 19.670 17.750 ;
        RECT 20.450 17.430 20.770 17.750 ;
        RECT 21.540 17.430 21.860 17.750 ;
        RECT 24.320 16.880 24.560 31.540 ;
        RECT 24.770 30.870 24.990 51.620 ;
        RECT 25.170 33.480 25.390 51.620 ;
        RECT 25.790 34.630 26.040 54.980 ;
        RECT 26.410 54.210 26.670 58.750 ;
        RECT 42.180 57.050 42.570 57.420 ;
        RECT 41.600 55.560 41.990 55.950 ;
        RECT 26.410 53.890 26.690 54.210 ;
        RECT 40.960 53.970 41.350 54.350 ;
        RECT 40.990 53.960 41.330 53.970 ;
        RECT 26.410 53.250 26.670 53.890 ;
        RECT 40.350 53.770 40.690 53.780 ;
        RECT 40.340 53.380 40.700 53.770 ;
        RECT 26.410 52.930 26.700 53.250 ;
        RECT 26.410 52.290 26.670 52.930 ;
        RECT 26.410 51.970 26.690 52.290 ;
        RECT 25.790 34.610 26.050 34.630 ;
        RECT 25.780 34.330 26.060 34.610 ;
        RECT 25.790 34.310 26.050 34.330 ;
        RECT 25.130 33.160 25.450 33.480 ;
        RECT 25.170 31.570 25.390 33.160 ;
        RECT 25.790 32.870 26.040 34.310 ;
        RECT 25.710 32.550 26.040 32.870 ;
        RECT 25.170 31.250 25.500 31.570 ;
        RECT 25.170 31.090 25.390 31.250 ;
        RECT 25.070 30.890 25.390 31.090 ;
        RECT 24.730 30.550 25.010 30.870 ;
        RECT 25.070 30.580 25.490 30.890 ;
        RECT 24.770 17.580 24.990 30.550 ;
        RECT 25.170 30.380 25.490 30.580 ;
        RECT 25.170 30.020 25.390 30.380 ;
        RECT 25.170 29.700 25.500 30.020 ;
        RECT 25.170 25.340 25.390 29.700 ;
        RECT 25.790 28.990 26.040 32.550 ;
        RECT 26.410 32.870 26.670 51.970 ;
        RECT 39.730 51.820 40.090 52.210 ;
        RECT 39.080 50.280 39.490 50.680 ;
        RECT 38.550 48.720 38.910 49.110 ;
        RECT 37.970 43.660 38.300 43.680 ;
        RECT 37.910 43.240 38.300 43.660 ;
        RECT 37.340 42.050 37.670 42.070 ;
        RECT 37.290 41.660 37.680 42.050 ;
        RECT 36.720 40.500 37.050 40.510 ;
        RECT 36.690 40.110 37.050 40.500 ;
        RECT 36.070 38.630 36.460 39.030 ;
        RECT 35.400 33.460 35.830 33.860 ;
        RECT 26.930 32.990 27.250 33.310 ;
        RECT 27.580 32.990 27.900 33.310 ;
        RECT 26.410 32.550 26.730 32.870 ;
        RECT 26.410 30.300 26.670 32.550 ;
        RECT 27.960 31.690 28.250 32.600 ;
        RECT 34.740 31.890 35.150 32.290 ;
        RECT 27.610 31.030 27.930 31.070 ;
        RECT 27.610 30.800 28.160 31.030 ;
        RECT 28.420 30.890 28.430 31.120 ;
        RECT 27.610 30.750 27.930 30.800 ;
        RECT 27.620 30.490 27.940 30.530 ;
        RECT 26.400 29.980 26.710 30.300 ;
        RECT 27.620 30.260 28.170 30.490 ;
        RECT 27.620 30.210 27.940 30.260 ;
        RECT 34.130 30.250 34.520 30.650 ;
        RECT 25.740 28.670 26.060 28.990 ;
        RECT 26.410 28.980 26.670 29.980 ;
        RECT 27.950 29.670 28.220 29.850 ;
        RECT 27.930 29.350 28.250 29.670 ;
        RECT 27.950 29.180 28.220 29.350 ;
        RECT 25.170 24.860 25.460 25.340 ;
        RECT 25.170 22.900 25.390 24.860 ;
        RECT 25.150 22.480 25.410 22.900 ;
        RECT 25.170 17.860 25.390 22.480 ;
        RECT 25.790 19.240 26.040 28.670 ;
        RECT 26.410 28.660 26.750 28.980 ;
        RECT 33.440 28.810 33.850 29.200 ;
        RECT 25.750 18.840 26.050 19.240 ;
        RECT 25.170 17.720 25.410 17.860 ;
        RECT 24.730 17.230 25.040 17.580 ;
        RECT 25.180 17.090 25.410 17.720 ;
        RECT 18.970 15.330 19.280 16.140 ;
        RECT 19.340 16.090 19.660 16.410 ;
        RECT 20.450 16.080 20.770 16.400 ;
        RECT 21.540 16.060 21.860 16.380 ;
        RECT 23.530 16.320 24.560 16.880 ;
        RECT 25.170 17.060 25.410 17.090 ;
        RECT 23.530 16.210 24.320 16.320 ;
        RECT 19.900 15.390 20.220 15.710 ;
        RECT 21.000 15.380 21.320 15.700 ;
        RECT 22.090 15.380 22.410 15.700 ;
        RECT 25.170 15.670 25.390 17.060 ;
        RECT 19.020 15.130 19.280 15.330 ;
        RECT 23.640 11.990 26.060 15.670 ;
        RECT 26.410 11.700 26.670 28.660 ;
        RECT 26.910 27.890 27.230 28.210 ;
        RECT 27.620 27.830 27.940 28.150 ;
        RECT 29.230 23.660 30.160 25.310 ;
        RECT 29.320 23.180 30.060 23.660 ;
        RECT 26.320 11.290 26.670 11.700 ;
        RECT 7.390 10.320 7.950 10.840 ;
        RECT 33.500 5.470 33.830 28.810 ;
        RECT 33.450 5.460 33.880 5.470 ;
        RECT 33.420 5.000 33.910 5.460 ;
        RECT 33.450 4.980 33.880 5.000 ;
        RECT 34.150 4.680 34.480 30.250 ;
        RECT 34.060 4.190 34.550 4.680 ;
        RECT 34.800 3.970 35.130 31.890 ;
        RECT 34.770 3.510 35.170 3.970 ;
        RECT 34.560 3.020 35.140 3.130 ;
        RECT 35.470 3.020 35.800 33.460 ;
        RECT 36.110 7.600 36.440 38.630 ;
        RECT 36.110 3.140 36.430 7.600 ;
        RECT 36.720 3.750 37.050 40.110 ;
        RECT 37.340 4.000 37.670 41.660 ;
        RECT 37.970 5.030 38.300 43.240 ;
        RECT 38.570 5.330 38.900 48.720 ;
        RECT 39.150 5.900 39.480 50.280 ;
        RECT 39.760 6.930 40.090 51.820 ;
        RECT 40.350 7.540 40.680 53.380 ;
        RECT 40.990 8.210 41.320 53.960 ;
        RECT 41.610 8.860 41.940 55.560 ;
        RECT 42.210 9.490 42.540 57.050 ;
        RECT 42.840 10.100 43.170 58.770 ;
        RECT 46.490 57.930 46.900 58.260 ;
        RECT 47.230 57.750 47.470 58.950 ;
        RECT 48.650 58.790 49.000 59.080 ;
        RECT 48.650 58.770 48.850 58.790 ;
        RECT 49.610 58.580 49.920 58.590 ;
        RECT 49.610 58.310 49.930 58.580 ;
        RECT 49.630 58.300 49.920 58.310 ;
        RECT 50.170 57.750 50.480 59.440 ;
        RECT 50.650 58.370 50.970 58.650 ;
        RECT 50.650 58.350 51.010 58.370 ;
        RECT 50.730 58.040 51.010 58.350 ;
        RECT 47.230 57.260 47.470 57.680 ;
        RECT 44.450 57.190 44.690 57.260 ;
        RECT 47.230 57.200 47.700 57.260 ;
        RECT 46.490 56.180 46.900 56.510 ;
        RECT 47.230 56.000 47.470 57.200 ;
        RECT 48.650 57.040 49.000 57.330 ;
        RECT 48.650 57.020 48.850 57.040 ;
        RECT 49.610 56.830 49.920 56.840 ;
        RECT 49.610 56.560 49.930 56.830 ;
        RECT 49.630 56.550 49.920 56.560 ;
        RECT 50.170 56.000 50.480 57.690 ;
        RECT 50.650 56.620 50.970 56.900 ;
        RECT 50.650 56.600 51.010 56.620 ;
        RECT 50.730 56.290 51.010 56.600 ;
        RECT 51.720 55.510 52.010 61.980 ;
        RECT 52.240 59.890 52.530 67.490 ;
        RECT 53.430 66.500 53.930 66.940 ;
        RECT 44.480 55.070 44.720 55.120 ;
        RECT 47.420 55.070 47.730 55.130 ;
        RECT 51.750 55.070 52.040 55.190 ;
        RECT 44.970 53.900 45.210 54.010 ;
        RECT 47.910 53.900 48.220 54.010 ;
        RECT 52.240 53.860 52.530 54.020 ;
        RECT 53.700 53.500 53.890 66.500 ;
        RECT 57.980 53.460 58.230 67.490 ;
        RECT 59.680 67.450 60.410 74.320 ;
        RECT 64.830 74.170 65.810 74.320 ;
        RECT 59.840 57.060 60.010 67.450 ;
        RECT 64.840 66.920 65.810 74.170 ;
        RECT 77.460 73.150 80.650 74.270 ;
        RECT 70.230 69.080 71.700 69.610 ;
        RECT 64.820 66.450 65.830 66.920 ;
        RECT 67.860 66.470 68.300 66.970 ;
        RECT 62.060 62.720 62.400 63.010 ;
        RECT 62.110 62.690 62.370 62.720 ;
        RECT 60.230 59.160 60.490 59.480 ;
        RECT 60.260 56.930 60.450 59.160 ;
        RECT 62.130 56.910 62.340 62.690 ;
        RECT 65.700 62.090 65.960 62.100 ;
        RECT 65.680 61.790 65.980 62.090 ;
        RECT 65.700 61.780 65.960 61.790 ;
        RECT 62.530 60.760 62.870 61.080 ;
        RECT 62.600 56.930 62.790 60.760 ;
        RECT 62.970 58.670 63.260 58.990 ;
        RECT 63.010 56.910 63.220 58.670 ;
        RECT 64.010 58.190 64.350 58.510 ;
        RECT 64.090 56.940 64.270 58.190 ;
        RECT 65.730 53.700 65.930 61.780 ;
        RECT 67.960 56.890 68.190 66.470 ;
        RECT 68.860 62.700 69.140 63.020 ;
        RECT 68.420 61.790 68.700 62.110 ;
        RECT 64.200 53.630 64.390 53.700 ;
        RECT 65.510 53.620 65.930 53.700 ;
        RECT 61.880 53.310 62.070 53.530 ;
        RECT 44.480 52.790 44.720 52.840 ;
        RECT 47.420 52.780 47.730 52.840 ;
        RECT 51.750 52.720 52.040 52.840 ;
        RECT 61.600 52.820 62.070 53.310 ;
        RECT 62.460 53.170 62.830 53.190 ;
        RECT 62.410 52.910 62.830 53.170 ;
        RECT 62.460 52.900 62.830 52.910 ;
        RECT 46.490 51.400 46.900 51.730 ;
        RECT 44.450 50.650 44.690 50.720 ;
        RECT 47.230 50.710 47.470 51.910 ;
        RECT 49.630 51.350 49.920 51.360 ;
        RECT 49.610 51.080 49.930 51.350 ;
        RECT 49.610 51.070 49.920 51.080 ;
        RECT 48.650 50.870 48.850 50.890 ;
        RECT 47.230 50.650 47.700 50.710 ;
        RECT 47.230 50.230 47.470 50.650 ;
        RECT 48.650 50.580 49.000 50.870 ;
        RECT 50.170 50.220 50.480 51.910 ;
        RECT 50.730 51.310 51.010 51.620 ;
        RECT 50.650 51.290 51.010 51.310 ;
        RECT 50.650 51.010 50.970 51.290 ;
        RECT 46.490 49.650 46.900 49.980 ;
        RECT 44.450 48.900 44.690 48.970 ;
        RECT 47.230 48.960 47.470 50.160 ;
        RECT 49.630 49.600 49.920 49.610 ;
        RECT 49.610 49.330 49.930 49.600 ;
        RECT 49.610 49.320 49.920 49.330 ;
        RECT 48.650 49.120 48.850 49.140 ;
        RECT 47.230 48.900 47.700 48.960 ;
        RECT 47.230 48.480 47.470 48.900 ;
        RECT 48.650 48.830 49.000 49.120 ;
        RECT 50.170 48.470 50.480 50.160 ;
        RECT 50.730 49.560 51.010 49.870 ;
        RECT 50.650 49.540 51.010 49.560 ;
        RECT 50.650 49.260 50.970 49.540 ;
        RECT 46.490 47.900 46.900 48.230 ;
        RECT 44.450 47.150 44.690 47.220 ;
        RECT 44.480 45.840 44.720 45.890 ;
        RECT 44.450 45.400 44.690 45.470 ;
        RECT 44.870 43.490 45.110 47.860 ;
        RECT 47.230 47.210 47.470 48.410 ;
        RECT 47.230 47.150 47.700 47.210 ;
        RECT 47.230 46.730 47.470 47.150 ;
        RECT 46.490 46.150 46.900 46.480 ;
        RECT 47.230 45.900 47.470 46.660 ;
        RECT 47.230 45.840 47.730 45.900 ;
        RECT 47.230 45.460 47.470 45.840 ;
        RECT 47.230 45.400 47.700 45.460 ;
        RECT 47.230 44.980 47.470 45.400 ;
        RECT 47.810 43.420 48.120 47.930 ;
        RECT 49.630 47.850 49.920 47.860 ;
        RECT 49.610 47.580 49.930 47.850 ;
        RECT 49.610 47.570 49.920 47.580 ;
        RECT 48.650 47.370 48.850 47.390 ;
        RECT 48.650 47.080 49.000 47.370 ;
        RECT 50.170 46.720 50.480 48.410 ;
        RECT 50.730 47.810 51.010 48.120 ;
        RECT 50.650 47.790 51.010 47.810 ;
        RECT 50.650 47.510 50.970 47.790 ;
        RECT 49.630 46.100 49.920 46.110 ;
        RECT 49.610 45.830 49.930 46.100 ;
        RECT 49.610 45.820 49.920 45.830 ;
        RECT 48.650 45.620 48.850 45.640 ;
        RECT 48.650 45.330 49.000 45.620 ;
        RECT 50.170 44.970 50.480 46.660 ;
        RECT 50.730 46.060 51.010 46.370 ;
        RECT 50.650 46.040 51.010 46.060 ;
        RECT 50.650 45.760 50.970 46.040 ;
        RECT 51.720 45.930 52.010 52.400 ;
        RECT 61.420 52.380 61.740 52.660 ;
        RECT 61.880 52.480 62.070 52.820 ;
        RECT 61.420 52.010 61.740 52.290 ;
        RECT 61.780 52.190 62.070 52.480 ;
        RECT 61.880 51.850 62.070 52.190 ;
        RECT 61.600 51.360 62.070 51.850 ;
        RECT 62.460 51.760 62.830 51.770 ;
        RECT 62.410 51.500 62.830 51.760 ;
        RECT 62.460 51.480 62.830 51.500 ;
        RECT 61.880 51.140 62.070 51.360 ;
        RECT 63.190 51.140 63.420 53.530 ;
        RECT 64.920 53.150 65.260 53.200 ;
        RECT 64.920 53.130 65.480 53.150 ;
        RECT 64.800 52.960 65.480 53.130 ;
        RECT 64.920 52.920 65.480 52.960 ;
        RECT 64.920 52.880 65.260 52.920 ;
        RECT 64.920 51.750 65.260 51.790 ;
        RECT 64.920 51.710 65.480 51.750 ;
        RECT 64.800 51.540 65.480 51.710 ;
        RECT 65.730 51.550 65.930 53.620 ;
        RECT 64.920 51.520 65.480 51.540 ;
        RECT 64.920 51.470 65.260 51.520 ;
        RECT 65.710 51.420 65.930 51.550 ;
        RECT 66.160 53.310 66.410 53.530 ;
        RECT 65.660 51.090 65.990 51.420 ;
        RECT 66.160 51.360 66.800 53.310 ;
        RECT 68.450 52.340 68.670 61.790 ;
        RECT 68.450 52.330 68.730 52.340 ;
        RECT 66.160 51.140 66.410 51.360 ;
        RECT 68.190 50.980 68.200 51.140 ;
        RECT 61.880 50.110 62.070 50.330 ;
        RECT 61.600 49.620 62.070 50.110 ;
        RECT 62.460 49.970 62.830 49.990 ;
        RECT 62.410 49.710 62.830 49.970 ;
        RECT 62.460 49.700 62.830 49.710 ;
        RECT 61.420 49.180 61.740 49.460 ;
        RECT 61.880 49.280 62.070 49.620 ;
        RECT 61.420 48.810 61.740 49.090 ;
        RECT 61.780 48.990 62.070 49.280 ;
        RECT 61.880 48.650 62.070 48.990 ;
        RECT 61.600 48.160 62.070 48.650 ;
        RECT 62.460 48.560 62.830 48.570 ;
        RECT 62.410 48.300 62.830 48.560 ;
        RECT 62.460 48.280 62.830 48.300 ;
        RECT 61.880 47.940 62.070 48.160 ;
        RECT 63.190 47.940 63.420 50.330 ;
        RECT 66.160 50.110 66.410 50.330 ;
        RECT 68.450 50.250 68.670 52.330 ;
        RECT 68.440 50.180 68.670 50.250 ;
        RECT 64.920 49.950 65.260 50.000 ;
        RECT 64.920 49.930 65.480 49.950 ;
        RECT 64.800 49.760 65.480 49.930 ;
        RECT 64.920 49.720 65.480 49.760 ;
        RECT 64.920 49.680 65.260 49.720 ;
        RECT 64.920 48.550 65.260 48.590 ;
        RECT 64.920 48.510 65.480 48.550 ;
        RECT 64.800 48.340 65.480 48.510 ;
        RECT 64.920 48.320 65.480 48.340 ;
        RECT 64.920 48.270 65.260 48.320 ;
        RECT 66.160 48.160 66.800 50.110 ;
        RECT 68.430 49.580 68.630 50.180 ;
        RECT 68.880 49.730 69.110 62.700 ;
        RECT 70.250 56.700 70.670 69.080 ;
        RECT 71.280 56.700 71.700 69.080 ;
        RECT 73.660 66.430 74.100 66.930 ;
        RECT 73.760 59.450 73.990 66.430 ;
        RECT 78.180 61.180 79.460 73.150 ;
        RECT 81.940 67.960 82.220 68.080 ;
        RECT 81.940 67.460 82.270 67.960 ;
        RECT 78.180 61.100 79.480 61.180 ;
        RECT 78.170 60.800 79.480 61.100 ;
        RECT 74.950 60.150 75.250 60.470 ;
        RECT 73.630 59.440 73.990 59.450 ;
        RECT 73.600 58.550 73.990 59.440 ;
        RECT 73.760 56.890 73.990 58.550 ;
        RECT 74.980 56.890 75.210 60.150 ;
        RECT 81.260 59.600 81.690 59.940 ;
        RECT 81.500 56.930 81.690 59.600 ;
        RECT 81.940 56.840 82.220 67.460 ;
        RECT 83.640 62.700 83.900 63.020 ;
        RECT 82.750 61.830 83.010 62.150 ;
        RECT 82.780 58.110 82.970 61.830 ;
        RECT 83.660 58.110 83.880 62.700 ;
        RECT 85.630 59.480 85.970 75.700 ;
        RECT 86.020 68.760 86.180 69.400 ;
        RECT 86.020 68.210 86.290 68.760 ;
        RECT 86.010 68.160 86.290 68.210 ;
        RECT 86.010 68.070 86.180 68.160 ;
        RECT 86.020 66.380 86.180 68.070 ;
        RECT 86.430 67.950 86.620 69.400 ;
        RECT 86.700 69.070 87.090 72.660 ;
        RECT 90.130 72.240 90.500 72.250 ;
        RECT 90.080 71.790 90.580 72.240 ;
        RECT 87.830 68.590 88.140 69.030 ;
        RECT 86.400 67.920 86.620 67.950 ;
        RECT 86.390 67.650 86.640 67.920 ;
        RECT 86.390 67.640 86.630 67.650 ;
        RECT 86.400 67.400 86.630 67.640 ;
        RECT 86.430 66.380 86.590 67.400 ;
        RECT 86.780 66.630 87.020 66.970 ;
        RECT 86.780 66.590 87.340 66.630 ;
        RECT 86.020 63.860 86.180 65.550 ;
        RECT 86.430 64.530 86.590 65.550 ;
        RECT 86.950 65.340 87.340 66.590 ;
        RECT 86.780 64.960 87.340 65.340 ;
        RECT 86.400 64.290 86.630 64.530 ;
        RECT 86.390 64.280 86.630 64.290 ;
        RECT 86.390 64.010 86.640 64.280 ;
        RECT 86.400 63.980 86.620 64.010 ;
        RECT 86.010 63.770 86.180 63.860 ;
        RECT 86.010 63.750 86.290 63.770 ;
        RECT 86.430 63.750 86.620 63.980 ;
        RECT 86.010 63.720 86.620 63.750 ;
        RECT 86.020 63.380 86.620 63.720 ;
        RECT 86.020 63.370 86.290 63.380 ;
        RECT 86.300 63.370 86.620 63.380 ;
        RECT 86.020 63.170 86.620 63.370 ;
        RECT 86.020 62.530 86.180 63.170 ;
        RECT 86.270 62.530 86.620 63.170 ;
        RECT 86.270 62.180 86.570 62.530 ;
        RECT 86.260 62.040 86.570 62.180 ;
        RECT 86.270 60.350 86.570 62.040 ;
        RECT 86.680 61.920 86.870 63.370 ;
        RECT 86.950 63.040 87.340 64.960 ;
        RECT 87.830 63.000 88.140 63.340 ;
        RECT 87.830 62.900 88.390 63.000 ;
        RECT 88.080 62.610 88.390 62.900 ;
        RECT 86.650 61.890 86.870 61.920 ;
        RECT 87.840 62.560 88.390 62.610 ;
        RECT 86.640 61.620 86.890 61.890 ;
        RECT 87.840 61.820 88.100 62.560 ;
        RECT 86.640 61.610 86.880 61.620 ;
        RECT 86.650 61.370 86.880 61.610 ;
        RECT 86.680 60.350 86.840 61.370 ;
        RECT 87.030 60.560 87.270 60.940 ;
        RECT 86.300 59.520 86.570 60.350 ;
        RECT 85.580 59.400 85.970 59.480 ;
        RECT 85.570 58.630 85.970 59.400 ;
        RECT 85.580 58.560 85.970 58.630 ;
        RECT 82.610 57.420 83.290 58.110 ;
        RECT 83.650 57.420 84.330 58.110 ;
        RECT 85.630 56.780 85.970 58.560 ;
        RECT 86.270 58.000 86.570 59.520 ;
        RECT 86.680 58.500 86.840 59.520 ;
        RECT 87.030 58.930 87.270 59.310 ;
        RECT 86.650 58.260 86.880 58.500 ;
        RECT 86.640 58.250 86.880 58.260 ;
        RECT 86.640 58.000 86.890 58.250 ;
        RECT 86.270 57.830 86.980 58.000 ;
        RECT 86.260 57.690 86.980 57.830 ;
        RECT 86.270 57.500 86.980 57.690 ;
        RECT 86.270 56.850 86.570 57.500 ;
        RECT 86.270 56.500 86.430 56.850 ;
        RECT 86.680 56.500 86.870 57.500 ;
        RECT 87.840 57.310 88.100 57.950 ;
        RECT 87.840 57.160 88.390 57.310 ;
        RECT 88.080 56.870 88.390 57.160 ;
        RECT 68.440 49.550 68.670 49.580 ;
        RECT 68.450 49.140 68.670 49.550 ;
        RECT 68.450 49.130 68.730 49.140 ;
        RECT 66.160 47.940 66.410 48.160 ;
        RECT 51.720 45.840 52.040 45.930 ;
        RECT 51.720 45.400 52.010 45.840 ;
        RECT 52.240 43.440 52.530 47.910 ;
        RECT 53.700 43.950 53.890 47.850 ;
        RECT 55.010 44.050 55.240 47.890 ;
        RECT 57.980 44.060 58.230 47.910 ;
        RECT 68.450 47.720 68.670 49.130 ;
        RECT 71.930 48.460 72.320 50.320 ;
        RECT 75.960 48.530 76.350 50.390 ;
        RECT 64.200 47.650 64.390 47.700 ;
        RECT 65.510 47.650 65.740 47.720 ;
        RECT 68.450 47.650 68.730 47.720 ;
        RECT 68.450 46.350 68.670 47.650 ;
        RECT 68.450 46.260 68.800 46.350 ;
        RECT 68.450 46.040 68.960 46.260 ;
        RECT 76.840 45.510 77.220 52.010 ;
        RECT 78.590 47.760 78.750 48.460 ;
        RECT 78.590 47.210 78.860 47.760 ;
        RECT 78.580 47.160 78.860 47.210 ;
        RECT 79.000 47.420 79.190 48.410 ;
        RECT 79.400 47.730 79.560 48.460 ;
        RECT 80.240 47.870 80.560 48.190 ;
        RECT 90.130 48.060 90.500 71.790 ;
        RECT 90.780 68.940 90.940 68.990 ;
        RECT 91.190 68.930 91.380 68.990 ;
        RECT 90.920 68.340 91.380 68.770 ;
        RECT 93.060 68.700 93.270 68.990 ;
        RECT 92.950 68.410 93.270 68.700 ;
        RECT 90.940 62.990 91.310 68.340 ;
        RECT 92.050 66.790 92.370 67.110 ;
        RECT 93.060 66.710 93.270 68.410 ;
        RECT 93.530 68.140 93.720 68.990 ;
        RECT 93.420 67.850 93.720 68.140 ;
        RECT 92.950 66.420 93.270 66.710 ;
        RECT 91.420 66.170 91.680 66.230 ;
        RECT 93.060 66.200 93.270 66.420 ;
        RECT 91.420 65.910 91.780 66.170 ;
        RECT 91.540 65.750 91.780 65.910 ;
        RECT 93.530 65.820 93.720 67.850 ;
        RECT 93.940 66.530 94.150 68.990 ;
        RECT 93.820 66.020 94.150 66.530 ;
        RECT 93.080 65.640 93.270 65.690 ;
        RECT 92.040 65.100 92.360 65.420 ;
        RECT 92.960 65.350 93.270 65.640 ;
        RECT 93.420 65.530 93.720 65.820 ;
        RECT 91.690 63.630 92.140 64.060 ;
        RECT 93.080 63.730 93.270 65.350 ;
        RECT 93.530 64.240 93.720 65.530 ;
        RECT 93.410 63.950 93.720 64.240 ;
        RECT 90.780 62.940 91.380 62.990 ;
        RECT 90.910 56.910 91.310 62.940 ;
        RECT 91.440 62.900 91.630 62.960 ;
        RECT 91.710 60.490 92.080 63.630 ;
        RECT 92.760 63.440 92.770 63.450 ;
        RECT 92.980 63.440 93.270 63.730 ;
        RECT 93.070 62.940 93.300 63.440 ;
        RECT 93.530 62.940 93.720 63.950 ;
        RECT 93.940 62.940 94.150 66.020 ;
        RECT 95.020 64.460 95.200 68.990 ;
        RECT 98.890 66.130 99.120 68.990 ;
        RECT 98.790 65.840 99.120 66.130 ;
        RECT 94.960 64.120 95.250 64.460 ;
        RECT 95.020 62.940 95.200 64.120 ;
        RECT 92.540 61.330 92.860 61.650 ;
        RECT 95.050 61.010 95.610 61.660 ;
        RECT 96.000 61.500 96.560 62.080 ;
        RECT 97.080 61.960 97.640 62.550 ;
        RECT 91.680 60.170 92.080 60.490 ;
        RECT 91.710 59.890 92.080 60.170 ;
        RECT 91.680 59.570 92.080 59.890 ;
        RECT 91.440 56.910 91.630 56.970 ;
        RECT 81.480 47.780 81.640 47.830 ;
        RECT 81.890 47.780 82.080 47.830 ;
        RECT 82.290 47.790 82.450 47.830 ;
        RECT 79.360 47.710 79.560 47.730 ;
        RECT 79.350 47.470 79.580 47.710 ;
        RECT 79.350 47.420 79.560 47.470 ;
        RECT 79.000 47.300 79.170 47.420 ;
        RECT 78.580 47.070 78.750 47.160 ;
        RECT 78.590 46.560 78.750 47.070 ;
        RECT 79.000 46.560 79.160 47.300 ;
        RECT 79.400 46.560 79.560 47.420 ;
        RECT 80.240 47.320 80.560 47.640 ;
        RECT 84.230 46.670 84.470 48.060 ;
        RECT 86.410 47.730 86.790 48.060 ;
        RECT 78.590 45.780 78.750 46.290 ;
        RECT 78.580 45.690 78.750 45.780 ;
        RECT 78.580 45.640 78.860 45.690 ;
        RECT 53.680 43.450 53.890 43.950 ;
        RECT 54.990 43.640 55.240 44.050 ;
        RECT 57.960 43.640 58.230 44.060 ;
        RECT 59.740 44.210 60.020 45.320 ;
        RECT 60.270 44.630 60.460 45.230 ;
        RECT 62.270 44.790 62.660 44.810 ;
        RECT 62.260 44.700 62.660 44.790 ;
        RECT 62.110 44.690 62.660 44.700 ;
        RECT 60.270 44.440 61.870 44.630 ;
        RECT 59.740 43.930 61.460 44.210 ;
        RECT 61.260 43.700 61.460 43.930 ;
        RECT 53.680 43.320 53.870 43.450 ;
        RECT 54.990 43.210 55.220 43.640 ;
        RECT 57.960 43.270 58.210 43.640 ;
        RECT 61.270 43.400 61.430 43.700 ;
        RECT 61.680 43.320 61.870 44.440 ;
        RECT 62.080 44.450 62.660 44.690 ;
        RECT 62.080 44.430 62.650 44.450 ;
        RECT 62.080 44.420 62.270 44.430 ;
        RECT 62.080 43.580 62.250 44.420 ;
        RECT 66.750 44.360 66.980 45.270 ;
        RECT 67.970 44.390 68.200 45.270 ;
        RECT 66.230 44.290 66.980 44.360 ;
        RECT 66.200 44.130 66.980 44.290 ;
        RECT 67.950 44.330 68.200 44.390 ;
        RECT 71.280 44.460 71.700 45.460 ;
        RECT 66.200 43.680 66.610 44.130 ;
        RECT 62.080 43.310 62.240 43.580 ;
        RECT 64.180 43.160 64.370 43.230 ;
        RECT 65.490 43.150 65.720 43.230 ;
        RECT 66.200 43.190 66.580 43.680 ;
        RECT 67.950 43.330 68.190 44.330 ;
        RECT 71.280 44.280 71.710 44.460 ;
        RECT 71.280 43.890 71.720 44.280 ;
        RECT 73.760 44.070 73.990 45.270 ;
        RECT 71.310 43.680 71.720 43.890 ;
        RECT 71.310 43.170 71.710 43.680 ;
        RECT 73.750 43.330 73.990 44.070 ;
        RECT 74.980 44.380 75.210 45.270 ;
        RECT 78.590 45.090 78.860 45.640 ;
        RECT 79.000 45.550 79.160 46.290 ;
        RECT 79.000 45.430 79.170 45.550 ;
        RECT 79.400 45.430 79.560 46.290 ;
        RECT 84.220 46.010 84.490 46.670 ;
        RECT 88.160 46.650 88.400 48.060 ;
        RECT 78.590 44.520 78.750 45.090 ;
        RECT 74.980 44.000 75.740 44.380 ;
        RECT 75.360 43.540 75.740 44.000 ;
        RECT 78.590 43.970 78.860 44.520 ;
        RECT 78.580 43.920 78.860 43.970 ;
        RECT 79.000 44.180 79.190 45.430 ;
        RECT 79.350 45.380 79.560 45.430 ;
        RECT 79.350 45.140 79.580 45.380 ;
        RECT 80.240 45.210 80.560 45.530 ;
        RECT 79.360 45.120 79.560 45.140 ;
        RECT 79.400 44.490 79.560 45.120 ;
        RECT 80.240 44.630 80.560 44.980 ;
        RECT 79.360 44.470 79.560 44.490 ;
        RECT 79.350 44.230 79.580 44.470 ;
        RECT 80.240 44.250 80.560 44.400 ;
        RECT 81.500 44.250 81.690 45.230 ;
        RECT 81.940 44.940 82.220 45.320 ;
        RECT 81.890 44.920 82.220 44.940 ;
        RECT 81.860 44.900 82.220 44.920 ;
        RECT 81.860 44.710 82.300 44.900 ;
        RECT 81.860 44.690 82.220 44.710 ;
        RECT 81.890 44.650 82.220 44.690 ;
        RECT 79.350 44.180 79.560 44.230 ;
        RECT 79.000 44.060 79.170 44.180 ;
        RECT 78.580 43.830 78.750 43.920 ;
        RECT 78.590 43.320 78.750 43.830 ;
        RECT 79.000 43.320 79.160 44.060 ;
        RECT 79.400 43.320 79.560 44.180 ;
        RECT 79.670 43.880 79.950 44.200 ;
        RECT 80.100 44.060 81.690 44.250 ;
        RECT 79.700 43.400 79.860 43.880 ;
        RECT 80.100 43.730 80.290 44.060 ;
        RECT 81.940 43.870 82.220 44.650 ;
        RECT 80.550 43.860 82.220 43.870 ;
        RECT 80.070 43.620 80.290 43.730 ;
        RECT 80.070 43.320 80.260 43.620 ;
        RECT 80.510 43.590 82.220 43.860 ;
        RECT 80.510 43.400 80.670 43.590 ;
        RECT 84.230 43.480 84.470 46.010 ;
        RECT 88.150 45.990 88.410 46.650 ;
        RECT 83.960 43.420 84.470 43.480 ;
        RECT 83.960 43.340 84.480 43.420 ;
        RECT 88.160 43.380 88.400 45.990 ;
        RECT 90.130 44.880 90.840 48.060 ;
        RECT 90.100 44.420 90.840 44.880 ;
        RECT 90.130 44.380 90.840 44.420 ;
        RECT 90.440 43.380 90.840 44.380 ;
        RECT 90.940 44.290 91.310 56.910 ;
        RECT 90.910 43.830 91.350 44.290 ;
        RECT 90.940 43.780 91.310 43.830 ;
        RECT 83.950 43.190 84.480 43.340 ;
        RECT 84.520 43.330 84.710 43.380 ;
        RECT 84.920 43.330 85.080 43.380 ;
        RECT 86.860 43.290 87.100 43.380 ;
        RECT 61.860 42.840 62.050 43.060 ;
        RECT 44.480 42.660 44.720 42.710 ;
        RECT 47.420 42.650 47.730 42.710 ;
        RECT 51.750 42.590 52.040 42.710 ;
        RECT 61.580 42.350 62.050 42.840 ;
        RECT 62.440 42.700 62.810 42.720 ;
        RECT 62.390 42.440 62.810 42.700 ;
        RECT 62.440 42.430 62.810 42.440 ;
        RECT 46.490 41.270 46.900 41.600 ;
        RECT 44.450 40.520 44.690 40.590 ;
        RECT 47.230 40.580 47.470 41.780 ;
        RECT 49.630 41.220 49.920 41.230 ;
        RECT 49.610 40.950 49.930 41.220 ;
        RECT 49.610 40.940 49.920 40.950 ;
        RECT 48.650 40.740 48.850 40.760 ;
        RECT 47.230 40.520 47.700 40.580 ;
        RECT 47.230 40.100 47.470 40.520 ;
        RECT 48.650 40.450 49.000 40.740 ;
        RECT 50.170 40.090 50.480 41.780 ;
        RECT 50.730 41.180 51.010 41.490 ;
        RECT 50.650 41.160 51.010 41.180 ;
        RECT 50.650 40.880 50.970 41.160 ;
        RECT 46.490 39.520 46.900 39.850 ;
        RECT 44.450 38.770 44.690 38.840 ;
        RECT 47.230 38.830 47.470 40.030 ;
        RECT 49.630 39.470 49.920 39.480 ;
        RECT 49.610 39.200 49.930 39.470 ;
        RECT 49.610 39.190 49.920 39.200 ;
        RECT 48.650 38.990 48.850 39.010 ;
        RECT 47.230 38.770 47.700 38.830 ;
        RECT 47.230 38.350 47.470 38.770 ;
        RECT 48.650 38.700 49.000 38.990 ;
        RECT 50.170 38.340 50.480 40.030 ;
        RECT 50.730 39.430 51.010 39.740 ;
        RECT 50.650 39.410 51.010 39.430 ;
        RECT 50.650 39.130 50.970 39.410 ;
        RECT 46.490 37.770 46.900 38.100 ;
        RECT 44.450 37.020 44.690 37.090 ;
        RECT 44.870 36.870 45.110 37.730 ;
        RECT 47.230 37.080 47.470 38.280 ;
        RECT 47.230 37.020 47.700 37.080 ;
        RECT 44.480 35.710 44.720 35.760 ;
        RECT 44.450 35.270 44.690 35.340 ;
        RECT 44.870 33.960 45.210 36.870 ;
        RECT 47.230 36.600 47.470 37.020 ;
        RECT 47.810 36.870 48.120 37.800 ;
        RECT 49.630 37.720 49.920 37.730 ;
        RECT 49.610 37.450 49.930 37.720 ;
        RECT 49.610 37.440 49.920 37.450 ;
        RECT 48.650 37.240 48.850 37.260 ;
        RECT 48.650 36.950 49.000 37.240 ;
        RECT 46.490 36.020 46.900 36.350 ;
        RECT 47.230 35.770 47.470 36.530 ;
        RECT 47.230 35.710 47.730 35.770 ;
        RECT 47.230 35.330 47.470 35.710 ;
        RECT 47.230 35.270 47.700 35.330 ;
        RECT 47.230 34.850 47.470 35.270 ;
        RECT 47.810 33.960 48.220 36.870 ;
        RECT 50.170 36.590 50.480 38.280 ;
        RECT 50.730 37.680 51.010 37.990 ;
        RECT 50.650 37.660 51.010 37.680 ;
        RECT 50.650 37.380 50.970 37.660 ;
        RECT 49.630 35.970 49.920 35.980 ;
        RECT 49.610 35.700 49.930 35.970 ;
        RECT 49.610 35.690 49.920 35.700 ;
        RECT 48.650 35.490 48.850 35.510 ;
        RECT 48.650 35.200 49.000 35.490 ;
        RECT 50.170 34.840 50.480 36.530 ;
        RECT 50.730 35.930 51.010 36.240 ;
        RECT 50.650 35.910 51.010 35.930 ;
        RECT 50.650 35.630 50.970 35.910 ;
        RECT 51.720 35.800 52.010 42.270 ;
        RECT 61.400 41.910 61.720 42.190 ;
        RECT 61.860 42.010 62.050 42.350 ;
        RECT 61.400 41.540 61.720 41.820 ;
        RECT 61.760 41.720 62.050 42.010 ;
        RECT 61.860 41.380 62.050 41.720 ;
        RECT 61.580 40.890 62.050 41.380 ;
        RECT 62.440 41.290 62.810 41.300 ;
        RECT 62.390 41.030 62.810 41.290 ;
        RECT 62.440 41.010 62.810 41.030 ;
        RECT 61.860 40.670 62.050 40.890 ;
        RECT 63.170 40.670 63.400 43.060 ;
        RECT 66.140 42.840 66.390 43.060 ;
        RECT 64.900 42.680 65.240 42.730 ;
        RECT 64.900 42.660 65.460 42.680 ;
        RECT 64.780 42.490 65.460 42.660 ;
        RECT 64.900 42.450 65.460 42.490 ;
        RECT 64.900 42.410 65.240 42.450 ;
        RECT 64.900 41.280 65.240 41.320 ;
        RECT 64.900 41.240 65.460 41.280 ;
        RECT 64.780 41.070 65.460 41.240 ;
        RECT 64.900 41.050 65.460 41.070 ;
        RECT 64.900 41.000 65.240 41.050 ;
        RECT 66.140 40.890 66.780 42.840 ;
        RECT 68.460 41.860 68.710 41.870 ;
        RECT 66.140 40.670 66.390 40.890 ;
        RECT 61.860 39.640 62.050 39.860 ;
        RECT 61.580 39.150 62.050 39.640 ;
        RECT 62.440 39.500 62.810 39.520 ;
        RECT 62.390 39.240 62.810 39.500 ;
        RECT 62.440 39.230 62.810 39.240 ;
        RECT 61.400 38.710 61.720 38.990 ;
        RECT 61.860 38.810 62.050 39.150 ;
        RECT 61.400 38.340 61.720 38.620 ;
        RECT 61.760 38.520 62.050 38.810 ;
        RECT 61.860 38.180 62.050 38.520 ;
        RECT 51.720 35.710 52.040 35.800 ;
        RECT 51.720 35.270 52.010 35.710 ;
        RECT 52.240 33.960 52.530 37.780 ;
        RECT 44.970 33.720 45.210 33.960 ;
        RECT 47.910 33.690 48.220 33.960 ;
        RECT 53.700 33.690 53.890 37.780 ;
        RECT 55.010 36.740 55.240 37.820 ;
        RECT 54.920 36.260 55.250 36.740 ;
        RECT 55.010 33.650 55.240 36.260 ;
        RECT 57.980 33.860 58.230 37.840 ;
        RECT 61.300 33.800 61.460 37.850 ;
        RECT 61.580 37.690 62.050 38.180 ;
        RECT 62.440 38.090 62.810 38.100 ;
        RECT 62.390 37.830 62.810 38.090 ;
        RECT 62.440 37.810 62.810 37.830 ;
        RECT 61.860 37.470 62.050 37.690 ;
        RECT 63.170 37.470 63.400 39.860 ;
        RECT 66.140 39.640 66.390 39.860 ;
        RECT 64.900 39.480 65.240 39.530 ;
        RECT 64.900 39.460 65.460 39.480 ;
        RECT 64.780 39.290 65.460 39.460 ;
        RECT 64.900 39.250 65.460 39.290 ;
        RECT 64.900 39.210 65.240 39.250 ;
        RECT 64.900 38.080 65.240 38.120 ;
        RECT 64.900 38.040 65.460 38.080 ;
        RECT 64.050 37.230 64.290 37.930 ;
        RECT 64.780 37.870 65.460 38.040 ;
        RECT 64.900 37.850 65.460 37.870 ;
        RECT 64.900 37.800 65.240 37.850 ;
        RECT 66.140 37.690 66.780 39.640 ;
        RECT 72.530 39.580 72.920 41.440 ;
        RECT 76.560 39.650 76.950 41.510 ;
        RECT 68.460 38.660 68.710 38.670 ;
        RECT 66.140 37.470 66.610 37.690 ;
        RECT 64.050 37.180 64.370 37.230 ;
        RECT 65.490 37.180 65.720 37.250 ;
        RECT 64.050 34.210 64.290 37.180 ;
        RECT 64.030 33.960 64.420 34.210 ;
        RECT 44.440 33.600 44.680 33.650 ;
        RECT 47.380 33.590 47.690 33.650 ;
        RECT 51.710 33.530 52.000 33.650 ;
        RECT 61.890 33.570 62.080 33.790 ;
        RECT 46.450 32.210 46.860 32.540 ;
        RECT 44.410 31.460 44.650 31.530 ;
        RECT 47.190 31.520 47.430 32.720 ;
        RECT 49.590 32.160 49.880 32.170 ;
        RECT 49.570 31.890 49.890 32.160 ;
        RECT 49.570 31.880 49.880 31.890 ;
        RECT 48.610 31.680 48.810 31.700 ;
        RECT 47.190 31.460 47.660 31.520 ;
        RECT 47.190 31.040 47.430 31.460 ;
        RECT 48.610 31.390 48.960 31.680 ;
        RECT 50.130 31.030 50.440 32.720 ;
        RECT 50.690 32.120 50.970 32.430 ;
        RECT 50.610 32.100 50.970 32.120 ;
        RECT 50.610 31.820 50.930 32.100 ;
        RECT 46.450 30.460 46.860 30.790 ;
        RECT 44.410 29.710 44.650 29.780 ;
        RECT 47.190 29.770 47.430 30.970 ;
        RECT 49.590 30.410 49.880 30.420 ;
        RECT 49.570 30.140 49.890 30.410 ;
        RECT 49.570 30.130 49.880 30.140 ;
        RECT 48.610 29.930 48.810 29.950 ;
        RECT 47.190 29.710 47.660 29.770 ;
        RECT 47.190 29.290 47.430 29.710 ;
        RECT 48.610 29.640 48.960 29.930 ;
        RECT 50.130 29.280 50.440 30.970 ;
        RECT 50.690 30.370 50.970 30.680 ;
        RECT 50.610 30.350 50.970 30.370 ;
        RECT 50.610 30.070 50.930 30.350 ;
        RECT 46.450 28.710 46.860 29.040 ;
        RECT 44.410 27.960 44.650 28.030 ;
        RECT 47.190 28.020 47.430 29.220 ;
        RECT 49.590 28.660 49.880 28.670 ;
        RECT 49.570 28.390 49.890 28.660 ;
        RECT 49.570 28.380 49.880 28.390 ;
        RECT 48.610 28.180 48.810 28.200 ;
        RECT 47.190 27.960 47.660 28.020 ;
        RECT 44.440 26.650 44.680 26.700 ;
        RECT 44.410 26.210 44.650 26.280 ;
        RECT 44.870 15.330 45.110 27.960 ;
        RECT 47.190 27.540 47.430 27.960 ;
        RECT 46.450 26.960 46.860 27.290 ;
        RECT 47.190 26.710 47.430 27.470 ;
        RECT 47.810 26.880 48.120 28.030 ;
        RECT 48.610 27.890 48.960 28.180 ;
        RECT 50.130 27.530 50.440 29.220 ;
        RECT 50.690 28.620 50.970 28.930 ;
        RECT 50.610 28.600 50.970 28.620 ;
        RECT 50.610 28.320 50.930 28.600 ;
        RECT 49.590 26.910 49.880 26.920 ;
        RECT 47.190 26.650 47.690 26.710 ;
        RECT 47.190 26.270 47.430 26.650 ;
        RECT 47.770 26.550 48.140 26.880 ;
        RECT 49.570 26.640 49.890 26.910 ;
        RECT 49.570 26.630 49.880 26.640 ;
        RECT 47.190 26.210 47.660 26.270 ;
        RECT 47.190 25.790 47.430 26.210 ;
        RECT 47.810 25.340 48.120 26.550 ;
        RECT 48.610 26.430 48.810 26.450 ;
        RECT 48.610 26.140 48.960 26.430 ;
        RECT 50.130 25.780 50.440 27.470 ;
        RECT 50.690 26.870 50.970 27.180 ;
        RECT 50.610 26.850 50.970 26.870 ;
        RECT 50.610 26.570 50.930 26.850 ;
        RECT 51.680 26.740 51.970 33.210 ;
        RECT 61.610 33.080 62.080 33.570 ;
        RECT 62.470 33.430 62.840 33.450 ;
        RECT 62.420 33.170 62.840 33.430 ;
        RECT 62.470 33.160 62.840 33.170 ;
        RECT 59.330 32.530 59.650 32.870 ;
        RECT 61.430 32.640 61.750 32.920 ;
        RECT 61.890 32.740 62.080 33.080 ;
        RECT 52.240 27.390 52.530 28.010 ;
        RECT 52.740 27.410 53.080 27.730 ;
        RECT 52.210 27.040 52.560 27.390 ;
        RECT 51.680 26.650 52.000 26.740 ;
        RECT 51.680 26.580 51.970 26.650 ;
        RECT 52.240 26.580 52.530 27.040 ;
        RECT 52.740 26.800 52.990 27.410 ;
        RECT 53.700 26.820 53.890 28.020 ;
        RECT 57.980 27.350 58.230 28.080 ;
        RECT 59.410 27.770 59.620 32.530 ;
        RECT 61.430 32.270 61.750 32.550 ;
        RECT 61.790 32.450 62.080 32.740 ;
        RECT 61.890 32.110 62.080 32.450 ;
        RECT 61.610 31.620 62.080 32.110 ;
        RECT 62.470 32.020 62.840 32.030 ;
        RECT 62.420 31.760 62.840 32.020 ;
        RECT 62.470 31.740 62.840 31.760 ;
        RECT 61.890 31.400 62.080 31.620 ;
        RECT 63.200 31.400 63.430 33.790 ;
        RECT 64.170 33.710 64.420 33.960 ;
        RECT 65.520 33.880 65.750 33.960 ;
        RECT 66.230 33.790 66.610 37.470 ;
        RECT 67.980 34.190 68.220 37.930 ;
        RECT 68.460 37.180 68.710 37.250 ;
        RECT 67.980 33.920 68.450 34.190 ;
        RECT 66.170 33.580 66.610 33.790 ;
        RECT 68.180 33.690 68.450 33.920 ;
        RECT 66.170 33.570 66.420 33.580 ;
        RECT 64.930 33.410 65.270 33.460 ;
        RECT 64.930 33.390 65.490 33.410 ;
        RECT 64.810 33.220 65.490 33.390 ;
        RECT 64.930 33.180 65.490 33.220 ;
        RECT 64.930 33.140 65.270 33.180 ;
        RECT 64.930 32.010 65.270 32.050 ;
        RECT 64.930 31.970 65.490 32.010 ;
        RECT 64.810 31.800 65.490 31.970 ;
        RECT 64.930 31.780 65.490 31.800 ;
        RECT 64.930 31.730 65.270 31.780 ;
        RECT 66.170 31.620 66.810 33.570 ;
        RECT 70.260 33.560 70.660 38.090 ;
        RECT 73.780 35.420 74.020 37.930 ;
        RECT 77.440 36.670 77.820 43.170 ;
        RECT 84.110 43.100 84.480 43.190 ;
        RECT 78.590 42.550 78.750 43.060 ;
        RECT 78.580 42.460 78.750 42.550 ;
        RECT 78.580 42.410 78.860 42.460 ;
        RECT 78.590 41.860 78.860 42.410 ;
        RECT 79.000 42.320 79.160 43.060 ;
        RECT 79.000 42.200 79.170 42.320 ;
        RECT 79.400 42.200 79.560 43.060 ;
        RECT 84.110 43.040 84.470 43.100 ;
        RECT 88.150 43.060 88.410 43.380 ;
        RECT 89.040 43.280 89.420 43.380 ;
        RECT 90.440 43.320 91.030 43.380 ;
        RECT 78.590 41.160 78.750 41.860 ;
        RECT 79.000 41.210 79.190 42.200 ;
        RECT 79.350 42.150 79.560 42.200 ;
        RECT 79.350 41.910 79.580 42.150 ;
        RECT 80.240 41.980 80.560 42.300 ;
        RECT 79.360 41.890 79.560 41.910 ;
        RECT 79.400 41.160 79.560 41.890 ;
        RECT 80.240 41.430 80.560 41.750 ;
        RECT 84.230 41.560 84.470 43.040 ;
        RECT 86.410 41.560 86.790 42.160 ;
        RECT 88.160 41.560 88.400 43.060 ;
        RECT 90.440 41.560 90.840 43.320 ;
        RECT 91.710 41.940 92.080 59.570 ;
        RECT 92.580 58.890 93.010 58.990 ;
        RECT 92.540 58.570 93.010 58.890 ;
        RECT 95.070 58.670 95.570 61.010 ;
        RECT 92.580 58.550 93.010 58.570 ;
        RECT 94.870 58.610 95.590 58.670 ;
        RECT 91.680 41.930 92.080 41.940 ;
        RECT 91.670 41.510 92.090 41.930 ;
        RECT 91.710 41.500 92.080 41.510 ;
        RECT 79.190 38.920 79.350 39.620 ;
        RECT 79.190 38.370 79.460 38.920 ;
        RECT 79.180 38.320 79.460 38.370 ;
        RECT 79.600 38.580 79.790 39.570 ;
        RECT 80.000 38.890 80.160 39.620 ;
        RECT 80.840 39.030 81.160 39.350 ;
        RECT 79.960 38.870 80.160 38.890 ;
        RECT 82.080 38.880 82.240 38.950 ;
        RECT 82.490 38.880 82.680 38.950 ;
        RECT 82.890 38.880 83.050 38.950 ;
        RECT 79.950 38.630 80.180 38.870 ;
        RECT 79.950 38.580 80.160 38.630 ;
        RECT 79.600 38.460 79.770 38.580 ;
        RECT 79.180 38.230 79.350 38.320 ;
        RECT 79.190 37.720 79.350 38.230 ;
        RECT 79.600 37.720 79.760 38.460 ;
        RECT 80.000 37.720 80.160 38.580 ;
        RECT 80.840 38.480 81.160 38.800 ;
        RECT 79.190 36.960 79.350 37.470 ;
        RECT 79.180 36.870 79.350 36.960 ;
        RECT 79.180 36.820 79.460 36.870 ;
        RECT 79.190 36.270 79.460 36.820 ;
        RECT 79.600 36.730 79.760 37.470 ;
        RECT 79.600 36.610 79.770 36.730 ;
        RECT 80.000 36.610 80.160 37.470 ;
        RECT 84.950 37.400 85.200 39.220 ;
        RECT 87.010 38.850 87.390 39.220 ;
        RECT 88.960 37.420 89.230 39.220 ;
        RECT 84.110 37.330 84.270 37.390 ;
        RECT 84.520 37.340 84.710 37.400 ;
        RECT 84.920 37.340 85.200 37.400 ;
        RECT 79.190 35.680 79.350 36.270 ;
        RECT 73.780 35.180 74.360 35.420 ;
        RECT 74.120 33.840 74.360 35.180 ;
        RECT 79.190 35.130 79.460 35.680 ;
        RECT 79.180 35.080 79.460 35.130 ;
        RECT 79.600 35.340 79.790 36.610 ;
        RECT 79.950 36.560 80.160 36.610 ;
        RECT 79.950 36.320 80.180 36.560 ;
        RECT 80.840 36.390 81.160 36.710 ;
        RECT 79.960 36.300 80.160 36.320 ;
        RECT 80.000 35.650 80.160 36.300 ;
        RECT 80.840 35.790 81.160 36.160 ;
        RECT 82.460 36.070 82.700 36.100 ;
        RECT 82.460 35.980 82.890 36.070 ;
        RECT 82.080 35.970 82.240 35.980 ;
        RECT 82.460 35.970 83.050 35.980 ;
        RECT 82.460 35.900 82.890 35.970 ;
        RECT 82.460 35.870 82.700 35.900 ;
        RECT 82.490 35.770 82.600 35.870 ;
        RECT 79.960 35.630 80.160 35.650 ;
        RECT 79.950 35.390 80.180 35.630 ;
        RECT 79.950 35.340 80.160 35.390 ;
        RECT 79.600 35.220 79.770 35.340 ;
        RECT 79.180 34.990 79.350 35.080 ;
        RECT 79.190 34.480 79.350 34.990 ;
        RECT 79.600 34.480 79.760 35.220 ;
        RECT 80.000 34.480 80.160 35.340 ;
        RECT 80.840 35.240 81.160 35.560 ;
        RECT 84.950 34.540 85.200 37.340 ;
        RECT 86.860 37.330 87.100 37.410 ;
        RECT 88.960 37.330 89.420 37.420 ;
        RECT 90.790 37.330 91.030 37.400 ;
        RECT 84.720 34.470 84.880 34.540 ;
        RECT 84.950 34.510 85.320 34.540 ;
        RECT 84.930 34.480 85.320 34.510 ;
        RECT 84.920 34.470 85.320 34.480 ;
        RECT 85.530 34.470 85.690 34.540 ;
        RECT 88.960 34.480 89.230 37.330 ;
        RECT 79.190 33.710 79.350 34.220 ;
        RECT 79.180 33.620 79.350 33.710 ;
        RECT 79.180 33.570 79.460 33.620 ;
        RECT 79.190 33.020 79.460 33.570 ;
        RECT 79.600 33.480 79.760 34.220 ;
        RECT 79.600 33.360 79.770 33.480 ;
        RECT 80.000 33.360 80.160 34.220 ;
        RECT 84.920 34.200 85.220 34.470 ;
        RECT 84.930 34.180 85.210 34.200 ;
        RECT 79.190 32.840 79.350 33.020 ;
        RECT 68.490 32.590 68.740 32.600 ;
        RECT 79.190 32.520 79.500 32.840 ;
        RECT 79.190 32.320 79.480 32.520 ;
        RECT 79.600 32.370 79.790 33.360 ;
        RECT 79.950 33.310 80.160 33.360 ;
        RECT 79.950 33.070 80.180 33.310 ;
        RECT 80.840 33.140 81.160 33.460 ;
        RECT 79.960 33.050 80.160 33.070 ;
        RECT 80.000 32.320 80.160 33.050 ;
        RECT 82.080 32.910 82.240 32.980 ;
        RECT 82.490 32.910 82.680 32.980 ;
        RECT 82.890 32.910 83.050 32.980 ;
        RECT 80.840 32.590 81.160 32.910 ;
        RECT 83.950 32.610 84.210 32.830 ;
        RECT 84.950 32.720 85.200 34.180 ;
        RECT 87.240 34.060 87.500 34.380 ;
        RECT 88.940 34.170 89.250 34.480 ;
        RECT 89.650 34.440 90.030 34.540 ;
        RECT 87.150 33.330 87.360 33.960 ;
        RECT 87.150 33.220 87.480 33.330 ;
        RECT 87.220 33.010 87.480 33.220 ;
        RECT 87.010 32.720 87.390 33.000 ;
        RECT 88.960 32.720 89.230 34.170 ;
        RECT 91.040 32.720 91.440 39.220 ;
        RECT 92.590 36.760 92.960 58.550 ;
        RECT 94.870 58.340 95.570 58.610 ;
        RECT 93.070 43.250 93.470 43.380 ;
        RECT 94.150 43.280 94.550 43.380 ;
        RECT 93.470 43.020 94.150 43.240 ;
        RECT 93.070 37.330 93.470 37.450 ;
        RECT 94.150 37.330 94.550 37.450 ;
        RECT 92.550 36.250 93.040 36.760 ;
        RECT 92.590 36.220 92.960 36.250 ;
        RECT 93.680 34.260 94.080 34.540 ;
        RECT 83.850 32.510 84.210 32.610 ;
        RECT 66.170 31.400 66.420 31.620 ;
        RECT 78.720 31.590 78.980 31.910 ;
        RECT 60.670 30.840 61.060 31.090 ;
        RECT 59.950 29.740 60.290 30.080 ;
        RECT 59.990 29.720 60.210 29.740 ;
        RECT 59.380 27.450 59.660 27.770 ;
        RECT 59.990 27.440 60.190 29.720 ;
        RECT 60.450 27.900 60.640 28.260 ;
        RECT 57.950 27.060 58.290 27.350 ;
        RECT 59.950 27.120 60.230 27.440 ;
        RECT 60.410 27.430 60.690 27.900 ;
        RECT 51.670 26.300 52.530 26.580 ;
        RECT 51.590 26.290 52.530 26.300 ;
        RECT 52.690 26.690 52.990 26.800 ;
        RECT 51.590 25.820 52.050 26.290 ;
        RECT 47.760 24.860 48.180 25.340 ;
        RECT 52.690 25.180 52.880 26.690 ;
        RECT 53.640 26.500 53.960 26.820 ;
        RECT 56.320 26.290 57.070 26.480 ;
        RECT 56.570 25.450 57.070 26.290 ;
        RECT 60.880 26.210 61.060 30.840 ;
        RECT 61.890 30.370 62.080 30.590 ;
        RECT 61.610 29.880 62.080 30.370 ;
        RECT 62.470 30.230 62.840 30.250 ;
        RECT 62.420 29.970 62.840 30.230 ;
        RECT 62.470 29.960 62.840 29.970 ;
        RECT 61.430 29.440 61.750 29.720 ;
        RECT 61.890 29.540 62.080 29.880 ;
        RECT 61.430 29.070 61.750 29.350 ;
        RECT 61.790 29.250 62.080 29.540 ;
        RECT 61.890 28.910 62.080 29.250 ;
        RECT 61.610 28.420 62.080 28.910 ;
        RECT 62.470 28.820 62.840 28.830 ;
        RECT 62.420 28.560 62.840 28.820 ;
        RECT 62.470 28.540 62.840 28.560 ;
        RECT 61.890 28.200 62.080 28.420 ;
        RECT 63.200 28.200 63.430 30.590 ;
        RECT 66.170 30.370 66.420 30.590 ;
        RECT 64.930 30.210 65.270 30.260 ;
        RECT 64.930 30.190 65.490 30.210 ;
        RECT 64.810 30.020 65.490 30.190 ;
        RECT 64.930 29.980 65.490 30.020 ;
        RECT 64.930 29.940 65.270 29.980 ;
        RECT 64.930 28.810 65.270 28.850 ;
        RECT 64.930 28.770 65.490 28.810 ;
        RECT 64.810 28.600 65.490 28.770 ;
        RECT 64.930 28.580 65.490 28.600 ;
        RECT 64.930 28.530 65.270 28.580 ;
        RECT 66.170 28.420 66.810 30.370 ;
        RECT 78.250 29.750 78.510 30.070 ;
        RECT 68.490 29.390 68.740 29.400 ;
        RECT 77.750 28.820 78.010 29.140 ;
        RECT 66.170 28.200 66.420 28.420 ;
        RECT 62.200 27.370 62.460 27.400 ;
        RECT 62.180 27.070 62.480 27.370 ;
        RECT 62.200 27.060 62.460 27.070 ;
        RECT 60.880 25.910 61.360 26.210 ;
        RECT 62.210 26.140 62.430 27.060 ;
        RECT 64.170 26.930 64.420 28.160 ;
        RECT 65.520 27.910 65.750 27.980 ;
        RECT 68.180 26.950 68.450 28.180 ;
        RECT 68.490 27.910 68.740 27.980 ;
        RECT 71.000 27.380 71.430 27.780 ;
        RECT 64.160 26.670 64.480 26.930 ;
        RECT 68.180 26.640 68.530 26.950 ;
        RECT 60.960 25.800 61.360 25.910 ;
        RECT 62.150 25.740 62.490 26.140 ;
        RECT 62.210 25.660 62.430 25.740 ;
        RECT 66.160 25.470 67.100 26.400 ;
        RECT 71.040 25.590 71.390 27.380 ;
        RECT 72.860 26.820 73.080 28.140 ;
        RECT 74.120 27.420 74.350 28.140 ;
        RECT 74.120 27.190 77.330 27.420 ;
        RECT 74.120 27.180 74.350 27.190 ;
        RECT 72.570 26.580 73.080 26.820 ;
        RECT 52.250 24.860 52.880 25.180 ;
        RECT 56.080 25.130 56.320 25.450 ;
        RECT 57.320 25.130 57.560 25.450 ;
        RECT 65.890 25.150 66.130 25.470 ;
        RECT 67.130 25.150 67.370 25.470 ;
        RECT 72.570 25.330 72.800 26.580 ;
        RECT 77.100 26.220 77.330 27.190 ;
        RECT 77.050 25.820 77.360 26.220 ;
        RECT 72.460 24.890 72.920 25.330 ;
        RECT 52.250 24.760 52.690 24.860 ;
        RECT 56.080 23.790 56.320 24.110 ;
        RECT 57.320 23.780 57.560 24.100 ;
        RECT 65.890 23.810 66.130 24.130 ;
        RECT 67.130 23.800 67.370 24.120 ;
        RECT 77.100 22.650 77.330 25.820 ;
        RECT 76.970 22.430 77.330 22.650 ;
        RECT 55.680 22.160 55.940 22.360 ;
        RECT 57.700 22.160 57.960 22.360 ;
        RECT 52.550 21.790 52.870 22.110 ;
        RECT 53.640 21.790 53.960 22.110 ;
        RECT 54.740 21.780 55.060 22.100 ;
        RECT 52.460 19.580 52.780 21.330 ;
        RECT 53.100 21.110 53.420 21.430 ;
        RECT 54.190 21.090 54.510 21.410 ;
        RECT 55.300 21.080 55.620 21.400 ;
        RECT 55.680 21.350 55.990 22.160 ;
        RECT 57.650 21.350 57.960 22.160 ;
        RECT 65.490 22.190 65.750 22.390 ;
        RECT 67.510 22.190 67.770 22.390 ;
        RECT 76.770 22.200 77.330 22.430 ;
        RECT 76.770 22.190 77.310 22.200 ;
        RECT 58.580 21.780 58.900 22.100 ;
        RECT 59.680 21.790 60.000 22.110 ;
        RECT 60.770 21.790 61.090 22.110 ;
        RECT 62.360 21.820 62.680 22.140 ;
        RECT 63.450 21.820 63.770 22.140 ;
        RECT 64.550 21.810 64.870 22.130 ;
        RECT 53.100 19.740 53.420 20.060 ;
        RECT 54.190 19.740 54.510 20.060 ;
        RECT 55.290 19.740 55.610 20.060 ;
        RECT 52.340 18.980 52.880 19.580 ;
        RECT 53.640 19.010 53.960 19.330 ;
        RECT 54.740 19.010 55.060 19.330 ;
        RECT 52.540 17.640 52.860 17.960 ;
        RECT 53.640 17.640 53.960 17.960 ;
        RECT 54.740 17.640 55.060 17.960 ;
        RECT 51.970 17.000 52.290 17.320 ;
        RECT 53.100 16.960 53.420 17.280 ;
        RECT 54.190 16.960 54.510 17.280 ;
        RECT 55.290 16.970 55.610 17.290 ;
        RECT 51.980 16.530 52.300 16.850 ;
        RECT 55.680 16.370 55.940 21.350 ;
        RECT 56.080 21.020 56.320 21.340 ;
        RECT 57.320 21.010 57.560 21.330 ;
        RECT 57.700 16.370 57.960 21.350 ;
        RECT 58.020 21.080 58.340 21.400 ;
        RECT 59.130 21.090 59.450 21.410 ;
        RECT 60.220 21.110 60.540 21.430 ;
        RECT 58.030 19.740 58.350 20.060 ;
        RECT 59.130 19.740 59.450 20.060 ;
        RECT 60.220 19.740 60.540 20.060 ;
        RECT 60.830 19.330 61.170 21.350 ;
        RECT 58.580 19.010 58.900 19.330 ;
        RECT 59.680 19.010 60.000 19.330 ;
        RECT 60.780 19.010 61.170 19.330 ;
        RECT 60.830 18.560 61.170 19.010 ;
        RECT 62.260 19.360 62.600 21.340 ;
        RECT 62.910 21.140 63.230 21.460 ;
        RECT 64.000 21.120 64.320 21.440 ;
        RECT 65.110 21.110 65.430 21.430 ;
        RECT 65.490 21.380 65.800 22.190 ;
        RECT 67.460 21.380 67.770 22.190 ;
        RECT 68.390 21.810 68.710 22.130 ;
        RECT 69.490 21.820 69.810 22.140 ;
        RECT 70.580 21.820 70.900 22.140 ;
        RECT 74.130 21.790 74.450 22.110 ;
        RECT 75.230 21.800 75.550 22.120 ;
        RECT 76.320 21.800 76.640 22.120 ;
        RECT 62.910 19.770 63.230 20.090 ;
        RECT 64.000 19.770 64.320 20.090 ;
        RECT 65.100 19.770 65.420 20.090 ;
        RECT 62.260 19.040 62.670 19.360 ;
        RECT 63.450 19.040 63.770 19.360 ;
        RECT 64.550 19.040 64.870 19.360 ;
        RECT 60.770 18.040 61.230 18.560 ;
        RECT 62.260 17.990 62.600 19.040 ;
        RECT 58.580 17.640 58.900 17.960 ;
        RECT 59.680 17.640 60.000 17.960 ;
        RECT 60.780 17.640 61.100 17.960 ;
        RECT 62.260 17.670 62.670 17.990 ;
        RECT 63.450 17.670 63.770 17.990 ;
        RECT 64.550 17.670 64.870 17.990 ;
        RECT 58.030 16.970 58.350 17.290 ;
        RECT 59.130 16.960 59.450 17.280 ;
        RECT 60.220 16.960 60.540 17.280 ;
        RECT 61.350 17.000 61.670 17.320 ;
        RECT 61.780 17.030 62.100 17.350 ;
        RECT 62.170 17.150 62.690 17.670 ;
        RECT 62.910 16.990 63.230 17.310 ;
        RECT 64.000 16.990 64.320 17.310 ;
        RECT 65.100 17.000 65.420 17.320 ;
        RECT 61.340 16.530 61.660 16.850 ;
        RECT 61.790 16.560 62.110 16.880 ;
        RECT 65.490 16.400 65.750 21.380 ;
        RECT 65.890 21.040 66.130 21.360 ;
        RECT 67.130 21.040 67.370 21.360 ;
        RECT 67.510 16.400 67.770 21.380 ;
        RECT 67.830 21.110 68.150 21.430 ;
        RECT 68.940 21.120 69.260 21.440 ;
        RECT 70.030 21.140 70.350 21.460 ;
        RECT 67.840 19.770 68.160 20.090 ;
        RECT 68.940 19.770 69.260 20.090 ;
        RECT 70.030 19.770 70.350 20.090 ;
        RECT 70.680 19.360 70.950 21.380 ;
        RECT 73.570 21.090 73.890 21.410 ;
        RECT 74.680 21.100 75.000 21.420 ;
        RECT 75.770 21.120 76.090 21.440 ;
        RECT 77.750 20.980 78.000 28.820 ;
        RECT 78.250 21.880 78.500 29.750 ;
        RECT 78.730 22.790 78.980 31.590 ;
        RECT 79.230 23.680 79.480 32.320 ;
        RECT 83.850 31.820 84.060 32.510 ;
        RECT 83.850 31.500 84.190 31.820 ;
        RECT 83.850 31.460 84.060 31.500 ;
        RECT 87.220 31.350 87.480 31.450 ;
        RECT 87.130 31.130 87.480 31.350 ;
        RECT 87.130 30.270 87.290 31.130 ;
        RECT 87.090 29.950 87.350 30.270 ;
        RECT 87.130 29.850 87.290 29.950 ;
        RECT 83.900 29.510 84.220 29.830 ;
        RECT 83.950 28.550 84.270 28.870 ;
        RECT 89.650 28.490 90.030 28.590 ;
        RECT 95.070 25.180 95.570 58.340 ;
        RECT 96.000 34.540 96.500 61.500 ;
        RECT 97.130 48.060 97.630 61.960 ;
        RECT 97.920 56.910 98.150 62.960 ;
        RECT 98.260 62.580 98.840 63.140 ;
        RECT 98.890 62.940 99.120 65.840 ;
        RECT 101.180 64.700 101.600 68.990 ;
        RECT 105.790 67.850 106.050 68.640 ;
        RECT 101.020 64.680 101.620 64.700 ;
        RECT 100.860 64.640 101.620 64.680 ;
        RECT 100.860 64.380 101.600 64.640 ;
        RECT 103.300 64.590 103.510 64.700 ;
        RECT 103.770 64.620 103.960 64.700 ;
        RECT 104.180 64.640 104.390 64.700 ;
        RECT 105.260 64.630 105.440 64.700 ;
        RECT 111.420 64.550 111.840 64.700 ;
        RECT 112.450 64.550 112.870 64.700 ;
        RECT 111.420 64.410 112.870 64.550 ;
        RECT 101.180 62.960 101.600 64.380 ;
        RECT 105.790 63.190 106.050 63.980 ;
        RECT 96.780 43.380 97.630 48.060 ;
        RECT 98.260 43.380 98.760 62.580 ;
        RECT 99.140 61.990 99.370 62.960 ;
        RECT 101.180 62.940 101.850 62.960 ;
        RECT 99.130 61.740 99.370 61.990 ;
        RECT 99.800 61.740 100.120 62.060 ;
        RECT 99.140 60.100 99.370 61.740 ;
        RECT 99.040 59.810 99.370 60.100 ;
        RECT 99.140 56.910 99.370 59.810 ;
        RECT 99.830 58.050 100.150 58.370 ;
        RECT 101.430 56.920 101.850 62.940 ;
        RECT 103.310 58.660 103.540 58.780 ;
        RECT 109.080 58.700 109.400 59.000 ;
        RECT 101.880 58.580 102.110 58.660 ;
        RECT 103.100 58.580 103.330 58.660 ;
        RECT 105.390 58.510 106.830 58.670 ;
        RECT 108.890 58.580 109.120 58.670 ;
        RECT 110.110 58.590 110.340 58.670 ;
        RECT 110.370 56.910 110.790 62.960 ;
        RECT 112.850 60.100 113.080 62.960 ;
        RECT 112.850 59.810 113.180 60.100 ;
        RECT 111.840 58.050 112.040 58.090 ;
        RECT 111.480 57.970 111.680 58.000 ;
        RECT 111.390 57.470 111.700 57.970 ;
        RECT 107.570 56.200 107.920 56.680 ;
        RECT 103.130 55.850 103.300 56.030 ;
        RECT 103.110 55.260 103.430 55.560 ;
        RECT 103.110 55.150 103.350 55.260 ;
        RECT 103.140 55.140 103.310 55.150 ;
        RECT 103.330 55.090 103.350 55.150 ;
        RECT 103.580 53.000 104.050 53.490 ;
        RECT 99.220 46.650 99.460 48.060 ;
        RECT 100.830 47.730 101.210 48.060 ;
        RECT 103.150 46.670 103.390 48.060 ;
        RECT 99.210 45.990 99.470 46.650 ;
        RECT 103.130 46.010 103.400 46.670 ;
        RECT 99.220 43.380 99.460 45.990 ;
        RECT 103.150 43.490 103.390 46.010 ;
        RECT 103.630 43.490 104.030 53.000 ;
        RECT 104.550 52.390 104.970 52.750 ;
        RECT 103.150 43.420 104.030 43.490 ;
        RECT 96.590 43.330 97.630 43.380 ;
        RECT 96.780 41.560 97.630 43.330 ;
        RECT 98.200 43.280 98.760 43.380 ;
        RECT 96.590 37.330 96.830 37.400 ;
        RECT 97.130 35.690 97.630 41.560 ;
        RECT 98.260 40.860 98.760 43.280 ;
        RECT 99.210 43.060 99.470 43.380 ;
        RECT 100.520 43.310 100.760 43.380 ;
        RECT 102.540 43.330 102.700 43.380 ;
        RECT 102.910 43.330 103.100 43.380 ;
        RECT 103.140 43.210 104.030 43.420 ;
        RECT 103.140 43.100 103.510 43.210 ;
        RECT 99.220 41.560 99.460 43.060 ;
        RECT 103.150 43.040 103.510 43.100 ;
        RECT 100.830 41.560 101.210 42.160 ;
        RECT 103.150 41.560 103.390 43.040 ;
        RECT 98.210 40.300 98.760 40.860 ;
        RECT 98.260 37.480 98.760 40.300 ;
        RECT 98.200 37.330 98.760 37.480 ;
        RECT 100.520 37.330 100.760 37.390 ;
        RECT 102.540 37.340 102.700 37.400 ;
        RECT 102.910 37.340 103.100 37.400 ;
        RECT 103.350 37.340 103.510 37.400 ;
        RECT 97.120 35.130 97.640 35.690 ;
        RECT 97.130 34.540 97.630 35.130 ;
        RECT 96.000 34.080 96.510 34.540 ;
        RECT 97.130 34.080 97.770 34.540 ;
        RECT 96.000 33.160 96.500 34.080 ;
        RECT 95.880 32.840 96.500 33.160 ;
        RECT 96.000 32.730 96.500 32.840 ;
        RECT 95.880 32.410 96.500 32.730 ;
        RECT 95.740 31.300 95.970 31.500 ;
        RECT 96.000 30.460 96.500 32.410 ;
        RECT 96.820 31.880 97.050 33.690 ;
        RECT 97.130 31.510 97.630 34.080 ;
        RECT 98.260 33.550 98.760 37.330 ;
        RECT 98.080 32.020 98.760 33.550 ;
        RECT 97.000 31.300 97.630 31.510 ;
        RECT 95.990 30.390 96.510 30.460 ;
        RECT 95.880 30.070 96.510 30.390 ;
        RECT 95.990 29.960 96.510 30.070 ;
        RECT 95.880 29.940 96.510 29.960 ;
        RECT 95.880 29.640 96.500 29.940 ;
        RECT 94.910 24.610 95.570 25.180 ;
        RECT 79.180 23.100 79.550 23.680 ;
        RECT 78.650 22.210 79.020 22.790 ;
        RECT 78.160 21.300 78.530 21.880 ;
        RECT 73.580 19.750 73.900 20.070 ;
        RECT 74.680 19.750 75.000 20.070 ;
        RECT 75.770 19.750 76.090 20.070 ;
        RECT 68.390 19.040 68.710 19.360 ;
        RECT 69.490 19.040 69.810 19.360 ;
        RECT 70.590 19.040 70.950 19.360 ;
        RECT 76.420 19.340 76.750 20.760 ;
        RECT 77.690 20.410 78.040 20.980 ;
        RECT 70.680 17.990 70.950 19.040 ;
        RECT 74.130 19.020 74.450 19.340 ;
        RECT 75.230 19.020 75.550 19.340 ;
        RECT 76.330 19.020 76.750 19.340 ;
        RECT 68.390 17.670 68.710 17.990 ;
        RECT 69.490 17.670 69.810 17.990 ;
        RECT 70.590 17.670 70.950 17.990 ;
        RECT 76.420 17.970 76.750 19.020 ;
        RECT 77.200 18.840 77.470 18.870 ;
        RECT 77.190 18.310 77.470 18.840 ;
        RECT 77.190 18.010 77.650 18.310 ;
        RECT 67.840 17.000 68.160 17.320 ;
        RECT 68.940 16.990 69.260 17.310 ;
        RECT 70.030 16.990 70.350 17.310 ;
        RECT 70.680 16.790 70.950 17.670 ;
        RECT 74.130 17.650 74.450 17.970 ;
        RECT 75.230 17.650 75.550 17.970 ;
        RECT 76.330 17.650 76.750 17.970 ;
        RECT 71.160 17.030 71.480 17.350 ;
        RECT 73.580 16.980 73.900 17.300 ;
        RECT 74.680 16.970 75.000 17.290 ;
        RECT 75.770 16.970 76.090 17.290 ;
        RECT 70.570 16.230 71.060 16.790 ;
        RECT 71.150 16.560 71.470 16.880 ;
        RECT 44.470 14.010 45.120 15.330 ;
        RECT 76.420 10.770 76.750 17.650 ;
        RECT 77.180 17.990 77.650 18.010 ;
        RECT 77.180 17.560 77.470 17.990 ;
        RECT 76.900 17.010 77.220 17.330 ;
        RECT 76.890 16.540 77.210 16.860 ;
        RECT 95.070 16.300 95.570 24.610 ;
        RECT 96.000 28.740 96.500 29.640 ;
        RECT 96.820 29.110 97.050 30.920 ;
        RECT 97.130 30.240 97.630 31.300 ;
        RECT 98.260 30.780 98.760 32.020 ;
        RECT 97.130 30.190 97.770 30.240 ;
        RECT 97.130 30.180 97.780 30.190 ;
        RECT 97.130 29.860 97.800 30.180 ;
        RECT 97.130 28.740 97.630 29.860 ;
        RECT 98.080 29.250 98.760 30.780 ;
        RECT 96.000 28.490 96.510 28.740 ;
        RECT 97.130 28.490 97.770 28.740 ;
        RECT 96.000 17.210 96.500 28.490 ;
        RECT 97.130 18.080 97.630 28.490 ;
        RECT 98.260 19.590 98.760 29.250 ;
        RECT 101.150 27.150 101.730 27.710 ;
        RECT 101.180 27.140 101.690 27.150 ;
        RECT 98.260 19.030 98.820 19.590 ;
        RECT 98.260 18.900 98.760 19.030 ;
        RECT 101.180 15.270 101.680 27.140 ;
        RECT 100.550 13.990 101.680 15.270 ;
        RECT 102.420 14.610 102.650 16.580 ;
        RECT 102.420 14.380 102.780 14.610 ;
        RECT 102.420 13.000 102.650 14.380 ;
        RECT 102.420 12.770 102.780 13.000 ;
        RECT 102.420 11.400 102.650 12.770 ;
        RECT 102.420 11.170 102.780 11.400 ;
        RECT 76.360 10.380 76.790 10.770 ;
        RECT 42.820 9.720 43.190 10.100 ;
        RECT 102.420 9.780 102.650 11.170 ;
        RECT 102.420 9.550 102.780 9.780 ;
        RECT 103.630 9.650 104.030 43.210 ;
        RECT 104.560 10.190 104.950 52.390 ;
        RECT 105.470 50.000 105.920 50.430 ;
        RECT 105.170 47.790 105.330 47.830 ;
        RECT 105.490 44.900 105.880 50.000 ;
        RECT 106.330 49.740 106.710 49.750 ;
        RECT 106.310 49.440 106.730 49.740 ;
        RECT 105.980 47.780 106.140 47.830 ;
        RECT 105.320 44.710 105.880 44.900 ;
        RECT 105.490 10.190 105.880 44.710 ;
        RECT 104.130 9.990 106.140 10.190 ;
        RECT 42.170 9.100 42.560 9.490 ;
        RECT 41.570 8.470 41.950 8.860 ;
        RECT 40.980 7.840 41.330 8.210 ;
        RECT 102.420 8.180 102.650 9.550 ;
        RECT 103.620 9.190 104.090 9.650 ;
        RECT 104.560 8.850 104.950 9.990 ;
        RECT 103.240 8.470 103.560 8.640 ;
        RECT 104.530 8.470 104.990 8.850 ;
        RECT 103.240 8.380 104.990 8.470 ;
        RECT 103.440 8.290 104.980 8.380 ;
        RECT 102.420 7.950 102.780 8.180 ;
        RECT 105.490 8.030 105.880 9.990 ;
        RECT 40.340 7.160 40.700 7.540 ;
        RECT 39.750 6.920 40.090 6.930 ;
        RECT 39.730 6.550 40.110 6.920 ;
        RECT 102.420 6.560 102.650 7.950 ;
        RECT 105.470 7.570 105.940 8.030 ;
        RECT 105.970 6.740 106.140 9.990 ;
        RECT 106.330 10.150 106.710 49.440 ;
        RECT 107.060 47.870 107.380 48.190 ;
        RECT 107.060 47.320 107.380 47.640 ;
        RECT 107.060 45.210 107.380 45.530 ;
        RECT 107.060 44.630 107.380 44.980 ;
        RECT 107.060 44.080 107.380 44.400 ;
        RECT 107.060 41.980 107.380 42.300 ;
        RECT 107.060 41.430 107.380 41.750 ;
        RECT 107.670 26.210 107.900 56.200 ;
        RECT 108.920 55.850 109.090 56.030 ;
        RECT 108.810 55.190 109.130 55.510 ;
        RECT 108.920 55.140 109.090 55.190 ;
        RECT 111.480 54.220 111.680 57.470 ;
        RECT 112.850 56.910 113.080 59.810 ;
        RECT 114.070 58.590 114.300 62.960 ;
        RECT 114.990 60.180 115.180 74.500 ;
        RECT 130.920 69.070 131.310 72.660 ;
        RECT 116.150 64.620 116.380 64.700 ;
        RECT 116.410 62.940 116.830 68.990 ;
        RECT 118.890 66.130 119.120 68.990 ;
        RECT 118.890 65.840 119.220 66.130 ;
        RECT 118.890 65.740 119.120 65.840 ;
        RECT 118.330 65.650 119.150 65.740 ;
        RECT 118.270 64.960 119.150 65.650 ;
        RECT 118.270 62.940 119.120 64.960 ;
        RECT 120.110 62.940 120.340 68.990 ;
        RECT 126.630 68.950 126.820 68.990 ;
        RECT 125.400 67.360 125.720 67.680 ;
        RECT 122.670 64.620 122.860 64.700 ;
        RECT 123.110 64.680 123.390 64.700 ;
        RECT 123.110 64.620 123.450 64.680 ;
        RECT 123.130 64.380 123.450 64.620 ;
        RECT 124.880 63.040 125.270 66.630 ;
        RECT 126.320 66.200 126.580 66.520 ;
        RECT 127.070 66.240 127.350 68.990 ;
        RECT 129.870 68.640 130.180 69.030 ;
        RECT 129.870 68.590 130.420 68.640 ;
        RECT 130.160 67.850 130.420 68.590 ;
        RECT 131.390 67.950 131.580 69.400 ;
        RECT 131.830 68.760 131.990 69.400 ;
        RECT 131.720 68.210 131.990 68.760 ;
        RECT 131.720 68.160 132.000 68.210 ;
        RECT 131.830 68.070 132.000 68.160 ;
        RECT 131.390 67.920 131.610 67.950 ;
        RECT 131.370 67.650 131.620 67.920 ;
        RECT 131.380 67.640 131.620 67.650 ;
        RECT 131.380 67.400 131.610 67.640 ;
        RECT 130.990 66.590 131.230 66.970 ;
        RECT 131.420 66.380 131.580 67.400 ;
        RECT 131.830 66.380 131.990 68.070 ;
        RECT 127.070 65.920 127.520 66.240 ;
        RECT 126.320 65.600 126.580 65.920 ;
        RECT 125.400 64.600 125.720 64.920 ;
        RECT 127.070 64.700 127.350 65.920 ;
        RECT 127.940 65.670 128.260 65.750 ;
        RECT 127.940 65.430 128.510 65.670 ;
        RECT 128.170 65.100 128.510 65.430 ;
        RECT 127.890 64.780 128.510 65.100 ;
        RECT 126.800 64.560 127.350 64.700 ;
        RECT 114.850 60.080 115.180 60.180 ;
        RECT 114.750 59.760 115.180 60.080 ;
        RECT 114.930 59.350 115.180 59.760 ;
        RECT 115.410 59.970 115.600 60.250 ;
        RECT 115.410 59.680 115.720 59.970 ;
        RECT 117.080 59.870 117.340 60.170 ;
        RECT 117.060 59.850 117.340 59.870 ;
        RECT 114.510 58.990 114.830 59.310 ;
        RECT 114.930 59.260 115.260 59.350 ;
        RECT 114.990 59.060 115.260 59.260 ;
        RECT 114.990 59.000 115.180 59.060 ;
        RECT 114.880 58.700 115.200 59.000 ;
        RECT 115.410 58.730 115.600 59.680 ;
        RECT 117.060 59.360 117.250 59.850 ;
        RECT 116.180 58.990 116.500 59.310 ;
        RECT 117.060 59.280 117.370 59.360 ;
        RECT 117.040 59.070 117.370 59.280 ;
        RECT 117.040 58.990 117.270 59.070 ;
        RECT 114.060 58.430 114.300 58.590 ;
        RECT 114.060 58.370 114.400 58.430 ;
        RECT 114.050 58.110 114.400 58.370 ;
        RECT 114.470 58.160 114.670 58.480 ;
        RECT 114.050 58.080 114.300 58.110 ;
        RECT 114.070 56.910 114.300 58.080 ;
        RECT 114.470 57.870 114.790 58.160 ;
        RECT 114.470 56.870 114.670 57.870 ;
        RECT 114.990 56.980 115.180 58.700 ;
        RECT 116.630 58.590 116.820 58.670 ;
        RECT 117.070 58.620 117.350 58.670 ;
        RECT 117.070 58.320 117.390 58.620 ;
        RECT 117.980 58.440 118.170 58.480 ;
        RECT 115.350 58.030 115.540 58.090 ;
        RECT 114.850 56.880 115.180 56.980 ;
        RECT 114.750 56.560 115.180 56.880 ;
        RECT 114.470 56.110 114.670 56.360 ;
        RECT 114.930 56.150 115.180 56.560 ;
        RECT 115.410 56.770 115.600 57.050 ;
        RECT 115.410 56.480 115.720 56.770 ;
        RECT 117.080 56.670 117.340 56.970 ;
        RECT 117.980 56.870 118.170 56.920 ;
        RECT 117.060 56.650 117.340 56.670 ;
        RECT 114.470 55.790 114.830 56.110 ;
        RECT 114.930 56.060 115.260 56.150 ;
        RECT 114.990 55.860 115.260 56.060 ;
        RECT 114.060 55.230 114.280 55.390 ;
        RECT 114.470 55.360 114.670 55.790 ;
        RECT 114.060 55.170 114.400 55.230 ;
        RECT 114.050 54.860 114.400 55.170 ;
        RECT 114.060 54.800 114.400 54.860 ;
        RECT 114.470 55.070 114.790 55.360 ;
        RECT 114.470 54.960 114.670 55.070 ;
        RECT 114.060 54.640 114.280 54.800 ;
        RECT 114.470 54.670 114.790 54.960 ;
        RECT 114.470 54.240 114.670 54.670 ;
        RECT 114.470 53.920 114.830 54.240 ;
        RECT 114.990 54.230 115.180 55.860 ;
        RECT 115.410 55.530 115.600 56.480 ;
        RECT 117.060 56.160 117.250 56.650 ;
        RECT 117.980 56.310 118.170 56.360 ;
        RECT 116.180 55.790 116.500 56.110 ;
        RECT 117.060 56.080 117.370 56.160 ;
        RECT 117.040 55.870 117.370 56.080 ;
        RECT 117.040 55.790 117.270 55.870 ;
        RECT 117.980 55.240 118.170 55.280 ;
        RECT 117.980 54.750 118.170 54.790 ;
        RECT 115.030 53.970 115.260 54.170 ;
        RECT 114.470 53.670 114.670 53.920 ;
        RECT 114.930 53.880 115.260 53.970 ;
        RECT 114.930 53.470 115.120 53.880 ;
        RECT 114.750 53.220 115.120 53.470 ;
        RECT 115.410 53.550 115.600 54.500 ;
        RECT 116.180 53.920 116.500 54.240 ;
        RECT 117.040 54.160 117.270 54.240 ;
        RECT 117.350 54.160 117.670 54.260 ;
        RECT 117.040 53.950 117.670 54.160 ;
        RECT 117.060 53.940 117.670 53.950 ;
        RECT 117.060 53.870 117.370 53.940 ;
        RECT 115.410 53.260 115.720 53.550 ;
        RECT 117.060 53.380 117.250 53.870 ;
        RECT 117.980 53.670 118.170 53.720 ;
        RECT 117.060 53.360 117.340 53.380 ;
        RECT 108.810 52.680 109.130 52.980 ;
        RECT 114.470 52.160 114.670 53.160 ;
        RECT 114.750 53.150 115.110 53.220 ;
        RECT 114.850 53.050 115.110 53.150 ;
        RECT 115.410 52.980 115.600 53.260 ;
        RECT 117.080 53.060 117.340 53.360 ;
        RECT 117.500 53.110 117.820 53.430 ;
        RECT 117.980 53.110 118.170 53.160 ;
        RECT 116.630 52.620 116.820 52.670 ;
        RECT 117.070 52.620 117.350 52.670 ;
        RECT 116.670 52.280 116.990 52.600 ;
        RECT 117.750 52.170 117.960 52.380 ;
        RECT 111.840 52.040 112.040 52.080 ;
        RECT 108.060 47.730 108.220 48.460 ;
        RECT 108.060 47.710 108.260 47.730 ;
        RECT 108.040 47.470 108.270 47.710 ;
        RECT 108.060 47.420 108.270 47.470 ;
        RECT 108.430 47.420 108.620 48.410 ;
        RECT 108.870 47.760 109.030 48.460 ;
        RECT 108.060 46.560 108.220 47.420 ;
        RECT 108.450 47.300 108.620 47.420 ;
        RECT 108.460 46.560 108.620 47.300 ;
        RECT 108.760 47.210 109.030 47.760 ;
        RECT 108.760 47.160 109.040 47.210 ;
        RECT 108.870 47.070 109.040 47.160 ;
        RECT 108.870 46.560 109.030 47.070 ;
        RECT 108.060 45.430 108.220 46.290 ;
        RECT 108.460 45.550 108.620 46.290 ;
        RECT 108.870 45.780 109.030 46.290 ;
        RECT 108.870 45.690 109.040 45.780 ;
        RECT 108.450 45.430 108.620 45.550 ;
        RECT 108.060 45.380 108.270 45.430 ;
        RECT 108.040 45.140 108.270 45.380 ;
        RECT 108.060 45.120 108.260 45.140 ;
        RECT 108.060 44.490 108.220 45.120 ;
        RECT 108.060 44.470 108.260 44.490 ;
        RECT 108.040 44.230 108.270 44.470 ;
        RECT 108.060 44.180 108.270 44.230 ;
        RECT 108.430 44.180 108.620 45.430 ;
        RECT 108.760 45.640 109.040 45.690 ;
        RECT 108.760 45.090 109.030 45.640 ;
        RECT 110.400 45.510 110.780 52.010 ;
        RECT 114.050 51.920 114.280 51.950 ;
        RECT 114.050 51.660 114.400 51.920 ;
        RECT 114.060 51.600 114.400 51.660 ;
        RECT 114.470 51.870 114.790 52.160 ;
        RECT 115.350 52.040 115.540 52.100 ;
        RECT 114.060 51.440 114.280 51.600 ;
        RECT 114.470 51.550 114.670 51.870 ;
        RECT 117.750 51.850 118.080 52.170 ;
        RECT 114.510 50.720 114.830 51.040 ;
        RECT 115.030 50.770 115.260 50.970 ;
        RECT 114.930 50.680 115.260 50.770 ;
        RECT 111.270 48.530 111.660 50.390 ;
        RECT 114.930 50.270 115.120 50.680 ;
        RECT 115.410 50.350 115.600 51.300 ;
        RECT 116.180 50.720 116.500 51.040 ;
        RECT 117.040 50.960 117.270 51.040 ;
        RECT 117.400 51.000 117.720 51.320 ;
        RECT 117.040 50.750 117.370 50.960 ;
        RECT 117.060 50.670 117.370 50.750 ;
        RECT 115.410 50.320 115.720 50.350 ;
        RECT 114.750 50.020 115.120 50.270 ;
        RECT 115.300 50.060 115.720 50.320 ;
        RECT 117.060 50.180 117.250 50.670 ;
        RECT 117.750 50.610 117.960 51.850 ;
        RECT 117.980 51.550 118.170 51.590 ;
        RECT 117.830 50.290 118.060 50.580 ;
        RECT 117.060 50.160 117.340 50.180 ;
        RECT 114.750 49.950 115.110 50.020 ;
        RECT 114.850 49.850 115.110 49.950 ;
        RECT 115.300 48.460 115.690 50.060 ;
        RECT 117.080 49.860 117.340 50.160 ;
        RECT 118.270 45.960 118.980 62.940 ;
        RECT 120.590 62.920 120.780 62.960 ;
        RECT 123.830 62.610 124.140 63.000 ;
        RECT 123.830 62.560 124.380 62.610 ;
        RECT 124.120 61.820 124.380 62.560 ;
        RECT 125.350 61.920 125.540 63.370 ;
        RECT 125.790 62.730 125.950 63.370 ;
        RECT 126.630 62.940 126.820 62.990 ;
        RECT 127.070 62.940 127.350 64.560 ;
        RECT 127.460 64.550 127.740 64.700 ;
        RECT 128.170 63.830 128.510 64.780 ;
        RECT 127.890 63.510 128.510 63.830 ;
        RECT 128.170 63.180 128.510 63.510 ;
        RECT 127.940 62.860 128.510 63.180 ;
        RECT 128.170 62.750 128.510 62.860 ;
        RECT 125.680 62.180 125.950 62.730 ;
        RECT 127.940 62.430 128.510 62.750 ;
        RECT 125.680 62.130 125.960 62.180 ;
        RECT 125.790 62.040 125.960 62.130 ;
        RECT 128.170 62.100 128.510 62.430 ;
        RECT 125.350 61.890 125.570 61.920 ;
        RECT 119.360 61.330 119.680 61.650 ;
        RECT 125.330 61.620 125.580 61.890 ;
        RECT 125.340 61.610 125.580 61.620 ;
        RECT 125.340 61.370 125.570 61.610 ;
        RECT 124.950 60.560 125.190 60.940 ;
        RECT 120.280 60.170 120.540 60.490 ;
        RECT 125.380 60.350 125.540 61.370 ;
        RECT 125.790 60.350 125.950 62.040 ;
        RECT 127.890 61.780 128.510 62.100 ;
        RECT 128.170 60.830 128.510 61.780 ;
        RECT 127.890 60.510 128.510 60.830 ;
        RECT 123.390 59.970 123.710 60.290 ;
        RECT 128.170 60.180 128.510 60.510 ;
        RECT 127.940 59.950 128.510 60.180 ;
        RECT 128.840 65.340 129.110 65.660 ;
        RECT 129.600 65.390 129.920 65.710 ;
        RECT 128.840 65.050 129.150 65.340 ;
        RECT 128.840 64.310 129.110 65.050 ;
        RECT 130.990 64.960 131.230 65.340 ;
        RECT 131.420 64.530 131.580 65.550 ;
        RECT 128.840 64.020 129.220 64.310 ;
        RECT 131.380 64.290 131.610 64.530 ;
        RECT 131.380 64.280 131.620 64.290 ;
        RECT 128.840 63.560 129.110 64.020 ;
        RECT 131.370 64.010 131.620 64.280 ;
        RECT 131.390 63.980 131.610 64.010 ;
        RECT 128.840 63.270 129.150 63.560 ;
        RECT 129.650 63.340 129.970 63.490 ;
        RECT 130.160 63.340 130.420 63.980 ;
        RECT 128.840 62.340 129.110 63.270 ;
        RECT 129.650 63.190 130.420 63.340 ;
        RECT 129.650 63.170 130.180 63.190 ;
        RECT 129.870 62.900 130.180 63.170 ;
        RECT 129.640 62.450 129.960 62.770 ;
        RECT 131.390 62.530 131.580 63.980 ;
        RECT 131.830 63.860 131.990 65.550 ;
        RECT 131.830 63.770 132.000 63.860 ;
        RECT 131.720 63.720 132.000 63.770 ;
        RECT 131.720 63.170 131.990 63.720 ;
        RECT 131.830 62.530 131.990 63.170 ;
        RECT 128.840 62.050 129.150 62.340 ;
        RECT 128.840 61.720 129.110 62.050 ;
        RECT 128.840 61.430 129.220 61.720 ;
        RECT 128.840 60.560 129.110 61.430 ;
        RECT 128.840 60.270 129.150 60.560 ;
        RECT 128.840 59.960 129.110 60.270 ;
        RECT 129.560 60.200 129.880 60.520 ;
        RECT 120.280 59.570 120.540 59.890 ;
        RECT 127.940 59.860 128.260 59.950 ;
        RECT 122.800 59.310 123.070 59.630 ;
        RECT 123.560 59.460 123.880 59.680 ;
        RECT 123.540 59.360 123.880 59.460 ;
        RECT 122.800 59.020 123.110 59.310 ;
        RECT 123.540 59.140 123.860 59.360 ;
        RECT 119.360 58.570 119.680 58.890 ;
        RECT 122.800 58.700 123.070 59.020 ;
        RECT 124.950 58.930 125.190 59.310 ;
        RECT 125.380 59.150 125.540 59.520 ;
        RECT 125.270 58.850 125.590 59.150 ;
        RECT 125.270 58.820 125.700 58.850 ;
        RECT 125.790 58.820 125.950 59.520 ;
        RECT 126.300 58.840 126.810 58.850 ;
        RECT 126.300 58.820 127.140 58.840 ;
        RECT 125.270 58.790 127.140 58.820 ;
        RECT 121.420 58.520 121.700 58.670 ;
        RECT 122.670 58.650 123.070 58.700 ;
        RECT 123.110 58.650 123.390 58.700 ;
        RECT 125.380 58.690 127.140 58.790 ;
        RECT 122.800 58.630 123.070 58.650 ;
        RECT 122.710 58.310 123.070 58.630 ;
        RECT 125.380 58.500 125.540 58.690 ;
        RECT 125.550 58.680 126.510 58.690 ;
        RECT 122.800 58.280 123.070 58.310 ;
        RECT 122.800 57.990 123.180 58.280 ;
        RECT 123.790 58.200 124.000 58.410 ;
        RECT 125.340 58.260 125.570 58.500 ;
        RECT 125.340 58.250 125.580 58.260 ;
        RECT 122.800 57.530 123.070 57.990 ;
        RECT 123.790 57.950 124.120 58.200 ;
        RECT 125.330 57.980 125.580 58.250 ;
        RECT 125.350 57.950 125.570 57.980 ;
        RECT 123.790 57.880 124.380 57.950 ;
        RECT 122.800 57.240 123.110 57.530 ;
        RECT 123.790 57.460 124.000 57.880 ;
        RECT 123.610 57.350 124.000 57.460 ;
        RECT 123.440 57.310 124.000 57.350 ;
        RECT 124.120 57.310 124.380 57.880 ;
        RECT 120.590 56.910 120.780 56.960 ;
        RECT 122.800 56.310 123.070 57.240 ;
        RECT 123.440 57.160 124.380 57.310 ;
        RECT 123.440 57.140 124.140 57.160 ;
        RECT 123.440 57.030 123.760 57.140 ;
        RECT 123.790 56.870 124.140 57.140 ;
        RECT 123.790 56.740 124.000 56.870 ;
        RECT 123.600 56.640 124.000 56.740 ;
        RECT 123.600 56.610 123.920 56.640 ;
        RECT 123.600 56.420 124.100 56.610 ;
        RECT 125.350 56.500 125.540 57.950 ;
        RECT 125.790 57.830 125.950 58.680 ;
        RECT 126.800 58.650 127.140 58.690 ;
        RECT 127.470 58.650 127.740 58.860 ;
        RECT 125.790 57.740 125.960 57.830 ;
        RECT 125.680 57.690 125.960 57.740 ;
        RECT 125.680 57.140 125.950 57.690 ;
        RECT 125.790 56.500 125.950 57.140 ;
        RECT 123.870 56.320 124.100 56.420 ;
        RECT 122.800 56.020 123.110 56.310 ;
        RECT 122.800 55.690 123.070 56.020 ;
        RECT 122.800 55.400 123.180 55.690 ;
        RECT 122.800 54.530 123.070 55.400 ;
        RECT 122.800 54.240 123.110 54.530 ;
        RECT 122.800 53.930 123.070 54.240 ;
        RECT 123.520 54.170 123.840 54.490 ;
        RECT 119.250 52.820 119.580 53.110 ;
        RECT 119.240 52.790 119.660 52.820 ;
        RECT 120.260 52.810 120.760 52.820 ;
        RECT 120.260 52.790 121.100 52.810 ;
        RECT 119.240 52.680 121.100 52.790 ;
        RECT 119.520 52.650 120.420 52.680 ;
        RECT 120.760 52.620 121.100 52.680 ;
        RECT 121.430 52.620 121.700 52.830 ;
        RECT 118.140 45.170 118.980 45.960 ;
        RECT 108.870 44.520 109.030 45.090 ;
        RECT 108.060 43.320 108.220 44.180 ;
        RECT 108.450 44.060 108.620 44.180 ;
        RECT 108.460 43.320 108.620 44.060 ;
        RECT 108.760 43.970 109.030 44.520 ;
        RECT 108.760 43.920 109.040 43.970 ;
        RECT 108.870 43.830 109.040 43.920 ;
        RECT 108.870 43.320 109.030 43.830 ;
        RECT 108.060 42.200 108.220 43.060 ;
        RECT 108.460 42.320 108.620 43.060 ;
        RECT 108.870 42.550 109.030 43.060 ;
        RECT 108.870 42.460 109.040 42.550 ;
        RECT 108.450 42.200 108.620 42.320 ;
        RECT 108.060 42.150 108.270 42.200 ;
        RECT 108.040 41.910 108.270 42.150 ;
        RECT 108.060 41.890 108.260 41.910 ;
        RECT 108.060 41.160 108.220 41.890 ;
        RECT 108.430 41.210 108.620 42.200 ;
        RECT 108.760 42.410 109.040 42.460 ;
        RECT 108.760 41.860 109.030 42.410 ;
        RECT 108.870 41.160 109.030 41.860 ;
        RECT 113.860 27.130 114.580 27.700 ;
        RECT 107.670 25.980 107.910 26.210 ;
        RECT 107.670 20.170 107.900 25.980 ;
        RECT 113.920 20.120 114.430 27.130 ;
        RECT 113.780 20.070 114.430 20.120 ;
        RECT 113.770 19.890 114.430 20.070 ;
        RECT 113.740 19.880 114.430 19.890 ;
        RECT 113.740 19.510 114.340 19.880 ;
        RECT 113.740 17.640 114.320 19.510 ;
        RECT 113.390 16.650 114.320 17.640 ;
        RECT 113.740 15.870 114.320 16.650 ;
        RECT 113.790 15.270 114.320 15.870 ;
        RECT 113.750 15.260 114.320 15.270 ;
        RECT 113.740 14.260 114.320 15.260 ;
        RECT 108.070 13.640 108.390 13.960 ;
        RECT 113.790 13.660 114.320 14.260 ;
        RECT 108.070 12.970 108.390 13.290 ;
        RECT 113.740 12.650 114.320 13.660 ;
        RECT 113.780 12.050 114.320 12.650 ;
        RECT 108.340 11.950 108.660 12.000 ;
        RECT 108.110 11.720 108.660 11.950 ;
        RECT 108.340 11.680 108.660 11.720 ;
        RECT 113.740 11.030 114.320 12.050 ;
        RECT 113.790 10.430 114.320 11.030 ;
        RECT 108.340 10.340 108.660 10.390 ;
        RECT 106.330 9.930 106.850 10.150 ;
        RECT 108.110 10.110 108.660 10.340 ;
        RECT 108.340 10.070 108.660 10.110 ;
        RECT 106.330 7.230 106.710 9.930 ;
        RECT 113.740 9.420 114.320 10.430 ;
        RECT 113.780 8.820 114.320 9.420 ;
        RECT 108.330 8.730 108.650 8.780 ;
        RECT 107.280 8.350 107.790 8.570 ;
        RECT 108.100 8.500 108.650 8.730 ;
        RECT 108.330 8.460 108.650 8.500 ;
        RECT 107.500 8.340 107.790 8.350 ;
        RECT 106.300 6.770 106.740 7.230 ;
        RECT 108.340 7.110 108.660 7.160 ;
        RECT 108.110 6.990 108.660 7.110 ;
        RECT 108.110 6.880 109.140 6.990 ;
        RECT 113.740 6.950 114.320 8.820 ;
        RECT 108.340 6.840 109.140 6.880 ;
        RECT 108.630 6.770 109.140 6.840 ;
        RECT 108.630 6.760 108.920 6.770 ;
        RECT 39.750 6.540 40.080 6.550 ;
        RECT 102.420 6.330 102.780 6.560 ;
        RECT 37.970 4.700 38.320 5.030 ;
        RECT 37.990 4.640 38.320 4.700 ;
        RECT 102.420 4.960 102.650 6.330 ;
        RECT 108.330 5.500 108.650 5.550 ;
        RECT 108.100 5.270 108.650 5.500 ;
        RECT 108.330 5.230 108.650 5.270 ;
        RECT 102.420 4.730 102.780 4.960 ;
        RECT 113.780 4.740 114.320 6.950 ;
        RECT 36.700 3.420 37.050 3.750 ;
        RECT 36.700 3.350 37.030 3.420 ;
        RECT 102.420 3.340 102.650 4.730 ;
        RECT 107.570 3.750 107.890 4.070 ;
        RECT 107.620 3.520 107.850 3.750 ;
        RECT 34.560 2.690 35.800 3.020 ;
        RECT 36.090 2.720 36.530 3.140 ;
        RECT 102.420 3.110 102.780 3.340 ;
        RECT 102.420 3.040 102.650 3.110 ;
        RECT 34.560 2.580 35.140 2.690 ;
        RECT 108.330 2.300 108.650 2.350 ;
        RECT 108.100 2.070 108.650 2.300 ;
        RECT 108.330 2.030 108.650 2.070 ;
        RECT 105.090 0.590 105.410 0.640 ;
        RECT 106.030 0.590 106.350 0.640 ;
        RECT 104.860 0.360 105.410 0.590 ;
        RECT 105.800 0.360 106.350 0.590 ;
        RECT 106.980 0.570 107.300 0.620 ;
        RECT 108.290 0.590 108.610 0.640 ;
        RECT 105.090 0.320 105.410 0.360 ;
        RECT 106.030 0.320 106.350 0.360 ;
        RECT 106.750 0.340 107.300 0.570 ;
        RECT 108.060 0.360 108.610 0.590 ;
        RECT 106.980 0.300 107.300 0.340 ;
        RECT 108.290 0.320 108.610 0.360 ;
      LAYER via ;
        RECT 7.510 72.460 7.900 72.850 ;
        RECT 1.000 69.050 1.260 69.310 ;
        RECT 3.860 69.100 4.120 69.360 ;
        RECT 7.590 69.010 7.980 69.400 ;
        RECT 0.990 68.020 1.250 68.280 ;
        RECT 1.660 68.040 1.920 68.300 ;
        RECT 2.400 68.030 2.660 68.290 ;
        RECT 0.990 67.570 1.250 67.830 ;
        RECT 2.400 67.590 2.660 67.850 ;
        RECT 0.990 67.150 1.250 67.410 ;
        RECT 1.660 67.200 1.920 67.460 ;
        RECT 2.420 67.170 2.680 67.430 ;
        RECT 0.990 65.800 1.250 66.060 ;
        RECT 3.550 67.720 3.810 67.980 ;
        RECT 3.360 65.300 3.620 65.560 ;
        RECT 1.640 64.400 1.900 64.660 ;
        RECT 3.070 64.420 3.330 64.680 ;
        RECT 0.850 63.820 1.110 64.080 ;
        RECT 1.780 63.820 2.040 64.080 ;
        RECT 2.480 63.820 2.740 64.080 ;
        RECT 3.220 63.820 3.480 64.080 ;
        RECT 3.930 63.810 4.190 64.070 ;
        RECT 8.970 67.840 9.230 68.100 ;
        RECT 17.050 67.300 17.310 67.560 ;
        RECT 18.410 67.380 18.670 67.640 ;
        RECT 19.100 67.370 19.360 67.630 ;
        RECT 8.890 65.140 9.310 65.560 ;
        RECT 14.840 63.740 15.130 64.320 ;
        RECT 16.330 63.640 16.590 63.900 ;
        RECT 26.190 63.660 26.450 63.920 ;
        RECT 28.130 62.680 28.390 62.940 ;
        RECT 22.550 59.000 22.810 59.260 ;
        RECT 23.640 59.010 23.900 59.270 ;
        RECT 21.010 58.090 21.270 58.350 ;
        RECT 22.560 58.010 22.820 58.270 ;
        RECT 20.990 57.170 21.250 57.430 ;
        RECT 20.970 56.180 21.230 56.440 ;
        RECT 22.560 57.020 22.820 57.280 ;
        RECT 22.050 56.430 22.310 56.690 ;
        RECT 22.470 56.290 22.730 56.550 ;
        RECT 22.020 55.510 22.280 55.770 ;
        RECT 22.560 55.590 22.820 55.850 ;
        RECT 22.470 55.300 22.730 55.560 ;
        RECT 22.030 54.590 22.290 54.850 ;
        RECT 22.560 54.600 22.820 54.860 ;
        RECT 21.380 53.570 21.640 53.830 ;
        RECT 21.340 52.610 21.600 52.870 ;
        RECT 21.380 51.650 21.640 51.910 ;
        RECT 22.470 54.310 22.730 54.570 ;
        RECT 23.650 58.020 23.910 58.280 ;
        RECT 22.560 53.610 22.820 53.870 ;
        RECT 23.650 57.030 23.910 57.290 ;
        RECT 33.920 62.250 34.230 62.560 ;
        RECT 50.500 69.890 50.920 70.310 ;
        RECT 46.650 69.130 47.070 69.550 ;
        RECT 52.170 67.520 52.610 67.960 ;
        RECT 57.890 67.520 58.330 67.960 ;
        RECT 59.710 67.490 60.150 67.930 ;
        RECT 47.750 66.500 48.190 66.940 ;
        RECT 44.990 63.480 45.250 63.740 ;
        RECT 37.920 62.790 38.180 63.050 ;
        RECT 36.750 61.800 37.020 62.060 ;
        RECT 25.420 61.020 25.770 61.370 ;
        RECT 30.670 61.330 30.930 61.590 ;
        RECT 46.600 61.460 46.860 61.720 ;
        RECT 46.600 59.710 46.860 59.970 ;
        RECT 48.700 62.300 48.960 62.560 ;
        RECT 49.640 61.820 49.900 62.080 ;
        RECT 50.680 61.860 50.940 62.120 ;
        RECT 50.740 61.580 51.000 61.840 ;
        RECT 48.700 60.550 48.960 60.810 ;
        RECT 49.640 60.070 49.900 60.330 ;
        RECT 50.680 60.110 50.940 60.370 ;
        RECT 50.740 59.830 51.000 60.090 ;
        RECT 26.440 58.780 26.700 59.170 ;
        RECT 42.840 58.790 43.170 59.050 ;
        RECT 25.800 57.960 26.060 58.360 ;
        RECT 25.820 56.850 26.080 57.110 ;
        RECT 23.770 56.190 24.030 56.450 ;
        RECT 25.820 55.930 26.080 56.190 ;
        RECT 23.770 55.200 24.030 55.460 ;
        RECT 25.790 55.010 26.050 55.270 ;
        RECT 23.770 54.210 24.030 54.470 ;
        RECT 21.340 36.370 21.600 36.840 ;
        RECT 21.980 36.370 22.240 36.840 ;
        RECT 19.980 35.340 20.240 35.600 ;
        RECT 19.460 34.940 19.720 35.200 ;
        RECT 10.180 33.690 10.840 34.350 ;
        RECT 22.060 35.320 22.320 35.580 ;
        RECT 23.820 35.330 24.090 35.600 ;
        RECT 21.400 34.960 21.660 35.220 ;
        RECT 19.480 31.030 19.740 31.290 ;
        RECT 15.390 29.170 15.760 29.540 ;
        RECT 10.220 27.830 10.880 28.490 ;
        RECT 19.340 27.790 19.600 28.050 ;
        RECT 24.320 34.940 24.580 35.200 ;
        RECT 22.650 28.230 22.910 28.490 ;
        RECT 20.440 27.800 20.700 28.060 ;
        RECT 21.530 27.800 21.790 28.060 ;
        RECT 22.660 27.760 22.920 28.020 ;
        RECT 19.890 27.120 20.150 27.380 ;
        RECT 20.990 27.120 21.250 27.380 ;
        RECT 22.090 27.120 22.350 27.380 ;
        RECT 19.890 25.750 20.150 26.010 ;
        RECT 20.990 25.750 21.250 26.010 ;
        RECT 22.090 25.750 22.350 26.010 ;
        RECT 19.340 25.020 19.600 25.280 ;
        RECT 20.440 25.020 20.700 25.280 ;
        RECT 21.530 25.020 21.790 25.280 ;
        RECT 19.330 23.680 19.590 23.940 ;
        RECT 20.440 23.670 20.700 23.930 ;
        RECT 21.530 23.650 21.790 23.910 ;
        RECT 15.380 22.930 15.750 23.300 ;
        RECT 19.890 22.980 20.150 23.240 ;
        RECT 20.990 22.970 21.250 23.230 ;
        RECT 22.080 22.970 22.340 23.230 ;
        RECT 22.920 22.510 23.180 22.870 ;
        RECT 18.370 17.270 18.660 17.560 ;
        RECT 22.690 20.670 22.950 20.930 ;
        RECT 19.380 20.230 19.640 20.490 ;
        RECT 20.480 20.240 20.740 20.500 ;
        RECT 21.570 20.240 21.830 20.500 ;
        RECT 22.700 20.200 22.960 20.460 ;
        RECT 19.930 19.560 20.190 19.820 ;
        RECT 21.030 19.560 21.290 19.820 ;
        RECT 22.130 19.560 22.390 19.820 ;
        RECT 19.930 18.190 20.190 18.450 ;
        RECT 21.030 18.190 21.290 18.450 ;
        RECT 22.130 18.190 22.390 18.450 ;
        RECT 19.380 17.460 19.640 17.720 ;
        RECT 20.480 17.460 20.740 17.720 ;
        RECT 21.570 17.460 21.830 17.720 ;
        RECT 42.210 57.070 42.540 57.400 ;
        RECT 41.640 55.590 41.970 55.920 ;
        RECT 26.430 53.920 26.690 54.180 ;
        RECT 41.000 53.990 41.330 54.320 ;
        RECT 40.360 53.420 40.690 53.750 ;
        RECT 26.440 52.960 26.700 53.220 ;
        RECT 26.430 52.000 26.690 52.260 ;
        RECT 25.790 34.340 26.050 34.600 ;
        RECT 25.170 33.190 25.430 33.450 ;
        RECT 25.740 32.580 26.000 32.840 ;
        RECT 25.240 31.280 25.500 31.540 ;
        RECT 24.750 30.580 25.010 30.840 ;
        RECT 25.240 29.730 25.500 29.990 ;
        RECT 39.750 51.850 40.080 52.180 ;
        RECT 39.120 50.320 39.450 50.650 ;
        RECT 38.560 48.750 38.890 49.080 ;
        RECT 37.940 43.280 38.270 43.610 ;
        RECT 37.310 41.690 37.640 42.020 ;
        RECT 36.690 40.140 37.020 40.470 ;
        RECT 36.090 38.660 36.420 38.990 ;
        RECT 35.450 33.490 35.780 33.820 ;
        RECT 26.960 33.020 27.220 33.280 ;
        RECT 27.610 33.020 27.870 33.280 ;
        RECT 26.440 32.580 26.700 32.840 ;
        RECT 27.980 32.000 28.240 32.260 ;
        RECT 34.780 31.920 35.110 32.250 ;
        RECT 27.640 30.780 27.900 31.040 ;
        RECT 26.430 30.010 26.690 30.270 ;
        RECT 27.650 30.240 27.910 30.500 ;
        RECT 34.160 30.280 34.490 30.610 ;
        RECT 25.770 28.700 26.030 28.960 ;
        RECT 27.960 29.380 28.220 29.640 ;
        RECT 26.460 28.690 26.720 28.950 ;
        RECT 33.480 28.840 33.810 29.170 ;
        RECT 25.190 24.890 25.450 25.310 ;
        RECT 25.150 22.510 25.410 22.870 ;
        RECT 25.770 18.880 26.030 19.210 ;
        RECT 24.740 17.260 25.030 17.550 ;
        RECT 19.370 16.120 19.630 16.380 ;
        RECT 20.480 16.110 20.740 16.370 ;
        RECT 21.570 16.090 21.830 16.350 ;
        RECT 23.580 16.250 24.180 16.850 ;
        RECT 19.930 15.420 20.190 15.680 ;
        RECT 21.030 15.410 21.290 15.670 ;
        RECT 22.120 15.410 22.380 15.670 ;
        RECT 26.940 27.920 27.200 28.180 ;
        RECT 27.650 27.860 27.910 28.120 ;
        RECT 29.440 24.480 30.020 25.190 ;
        RECT 26.360 11.320 26.620 11.660 ;
        RECT 7.450 10.380 7.840 10.770 ;
        RECT 33.450 5.010 33.880 5.440 ;
        RECT 34.100 4.220 34.530 4.650 ;
        RECT 34.770 3.540 35.170 3.940 ;
        RECT 34.600 2.600 35.110 3.110 ;
        RECT 46.600 57.960 46.860 58.220 ;
        RECT 48.700 58.800 48.960 59.060 ;
        RECT 49.640 58.320 49.900 58.580 ;
        RECT 50.680 58.360 50.940 58.620 ;
        RECT 50.740 58.080 51.000 58.340 ;
        RECT 46.600 56.210 46.860 56.470 ;
        RECT 48.700 57.050 48.960 57.310 ;
        RECT 49.640 56.570 49.900 56.830 ;
        RECT 50.680 56.610 50.940 56.870 ;
        RECT 50.740 56.330 51.000 56.590 ;
        RECT 53.460 66.500 53.900 66.940 ;
        RECT 70.270 69.130 71.620 69.550 ;
        RECT 64.850 66.490 65.800 66.900 ;
        RECT 67.860 66.500 68.300 66.940 ;
        RECT 62.110 62.720 62.370 62.980 ;
        RECT 60.230 59.190 60.490 59.450 ;
        RECT 65.700 61.810 65.960 62.070 ;
        RECT 62.570 60.790 62.830 61.050 ;
        RECT 62.990 58.700 63.250 58.960 ;
        RECT 64.050 58.220 64.310 58.480 ;
        RECT 68.870 62.730 69.130 62.990 ;
        RECT 68.430 61.820 68.690 62.080 ;
        RECT 62.540 52.910 62.800 53.170 ;
        RECT 46.600 51.440 46.860 51.700 ;
        RECT 49.640 51.080 49.900 51.340 ;
        RECT 48.700 50.600 48.960 50.860 ;
        RECT 50.740 51.320 51.000 51.580 ;
        RECT 50.680 51.040 50.940 51.300 ;
        RECT 46.600 49.690 46.860 49.950 ;
        RECT 49.640 49.330 49.900 49.590 ;
        RECT 48.700 48.850 48.960 49.110 ;
        RECT 50.740 49.570 51.000 49.830 ;
        RECT 50.680 49.290 50.940 49.550 ;
        RECT 46.600 47.940 46.860 48.200 ;
        RECT 46.600 46.190 46.860 46.450 ;
        RECT 49.640 47.580 49.900 47.840 ;
        RECT 48.700 47.100 48.960 47.360 ;
        RECT 50.740 47.820 51.000 48.080 ;
        RECT 50.680 47.540 50.940 47.800 ;
        RECT 49.640 45.830 49.900 46.090 ;
        RECT 48.700 45.350 48.960 45.610 ;
        RECT 50.740 46.070 51.000 46.330 ;
        RECT 50.680 45.790 50.940 46.050 ;
        RECT 61.450 52.390 61.710 52.650 ;
        RECT 61.450 52.020 61.710 52.280 ;
        RECT 62.540 51.500 62.800 51.760 ;
        RECT 64.950 52.910 65.210 53.170 ;
        RECT 64.950 51.500 65.210 51.760 ;
        RECT 65.690 51.120 65.960 51.390 ;
        RECT 62.540 49.710 62.800 49.970 ;
        RECT 61.450 49.190 61.710 49.450 ;
        RECT 61.450 48.820 61.710 49.080 ;
        RECT 62.540 48.300 62.800 48.560 ;
        RECT 64.950 49.710 65.210 49.970 ;
        RECT 64.950 48.300 65.210 48.560 ;
        RECT 73.660 66.460 74.100 66.900 ;
        RECT 81.990 67.490 82.270 67.930 ;
        RECT 78.210 60.830 79.430 61.090 ;
        RECT 74.970 60.180 75.230 60.440 ;
        RECT 81.300 59.640 81.560 59.900 ;
        RECT 83.640 62.730 83.900 62.990 ;
        RECT 82.750 61.860 83.010 62.120 ;
        RECT 90.160 71.830 90.530 72.200 ;
        RECT 87.850 68.620 88.110 68.880 ;
        RECT 86.310 63.440 86.570 63.710 ;
        RECT 87.850 63.050 88.110 63.310 ;
        RECT 88.100 62.590 88.360 62.850 ;
        RECT 82.750 57.650 83.010 57.910 ;
        RECT 83.770 57.660 84.030 57.920 ;
        RECT 86.520 57.540 86.950 57.970 ;
        RECT 88.100 57.020 88.360 57.280 ;
        RECT 80.270 47.900 80.530 48.160 ;
        RECT 90.980 68.370 91.350 68.740 ;
        RECT 92.080 66.820 92.340 67.080 ;
        RECT 91.420 65.940 91.680 66.200 ;
        RECT 92.070 65.130 92.330 65.390 ;
        RECT 91.750 63.660 92.120 64.030 ;
        RECT 92.570 61.360 92.830 61.620 ;
        RECT 95.080 61.050 95.580 61.550 ;
        RECT 96.030 61.540 96.530 62.040 ;
        RECT 97.110 62.010 97.610 62.510 ;
        RECT 91.680 60.200 91.940 60.460 ;
        RECT 91.680 59.600 91.940 59.860 ;
        RECT 80.270 47.350 80.530 47.610 ;
        RECT 62.330 44.480 62.610 44.760 ;
        RECT 80.270 45.240 80.530 45.500 ;
        RECT 80.270 44.660 80.530 44.950 ;
        RECT 79.680 43.910 79.940 44.170 ;
        RECT 80.270 44.110 80.530 44.370 ;
        RECT 83.990 43.390 84.250 43.470 ;
        RECT 83.990 43.210 84.480 43.390 ;
        RECT 90.170 44.460 90.540 44.830 ;
        RECT 90.940 43.870 91.310 44.240 ;
        RECT 62.520 42.440 62.780 42.700 ;
        RECT 46.600 41.310 46.860 41.570 ;
        RECT 49.640 40.950 49.900 41.210 ;
        RECT 48.700 40.470 48.960 40.730 ;
        RECT 50.740 41.190 51.000 41.450 ;
        RECT 50.680 40.910 50.940 41.170 ;
        RECT 46.600 39.560 46.860 39.820 ;
        RECT 49.640 39.200 49.900 39.460 ;
        RECT 48.700 38.720 48.960 38.980 ;
        RECT 50.740 39.440 51.000 39.700 ;
        RECT 50.680 39.160 50.940 39.420 ;
        RECT 46.600 37.810 46.860 38.070 ;
        RECT 49.640 37.450 49.900 37.710 ;
        RECT 48.700 36.970 48.960 37.230 ;
        RECT 46.600 36.060 46.860 36.320 ;
        RECT 50.740 37.690 51.000 37.950 ;
        RECT 50.680 37.410 50.940 37.670 ;
        RECT 49.640 35.700 49.900 35.960 ;
        RECT 48.700 35.220 48.960 35.480 ;
        RECT 50.740 35.940 51.000 36.200 ;
        RECT 50.680 35.660 50.940 35.920 ;
        RECT 61.430 41.920 61.690 42.180 ;
        RECT 61.430 41.550 61.690 41.810 ;
        RECT 62.520 41.030 62.780 41.290 ;
        RECT 64.930 42.440 65.190 42.700 ;
        RECT 64.930 41.030 65.190 41.290 ;
        RECT 62.520 39.240 62.780 39.500 ;
        RECT 61.430 38.720 61.690 38.980 ;
        RECT 61.430 38.350 61.690 38.610 ;
        RECT 54.960 36.290 55.220 36.700 ;
        RECT 62.520 37.830 62.780 38.090 ;
        RECT 64.930 39.240 65.190 39.500 ;
        RECT 64.930 37.830 65.190 38.090 ;
        RECT 46.560 32.250 46.820 32.510 ;
        RECT 49.600 31.890 49.860 32.150 ;
        RECT 48.660 31.410 48.920 31.670 ;
        RECT 50.700 32.130 50.960 32.390 ;
        RECT 50.640 31.850 50.900 32.110 ;
        RECT 46.560 30.500 46.820 30.760 ;
        RECT 49.600 30.140 49.860 30.400 ;
        RECT 48.660 29.660 48.920 29.920 ;
        RECT 50.700 30.380 50.960 30.640 ;
        RECT 50.640 30.100 50.900 30.360 ;
        RECT 46.560 28.750 46.820 29.010 ;
        RECT 49.600 28.390 49.860 28.650 ;
        RECT 46.560 27.000 46.820 27.260 ;
        RECT 48.660 27.910 48.920 28.170 ;
        RECT 50.700 28.630 50.960 28.890 ;
        RECT 50.640 28.350 50.900 28.610 ;
        RECT 47.800 26.560 48.110 26.870 ;
        RECT 49.600 26.640 49.860 26.900 ;
        RECT 48.660 26.160 48.920 26.420 ;
        RECT 50.700 26.880 50.960 27.140 ;
        RECT 50.640 26.600 50.900 26.860 ;
        RECT 62.550 33.170 62.810 33.430 ;
        RECT 59.360 32.570 59.620 32.830 ;
        RECT 61.460 32.650 61.720 32.910 ;
        RECT 52.780 27.440 53.040 27.700 ;
        RECT 52.240 27.070 52.530 27.360 ;
        RECT 61.460 32.280 61.720 32.540 ;
        RECT 62.550 31.760 62.810 32.020 ;
        RECT 64.960 33.170 65.220 33.430 ;
        RECT 64.960 31.760 65.220 32.020 ;
        RECT 84.220 43.130 84.480 43.210 ;
        RECT 88.150 43.090 88.410 43.350 ;
        RECT 80.270 42.010 80.530 42.270 ;
        RECT 80.270 41.460 80.530 41.720 ;
        RECT 92.630 58.860 93.000 58.960 ;
        RECT 92.570 58.600 93.000 58.860 ;
        RECT 92.630 58.590 93.000 58.600 ;
        RECT 91.680 41.540 92.050 41.910 ;
        RECT 80.870 39.060 81.130 39.320 ;
        RECT 80.870 38.510 81.130 38.770 ;
        RECT 80.870 36.420 81.130 36.680 ;
        RECT 80.870 35.820 81.130 36.130 ;
        RECT 80.870 35.270 81.130 35.530 ;
        RECT 84.940 34.210 85.200 34.470 ;
        RECT 79.240 32.550 79.500 32.810 ;
        RECT 80.870 33.170 81.130 33.430 ;
        RECT 80.870 32.620 81.130 32.880 ;
        RECT 83.950 32.540 84.210 32.800 ;
        RECT 87.240 34.090 87.500 34.350 ;
        RECT 88.960 34.190 89.230 34.450 ;
        RECT 87.220 33.040 87.480 33.300 ;
        RECT 94.900 58.350 95.160 58.610 ;
        RECT 92.610 36.290 92.980 36.700 ;
        RECT 78.720 31.620 78.980 31.880 ;
        RECT 59.990 29.790 60.250 30.050 ;
        RECT 59.390 27.480 59.650 27.740 ;
        RECT 60.420 27.470 60.680 27.730 ;
        RECT 57.990 27.070 58.250 27.330 ;
        RECT 59.960 27.150 60.220 27.410 ;
        RECT 51.610 25.850 52.030 26.270 ;
        RECT 47.760 24.890 48.180 25.310 ;
        RECT 53.670 26.530 53.930 26.790 ;
        RECT 62.550 29.970 62.810 30.230 ;
        RECT 61.460 29.450 61.720 29.710 ;
        RECT 61.460 29.080 61.720 29.340 ;
        RECT 62.550 28.560 62.810 28.820 ;
        RECT 64.960 29.970 65.220 30.230 ;
        RECT 64.960 28.560 65.220 28.820 ;
        RECT 78.250 29.780 78.510 30.040 ;
        RECT 77.750 28.850 78.010 29.110 ;
        RECT 62.200 27.090 62.460 27.350 ;
        RECT 61.000 25.840 61.330 26.170 ;
        RECT 71.040 27.400 71.390 27.750 ;
        RECT 64.190 26.670 64.450 26.930 ;
        RECT 68.230 26.640 68.500 26.910 ;
        RECT 62.150 25.770 62.490 26.110 ;
        RECT 71.080 25.630 71.340 25.950 ;
        RECT 77.070 25.850 77.330 26.190 ;
        RECT 52.290 24.800 52.610 25.120 ;
        RECT 72.500 24.920 72.880 25.300 ;
        RECT 52.580 21.820 52.840 22.080 ;
        RECT 53.670 21.820 53.930 22.080 ;
        RECT 54.770 21.810 55.030 22.070 ;
        RECT 53.130 21.140 53.390 21.400 ;
        RECT 54.220 21.120 54.480 21.380 ;
        RECT 55.330 21.110 55.590 21.370 ;
        RECT 58.610 21.810 58.870 22.070 ;
        RECT 59.710 21.820 59.970 22.080 ;
        RECT 60.800 21.820 61.060 22.080 ;
        RECT 62.390 21.850 62.650 22.110 ;
        RECT 63.480 21.850 63.740 22.110 ;
        RECT 64.580 21.840 64.840 22.100 ;
        RECT 53.130 19.770 53.390 20.030 ;
        RECT 54.220 19.770 54.480 20.030 ;
        RECT 55.320 19.770 55.580 20.030 ;
        RECT 52.390 19.020 52.850 19.480 ;
        RECT 53.670 19.040 53.930 19.300 ;
        RECT 54.770 19.040 55.030 19.300 ;
        RECT 52.570 17.670 52.830 17.930 ;
        RECT 53.670 17.670 53.930 17.930 ;
        RECT 54.770 17.670 55.030 17.930 ;
        RECT 52.000 17.030 52.260 17.290 ;
        RECT 53.130 16.990 53.390 17.250 ;
        RECT 54.220 16.990 54.480 17.250 ;
        RECT 55.320 17.000 55.580 17.260 ;
        RECT 52.010 16.560 52.270 16.820 ;
        RECT 58.050 21.110 58.310 21.370 ;
        RECT 59.160 21.120 59.420 21.380 ;
        RECT 60.250 21.140 60.510 21.400 ;
        RECT 58.060 19.770 58.320 20.030 ;
        RECT 59.160 19.770 59.420 20.030 ;
        RECT 60.250 19.770 60.510 20.030 ;
        RECT 58.610 19.040 58.870 19.300 ;
        RECT 59.710 19.040 59.970 19.300 ;
        RECT 60.810 19.040 61.070 19.300 ;
        RECT 62.940 21.170 63.200 21.430 ;
        RECT 64.030 21.150 64.290 21.410 ;
        RECT 65.140 21.140 65.400 21.400 ;
        RECT 68.420 21.840 68.680 22.100 ;
        RECT 69.520 21.850 69.780 22.110 ;
        RECT 70.610 21.850 70.870 22.110 ;
        RECT 74.160 21.820 74.420 22.080 ;
        RECT 75.260 21.830 75.520 22.090 ;
        RECT 76.350 21.830 76.610 22.090 ;
        RECT 62.940 19.800 63.200 20.060 ;
        RECT 64.030 19.800 64.290 20.060 ;
        RECT 65.130 19.800 65.390 20.060 ;
        RECT 62.380 19.070 62.640 19.330 ;
        RECT 63.480 19.070 63.740 19.330 ;
        RECT 64.580 19.070 64.840 19.330 ;
        RECT 60.770 18.070 61.230 18.530 ;
        RECT 58.610 17.670 58.870 17.930 ;
        RECT 59.710 17.670 59.970 17.930 ;
        RECT 60.810 17.670 61.070 17.930 ;
        RECT 62.380 17.700 62.640 17.960 ;
        RECT 63.480 17.700 63.740 17.960 ;
        RECT 64.580 17.700 64.840 17.960 ;
        RECT 58.060 17.000 58.320 17.260 ;
        RECT 59.160 16.990 59.420 17.250 ;
        RECT 60.250 16.990 60.510 17.250 ;
        RECT 61.380 17.030 61.640 17.290 ;
        RECT 61.810 17.060 62.070 17.320 ;
        RECT 62.200 17.180 62.660 17.640 ;
        RECT 62.940 17.020 63.200 17.280 ;
        RECT 64.030 17.020 64.290 17.280 ;
        RECT 65.130 17.030 65.390 17.290 ;
        RECT 61.370 16.560 61.630 16.820 ;
        RECT 61.820 16.590 62.080 16.850 ;
        RECT 67.860 21.140 68.120 21.400 ;
        RECT 68.970 21.150 69.230 21.410 ;
        RECT 70.060 21.170 70.320 21.430 ;
        RECT 67.870 19.800 68.130 20.060 ;
        RECT 68.970 19.800 69.230 20.060 ;
        RECT 70.060 19.800 70.320 20.060 ;
        RECT 73.600 21.120 73.860 21.380 ;
        RECT 74.710 21.130 74.970 21.390 ;
        RECT 75.800 21.150 76.060 21.410 ;
        RECT 83.930 31.530 84.190 31.790 ;
        RECT 87.220 31.160 87.480 31.420 ;
        RECT 87.090 29.980 87.350 30.240 ;
        RECT 83.930 29.540 84.190 29.800 ;
        RECT 83.980 28.580 84.240 28.840 ;
        RECT 98.300 62.610 98.800 63.110 ;
        RECT 100.890 64.400 101.150 64.660 ;
        RECT 99.830 61.770 100.090 62.030 ;
        RECT 99.860 58.080 100.120 58.340 ;
        RECT 109.110 58.720 109.370 58.980 ;
        RECT 111.430 57.510 111.690 57.940 ;
        RECT 107.600 56.230 107.860 56.650 ;
        RECT 103.140 55.280 103.400 55.540 ;
        RECT 103.600 53.030 104.000 53.430 ;
        RECT 104.580 52.390 104.940 52.750 ;
        RECT 103.390 43.390 103.650 43.480 ;
        RECT 99.210 43.090 99.470 43.350 ;
        RECT 103.140 43.220 103.650 43.390 ;
        RECT 103.140 43.130 103.400 43.220 ;
        RECT 98.210 40.330 98.710 40.830 ;
        RECT 97.130 35.140 97.630 35.610 ;
        RECT 96.060 33.130 96.320 33.380 ;
        RECT 95.910 33.120 96.320 33.130 ;
        RECT 95.910 32.870 96.170 33.120 ;
        RECT 95.910 32.450 96.170 32.700 ;
        RECT 95.910 32.440 96.320 32.450 ;
        RECT 96.060 32.190 96.320 32.440 ;
        RECT 96.060 30.450 96.320 30.610 ;
        RECT 96.000 30.360 96.500 30.450 ;
        RECT 95.910 30.100 96.500 30.360 ;
        RECT 96.000 29.950 96.500 30.100 ;
        RECT 95.910 29.680 96.170 29.930 ;
        RECT 95.910 29.670 96.320 29.680 ;
        RECT 94.950 24.650 95.450 25.150 ;
        RECT 79.220 23.140 79.480 23.640 ;
        RECT 78.680 22.240 78.940 22.740 ;
        RECT 78.210 21.340 78.470 21.840 ;
        RECT 73.610 19.780 73.870 20.040 ;
        RECT 74.710 19.780 74.970 20.040 ;
        RECT 75.800 19.780 76.060 20.040 ;
        RECT 68.420 19.070 68.680 19.330 ;
        RECT 69.520 19.070 69.780 19.330 ;
        RECT 77.730 20.440 77.990 20.940 ;
        RECT 70.620 19.070 70.880 19.330 ;
        RECT 74.160 19.050 74.420 19.310 ;
        RECT 75.260 19.050 75.520 19.310 ;
        RECT 76.360 19.050 76.620 19.310 ;
        RECT 68.420 17.700 68.680 17.960 ;
        RECT 69.520 17.700 69.780 17.960 ;
        RECT 70.620 17.700 70.880 17.960 ;
        RECT 67.870 17.030 68.130 17.290 ;
        RECT 68.970 17.020 69.230 17.280 ;
        RECT 70.060 17.020 70.320 17.280 ;
        RECT 74.160 17.680 74.420 17.940 ;
        RECT 75.260 17.680 75.520 17.940 ;
        RECT 76.360 17.680 76.620 17.940 ;
        RECT 71.190 17.060 71.450 17.320 ;
        RECT 73.610 17.010 73.870 17.270 ;
        RECT 74.710 17.000 74.970 17.260 ;
        RECT 75.800 17.000 76.060 17.260 ;
        RECT 70.590 16.270 71.050 16.730 ;
        RECT 71.180 16.590 71.440 16.850 ;
        RECT 44.520 14.040 44.780 15.160 ;
        RECT 76.930 17.040 77.190 17.300 ;
        RECT 76.920 16.570 77.180 16.830 ;
        RECT 96.060 29.420 96.320 29.670 ;
        RECT 97.510 29.890 97.780 30.160 ;
        RECT 101.190 27.170 101.690 27.670 ;
        RECT 98.320 19.060 98.820 19.560 ;
        RECT 97.130 18.110 97.630 18.570 ;
        RECT 96.000 17.240 96.500 17.700 ;
        RECT 95.070 16.330 95.570 16.790 ;
        RECT 100.610 14.040 101.550 15.160 ;
        RECT 76.400 10.410 76.730 10.740 ;
        RECT 42.840 9.750 43.170 10.080 ;
        RECT 105.500 50.020 105.890 50.410 ;
        RECT 106.330 49.460 106.710 49.720 ;
        RECT 42.220 9.130 42.550 9.460 ;
        RECT 41.590 8.500 41.920 8.830 ;
        RECT 40.990 7.870 41.320 8.200 ;
        RECT 103.660 9.220 104.060 9.620 ;
        RECT 103.270 8.380 103.530 8.640 ;
        RECT 104.570 8.420 104.960 8.810 ;
        RECT 40.350 7.190 40.680 7.520 ;
        RECT 39.750 6.570 40.080 6.900 ;
        RECT 105.500 7.600 105.890 7.990 ;
        RECT 107.090 47.900 107.350 48.160 ;
        RECT 107.090 47.350 107.350 47.610 ;
        RECT 107.090 45.240 107.350 45.500 ;
        RECT 107.090 44.660 107.350 44.950 ;
        RECT 107.090 44.110 107.350 44.370 ;
        RECT 107.090 42.010 107.350 42.270 ;
        RECT 107.090 41.460 107.350 41.720 ;
        RECT 108.840 55.220 109.100 55.480 ;
        RECT 118.380 65.000 119.090 65.710 ;
        RECT 125.430 67.390 125.690 67.650 ;
        RECT 123.160 64.400 123.420 64.660 ;
        RECT 126.320 66.230 126.580 66.490 ;
        RECT 129.900 68.620 130.160 68.880 ;
        RECT 127.260 65.950 127.520 66.210 ;
        RECT 126.320 65.630 126.580 65.890 ;
        RECT 125.430 64.630 125.690 64.890 ;
        RECT 127.970 65.460 128.230 65.720 ;
        RECT 127.920 64.810 128.180 65.070 ;
        RECT 114.850 59.890 115.110 60.150 ;
        RECT 117.080 59.880 117.340 60.140 ;
        RECT 114.540 59.020 114.800 59.280 ;
        RECT 114.910 58.720 115.170 58.980 ;
        RECT 116.210 59.020 116.470 59.280 ;
        RECT 114.140 58.140 114.400 58.400 ;
        RECT 117.100 58.340 117.360 58.600 ;
        RECT 114.850 56.690 115.110 56.950 ;
        RECT 117.080 56.680 117.340 56.940 ;
        RECT 114.540 55.820 114.800 56.080 ;
        RECT 114.140 54.830 114.400 55.200 ;
        RECT 116.210 55.820 116.470 56.080 ;
        RECT 114.540 53.950 114.800 54.210 ;
        RECT 108.840 52.700 109.100 52.960 ;
        RECT 114.850 53.080 115.110 53.340 ;
        RECT 116.210 53.950 116.470 54.210 ;
        RECT 117.380 53.970 117.640 54.230 ;
        RECT 117.080 53.090 117.340 53.350 ;
        RECT 117.530 53.140 117.790 53.400 ;
        RECT 116.700 52.310 116.960 52.570 ;
        RECT 114.140 51.630 114.400 51.890 ;
        RECT 117.820 51.880 118.080 52.140 ;
        RECT 114.540 50.750 114.800 51.010 ;
        RECT 116.210 50.750 116.470 51.010 ;
        RECT 117.430 51.030 117.690 51.290 ;
        RECT 114.850 49.880 115.110 50.140 ;
        RECT 117.080 49.890 117.340 50.150 ;
        RECT 123.860 62.590 124.120 62.850 ;
        RECT 127.920 63.540 128.180 63.800 ;
        RECT 127.970 62.890 128.230 63.150 ;
        RECT 127.970 62.460 128.230 62.720 ;
        RECT 119.390 61.360 119.650 61.620 ;
        RECT 120.280 60.200 120.540 60.460 ;
        RECT 127.920 61.810 128.180 62.070 ;
        RECT 127.920 60.540 128.180 60.800 ;
        RECT 123.420 60.000 123.680 60.260 ;
        RECT 127.970 59.890 128.230 60.150 ;
        RECT 129.630 65.420 129.890 65.680 ;
        RECT 129.680 63.310 129.940 63.460 ;
        RECT 129.680 63.200 130.160 63.310 ;
        RECT 129.900 63.050 130.160 63.200 ;
        RECT 129.670 62.480 129.930 62.740 ;
        RECT 129.590 60.230 129.850 60.490 ;
        RECT 120.280 59.600 120.540 59.860 ;
        RECT 123.590 59.430 123.850 59.650 ;
        RECT 123.570 59.390 123.850 59.430 ;
        RECT 123.570 59.170 123.830 59.390 ;
        RECT 119.390 58.600 119.650 58.860 ;
        RECT 125.300 58.870 125.560 59.130 ;
        RECT 122.740 58.340 123.000 58.600 ;
        RECT 123.860 57.910 124.120 58.170 ;
        RECT 123.640 57.320 123.900 57.430 ;
        RECT 123.470 57.280 123.900 57.320 ;
        RECT 123.470 57.170 124.120 57.280 ;
        RECT 123.470 57.060 123.730 57.170 ;
        RECT 123.860 57.020 124.120 57.170 ;
        RECT 123.630 56.450 123.890 56.710 ;
        RECT 123.550 54.200 123.810 54.460 ;
        RECT 119.280 52.830 119.550 53.090 ;
        RECT 118.190 45.210 118.900 45.920 ;
        RECT 113.990 27.160 114.500 27.670 ;
        RECT 108.100 13.670 108.360 13.930 ;
        RECT 108.100 13.000 108.360 13.260 ;
        RECT 108.370 11.710 108.630 11.970 ;
        RECT 108.370 10.100 108.630 10.360 ;
        RECT 108.360 8.490 108.620 8.750 ;
        RECT 106.320 6.810 106.700 7.190 ;
        RECT 108.370 6.870 108.630 7.130 ;
        RECT 39.150 5.930 39.480 6.260 ;
        RECT 38.570 5.360 38.900 5.690 ;
        RECT 37.990 4.670 38.320 5.000 ;
        RECT 108.360 5.260 108.620 5.520 ;
        RECT 37.340 4.030 37.670 4.360 ;
        RECT 36.700 3.380 37.030 3.720 ;
        RECT 107.600 3.780 107.860 4.040 ;
        RECT 36.120 2.740 36.490 3.110 ;
        RECT 108.360 2.060 108.620 2.320 ;
        RECT 105.120 0.350 105.380 0.610 ;
        RECT 106.060 0.350 106.320 0.610 ;
        RECT 107.010 0.330 107.270 0.590 ;
        RECT 108.320 0.350 108.580 0.610 ;
      LAYER met2 ;
        RECT 26.030 70.480 26.780 70.490 ;
        RECT 26.030 70.180 27.650 70.480 ;
        RECT 26.030 70.010 26.270 70.180 ;
        RECT 27.350 69.960 27.650 70.180 ;
        RECT 0.970 69.050 1.290 69.310 ;
        RECT 3.830 69.210 4.150 69.360 ;
        RECT 1.350 68.970 4.240 69.210 ;
        RECT 87.830 68.910 88.140 68.920 ;
        RECT 85.660 68.730 88.140 68.910 ;
        RECT 87.830 68.590 88.140 68.730 ;
        RECT 129.870 68.910 130.180 68.920 ;
        RECT 129.870 68.730 132.350 68.910 ;
        RECT 129.870 68.590 130.180 68.730 ;
        RECT 90.420 68.310 90.500 68.490 ;
        RECT 18.390 67.670 18.700 67.680 ;
        RECT 3.630 66.390 3.900 67.670 ;
        RECT 18.390 67.350 18.810 67.670 ;
        RECT 18.510 67.210 18.810 67.350 ;
        RECT 19.080 67.660 19.390 67.670 ;
        RECT 19.080 67.340 19.540 67.660 ;
        RECT 125.400 67.470 125.710 67.690 ;
        RECT 125.400 67.360 127.590 67.470 ;
        RECT 19.240 67.200 19.540 67.340 ;
        RECT 125.560 67.250 127.590 67.360 ;
        RECT 92.060 66.950 92.370 67.120 ;
        RECT 92.060 66.790 101.940 66.950 ;
        RECT 92.230 66.760 101.940 66.790 ;
        RECT 1.110 66.380 3.900 66.390 ;
        RECT 0.450 66.160 3.900 66.380 ;
        RECT 126.290 66.230 126.610 66.490 ;
        RECT 0.450 66.150 3.380 66.160 ;
        RECT 0.960 65.990 1.280 66.060 ;
        RECT 0.450 65.800 1.280 65.990 ;
        RECT 91.390 65.940 91.710 66.200 ;
        RECT 127.230 66.130 127.550 66.210 ;
        RECT 91.780 66.030 101.940 66.070 ;
        RECT 91.770 65.840 101.940 66.030 ;
        RECT 126.240 65.950 127.550 66.130 ;
        RECT 0.450 65.670 1.070 65.800 ;
        RECT 126.240 65.780 127.420 65.950 ;
        RECT 126.290 65.630 126.610 65.780 ;
        RECT 3.330 65.510 3.640 65.590 ;
        RECT 0.450 65.280 3.640 65.510 ;
        RECT 127.940 65.470 128.250 65.760 ;
        RECT 129.600 65.470 129.910 65.720 ;
        RECT 3.330 65.260 3.640 65.280 ;
        RECT 127.220 65.390 129.910 65.470 ;
        RECT 127.220 65.240 129.760 65.390 ;
        RECT 92.220 64.900 101.940 65.090 ;
        RECT 1.620 64.370 1.930 64.700 ;
        RECT 3.050 64.390 3.360 64.720 ;
        RECT 125.400 64.710 125.710 64.930 ;
        RECT 127.450 64.710 127.780 64.880 ;
        RECT 127.890 64.780 128.200 65.110 ;
        RECT 125.400 64.670 127.780 64.710 ;
        RECT 124.230 64.430 124.540 64.670 ;
        RECT 125.400 64.600 127.590 64.670 ;
        RECT 125.550 64.500 127.590 64.600 ;
        RECT 125.340 63.800 125.560 63.820 ;
        RECT 90.420 63.440 90.500 63.620 ;
        RECT 92.730 63.610 92.890 63.630 ;
        RECT 92.730 63.560 101.940 63.610 ;
        RECT 92.850 63.460 101.940 63.560 ;
        RECT 125.290 63.460 125.560 63.800 ;
        RECT 127.450 63.730 127.780 63.940 ;
        RECT 127.890 63.500 128.200 63.830 ;
        RECT 129.650 63.340 129.960 63.500 ;
        RECT 129.650 63.330 130.180 63.340 ;
        RECT 127.480 63.200 130.180 63.330 ;
        RECT 123.550 62.960 123.900 63.180 ;
        RECT 127.480 63.100 132.350 63.200 ;
        RECT 125.360 62.890 125.560 62.900 ;
        RECT 123.830 62.880 124.140 62.890 ;
        RECT 125.360 62.880 125.580 62.890 ;
        RECT 123.830 62.700 126.310 62.880 ;
        RECT 127.940 62.850 128.250 63.100 ;
        RECT 129.870 63.020 132.350 63.100 ;
        RECT 129.870 63.010 130.180 63.020 ;
        RECT 123.830 62.560 124.140 62.700 ;
        RECT 125.360 62.560 125.580 62.700 ;
        RECT 125.380 62.550 125.580 62.560 ;
        RECT 127.940 62.500 128.250 62.760 ;
        RECT 129.640 62.500 129.950 62.780 ;
        RECT 110.020 62.280 119.140 62.460 ;
        RECT 127.220 62.280 130.130 62.500 ;
        RECT 99.810 61.870 100.120 62.070 ;
        RECT 99.810 61.860 100.410 61.870 ;
        RECT 99.810 61.740 102.200 61.860 ;
        RECT 124.310 61.760 124.630 62.000 ;
        RECT 99.950 61.700 102.200 61.740 ;
        RECT 100.260 61.680 102.200 61.700 ;
        RECT 127.450 61.670 127.780 61.880 ;
        RECT 127.890 61.780 128.200 62.110 ;
        RECT 128.650 61.990 128.760 62.220 ;
        RECT 128.650 61.170 128.760 61.390 ;
        RECT 43.680 60.500 43.780 60.820 ;
        RECT 127.450 60.730 127.780 60.940 ;
        RECT 52.600 60.370 55.450 60.570 ;
        RECT 127.890 60.500 128.200 60.830 ;
        RECT 52.210 59.680 52.380 59.880 ;
        RECT 55.250 59.870 55.450 60.370 ;
        RECT 129.560 60.340 129.870 60.530 ;
        RECT 127.210 60.110 129.920 60.340 ;
        RECT 81.270 59.870 81.580 59.930 ;
        RECT 55.250 59.670 81.580 59.870 ;
        RECT 127.940 59.850 128.250 60.110 ;
        RECT 81.270 59.610 81.580 59.670 ;
        RECT 60.200 59.400 60.520 59.450 ;
        RECT 55.200 59.200 60.570 59.400 ;
        RECT 55.200 58.820 55.400 59.200 ;
        RECT 60.200 59.190 60.520 59.200 ;
        RECT 100.660 59.150 100.740 59.330 ;
        RECT 62.960 58.960 63.270 58.970 ;
        RECT 62.960 58.930 63.280 58.960 ;
        RECT 20.680 58.610 20.750 58.650 ;
        RECT 52.600 58.620 55.400 58.820 ;
        RECT 55.710 58.730 63.280 58.930 ;
        RECT 20.680 58.380 20.820 58.610 ;
        RECT 22.660 58.390 23.480 58.560 ;
        RECT 52.190 57.930 52.380 58.130 ;
        RECT 20.680 57.460 20.820 57.630 ;
        RECT 22.660 57.470 23.480 57.640 ;
        RECT 20.960 57.140 21.270 57.470 ;
        RECT 23.620 57.090 23.930 57.330 ;
        RECT 23.620 57.000 23.940 57.090 ;
        RECT 55.710 57.070 55.910 58.730 ;
        RECT 62.960 58.700 63.280 58.730 ;
        RECT 62.960 58.690 63.270 58.700 ;
        RECT 64.020 58.450 64.340 58.490 ;
        RECT 23.720 56.920 23.940 57.000 ;
        RECT 52.600 56.870 55.910 57.070 ;
        RECT 56.260 58.250 64.420 58.450 ;
        RECT 122.710 58.300 123.020 58.630 ;
        RECT 20.680 56.680 20.820 56.710 ;
        RECT 20.680 56.540 20.890 56.680 ;
        RECT 20.940 56.150 21.250 56.480 ;
        RECT 21.960 56.140 22.330 56.330 ;
        RECT 23.740 56.160 24.050 56.490 ;
        RECT 52.220 56.180 52.380 56.380 ;
        RECT 20.680 55.520 20.820 55.710 ;
        RECT 23.740 55.170 24.050 55.500 ;
        RECT 43.680 55.250 43.780 55.570 ;
        RECT 56.260 55.320 56.460 58.250 ;
        RECT 64.020 58.210 64.340 58.250 ;
        RECT 94.630 57.990 94.700 58.170 ;
        RECT 118.420 58.010 118.490 58.210 ;
        RECT 115.790 56.880 115.860 57.080 ;
        RECT 117.510 56.930 117.860 57.150 ;
        RECT 52.560 55.120 56.460 55.320 ;
        RECT 59.410 56.450 59.700 56.630 ;
        RECT 20.680 54.730 20.820 54.750 ;
        RECT 20.680 54.560 20.750 54.730 ;
        RECT 23.740 54.180 24.050 54.510 ;
        RECT 20.680 53.740 20.820 53.790 ;
        RECT 20.680 53.600 20.750 53.740 ;
        RECT 59.410 53.610 59.590 56.450 ;
        RECT 115.650 55.840 115.870 55.850 ;
        RECT 116.180 55.840 116.490 56.120 ;
        RECT 115.650 55.640 117.280 55.840 ;
        RECT 118.270 55.730 118.590 55.970 ;
        RECT 122.610 55.960 122.720 56.190 ;
        RECT 115.650 55.630 115.870 55.640 ;
        RECT 103.110 55.510 103.430 55.560 ;
        RECT 103.110 55.260 109.130 55.510 ;
        RECT 108.810 55.190 109.130 55.260 ;
        RECT 111.100 55.170 111.150 55.370 ;
        RECT 118.420 55.020 118.490 55.220 ;
        RECT 122.610 55.140 122.720 55.360 ;
        RECT 111.100 54.660 111.150 54.860 ;
        RECT 118.420 54.810 118.490 55.010 ;
        RECT 83.760 54.020 84.360 54.580 ;
        RECT 87.360 54.410 92.590 54.640 ;
        RECT 115.650 54.390 115.870 54.400 ;
        RECT 115.650 54.190 117.280 54.390 ;
        RECT 115.650 54.180 115.870 54.190 ;
        RECT 116.180 53.910 116.490 54.190 ;
        RECT 103.480 53.870 103.960 53.880 ;
        RECT 58.640 53.440 59.590 53.610 ;
        RECT 67.530 53.430 69.310 53.600 ;
        RECT 87.370 53.590 92.590 53.810 ;
        RECT 92.960 53.590 101.170 53.810 ;
        RECT 103.480 53.630 104.370 53.870 ;
        RECT 62.510 53.150 62.830 53.200 ;
        RECT 64.920 53.150 65.240 53.170 ;
        RECT 52.980 53.010 53.180 53.130 ;
        RECT 52.980 52.810 53.330 53.010 ;
        RECT 62.510 52.960 65.240 53.150 ;
        RECT 94.630 53.120 94.710 53.300 ;
        RECT 62.510 52.880 62.830 52.960 ;
        RECT 63.590 52.890 63.680 52.960 ;
        RECT 64.920 52.910 65.240 52.960 ;
        RECT 52.980 52.790 53.180 52.810 ;
        RECT 43.680 52.340 43.780 52.660 ;
        RECT 52.600 52.590 53.180 52.790 ;
        RECT 61.310 52.440 61.750 52.670 ;
        RECT 61.410 52.370 61.750 52.440 ;
        RECT 61.410 52.230 61.750 52.300 ;
        RECT 61.310 52.000 61.750 52.230 ;
        RECT 46.430 51.410 46.890 51.730 ;
        RECT 48.600 51.370 51.040 51.590 ;
        RECT 52.220 51.530 52.380 51.730 ;
        RECT 52.930 51.590 53.300 51.790 ;
        RECT 43.680 50.590 43.780 50.910 ;
        RECT 48.700 50.570 48.960 51.370 ;
        RECT 49.620 51.340 49.940 51.360 ;
        RECT 49.610 51.290 49.940 51.340 ;
        RECT 50.700 51.310 51.040 51.370 ;
        RECT 50.650 51.290 50.970 51.300 ;
        RECT 49.610 51.090 52.280 51.290 ;
        RECT 49.610 51.080 49.940 51.090 ;
        RECT 49.620 51.070 49.940 51.080 ;
        RECT 50.650 51.040 50.970 51.090 ;
        RECT 52.930 51.040 53.130 51.590 ;
        RECT 58.970 51.560 59.700 51.740 ;
        RECT 62.510 51.710 62.830 51.790 ;
        RECT 63.590 51.710 63.670 51.780 ;
        RECT 64.920 51.710 65.240 51.760 ;
        RECT 58.970 51.350 59.150 51.560 ;
        RECT 62.510 51.520 65.240 51.710 ;
        RECT 62.510 51.470 62.830 51.520 ;
        RECT 64.920 51.500 65.240 51.520 ;
        RECT 100.950 51.710 101.170 53.590 ;
        RECT 117.510 53.250 117.820 53.440 ;
        RECT 117.470 53.000 118.020 53.250 ;
        RECT 111.100 51.970 111.150 52.170 ;
        RECT 113.730 51.890 114.340 52.020 ;
        RECT 117.650 51.970 118.120 52.220 ;
        RECT 113.730 51.820 114.430 51.890 ;
        RECT 117.790 51.880 118.110 51.970 ;
        RECT 118.420 51.820 118.490 52.020 ;
        RECT 100.950 51.700 102.550 51.710 ;
        RECT 100.950 51.500 110.940 51.700 ;
        RECT 114.110 51.630 114.430 51.820 ;
        RECT 100.950 51.490 102.550 51.500 ;
        RECT 58.580 51.170 59.150 51.350 ;
        RECT 67.310 51.180 69.310 51.340 ;
        RECT 68.040 51.170 69.310 51.180 ;
        RECT 68.740 51.160 69.310 51.170 ;
        RECT 88.140 51.130 92.590 51.290 ;
        RECT 88.110 51.090 92.590 51.130 ;
        RECT 92.960 51.190 110.150 51.290 ;
        RECT 92.960 51.090 110.940 51.190 ;
        RECT 52.600 50.840 53.130 51.040 ;
        RECT 59.070 50.410 59.620 50.590 ;
        RECT 82.700 50.550 83.260 51.090 ;
        RECT 59.070 50.390 59.250 50.410 ;
        RECT 58.650 50.230 59.250 50.390 ;
        RECT 67.530 50.220 69.310 50.380 ;
        RECT 46.430 49.660 46.890 49.980 ;
        RECT 48.600 49.620 51.040 49.840 ;
        RECT 52.190 49.780 52.380 49.980 ;
        RECT 62.510 49.950 62.830 50.000 ;
        RECT 64.920 49.950 65.240 49.970 ;
        RECT 48.700 48.820 48.960 49.620 ;
        RECT 49.620 49.590 49.940 49.610 ;
        RECT 49.610 49.540 49.940 49.590 ;
        RECT 50.700 49.560 51.040 49.620 ;
        RECT 50.650 49.540 50.970 49.550 ;
        RECT 49.610 49.340 52.280 49.540 ;
        RECT 52.960 49.480 53.280 49.920 ;
        RECT 62.510 49.760 65.240 49.950 ;
        RECT 62.510 49.680 62.830 49.760 ;
        RECT 63.590 49.680 63.740 49.760 ;
        RECT 64.920 49.710 65.240 49.760 ;
        RECT 49.610 49.330 49.940 49.340 ;
        RECT 49.620 49.320 49.940 49.330 ;
        RECT 50.650 49.290 50.970 49.340 ;
        RECT 52.960 49.290 53.160 49.480 ;
        RECT 52.600 49.090 53.160 49.290 ;
        RECT 61.310 49.240 61.750 49.470 ;
        RECT 61.410 49.170 61.750 49.240 ;
        RECT 61.410 49.030 61.750 49.100 ;
        RECT 61.310 48.800 61.750 49.030 ;
        RECT 88.110 48.610 88.340 51.090 ;
        RECT 109.850 50.990 110.940 51.090 ;
        RECT 114.040 51.040 114.610 51.190 ;
        RECT 114.040 50.990 114.820 51.040 ;
        RECT 114.510 50.710 114.820 50.990 ;
        RECT 52.890 48.360 53.270 48.540 ;
        RECT 62.510 48.510 62.830 48.590 ;
        RECT 63.590 48.510 63.670 48.580 ;
        RECT 64.920 48.510 65.240 48.560 ;
        RECT 46.430 47.910 46.890 48.230 ;
        RECT 48.600 47.870 51.040 48.090 ;
        RECT 52.210 48.030 52.380 48.230 ;
        RECT 43.680 47.090 43.780 47.410 ;
        RECT 48.700 47.070 48.960 47.870 ;
        RECT 49.620 47.840 49.940 47.860 ;
        RECT 49.610 47.790 49.940 47.840 ;
        RECT 50.700 47.810 51.040 47.870 ;
        RECT 50.650 47.790 50.970 47.800 ;
        RECT 49.610 47.590 52.280 47.790 ;
        RECT 49.610 47.580 49.940 47.590 ;
        RECT 49.620 47.570 49.940 47.580 ;
        RECT 50.650 47.540 50.970 47.590 ;
        RECT 52.890 47.540 53.070 48.360 ;
        RECT 62.510 48.320 65.240 48.510 ;
        RECT 62.510 48.270 62.830 48.320 ;
        RECT 64.920 48.300 65.240 48.320 ;
        RECT 58.630 47.910 59.350 48.090 ;
        RECT 52.600 47.340 53.080 47.540 ;
        RECT 46.430 46.160 46.890 46.480 ;
        RECT 48.600 46.120 51.040 46.340 ;
        RECT 52.220 46.280 52.380 46.480 ;
        RECT 48.700 45.320 48.960 46.120 ;
        RECT 49.620 46.090 49.940 46.110 ;
        RECT 49.610 46.040 49.940 46.090 ;
        RECT 50.700 46.060 51.040 46.120 ;
        RECT 50.650 46.040 50.970 46.050 ;
        RECT 49.610 45.840 52.280 46.040 ;
        RECT 49.610 45.830 49.940 45.840 ;
        RECT 49.620 45.820 49.940 45.830 ;
        RECT 50.650 45.790 50.970 45.840 ;
        RECT 59.170 45.720 59.350 47.910 ;
        RECT 67.530 47.900 69.310 48.080 ;
        RECT 80.250 47.910 80.560 48.200 ;
        RECT 83.740 48.000 84.360 48.530 ;
        RECT 87.360 48.380 88.340 48.610 ;
        RECT 88.950 48.480 92.590 48.680 ;
        RECT 92.960 48.500 110.150 48.680 ;
        RECT 92.960 48.480 110.940 48.500 ;
        RECT 78.230 47.870 80.560 47.910 ;
        RECT 78.230 47.730 80.410 47.870 ;
        RECT 88.950 47.780 89.150 48.480 ;
        RECT 109.890 48.300 110.940 48.480 ;
        RECT 107.060 47.910 107.370 48.200 ;
        RECT 107.060 47.870 109.390 47.910 ;
        RECT 80.250 47.480 80.560 47.650 ;
        RECT 87.370 47.630 89.150 47.780 ;
        RECT 107.210 47.730 109.390 47.870 ;
        RECT 87.370 47.560 89.120 47.630 ;
        RECT 78.230 47.320 80.560 47.480 ;
        RECT 78.230 47.300 80.400 47.320 ;
        RECT 80.700 47.300 80.790 47.480 ;
        RECT 83.560 47.320 91.190 47.500 ;
        RECT 96.430 47.320 104.060 47.500 ;
        RECT 107.060 47.480 107.370 47.650 ;
        RECT 106.830 47.300 106.920 47.480 ;
        RECT 107.060 47.320 109.390 47.480 ;
        RECT 107.220 47.300 109.390 47.320 ;
        RECT 83.560 46.880 91.190 47.060 ;
        RECT 96.430 46.880 104.060 47.060 ;
        RECT 83.560 45.780 91.190 45.960 ;
        RECT 96.430 45.780 104.060 45.960 ;
        RECT 59.170 45.540 59.710 45.720 ;
        RECT 78.230 45.530 80.400 45.550 ;
        RECT 78.230 45.370 80.560 45.530 ;
        RECT 80.700 45.370 80.790 45.550 ;
        RECT 80.250 45.200 80.560 45.370 ;
        RECT 83.560 45.350 91.190 45.530 ;
        RECT 96.430 45.350 104.060 45.530 ;
        RECT 106.830 45.370 106.920 45.550 ;
        RECT 107.220 45.530 109.390 45.550 ;
        RECT 107.060 45.370 109.390 45.530 ;
        RECT 107.060 45.200 107.370 45.370 ;
        RECT 107.210 44.980 109.390 45.120 ;
        RECT 107.060 44.940 109.390 44.980 ;
        RECT 107.060 44.670 107.370 44.940 ;
        RECT 107.060 44.630 109.390 44.670 ;
        RECT 107.210 44.490 109.390 44.630 ;
        RECT 96.430 44.080 104.050 44.260 ;
        RECT 107.060 44.240 107.370 44.410 ;
        RECT 106.830 44.060 106.920 44.240 ;
        RECT 107.060 44.080 109.390 44.240 ;
        RECT 107.220 44.060 109.390 44.080 ;
        RECT 83.560 43.650 91.190 43.830 ;
        RECT 96.430 43.650 104.060 43.830 ;
        RECT 59.090 43.120 59.270 43.130 ;
        RECT 58.750 43.010 59.270 43.120 ;
        RECT 58.750 42.940 61.100 43.010 ;
        RECT 67.510 42.960 69.290 43.130 ;
        RECT 59.090 42.830 61.100 42.940 ;
        RECT 83.750 42.870 83.810 43.050 ;
        RECT 103.780 42.870 103.870 43.050 ;
        RECT 62.490 42.680 62.810 42.730 ;
        RECT 64.900 42.680 65.220 42.700 ;
        RECT 43.680 42.210 43.780 42.530 ;
        RECT 52.670 42.460 53.270 42.660 ;
        RECT 62.490 42.490 65.220 42.680 ;
        RECT 83.570 42.550 91.190 42.730 ;
        RECT 96.430 42.550 104.050 42.730 ;
        RECT 62.490 42.410 62.810 42.490 ;
        RECT 63.570 42.420 63.660 42.490 ;
        RECT 64.900 42.440 65.220 42.490 ;
        RECT 83.750 42.440 83.820 42.550 ;
        RECT 103.780 42.440 103.870 42.550 ;
        RECT 78.230 42.300 80.400 42.320 ;
        RECT 61.290 41.970 61.730 42.200 ;
        RECT 78.230 42.140 80.560 42.300 ;
        RECT 80.700 42.140 80.790 42.320 ;
        RECT 80.250 41.970 80.560 42.140 ;
        RECT 83.590 42.130 91.190 42.300 ;
        RECT 96.430 42.130 104.030 42.300 ;
        RECT 106.830 42.140 106.920 42.320 ;
        RECT 107.220 42.300 109.390 42.320 ;
        RECT 107.060 42.140 109.390 42.300 ;
        RECT 107.060 41.970 107.370 42.140 ;
        RECT 61.390 41.900 61.730 41.970 ;
        RECT 61.390 41.760 61.730 41.830 ;
        RECT 52.220 41.400 52.380 41.600 ;
        RECT 61.290 41.530 61.730 41.760 ;
        RECT 78.230 41.750 80.410 41.890 ;
        RECT 107.210 41.750 109.390 41.890 ;
        RECT 78.230 41.710 80.560 41.750 ;
        RECT 80.250 41.420 80.560 41.710 ;
        RECT 107.060 41.710 109.390 41.750 ;
        RECT 103.810 41.330 103.870 41.510 ;
        RECT 107.060 41.420 107.370 41.710 ;
        RECT 52.870 41.260 53.250 41.270 ;
        RECT 52.850 41.090 53.250 41.260 ;
        RECT 62.490 41.240 62.810 41.320 ;
        RECT 63.570 41.240 63.650 41.310 ;
        RECT 64.900 41.240 65.220 41.290 ;
        RECT 52.850 40.910 53.050 41.090 ;
        RECT 62.490 41.050 65.220 41.240 ;
        RECT 43.680 40.460 43.780 40.780 ;
        RECT 52.600 40.710 53.050 40.910 ;
        RECT 58.830 40.880 61.160 41.040 ;
        RECT 62.490 41.000 62.810 41.050 ;
        RECT 64.900 41.030 65.220 41.050 ;
        RECT 83.750 40.900 83.880 41.080 ;
        RECT 103.810 40.900 103.870 41.080 ;
        RECT 58.610 40.860 61.160 40.880 ;
        RECT 58.610 40.700 59.010 40.860 ;
        RECT 67.290 40.710 69.290 40.870 ;
        RECT 68.020 40.700 69.290 40.710 ;
        RECT 68.720 40.690 69.290 40.700 ;
        RECT 58.630 39.910 59.030 39.920 ;
        RECT 52.190 39.650 52.380 39.850 ;
        RECT 58.630 39.770 59.040 39.910 ;
        RECT 58.630 39.760 61.140 39.770 ;
        RECT 58.860 39.590 61.140 39.760 ;
        RECT 67.510 39.750 69.290 39.910 ;
        RECT 83.750 39.630 83.820 39.810 ;
        RECT 103.780 39.630 103.870 39.810 ;
        RECT 62.490 39.480 62.810 39.530 ;
        RECT 64.900 39.480 65.220 39.500 ;
        RECT 52.800 39.310 53.250 39.440 ;
        RECT 52.800 39.160 53.290 39.310 ;
        RECT 62.490 39.290 65.220 39.480 ;
        RECT 62.490 39.210 62.810 39.290 ;
        RECT 63.570 39.210 63.720 39.290 ;
        RECT 64.900 39.240 65.220 39.290 ;
        RECT 52.600 39.110 53.290 39.160 ;
        RECT 52.600 38.960 53.150 39.110 ;
        RECT 80.850 39.070 81.160 39.360 ;
        RECT 83.750 39.200 83.820 39.380 ;
        RECT 103.780 39.200 103.870 39.380 ;
        RECT 78.830 39.030 81.160 39.070 ;
        RECT 61.290 38.770 61.730 39.000 ;
        RECT 78.830 38.890 81.010 39.030 ;
        RECT 61.390 38.700 61.730 38.770 ;
        RECT 80.850 38.640 81.160 38.810 ;
        RECT 90.450 38.710 97.210 38.890 ;
        RECT 61.390 38.560 61.730 38.630 ;
        RECT 61.290 38.330 61.730 38.560 ;
        RECT 78.830 38.480 81.160 38.640 ;
        RECT 78.830 38.460 81.000 38.480 ;
        RECT 81.300 38.460 81.390 38.640 ;
        RECT 81.720 38.480 81.810 38.660 ;
        RECT 52.210 37.900 52.380 38.100 ;
        RECT 52.840 37.890 53.270 38.120 ;
        RECT 62.490 38.040 62.810 38.120 ;
        RECT 63.570 38.040 63.650 38.110 ;
        RECT 64.900 38.040 65.220 38.090 ;
        RECT 81.720 38.050 81.810 38.230 ;
        RECT 83.750 38.100 83.820 38.280 ;
        RECT 84.180 38.040 91.790 38.230 ;
        RECT 103.780 38.100 103.870 38.280 ;
        RECT 52.840 37.410 53.040 37.890 ;
        RECT 62.490 37.850 65.220 38.040 ;
        RECT 58.820 37.630 61.120 37.810 ;
        RECT 62.490 37.800 62.810 37.850 ;
        RECT 64.900 37.830 65.220 37.850 ;
        RECT 83.750 37.670 83.820 37.850 ;
        RECT 103.780 37.670 103.870 37.850 ;
        RECT 58.820 37.620 59.020 37.630 ;
        RECT 58.610 37.440 59.020 37.620 ;
        RECT 67.510 37.430 69.290 37.610 ;
        RECT 43.680 36.960 43.780 37.280 ;
        RECT 52.600 37.210 53.040 37.410 ;
        RECT 81.720 36.960 81.810 37.140 ;
        RECT 84.160 36.960 91.790 37.140 ;
        RECT 52.220 36.150 52.380 36.350 ;
        RECT 81.720 34.810 81.830 34.990 ;
        RECT 84.160 34.820 91.020 34.990 ;
        RECT 91.320 34.850 91.790 35.010 ;
        RECT 91.320 34.840 91.780 34.850 ;
        RECT 84.910 34.420 85.230 34.480 ;
        RECT 88.930 34.420 89.260 34.450 ;
        RECT 84.910 34.250 89.260 34.420 ;
        RECT 83.810 34.070 84.540 34.250 ;
        RECT 84.910 34.200 85.230 34.250 ;
        RECT 87.210 34.230 87.530 34.250 ;
        RECT 88.930 34.230 89.260 34.250 ;
        RECT 87.210 34.090 95.040 34.230 ;
        RECT 87.390 34.040 95.040 34.090 ;
        RECT 87.390 34.030 95.210 34.040 ;
        RECT 84.160 34.020 95.210 34.030 ;
        RECT 58.640 33.680 58.950 33.860 ;
        RECT 67.540 33.690 69.320 33.860 ;
        RECT 81.720 33.710 81.830 33.890 ;
        RECT 84.160 33.860 91.790 34.020 ;
        RECT 94.830 33.830 95.210 34.020 ;
        RECT 94.320 33.820 94.460 33.830 ;
        RECT 26.930 32.980 27.240 33.310 ;
        RECT 43.640 33.150 43.740 33.470 ;
        RECT 52.560 33.400 53.170 33.600 ;
        RECT 58.770 33.500 61.120 33.680 ;
        RECT 78.830 33.460 81.000 33.480 ;
        RECT 52.970 33.360 53.170 33.400 ;
        RECT 62.520 33.410 62.840 33.460 ;
        RECT 64.930 33.410 65.250 33.430 ;
        RECT 52.970 33.160 53.390 33.360 ;
        RECT 62.520 33.220 65.250 33.410 ;
        RECT 78.830 33.300 81.160 33.460 ;
        RECT 81.300 33.300 81.390 33.480 ;
        RECT 62.520 33.140 62.840 33.220 ;
        RECT 63.600 33.150 63.690 33.220 ;
        RECT 64.930 33.170 65.250 33.220 ;
        RECT 80.850 33.130 81.160 33.300 ;
        RECT 81.720 33.280 81.830 33.460 ;
        RECT 83.850 33.190 84.000 33.610 ;
        RECT 94.320 33.490 94.470 33.820 ;
        RECT 83.850 33.100 87.120 33.190 ;
        RECT 87.190 33.100 87.510 33.300 ;
        RECT 94.320 33.290 95.530 33.490 ;
        RECT 24.900 32.760 25.610 32.970 ;
        RECT 59.410 32.870 60.580 33.020 ;
        RECT 59.350 32.540 59.630 32.870 ;
        RECT 61.320 32.700 61.760 32.930 ;
        RECT 78.830 32.910 81.010 33.050 ;
        RECT 83.850 33.040 87.510 33.100 ;
        RECT 95.640 33.060 95.760 33.270 ;
        RECT 96.670 33.180 97.930 33.340 ;
        RECT 86.980 32.940 87.280 33.040 ;
        RECT 78.830 32.870 81.160 32.910 ;
        RECT 61.420 32.630 61.760 32.700 ;
        RECT 80.850 32.580 81.160 32.870 ;
        RECT 83.920 32.710 84.240 32.800 ;
        RECT 52.180 32.340 52.340 32.540 ;
        RECT 61.420 32.490 61.760 32.560 ;
        RECT 27.950 32.230 28.270 32.290 ;
        RECT 61.320 32.260 61.760 32.490 ;
        RECT 83.830 32.540 84.240 32.710 ;
        RECT 94.430 32.630 95.630 32.730 ;
        RECT 94.420 32.550 95.630 32.630 ;
        RECT 83.830 32.440 84.150 32.540 ;
        RECT 95.350 32.430 95.630 32.550 ;
        RECT 95.350 32.410 95.380 32.430 ;
        RECT 95.640 32.300 95.760 32.510 ;
        RECT 27.950 32.020 28.430 32.230 ;
        RECT 83.780 32.120 84.360 32.300 ;
        RECT 27.950 31.970 28.270 32.020 ;
        RECT 52.960 31.850 53.280 32.010 ;
        RECT 24.900 31.400 25.150 31.620 ;
        RECT 43.640 31.400 43.740 31.720 ;
        RECT 52.560 31.650 53.280 31.850 ;
        RECT 62.520 31.970 62.840 32.050 ;
        RECT 63.600 31.970 63.680 32.040 ;
        RECT 64.930 31.970 65.250 32.020 ;
        RECT 62.520 31.780 65.250 31.970 ;
        RECT 87.060 31.960 87.290 31.970 ;
        RECT 87.060 31.930 94.630 31.960 ;
        RECT 62.520 31.730 62.840 31.780 ;
        RECT 64.930 31.760 65.250 31.780 ;
        RECT 58.750 31.600 60.540 31.730 ;
        RECT 83.900 31.660 84.220 31.790 ;
        RECT 87.060 31.760 94.690 31.930 ;
        RECT 87.060 31.660 87.300 31.760 ;
        RECT 58.610 31.550 60.540 31.600 ;
        RECT 58.610 31.400 58.930 31.550 ;
        RECT 67.320 31.440 69.320 31.600 ;
        RECT 83.850 31.480 87.300 31.660 ;
        RECT 94.500 31.560 95.210 31.760 ;
        RECT 83.850 31.460 87.220 31.480 ;
        RECT 68.050 31.430 69.320 31.440 ;
        RECT 68.750 31.420 69.320 31.430 ;
        RECT 58.610 31.320 58.790 31.400 ;
        RECT 87.190 31.280 87.510 31.420 ;
        RECT 87.190 31.260 94.650 31.280 ;
        RECT 87.190 31.160 95.210 31.260 ;
        RECT 87.200 31.060 95.210 31.160 ;
        RECT 87.200 31.050 87.520 31.060 ;
        RECT 83.810 30.830 84.360 31.010 ;
        RECT 52.150 30.590 52.340 30.790 ;
        RECT 58.660 30.490 58.860 30.650 ;
        RECT 58.680 30.440 58.860 30.490 ;
        RECT 67.540 30.480 69.320 30.640 ;
        RECT 58.680 30.260 60.570 30.440 ;
        RECT 62.520 30.210 62.840 30.260 ;
        RECT 64.930 30.210 65.250 30.230 ;
        RECT 52.560 30.080 53.250 30.100 ;
        RECT 27.930 29.620 28.250 29.670 ;
        RECT 43.640 29.650 43.740 29.970 ;
        RECT 52.560 29.900 53.330 30.080 ;
        RECT 53.040 29.810 53.330 29.900 ;
        RECT 59.960 30.030 60.280 30.070 ;
        RECT 59.960 29.820 60.570 30.030 ;
        RECT 62.520 30.020 65.250 30.210 ;
        RECT 62.520 29.940 62.840 30.020 ;
        RECT 63.600 29.940 63.750 30.020 ;
        RECT 64.930 29.970 65.250 30.020 ;
        RECT 83.790 30.100 83.990 30.600 ;
        RECT 94.410 30.440 95.410 30.600 ;
        RECT 95.640 30.290 95.760 30.500 ;
        RECT 87.060 30.100 87.380 30.240 ;
        RECT 83.790 29.980 87.380 30.100 ;
        RECT 83.790 29.900 87.340 29.980 ;
        RECT 59.960 29.750 60.420 29.820 ;
        RECT 27.930 29.410 28.430 29.620 ;
        RECT 61.320 29.500 61.760 29.730 ;
        RECT 83.900 29.660 84.210 29.840 ;
        RECT 61.420 29.430 61.760 29.500 ;
        RECT 83.780 29.510 84.210 29.660 ;
        RECT 27.930 29.350 28.250 29.410 ;
        RECT 83.780 29.390 84.060 29.510 ;
        RECT 94.420 29.460 95.420 29.630 ;
        RECT 95.640 29.530 95.760 29.740 ;
        RECT 94.420 29.450 95.360 29.460 ;
        RECT 61.420 29.290 61.760 29.360 ;
        RECT 24.900 29.080 25.170 29.090 ;
        RECT 24.900 28.870 25.650 29.080 ;
        RECT 61.320 29.060 61.760 29.290 ;
        RECT 52.170 28.840 52.340 29.040 ;
        RECT 53.020 28.930 53.320 28.970 ;
        RECT 53.010 28.690 53.320 28.930 ;
        RECT 83.790 28.870 84.360 29.050 ;
        RECT 94.650 29.000 95.200 29.010 ;
        RECT 62.520 28.770 62.840 28.850 ;
        RECT 63.600 28.770 63.680 28.840 ;
        RECT 64.930 28.770 65.250 28.820 ;
        RECT 22.780 28.520 23.380 28.670 ;
        RECT 22.630 28.190 23.380 28.520 ;
        RECT 53.010 28.350 53.210 28.690 ;
        RECT 62.520 28.580 65.250 28.770 ;
        RECT 83.950 28.720 84.260 28.870 ;
        RECT 62.520 28.530 62.840 28.580 ;
        RECT 64.930 28.560 65.250 28.580 ;
        RECT 83.830 28.590 84.260 28.720 ;
        RECT 87.070 28.780 95.200 29.000 ;
        RECT 87.070 28.770 94.660 28.780 ;
        RECT 87.070 28.760 87.840 28.770 ;
        RECT 87.070 28.590 87.310 28.760 ;
        RECT 83.830 28.510 87.310 28.590 ;
        RECT 58.920 28.350 60.550 28.480 ;
        RECT 83.940 28.350 87.310 28.510 ;
        RECT 22.780 28.050 23.380 28.190 ;
        RECT 24.900 28.090 26.860 28.310 ;
        RECT 22.640 27.850 23.380 28.050 ;
        RECT 26.910 27.880 27.220 28.210 ;
        RECT 27.750 28.150 28.430 28.230 ;
        RECT 27.620 28.020 28.430 28.150 ;
        RECT 22.640 27.720 22.950 27.850 ;
        RECT 27.620 27.820 27.930 28.020 ;
        RECT 43.640 27.900 43.740 28.220 ;
        RECT 52.560 28.150 53.210 28.350 ;
        RECT 58.610 28.300 60.550 28.350 ;
        RECT 58.610 28.170 59.100 28.300 ;
        RECT 67.540 28.160 69.320 28.340 ;
        RECT 52.750 27.650 53.070 27.700 ;
        RECT 59.360 27.650 59.680 27.750 ;
        RECT 52.750 27.490 59.680 27.650 ;
        RECT 52.750 27.440 53.070 27.490 ;
        RECT 59.360 27.470 59.680 27.490 ;
        RECT 60.390 27.630 60.710 27.940 ;
        RECT 71.010 27.650 71.420 27.760 ;
        RECT 64.040 27.630 71.420 27.650 ;
        RECT 60.390 27.490 71.420 27.630 ;
        RECT 60.390 27.460 60.710 27.490 ;
        RECT 63.960 27.420 71.420 27.490 ;
        RECT 59.950 27.410 60.230 27.420 ;
        RECT 59.930 27.320 60.250 27.410 ;
        RECT 71.010 27.390 71.420 27.420 ;
        RECT 62.170 27.320 62.490 27.350 ;
        RECT 59.900 27.160 62.490 27.320 ;
        RECT 59.930 27.150 60.250 27.160 ;
        RECT 59.950 27.140 60.230 27.150 ;
        RECT 62.170 27.090 62.490 27.160 ;
        RECT 62.190 27.080 62.470 27.090 ;
        RECT 60.970 25.810 61.350 26.200 ;
        RECT 77.050 26.190 77.350 26.210 ;
        RECT 62.120 25.770 62.520 26.110 ;
        RECT 70.710 25.610 71.370 25.970 ;
        RECT 76.340 25.850 77.360 26.190 ;
        RECT 77.050 25.830 77.360 25.850 ;
        RECT 52.270 24.770 52.650 25.150 ;
        RECT 72.460 24.890 72.910 25.320 ;
        RECT 22.820 20.960 23.420 21.110 ;
        RECT 22.670 20.630 23.420 20.960 ;
        RECT 22.820 20.490 23.420 20.630 ;
        RECT 22.680 20.290 23.420 20.490 ;
        RECT 22.680 20.160 22.990 20.290 ;
        RECT 51.970 17.200 52.280 17.330 ;
        RECT 51.540 17.000 52.280 17.200 ;
        RECT 51.540 16.860 52.140 17.000 ;
        RECT 51.540 16.530 52.290 16.860 ;
        RECT 51.540 16.380 52.140 16.530 ;
        RECT 108.070 13.640 108.400 13.950 ;
        RECT 108.090 13.460 108.380 13.640 ;
        RECT 108.100 13.280 108.380 13.460 ;
        RECT 108.070 12.970 108.400 13.280 ;
        RECT 108.100 12.710 108.380 12.970 ;
        RECT 6.070 7.350 7.340 9.230 ;
        RECT 6.140 2.600 7.410 4.480 ;
        RECT 106.030 0.320 106.350 0.640 ;
      LAYER via2 ;
        RECT 83.890 54.130 84.230 54.470 ;
        RECT 82.820 50.650 83.150 51.000 ;
        RECT 83.910 48.080 84.250 48.440 ;
  END
END sky130_hilas_TopLevelTextStructure

MACRO sky130_hilas_pFETLarge
  CLASS CORE ;
  FOREIGN sky130_hilas_pFETLarge ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.640 BY 5.990 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA 6.540500 ;
    PORT
      LAYER met2 ;
        RECT 0.430 0.830 0.740 0.960 ;
        RECT 0.000 0.630 0.740 0.830 ;
        RECT 0.000 0.490 0.600 0.630 ;
        RECT 0.000 0.160 0.750 0.490 ;
        RECT 0.000 0.010 0.600 0.160 ;
    END
  END GATE
  PIN SOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 4.358700 ;
    PORT
      LAYER met2 ;
        RECT 1.010 5.610 1.320 5.750 ;
        RECT 2.100 5.610 2.410 5.750 ;
        RECT 3.200 5.610 3.510 5.740 ;
        RECT 0.330 5.600 3.510 5.610 ;
        RECT 0.240 5.410 3.510 5.600 ;
        RECT 0.240 5.270 3.390 5.410 ;
        RECT 0.240 2.820 0.560 5.270 ;
        RECT 1.000 2.820 1.310 2.970 ;
        RECT 2.100 2.820 2.410 2.970 ;
        RECT 3.200 2.820 3.510 2.970 ;
        RECT 0.240 2.640 3.510 2.820 ;
        RECT 0.240 2.490 3.400 2.640 ;
        RECT 0.240 1.450 0.560 2.490 ;
        RECT 1.000 1.450 1.310 1.600 ;
        RECT 2.100 1.450 2.410 1.600 ;
        RECT 3.200 1.450 3.510 1.600 ;
        RECT 0.240 1.270 3.510 1.450 ;
        RECT 0.240 1.130 3.400 1.270 ;
    END
  END SOURCE
  PIN DRAIN
    USE ANALOG ;
    ANTENNADIFFAREA 4.311400 ;
    PORT
      LAYER met2 ;
        RECT 1.560 4.890 1.870 5.070 ;
        RECT 2.650 4.890 2.960 5.050 ;
        RECT 3.760 4.890 4.070 5.040 ;
        RECT 1.430 4.590 4.370 4.890 ;
        RECT 3.620 4.550 4.370 4.590 ;
        RECT 3.990 4.420 4.370 4.550 ;
        RECT 4.020 3.700 4.370 4.420 ;
        RECT 1.560 3.550 1.870 3.700 ;
        RECT 2.650 3.550 2.960 3.700 ;
        RECT 3.750 3.550 4.370 3.700 ;
        RECT 1.420 3.220 4.370 3.550 ;
        RECT 4.020 0.930 4.370 3.220 ;
        RECT 1.560 0.780 1.870 0.920 ;
        RECT 2.650 0.780 2.960 0.920 ;
        RECT 3.750 0.780 4.370 0.930 ;
        RECT 1.430 0.460 4.370 0.780 ;
        RECT 1.430 0.450 4.140 0.460 ;
    END
  END DRAIN
  PIN WELL
    USE ANALOG ;
    ANTENNADIFFAREA 0.213200 ;
    PORT
      LAYER nwell ;
        RECT 0.780 5.880 4.170 5.970 ;
        RECT 0.780 0.270 4.640 5.880 ;
        RECT 4.020 0.180 4.640 0.270 ;
      LAYER met1 ;
        RECT 4.140 5.790 4.400 5.990 ;
        RECT 4.140 4.980 4.450 5.790 ;
        RECT 4.140 0.000 4.400 4.980 ;
    END
  END WELL
  OBS
      LAYER li1 ;
        RECT 1.020 5.710 1.190 5.740 ;
        RECT 1.020 5.670 1.340 5.710 ;
        RECT 1.020 5.480 1.350 5.670 ;
        RECT 1.020 5.450 1.340 5.480 ;
        RECT 1.020 3.250 1.190 5.450 ;
        RECT 1.570 5.030 1.740 5.740 ;
        RECT 2.120 5.710 2.290 5.740 ;
        RECT 2.110 5.670 2.430 5.710 ;
        RECT 2.110 5.480 2.440 5.670 ;
        RECT 2.110 5.450 2.430 5.480 ;
        RECT 1.570 4.990 1.890 5.030 ;
        RECT 1.570 4.800 1.900 4.990 ;
        RECT 1.570 4.770 1.890 4.800 ;
        RECT 1.570 3.660 1.740 4.770 ;
        RECT 1.570 3.620 1.890 3.660 ;
        RECT 1.570 3.430 1.900 3.620 ;
        RECT 1.570 3.400 1.890 3.430 ;
        RECT 1.570 3.240 1.740 3.400 ;
        RECT 2.120 3.240 2.290 5.450 ;
        RECT 2.670 5.010 2.840 5.740 ;
        RECT 3.220 5.700 3.390 5.740 ;
        RECT 3.210 5.660 3.530 5.700 ;
        RECT 3.210 5.470 3.540 5.660 ;
        RECT 3.210 5.440 3.530 5.470 ;
        RECT 2.660 4.970 2.980 5.010 ;
        RECT 2.660 4.780 2.990 4.970 ;
        RECT 2.660 4.750 2.980 4.780 ;
        RECT 2.670 3.660 2.840 4.750 ;
        RECT 2.660 3.620 2.980 3.660 ;
        RECT 2.660 3.430 2.990 3.620 ;
        RECT 2.660 3.400 2.980 3.430 ;
        RECT 2.670 3.240 2.840 3.400 ;
        RECT 3.220 3.240 3.390 5.440 ;
        RECT 3.770 5.000 3.940 5.740 ;
        RECT 3.770 4.960 4.090 5.000 ;
        RECT 3.770 4.770 4.100 4.960 ;
        RECT 4.250 4.920 4.420 5.680 ;
        RECT 3.770 4.740 4.090 4.770 ;
        RECT 3.770 3.660 3.940 4.740 ;
        RECT 3.760 3.620 4.080 3.660 ;
        RECT 3.760 3.430 4.090 3.620 ;
        RECT 3.760 3.400 4.080 3.430 ;
        RECT 3.770 3.240 3.940 3.400 ;
        RECT 0.960 3.160 1.120 3.190 ;
        RECT 0.960 2.930 1.130 3.160 ;
        RECT 1.510 3.150 1.670 3.190 ;
        RECT 0.960 2.890 1.330 2.930 ;
        RECT 1.510 2.910 1.680 3.150 ;
        RECT 2.060 2.930 2.230 3.220 ;
        RECT 2.610 3.150 2.770 3.190 ;
        RECT 3.160 3.150 3.320 3.190 ;
        RECT 3.710 3.170 3.870 3.190 ;
        RECT 0.960 2.810 1.340 2.890 ;
        RECT 1.510 2.810 1.740 2.910 ;
        RECT 2.060 2.890 2.430 2.930 ;
        RECT 2.610 2.910 2.780 3.150 ;
        RECT 3.160 2.930 3.330 3.150 ;
        RECT 2.060 2.810 2.440 2.890 ;
        RECT 2.610 2.810 2.840 2.910 ;
        RECT 3.160 2.890 3.530 2.930 ;
        RECT 3.710 2.910 3.880 3.170 ;
        RECT 3.160 2.810 3.540 2.890 ;
        RECT 3.710 2.810 3.940 2.910 ;
        RECT 1.010 2.700 1.340 2.810 ;
        RECT 1.010 2.670 1.330 2.700 ;
        RECT 1.020 1.560 1.190 2.670 ;
        RECT 1.010 1.520 1.330 1.560 ;
        RECT 1.010 1.330 1.340 1.520 ;
        RECT 1.010 1.300 1.330 1.330 ;
        RECT 0.190 0.940 0.700 1.020 ;
        RECT 0.190 0.920 0.710 0.940 ;
        RECT 0.190 0.880 0.760 0.920 ;
        RECT 0.190 0.690 0.770 0.880 ;
        RECT 0.200 0.660 0.760 0.690 ;
        RECT 0.200 0.450 0.710 0.660 ;
        RECT 0.200 0.410 0.770 0.450 ;
        RECT 1.020 0.420 1.190 1.300 ;
        RECT 1.570 0.880 1.740 2.810 ;
        RECT 2.110 2.700 2.440 2.810 ;
        RECT 2.110 2.670 2.430 2.700 ;
        RECT 2.120 1.560 2.290 2.670 ;
        RECT 2.110 1.520 2.430 1.560 ;
        RECT 2.110 1.330 2.440 1.520 ;
        RECT 2.110 1.300 2.430 1.330 ;
        RECT 1.570 0.840 1.890 0.880 ;
        RECT 1.570 0.650 1.900 0.840 ;
        RECT 1.570 0.620 1.890 0.650 ;
        RECT 1.570 0.410 1.740 0.620 ;
        RECT 2.120 0.410 2.290 1.300 ;
        RECT 2.670 0.880 2.840 2.810 ;
        RECT 3.210 2.700 3.540 2.810 ;
        RECT 3.210 2.670 3.530 2.700 ;
        RECT 3.220 1.560 3.390 2.670 ;
        RECT 3.210 1.520 3.530 1.560 ;
        RECT 3.210 1.330 3.540 1.520 ;
        RECT 3.210 1.300 3.530 1.330 ;
        RECT 2.660 0.840 2.980 0.880 ;
        RECT 2.660 0.650 2.990 0.840 ;
        RECT 2.660 0.620 2.980 0.650 ;
        RECT 2.670 0.410 2.840 0.620 ;
        RECT 3.220 0.410 3.390 1.300 ;
        RECT 3.770 0.890 3.940 2.810 ;
        RECT 3.760 0.850 4.080 0.890 ;
        RECT 3.760 0.660 4.090 0.850 ;
        RECT 3.760 0.630 4.080 0.660 ;
        RECT 3.770 0.410 3.940 0.630 ;
        RECT 0.200 0.220 0.780 0.410 ;
        RECT 0.200 0.190 0.770 0.220 ;
        RECT 0.200 0.010 0.710 0.190 ;
      LAYER mcon ;
        RECT 1.080 5.490 1.250 5.660 ;
        RECT 2.170 5.490 2.340 5.660 ;
        RECT 1.630 4.810 1.800 4.980 ;
        RECT 1.630 3.440 1.800 3.610 ;
        RECT 3.270 5.480 3.440 5.650 ;
        RECT 2.720 4.790 2.890 4.960 ;
        RECT 2.720 3.440 2.890 3.610 ;
        RECT 4.250 5.510 4.420 5.680 ;
        RECT 4.250 5.150 4.420 5.320 ;
        RECT 3.830 4.780 4.000 4.950 ;
        RECT 3.820 3.440 3.990 3.610 ;
        RECT 1.070 2.710 1.240 2.880 ;
        RECT 1.070 1.340 1.240 1.510 ;
        RECT 0.500 0.700 0.670 0.870 ;
        RECT 2.170 2.710 2.340 2.880 ;
        RECT 2.170 1.340 2.340 1.510 ;
        RECT 1.630 0.660 1.800 0.830 ;
        RECT 3.270 2.710 3.440 2.880 ;
        RECT 3.270 1.340 3.440 1.510 ;
        RECT 2.720 0.660 2.890 0.830 ;
        RECT 3.820 0.670 3.990 0.840 ;
        RECT 0.510 0.230 0.680 0.400 ;
      LAYER met1 ;
        RECT 1.010 5.420 1.330 5.740 ;
        RECT 2.100 5.420 2.420 5.740 ;
        RECT 3.200 5.410 3.520 5.730 ;
        RECT 1.560 4.740 1.880 5.060 ;
        RECT 2.650 4.720 2.970 5.040 ;
        RECT 3.760 4.710 4.080 5.030 ;
        RECT 1.560 3.370 1.880 3.690 ;
        RECT 2.650 3.370 2.970 3.690 ;
        RECT 3.750 3.370 4.070 3.690 ;
        RECT 1.000 2.640 1.320 2.960 ;
        RECT 2.100 2.640 2.420 2.960 ;
        RECT 3.200 2.640 3.520 2.960 ;
        RECT 1.000 1.270 1.320 1.590 ;
        RECT 2.100 1.270 2.420 1.590 ;
        RECT 3.200 1.270 3.520 1.590 ;
        RECT 0.430 0.630 0.750 0.950 ;
        RECT 1.560 0.590 1.880 0.910 ;
        RECT 2.650 0.590 2.970 0.910 ;
        RECT 3.750 0.600 4.070 0.920 ;
        RECT 0.440 0.160 0.760 0.480 ;
      LAYER via ;
        RECT 1.040 5.450 1.300 5.710 ;
        RECT 2.130 5.450 2.390 5.710 ;
        RECT 3.230 5.440 3.490 5.700 ;
        RECT 1.590 4.770 1.850 5.030 ;
        RECT 2.680 4.750 2.940 5.010 ;
        RECT 3.790 4.740 4.050 5.000 ;
        RECT 1.590 3.400 1.850 3.660 ;
        RECT 2.680 3.400 2.940 3.660 ;
        RECT 3.780 3.400 4.040 3.660 ;
        RECT 1.030 2.670 1.290 2.930 ;
        RECT 2.130 2.670 2.390 2.930 ;
        RECT 3.230 2.670 3.490 2.930 ;
        RECT 1.030 1.300 1.290 1.560 ;
        RECT 2.130 1.300 2.390 1.560 ;
        RECT 3.230 1.300 3.490 1.560 ;
        RECT 0.460 0.660 0.720 0.920 ;
        RECT 1.590 0.620 1.850 0.880 ;
        RECT 2.680 0.620 2.940 0.880 ;
        RECT 3.780 0.630 4.040 0.890 ;
        RECT 0.470 0.190 0.730 0.450 ;
  END
END sky130_hilas_pFETLarge

MACRO sky130_hilas_VinjInv2
  CLASS CORE ;
  FOREIGN sky130_hilas_VinjInv2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.610 BY 1.640 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 0.000 0.000 1.980 1.640 ;
      LAYER li1 ;
        RECT 0.620 1.210 0.790 1.350 ;
        RECT 0.620 1.040 0.810 1.210 ;
        RECT 0.620 0.940 0.790 1.040 ;
        RECT 0.190 0.560 0.360 0.660 ;
        RECT 0.170 0.390 0.360 0.560 ;
        RECT 0.190 0.330 0.360 0.390 ;
        RECT 0.610 0.600 0.780 0.660 ;
        RECT 0.610 0.330 0.860 0.600 ;
        RECT 1.350 0.580 1.600 0.660 ;
        RECT 1.350 0.410 2.650 0.580 ;
        RECT 3.210 0.570 3.380 1.200 ;
        RECT 0.620 0.310 0.860 0.330 ;
        RECT 1.430 0.320 1.600 0.410 ;
        RECT 3.130 0.400 3.460 0.570 ;
      LAYER mcon ;
        RECT 0.640 1.040 0.810 1.210 ;
        RECT 3.210 0.680 3.380 0.850 ;
        RECT 0.650 0.360 0.820 0.530 ;
        RECT 1.990 0.410 2.160 0.580 ;
      LAYER met1 ;
        RECT 0.610 1.260 0.830 1.600 ;
        RECT 0.610 1.000 0.840 1.260 ;
        RECT 0.080 0.320 0.390 0.670 ;
        RECT 0.610 0.600 0.830 1.000 ;
        RECT 0.610 0.290 0.860 0.600 ;
        RECT 1.910 0.360 2.230 0.620 ;
        RECT 0.610 0.090 0.830 0.290 ;
        RECT 3.180 0.090 3.410 1.600 ;
      LAYER via ;
        RECT 0.110 0.350 0.370 0.610 ;
        RECT 1.940 0.360 2.200 0.620 ;
      LAYER met2 ;
        RECT 0.000 1.030 3.610 1.210 ;
        RECT 0.080 0.510 0.400 0.610 ;
        RECT 0.070 0.350 0.400 0.510 ;
        RECT 1.910 0.540 2.230 0.620 ;
        RECT 1.910 0.360 3.610 0.540 ;
  END
END sky130_hilas_VinjInv2

MACRO sky130_hilas_capacitorSize03
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize03 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.720 BY 7.900 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.420 2.410 5.790 2.690 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.020 2.370 0.290 2.650 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 0.000 4.850 5.780 5.030 ;
        RECT 0.000 4.420 5.780 4.600 ;
        RECT 0.030 3.420 5.780 3.600 ;
        RECT 0.030 3.110 5.780 3.170 ;
        RECT 0.030 2.990 5.820 3.110 ;
        RECT 0.600 2.670 0.970 2.990 ;
        RECT 5.450 2.710 5.820 2.990 ;
        RECT 0.030 1.840 5.780 2.010 ;
        RECT 0.030 1.420 5.780 1.590 ;
        RECT 0.030 0.440 5.780 0.610 ;
        RECT 0.030 0.000 5.780 0.170 ;
      LAYER via2 ;
        RECT 0.650 2.730 0.930 3.010 ;
        RECT 5.500 2.770 5.780 3.050 ;
      LAYER met3 ;
        RECT 5.880 5.040 8.720 7.900 ;
        RECT 5.880 3.260 8.720 4.890 ;
        RECT 0.380 2.470 1.170 3.220 ;
        RECT 1.450 2.900 1.720 2.910 ;
        RECT 5.230 2.900 8.720 3.260 ;
        RECT 1.450 2.510 8.720 2.900 ;
        RECT 1.450 2.150 5.590 2.510 ;
        RECT 5.880 2.030 8.720 2.510 ;
      LAYER via3 ;
        RECT 0.570 2.620 1.000 3.100 ;
        RECT 5.420 2.660 5.850 3.140 ;
      LAYER met4 ;
        RECT 7.000 6.560 7.450 6.570 ;
        RECT 6.980 6.070 7.500 6.560 ;
        RECT 0.470 2.770 1.130 3.190 ;
        RECT 2.580 2.780 3.020 3.620 ;
        RECT 7.000 3.550 7.450 3.560 ;
        RECT 1.160 2.770 2.170 2.780 ;
        RECT 2.570 2.770 3.030 2.780 ;
        RECT 0.450 2.270 3.030 2.770 ;
        RECT 5.320 2.570 5.980 3.230 ;
        RECT 6.980 3.060 7.500 3.550 ;
        RECT 0.450 2.260 1.520 2.270 ;
        RECT 2.570 1.610 3.030 2.270 ;
        RECT 2.570 1.110 3.050 1.610 ;
        RECT 3.020 0.810 3.050 1.110 ;
  END
END sky130_hilas_capacitorSize03

MACRO sky130_hilas_swc4x1BiasCell
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x1BiasCell ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.250 BY 10.910 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN ROW1
    PORT
      LAYER met2 ;
        RECT 9.990 5.740 10.080 5.920 ;
    END
  END ROW1
  PIN ROW2
    PORT
      LAYER met2 ;
        RECT 9.990 4.650 10.080 4.830 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.010 4.650 7.640 4.830 ;
    END
  END ROW2
  PIN ROW3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.010 2.540 0.480 2.700 ;
        RECT 0.020 2.530 0.480 2.540 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.970 2.500 10.080 2.680 ;
    END
  END ROW3
  PIN ROW4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.010 1.550 7.640 1.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.970 1.400 10.080 1.580 ;
    END
  END ROW4
  PIN VTUN
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 0.360 0.410 0.760 6.910 ;
    END
  END VTUN
  PIN GATE1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 4.410 0.410 4.790 0.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.410 6.540 4.790 6.910 ;
    END
  END GATE1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 9.560 6.570 9.720 6.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 9.560 0.600 9.720 0.670 ;
    END
  END VINJ
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 8.750 6.570 8.910 6.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.750 0.600 8.910 0.670 ;
    END
  END VPWR
  PIN COLSEL1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 9.120 0.600 9.310 0.670 ;
    END
  END COLSEL1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 2.540 2.110 2.870 2.140 ;
        RECT 6.570 2.110 6.890 2.170 ;
        RECT 2.540 1.940 6.890 2.110 ;
        RECT 2.540 1.880 2.870 1.940 ;
        RECT 6.570 1.890 6.890 1.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.600 2.200 6.850 6.910 ;
        RECT 6.590 2.170 6.870 2.200 ;
        RECT 6.580 1.890 6.880 2.170 ;
        RECT 6.590 1.870 6.870 1.890 ;
        RECT 6.600 0.410 6.850 1.870 ;
      LAYER via ;
        RECT 6.600 1.900 6.860 2.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.570 2.170 2.840 6.910 ;
        RECT 2.550 1.860 2.860 2.170 ;
        RECT 2.570 0.410 2.840 1.860 ;
      LAYER via ;
        RECT 2.570 1.880 2.840 2.140 ;
    END
  END VGND
  PIN DRAIN3
    PORT
      LAYER met2 ;
        RECT 9.970 2.930 10.080 3.110 ;
    END
  END DRAIN3
  PIN DRAIN4
    PORT
      LAYER met2 ;
        RECT 9.970 0.970 10.080 1.150 ;
    END
  END DRAIN4
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 9.990 6.170 10.080 6.350 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 9.990 4.220 10.080 4.400 ;
    END
  END DRAIN2
  OBS
      LAYER nwell ;
        RECT 14.520 10.850 16.250 10.910 ;
        RECT 10.410 5.410 12.970 7.320 ;
        RECT 0.580 5.180 1.170 5.340 ;
        RECT 4.320 5.120 5.430 5.390 ;
        RECT 7.520 4.200 7.610 4.280 ;
        RECT 8.960 3.700 9.130 3.760 ;
        RECT 8.960 3.690 9.310 3.700 ;
        RECT 8.960 3.590 9.130 3.690 ;
        RECT 9.300 3.590 9.310 3.690 ;
        RECT 10.410 2.170 12.970 5.160 ;
        RECT 13.330 4.410 16.250 10.850 ;
        RECT 18.520 7.280 20.250 9.120 ;
        RECT 13.330 4.360 15.560 4.410 ;
        RECT 0.580 1.940 1.170 2.090 ;
        RECT 4.320 1.920 5.430 2.110 ;
        RECT 10.410 0.000 12.970 1.910 ;
      LAYER li1 ;
        RECT 14.910 7.800 15.460 8.230 ;
        RECT 18.940 7.730 19.490 8.160 ;
        RECT 10.650 6.970 10.970 7.010 ;
        RECT 10.650 6.850 10.980 6.970 ;
        RECT 10.650 6.750 11.090 6.850 ;
        RECT 10.750 6.680 11.090 6.750 ;
        RECT 12.370 6.580 12.570 6.930 ;
        RECT 10.650 6.420 10.970 6.460 ;
        RECT 10.650 6.230 10.980 6.420 ;
        RECT 10.650 6.200 11.090 6.230 ;
        RECT 10.750 6.060 11.090 6.200 ;
        RECT 11.640 5.960 11.840 6.560 ;
        RECT 12.370 6.550 12.580 6.580 ;
        RECT 12.360 5.960 12.580 6.550 ;
        RECT 2.620 4.890 2.790 5.420 ;
        RECT 6.640 4.860 6.810 5.390 ;
        RECT 10.750 4.370 11.090 4.510 ;
        RECT 10.650 4.340 11.090 4.370 ;
        RECT 2.630 2.960 2.800 4.130 ;
        RECT 6.650 3.000 6.820 4.190 ;
        RECT 10.650 4.150 10.980 4.340 ;
        RECT 10.650 4.110 10.970 4.150 ;
        RECT 11.640 4.010 11.840 4.610 ;
        RECT 12.360 4.020 12.580 4.610 ;
        RECT 12.370 3.990 12.580 4.020 ;
        RECT 10.750 3.820 11.090 3.890 ;
        RECT 8.870 3.590 9.310 3.760 ;
        RECT 10.650 3.720 11.090 3.820 ;
        RECT 10.650 3.610 10.980 3.720 ;
        RECT 10.650 3.510 11.090 3.610 ;
        RECT 10.750 3.440 11.090 3.510 ;
        RECT 12.370 3.340 12.570 3.990 ;
        RECT 10.650 3.180 10.970 3.220 ;
        RECT 10.650 2.990 10.980 3.180 ;
        RECT 10.650 2.960 11.090 2.990 ;
        RECT 10.750 2.820 11.090 2.960 ;
        RECT 11.640 2.720 11.840 3.320 ;
        RECT 12.370 3.310 12.580 3.340 ;
        RECT 12.360 2.720 12.580 3.310 ;
        RECT 10.750 1.120 11.090 1.260 ;
        RECT 10.650 1.090 11.090 1.120 ;
        RECT 10.650 0.900 10.980 1.090 ;
        RECT 10.650 0.860 10.970 0.900 ;
        RECT 11.640 0.760 11.840 1.360 ;
        RECT 12.360 0.770 12.580 1.360 ;
        RECT 12.370 0.740 12.580 0.770 ;
        RECT 10.750 0.570 11.090 0.640 ;
        RECT 10.650 0.470 11.090 0.570 ;
        RECT 10.650 0.350 10.980 0.470 ;
        RECT 12.370 0.390 12.570 0.740 ;
        RECT 10.650 0.310 10.970 0.350 ;
      LAYER mcon ;
        RECT 14.910 7.880 15.180 8.150 ;
        RECT 18.940 7.810 19.210 8.080 ;
        RECT 10.710 6.790 10.880 6.960 ;
        RECT 10.710 6.240 10.880 6.410 ;
        RECT 11.650 6.350 11.820 6.520 ;
        RECT 12.380 6.380 12.550 6.550 ;
        RECT 2.620 5.250 2.790 5.420 ;
        RECT 6.640 5.220 6.810 5.390 ;
        RECT 2.630 3.960 2.800 4.130 ;
        RECT 2.630 3.320 2.800 3.490 ;
        RECT 6.650 4.020 6.820 4.190 ;
        RECT 10.710 4.160 10.880 4.330 ;
        RECT 11.650 4.050 11.820 4.220 ;
        RECT 12.380 4.020 12.550 4.190 ;
        RECT 9.130 3.590 9.310 3.760 ;
        RECT 6.650 3.360 6.820 3.530 ;
        RECT 10.710 3.550 10.880 3.780 ;
        RECT 10.710 3.000 10.880 3.170 ;
        RECT 11.650 3.110 11.820 3.280 ;
        RECT 12.380 3.140 12.550 3.310 ;
        RECT 10.710 0.910 10.880 1.080 ;
        RECT 11.650 0.800 11.820 0.970 ;
        RECT 12.380 0.770 12.550 0.940 ;
        RECT 10.710 0.360 10.880 0.530 ;
      LAYER met1 ;
        RECT 10.640 6.720 10.960 7.040 ;
        RECT 9.120 6.570 9.310 6.640 ;
        RECT 11.640 6.580 11.800 7.310 ;
        RECT 11.640 6.560 11.840 6.580 ;
        RECT 10.640 6.170 10.960 6.490 ;
        RECT 11.620 6.320 11.850 6.560 ;
        RECT 11.640 6.270 11.850 6.320 ;
        RECT 12.010 6.270 12.200 7.260 ;
        RECT 12.450 6.610 12.610 7.310 ;
        RECT 11.640 5.410 11.800 6.270 ;
        RECT 12.030 6.150 12.200 6.270 ;
        RECT 12.040 5.410 12.200 6.150 ;
        RECT 12.340 6.060 12.610 6.610 ;
        RECT 12.340 6.010 12.620 6.060 ;
        RECT 12.450 5.920 12.620 6.010 ;
        RECT 12.450 5.410 12.610 5.920 ;
        RECT 10.640 4.080 10.960 4.400 ;
        RECT 11.640 4.300 11.800 5.160 ;
        RECT 12.040 4.420 12.200 5.160 ;
        RECT 12.450 4.650 12.610 5.160 ;
        RECT 12.450 4.560 12.620 4.650 ;
        RECT 12.030 4.300 12.200 4.420 ;
        RECT 11.640 4.250 11.850 4.300 ;
        RECT 11.620 4.010 11.850 4.250 ;
        RECT 11.640 3.990 11.840 4.010 ;
        RECT 9.100 3.760 9.340 3.790 ;
        RECT 8.910 3.670 9.340 3.760 ;
        RECT 8.750 3.660 9.340 3.670 ;
        RECT 9.560 3.660 9.720 3.670 ;
        RECT 8.910 3.590 9.340 3.660 ;
        RECT 9.100 3.560 9.340 3.590 ;
        RECT 9.200 3.460 9.310 3.560 ;
        RECT 10.640 3.480 10.960 3.850 ;
        RECT 11.640 3.340 11.800 3.990 ;
        RECT 11.640 3.320 11.840 3.340 ;
        RECT 10.640 2.930 10.960 3.250 ;
        RECT 11.620 3.080 11.850 3.320 ;
        RECT 11.640 3.030 11.850 3.080 ;
        RECT 12.010 3.030 12.200 4.300 ;
        RECT 12.340 4.510 12.620 4.560 ;
        RECT 12.340 3.960 12.610 4.510 ;
        RECT 13.980 4.360 14.360 10.860 ;
        RECT 14.850 7.340 15.240 9.200 ;
        RECT 18.880 7.270 19.270 9.130 ;
        RECT 12.450 3.370 12.610 3.960 ;
        RECT 11.640 2.170 11.800 3.030 ;
        RECT 12.030 2.910 12.200 3.030 ;
        RECT 12.040 2.170 12.200 2.910 ;
        RECT 12.340 2.820 12.610 3.370 ;
        RECT 12.340 2.770 12.620 2.820 ;
        RECT 12.450 2.680 12.620 2.770 ;
        RECT 12.450 2.170 12.610 2.680 ;
        RECT 10.640 0.830 10.960 1.150 ;
        RECT 11.640 1.050 11.800 1.910 ;
        RECT 12.040 1.170 12.200 1.910 ;
        RECT 12.450 1.400 12.610 1.910 ;
        RECT 12.450 1.310 12.620 1.400 ;
        RECT 12.030 1.050 12.200 1.170 ;
        RECT 11.640 1.000 11.850 1.050 ;
        RECT 11.620 0.760 11.850 1.000 ;
        RECT 11.640 0.740 11.840 0.760 ;
        RECT 10.640 0.280 10.960 0.600 ;
        RECT 11.640 0.010 11.800 0.740 ;
        RECT 12.010 0.060 12.200 1.050 ;
        RECT 12.340 1.260 12.620 1.310 ;
        RECT 12.340 0.710 12.610 1.260 ;
        RECT 12.450 0.010 12.610 0.710 ;
      LAYER via ;
        RECT 10.670 6.750 10.930 7.010 ;
        RECT 10.670 6.200 10.930 6.460 ;
        RECT 10.670 4.110 10.930 4.370 ;
        RECT 10.670 3.510 10.930 3.820 ;
        RECT 10.670 2.960 10.930 3.220 ;
        RECT 10.670 0.860 10.930 1.120 ;
        RECT 10.670 0.310 10.930 0.570 ;
      LAYER met2 ;
        RECT 10.640 6.760 10.950 7.050 ;
        RECT 10.640 6.720 12.970 6.760 ;
        RECT 10.790 6.580 12.970 6.720 ;
        RECT 10.640 6.330 10.950 6.500 ;
        RECT 10.410 6.150 10.500 6.330 ;
        RECT 10.640 6.170 12.970 6.330 ;
        RECT 10.800 6.150 12.970 6.170 ;
        RECT 0.010 5.730 7.620 5.920 ;
        RECT 10.410 4.240 10.500 4.420 ;
        RECT 10.800 4.400 12.970 4.420 ;
        RECT 10.640 4.240 12.970 4.400 ;
        RECT 7.520 4.210 7.610 4.240 ;
        RECT 7.520 4.100 7.640 4.210 ;
        RECT 10.640 4.070 10.950 4.240 ;
        RECT 10.790 3.850 12.970 3.990 ;
        RECT 10.640 3.810 12.970 3.850 ;
        RECT 10.640 3.520 10.950 3.810 ;
        RECT 10.640 3.480 12.970 3.520 ;
        RECT 10.790 3.340 12.970 3.480 ;
        RECT 7.490 2.950 7.640 3.120 ;
        RECT 10.640 3.090 10.950 3.260 ;
        RECT 10.410 2.910 10.500 3.090 ;
        RECT 10.640 2.930 12.970 3.090 ;
        RECT 10.800 2.910 12.970 2.930 ;
        RECT 0.780 2.510 7.640 2.680 ;
        RECT 10.410 0.990 10.500 1.170 ;
        RECT 10.800 1.150 12.970 1.170 ;
        RECT 10.640 0.990 12.970 1.150 ;
        RECT 10.640 0.820 10.950 0.990 ;
        RECT 10.790 0.600 12.970 0.740 ;
        RECT 10.640 0.560 12.970 0.600 ;
        RECT 10.640 0.270 10.950 0.560 ;
  END
END sky130_hilas_swc4x1BiasCell

MACRO sky130_hilas_FGtrans2x1cell
  CLASS CORE ;
  FOREIGN sky130_hilas_FGtrans2x1cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.570 BY 10.520 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN COLSEL1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 16.850 6.460 17.040 6.520 ;
    END
    PORT
      LAYER met1 ;
        RECT 16.850 0.470 17.040 0.520 ;
    END
  END COLSEL1
  PIN VINJ
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 17.290 0.470 17.450 0.520 ;
    END
  END VINJ
  PIN DRAIN1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 17.730 5.840 17.810 6.020 ;
    END
  END DRAIN1
  PIN DRAIN2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 17.730 0.970 17.810 1.150 ;
    END
  END DRAIN2
  PIN PROG
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 14.080 4.060 14.290 6.520 ;
        RECT 14.080 3.550 14.410 4.060 ;
        RECT 14.080 0.470 14.290 3.550 ;
    END
  END PROG
  PIN RUN
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 13.030 1.990 13.210 6.520 ;
        RECT 12.980 1.650 13.270 1.990 ;
        RECT 13.030 0.470 13.210 1.650 ;
    END
  END RUN
  PIN VIN2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 14.960 3.170 15.150 3.220 ;
        RECT 14.960 2.880 15.270 3.170 ;
        RECT 14.960 1.260 15.150 2.880 ;
        RECT 14.960 0.970 15.250 1.260 ;
        RECT 14.930 0.470 15.160 0.970 ;
    END
  END VIN2
  PIN VIN1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 14.960 6.230 15.170 6.520 ;
        RECT 14.960 5.940 15.280 6.230 ;
        RECT 14.960 4.240 15.170 5.940 ;
        RECT 14.960 3.950 15.280 4.240 ;
        RECT 14.960 3.730 15.170 3.950 ;
    END
  END VIN1
  PIN GATE1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 14.510 5.670 14.700 6.520 ;
        RECT 14.510 5.380 14.810 5.670 ;
        RECT 14.510 3.350 14.700 5.380 ;
        RECT 14.510 3.060 14.810 3.350 ;
        RECT 14.510 1.770 14.700 3.060 ;
        RECT 14.510 1.480 14.820 1.770 ;
        RECT 14.510 0.470 14.700 1.480 ;
    END
  END GATE1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 9.110 3.660 9.340 6.520 ;
        RECT 9.110 3.370 9.440 3.660 ;
        RECT 9.110 0.470 9.340 3.370 ;
    END
  END VGND
  PIN VTUN
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 6.630 0.470 7.050 6.520 ;
    END
  END VTUN
  PIN DRAIN2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 15.340 1.140 15.500 1.160 ;
        RECT 6.290 1.090 15.500 1.140 ;
        RECT 6.290 0.990 15.380 1.090 ;
    END
  END DRAIN2
  PIN DRAIN1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 15.080 6.020 15.400 6.040 ;
        RECT 6.290 5.840 15.400 6.020 ;
    END
  END DRAIN1
  PIN COL1
    PORT
      LAYER met2 ;
        RECT 6.290 3.560 16.450 3.600 ;
        RECT 6.290 3.370 16.460 3.560 ;
    END
  END COL1
  PIN ROW1
    PORT
      LAYER met2 ;
        RECT 15.860 4.480 16.170 4.650 ;
        RECT 6.290 4.320 16.170 4.480 ;
        RECT 6.290 4.290 16.000 4.320 ;
    END
  END ROW1
  PIN ROW2
    PORT
      LAYER met2 ;
        RECT 6.290 2.430 16.010 2.620 ;
    END
  END ROW2
  OBS
      LAYER nwell ;
        RECT 20.800 10.180 22.530 10.520 ;
        RECT 20.780 8.620 22.530 10.180 ;
        RECT 20.780 6.990 22.510 8.620 ;
        RECT 0.010 6.560 2.720 6.600 ;
        RECT 0.000 4.910 2.720 6.560 ;
        RECT 0.000 0.330 2.720 1.980 ;
        RECT 6.870 1.870 7.430 4.290 ;
        RECT 19.260 3.820 22.570 6.990 ;
        RECT 6.630 0.480 7.050 0.550 ;
        RECT 0.010 0.290 2.720 0.330 ;
        RECT 19.260 0.000 22.570 3.170 ;
      LAYER li1 ;
        RECT 21.200 8.790 21.750 9.220 ;
        RECT 21.200 7.060 21.750 7.490 ;
        RECT 20.160 6.360 20.690 6.530 ;
        RECT 21.970 6.260 22.170 6.610 ;
        RECT 21.970 6.230 22.180 6.260 ;
        RECT 2.190 5.430 2.420 6.120 ;
        RECT 14.100 5.920 14.980 6.090 ;
        RECT 15.070 5.970 15.260 6.200 ;
        RECT 14.100 5.530 14.270 5.920 ;
        RECT 18.290 5.780 18.640 5.950 ;
        RECT 19.660 5.780 19.990 5.950 ;
        RECT 13.880 5.360 14.270 5.530 ;
        RECT 14.600 5.530 14.790 5.640 ;
        RECT 14.600 5.410 14.900 5.530 ;
        RECT 14.680 5.360 14.900 5.410 ;
        RECT 18.290 4.990 18.640 5.160 ;
        RECT 19.660 4.990 19.990 5.160 ;
        RECT 12.450 4.570 13.530 4.740 ;
        RECT 13.860 4.570 14.940 4.740 ;
        RECT 15.870 4.570 16.190 4.610 ;
        RECT 15.870 4.380 16.200 4.570 ;
        RECT 15.870 4.350 16.190 4.380 ;
        RECT 9.320 3.630 9.510 3.950 ;
        RECT 9.230 3.540 9.510 3.630 ;
        RECT 9.230 3.400 12.870 3.540 ;
        RECT 9.320 3.360 12.870 3.400 ;
        RECT 9.320 2.940 9.510 3.360 ;
        RECT 13.620 3.210 13.790 3.780 ;
        RECT 14.190 3.630 14.400 4.060 ;
        RECT 15.070 3.980 15.260 4.210 ;
        RECT 18.300 4.200 18.640 4.370 ;
        RECT 19.660 4.200 19.990 4.370 ;
        RECT 20.410 4.280 20.580 5.970 ;
        RECT 21.240 4.370 21.410 5.980 ;
        RECT 21.960 5.650 22.180 6.230 ;
        RECT 21.970 5.640 22.180 5.650 ;
        RECT 21.610 5.470 21.800 5.480 ;
        RECT 21.610 5.180 21.810 5.470 ;
        RECT 21.600 4.850 21.870 5.180 ;
        RECT 21.240 4.180 21.420 4.370 ;
        RECT 14.880 3.780 14.960 3.950 ;
        RECT 14.210 3.610 14.380 3.630 ;
        RECT 13.800 3.180 13.880 3.190 ;
        RECT 14.460 3.180 14.510 3.190 ;
        RECT 13.800 3.140 14.510 3.180 ;
        RECT 13.780 3.100 14.510 3.140 ;
        RECT 13.710 2.980 14.550 3.100 ;
        RECT 14.600 3.090 14.790 3.320 ;
        RECT 14.880 3.040 14.930 3.210 ;
        RECT 15.060 2.910 15.250 3.140 ;
        RECT 15.880 2.880 16.200 2.920 ;
        RECT 15.880 2.690 16.210 2.880 ;
        RECT 15.880 2.660 16.200 2.690 ;
        RECT 18.300 2.620 18.640 2.790 ;
        RECT 19.660 2.620 19.990 2.790 ;
        RECT 12.300 2.250 13.540 2.420 ;
        RECT 13.860 2.250 14.940 2.420 ;
        RECT 13.040 1.930 13.210 1.990 ;
        RECT 13.020 1.720 13.230 1.930 ;
        RECT 18.290 1.830 18.640 2.000 ;
        RECT 19.660 1.830 19.990 2.000 ;
        RECT 13.040 1.650 13.210 1.720 ;
        RECT 14.610 1.630 14.800 1.740 ;
        RECT 13.880 1.620 14.340 1.630 ;
        RECT 13.870 1.470 14.340 1.620 ;
        RECT 14.610 1.510 14.900 1.630 ;
        RECT 13.880 1.460 14.340 1.470 ;
        RECT 14.690 1.460 14.900 1.510 ;
        RECT 2.190 0.770 2.420 1.460 ;
        RECT 14.150 1.120 14.340 1.460 ;
        RECT 15.040 1.120 15.230 1.230 ;
        RECT 14.150 1.000 15.230 1.120 ;
        RECT 18.290 1.040 18.640 1.210 ;
        RECT 19.660 1.040 19.990 1.210 ;
        RECT 20.410 1.020 20.580 2.710 ;
        RECT 21.240 2.620 21.420 2.810 ;
        RECT 21.240 1.010 21.410 2.620 ;
        RECT 21.600 1.810 21.870 2.140 ;
        RECT 21.610 1.520 21.810 1.810 ;
        RECT 21.610 1.510 21.800 1.520 ;
        RECT 21.970 1.340 22.180 1.350 ;
        RECT 14.150 0.940 15.110 1.000 ;
        RECT 21.960 0.760 22.180 1.340 ;
        RECT 21.970 0.730 22.180 0.760 ;
        RECT 20.160 0.460 20.690 0.630 ;
        RECT 21.970 0.380 22.170 0.730 ;
      LAYER mcon ;
        RECT 21.200 8.870 21.470 9.140 ;
        RECT 21.200 7.140 21.470 7.410 ;
        RECT 2.220 5.910 2.390 6.080 ;
        RECT 2.220 5.460 2.390 5.630 ;
        RECT 15.080 6.000 15.250 6.170 ;
        RECT 21.980 6.060 22.150 6.230 ;
        RECT 14.610 5.440 14.780 5.610 ;
        RECT 15.930 4.390 16.100 4.560 ;
        RECT 21.620 5.220 21.800 5.410 ;
        RECT 15.080 4.010 15.250 4.180 ;
        RECT 9.240 3.430 9.410 3.600 ;
        RECT 14.610 3.120 14.780 3.290 ;
        RECT 15.070 2.940 15.240 3.110 ;
        RECT 15.940 2.700 16.110 2.870 ;
        RECT 14.620 1.540 14.790 1.710 ;
        RECT 2.220 1.260 2.390 1.430 ;
        RECT 2.220 0.810 2.390 0.980 ;
        RECT 15.050 1.030 15.220 1.200 ;
        RECT 21.620 1.580 21.800 1.770 ;
        RECT 21.980 0.760 22.150 0.930 ;
      LAYER met1 ;
        RECT 21.140 6.600 21.530 10.190 ;
        RECT 17.290 6.470 17.450 6.520 ;
        RECT 2.180 5.380 2.440 6.170 ;
        RECT 20.090 6.120 20.400 6.560 ;
        RECT 21.610 5.480 21.800 6.930 ;
        RECT 22.050 6.290 22.210 6.930 ;
        RECT 21.940 5.740 22.210 6.290 ;
        RECT 21.940 5.690 22.220 5.740 ;
        RECT 22.050 5.600 22.220 5.690 ;
        RECT 21.610 5.450 21.830 5.480 ;
        RECT 21.590 5.180 21.840 5.450 ;
        RECT 21.600 5.170 21.840 5.180 ;
        RECT 21.600 4.930 21.830 5.170 ;
        RECT 15.860 4.320 16.180 4.640 ;
        RECT 21.210 4.120 21.450 4.500 ;
        RECT 21.640 3.910 21.800 4.930 ;
        RECT 22.050 3.910 22.210 5.600 ;
        RECT 16.550 3.700 16.810 3.760 ;
        RECT 16.450 3.440 16.810 3.700 ;
        RECT 16.450 3.280 16.690 3.440 ;
        RECT 15.870 2.630 16.190 2.950 ;
        RECT 21.210 2.490 21.450 2.870 ;
        RECT 21.640 2.060 21.800 3.080 ;
        RECT 21.600 1.820 21.830 2.060 ;
        RECT 21.600 1.810 21.840 1.820 ;
        RECT 21.590 1.540 21.840 1.810 ;
        RECT 21.610 1.510 21.830 1.540 ;
        RECT 2.180 0.720 2.440 1.510 ;
        RECT 15.460 0.970 15.470 0.980 ;
        RECT 20.090 0.430 20.400 0.870 ;
        RECT 21.610 0.060 21.800 1.510 ;
        RECT 22.050 1.390 22.210 3.080 ;
        RECT 22.050 1.300 22.220 1.390 ;
        RECT 21.940 1.250 22.220 1.300 ;
        RECT 21.940 0.700 22.210 1.250 ;
        RECT 22.050 0.060 22.210 0.700 ;
      LAYER via ;
        RECT 20.120 6.150 20.380 6.410 ;
        RECT 15.890 4.350 16.150 4.610 ;
        RECT 16.550 3.470 16.810 3.730 ;
        RECT 15.900 2.660 16.160 2.920 ;
        RECT 20.120 0.580 20.380 0.840 ;
      LAYER met2 ;
        RECT 20.090 6.440 20.400 6.450 ;
        RECT 20.090 6.260 22.570 6.440 ;
        RECT 20.090 6.120 20.400 6.260 ;
        RECT 16.520 3.470 16.840 3.730 ;
        RECT 15.870 2.630 16.180 2.960 ;
        RECT 20.090 0.730 20.400 0.870 ;
        RECT 20.090 0.550 22.570 0.730 ;
        RECT 20.090 0.540 20.400 0.550 ;
  END
END sky130_hilas_FGtrans2x1cell

MACRO sky130_hilas_capacitorSize01
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.090 BY 7.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 10.060 2.380 10.420 2.660 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.020 2.370 0.290 2.650 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 0.000 4.850 10.420 5.030 ;
        RECT 0.000 4.420 10.420 4.600 ;
        RECT 0.030 3.420 10.420 3.600 ;
        RECT 8.510 3.170 10.420 3.180 ;
        RECT 0.030 3.080 10.420 3.170 ;
        RECT 0.030 2.990 10.460 3.080 ;
        RECT 0.600 2.670 0.970 2.990 ;
        RECT 10.090 2.680 10.460 2.990 ;
        RECT 0.030 1.840 10.420 2.010 ;
        RECT 0.030 1.420 10.420 1.590 ;
        RECT 0.030 0.440 10.420 0.610 ;
        RECT 0.030 0.000 10.420 0.170 ;
      LAYER via2 ;
        RECT 0.650 2.730 0.930 3.010 ;
        RECT 10.140 2.740 10.420 3.020 ;
      LAYER met3 ;
        RECT 5.890 7.840 8.710 7.870 ;
        RECT 0.380 2.470 1.170 3.220 ;
        RECT 5.890 2.060 13.090 7.840 ;
        RECT 8.680 2.040 13.090 2.060 ;
      LAYER via3 ;
        RECT 0.570 2.620 1.000 3.100 ;
        RECT 10.060 2.630 10.490 3.110 ;
      LAYER met4 ;
        RECT 0.470 2.770 1.130 3.190 ;
        RECT 6.780 3.140 9.820 3.610 ;
        RECT 1.160 2.770 2.170 2.780 ;
        RECT 0.450 2.270 3.800 2.770 ;
        RECT 9.960 2.540 10.620 3.200 ;
        RECT 0.450 2.260 1.520 2.270 ;
        RECT 3.160 1.150 3.790 2.270 ;
        RECT 3.160 0.850 5.310 1.150 ;
        RECT 3.490 0.840 5.310 0.850 ;
  END
END sky130_hilas_capacitorSize01

MACRO sky130_hilas_Tgate4Double01
  CLASS CORE ;
  FOREIGN sky130_hilas_Tgate4Double01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.710 BY 6.950 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.740 6.460 0.940 6.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.570 0.450 6.760 0.490 ;
    END
  END VGND
  PIN INPUT1_1
    PORT
      LAYER met2 ;
        RECT 0.000 6.190 0.050 6.390 ;
    END
  END INPUT1_1
  PIN SELECT1
    PORT
      LAYER met2 ;
        RECT 0.000 5.210 0.060 5.410 ;
    END
  END SELECT1
  PIN SELECT2
    PORT
      LAYER met2 ;
        RECT 0.000 4.560 0.060 4.760 ;
    END
  END SELECT2
  PIN INPUT2_2
    PORT
      LAYER met2 ;
        RECT 0.000 4.060 0.050 4.260 ;
    END
  END INPUT2_2
  PIN INPUT1_2
    PORT
      LAYER met2 ;
        RECT 0.000 3.580 0.050 3.780 ;
    END
  END INPUT1_2
  PIN SELECT3
    PORT
      LAYER met2 ;
        RECT 0.000 2.190 0.060 2.390 ;
    END
  END SELECT3
  PIN INPUT2_3
    PORT
      LAYER met2 ;
        RECT 0.000 2.690 0.050 2.890 ;
    END
  END INPUT2_3
  PIN SELECT4
    PORT
      LAYER met2 ;
        RECT 0.000 1.540 0.060 1.740 ;
    END
  END SELECT4
  PIN INPUT2_4
    PORT
      LAYER met2 ;
        RECT 0.000 1.040 0.050 1.240 ;
    END
  END INPUT2_4
  PIN INPUT1_4
    PORT
      LAYER met2 ;
        RECT 0.000 0.560 0.050 0.760 ;
    END
  END INPUT1_4
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 6.570 6.460 6.760 6.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.740 0.450 0.940 0.490 ;
    END
  END VPWR
  PIN OUTPUT4
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 7.020 1.560 7.080 1.740 ;
        RECT 2.630 1.410 8.400 1.560 ;
        RECT 2.630 1.360 8.610 1.410 ;
        RECT 5.220 1.090 5.530 1.360 ;
        RECT 8.300 1.080 8.610 1.360 ;
    END
  END OUTPUT4
  PIN OUTPUT3
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 5.220 2.570 5.530 2.840 ;
        RECT 8.300 2.570 8.610 2.850 ;
        RECT 2.630 2.520 8.610 2.570 ;
        RECT 2.630 2.370 8.400 2.520 ;
        RECT 7.020 2.190 7.080 2.370 ;
    END
  END OUTPUT3
  PIN OUTPUT2
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 7.020 4.580 7.080 4.760 ;
        RECT 2.630 4.430 8.400 4.580 ;
        RECT 2.630 4.380 8.610 4.430 ;
        RECT 5.220 4.110 5.530 4.380 ;
        RECT 8.300 4.100 8.610 4.380 ;
    END
  END OUTPUT2
  PIN OUTPUT1
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 5.220 5.590 5.530 5.860 ;
        RECT 8.300 5.590 8.610 5.870 ;
        RECT 2.630 5.540 8.610 5.590 ;
        RECT 2.630 5.390 8.400 5.540 ;
        RECT 7.010 5.210 7.080 5.390 ;
    END
  END OUTPUT1
  PIN INPUT2_1
    PORT
      LAYER met2 ;
        RECT 0.000 5.710 0.050 5.910 ;
    END
  END INPUT2_1
  PIN INPUT1_3
    PORT
      LAYER met2 ;
        RECT 0.000 3.170 0.050 3.370 ;
    END
  END INPUT1_3
  OBS
      LAYER nwell ;
        RECT 2.750 5.280 6.220 6.800 ;
        RECT 2.750 2.260 6.220 4.690 ;
        RECT 2.750 0.150 6.220 1.670 ;
      LAYER li1 ;
        RECT 2.960 6.520 3.170 6.950 ;
        RECT 2.980 6.500 3.150 6.520 ;
        RECT 3.480 6.380 3.670 6.490 ;
        RECT 3.480 6.260 3.900 6.380 ;
        RECT 3.380 6.210 3.900 6.260 ;
        RECT 4.250 6.210 8.470 6.390 ;
        RECT 8.850 6.220 9.200 6.390 ;
        RECT 9.300 6.380 9.490 6.490 ;
        RECT 9.300 6.260 9.630 6.380 ;
        RECT 3.380 6.130 3.570 6.210 ;
        RECT 3.360 6.100 3.570 6.130 ;
        RECT 3.350 6.090 3.570 6.100 ;
        RECT 3.230 6.040 3.570 6.090 ;
        RECT 3.100 6.010 3.570 6.040 ;
        RECT 3.060 5.980 3.570 6.010 ;
        RECT 3.880 6.150 4.200 6.190 ;
        RECT 3.060 5.920 3.550 5.980 ;
        RECT 3.880 5.960 4.210 6.150 ;
        RECT 4.740 6.090 5.070 6.210 ;
        RECT 6.800 6.150 7.120 6.190 ;
        RECT 9.380 6.180 9.630 6.260 ;
        RECT 4.450 5.990 4.640 6.080 ;
        RECT 3.880 5.930 4.200 5.960 ;
        RECT 3.060 5.870 3.400 5.920 ;
        RECT 3.060 5.850 3.320 5.870 ;
        RECT 4.340 5.850 4.640 5.990 ;
        RECT 5.900 5.870 6.090 6.100 ;
        RECT 6.800 5.960 7.130 6.150 ;
        RECT 6.800 5.930 7.120 5.960 ;
        RECT 7.610 5.870 7.800 6.090 ;
        RECT 7.510 5.860 7.800 5.870 ;
        RECT 3.060 5.830 3.290 5.850 ;
        RECT 3.060 5.790 3.270 5.830 ;
        RECT 3.060 5.510 3.230 5.790 ;
        RECT 3.740 5.750 3.920 5.790 ;
        RECT 3.570 5.580 3.920 5.750 ;
        RECT 4.340 5.500 4.510 5.850 ;
        RECT 5.120 5.820 5.290 5.840 ;
        RECT 5.120 5.780 5.550 5.820 ;
        RECT 5.120 5.590 5.560 5.780 ;
        RECT 5.120 5.560 5.550 5.590 ;
        RECT 5.120 5.540 5.290 5.560 ;
        RECT 5.810 5.500 5.980 5.850 ;
        RECT 6.770 5.500 6.940 5.800 ;
        RECT 7.510 5.490 7.680 5.860 ;
        RECT 8.230 5.830 8.400 5.840 ;
        RECT 8.230 5.790 8.630 5.830 ;
        RECT 8.230 5.600 8.640 5.790 ;
        RECT 8.840 5.760 9.030 5.870 ;
        RECT 8.840 5.640 9.180 5.760 ;
        RECT 8.230 5.570 8.630 5.600 ;
        RECT 8.890 5.590 9.180 5.640 ;
        RECT 8.230 5.540 8.400 5.570 ;
        RECT 9.460 5.500 9.630 6.180 ;
        RECT 3.060 4.180 3.230 4.460 ;
        RECT 3.570 4.220 3.920 4.390 ;
        RECT 3.740 4.180 3.920 4.220 ;
        RECT 3.060 4.140 3.270 4.180 ;
        RECT 3.060 4.120 3.290 4.140 ;
        RECT 4.340 4.120 4.510 4.470 ;
        RECT 5.120 4.410 5.290 4.430 ;
        RECT 5.120 4.380 5.550 4.410 ;
        RECT 5.120 4.190 5.560 4.380 ;
        RECT 5.120 4.150 5.550 4.190 ;
        RECT 5.120 4.130 5.290 4.150 ;
        RECT 5.810 4.120 5.980 4.470 ;
        RECT 6.770 4.170 6.940 4.470 ;
        RECT 3.060 4.100 3.320 4.120 ;
        RECT 3.060 4.050 3.400 4.100 ;
        RECT 3.060 3.990 3.550 4.050 ;
        RECT 3.880 4.010 4.200 4.040 ;
        RECT 3.060 3.960 3.570 3.990 ;
        RECT 3.100 3.930 3.570 3.960 ;
        RECT 2.960 3.500 3.170 3.930 ;
        RECT 3.230 3.880 3.570 3.930 ;
        RECT 3.350 3.870 3.570 3.880 ;
        RECT 3.360 3.840 3.570 3.870 ;
        RECT 3.380 3.760 3.570 3.840 ;
        RECT 3.880 3.820 4.210 4.010 ;
        RECT 4.340 3.980 4.640 4.120 ;
        RECT 7.510 4.110 7.680 4.480 ;
        RECT 8.230 4.400 8.400 4.430 ;
        RECT 8.230 4.370 8.630 4.400 ;
        RECT 8.230 4.180 8.640 4.370 ;
        RECT 8.890 4.330 9.180 4.380 ;
        RECT 8.840 4.210 9.180 4.330 ;
        RECT 8.230 4.140 8.630 4.180 ;
        RECT 8.230 4.130 8.400 4.140 ;
        RECT 7.510 4.100 7.800 4.110 ;
        RECT 8.840 4.100 9.030 4.210 ;
        RECT 4.450 3.890 4.640 3.980 ;
        RECT 3.880 3.780 4.200 3.820 ;
        RECT 4.740 3.760 5.070 3.880 ;
        RECT 5.900 3.870 6.090 4.100 ;
        RECT 6.800 4.010 7.120 4.040 ;
        RECT 6.800 3.820 7.130 4.010 ;
        RECT 7.610 3.880 7.800 4.100 ;
        RECT 6.800 3.780 7.120 3.820 ;
        RECT 9.460 3.790 9.630 4.470 ;
        RECT 3.380 3.710 3.900 3.760 ;
        RECT 3.480 3.590 3.900 3.710 ;
        RECT 2.980 3.480 3.150 3.500 ;
        RECT 3.480 3.480 3.670 3.590 ;
        RECT 4.250 3.580 8.470 3.760 ;
        RECT 8.850 3.580 9.200 3.750 ;
        RECT 9.380 3.710 9.630 3.790 ;
        RECT 9.300 3.590 9.630 3.710 ;
        RECT 9.300 3.480 9.490 3.590 ;
        RECT 2.980 3.450 3.150 3.470 ;
        RECT 2.960 3.020 3.170 3.450 ;
        RECT 3.480 3.360 3.670 3.470 ;
        RECT 3.480 3.240 3.900 3.360 ;
        RECT 3.380 3.190 3.900 3.240 ;
        RECT 4.250 3.190 8.470 3.370 ;
        RECT 8.850 3.200 9.200 3.370 ;
        RECT 9.300 3.360 9.490 3.470 ;
        RECT 9.300 3.240 9.630 3.360 ;
        RECT 3.380 3.110 3.570 3.190 ;
        RECT 3.360 3.080 3.570 3.110 ;
        RECT 3.350 3.070 3.570 3.080 ;
        RECT 3.230 3.020 3.570 3.070 ;
        RECT 3.100 2.990 3.570 3.020 ;
        RECT 3.060 2.960 3.570 2.990 ;
        RECT 3.880 3.130 4.200 3.170 ;
        RECT 3.060 2.900 3.550 2.960 ;
        RECT 3.880 2.940 4.210 3.130 ;
        RECT 4.740 3.070 5.070 3.190 ;
        RECT 6.800 3.130 7.120 3.170 ;
        RECT 9.380 3.160 9.630 3.240 ;
        RECT 4.450 2.970 4.640 3.060 ;
        RECT 3.880 2.910 4.200 2.940 ;
        RECT 3.060 2.850 3.400 2.900 ;
        RECT 3.060 2.830 3.320 2.850 ;
        RECT 4.340 2.830 4.640 2.970 ;
        RECT 5.900 2.850 6.090 3.080 ;
        RECT 6.800 2.940 7.130 3.130 ;
        RECT 6.800 2.910 7.120 2.940 ;
        RECT 7.610 2.850 7.800 3.070 ;
        RECT 7.510 2.840 7.800 2.850 ;
        RECT 3.060 2.810 3.290 2.830 ;
        RECT 3.060 2.770 3.270 2.810 ;
        RECT 3.060 2.490 3.230 2.770 ;
        RECT 3.740 2.730 3.920 2.770 ;
        RECT 3.570 2.560 3.920 2.730 ;
        RECT 4.340 2.480 4.510 2.830 ;
        RECT 5.120 2.800 5.290 2.820 ;
        RECT 5.120 2.760 5.550 2.800 ;
        RECT 5.120 2.570 5.560 2.760 ;
        RECT 5.120 2.540 5.550 2.570 ;
        RECT 5.120 2.520 5.290 2.540 ;
        RECT 5.810 2.480 5.980 2.830 ;
        RECT 6.770 2.480 6.940 2.780 ;
        RECT 7.510 2.470 7.680 2.840 ;
        RECT 8.230 2.810 8.400 2.820 ;
        RECT 8.230 2.770 8.630 2.810 ;
        RECT 8.230 2.580 8.640 2.770 ;
        RECT 8.840 2.740 9.030 2.850 ;
        RECT 8.840 2.620 9.180 2.740 ;
        RECT 8.230 2.550 8.630 2.580 ;
        RECT 8.890 2.570 9.180 2.620 ;
        RECT 8.230 2.520 8.400 2.550 ;
        RECT 9.460 2.480 9.630 3.160 ;
        RECT 3.060 1.160 3.230 1.440 ;
        RECT 3.570 1.200 3.920 1.370 ;
        RECT 3.740 1.160 3.920 1.200 ;
        RECT 3.060 1.120 3.270 1.160 ;
        RECT 3.060 1.100 3.290 1.120 ;
        RECT 4.340 1.100 4.510 1.450 ;
        RECT 5.120 1.390 5.290 1.410 ;
        RECT 5.120 1.360 5.550 1.390 ;
        RECT 5.120 1.170 5.560 1.360 ;
        RECT 5.120 1.130 5.550 1.170 ;
        RECT 5.120 1.110 5.290 1.130 ;
        RECT 5.810 1.100 5.980 1.450 ;
        RECT 6.770 1.150 6.940 1.450 ;
        RECT 3.060 1.080 3.320 1.100 ;
        RECT 3.060 1.030 3.400 1.080 ;
        RECT 3.060 0.970 3.550 1.030 ;
        RECT 3.880 0.990 4.200 1.020 ;
        RECT 3.060 0.940 3.570 0.970 ;
        RECT 3.100 0.910 3.570 0.940 ;
        RECT 3.230 0.860 3.570 0.910 ;
        RECT 3.350 0.850 3.570 0.860 ;
        RECT 3.360 0.820 3.570 0.850 ;
        RECT 3.380 0.740 3.570 0.820 ;
        RECT 3.880 0.800 4.210 0.990 ;
        RECT 4.340 0.960 4.640 1.100 ;
        RECT 7.510 1.090 7.680 1.460 ;
        RECT 8.230 1.380 8.400 1.410 ;
        RECT 8.230 1.350 8.630 1.380 ;
        RECT 8.230 1.160 8.640 1.350 ;
        RECT 8.890 1.310 9.180 1.360 ;
        RECT 8.840 1.190 9.180 1.310 ;
        RECT 8.230 1.120 8.630 1.160 ;
        RECT 8.230 1.110 8.400 1.120 ;
        RECT 7.510 1.080 7.800 1.090 ;
        RECT 8.840 1.080 9.030 1.190 ;
        RECT 4.450 0.870 4.640 0.960 ;
        RECT 3.880 0.760 4.200 0.800 ;
        RECT 4.740 0.740 5.070 0.860 ;
        RECT 5.900 0.850 6.090 1.080 ;
        RECT 6.800 0.990 7.120 1.020 ;
        RECT 6.800 0.800 7.130 0.990 ;
        RECT 7.610 0.860 7.800 1.080 ;
        RECT 6.800 0.760 7.120 0.800 ;
        RECT 9.460 0.770 9.630 1.450 ;
        RECT 3.380 0.690 3.900 0.740 ;
        RECT 3.480 0.570 3.900 0.690 ;
        RECT 3.480 0.460 3.670 0.570 ;
        RECT 4.250 0.560 8.470 0.740 ;
        RECT 8.850 0.560 9.200 0.730 ;
        RECT 9.380 0.690 9.630 0.770 ;
        RECT 9.300 0.570 9.630 0.690 ;
        RECT 9.300 0.460 9.490 0.570 ;
        RECT 2.980 0.430 3.150 0.450 ;
        RECT 2.960 0.000 3.170 0.430 ;
      LAYER mcon ;
        RECT 3.490 6.290 3.660 6.460 ;
        RECT 9.310 6.290 9.480 6.460 ;
        RECT 3.940 5.970 4.110 6.140 ;
        RECT 4.460 5.880 4.630 6.050 ;
        RECT 5.910 5.900 6.080 6.070 ;
        RECT 6.860 5.970 7.030 6.140 ;
        RECT 7.620 5.890 7.790 6.060 ;
        RECT 5.290 5.600 5.460 5.770 ;
        RECT 8.370 5.610 8.540 5.780 ;
        RECT 8.850 5.670 9.020 5.840 ;
        RECT 5.290 4.200 5.460 4.370 ;
        RECT 8.370 4.190 8.540 4.360 ;
        RECT 8.850 4.130 9.020 4.300 ;
        RECT 3.940 3.830 4.110 4.000 ;
        RECT 4.460 3.920 4.630 4.090 ;
        RECT 5.910 3.900 6.080 4.070 ;
        RECT 6.860 3.830 7.030 4.000 ;
        RECT 7.620 3.910 7.790 4.080 ;
        RECT 3.490 3.510 3.660 3.680 ;
        RECT 9.310 3.510 9.480 3.680 ;
        RECT 2.980 3.300 3.150 3.470 ;
        RECT 3.490 3.270 3.660 3.440 ;
        RECT 9.310 3.270 9.480 3.440 ;
        RECT 3.940 2.950 4.110 3.120 ;
        RECT 4.460 2.860 4.630 3.030 ;
        RECT 5.910 2.880 6.080 3.050 ;
        RECT 6.860 2.950 7.030 3.120 ;
        RECT 7.620 2.870 7.790 3.040 ;
        RECT 5.290 2.580 5.460 2.750 ;
        RECT 8.370 2.590 8.540 2.760 ;
        RECT 8.850 2.650 9.020 2.820 ;
        RECT 5.290 1.180 5.460 1.350 ;
        RECT 8.370 1.170 8.540 1.340 ;
        RECT 8.850 1.110 9.020 1.280 ;
        RECT 3.940 0.810 4.110 0.980 ;
        RECT 4.460 0.900 4.630 1.070 ;
        RECT 5.910 0.880 6.080 1.050 ;
        RECT 6.860 0.810 7.030 0.980 ;
        RECT 7.620 0.890 7.790 1.060 ;
        RECT 3.490 0.490 3.660 0.660 ;
        RECT 9.310 0.490 9.480 0.660 ;
        RECT 2.980 0.280 3.150 0.450 ;
      LAYER met1 ;
        RECT 2.960 6.790 3.180 6.950 ;
        RECT 2.960 6.730 3.300 6.790 ;
        RECT 2.950 6.470 3.300 6.730 ;
        RECT 3.370 6.520 3.570 6.800 ;
        RECT 2.950 6.440 3.180 6.470 ;
        RECT 3.370 6.230 3.690 6.520 ;
        RECT 4.430 6.390 4.690 6.710 ;
        RECT 5.850 6.400 6.110 6.720 ;
        RECT 7.600 6.420 7.860 6.740 ;
        RECT 8.640 6.560 8.900 6.730 ;
        RECT 8.640 6.410 8.910 6.560 ;
        RECT 3.370 5.280 3.570 6.230 ;
        RECT 3.870 5.900 4.190 6.220 ;
        RECT 4.350 6.110 4.520 6.290 ;
        RECT 5.800 6.130 5.970 6.310 ;
        RECT 4.350 6.020 4.660 6.110 ;
        RECT 5.800 6.040 6.110 6.130 ;
        RECT 4.430 5.820 4.660 6.020 ;
        RECT 5.220 5.530 5.540 5.850 ;
        RECT 5.880 5.840 6.110 6.040 ;
        RECT 6.790 5.900 7.110 6.220 ;
        RECT 7.520 6.120 7.690 6.350 ;
        RECT 7.520 6.010 7.820 6.120 ;
        RECT 7.590 5.830 7.820 6.010 ;
        RECT 8.720 5.900 8.910 6.410 ;
        RECT 9.200 6.520 9.390 6.800 ;
        RECT 9.200 6.230 9.510 6.520 ;
        RECT 8.300 5.540 8.620 5.860 ;
        RECT 8.720 5.810 9.050 5.900 ;
        RECT 8.820 5.610 9.050 5.810 ;
        RECT 9.200 5.280 9.390 6.230 ;
        RECT 2.960 3.770 3.180 3.930 ;
        RECT 2.960 3.710 3.300 3.770 ;
        RECT 2.950 3.240 3.300 3.710 ;
        RECT 2.960 3.180 3.300 3.240 ;
        RECT 3.370 3.740 3.570 4.690 ;
        RECT 3.870 3.750 4.190 4.070 ;
        RECT 4.430 3.950 4.660 4.150 ;
        RECT 5.220 4.120 5.540 4.440 ;
        RECT 4.350 3.860 4.660 3.950 ;
        RECT 5.880 3.930 6.110 4.130 ;
        RECT 3.370 3.210 3.690 3.740 ;
        RECT 4.350 3.690 4.520 3.860 ;
        RECT 5.800 3.840 6.110 3.930 ;
        RECT 5.800 3.700 5.970 3.840 ;
        RECT 6.790 3.750 7.110 4.070 ;
        RECT 7.590 3.960 7.820 4.140 ;
        RECT 8.300 4.110 8.620 4.430 ;
        RECT 8.820 4.160 9.050 4.360 ;
        RECT 7.520 3.850 7.820 3.960 ;
        RECT 8.720 4.070 9.050 4.160 ;
        RECT 7.520 3.720 7.690 3.850 ;
        RECT 4.350 3.680 4.690 3.690 ;
        RECT 4.430 3.270 4.690 3.680 ;
        RECT 5.800 3.660 6.110 3.700 ;
        RECT 5.850 3.290 6.110 3.660 ;
        RECT 7.520 3.620 7.860 3.720 ;
        RECT 8.720 3.710 8.910 4.070 ;
        RECT 7.600 3.330 7.860 3.620 ;
        RECT 4.350 3.260 4.690 3.270 ;
        RECT 2.960 3.020 3.180 3.180 ;
        RECT 3.370 2.260 3.570 3.210 ;
        RECT 3.870 2.880 4.190 3.200 ;
        RECT 4.350 3.090 4.520 3.260 ;
        RECT 5.800 3.250 6.110 3.290 ;
        RECT 5.800 3.110 5.970 3.250 ;
        RECT 7.520 3.230 7.860 3.330 ;
        RECT 8.640 3.240 8.910 3.710 ;
        RECT 4.350 3.000 4.660 3.090 ;
        RECT 5.800 3.020 6.110 3.110 ;
        RECT 4.430 2.800 4.660 3.000 ;
        RECT 5.220 2.510 5.540 2.830 ;
        RECT 5.880 2.820 6.110 3.020 ;
        RECT 6.790 2.880 7.110 3.200 ;
        RECT 7.520 3.100 7.690 3.230 ;
        RECT 7.520 2.990 7.820 3.100 ;
        RECT 7.590 2.810 7.820 2.990 ;
        RECT 8.720 2.880 8.910 3.240 ;
        RECT 9.200 3.740 9.390 4.690 ;
        RECT 9.200 3.210 9.510 3.740 ;
        RECT 8.300 2.520 8.620 2.840 ;
        RECT 8.720 2.790 9.050 2.880 ;
        RECT 8.820 2.590 9.050 2.790 ;
        RECT 9.200 2.260 9.390 3.210 ;
        RECT 3.370 0.720 3.570 1.670 ;
        RECT 3.870 0.730 4.190 1.050 ;
        RECT 4.430 0.930 4.660 1.130 ;
        RECT 5.220 1.100 5.540 1.420 ;
        RECT 4.350 0.840 4.660 0.930 ;
        RECT 5.880 0.910 6.110 1.110 ;
        RECT 2.950 0.480 3.180 0.510 ;
        RECT 2.950 0.220 3.300 0.480 ;
        RECT 2.960 0.160 3.300 0.220 ;
        RECT 3.370 0.430 3.690 0.720 ;
        RECT 4.350 0.660 4.520 0.840 ;
        RECT 5.800 0.820 6.110 0.910 ;
        RECT 5.800 0.640 5.970 0.820 ;
        RECT 6.790 0.730 7.110 1.050 ;
        RECT 7.590 0.940 7.820 1.120 ;
        RECT 8.300 1.090 8.620 1.410 ;
        RECT 8.820 1.140 9.050 1.340 ;
        RECT 7.520 0.830 7.820 0.940 ;
        RECT 8.720 1.050 9.050 1.140 ;
        RECT 7.520 0.600 7.690 0.830 ;
        RECT 2.960 0.000 3.180 0.160 ;
        RECT 3.370 0.150 3.570 0.430 ;
        RECT 4.430 0.240 4.690 0.560 ;
        RECT 5.850 0.230 6.110 0.550 ;
        RECT 8.720 0.540 8.910 1.050 ;
        RECT 7.600 0.210 7.860 0.530 ;
        RECT 8.640 0.390 8.910 0.540 ;
        RECT 9.200 0.720 9.390 1.670 ;
        RECT 9.200 0.430 9.510 0.720 ;
        RECT 8.640 0.220 8.900 0.390 ;
        RECT 9.200 0.150 9.390 0.430 ;
      LAYER via ;
        RECT 3.040 6.500 3.300 6.760 ;
        RECT 4.430 6.420 4.690 6.680 ;
        RECT 5.850 6.430 6.110 6.690 ;
        RECT 7.600 6.450 7.860 6.710 ;
        RECT 8.640 6.440 8.900 6.700 ;
        RECT 3.900 5.930 4.160 6.190 ;
        RECT 6.820 5.930 7.080 6.190 ;
        RECT 5.250 5.560 5.510 5.820 ;
        RECT 8.330 5.570 8.590 5.830 ;
        RECT 3.040 3.480 3.300 3.740 ;
        RECT 3.040 3.210 3.300 3.470 ;
        RECT 5.250 4.150 5.510 4.410 ;
        RECT 3.900 3.780 4.160 4.040 ;
        RECT 8.330 4.140 8.590 4.400 ;
        RECT 6.820 3.780 7.080 4.040 ;
        RECT 4.430 3.290 4.690 3.660 ;
        RECT 5.850 3.280 6.110 3.670 ;
        RECT 3.900 2.910 4.160 3.170 ;
        RECT 7.600 3.260 7.860 3.690 ;
        RECT 8.640 3.270 8.900 3.680 ;
        RECT 6.820 2.910 7.080 3.170 ;
        RECT 5.250 2.540 5.510 2.800 ;
        RECT 8.330 2.550 8.590 2.810 ;
        RECT 5.250 1.130 5.510 1.390 ;
        RECT 3.900 0.760 4.160 1.020 ;
        RECT 8.330 1.120 8.590 1.380 ;
        RECT 3.040 0.190 3.300 0.450 ;
        RECT 6.820 0.760 7.080 1.020 ;
        RECT 4.430 0.270 4.690 0.530 ;
        RECT 5.850 0.260 6.110 0.520 ;
        RECT 7.600 0.240 7.860 0.500 ;
        RECT 8.640 0.250 8.900 0.510 ;
      LAYER met2 ;
        RECT 3.010 6.570 3.330 6.760 ;
        RECT 4.400 6.570 4.720 6.680 ;
        RECT 5.820 6.570 6.140 6.690 ;
        RECT 7.570 6.570 7.890 6.710 ;
        RECT 8.610 6.570 8.930 6.700 ;
        RECT 2.630 6.500 3.330 6.570 ;
        RECT 2.630 6.370 3.240 6.500 ;
        RECT 4.330 6.370 9.710 6.570 ;
        RECT 3.870 6.070 4.180 6.230 ;
        RECT 6.790 6.070 7.100 6.230 ;
        RECT 2.630 5.900 7.100 6.070 ;
        RECT 2.630 5.870 7.000 5.900 ;
        RECT 2.630 4.070 7.000 4.100 ;
        RECT 2.630 3.900 7.100 4.070 ;
        RECT 3.870 3.740 4.180 3.900 ;
        RECT 6.790 3.740 7.100 3.900 ;
        RECT 3.010 3.600 3.330 3.740 ;
        RECT 4.400 3.600 4.720 3.660 ;
        RECT 5.820 3.600 6.140 3.670 ;
        RECT 7.570 3.600 7.890 3.690 ;
        RECT 8.610 3.600 8.930 3.680 ;
        RECT 2.630 3.480 3.330 3.600 ;
        RECT 2.630 3.470 3.240 3.480 ;
        RECT 2.630 3.350 3.330 3.470 ;
        RECT 4.330 3.350 9.710 3.600 ;
        RECT 3.010 3.210 3.330 3.350 ;
        RECT 4.400 3.290 4.720 3.350 ;
        RECT 5.820 3.280 6.140 3.350 ;
        RECT 7.570 3.260 7.890 3.350 ;
        RECT 8.610 3.270 8.930 3.350 ;
        RECT 3.870 3.050 4.180 3.210 ;
        RECT 6.790 3.050 7.100 3.210 ;
        RECT 2.630 2.880 7.100 3.050 ;
        RECT 2.630 2.850 7.000 2.880 ;
        RECT 2.630 1.050 7.000 1.080 ;
        RECT 2.630 0.880 7.100 1.050 ;
        RECT 3.870 0.720 4.180 0.880 ;
        RECT 6.790 0.720 7.100 0.880 ;
        RECT 2.630 0.450 3.240 0.580 ;
        RECT 2.630 0.380 3.330 0.450 ;
        RECT 4.330 0.380 9.710 0.580 ;
        RECT 3.010 0.190 3.330 0.380 ;
        RECT 4.400 0.270 4.720 0.380 ;
        RECT 5.820 0.260 6.140 0.380 ;
        RECT 7.570 0.240 7.890 0.380 ;
        RECT 8.610 0.250 8.930 0.380 ;
  END
END sky130_hilas_Tgate4Double01

MACRO sky130_hilas_cellAttempt01
  CLASS CORE ;
  FOREIGN sky130_hilas_cellAttempt01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.240 BY 10.900 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 0.350 0.410 0.750 6.910 ;
    END
  END VTUN
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 9.550 6.630 9.710 6.680 ;
    END
  END VINJ
  PIN COLSEL1
    PORT
      LAYER met1 ;
        RECT 9.110 6.630 9.300 6.680 ;
    END
  END COLSEL1
  PIN COL1
    PORT
      LAYER met1 ;
        RECT 8.740 6.640 8.900 6.680 ;
    END
  END COL1
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT 4.400 6.580 4.780 6.910 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.400 0.410 4.780 1.010 ;
    END
  END GATE1
  PIN ROW4
    PORT
      LAYER met2 ;
        RECT 0.000 1.400 7.620 1.580 ;
    END
  END ROW4
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 2.750 2.190 3.070 2.200 ;
        RECT 6.680 2.190 7.000 2.250 ;
        RECT 2.750 2.010 7.000 2.190 ;
        RECT 2.750 1.940 3.070 2.010 ;
        RECT 6.680 1.960 7.000 2.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.720 5.520 6.960 6.910 ;
        RECT 6.700 4.860 6.970 5.520 ;
        RECT 6.720 2.270 6.960 4.860 ;
        RECT 6.710 1.950 6.970 2.270 ;
        RECT 6.720 0.410 6.960 1.950 ;
      LAYER via ;
        RECT 6.710 1.980 6.970 2.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.790 5.500 3.030 6.910 ;
        RECT 2.780 4.840 3.040 5.500 ;
        RECT 2.790 2.230 3.030 4.840 ;
        RECT 2.780 1.910 3.040 2.230 ;
        RECT 2.790 0.410 3.030 1.910 ;
      LAYER via ;
        RECT 2.780 1.940 3.040 2.200 ;
    END
  END VGND
  PIN DRAIN4
    PORT
      LAYER met2 ;
        RECT 0.000 0.980 7.600 1.150 ;
    END
  END DRAIN4
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 0.000 6.170 7.630 6.350 ;
    END
  END DRAIN1
  PIN ROW1
    PORT
      LAYER met2 ;
        RECT 0.000 5.730 7.630 5.910 ;
    END
  END ROW1
  PIN ROW3
    PORT
      LAYER met2 ;
        RECT 0.000 2.500 7.630 2.680 ;
    END
  END ROW3
  PIN DRAIN3
    PORT
      LAYER met2 ;
        RECT 0.000 2.930 7.620 3.110 ;
    END
  END DRAIN3
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 0.000 4.200 7.630 4.380 ;
    END
  END DRAIN2
  PIN ROW2
    PORT
      LAYER met2 ;
        RECT 0.000 4.630 7.630 4.810 ;
    END
  END ROW2
  OBS
      LAYER nwell ;
        RECT 14.510 10.850 16.240 10.900 ;
        RECT 0.000 5.570 0.070 5.750 ;
        RECT 10.400 5.410 12.960 7.320 ;
        RECT 0.570 5.220 1.160 5.330 ;
        RECT 4.310 5.160 5.420 5.390 ;
        RECT 8.950 3.730 9.300 3.740 ;
        RECT 8.950 3.570 9.120 3.730 ;
        RECT 9.290 3.570 9.300 3.730 ;
        RECT 0.570 1.940 1.160 2.130 ;
        RECT 4.310 1.920 5.420 2.190 ;
        RECT 10.400 2.170 12.960 5.140 ;
        RECT 13.320 4.410 16.240 10.850 ;
        RECT 18.510 7.320 20.240 9.160 ;
        RECT 13.320 4.360 15.550 4.410 ;
        RECT 10.400 0.000 12.960 1.910 ;
      LAYER li1 ;
        RECT 14.900 7.840 15.450 8.270 ;
        RECT 18.930 7.770 19.480 8.200 ;
        RECT 10.640 6.970 10.960 7.010 ;
        RECT 10.640 6.850 10.970 6.970 ;
        RECT 10.640 6.750 11.080 6.850 ;
        RECT 10.740 6.680 11.080 6.750 ;
        RECT 12.360 6.580 12.560 6.930 ;
        RECT 10.640 6.420 10.960 6.460 ;
        RECT 10.640 6.230 10.970 6.420 ;
        RECT 10.640 6.200 11.080 6.230 ;
        RECT 10.740 6.060 11.080 6.200 ;
        RECT 11.630 5.960 11.830 6.560 ;
        RECT 12.360 6.550 12.570 6.580 ;
        RECT 12.350 5.960 12.570 6.550 ;
        RECT 2.820 4.930 2.990 5.460 ;
        RECT 6.760 4.920 6.930 5.450 ;
        RECT 10.740 4.350 11.080 4.490 ;
        RECT 10.640 4.320 11.080 4.350 ;
        RECT 2.830 3.220 3.000 4.230 ;
        RECT 10.640 4.130 10.970 4.320 ;
        RECT 10.640 4.090 10.960 4.130 ;
        RECT 6.760 3.080 6.930 4.090 ;
        RECT 11.630 3.990 11.830 4.590 ;
        RECT 12.350 4.000 12.570 4.590 ;
        RECT 12.360 3.970 12.570 4.000 ;
        RECT 10.740 3.800 11.080 3.870 ;
        RECT 8.860 3.570 9.300 3.740 ;
        RECT 10.640 3.700 11.080 3.800 ;
        RECT 10.640 3.610 10.970 3.700 ;
        RECT 10.640 3.510 11.080 3.610 ;
        RECT 10.740 3.440 11.080 3.510 ;
        RECT 12.360 3.340 12.560 3.970 ;
        RECT 10.640 3.180 10.960 3.220 ;
        RECT 10.640 2.990 10.970 3.180 ;
        RECT 10.640 2.960 11.080 2.990 ;
        RECT 10.740 2.820 11.080 2.960 ;
        RECT 11.630 2.720 11.830 3.320 ;
        RECT 12.360 3.310 12.570 3.340 ;
        RECT 12.350 2.720 12.570 3.310 ;
        RECT 10.740 1.120 11.080 1.260 ;
        RECT 10.640 1.090 11.080 1.120 ;
        RECT 10.640 0.900 10.970 1.090 ;
        RECT 10.640 0.860 10.960 0.900 ;
        RECT 11.630 0.760 11.830 1.360 ;
        RECT 12.350 0.770 12.570 1.360 ;
        RECT 12.360 0.740 12.570 0.770 ;
        RECT 10.740 0.570 11.080 0.640 ;
        RECT 10.640 0.470 11.080 0.570 ;
        RECT 10.640 0.350 10.970 0.470 ;
        RECT 12.360 0.390 12.560 0.740 ;
        RECT 10.640 0.310 10.960 0.350 ;
      LAYER mcon ;
        RECT 14.900 7.920 15.170 8.190 ;
        RECT 18.930 7.850 19.200 8.120 ;
        RECT 10.700 6.790 10.870 6.960 ;
        RECT 10.700 6.240 10.870 6.410 ;
        RECT 11.640 6.350 11.810 6.520 ;
        RECT 12.370 6.380 12.540 6.550 ;
        RECT 2.820 5.290 2.990 5.460 ;
        RECT 6.760 5.280 6.930 5.450 ;
        RECT 10.700 4.140 10.870 4.310 ;
        RECT 2.830 3.830 3.000 4.000 ;
        RECT 2.830 3.470 3.000 3.640 ;
        RECT 11.640 4.030 11.810 4.200 ;
        RECT 12.370 4.000 12.540 4.170 ;
        RECT 6.760 3.690 6.930 3.860 ;
        RECT 9.120 3.570 9.300 3.740 ;
        RECT 10.700 3.550 10.870 3.760 ;
        RECT 6.760 3.330 6.930 3.500 ;
        RECT 10.700 3.000 10.870 3.170 ;
        RECT 11.640 3.110 11.810 3.280 ;
        RECT 12.370 3.140 12.540 3.310 ;
        RECT 10.700 0.910 10.870 1.080 ;
        RECT 11.640 0.800 11.810 0.970 ;
        RECT 12.370 0.770 12.540 0.940 ;
        RECT 10.700 0.360 10.870 0.530 ;
      LAYER met1 ;
        RECT 10.630 6.720 10.950 7.040 ;
        RECT 11.630 6.580 11.790 7.310 ;
        RECT 11.630 6.560 11.830 6.580 ;
        RECT 10.630 6.170 10.950 6.490 ;
        RECT 11.610 6.320 11.840 6.560 ;
        RECT 11.630 6.270 11.840 6.320 ;
        RECT 12.000 6.270 12.190 7.260 ;
        RECT 12.440 6.610 12.600 7.310 ;
        RECT 11.630 5.410 11.790 6.270 ;
        RECT 12.020 6.150 12.190 6.270 ;
        RECT 12.030 5.410 12.190 6.150 ;
        RECT 12.330 6.060 12.600 6.610 ;
        RECT 12.330 6.010 12.610 6.060 ;
        RECT 12.440 5.920 12.610 6.010 ;
        RECT 12.440 5.410 12.600 5.920 ;
        RECT 10.630 4.060 10.950 4.380 ;
        RECT 11.630 4.280 11.790 5.140 ;
        RECT 12.030 4.400 12.190 5.140 ;
        RECT 12.440 4.630 12.600 5.140 ;
        RECT 12.440 4.540 12.610 4.630 ;
        RECT 12.020 4.280 12.190 4.400 ;
        RECT 11.630 4.230 11.840 4.280 ;
        RECT 11.610 3.990 11.840 4.230 ;
        RECT 11.630 3.970 11.830 3.990 ;
        RECT 9.170 3.770 9.300 3.790 ;
        RECT 9.090 3.750 9.330 3.770 ;
        RECT 8.890 3.560 9.330 3.750 ;
        RECT 9.090 3.540 9.330 3.560 ;
        RECT 9.190 3.500 9.300 3.540 ;
        RECT 10.630 3.480 10.950 3.830 ;
        RECT 11.630 3.340 11.790 3.970 ;
        RECT 11.630 3.320 11.830 3.340 ;
        RECT 10.630 2.930 10.950 3.250 ;
        RECT 11.610 3.080 11.840 3.320 ;
        RECT 11.630 3.030 11.840 3.080 ;
        RECT 12.000 3.030 12.190 4.280 ;
        RECT 12.330 4.490 12.610 4.540 ;
        RECT 12.330 3.940 12.600 4.490 ;
        RECT 13.970 4.360 14.350 10.860 ;
        RECT 14.840 7.380 15.230 9.240 ;
        RECT 18.870 7.310 19.260 9.170 ;
        RECT 12.440 3.370 12.600 3.940 ;
        RECT 11.630 2.170 11.790 3.030 ;
        RECT 12.020 2.910 12.190 3.030 ;
        RECT 12.030 2.170 12.190 2.910 ;
        RECT 12.330 2.820 12.600 3.370 ;
        RECT 12.330 2.770 12.610 2.820 ;
        RECT 12.440 2.680 12.610 2.770 ;
        RECT 12.440 2.170 12.600 2.680 ;
        RECT 10.630 0.830 10.950 1.150 ;
        RECT 11.630 1.050 11.790 1.910 ;
        RECT 12.030 1.170 12.190 1.910 ;
        RECT 12.440 1.400 12.600 1.910 ;
        RECT 12.440 1.310 12.610 1.400 ;
        RECT 12.020 1.050 12.190 1.170 ;
        RECT 11.630 1.000 11.840 1.050 ;
        RECT 11.610 0.760 11.840 1.000 ;
        RECT 11.630 0.740 11.830 0.760 ;
        RECT 10.630 0.280 10.950 0.600 ;
        RECT 11.630 0.010 11.790 0.740 ;
        RECT 12.000 0.060 12.190 1.050 ;
        RECT 12.330 1.260 12.610 1.310 ;
        RECT 12.330 0.710 12.600 1.260 ;
        RECT 12.440 0.010 12.600 0.710 ;
      LAYER via ;
        RECT 10.660 6.750 10.920 7.010 ;
        RECT 10.660 6.200 10.920 6.460 ;
        RECT 10.660 4.090 10.920 4.350 ;
        RECT 10.660 3.510 10.920 3.800 ;
        RECT 10.660 2.960 10.920 3.220 ;
        RECT 10.660 0.860 10.920 1.120 ;
        RECT 10.660 0.310 10.920 0.570 ;
      LAYER met2 ;
        RECT 10.630 6.760 10.940 7.050 ;
        RECT 10.630 6.720 12.960 6.760 ;
        RECT 10.780 6.580 12.960 6.720 ;
        RECT 10.630 6.330 10.940 6.500 ;
        RECT 10.400 6.150 10.490 6.330 ;
        RECT 10.630 6.170 12.960 6.330 ;
        RECT 10.790 6.150 12.960 6.170 ;
        RECT 10.400 4.220 10.490 4.400 ;
        RECT 10.790 4.380 12.960 4.400 ;
        RECT 10.630 4.220 12.960 4.380 ;
        RECT 10.630 4.050 10.940 4.220 ;
        RECT 10.780 3.830 12.960 3.970 ;
        RECT 10.630 3.790 12.960 3.830 ;
        RECT 10.630 3.520 10.940 3.790 ;
        RECT 10.630 3.480 12.960 3.520 ;
        RECT 10.780 3.340 12.960 3.480 ;
        RECT 10.630 3.090 10.940 3.260 ;
        RECT 10.400 2.910 10.490 3.090 ;
        RECT 10.630 2.930 12.960 3.090 ;
        RECT 10.790 2.910 12.960 2.930 ;
        RECT 10.400 0.990 10.490 1.170 ;
        RECT 10.790 1.150 12.960 1.170 ;
        RECT 10.630 0.990 12.960 1.150 ;
        RECT 10.630 0.820 10.940 0.990 ;
        RECT 10.780 0.600 12.960 0.740 ;
        RECT 10.630 0.560 12.960 0.600 ;
        RECT 10.630 0.270 10.940 0.560 ;
  END
END sky130_hilas_cellAttempt01

MACRO sky130_hilas_StepUpDigital
  CLASS CORE ;
  FOREIGN sky130_hilas_StepUpDigital ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.360 BY 2.180 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 0.220 0.000 2.720 1.750 ;
        RECT 3.810 0.580 5.580 2.170 ;
        RECT 6.590 1.680 8.360 1.750 ;
        RECT 6.590 0.000 8.360 0.090 ;
      LAYER li1 ;
        RECT 0.160 1.750 0.330 1.790 ;
        RECT 0.160 1.730 1.310 1.750 ;
        RECT 0.160 1.560 1.350 1.730 ;
        RECT 1.800 1.700 2.260 1.730 ;
        RECT 3.570 1.700 3.920 1.800 ;
        RECT 1.800 1.560 2.910 1.700 ;
        RECT 2.090 1.530 2.910 1.560 ;
        RECT 3.150 1.530 4.320 1.700 ;
        RECT 4.570 1.530 5.330 1.700 ;
        RECT 2.090 1.390 2.350 1.530 ;
        RECT 0.560 1.060 0.890 1.230 ;
        RECT 1.170 1.220 2.350 1.390 ;
        RECT 5.100 1.520 5.330 1.530 ;
        RECT 1.170 1.070 1.950 1.220 ;
        RECT 2.090 1.080 2.350 1.220 ;
        RECT 2.650 1.290 2.940 1.320 ;
        RECT 2.650 1.120 2.980 1.290 ;
        RECT 2.650 1.080 2.940 1.120 ;
        RECT 3.560 1.080 3.890 1.340 ;
        RECT 5.100 1.080 5.370 1.520 ;
        RECT 0.000 0.880 0.620 1.050 ;
        RECT 0.630 0.600 0.810 1.060 ;
        RECT 1.170 0.780 1.350 1.070 ;
        RECT 1.590 0.720 1.800 1.050 ;
        RECT 2.090 0.910 2.420 1.080 ;
        RECT 2.660 0.910 4.820 1.080 ;
        RECT 2.090 0.860 2.320 0.910 ;
        RECT 5.070 0.900 5.400 1.080 ;
        RECT 5.750 0.940 5.920 1.000 ;
        RECT 2.150 0.630 2.320 0.860 ;
        RECT 5.730 0.720 5.950 0.940 ;
        RECT 5.750 0.670 5.920 0.720 ;
        RECT 2.150 0.620 2.530 0.630 ;
        RECT 0.630 0.430 1.590 0.600 ;
        RECT 2.060 0.560 2.530 0.620 ;
        RECT 2.060 0.510 2.870 0.560 ;
        RECT 2.060 0.450 2.880 0.510 ;
        RECT 2.140 0.390 2.880 0.450 ;
        RECT 2.140 0.340 2.530 0.390 ;
      LAYER mcon ;
        RECT 3.630 1.570 3.840 1.780 ;
        RECT 1.670 1.140 1.840 1.310 ;
        RECT 2.710 1.100 2.880 1.270 ;
        RECT 5.140 1.200 5.310 1.370 ;
        RECT 0.630 0.800 0.800 0.970 ;
        RECT 0.630 0.440 0.800 0.610 ;
      LAYER met1 ;
        RECT 0.560 0.000 0.850 1.750 ;
        RECT 1.600 1.110 1.920 1.390 ;
        RECT 1.560 1.090 1.920 1.110 ;
        RECT 1.560 0.780 1.840 1.090 ;
        RECT 2.090 0.490 2.400 2.180 ;
        RECT 3.570 1.530 3.920 1.820 ;
        RECT 5.100 1.750 5.340 2.170 ;
        RECT 4.870 1.690 5.340 1.750 ;
        RECT 3.720 1.510 3.920 1.530 ;
        RECT 2.650 1.320 2.960 1.330 ;
        RECT 2.640 1.050 2.960 1.320 ;
        RECT 2.650 1.040 2.940 1.050 ;
        RECT 5.100 0.490 5.340 1.690 ;
        RECT 7.880 1.680 8.120 1.750 ;
        RECT 5.670 0.670 6.080 1.000 ;
      LAYER via ;
        RECT 1.630 1.100 1.890 1.360 ;
        RECT 1.570 0.820 1.830 1.080 ;
        RECT 3.610 1.540 3.870 1.800 ;
        RECT 2.670 1.060 2.930 1.320 ;
        RECT 5.710 0.700 5.970 0.960 ;
      LAYER met2 ;
        RECT 1.600 1.310 1.920 1.360 ;
        RECT 2.630 1.320 2.950 1.330 ;
        RECT 2.630 1.310 2.960 1.320 ;
        RECT 0.290 1.110 2.960 1.310 ;
        RECT 1.600 1.100 1.920 1.110 ;
        RECT 1.530 1.030 1.870 1.090 ;
        RECT 2.630 1.060 2.960 1.110 ;
        RECT 2.630 1.040 2.950 1.060 ;
        RECT 3.610 1.030 3.870 1.830 ;
        RECT 1.530 0.810 3.970 1.030 ;
        RECT 5.680 0.670 6.140 0.990 ;
  END
END sky130_hilas_StepUpDigital

MACRO sky130_hilas_VinjNOR3
  CLASS CORE ;
  FOREIGN sky130_hilas_VinjNOR3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.880 BY 1.640 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 0.010 0.000 3.450 1.640 ;
      LAYER li1 ;
        RECT 0.630 1.210 0.800 1.350 ;
        RECT 1.360 1.230 1.530 1.310 ;
        RECT 2.170 1.230 2.340 1.310 ;
        RECT 3.710 1.270 3.880 1.390 ;
        RECT 0.630 1.040 0.820 1.210 ;
        RECT 0.630 0.940 0.800 1.040 ;
        RECT 1.360 0.660 1.570 1.230 ;
        RECT 2.130 0.980 2.340 1.230 ;
        RECT 2.730 1.050 2.900 1.150 ;
        RECT 3.670 1.100 3.880 1.270 ;
        RECT 5.600 1.200 5.860 1.270 ;
        RECT 6.400 1.200 6.580 1.330 ;
        RECT 3.710 1.060 3.880 1.100 ;
        RECT 2.130 0.660 2.300 0.980 ;
        RECT 2.700 0.880 2.900 1.050 ;
        RECT 2.730 0.780 2.900 0.880 ;
        RECT 4.270 1.020 5.140 1.190 ;
        RECT 5.600 1.020 6.580 1.200 ;
        RECT 0.200 0.560 0.370 0.660 ;
        RECT 0.180 0.390 0.370 0.560 ;
        RECT 0.200 0.330 0.370 0.390 ;
        RECT 0.620 0.600 0.790 0.660 ;
        RECT 0.620 0.330 0.870 0.600 ;
        RECT 1.360 0.410 1.610 0.660 ;
        RECT 0.630 0.310 0.870 0.330 ;
        RECT 1.440 0.320 1.610 0.410 ;
        RECT 2.090 0.410 2.300 0.660 ;
        RECT 4.270 0.580 4.440 1.020 ;
        RECT 5.600 0.580 5.860 1.020 ;
        RECT 6.400 0.910 6.580 1.020 ;
        RECT 2.810 0.410 4.440 0.580 ;
        RECT 4.890 0.410 5.860 0.580 ;
        RECT 6.310 0.410 6.650 0.580 ;
        RECT 2.090 0.330 2.260 0.410 ;
        RECT 3.580 0.370 3.750 0.410 ;
      LAYER mcon ;
        RECT 0.650 1.040 0.820 1.210 ;
        RECT 0.660 0.360 0.830 0.530 ;
        RECT 5.630 0.700 5.810 0.880 ;
      LAYER met1 ;
        RECT 0.620 1.260 0.840 1.600 ;
        RECT 0.620 1.000 0.850 1.260 ;
        RECT 0.090 0.320 0.400 0.670 ;
        RECT 0.620 0.600 0.840 1.000 ;
        RECT 2.640 0.840 2.970 1.100 ;
        RECT 3.610 1.060 4.040 1.350 ;
        RECT 0.620 0.290 0.870 0.600 ;
        RECT 3.480 0.310 3.870 0.580 ;
        RECT 0.620 0.090 0.840 0.290 ;
        RECT 5.590 0.090 5.860 1.610 ;
        RECT 6.410 0.320 6.720 0.640 ;
      LAYER via ;
        RECT 0.120 0.350 0.380 0.610 ;
        RECT 2.680 0.840 2.940 1.100 ;
        RECT 3.670 1.090 3.930 1.350 ;
        RECT 3.540 0.310 3.800 0.570 ;
        RECT 6.440 0.350 6.700 0.610 ;
      LAYER met2 ;
        RECT 0.000 1.290 4.040 1.450 ;
        RECT 2.640 1.020 2.970 1.100 ;
        RECT 3.620 1.060 4.040 1.290 ;
        RECT 2.370 1.000 2.970 1.020 ;
        RECT 0.010 0.840 2.970 1.000 ;
        RECT 0.090 0.510 0.410 0.610 ;
        RECT 0.010 0.350 0.410 0.510 ;
        RECT 3.500 0.490 3.870 0.570 ;
        RECT 3.500 0.480 4.530 0.490 ;
        RECT 6.410 0.480 6.720 0.640 ;
        RECT 3.500 0.310 6.880 0.480 ;
  END
END sky130_hilas_VinjNOR3

MACRO sky130_hilas_VinjDiodeProtect01
  CLASS CORE ;
  FOREIGN sky130_hilas_VinjDiodeProtect01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.590 BY 10.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN OUTPUT 
    ANTENNADIFFAREA 58.900799 ;
    PORT
      LAYER met1 ;
        RECT 14.350 10.250 14.700 10.410 ;
        RECT 14.340 9.300 14.710 10.250 ;
        RECT 13.990 8.930 16.460 9.300 ;
        RECT 12.550 7.470 16.460 8.930 ;
        RECT 2.840 7.460 16.460 7.470 ;
        RECT 2.170 6.900 16.460 7.460 ;
        RECT 2.170 2.600 25.520 6.900 ;
        RECT 2.170 2.320 16.460 2.600 ;
        RECT 12.550 0.770 16.460 2.320 ;
        RECT 12.530 0.000 16.480 0.770 ;
    END
  END OUTPUT 
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.000 7.380 28.590 8.780 ;
        RECT 0.470 7.370 1.400 7.380 ;
        RECT 0.720 6.260 0.890 7.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.440 8.130 2.810 8.760 ;
        RECT 23.780 8.280 27.910 8.680 ;
        RECT 23.780 8.190 27.920 8.280 ;
        RECT 0.470 6.170 1.420 8.130 ;
        RECT 2.170 8.110 2.750 8.130 ;
        RECT 27.390 7.290 27.920 8.190 ;
        RECT 0.700 0.500 1.420 6.170 ;
      LAYER via ;
        RECT 0.660 8.280 2.690 8.610 ;
        RECT 24.050 8.280 27.040 8.630 ;
        RECT 0.600 7.420 1.300 8.040 ;
        RECT 27.480 7.480 27.830 8.240 ;
    END
  END VGND
  PIN VINJ
    ANTENNADIFFAREA 9.088799 ;
    PORT
      LAYER nwell ;
        RECT 14.870 1.910 26.920 7.850 ;
      LAYER met2 ;
        RECT 26.340 2.480 26.980 5.490 ;
        RECT 0.000 1.080 28.590 2.480 ;
        RECT 25.440 0.950 28.070 1.080 ;
        RECT 25.440 0.440 27.990 0.950 ;
        RECT 25.440 0.370 26.060 0.440 ;
    END
  END VINJ
  PIN INPUT
    PORT
      LAYER met1 ;
        RECT 7.710 10.280 11.610 10.870 ;
        RECT 7.710 8.930 8.000 10.280 ;
    END
  END INPUT
  OBS
      LAYER li1 ;
        RECT 7.730 8.930 7.980 10.390 ;
        RECT 7.770 8.920 7.940 8.930 ;
        RECT 14.410 8.900 14.660 10.380 ;
        RECT 0.550 8.180 27.930 8.690 ;
        RECT 0.550 6.250 1.350 8.180 ;
        RECT 1.930 7.730 2.100 7.810 ;
        RECT 13.170 7.730 13.400 7.820 ;
        RECT 1.930 7.720 13.400 7.730 ;
        RECT 0.550 1.670 1.060 6.250 ;
        RECT 1.920 2.250 13.400 7.720 ;
        RECT 1.850 2.080 13.400 2.250 ;
        RECT 1.920 2.020 2.110 2.080 ;
        RECT 13.170 1.840 13.400 2.080 ;
        RECT 1.800 1.670 3.600 1.680 ;
        RECT 13.960 1.670 14.470 8.180 ;
        RECT 15.230 7.290 26.480 7.460 ;
        RECT 15.230 2.420 15.400 7.290 ;
        RECT 15.790 6.960 25.900 6.980 ;
        RECT 15.790 6.920 25.920 6.960 ;
        RECT 15.740 6.750 25.920 6.920 ;
        RECT 15.790 2.730 25.920 6.750 ;
        RECT 26.310 5.530 26.480 7.290 ;
        RECT 15.790 2.650 25.900 2.730 ;
        RECT 15.220 2.350 15.400 2.420 ;
        RECT 26.310 2.350 26.920 5.530 ;
        RECT 15.220 2.180 26.920 2.350 ;
        RECT 26.380 2.070 26.920 2.180 ;
        RECT 27.380 1.830 27.930 8.180 ;
        RECT 27.370 1.670 27.930 1.830 ;
        RECT 0.550 1.330 27.930 1.670 ;
        RECT 0.580 1.160 27.930 1.330 ;
        RECT 0.580 1.140 1.270 1.160 ;
        RECT 1.780 1.150 3.580 1.160 ;
      LAYER mcon ;
        RECT 7.770 9.870 7.940 10.040 ;
        RECT 7.770 9.510 7.940 9.680 ;
        RECT 7.770 9.140 7.940 9.310 ;
        RECT 14.450 10.190 14.620 10.360 ;
        RECT 14.450 9.830 14.620 10.000 ;
        RECT 14.450 9.470 14.620 9.640 ;
        RECT 14.450 9.110 14.620 9.280 ;
        RECT 0.630 8.520 2.490 8.530 ;
        RECT 0.630 8.350 2.500 8.520 ;
        RECT 23.990 8.340 27.150 8.520 ;
        RECT 0.670 6.260 0.850 8.160 ;
        RECT 1.070 6.250 1.250 8.160 ;
        RECT 2.260 7.220 13.240 7.390 ;
        RECT 2.260 6.600 13.240 6.770 ;
        RECT 2.270 5.980 13.250 6.150 ;
        RECT 2.290 5.400 13.270 5.570 ;
        RECT 2.300 4.810 13.280 4.980 ;
        RECT 2.300 4.210 13.280 4.380 ;
        RECT 2.250 3.610 13.230 3.780 ;
        RECT 2.260 3.000 13.240 3.170 ;
        RECT 2.250 2.400 13.230 2.570 ;
        RECT 15.990 6.460 25.440 6.630 ;
        RECT 15.980 5.710 25.370 5.880 ;
        RECT 16.010 4.990 25.410 5.160 ;
        RECT 16.020 4.330 25.390 4.500 ;
        RECT 16.010 3.680 25.460 3.850 ;
        RECT 16.020 3.040 25.410 3.210 ;
        RECT 27.560 7.360 27.760 8.290 ;
        RECT 26.490 2.120 26.840 5.420 ;
      LAYER met1 ;
        RECT 26.290 5.480 26.860 5.490 ;
        RECT 26.290 2.060 26.910 5.480 ;
        RECT 26.290 2.050 26.860 2.060 ;
        RECT 25.460 0.420 26.020 0.920 ;
        RECT 25.470 0.200 26.020 0.420 ;
      LAYER via ;
        RECT 26.450 2.190 26.870 5.360 ;
        RECT 25.480 0.370 26.000 0.890 ;
  END
END sky130_hilas_VinjDiodeProtect01

MACRO sky130_hilas_LevelShift4InputUp
  CLASS CORE ;
  FOREIGN sky130_hilas_LevelShift4InputUp ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.890 BY 7.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 7.850 6.950 8.090 7.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 7.850 0.000 8.090 0.050 ;
    END
  END VPWR
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 0.530 0.000 0.820 0.120 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.220 5.960 2.720 7.440 ;
        RECT 0.190 5.760 2.720 5.960 ;
        RECT 0.220 0.440 2.720 5.760 ;
      LAYER met1 ;
        RECT 0.560 7.000 0.850 7.440 ;
        RECT 0.530 6.910 0.850 7.000 ;
        RECT 0.560 0.440 0.850 6.910 ;
    END
  END VINJ
  PIN OUTPUT1
    PORT
      LAYER met2 ;
        RECT 0.190 6.360 0.350 6.560 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    PORT
      LAYER met2 ;
        RECT 0.190 4.610 0.360 4.810 ;
    END
  END OUTPUT2
  PIN OUTPUT3
    PORT
      LAYER met2 ;
        RECT 0.190 2.860 0.380 3.060 ;
    END
  END OUTPUT3
  PIN OUTPUT4
    PORT
      LAYER met2 ;
        RECT 0.190 1.110 0.350 1.310 ;
    END
  END OUTPUT4
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 4.840 0.000 5.150 0.060 ;
    END
    PORT
      LAYER nwell ;
        RECT 3.810 6.270 5.580 7.860 ;
      LAYER met1 ;
        RECT 5.100 7.440 5.340 7.860 ;
        RECT 4.870 7.380 5.340 7.440 ;
        RECT 5.100 7.000 5.340 7.380 ;
        RECT 4.840 6.940 5.340 7.000 ;
        RECT 5.100 6.180 5.340 6.940 ;
    END
  END VGND
  PIN INPUT1
    PORT
      LAYER met2 ;
        RECT 8.790 5.430 8.890 5.750 ;
    END
  END INPUT1
  PIN INPUT2
    PORT
      LAYER met2 ;
        RECT 8.790 3.680 8.890 4.000 ;
    END
  END INPUT2
  PIN INPUT3
    PORT
      LAYER met2 ;
        RECT 8.790 1.930 8.890 2.250 ;
    END
  END INPUT3
  PIN INPUT4
    PORT
      LAYER met2 ;
        RECT 8.790 0.180 8.890 0.500 ;
    END
  END INPUT4
  OBS
      LAYER nwell ;
        RECT 6.590 7.370 8.360 7.440 ;
        RECT 3.810 4.520 5.580 6.110 ;
        RECT 6.590 5.620 8.360 5.780 ;
        RECT 3.810 2.770 5.580 4.360 ;
        RECT 6.590 3.870 8.360 4.030 ;
        RECT 3.810 1.020 5.580 2.610 ;
        RECT 6.590 2.120 8.360 2.280 ;
        RECT 6.590 0.440 8.360 0.530 ;
      LAYER li1 ;
        RECT 0.160 7.440 0.330 7.480 ;
        RECT 0.160 7.420 1.310 7.440 ;
        RECT 0.160 7.250 1.350 7.420 ;
        RECT 1.800 7.390 2.260 7.420 ;
        RECT 3.570 7.390 3.920 7.490 ;
        RECT 1.800 7.250 2.910 7.390 ;
        RECT 2.090 7.220 2.910 7.250 ;
        RECT 3.150 7.220 4.320 7.390 ;
        RECT 4.570 7.220 5.330 7.390 ;
        RECT 2.090 7.080 2.350 7.220 ;
        RECT 0.560 6.750 0.890 6.920 ;
        RECT 1.170 6.910 2.350 7.080 ;
        RECT 5.100 7.210 5.330 7.220 ;
        RECT 1.170 6.760 1.950 6.910 ;
        RECT 2.090 6.770 2.350 6.910 ;
        RECT 2.650 6.980 2.940 7.010 ;
        RECT 2.650 6.810 2.980 6.980 ;
        RECT 2.650 6.770 2.940 6.810 ;
        RECT 3.560 6.770 3.890 7.030 ;
        RECT 5.100 6.770 5.370 7.210 ;
        RECT 0.000 6.570 0.620 6.740 ;
        RECT 0.630 6.290 0.810 6.750 ;
        RECT 1.170 6.470 1.350 6.760 ;
        RECT 1.590 6.410 1.800 6.740 ;
        RECT 2.090 6.600 2.420 6.770 ;
        RECT 2.660 6.600 4.820 6.770 ;
        RECT 2.090 6.550 2.320 6.600 ;
        RECT 5.070 6.590 5.400 6.770 ;
        RECT 5.750 6.630 5.920 6.690 ;
        RECT 2.150 6.320 2.320 6.550 ;
        RECT 5.730 6.410 5.950 6.630 ;
        RECT 5.750 6.360 5.920 6.410 ;
        RECT 2.150 6.310 2.530 6.320 ;
        RECT 0.630 6.120 1.590 6.290 ;
        RECT 2.060 6.250 2.530 6.310 ;
        RECT 2.060 6.200 2.870 6.250 ;
        RECT 2.060 6.140 2.880 6.200 ;
        RECT 2.140 6.080 2.880 6.140 ;
        RECT 2.140 6.030 2.530 6.080 ;
        RECT 0.160 5.690 0.330 5.730 ;
        RECT 0.160 5.670 1.310 5.690 ;
        RECT 0.160 5.500 1.350 5.670 ;
        RECT 1.800 5.640 2.260 5.670 ;
        RECT 3.570 5.640 3.920 5.740 ;
        RECT 1.800 5.500 2.910 5.640 ;
        RECT 2.090 5.470 2.910 5.500 ;
        RECT 3.150 5.470 4.320 5.640 ;
        RECT 4.570 5.470 5.330 5.640 ;
        RECT 2.090 5.330 2.350 5.470 ;
        RECT 0.560 5.000 0.890 5.170 ;
        RECT 1.170 5.160 2.350 5.330 ;
        RECT 5.100 5.460 5.330 5.470 ;
        RECT 1.170 5.010 1.950 5.160 ;
        RECT 2.090 5.020 2.350 5.160 ;
        RECT 2.650 5.230 2.940 5.260 ;
        RECT 2.650 5.060 2.980 5.230 ;
        RECT 2.650 5.020 2.940 5.060 ;
        RECT 3.560 5.020 3.890 5.280 ;
        RECT 5.100 5.020 5.370 5.460 ;
        RECT 0.000 4.820 0.620 4.990 ;
        RECT 0.630 4.540 0.810 5.000 ;
        RECT 1.170 4.720 1.350 5.010 ;
        RECT 1.590 4.660 1.800 4.990 ;
        RECT 2.090 4.850 2.420 5.020 ;
        RECT 2.660 4.850 4.820 5.020 ;
        RECT 2.090 4.800 2.320 4.850 ;
        RECT 5.070 4.840 5.400 5.020 ;
        RECT 5.750 4.880 5.920 4.940 ;
        RECT 2.150 4.570 2.320 4.800 ;
        RECT 5.730 4.660 5.950 4.880 ;
        RECT 5.750 4.610 5.920 4.660 ;
        RECT 2.150 4.560 2.530 4.570 ;
        RECT 0.630 4.370 1.590 4.540 ;
        RECT 2.060 4.500 2.530 4.560 ;
        RECT 2.060 4.450 2.870 4.500 ;
        RECT 2.060 4.390 2.880 4.450 ;
        RECT 2.140 4.330 2.880 4.390 ;
        RECT 2.140 4.280 2.530 4.330 ;
        RECT 0.160 3.940 0.330 3.980 ;
        RECT 0.160 3.920 1.310 3.940 ;
        RECT 0.160 3.750 1.350 3.920 ;
        RECT 1.800 3.890 2.260 3.920 ;
        RECT 3.570 3.890 3.920 3.990 ;
        RECT 1.800 3.750 2.910 3.890 ;
        RECT 2.090 3.720 2.910 3.750 ;
        RECT 3.150 3.720 4.320 3.890 ;
        RECT 4.570 3.720 5.330 3.890 ;
        RECT 2.090 3.580 2.350 3.720 ;
        RECT 0.560 3.250 0.890 3.420 ;
        RECT 1.170 3.410 2.350 3.580 ;
        RECT 5.100 3.710 5.330 3.720 ;
        RECT 1.170 3.260 1.950 3.410 ;
        RECT 2.090 3.270 2.350 3.410 ;
        RECT 2.650 3.480 2.940 3.510 ;
        RECT 2.650 3.310 2.980 3.480 ;
        RECT 2.650 3.270 2.940 3.310 ;
        RECT 3.560 3.270 3.890 3.530 ;
        RECT 5.100 3.270 5.370 3.710 ;
        RECT 0.000 3.070 0.620 3.240 ;
        RECT 0.630 2.790 0.810 3.250 ;
        RECT 1.170 2.970 1.350 3.260 ;
        RECT 1.590 2.910 1.800 3.240 ;
        RECT 2.090 3.100 2.420 3.270 ;
        RECT 2.660 3.100 4.820 3.270 ;
        RECT 2.090 3.050 2.320 3.100 ;
        RECT 5.070 3.090 5.400 3.270 ;
        RECT 5.750 3.130 5.920 3.190 ;
        RECT 2.150 2.820 2.320 3.050 ;
        RECT 5.730 2.910 5.950 3.130 ;
        RECT 5.750 2.860 5.920 2.910 ;
        RECT 2.150 2.810 2.530 2.820 ;
        RECT 0.630 2.620 1.590 2.790 ;
        RECT 2.060 2.750 2.530 2.810 ;
        RECT 2.060 2.700 2.870 2.750 ;
        RECT 2.060 2.640 2.880 2.700 ;
        RECT 2.140 2.580 2.880 2.640 ;
        RECT 2.140 2.530 2.530 2.580 ;
        RECT 0.160 2.190 0.330 2.230 ;
        RECT 0.160 2.170 1.310 2.190 ;
        RECT 0.160 2.000 1.350 2.170 ;
        RECT 1.800 2.140 2.260 2.170 ;
        RECT 3.570 2.140 3.920 2.240 ;
        RECT 1.800 2.000 2.910 2.140 ;
        RECT 2.090 1.970 2.910 2.000 ;
        RECT 3.150 1.970 4.320 2.140 ;
        RECT 4.570 1.970 5.330 2.140 ;
        RECT 2.090 1.830 2.350 1.970 ;
        RECT 0.560 1.500 0.890 1.670 ;
        RECT 1.170 1.660 2.350 1.830 ;
        RECT 5.100 1.960 5.330 1.970 ;
        RECT 1.170 1.510 1.950 1.660 ;
        RECT 2.090 1.520 2.350 1.660 ;
        RECT 2.650 1.730 2.940 1.760 ;
        RECT 2.650 1.560 2.980 1.730 ;
        RECT 2.650 1.520 2.940 1.560 ;
        RECT 3.560 1.520 3.890 1.780 ;
        RECT 5.100 1.520 5.370 1.960 ;
        RECT 0.000 1.320 0.620 1.490 ;
        RECT 0.630 1.040 0.810 1.500 ;
        RECT 1.170 1.220 1.350 1.510 ;
        RECT 1.590 1.160 1.800 1.490 ;
        RECT 2.090 1.350 2.420 1.520 ;
        RECT 2.660 1.350 4.820 1.520 ;
        RECT 2.090 1.300 2.320 1.350 ;
        RECT 5.070 1.340 5.400 1.520 ;
        RECT 5.750 1.380 5.920 1.440 ;
        RECT 2.150 1.070 2.320 1.300 ;
        RECT 5.730 1.160 5.950 1.380 ;
        RECT 5.750 1.110 5.920 1.160 ;
        RECT 2.150 1.060 2.530 1.070 ;
        RECT 0.630 0.870 1.590 1.040 ;
        RECT 2.060 1.000 2.530 1.060 ;
        RECT 2.060 0.950 2.870 1.000 ;
        RECT 2.060 0.890 2.880 0.950 ;
        RECT 2.140 0.830 2.880 0.890 ;
        RECT 2.140 0.780 2.530 0.830 ;
      LAYER mcon ;
        RECT 3.630 7.260 3.840 7.470 ;
        RECT 1.670 6.830 1.840 7.000 ;
        RECT 2.710 6.790 2.880 6.960 ;
        RECT 5.140 6.890 5.310 7.060 ;
        RECT 0.630 6.490 0.800 6.660 ;
        RECT 0.630 6.130 0.800 6.300 ;
        RECT 3.630 5.510 3.840 5.720 ;
        RECT 1.670 5.080 1.840 5.250 ;
        RECT 2.710 5.040 2.880 5.210 ;
        RECT 5.140 5.140 5.310 5.310 ;
        RECT 0.630 4.740 0.800 4.910 ;
        RECT 0.630 4.380 0.800 4.550 ;
        RECT 3.630 3.760 3.840 3.970 ;
        RECT 1.670 3.330 1.840 3.500 ;
        RECT 2.710 3.290 2.880 3.460 ;
        RECT 5.140 3.390 5.310 3.560 ;
        RECT 0.630 2.990 0.800 3.160 ;
        RECT 0.630 2.630 0.800 2.800 ;
        RECT 3.630 2.010 3.840 2.220 ;
        RECT 1.670 1.580 1.840 1.750 ;
        RECT 2.710 1.540 2.880 1.710 ;
        RECT 5.140 1.640 5.310 1.810 ;
        RECT 0.630 1.240 0.800 1.410 ;
        RECT 0.630 0.880 0.800 1.050 ;
      LAYER met1 ;
        RECT 1.600 6.800 1.920 7.080 ;
        RECT 1.560 6.780 1.920 6.800 ;
        RECT 1.560 6.470 1.840 6.780 ;
        RECT 2.090 6.180 2.400 7.870 ;
        RECT 3.570 7.220 3.920 7.510 ;
        RECT 7.880 7.370 8.120 7.440 ;
        RECT 3.720 7.200 3.920 7.220 ;
        RECT 2.650 7.010 2.960 7.020 ;
        RECT 2.640 6.740 2.960 7.010 ;
        RECT 2.650 6.730 2.940 6.740 ;
        RECT 5.670 6.360 6.080 6.690 ;
        RECT 1.600 5.050 1.920 5.330 ;
        RECT 1.560 5.030 1.920 5.050 ;
        RECT 1.560 4.720 1.840 5.030 ;
        RECT 2.090 4.430 2.400 6.120 ;
        RECT 3.570 5.470 3.920 5.760 ;
        RECT 5.100 5.690 5.340 6.110 ;
        RECT 4.870 5.630 5.340 5.690 ;
        RECT 3.720 5.450 3.920 5.470 ;
        RECT 2.650 5.260 2.960 5.270 ;
        RECT 2.640 4.990 2.960 5.260 ;
        RECT 2.650 4.980 2.940 4.990 ;
        RECT 5.100 4.430 5.340 5.630 ;
        RECT 7.880 5.620 8.120 5.690 ;
        RECT 5.670 4.610 6.080 4.940 ;
        RECT 1.600 3.300 1.920 3.580 ;
        RECT 1.560 3.280 1.920 3.300 ;
        RECT 1.560 2.970 1.840 3.280 ;
        RECT 2.090 2.680 2.400 4.370 ;
        RECT 3.570 3.720 3.920 4.010 ;
        RECT 5.100 3.940 5.340 4.360 ;
        RECT 4.870 3.880 5.340 3.940 ;
        RECT 3.720 3.700 3.920 3.720 ;
        RECT 2.650 3.510 2.960 3.520 ;
        RECT 2.640 3.240 2.960 3.510 ;
        RECT 2.650 3.230 2.940 3.240 ;
        RECT 5.100 2.680 5.340 3.880 ;
        RECT 7.880 3.870 8.120 3.940 ;
        RECT 5.670 2.860 6.080 3.190 ;
        RECT 1.600 1.550 1.920 1.830 ;
        RECT 1.560 1.530 1.920 1.550 ;
        RECT 1.560 1.220 1.840 1.530 ;
        RECT 2.090 0.930 2.400 2.620 ;
        RECT 3.570 1.970 3.920 2.260 ;
        RECT 5.100 2.190 5.340 2.610 ;
        RECT 4.870 2.130 5.340 2.190 ;
        RECT 3.720 1.950 3.920 1.970 ;
        RECT 2.650 1.760 2.960 1.770 ;
        RECT 2.640 1.490 2.960 1.760 ;
        RECT 2.650 1.480 2.940 1.490 ;
        RECT 5.100 0.930 5.340 2.130 ;
        RECT 7.880 2.120 8.120 2.190 ;
        RECT 5.670 1.110 6.080 1.440 ;
      LAYER via ;
        RECT 1.630 6.790 1.890 7.050 ;
        RECT 1.570 6.510 1.830 6.770 ;
        RECT 3.610 7.230 3.870 7.490 ;
        RECT 2.670 6.750 2.930 7.010 ;
        RECT 5.710 6.390 5.970 6.650 ;
        RECT 1.630 5.040 1.890 5.300 ;
        RECT 1.570 4.760 1.830 5.020 ;
        RECT 3.610 5.480 3.870 5.740 ;
        RECT 2.670 5.000 2.930 5.260 ;
        RECT 5.710 4.640 5.970 4.900 ;
        RECT 1.630 3.290 1.890 3.550 ;
        RECT 1.570 3.010 1.830 3.270 ;
        RECT 3.610 3.730 3.870 3.990 ;
        RECT 2.670 3.250 2.930 3.510 ;
        RECT 5.710 2.890 5.970 3.150 ;
        RECT 1.630 1.540 1.890 1.800 ;
        RECT 1.570 1.260 1.830 1.520 ;
        RECT 3.610 1.980 3.870 2.240 ;
        RECT 2.670 1.500 2.930 1.760 ;
        RECT 5.710 1.140 5.970 1.400 ;
      LAYER met2 ;
        RECT 1.600 7.000 1.920 7.050 ;
        RECT 2.630 7.010 2.950 7.020 ;
        RECT 2.630 7.000 2.960 7.010 ;
        RECT 0.290 6.800 2.960 7.000 ;
        RECT 1.600 6.790 1.920 6.800 ;
        RECT 1.530 6.720 1.870 6.780 ;
        RECT 2.630 6.750 2.960 6.800 ;
        RECT 2.630 6.730 2.950 6.750 ;
        RECT 3.610 6.720 3.870 7.520 ;
        RECT 1.530 6.500 3.970 6.720 ;
        RECT 5.680 6.360 6.140 6.680 ;
        RECT 1.600 5.250 1.920 5.300 ;
        RECT 2.630 5.260 2.950 5.270 ;
        RECT 2.630 5.250 2.960 5.260 ;
        RECT 0.290 5.050 2.960 5.250 ;
        RECT 1.600 5.040 1.920 5.050 ;
        RECT 1.530 4.970 1.870 5.030 ;
        RECT 2.630 5.000 2.960 5.050 ;
        RECT 2.630 4.980 2.950 5.000 ;
        RECT 3.610 4.970 3.870 5.770 ;
        RECT 1.530 4.750 3.970 4.970 ;
        RECT 5.680 4.610 6.140 4.930 ;
        RECT 1.600 3.500 1.920 3.550 ;
        RECT 2.630 3.510 2.950 3.520 ;
        RECT 2.630 3.500 2.960 3.510 ;
        RECT 0.290 3.300 2.960 3.500 ;
        RECT 1.600 3.290 1.920 3.300 ;
        RECT 1.530 3.220 1.870 3.280 ;
        RECT 2.630 3.250 2.960 3.300 ;
        RECT 2.630 3.230 2.950 3.250 ;
        RECT 3.610 3.220 3.870 4.020 ;
        RECT 1.530 3.000 3.970 3.220 ;
        RECT 5.680 2.860 6.140 3.180 ;
        RECT 1.600 1.750 1.920 1.800 ;
        RECT 2.630 1.760 2.950 1.770 ;
        RECT 2.630 1.750 2.960 1.760 ;
        RECT 0.290 1.550 2.960 1.750 ;
        RECT 1.600 1.540 1.920 1.550 ;
        RECT 1.530 1.470 1.870 1.530 ;
        RECT 2.630 1.500 2.960 1.550 ;
        RECT 2.630 1.480 2.950 1.500 ;
        RECT 3.610 1.470 3.870 2.270 ;
        RECT 1.530 1.250 3.970 1.470 ;
        RECT 5.680 1.110 6.140 1.430 ;
  END
END sky130_hilas_LevelShift4InputUp

MACRO sky130_hilas_WTA4Stage01
  CLASS CORE ;
  FOREIGN sky130_hilas_WTA4Stage01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.920 BY 14.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 25.990 5.730 26.220 6.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.990 0.140 26.220 0.390 ;
    END
  END VGND
  PIN OUTPUT1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 25.120 4.830 26.380 4.990 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.476800 ;
    ANTENNADIFFAREA 0.725100 ;
    PORT
      LAYER met2 ;
        RECT 24.480 4.810 24.790 5.070 ;
        RECT 24.330 4.650 26.920 4.810 ;
        RECT 24.330 4.480 24.640 4.650 ;
        RECT 24.330 4.220 24.640 4.390 ;
        RECT 24.330 4.060 26.920 4.220 ;
        RECT 24.480 3.800 24.790 4.060 ;
        RECT 25.120 3.900 26.380 4.060 ;
    END
  END OUTPUT2
  PIN OUTPUT3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 25.120 2.060 26.380 2.220 ;
    END
  END OUTPUT3
  PIN OUTPUT4
    USE ANALOG ;
    ANTENNAGATEAREA 0.476800 ;
    ANTENNADIFFAREA 0.725100 ;
    PORT
      LAYER met2 ;
        RECT 24.480 2.040 24.790 2.300 ;
        RECT 24.330 1.880 26.920 2.040 ;
        RECT 24.330 1.730 24.640 1.880 ;
        RECT 25.930 1.730 26.260 1.820 ;
        RECT 19.580 1.560 26.260 1.730 ;
        RECT 24.330 1.450 24.640 1.560 ;
        RECT 25.930 1.530 26.260 1.560 ;
        RECT 24.330 1.290 26.920 1.450 ;
        RECT 24.480 1.030 24.790 1.290 ;
        RECT 25.140 1.130 26.380 1.290 ;
    END
  END OUTPUT4
  PIN INPUT1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 12.300 4.840 12.450 5.260 ;
        RECT 12.300 4.750 15.570 4.840 ;
        RECT 15.640 4.750 15.960 4.950 ;
        RECT 12.300 4.690 15.960 4.750 ;
        RECT 15.430 4.590 15.730 4.690 ;
    END
  END INPUT1
  PIN INPUT2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 12.370 4.360 12.690 4.450 ;
        RECT 12.280 4.190 12.690 4.360 ;
        RECT 12.280 4.090 12.600 4.190 ;
        RECT 15.510 3.610 15.740 3.620 ;
        RECT 15.510 3.580 23.080 3.610 ;
        RECT 12.350 3.310 12.670 3.440 ;
        RECT 15.510 3.410 23.140 3.580 ;
        RECT 15.510 3.310 15.750 3.410 ;
        RECT 12.300 3.130 15.750 3.310 ;
        RECT 22.950 3.210 23.660 3.410 ;
        RECT 12.300 3.110 15.670 3.130 ;
    END
  END INPUT2
  PIN INPUT3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 15.640 2.930 15.960 3.070 ;
        RECT 15.640 2.910 23.100 2.930 ;
        RECT 15.640 2.810 23.660 2.910 ;
        RECT 15.650 2.710 23.660 2.810 ;
        RECT 15.650 2.700 15.970 2.710 ;
        RECT 12.240 1.750 12.440 2.250 ;
        RECT 15.510 1.750 15.830 1.890 ;
        RECT 12.240 1.630 15.830 1.750 ;
        RECT 12.240 1.550 15.790 1.630 ;
    END
  END INPUT3
  PIN INPUT4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 12.350 1.310 12.660 1.490 ;
        RECT 12.230 1.160 12.660 1.310 ;
        RECT 12.230 1.040 12.510 1.160 ;
        RECT 12.240 0.520 12.810 0.700 ;
        RECT 23.100 0.650 23.650 0.660 ;
        RECT 12.400 0.370 12.710 0.520 ;
        RECT 12.280 0.240 12.710 0.370 ;
        RECT 15.520 0.430 23.650 0.650 ;
        RECT 15.520 0.420 23.110 0.430 ;
        RECT 15.520 0.410 16.290 0.420 ;
        RECT 15.520 0.240 15.760 0.410 ;
        RECT 12.280 0.160 15.760 0.240 ;
        RECT 12.390 0.000 15.760 0.160 ;
    END
  END INPUT4
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 12.260 5.720 12.990 5.900 ;
    END
  END DRAIN1
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT 18.100 6.090 18.480 6.190 ;
    END
  END GATE1
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 22.130 5.910 22.530 6.190 ;
    END
  END VTUN
  PIN WTAMIDDLENODE
    PORT
      LAYER met1 ;
        RECT 24.730 0.140 24.960 0.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 24.730 5.730 24.960 6.190 ;
    END
  END WTAMIDDLENODE
  PIN COLSEL1
    ANTENNADIFFAREA 1.047900 ;
    PORT
      LAYER met2 ;
        RECT 13.360 6.070 13.680 6.130 ;
        RECT 17.380 6.070 17.710 6.100 ;
        RECT 13.360 5.900 17.710 6.070 ;
        RECT 13.360 5.850 13.680 5.900 ;
        RECT 15.660 5.880 15.980 5.900 ;
        RECT 17.380 5.880 17.710 5.900 ;
        RECT 15.660 5.740 23.490 5.880 ;
        RECT 15.840 5.690 23.490 5.740 ;
        RECT 15.840 5.680 23.660 5.690 ;
        RECT 12.610 5.670 23.660 5.680 ;
        RECT 12.610 5.510 20.240 5.670 ;
        RECT 23.280 5.480 23.660 5.670 ;
    END
  END COLSEL1
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 13.980 6.120 14.140 6.190 ;
    END
  END VPWR
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 13.170 6.120 13.330 6.190 ;
    END
  END VINJ
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 12.230 3.770 12.810 3.950 ;
    END
  END DRAIN2
  PIN DRAIN3
    PORT
      LAYER met2 ;
        RECT 12.260 2.480 12.810 2.660 ;
    END
  END DRAIN3
  OBS
      LAYER nwell ;
        RECT 4.000 14.810 5.730 14.870 ;
        RECT 0.000 11.240 1.730 13.080 ;
        RECT 4.000 8.370 6.920 14.810 ;
        RECT 7.280 9.370 9.840 11.280 ;
        RECT 4.690 8.320 6.920 8.370 ;
        RECT 7.280 6.130 9.840 9.120 ;
        RECT 14.820 9.080 15.930 9.350 ;
        RECT 19.080 9.140 19.670 9.300 ;
        RECT 12.640 8.160 12.730 8.240 ;
        RECT 11.120 7.660 11.290 7.720 ;
        RECT 10.940 7.650 11.290 7.660 ;
        RECT 10.940 7.550 10.950 7.650 ;
        RECT 11.120 7.550 11.290 7.650 ;
        RECT 12.410 6.180 15.370 6.190 ;
        RECT 12.410 6.030 12.820 6.180 ;
        RECT 18.100 6.090 18.480 6.190 ;
        RECT 12.410 6.020 13.000 6.030 ;
        RECT 7.280 3.960 9.840 5.870 ;
        RECT 12.410 4.260 12.820 6.020 ;
        RECT 14.820 5.880 15.930 6.070 ;
        RECT 22.130 6.050 22.530 6.190 ;
        RECT 19.080 5.900 19.670 6.050 ;
        RECT 12.300 3.840 12.820 4.260 ;
        RECT 12.300 3.640 12.810 3.840 ;
        RECT 12.300 3.110 12.820 3.640 ;
        RECT 12.410 0.150 12.820 3.110 ;
      LAYER li1 ;
        RECT 0.760 11.690 1.310 12.120 ;
        RECT 4.790 11.760 5.340 12.190 ;
        RECT 9.280 10.930 9.600 10.970 ;
        RECT 7.680 10.540 7.880 10.890 ;
        RECT 9.270 10.810 9.600 10.930 ;
        RECT 9.160 10.710 9.600 10.810 ;
        RECT 9.160 10.640 9.500 10.710 ;
        RECT 7.670 10.510 7.880 10.540 ;
        RECT 7.670 9.920 7.890 10.510 ;
        RECT 8.410 9.920 8.610 10.520 ;
        RECT 9.280 10.380 9.600 10.420 ;
        RECT 9.270 10.190 9.600 10.380 ;
        RECT 9.160 10.160 9.600 10.190 ;
        RECT 9.160 10.020 9.500 10.160 ;
        RECT 13.440 8.820 13.610 9.350 ;
        RECT 17.460 8.850 17.630 9.380 ;
        RECT 7.670 7.980 7.890 8.570 ;
        RECT 7.670 7.950 7.880 7.980 ;
        RECT 8.410 7.970 8.610 8.570 ;
        RECT 9.160 8.330 9.500 8.470 ;
        RECT 9.160 8.300 9.600 8.330 ;
        RECT 9.270 8.110 9.600 8.300 ;
        RECT 9.280 8.070 9.600 8.110 ;
        RECT 7.680 7.300 7.880 7.950 ;
        RECT 9.160 7.780 9.500 7.850 ;
        RECT 9.160 7.680 9.600 7.780 ;
        RECT 9.270 7.570 9.600 7.680 ;
        RECT 9.160 7.470 9.600 7.570 ;
        RECT 10.940 7.550 11.380 7.720 ;
        RECT 9.160 7.400 9.500 7.470 ;
        RECT 7.670 7.270 7.880 7.300 ;
        RECT 7.670 6.680 7.890 7.270 ;
        RECT 8.410 6.680 8.610 7.280 ;
        RECT 9.280 7.140 9.600 7.180 ;
        RECT 9.270 6.950 9.600 7.140 ;
        RECT 13.430 6.960 13.600 8.150 ;
        RECT 9.160 6.920 9.600 6.950 ;
        RECT 17.450 6.920 17.620 8.090 ;
        RECT 9.160 6.780 9.500 6.920 ;
        RECT 7.670 4.730 7.890 5.320 ;
        RECT 7.670 4.700 7.880 4.730 ;
        RECT 8.410 4.720 8.610 5.320 ;
        RECT 25.280 5.280 25.490 5.300 ;
        RECT 9.160 5.080 9.500 5.220 ;
        RECT 25.260 5.110 25.930 5.280 ;
        RECT 9.160 5.050 9.600 5.080 ;
        RECT 9.270 4.860 9.600 5.050 ;
        RECT 9.280 4.820 9.600 4.860 ;
        RECT 24.490 4.990 24.810 5.030 ;
        RECT 24.490 4.900 24.820 4.990 ;
        RECT 25.260 4.900 25.510 5.110 ;
        RECT 24.490 4.880 25.990 4.900 ;
        RECT 24.490 4.780 26.070 4.880 ;
        RECT 24.340 4.730 26.070 4.780 ;
        RECT 7.680 4.350 7.880 4.700 ;
        RECT 9.160 4.530 9.500 4.600 ;
        RECT 24.340 4.560 25.010 4.730 ;
        RECT 25.180 4.710 25.510 4.730 ;
        RECT 25.730 4.710 26.070 4.730 ;
        RECT 9.160 4.430 9.600 4.530 ;
        RECT 24.340 4.520 24.660 4.560 ;
        RECT 9.270 4.310 9.600 4.430 ;
        RECT 9.280 4.270 9.600 4.310 ;
        RECT 24.340 4.310 24.660 4.350 ;
        RECT 24.670 4.310 25.010 4.560 ;
        RECT 25.260 4.540 25.430 4.710 ;
        RECT 25.820 4.540 25.990 4.710 ;
        RECT 25.180 4.330 25.510 4.540 ;
        RECT 25.730 4.330 26.070 4.540 ;
        RECT 24.340 4.140 25.010 4.310 ;
        RECT 25.260 4.160 25.430 4.330 ;
        RECT 25.820 4.160 25.990 4.330 ;
        RECT 25.180 4.140 25.510 4.160 ;
        RECT 25.730 4.140 26.070 4.160 ;
        RECT 24.340 4.090 26.070 4.140 ;
        RECT 24.490 3.990 26.070 4.090 ;
        RECT 24.490 3.970 25.990 3.990 ;
        RECT 24.490 3.880 24.820 3.970 ;
        RECT 24.490 3.840 24.810 3.880 ;
        RECT 25.260 3.760 25.510 3.970 ;
        RECT 26.390 3.910 26.900 4.960 ;
        RECT 25.260 3.590 25.930 3.760 ;
        RECT 25.280 3.570 25.490 3.590 ;
        RECT 25.280 2.510 25.490 2.530 ;
        RECT 25.260 2.340 25.930 2.510 ;
        RECT 24.490 2.220 24.810 2.260 ;
        RECT 24.490 2.130 24.820 2.220 ;
        RECT 25.260 2.130 25.510 2.340 ;
        RECT 24.490 2.110 25.990 2.130 ;
        RECT 24.490 2.010 26.070 2.110 ;
        RECT 24.340 1.960 26.070 2.010 ;
        RECT 24.340 1.790 25.010 1.960 ;
        RECT 25.180 1.940 25.510 1.960 ;
        RECT 25.730 1.940 26.070 1.960 ;
        RECT 24.340 1.750 24.660 1.790 ;
        RECT 24.340 1.540 24.660 1.580 ;
        RECT 24.670 1.540 25.010 1.790 ;
        RECT 25.260 1.770 25.430 1.940 ;
        RECT 25.820 1.770 25.990 1.940 ;
        RECT 25.180 1.560 25.510 1.770 ;
        RECT 25.730 1.560 26.070 1.770 ;
        RECT 12.360 1.410 12.680 1.450 ;
        RECT 12.360 1.240 12.690 1.410 ;
        RECT 24.340 1.370 25.010 1.540 ;
        RECT 25.260 1.390 25.430 1.560 ;
        RECT 25.820 1.390 25.990 1.560 ;
        RECT 25.180 1.370 25.510 1.390 ;
        RECT 25.730 1.370 26.070 1.390 ;
        RECT 24.340 1.320 26.070 1.370 ;
        RECT 12.270 1.220 12.690 1.240 ;
        RECT 24.490 1.220 26.070 1.320 ;
        RECT 12.270 1.190 12.680 1.220 ;
        RECT 24.490 1.200 25.990 1.220 ;
        RECT 12.270 0.490 12.450 1.190 ;
        RECT 24.490 1.110 24.820 1.200 ;
        RECT 24.490 1.070 24.810 1.110 ;
        RECT 25.260 0.990 25.510 1.200 ;
        RECT 26.390 1.140 26.900 2.190 ;
        RECT 25.260 0.820 25.930 0.990 ;
        RECT 25.280 0.800 25.490 0.820 ;
        RECT 12.270 0.450 12.730 0.490 ;
        RECT 12.270 0.320 12.740 0.450 ;
        RECT 12.410 0.260 12.740 0.320 ;
        RECT 12.410 0.230 12.730 0.260 ;
      LAYER mcon ;
        RECT 1.040 11.770 1.310 12.040 ;
        RECT 5.070 11.840 5.340 12.110 ;
        RECT 9.370 10.750 9.540 10.920 ;
        RECT 7.700 10.340 7.870 10.510 ;
        RECT 8.430 10.310 8.600 10.480 ;
        RECT 9.370 10.200 9.540 10.370 ;
        RECT 13.440 9.180 13.610 9.350 ;
        RECT 17.460 9.210 17.630 9.380 ;
        RECT 7.700 7.980 7.870 8.150 ;
        RECT 8.430 8.010 8.600 8.180 ;
        RECT 9.370 8.120 9.540 8.290 ;
        RECT 13.430 7.980 13.600 8.150 ;
        RECT 9.370 7.510 9.540 7.740 ;
        RECT 13.430 7.320 13.600 7.490 ;
        RECT 7.700 7.100 7.870 7.270 ;
        RECT 8.430 7.070 8.600 7.240 ;
        RECT 9.370 6.960 9.540 7.130 ;
        RECT 17.450 7.920 17.620 8.090 ;
        RECT 17.450 7.280 17.620 7.450 ;
        RECT 7.700 4.730 7.870 4.900 ;
        RECT 25.300 5.110 25.470 5.280 ;
        RECT 8.430 4.760 8.600 4.930 ;
        RECT 9.370 4.870 9.540 5.040 ;
        RECT 24.550 4.810 24.720 4.980 ;
        RECT 24.400 4.570 24.570 4.740 ;
        RECT 9.370 4.320 9.540 4.490 ;
        RECT 26.560 4.540 26.730 4.710 ;
        RECT 24.400 4.130 24.570 4.300 ;
        RECT 26.560 4.160 26.730 4.330 ;
        RECT 24.550 3.890 24.720 4.060 ;
        RECT 25.300 3.590 25.470 3.760 ;
        RECT 25.300 2.340 25.470 2.510 ;
        RECT 24.550 2.040 24.720 2.210 ;
        RECT 24.400 1.800 24.570 1.970 ;
        RECT 26.560 1.770 26.730 1.940 ;
        RECT 12.420 1.230 12.590 1.400 ;
        RECT 24.400 1.360 24.570 1.530 ;
        RECT 26.560 1.390 26.730 1.560 ;
        RECT 24.550 1.120 24.720 1.290 ;
        RECT 25.300 0.820 25.470 0.990 ;
        RECT 12.470 0.270 12.640 0.440 ;
      LAYER met1 ;
        RECT 0.980 11.230 1.370 13.090 ;
        RECT 5.010 11.300 5.400 13.160 ;
        RECT 5.890 8.320 6.270 14.820 ;
        RECT 7.640 10.570 7.800 11.270 ;
        RECT 7.640 10.020 7.910 10.570 ;
        RECT 7.630 9.970 7.910 10.020 ;
        RECT 8.050 10.230 8.240 11.220 ;
        RECT 8.450 10.540 8.610 11.270 ;
        RECT 9.290 10.680 9.610 11.000 ;
        RECT 8.410 10.520 8.610 10.540 ;
        RECT 10.530 10.530 10.690 10.600 ;
        RECT 10.940 10.530 11.130 10.600 ;
        RECT 11.340 10.530 11.500 10.600 ;
        RECT 8.400 10.280 8.630 10.520 ;
        RECT 8.400 10.230 8.610 10.280 ;
        RECT 8.050 10.110 8.220 10.230 ;
        RECT 7.630 9.880 7.800 9.970 ;
        RECT 7.640 9.370 7.800 9.880 ;
        RECT 8.050 9.370 8.210 10.110 ;
        RECT 8.450 9.370 8.610 10.230 ;
        RECT 9.290 10.130 9.610 10.450 ;
        RECT 7.640 8.610 7.800 9.120 ;
        RECT 7.630 8.520 7.800 8.610 ;
        RECT 7.630 8.470 7.910 8.520 ;
        RECT 7.640 7.920 7.910 8.470 ;
        RECT 8.050 8.380 8.210 9.120 ;
        RECT 8.050 8.260 8.220 8.380 ;
        RECT 8.450 8.260 8.610 9.120 ;
        RECT 7.640 7.330 7.800 7.920 ;
        RECT 7.640 6.780 7.910 7.330 ;
        RECT 7.630 6.730 7.910 6.780 ;
        RECT 8.050 6.990 8.240 8.260 ;
        RECT 8.400 8.210 8.610 8.260 ;
        RECT 8.400 7.970 8.630 8.210 ;
        RECT 9.290 8.040 9.610 8.360 ;
        RECT 8.410 7.950 8.610 7.970 ;
        RECT 8.450 7.300 8.610 7.950 ;
        RECT 9.290 7.440 9.610 7.810 ;
        RECT 10.910 7.720 11.150 7.750 ;
        RECT 10.910 7.630 11.340 7.720 ;
        RECT 10.530 7.620 10.690 7.630 ;
        RECT 10.910 7.620 11.500 7.630 ;
        RECT 10.910 7.550 11.340 7.620 ;
        RECT 10.910 7.520 11.150 7.550 ;
        RECT 10.940 7.420 11.050 7.520 ;
        RECT 8.410 7.280 8.610 7.300 ;
        RECT 8.400 7.040 8.630 7.280 ;
        RECT 8.400 6.990 8.610 7.040 ;
        RECT 8.050 6.870 8.220 6.990 ;
        RECT 7.630 6.640 7.800 6.730 ;
        RECT 7.640 6.130 7.800 6.640 ;
        RECT 8.050 6.130 8.210 6.870 ;
        RECT 8.450 6.130 8.610 6.990 ;
        RECT 9.290 6.890 9.610 7.210 ;
        RECT 13.400 6.190 13.650 10.870 ;
        RECT 15.460 10.500 15.840 10.870 ;
        RECT 13.400 6.160 13.770 6.190 ;
        RECT 13.380 6.130 13.770 6.160 ;
        RECT 17.410 6.130 17.680 10.870 ;
        RECT 13.370 6.120 13.770 6.130 ;
        RECT 7.640 5.360 7.800 5.870 ;
        RECT 7.630 5.270 7.800 5.360 ;
        RECT 7.630 5.220 7.910 5.270 ;
        RECT 7.640 4.670 7.910 5.220 ;
        RECT 8.050 5.130 8.210 5.870 ;
        RECT 8.050 5.010 8.220 5.130 ;
        RECT 8.450 5.010 8.610 5.870 ;
        RECT 13.370 5.850 13.670 6.120 ;
        RECT 13.380 5.830 13.660 5.850 ;
        RECT 7.640 3.970 7.800 4.670 ;
        RECT 8.050 4.020 8.240 5.010 ;
        RECT 8.400 4.960 8.610 5.010 ;
        RECT 8.400 4.720 8.630 4.960 ;
        RECT 9.290 4.790 9.610 5.110 ;
        RECT 8.410 4.700 8.610 4.720 ;
        RECT 8.450 3.970 8.610 4.700 ;
        RECT 10.530 4.560 10.690 4.630 ;
        RECT 10.940 4.560 11.130 4.630 ;
        RECT 11.340 4.560 11.500 4.630 ;
        RECT 9.290 4.240 9.610 4.560 ;
        RECT 12.400 4.260 12.660 4.480 ;
        RECT 13.400 4.370 13.650 5.830 ;
        RECT 15.690 5.710 15.950 6.030 ;
        RECT 17.390 5.820 17.700 6.130 ;
        RECT 15.600 4.980 15.810 5.610 ;
        RECT 15.600 4.870 15.930 4.980 ;
        RECT 15.670 4.660 15.930 4.870 ;
        RECT 15.460 4.370 15.840 4.650 ;
        RECT 17.410 4.370 17.680 5.820 ;
        RECT 19.490 4.370 19.890 10.870 ;
        RECT 24.480 4.810 24.800 5.060 ;
        RECT 24.330 4.740 24.800 4.810 ;
        RECT 24.330 4.490 24.650 4.740 ;
        RECT 12.300 4.160 12.660 4.260 ;
        RECT 12.300 3.470 12.510 4.160 ;
        RECT 24.330 4.130 24.650 4.380 ;
        RECT 24.330 4.060 24.800 4.130 ;
        RECT 24.480 3.810 24.800 4.060 ;
        RECT 25.270 3.530 25.500 5.340 ;
        RECT 26.530 3.670 26.760 5.200 ;
        RECT 12.300 3.150 12.640 3.470 ;
        RECT 12.300 3.110 12.510 3.150 ;
        RECT 15.670 3.000 15.930 3.100 ;
        RECT 15.580 2.780 15.930 3.000 ;
        RECT 24.190 2.950 24.420 3.150 ;
        RECT 25.450 2.950 25.680 3.160 ;
        RECT 15.580 1.920 15.740 2.780 ;
        RECT 24.480 2.040 24.800 2.290 ;
        RECT 24.330 1.970 24.800 2.040 ;
        RECT 15.540 1.600 15.800 1.920 ;
        RECT 24.330 1.720 24.650 1.970 ;
        RECT 15.580 1.500 15.740 1.600 ;
        RECT 12.350 1.160 12.670 1.480 ;
        RECT 24.330 1.360 24.650 1.610 ;
        RECT 24.330 1.290 24.800 1.360 ;
        RECT 24.480 1.040 24.800 1.290 ;
        RECT 25.270 0.760 25.500 2.570 ;
        RECT 25.990 1.840 26.220 1.890 ;
        RECT 25.950 1.830 26.230 1.840 ;
        RECT 25.950 1.510 26.250 1.830 ;
        RECT 26.530 0.900 26.760 2.430 ;
        RECT 12.400 0.200 12.720 0.520 ;
        RECT 18.100 0.140 18.480 0.240 ;
      LAYER via ;
        RECT 9.320 10.710 9.580 10.970 ;
        RECT 9.320 10.160 9.580 10.420 ;
        RECT 9.320 8.070 9.580 8.330 ;
        RECT 9.320 7.470 9.580 7.780 ;
        RECT 9.320 6.920 9.580 7.180 ;
        RECT 13.390 5.860 13.650 6.120 ;
        RECT 9.320 4.820 9.580 5.080 ;
        RECT 9.320 4.270 9.580 4.530 ;
        RECT 12.400 4.190 12.660 4.450 ;
        RECT 15.690 5.740 15.950 6.000 ;
        RECT 17.410 5.840 17.680 6.100 ;
        RECT 15.670 4.690 15.930 4.950 ;
        RECT 24.510 4.780 24.770 5.030 ;
        RECT 24.360 4.770 24.770 4.780 ;
        RECT 24.360 4.520 24.620 4.770 ;
        RECT 24.360 4.100 24.620 4.350 ;
        RECT 24.360 4.090 24.770 4.100 ;
        RECT 24.510 3.840 24.770 4.090 ;
        RECT 12.380 3.180 12.640 3.440 ;
        RECT 15.670 2.810 15.930 3.070 ;
        RECT 24.510 2.010 24.770 2.260 ;
        RECT 15.540 1.630 15.800 1.890 ;
        RECT 24.360 2.000 24.770 2.010 ;
        RECT 24.360 1.750 24.620 2.000 ;
        RECT 12.380 1.190 12.640 1.450 ;
        RECT 24.360 1.330 24.620 1.580 ;
        RECT 24.360 1.320 24.770 1.330 ;
        RECT 24.510 1.070 24.770 1.320 ;
        RECT 25.960 1.540 26.230 1.810 ;
        RECT 12.430 0.230 12.690 0.490 ;
      LAYER met2 ;
        RECT 9.300 10.720 9.610 11.010 ;
        RECT 7.280 10.680 9.610 10.720 ;
        RECT 7.280 10.540 9.460 10.680 ;
        RECT 9.300 10.290 9.610 10.460 ;
        RECT 7.280 10.130 9.610 10.290 ;
        RECT 7.280 10.110 9.450 10.130 ;
        RECT 9.750 10.110 9.840 10.290 ;
        RECT 10.170 10.130 10.260 10.310 ;
        RECT 10.170 9.700 10.260 9.880 ;
        RECT 12.630 9.690 20.240 9.880 ;
        RECT 10.170 8.610 10.260 8.790 ;
        RECT 12.610 8.610 20.240 8.790 ;
        RECT 7.280 8.360 9.450 8.380 ;
        RECT 7.280 8.200 9.610 8.360 ;
        RECT 9.750 8.200 9.840 8.380 ;
        RECT 9.300 8.030 9.610 8.200 ;
        RECT 10.170 8.180 10.260 8.360 ;
        RECT 12.640 8.170 12.730 8.200 ;
        RECT 12.610 8.060 12.730 8.170 ;
        RECT 7.280 7.810 9.460 7.950 ;
        RECT 7.280 7.770 9.610 7.810 ;
        RECT 9.300 7.480 9.610 7.770 ;
        RECT 7.280 7.440 9.610 7.480 ;
        RECT 7.280 7.300 9.460 7.440 ;
        RECT 9.300 7.050 9.610 7.220 ;
        RECT 7.280 6.890 9.610 7.050 ;
        RECT 7.280 6.870 9.450 6.890 ;
        RECT 9.750 6.870 9.840 7.050 ;
        RECT 10.170 6.890 10.280 7.070 ;
        RECT 12.610 6.910 12.760 7.080 ;
        RECT 10.170 6.460 10.280 6.640 ;
        RECT 12.610 6.470 19.470 6.640 ;
        RECT 19.770 6.500 20.240 6.660 ;
        RECT 19.770 6.490 20.230 6.500 ;
        RECT 10.170 5.360 10.280 5.540 ;
        RECT 22.770 5.470 22.910 5.480 ;
        RECT 22.770 5.140 22.920 5.470 ;
        RECT 7.280 5.110 9.450 5.130 ;
        RECT 7.280 4.950 9.610 5.110 ;
        RECT 9.750 4.950 9.840 5.130 ;
        RECT 9.300 4.780 9.610 4.950 ;
        RECT 10.170 4.930 10.280 5.110 ;
        RECT 22.770 4.940 23.980 5.140 ;
        RECT 24.090 4.710 24.210 4.920 ;
        RECT 7.280 4.560 9.460 4.700 ;
        RECT 7.280 4.520 9.610 4.560 ;
        RECT 9.300 4.230 9.610 4.520 ;
        RECT 22.880 4.280 24.080 4.380 ;
        RECT 22.870 4.200 24.080 4.280 ;
        RECT 23.800 4.080 24.080 4.200 ;
        RECT 23.800 4.060 23.830 4.080 ;
        RECT 24.090 3.950 24.210 4.160 ;
        RECT 22.860 2.090 23.860 2.250 ;
        RECT 24.090 1.940 24.210 2.150 ;
        RECT 22.870 1.110 23.870 1.280 ;
        RECT 24.090 1.180 24.210 1.390 ;
        RECT 22.870 1.100 23.810 1.110 ;
  END
END sky130_hilas_WTA4Stage01

MACRO sky130_hilas_Trans4small
  CLASS CORE ;
  FOREIGN sky130_hilas_Trans4small ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.400 BY 6.460 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN NFET_SOURCE1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 5.710 0.070 5.750 ;
        RECT 0.000 5.480 0.140 5.710 ;
    END
  END NFET_SOURCE1
  PIN NFET_GATE1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 5.070 0.160 5.240 ;
    END
  END NFET_GATE1
  PIN NFET_SOURCE2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 4.560 0.140 4.730 ;
    END
  END NFET_SOURCE2
  PIN NFET_GATE2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 4.150 0.170 4.320 ;
    END
  END NFET_GATE2
  PIN NFET_SOURCE3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 3.780 0.140 3.810 ;
        RECT 0.000 3.640 0.210 3.780 ;
    END
  END NFET_SOURCE3
  PIN NFET_GATE3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 3.230 0.160 3.400 ;
    END
  END NFET_GATE3
  PIN PFET_SOURCE1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 2.620 0.140 2.810 ;
    END
  END PFET_SOURCE1
  PIN PFET_GATE1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 2.200 0.140 2.390 ;
    END
  END PFET_GATE1
  PIN PFET_SOURCE2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 1.830 0.140 1.850 ;
        RECT 0.000 1.660 0.070 1.830 ;
    END
  END PFET_SOURCE2
  PIN PFET_GATE2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 1.410 0.140 1.430 ;
        RECT 0.000 1.240 0.070 1.410 ;
    END
  END PFET_GATE2
  PIN PFET_SOURCE3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 0.840 0.140 0.890 ;
        RECT 0.000 0.700 0.070 0.840 ;
    END
  END PFET_SOURCE3
  PIN PFET_GATE3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 0.450 0.140 0.470 ;
        RECT 0.000 0.280 0.150 0.450 ;
    END
  END PFET_GATE3
  PIN WELL
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 1.280 0.740 3.310 3.710 ;
        RECT 2.100 0.630 2.640 0.740 ;
        RECT 1.920 0.180 2.640 0.630 ;
        RECT 0.070 0.000 2.640 0.180 ;
      LAYER met2 ;
        RECT 1.850 1.790 2.170 1.990 ;
        RECT 1.850 1.710 2.800 1.790 ;
        RECT 1.760 1.590 2.800 1.710 ;
        RECT 1.760 1.380 2.070 1.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.850 1.950 2.170 1.990 ;
        RECT 1.620 1.720 2.170 1.950 ;
        RECT 1.850 1.700 2.170 1.720 ;
        RECT 1.760 1.670 2.170 1.700 ;
        RECT 1.760 1.380 2.080 1.670 ;
        RECT 2.180 1.270 2.400 5.880 ;
        RECT 2.160 1.200 2.400 1.270 ;
        RECT 2.160 1.100 2.500 1.200 ;
        RECT 2.180 0.970 2.500 1.100 ;
        RECT 2.180 0.000 2.400 0.970 ;
      LAYER via ;
        RECT 1.880 1.700 2.140 1.960 ;
        RECT 1.790 1.410 2.050 1.670 ;
    END
  END WELL
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 1.850 5.080 2.160 5.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.850 5.080 2.170 5.400 ;
        RECT 2.580 5.330 2.800 5.880 ;
        RECT 2.580 5.040 2.900 5.330 ;
        RECT 2.580 0.000 2.800 5.040 ;
      LAYER via ;
        RECT 1.880 5.110 2.140 5.370 ;
    END
  END VGND
  PIN PFET_DRAIN3
    USE ANALOG ;
    ANTENNAGATEAREA 0.163800 ;
    PORT
      LAYER met2 ;
        RECT 1.850 0.830 2.170 1.000 ;
        RECT 1.850 0.680 2.800 0.830 ;
        RECT 1.990 0.630 2.800 0.680 ;
    END
  END PFET_DRAIN3
  PIN PFET_DRAIN1
    USE ANALOG ;
    ANTENNAGATEAREA 0.163800 ;
    ANTENNADIFFAREA 0.117600 ;
    PORT
      LAYER met2 ;
        RECT 1.850 2.750 2.170 2.980 ;
        RECT 1.850 2.700 2.800 2.750 ;
        RECT 1.760 2.550 2.800 2.700 ;
        RECT 1.760 2.370 2.070 2.550 ;
    END
  END PFET_DRAIN1
  PIN NFET_DRAIN3
    USE ANALOG ;
    ANTENNAGATEAREA 0.113400 ;
    ANTENNADIFFAREA 0.117600 ;
    PORT
      LAYER met2 ;
        RECT 1.980 3.690 2.800 3.820 ;
        RECT 1.760 3.650 2.800 3.690 ;
        RECT 1.760 3.360 2.070 3.650 ;
    END
  END NFET_DRAIN3
  PIN NFET_DRAIN2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.980 4.570 2.800 4.740 ;
    END
  END NFET_DRAIN2
  PIN NFET_DRAIN1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.980 5.490 2.800 5.660 ;
    END
  END NFET_DRAIN1
  OBS
      LAYER li1 ;
        RECT 1.850 6.320 2.170 6.360 ;
        RECT 2.940 6.330 3.260 6.370 ;
        RECT 1.850 6.250 2.180 6.320 ;
        RECT 1.850 6.100 2.220 6.250 ;
        RECT 2.020 5.920 2.220 6.100 ;
        RECT 2.610 5.920 2.810 6.250 ;
        RECT 2.940 6.140 3.270 6.330 ;
        RECT 2.940 6.110 3.260 6.140 ;
        RECT 1.470 5.610 1.800 5.780 ;
        RECT 0.310 5.410 0.630 5.450 ;
        RECT 0.310 5.220 0.640 5.410 ;
        RECT 1.860 5.330 2.180 5.370 ;
        RECT 2.950 5.340 3.270 5.380 ;
        RECT 1.860 5.260 2.190 5.330 ;
        RECT 2.200 5.260 2.370 5.310 ;
        RECT 2.690 5.260 2.880 5.300 ;
        RECT 1.860 5.230 2.370 5.260 ;
        RECT 2.620 5.230 2.880 5.260 ;
        RECT 0.310 5.190 0.630 5.220 ;
        RECT 0.330 5.120 0.540 5.190 ;
        RECT 1.860 5.110 2.880 5.230 ;
        RECT 2.950 5.150 3.280 5.340 ;
        RECT 2.950 5.120 3.270 5.150 ;
        RECT 2.030 5.070 2.880 5.110 ;
        RECT 2.030 4.980 2.820 5.070 ;
        RECT 2.030 4.930 2.380 4.980 ;
        RECT 2.620 4.930 2.820 4.980 ;
        RECT 2.200 4.920 2.380 4.930 ;
        RECT 1.480 4.620 1.810 4.790 ;
        RECT 0.290 4.490 0.610 4.530 ;
        RECT 0.290 4.300 0.620 4.490 ;
        RECT 1.860 4.340 2.180 4.380 ;
        RECT 2.950 4.350 3.270 4.390 ;
        RECT 0.290 4.270 0.610 4.300 ;
        RECT 1.860 4.270 2.190 4.340 ;
        RECT 1.860 4.120 2.230 4.270 ;
        RECT 2.030 3.940 2.230 4.120 ;
        RECT 2.620 3.940 2.820 4.270 ;
        RECT 2.950 4.160 3.280 4.350 ;
        RECT 2.950 4.130 3.270 4.160 ;
        RECT 1.480 3.650 1.810 3.800 ;
        RECT 1.480 3.630 2.090 3.650 ;
        RECT 1.770 3.610 2.090 3.630 ;
        RECT 0.270 3.500 0.590 3.540 ;
        RECT 0.270 3.310 0.600 3.500 ;
        RECT 1.770 3.440 2.100 3.610 ;
        RECT 3.070 3.510 3.390 3.550 ;
        RECT 1.770 3.390 2.250 3.440 ;
        RECT 0.270 3.280 0.590 3.310 ;
        RECT 1.940 3.260 2.250 3.390 ;
        RECT 1.920 3.240 2.250 3.260 ;
        RECT 2.080 3.110 2.250 3.240 ;
        RECT 2.760 3.110 2.930 3.440 ;
        RECT 3.070 3.320 3.400 3.510 ;
        RECT 3.070 3.290 3.390 3.320 ;
        RECT 1.700 2.910 2.130 2.930 ;
        RECT 1.680 2.740 2.130 2.910 ;
        RECT 1.700 2.720 2.130 2.740 ;
        RECT 1.770 2.620 2.090 2.660 ;
        RECT 1.770 2.450 2.100 2.620 ;
        RECT 3.070 2.520 3.390 2.560 ;
        RECT 1.770 2.400 2.250 2.450 ;
        RECT 1.940 2.270 2.250 2.400 ;
        RECT 1.920 2.250 2.250 2.270 ;
        RECT 2.080 2.120 2.250 2.250 ;
        RECT 2.760 2.120 2.930 2.450 ;
        RECT 3.070 2.330 3.400 2.520 ;
        RECT 3.070 2.300 3.390 2.330 ;
        RECT 1.700 1.920 2.130 1.940 ;
        RECT 1.680 1.750 2.130 1.920 ;
        RECT 1.700 1.730 2.130 1.750 ;
        RECT 1.770 1.630 2.090 1.670 ;
        RECT 1.770 1.460 2.100 1.630 ;
        RECT 3.070 1.530 3.390 1.570 ;
        RECT 1.770 1.410 2.250 1.460 ;
        RECT 1.940 1.280 2.250 1.410 ;
        RECT 1.920 1.270 2.250 1.280 ;
        RECT 1.920 1.260 2.410 1.270 ;
        RECT 2.080 1.180 2.410 1.260 ;
        RECT 2.080 1.100 2.470 1.180 ;
        RECT 2.760 1.130 2.930 1.460 ;
        RECT 3.070 1.340 3.400 1.530 ;
        RECT 3.070 1.310 3.390 1.340 ;
        RECT 2.240 0.990 2.470 1.100 ;
        RECT 1.700 0.930 2.130 0.950 ;
        RECT 1.680 0.760 2.130 0.930 ;
        RECT 1.700 0.740 2.130 0.760 ;
      LAYER mcon ;
        RECT 1.910 6.140 2.080 6.310 ;
        RECT 3.000 6.150 3.170 6.320 ;
        RECT 0.370 5.230 0.540 5.400 ;
        RECT 1.920 5.150 2.090 5.320 ;
        RECT 2.700 5.100 2.870 5.270 ;
        RECT 3.010 5.160 3.180 5.330 ;
        RECT 0.350 4.310 0.520 4.480 ;
        RECT 1.920 4.160 2.090 4.330 ;
        RECT 3.010 4.170 3.180 4.340 ;
        RECT 0.330 3.320 0.500 3.490 ;
        RECT 1.830 3.430 2.000 3.600 ;
        RECT 3.130 3.330 3.300 3.500 ;
        RECT 1.830 2.440 2.000 2.610 ;
        RECT 3.130 2.340 3.300 2.510 ;
        RECT 1.830 1.450 2.000 1.620 ;
        RECT 2.270 1.000 2.440 1.170 ;
        RECT 3.130 1.350 3.300 1.520 ;
      LAYER met1 ;
        RECT 1.840 6.070 2.160 6.390 ;
        RECT 2.930 6.080 3.250 6.400 ;
        RECT 0.300 5.160 0.620 5.480 ;
        RECT 2.940 5.090 3.260 5.410 ;
        RECT 0.280 4.240 0.600 4.560 ;
        RECT 1.850 4.090 2.170 4.410 ;
        RECT 2.940 4.100 3.260 4.420 ;
        RECT 0.260 3.250 0.580 3.570 ;
        RECT 1.760 3.360 2.080 3.680 ;
        RECT 3.060 3.260 3.380 3.580 ;
        RECT 1.850 2.940 2.170 2.980 ;
        RECT 1.620 2.710 2.170 2.940 ;
        RECT 1.850 2.690 2.170 2.710 ;
        RECT 1.760 2.660 2.170 2.690 ;
        RECT 1.760 2.370 2.080 2.660 ;
        RECT 3.060 2.270 3.380 2.590 ;
        RECT 3.060 1.280 3.380 1.600 ;
        RECT 1.850 0.960 2.170 1.000 ;
        RECT 1.620 0.730 2.170 0.960 ;
        RECT 1.850 0.680 2.170 0.730 ;
      LAYER via ;
        RECT 1.870 6.100 2.130 6.360 ;
        RECT 2.960 6.110 3.220 6.370 ;
        RECT 0.330 5.190 0.590 5.450 ;
        RECT 2.970 5.120 3.230 5.380 ;
        RECT 0.310 4.270 0.570 4.530 ;
        RECT 1.880 4.120 2.140 4.380 ;
        RECT 2.970 4.130 3.230 4.390 ;
        RECT 0.290 3.280 0.550 3.540 ;
        RECT 1.790 3.390 2.050 3.650 ;
        RECT 3.090 3.290 3.350 3.550 ;
        RECT 1.880 2.690 2.140 2.950 ;
        RECT 1.790 2.400 2.050 2.660 ;
        RECT 3.090 2.300 3.350 2.560 ;
        RECT 3.090 1.310 3.350 1.570 ;
        RECT 1.880 0.710 2.140 0.970 ;
      LAYER met2 ;
        RECT 1.170 5.990 1.770 6.160 ;
        RECT 1.840 6.070 2.150 6.400 ;
        RECT 2.930 6.170 3.240 6.410 ;
        RECT 2.930 6.080 3.250 6.170 ;
        RECT 3.030 6.000 3.250 6.080 ;
        RECT 0.300 5.160 0.610 5.490 ;
        RECT 2.940 5.180 3.250 5.420 ;
        RECT 1.180 5.000 1.780 5.170 ;
        RECT 2.940 5.090 3.260 5.180 ;
        RECT 3.040 5.010 3.260 5.090 ;
        RECT 0.280 4.240 0.590 4.570 ;
        RECT 1.180 4.010 1.780 4.180 ;
        RECT 1.850 4.090 2.160 4.420 ;
        RECT 2.940 4.190 3.250 4.430 ;
        RECT 2.940 4.100 3.260 4.190 ;
        RECT 3.040 4.020 3.260 4.100 ;
        RECT 0.260 3.250 0.570 3.580 ;
        RECT 1.280 3.240 1.650 3.430 ;
        RECT 3.060 3.260 3.370 3.590 ;
        RECT 1.280 2.820 1.660 3.010 ;
        RECT 1.280 2.250 1.650 2.440 ;
        RECT 3.060 2.270 3.370 2.600 ;
        RECT 1.280 1.830 1.660 2.020 ;
        RECT 1.280 1.260 1.650 1.450 ;
        RECT 3.060 1.280 3.370 1.610 ;
        RECT 1.280 0.840 1.660 1.030 ;
  END
END sky130_hilas_Trans4small

MACRO sky130_hilas_FGBiasWeakGate2x1cell
  CLASS CORE ;
  FOREIGN sky130_hilas_FGBiasWeakGate2x1cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.540 BY 10.520 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DRAIN1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 5.840 9.120 6.020 ;
    END
  END DRAIN1
  PIN VIN11
    PORT
      LAYER met2 ;
        RECT 2.080 5.430 2.390 5.630 ;
        RECT 1.790 5.420 2.390 5.430 ;
        RECT 0.000 5.300 2.390 5.420 ;
        RECT 0.000 5.260 2.250 5.300 ;
        RECT 0.000 5.240 1.940 5.260 ;
    END
  END VIN11
  PIN ROW1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 9.340 5.000 9.650 5.220 ;
        RECT 9.340 4.990 11.530 5.000 ;
        RECT 0.000 4.780 11.530 4.990 ;
        RECT 0.000 4.770 10.220 4.780 ;
    END
  END ROW1
  PIN ROW2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 9.340 2.240 9.650 2.460 ;
        RECT 0.000 2.030 11.530 2.240 ;
        RECT 0.000 2.020 10.220 2.030 ;
    END
  END ROW2
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 11.010 0.470 11.290 6.520 ;
    END
  END VINJ
  PIN COLSEL1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 10.570 6.460 10.760 6.520 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.570 0.470 10.760 0.530 ;
    END
  END COLSEL1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2.830 5.550 3.060 6.520 ;
        RECT 2.830 5.300 3.070 5.550 ;
        RECT 2.830 3.660 3.060 5.300 ;
        RECT 2.830 3.370 3.160 3.660 ;
        RECT 2.830 0.470 3.060 3.370 ;
    END
  END VGND
  PIN GATE1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 4.050 0.470 4.280 6.520 ;
    END
  END GATE1
  PIN VTUN
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 0.350 0.480 0.770 6.520 ;
    END
  END VTUN
  PIN DRAIN2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 9.060 1.140 9.220 1.160 ;
        RECT 0.000 1.090 9.220 1.140 ;
        RECT 0.000 0.990 9.100 1.090 ;
    END
  END DRAIN2
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 1.500 1.950 1.710 ;
    END
  END VIN12
  PIN COMMONSOURCE
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 3.800 10.550 4.020 ;
        RECT 10.230 3.760 10.550 3.800 ;
    END
  END COMMONSOURCE
  OBS
      LAYER nwell ;
        RECT 14.520 10.180 16.250 10.520 ;
        RECT 14.500 8.620 16.250 10.180 ;
        RECT 14.500 6.990 16.230 8.620 ;
        RECT 12.980 6.600 16.290 6.990 ;
        RECT 12.980 6.560 16.530 6.600 ;
        RECT 12.980 4.910 16.540 6.560 ;
        RECT 0.590 1.870 1.150 4.290 ;
        RECT 12.980 3.820 16.290 4.910 ;
        RECT 12.980 1.980 16.290 3.170 ;
        RECT 12.980 0.330 16.540 1.980 ;
        RECT 12.980 0.290 16.530 0.330 ;
        RECT 12.980 0.000 16.290 0.290 ;
      LAYER li1 ;
        RECT 14.920 8.790 15.470 9.220 ;
        RECT 14.920 7.060 15.470 7.490 ;
        RECT 13.880 6.360 14.410 6.530 ;
        RECT 1.870 5.510 6.930 6.340 ;
        RECT 15.690 6.260 15.890 6.610 ;
        RECT 15.690 6.230 15.900 6.260 ;
        RECT 1.940 5.430 2.420 5.510 ;
        RECT 14.120 5.430 14.350 6.120 ;
        RECT 2.090 5.330 2.420 5.430 ;
        RECT 2.270 5.180 2.420 5.330 ;
        RECT 9.350 5.140 9.670 5.180 ;
        RECT 9.350 4.950 9.680 5.140 ;
        RECT 9.350 4.920 9.670 4.950 ;
        RECT 14.130 4.280 14.300 5.430 ;
        RECT 14.960 4.370 15.130 5.980 ;
        RECT 15.680 5.650 15.900 6.230 ;
        RECT 15.690 5.640 15.900 5.650 ;
        RECT 15.330 5.470 15.520 5.480 ;
        RECT 15.330 5.180 15.530 5.470 ;
        RECT 15.320 4.850 15.610 5.180 ;
        RECT 14.960 4.180 15.140 4.370 ;
        RECT 3.040 3.630 3.230 3.950 ;
        RECT 2.950 3.540 3.230 3.630 ;
        RECT 2.950 3.400 6.590 3.540 ;
        RECT 3.040 3.360 6.590 3.400 ;
        RECT 3.040 2.940 3.230 3.360 ;
        RECT 9.350 2.380 9.670 2.420 ;
        RECT 4.070 2.320 4.300 2.360 ;
        RECT 9.350 2.190 9.680 2.380 ;
        RECT 9.350 2.160 9.670 2.190 ;
        RECT 2.060 1.860 2.380 1.900 ;
        RECT 2.060 1.670 2.390 1.860 ;
        RECT 2.060 1.640 2.380 1.670 ;
        RECT 2.240 1.500 2.260 1.640 ;
        RECT 1.910 1.420 2.260 1.500 ;
        RECT 14.130 1.460 14.300 2.710 ;
        RECT 14.960 2.620 15.140 2.810 ;
        RECT 1.910 0.570 6.960 1.420 ;
        RECT 14.120 0.770 14.350 1.460 ;
        RECT 14.960 1.010 15.130 2.620 ;
        RECT 15.320 1.810 15.610 2.140 ;
        RECT 15.330 1.520 15.530 1.810 ;
        RECT 15.330 1.510 15.520 1.520 ;
        RECT 15.690 1.340 15.900 1.350 ;
        RECT 15.680 0.760 15.900 1.340 ;
        RECT 15.690 0.730 15.900 0.760 ;
        RECT 13.880 0.460 14.410 0.630 ;
        RECT 15.690 0.380 15.890 0.730 ;
      LAYER mcon ;
        RECT 14.920 8.870 15.190 9.140 ;
        RECT 14.920 7.140 15.190 7.410 ;
        RECT 2.150 5.370 2.320 5.540 ;
        RECT 14.150 5.910 14.320 6.080 ;
        RECT 15.700 6.060 15.870 6.230 ;
        RECT 14.150 5.460 14.320 5.630 ;
        RECT 9.410 4.960 9.580 5.130 ;
        RECT 15.340 5.220 15.520 5.410 ;
        RECT 2.960 3.430 3.130 3.600 ;
        RECT 9.410 2.200 9.580 2.370 ;
        RECT 2.120 1.680 2.290 1.850 ;
        RECT 14.150 1.260 14.320 1.430 ;
        RECT 15.340 1.580 15.520 1.770 ;
        RECT 14.150 0.810 14.320 0.980 ;
        RECT 15.700 0.760 15.870 0.930 ;
      LAYER met1 ;
        RECT 14.860 6.600 15.250 10.190 ;
        RECT 13.810 6.170 14.120 6.560 ;
        RECT 13.810 6.120 14.360 6.170 ;
        RECT 2.080 5.300 2.400 5.620 ;
        RECT 14.100 5.380 14.360 6.120 ;
        RECT 15.330 5.480 15.520 6.930 ;
        RECT 15.770 6.290 15.930 6.930 ;
        RECT 15.660 5.740 15.930 6.290 ;
        RECT 15.660 5.690 15.940 5.740 ;
        RECT 15.770 5.600 15.940 5.690 ;
        RECT 15.330 5.450 15.550 5.480 ;
        RECT 9.340 4.890 9.660 5.210 ;
        RECT 15.310 5.180 15.560 5.450 ;
        RECT 15.320 5.170 15.560 5.180 ;
        RECT 15.320 4.930 15.550 5.170 ;
        RECT 14.930 4.120 15.170 4.500 ;
        RECT 10.260 3.730 10.520 4.050 ;
        RECT 15.360 3.910 15.520 4.930 ;
        RECT 15.770 3.910 15.930 5.600 ;
        RECT 10.260 3.130 10.520 3.450 ;
        RECT 14.930 2.490 15.170 2.870 ;
        RECT 9.340 2.130 9.660 2.450 ;
        RECT 15.360 2.060 15.520 3.080 ;
        RECT 2.050 1.610 2.370 1.930 ;
        RECT 15.320 1.820 15.550 2.060 ;
        RECT 15.320 1.810 15.560 1.820 ;
        RECT 15.310 1.540 15.560 1.810 ;
        RECT 15.330 1.510 15.550 1.540 ;
        RECT 14.100 0.870 14.360 1.510 ;
        RECT 13.810 0.720 14.360 0.870 ;
        RECT 13.810 0.430 14.120 0.720 ;
        RECT 15.330 0.060 15.520 1.510 ;
        RECT 15.770 1.390 15.930 3.080 ;
        RECT 15.770 1.300 15.940 1.390 ;
        RECT 15.660 1.250 15.940 1.300 ;
        RECT 15.660 0.700 15.930 1.250 ;
        RECT 15.770 0.060 15.930 0.700 ;
      LAYER via ;
        RECT 13.840 6.150 14.100 6.410 ;
        RECT 2.110 5.330 2.370 5.590 ;
        RECT 9.370 4.920 9.630 5.180 ;
        RECT 10.260 3.760 10.520 4.020 ;
        RECT 10.260 3.160 10.520 3.420 ;
        RECT 9.370 2.160 9.630 2.420 ;
        RECT 2.080 1.640 2.340 1.900 ;
        RECT 13.840 0.580 14.100 0.840 ;
      LAYER met2 ;
        RECT 13.810 6.440 14.120 6.450 ;
        RECT 13.810 6.260 16.290 6.440 ;
        RECT 13.810 6.120 14.120 6.260 ;
        RECT 10.180 3.420 10.440 3.660 ;
        RECT 10.180 3.310 10.550 3.420 ;
        RECT 10.230 3.160 10.550 3.310 ;
        RECT 2.050 1.610 2.360 1.940 ;
        RECT 13.810 0.730 14.120 0.870 ;
        RECT 13.810 0.550 16.290 0.730 ;
        RECT 13.810 0.540 14.120 0.550 ;
  END
END sky130_hilas_FGBiasWeakGate2x1cell

MACRO sky130_hilas_swc4x2cell
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x2cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 45.720 BY 14.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 27.250 5.950 27.630 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.250 0.000 27.630 0.150 ;
    END
  END GATE2
  PIN VTUN
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 22.120 0.000 22.520 0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.200 0.000 23.600 0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.200 5.950 23.600 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 22.120 5.920 22.520 6.050 ;
    END
  END VTUN
  PIN GATE1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 18.090 5.950 18.470 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 18.090 0.000 18.470 0.090 ;
    END
  END GATE1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 32.400 0.010 32.560 0.070 ;
    END
  END VINJ
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 13.000 6.000 32.740 6.180 ;
        RECT 13.000 5.860 17.490 6.000 ;
        RECT 13.240 5.830 17.490 5.860 ;
        RECT 13.240 5.780 13.560 5.830 ;
        RECT 17.170 5.760 17.490 5.830 ;
        RECT 28.230 5.870 32.740 6.000 ;
        RECT 28.230 5.830 32.480 5.870 ;
        RECT 28.230 5.760 28.550 5.830 ;
        RECT 32.160 5.780 32.480 5.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.280 9.340 13.520 10.730 ;
        RECT 13.270 8.680 13.540 9.340 ;
        RECT 13.280 6.150 13.520 8.680 ;
        RECT 13.010 6.090 13.520 6.150 ;
        RECT 13.010 6.010 13.530 6.090 ;
        RECT 13.000 5.860 13.530 6.010 ;
        RECT 13.160 5.770 13.530 5.860 ;
        RECT 13.160 5.710 13.520 5.770 ;
        RECT 13.280 4.230 13.520 5.710 ;
      LAYER via ;
        RECT 13.040 6.060 13.300 6.140 ;
        RECT 13.040 5.880 13.530 6.060 ;
        RECT 13.270 5.800 13.530 5.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.160 0.000 13.320 0.060 ;
    END
  END VINJ
  PIN GATESELECT1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 13.570 6.000 13.760 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.570 0.010 13.760 0.070 ;
    END
  END GATESELECT1
  PIN GATESELECT2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 31.960 0.010 32.150 0.070 ;
    END
  END GATESELECT2
  PIN COL1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 13.970 6.000 14.130 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.970 0.010 14.130 0.070 ;
    END
  END COL1
  PIN COL2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 31.590 0.010 31.750 0.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.590 6.000 31.750 6.050 ;
    END
  END COL2
  PIN ROW1
    PORT
      LAYER met2 ;
        RECT 12.620 5.220 20.240 5.400 ;
        RECT 12.800 5.110 12.870 5.220 ;
    END
    PORT
      LAYER met2 ;
        RECT 25.480 5.220 33.100 5.400 ;
        RECT 32.830 5.110 32.920 5.220 ;
    END
  END ROW1
  PIN ROW2
    PORT
      LAYER met2 ;
        RECT 12.800 4.000 12.860 4.180 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.860 4.000 32.920 4.180 ;
    END
  END ROW2
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 12.800 5.540 12.860 5.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.830 5.540 32.920 5.720 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 12.800 3.570 12.930 3.750 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.860 3.570 32.920 3.750 ;
    END
  END DRAIN2
  PIN DRAIN3
    PORT
      LAYER met2 ;
        RECT 12.800 2.300 12.870 2.480 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.830 2.300 32.920 2.480 ;
    END
  END DRAIN3
  PIN ROW3
    PORT
      LAYER met2 ;
        RECT 12.800 1.870 12.870 2.050 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.830 1.870 32.920 2.050 ;
    END
  END ROW3
  PIN ROW4
    PORT
      LAYER met2 ;
        RECT 12.800 0.770 12.870 0.950 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.830 0.770 32.920 0.950 ;
    END
  END ROW4
  PIN DRAIN4
    PORT
      LAYER met2 ;
        RECT 12.800 0.340 12.870 0.520 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.830 0.340 32.920 0.520 ;
    END
  END DRAIN4
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 15.910 5.960 16.150 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.910 0.000 16.150 0.080 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.840 0.000 20.080 0.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.490 6.050 19.890 10.730 ;
        RECT 19.490 5.990 20.080 6.050 ;
        RECT 19.490 4.230 19.890 5.990 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.640 0.000 25.880 0.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.570 0.000 29.810 0.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.830 6.050 26.230 10.730 ;
        RECT 25.640 6.000 26.230 6.050 ;
        RECT 25.830 4.230 26.230 6.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.570 5.980 29.810 6.050 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 4.000 14.670 5.730 14.720 ;
        RECT 39.990 14.670 41.720 14.720 ;
        RECT 0.000 11.140 1.730 12.980 ;
        RECT 4.000 8.230 6.920 14.670 ;
        RECT 7.280 9.230 9.840 11.140 ;
        RECT 20.170 9.390 20.240 9.570 ;
        RECT 25.480 9.390 25.550 9.570 ;
        RECT 35.880 9.230 38.440 11.140 ;
        RECT 14.820 8.980 15.930 9.210 ;
        RECT 19.080 9.040 19.670 9.150 ;
        RECT 26.050 9.040 26.640 9.150 ;
        RECT 29.790 8.980 30.900 9.210 ;
        RECT 4.690 8.180 6.920 8.230 ;
        RECT 7.280 5.990 9.840 8.960 ;
        RECT 10.940 7.550 11.290 7.560 ;
        RECT 10.940 7.390 10.950 7.550 ;
        RECT 11.120 7.390 11.290 7.550 ;
        RECT 34.430 7.550 34.780 7.560 ;
        RECT 34.430 7.390 34.600 7.550 ;
        RECT 34.770 7.390 34.780 7.550 ;
        RECT 14.820 5.740 15.930 6.010 ;
        RECT 19.080 5.760 19.670 5.950 ;
        RECT 26.050 5.760 26.640 5.950 ;
        RECT 29.790 5.740 30.900 6.010 ;
        RECT 32.640 5.870 32.730 6.170 ;
        RECT 35.880 5.990 38.440 8.960 ;
        RECT 38.800 8.230 41.720 14.670 ;
        RECT 43.990 11.140 45.720 12.980 ;
        RECT 38.800 8.180 41.030 8.230 ;
        RECT 7.280 3.820 9.840 5.730 ;
        RECT 35.880 3.820 38.440 5.730 ;
        RECT 12.800 3.690 12.930 3.750 ;
        RECT 12.800 3.570 12.870 3.690 ;
      LAYER li1 ;
        RECT 0.760 11.590 1.310 12.020 ;
        RECT 4.790 11.660 5.340 12.090 ;
        RECT 40.380 11.660 40.930 12.090 ;
        RECT 44.410 11.590 44.960 12.020 ;
        RECT 9.280 10.790 9.600 10.830 ;
        RECT 7.680 10.400 7.880 10.750 ;
        RECT 9.270 10.670 9.600 10.790 ;
        RECT 9.160 10.570 9.600 10.670 ;
        RECT 36.120 10.790 36.440 10.830 ;
        RECT 36.120 10.670 36.450 10.790 ;
        RECT 36.120 10.570 36.560 10.670 ;
        RECT 9.160 10.500 9.500 10.570 ;
        RECT 36.220 10.500 36.560 10.570 ;
        RECT 7.670 10.370 7.880 10.400 ;
        RECT 37.840 10.400 38.040 10.750 ;
        RECT 7.670 9.780 7.890 10.370 ;
        RECT 8.410 9.780 8.610 10.380 ;
        RECT 9.280 10.240 9.600 10.280 ;
        RECT 9.270 10.050 9.600 10.240 ;
        RECT 9.160 10.020 9.600 10.050 ;
        RECT 36.120 10.240 36.440 10.280 ;
        RECT 36.120 10.050 36.450 10.240 ;
        RECT 36.120 10.020 36.560 10.050 ;
        RECT 9.160 9.880 9.500 10.020 ;
        RECT 36.220 9.880 36.560 10.020 ;
        RECT 37.110 9.780 37.310 10.380 ;
        RECT 37.840 10.370 38.050 10.400 ;
        RECT 37.830 9.780 38.050 10.370 ;
        RECT 13.310 8.740 13.480 9.270 ;
        RECT 17.250 8.750 17.420 9.280 ;
        RECT 28.300 8.750 28.470 9.280 ;
        RECT 32.240 8.740 32.410 9.270 ;
        RECT 7.670 7.820 7.890 8.410 ;
        RECT 7.670 7.790 7.880 7.820 ;
        RECT 8.410 7.810 8.610 8.410 ;
        RECT 9.160 8.170 9.500 8.310 ;
        RECT 36.220 8.170 36.560 8.310 ;
        RECT 9.160 8.140 9.600 8.170 ;
        RECT 9.270 7.950 9.600 8.140 ;
        RECT 36.120 8.140 36.560 8.170 ;
        RECT 9.280 7.910 9.600 7.950 ;
        RECT 7.680 7.160 7.880 7.790 ;
        RECT 9.160 7.620 9.500 7.690 ;
        RECT 9.160 7.520 9.600 7.620 ;
        RECT 9.270 7.430 9.600 7.520 ;
        RECT 9.160 7.330 9.600 7.430 ;
        RECT 10.940 7.390 11.380 7.560 ;
        RECT 9.160 7.260 9.500 7.330 ;
        RECT 7.670 7.130 7.880 7.160 ;
        RECT 7.670 6.540 7.890 7.130 ;
        RECT 8.410 6.540 8.610 7.140 ;
        RECT 9.280 7.000 9.600 7.040 ;
        RECT 9.270 6.810 9.600 7.000 ;
        RECT 13.310 6.900 13.480 7.910 ;
        RECT 17.240 7.040 17.410 8.050 ;
        RECT 28.310 7.040 28.480 8.050 ;
        RECT 36.120 7.950 36.450 8.140 ;
        RECT 36.120 7.910 36.440 7.950 ;
        RECT 32.240 6.900 32.410 7.910 ;
        RECT 37.110 7.810 37.310 8.410 ;
        RECT 37.830 7.820 38.050 8.410 ;
        RECT 37.840 7.790 38.050 7.820 ;
        RECT 36.220 7.620 36.560 7.690 ;
        RECT 34.340 7.390 34.780 7.560 ;
        RECT 36.120 7.520 36.560 7.620 ;
        RECT 36.120 7.430 36.450 7.520 ;
        RECT 36.120 7.330 36.560 7.430 ;
        RECT 36.220 7.260 36.560 7.330 ;
        RECT 37.840 7.160 38.040 7.790 ;
        RECT 36.120 7.000 36.440 7.040 ;
        RECT 9.160 6.780 9.600 6.810 ;
        RECT 36.120 6.810 36.450 7.000 ;
        RECT 36.120 6.780 36.560 6.810 ;
        RECT 9.160 6.640 9.500 6.780 ;
        RECT 36.220 6.640 36.560 6.780 ;
        RECT 37.110 6.540 37.310 7.140 ;
        RECT 37.840 7.130 38.050 7.160 ;
        RECT 37.830 6.540 38.050 7.130 ;
        RECT 7.670 4.590 7.890 5.180 ;
        RECT 7.670 4.560 7.880 4.590 ;
        RECT 8.410 4.580 8.610 5.180 ;
        RECT 9.160 4.940 9.500 5.080 ;
        RECT 36.220 4.940 36.560 5.080 ;
        RECT 9.160 4.910 9.600 4.940 ;
        RECT 9.270 4.720 9.600 4.910 ;
        RECT 9.280 4.680 9.600 4.720 ;
        RECT 36.120 4.910 36.560 4.940 ;
        RECT 36.120 4.720 36.450 4.910 ;
        RECT 36.120 4.680 36.440 4.720 ;
        RECT 37.110 4.580 37.310 5.180 ;
        RECT 37.830 4.590 38.050 5.180 ;
        RECT 7.680 4.210 7.880 4.560 ;
        RECT 37.840 4.560 38.050 4.590 ;
        RECT 9.160 4.390 9.500 4.460 ;
        RECT 36.220 4.390 36.560 4.460 ;
        RECT 9.160 4.290 9.600 4.390 ;
        RECT 9.270 4.170 9.600 4.290 ;
        RECT 9.280 4.130 9.600 4.170 ;
        RECT 36.120 4.290 36.560 4.390 ;
        RECT 36.120 4.170 36.450 4.290 ;
        RECT 37.840 4.210 38.040 4.560 ;
        RECT 36.120 4.130 36.440 4.170 ;
      LAYER mcon ;
        RECT 1.040 11.670 1.310 11.940 ;
        RECT 5.070 11.740 5.340 12.010 ;
        RECT 40.380 11.740 40.650 12.010 ;
        RECT 44.410 11.670 44.680 11.940 ;
        RECT 9.370 10.610 9.540 10.780 ;
        RECT 36.180 10.610 36.350 10.780 ;
        RECT 7.700 10.200 7.870 10.370 ;
        RECT 8.430 10.170 8.600 10.340 ;
        RECT 9.370 10.060 9.540 10.230 ;
        RECT 36.180 10.060 36.350 10.230 ;
        RECT 37.120 10.170 37.290 10.340 ;
        RECT 37.850 10.200 38.020 10.370 ;
        RECT 13.310 9.100 13.480 9.270 ;
        RECT 17.250 9.110 17.420 9.280 ;
        RECT 28.300 9.110 28.470 9.280 ;
        RECT 32.240 9.100 32.410 9.270 ;
        RECT 7.700 7.820 7.870 7.990 ;
        RECT 8.430 7.850 8.600 8.020 ;
        RECT 9.370 7.960 9.540 8.130 ;
        RECT 9.370 7.370 9.540 7.580 ;
        RECT 13.310 7.510 13.480 7.680 ;
        RECT 13.310 7.150 13.480 7.320 ;
        RECT 7.700 6.960 7.870 7.130 ;
        RECT 8.430 6.930 8.600 7.100 ;
        RECT 9.370 6.820 9.540 6.990 ;
        RECT 17.240 7.650 17.410 7.820 ;
        RECT 17.240 7.290 17.410 7.460 ;
        RECT 36.180 7.960 36.350 8.130 ;
        RECT 28.310 7.650 28.480 7.820 ;
        RECT 28.310 7.290 28.480 7.460 ;
        RECT 37.120 7.850 37.290 8.020 ;
        RECT 37.850 7.820 38.020 7.990 ;
        RECT 32.240 7.510 32.410 7.680 ;
        RECT 34.600 7.390 34.780 7.560 ;
        RECT 36.180 7.370 36.350 7.580 ;
        RECT 32.240 7.150 32.410 7.320 ;
        RECT 36.180 6.820 36.350 6.990 ;
        RECT 37.120 6.930 37.290 7.100 ;
        RECT 37.850 6.960 38.020 7.130 ;
        RECT 7.700 4.590 7.870 4.760 ;
        RECT 8.430 4.620 8.600 4.790 ;
        RECT 9.370 4.730 9.540 4.900 ;
        RECT 36.180 4.730 36.350 4.900 ;
        RECT 37.120 4.620 37.290 4.790 ;
        RECT 37.850 4.590 38.020 4.760 ;
        RECT 9.370 4.180 9.540 4.350 ;
        RECT 36.180 4.180 36.350 4.350 ;
      LAYER met1 ;
        RECT 0.980 11.130 1.370 12.990 ;
        RECT 5.010 11.200 5.400 13.060 ;
        RECT 5.890 8.180 6.270 14.680 ;
        RECT 7.640 10.430 7.800 11.130 ;
        RECT 7.640 9.880 7.910 10.430 ;
        RECT 7.630 9.830 7.910 9.880 ;
        RECT 8.050 10.090 8.240 11.080 ;
        RECT 8.450 10.400 8.610 11.130 ;
        RECT 9.290 10.540 9.610 10.860 ;
        RECT 10.530 10.450 10.690 10.500 ;
        RECT 10.940 10.450 11.130 10.500 ;
        RECT 11.340 10.460 11.500 10.500 ;
        RECT 15.460 10.400 15.840 10.730 ;
        RECT 8.410 10.380 8.610 10.400 ;
        RECT 8.400 10.140 8.630 10.380 ;
        RECT 8.400 10.090 8.610 10.140 ;
        RECT 8.050 9.970 8.220 10.090 ;
        RECT 7.630 9.740 7.800 9.830 ;
        RECT 7.640 9.230 7.800 9.740 ;
        RECT 8.050 9.230 8.210 9.970 ;
        RECT 8.450 9.230 8.610 10.090 ;
        RECT 9.290 9.990 9.610 10.310 ;
        RECT 17.210 9.320 17.450 10.730 ;
        RECT 28.270 9.320 28.510 10.730 ;
        RECT 29.880 10.400 30.260 10.730 ;
        RECT 32.200 9.340 32.440 10.730 ;
        RECT 36.110 10.540 36.430 10.860 ;
        RECT 34.220 10.460 34.380 10.500 ;
        RECT 34.590 10.450 34.780 10.500 ;
        RECT 35.030 10.450 35.190 10.500 ;
        RECT 37.110 10.400 37.270 11.130 ;
        RECT 37.110 10.380 37.310 10.400 ;
        RECT 36.110 9.990 36.430 10.310 ;
        RECT 37.090 10.140 37.320 10.380 ;
        RECT 37.110 10.090 37.320 10.140 ;
        RECT 37.480 10.090 37.670 11.080 ;
        RECT 37.920 10.430 38.080 11.130 ;
        RECT 7.640 8.450 7.800 8.960 ;
        RECT 7.630 8.360 7.800 8.450 ;
        RECT 7.630 8.310 7.910 8.360 ;
        RECT 7.640 7.760 7.910 8.310 ;
        RECT 8.050 8.220 8.210 8.960 ;
        RECT 8.050 8.100 8.220 8.220 ;
        RECT 8.450 8.100 8.610 8.960 ;
        RECT 17.200 8.660 17.460 9.320 ;
        RECT 28.260 8.660 28.520 9.320 ;
        RECT 32.180 8.680 32.450 9.340 ;
        RECT 37.110 9.230 37.270 10.090 ;
        RECT 37.500 9.970 37.670 10.090 ;
        RECT 37.510 9.230 37.670 9.970 ;
        RECT 37.810 9.880 38.080 10.430 ;
        RECT 37.810 9.830 38.090 9.880 ;
        RECT 37.920 9.740 38.090 9.830 ;
        RECT 37.920 9.230 38.080 9.740 ;
        RECT 7.640 7.190 7.800 7.760 ;
        RECT 7.640 6.640 7.910 7.190 ;
        RECT 7.630 6.590 7.910 6.640 ;
        RECT 8.050 6.850 8.240 8.100 ;
        RECT 8.400 8.050 8.610 8.100 ;
        RECT 8.400 7.810 8.630 8.050 ;
        RECT 9.290 7.880 9.610 8.200 ;
        RECT 8.410 7.790 8.610 7.810 ;
        RECT 8.450 7.160 8.610 7.790 ;
        RECT 9.290 7.300 9.610 7.650 ;
        RECT 10.940 7.590 11.070 7.610 ;
        RECT 10.910 7.570 11.150 7.590 ;
        RECT 10.910 7.380 11.350 7.570 ;
        RECT 10.910 7.360 11.150 7.380 ;
        RECT 10.940 7.320 11.050 7.360 ;
        RECT 8.410 7.140 8.610 7.160 ;
        RECT 8.400 6.900 8.630 7.140 ;
        RECT 8.400 6.850 8.610 6.900 ;
        RECT 8.050 6.730 8.220 6.850 ;
        RECT 7.630 6.500 7.800 6.590 ;
        RECT 7.640 5.990 7.800 6.500 ;
        RECT 8.050 5.990 8.210 6.730 ;
        RECT 8.450 5.990 8.610 6.850 ;
        RECT 9.290 6.750 9.610 7.070 ;
        RECT 17.210 6.050 17.450 8.660 ;
        RECT 28.270 6.050 28.510 8.660 ;
        RECT 32.200 6.160 32.440 8.680 ;
        RECT 36.110 7.880 36.430 8.200 ;
        RECT 37.110 8.100 37.270 8.960 ;
        RECT 37.510 8.220 37.670 8.960 ;
        RECT 37.920 8.450 38.080 8.960 ;
        RECT 37.920 8.360 38.090 8.450 ;
        RECT 37.500 8.100 37.670 8.220 ;
        RECT 37.110 8.050 37.320 8.100 ;
        RECT 37.090 7.810 37.320 8.050 ;
        RECT 37.110 7.790 37.310 7.810 ;
        RECT 34.650 7.590 34.780 7.610 ;
        RECT 34.570 7.570 34.810 7.590 ;
        RECT 34.370 7.380 34.810 7.570 ;
        RECT 34.570 7.360 34.810 7.380 ;
        RECT 34.670 7.320 34.780 7.360 ;
        RECT 36.110 7.300 36.430 7.650 ;
        RECT 37.110 7.160 37.270 7.790 ;
        RECT 37.110 7.140 37.310 7.160 ;
        RECT 36.110 6.750 36.430 7.070 ;
        RECT 37.090 6.900 37.320 7.140 ;
        RECT 37.110 6.850 37.320 6.900 ;
        RECT 37.480 6.850 37.670 8.100 ;
        RECT 37.810 8.310 38.090 8.360 ;
        RECT 37.810 7.760 38.080 8.310 ;
        RECT 39.450 8.180 39.830 14.680 ;
        RECT 40.320 11.200 40.710 13.060 ;
        RECT 44.350 11.130 44.740 12.990 ;
        RECT 37.920 7.190 38.080 7.760 ;
        RECT 32.200 6.090 32.730 6.160 ;
        RECT 17.200 5.730 17.460 6.050 ;
        RECT 7.640 5.220 7.800 5.730 ;
        RECT 7.630 5.130 7.800 5.220 ;
        RECT 7.630 5.080 7.910 5.130 ;
        RECT 7.640 4.530 7.910 5.080 ;
        RECT 8.050 4.990 8.210 5.730 ;
        RECT 8.050 4.870 8.220 4.990 ;
        RECT 8.450 4.870 8.610 5.730 ;
        RECT 7.640 3.830 7.800 4.530 ;
        RECT 8.050 3.880 8.240 4.870 ;
        RECT 8.400 4.820 8.610 4.870 ;
        RECT 8.400 4.580 8.630 4.820 ;
        RECT 9.290 4.650 9.610 4.970 ;
        RECT 8.410 4.560 8.610 4.580 ;
        RECT 8.450 3.830 8.610 4.560 ;
        RECT 9.290 4.100 9.610 4.420 ;
        RECT 15.460 4.230 15.840 4.830 ;
        RECT 17.210 4.230 17.450 5.730 ;
        RECT 22.520 5.690 23.200 5.910 ;
        RECT 28.260 5.730 28.520 6.050 ;
        RECT 31.960 6.000 32.150 6.050 ;
        RECT 32.190 5.880 32.730 6.090 ;
        RECT 37.110 5.990 37.270 6.850 ;
        RECT 37.500 6.730 37.670 6.850 ;
        RECT 37.510 5.990 37.670 6.730 ;
        RECT 37.810 6.640 38.080 7.190 ;
        RECT 37.810 6.590 38.090 6.640 ;
        RECT 37.920 6.500 38.090 6.590 ;
        RECT 37.920 5.990 38.080 6.500 ;
        RECT 32.190 5.770 32.560 5.880 ;
        RECT 28.270 4.230 28.510 5.730 ;
        RECT 32.200 5.710 32.560 5.770 ;
        RECT 29.880 4.230 30.260 4.830 ;
        RECT 32.200 4.230 32.440 5.710 ;
        RECT 36.110 4.650 36.430 4.970 ;
        RECT 37.110 4.870 37.270 5.730 ;
        RECT 37.510 4.990 37.670 5.730 ;
        RECT 37.920 5.220 38.080 5.730 ;
        RECT 37.920 5.130 38.090 5.220 ;
        RECT 37.500 4.870 37.670 4.990 ;
        RECT 37.110 4.820 37.320 4.870 ;
        RECT 37.090 4.580 37.320 4.820 ;
        RECT 37.110 4.560 37.310 4.580 ;
        RECT 36.110 4.100 36.430 4.420 ;
        RECT 37.110 3.830 37.270 4.560 ;
        RECT 37.480 3.880 37.670 4.870 ;
        RECT 37.810 5.080 38.090 5.130 ;
        RECT 37.810 4.530 38.080 5.080 ;
        RECT 37.920 3.830 38.080 4.530 ;
      LAYER via ;
        RECT 9.320 10.570 9.580 10.830 ;
        RECT 9.320 10.020 9.580 10.280 ;
        RECT 36.140 10.570 36.400 10.830 ;
        RECT 36.140 10.020 36.400 10.280 ;
        RECT 9.320 7.910 9.580 8.170 ;
        RECT 9.320 7.330 9.580 7.620 ;
        RECT 9.320 6.780 9.580 7.040 ;
        RECT 36.140 7.910 36.400 8.170 ;
        RECT 36.140 7.330 36.400 7.620 ;
        RECT 36.140 6.780 36.400 7.040 ;
        RECT 32.440 6.060 32.700 6.150 ;
        RECT 17.200 5.760 17.460 6.020 ;
        RECT 9.320 4.680 9.580 4.940 ;
        RECT 9.320 4.130 9.580 4.390 ;
        RECT 28.260 5.760 28.520 6.020 ;
        RECT 32.190 5.890 32.700 6.060 ;
        RECT 32.190 5.800 32.450 5.890 ;
        RECT 36.140 4.680 36.400 4.940 ;
        RECT 36.140 4.130 36.400 4.390 ;
      LAYER met2 ;
        RECT 9.300 10.580 9.610 10.870 ;
        RECT 7.280 10.540 9.610 10.580 ;
        RECT 36.110 10.580 36.420 10.870 ;
        RECT 36.110 10.540 38.440 10.580 ;
        RECT 7.280 10.400 9.460 10.540 ;
        RECT 36.260 10.400 38.440 10.540 ;
        RECT 9.300 10.150 9.610 10.320 ;
        RECT 7.280 9.990 9.610 10.150 ;
        RECT 7.280 9.970 9.450 9.990 ;
        RECT 9.750 9.970 9.840 10.150 ;
        RECT 12.610 9.990 20.240 10.170 ;
        RECT 25.480 9.990 33.110 10.170 ;
        RECT 36.110 10.150 36.420 10.320 ;
        RECT 35.880 9.970 35.970 10.150 ;
        RECT 36.110 9.990 38.440 10.150 ;
        RECT 36.270 9.970 38.440 9.990 ;
        RECT 12.610 9.550 20.240 9.730 ;
        RECT 25.480 9.550 33.110 9.730 ;
        RECT 12.610 8.450 20.240 8.630 ;
        RECT 25.480 8.450 33.110 8.630 ;
        RECT 7.280 8.200 9.450 8.220 ;
        RECT 7.280 8.040 9.610 8.200 ;
        RECT 9.750 8.040 9.840 8.220 ;
        RECT 9.300 7.870 9.610 8.040 ;
        RECT 12.610 8.020 20.240 8.200 ;
        RECT 25.480 8.020 33.110 8.200 ;
        RECT 35.880 8.040 35.970 8.220 ;
        RECT 36.270 8.200 38.440 8.220 ;
        RECT 36.110 8.040 38.440 8.200 ;
        RECT 36.110 7.870 36.420 8.040 ;
        RECT 7.280 7.650 9.460 7.790 ;
        RECT 36.260 7.650 38.440 7.790 ;
        RECT 7.280 7.610 9.610 7.650 ;
        RECT 9.300 7.340 9.610 7.610 ;
        RECT 7.280 7.300 9.610 7.340 ;
        RECT 36.110 7.610 38.440 7.650 ;
        RECT 36.110 7.340 36.420 7.610 ;
        RECT 36.110 7.300 38.440 7.340 ;
        RECT 7.280 7.160 9.460 7.300 ;
        RECT 36.260 7.160 38.440 7.300 ;
        RECT 9.300 6.910 9.610 7.080 ;
        RECT 7.280 6.750 9.610 6.910 ;
        RECT 7.280 6.730 9.450 6.750 ;
        RECT 9.750 6.730 9.840 6.910 ;
        RECT 12.620 6.750 20.240 6.930 ;
        RECT 25.480 6.750 33.100 6.930 ;
        RECT 36.110 6.910 36.420 7.080 ;
        RECT 35.880 6.730 35.970 6.910 ;
        RECT 36.110 6.750 38.440 6.910 ;
        RECT 36.270 6.730 38.440 6.750 ;
        RECT 12.610 6.320 20.240 6.500 ;
        RECT 25.480 6.320 33.110 6.500 ;
        RECT 7.280 4.970 9.450 4.990 ;
        RECT 7.280 4.810 9.610 4.970 ;
        RECT 9.750 4.810 9.840 4.990 ;
        RECT 9.300 4.640 9.610 4.810 ;
        RECT 12.640 4.800 20.240 4.970 ;
        RECT 25.480 4.800 33.080 4.970 ;
        RECT 35.880 4.810 35.970 4.990 ;
        RECT 36.270 4.970 38.440 4.990 ;
        RECT 36.110 4.810 38.440 4.970 ;
        RECT 36.110 4.640 36.420 4.810 ;
        RECT 7.280 4.420 9.460 4.560 ;
        RECT 36.260 4.420 38.440 4.560 ;
        RECT 7.280 4.380 9.610 4.420 ;
        RECT 9.300 4.090 9.610 4.380 ;
        RECT 36.110 4.380 38.440 4.420 ;
        RECT 36.110 4.090 36.420 4.380 ;
        RECT 19.500 1.380 26.260 1.560 ;
  END
END sky130_hilas_swc4x2cell

MACRO sky130_hilas_polyresistorGND
  CLASS CORE ;
  FOREIGN sky130_hilas_polyresistorGND ;
  ORIGIN 0.000 0.000 ;
  SIZE 55.470 BY 10.890 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN INPUT
    PORT
      LAYER met1 ;
        RECT 21.060 10.250 23.470 10.890 ;
        RECT 21.080 8.900 21.490 10.250 ;
    END
  END INPUT
  PIN OUTPUT
    ANTENNADIFFAREA 16.452000 ;
    PORT
      LAYER met2 ;
        RECT 0.000 7.380 55.470 8.770 ;
    END
  END OUTPUT
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 27.810 9.590 28.220 10.360 ;
        RECT 27.540 9.320 28.220 9.590 ;
        RECT 27.540 8.890 29.230 9.320 ;
        RECT 0.330 8.710 24.700 8.730 ;
        RECT 0.270 8.320 24.700 8.710 ;
        RECT 0.270 0.070 0.680 8.320 ;
        RECT 26.870 0.820 29.230 8.890 ;
        RECT 33.500 8.720 54.860 8.730 ;
        RECT 33.440 8.330 54.860 8.720 ;
        RECT 33.440 8.320 54.700 8.330 ;
        RECT 26.750 0.000 29.230 0.820 ;
      LAYER via ;
        RECT 0.820 8.410 24.620 8.670 ;
        RECT 33.500 8.410 54.360 8.670 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 21.140 9.120 21.360 10.240 ;
        RECT 21.090 8.930 21.420 9.120 ;
        RECT 27.880 8.930 28.120 10.280 ;
        RECT 0.380 8.460 55.120 8.730 ;
        RECT 0.380 8.330 24.720 8.460 ;
        RECT 33.410 8.330 55.120 8.460 ;
        RECT 0.380 0.730 0.550 8.330 ;
        RECT 54.950 1.250 55.120 8.330 ;
        RECT 26.820 0.390 29.180 0.560 ;
      LAYER mcon ;
        RECT 21.170 10.040 21.340 10.210 ;
        RECT 21.170 9.680 21.340 9.850 ;
        RECT 21.170 9.320 21.340 9.490 ;
        RECT 21.170 8.960 21.340 9.130 ;
        RECT 27.920 9.870 28.090 10.040 ;
        RECT 27.920 9.510 28.090 9.680 ;
        RECT 27.920 9.150 28.090 9.320 ;
        RECT 0.720 8.350 24.620 8.520 ;
        RECT 33.500 8.350 54.670 8.520 ;
        RECT 27.190 0.390 27.360 0.560 ;
        RECT 27.560 0.390 27.730 0.560 ;
        RECT 27.920 0.390 28.090 0.560 ;
        RECT 28.280 0.390 28.450 0.560 ;
        RECT 28.640 0.390 28.820 0.560 ;
        RECT 29.010 0.390 29.180 0.560 ;
      LAYER met2 ;
        RECT 0.000 1.080 55.470 2.480 ;
  END
END sky130_hilas_polyresistorGND

MACRO sky130_hilas_swc4x2cellOverlap
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x2cellOverlap ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.570 BY 10.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VERT1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 5.970 5.990 6.130 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.970 0.010 6.130 0.080 ;
    END
  END VERT1
  PIN HORIZ1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.800 4.940 4.880 5.120 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.670 4.940 22.780 5.120 ;
    END
  END HORIZ1
  PIN DRAIN1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.800 5.370 4.880 5.550 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.660 5.370 22.770 5.550 ;
    END
  END DRAIN1
  PIN HORIZ2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.800 3.940 4.880 4.120 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.670 3.940 22.780 4.120 ;
    END
  END HORIZ2
  PIN DRAIN2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.800 3.510 4.880 3.690 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.670 3.510 22.780 3.690 ;
    END
  END DRAIN2
  PIN DRAIN3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.800 2.360 4.870 2.540 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.660 2.360 22.770 2.540 ;
    END
  END DRAIN3
  PIN HORIZ3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.800 1.930 4.870 2.110 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.660 1.930 22.770 2.110 ;
    END
  END HORIZ3
  PIN HORIZ4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.800 0.940 4.870 1.120 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.660 0.940 22.770 1.120 ;
    END
  END HORIZ4
  PIN DRAIN4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.800 0.510 4.870 0.690 ;
    END
  END DRAIN4
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 5.160 5.990 5.320 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.160 0.010 5.320 0.080 ;
    END
    PORT
      LAYER met1 ;
        RECT 22.250 0.010 22.410 0.080 ;
    END
    PORT
      LAYER met1 ;
        RECT 22.250 5.980 22.410 6.050 ;
    END
  END VINJ
  PIN GATESELECT1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 5.570 5.990 5.760 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.570 0.010 5.760 0.080 ;
    END
  END GATESELECT1
  PIN VERT2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 21.440 5.980 21.600 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.440 0.010 21.600 0.080 ;
    END
  END VERT2
  PIN GATESELECT2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 21.810 5.980 22.000 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.810 0.010 22.000 0.080 ;
    END
  END GATESELECT2
  PIN DRAIN
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 22.660 0.510 22.770 0.690 ;
    END
  END DRAIN
  PIN GATE2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 18.090 0.000 18.330 6.050 ;
    END
  END GATE2
  PIN GATE1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 9.240 0.000 9.490 6.050 ;
    END
  END GATE1
  PIN VTUN
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 12.850 0.000 13.150 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 14.430 0.000 14.730 6.050 ;
    END
  END VTUN
  OBS
      LAYER nwell ;
        RECT 0.240 10.800 4.240 10.870 ;
        RECT 0.000 8.890 4.240 10.800 ;
        RECT 0.240 8.730 4.240 8.890 ;
        RECT 0.000 5.880 4.240 8.730 ;
        RECT 0.240 5.730 4.240 5.880 ;
        RECT 0.000 4.820 4.240 5.730 ;
        RECT 23.330 10.800 27.330 10.870 ;
        RECT 23.330 8.890 27.570 10.800 ;
        RECT 23.330 8.730 27.330 8.890 ;
        RECT 23.330 5.880 27.570 8.730 ;
        RECT 23.330 5.730 27.330 5.880 ;
        RECT 23.330 4.820 27.570 5.730 ;
        RECT 0.000 3.820 2.560 4.820 ;
        RECT 25.010 3.820 27.570 4.820 ;
      LAYER li1 ;
        RECT 0.580 10.410 3.890 10.540 ;
        RECT 0.400 10.060 3.890 10.410 ;
        RECT 0.390 9.560 3.890 10.060 ;
        RECT 0.390 9.440 0.610 9.560 ;
        RECT 1.130 9.440 1.330 9.560 ;
        RECT 1.880 9.540 2.220 9.560 ;
        RECT 10.390 9.550 10.560 10.440 ;
        RECT 17.010 9.550 17.180 10.440 ;
        RECT 23.680 10.410 26.990 10.540 ;
        RECT 23.680 10.060 27.170 10.410 ;
        RECT 23.680 9.560 27.180 10.060 ;
        RECT 25.350 9.540 25.690 9.560 ;
        RECT 26.240 9.440 26.440 9.560 ;
        RECT 26.960 9.440 27.180 9.560 ;
        RECT 0.580 8.180 3.890 9.070 ;
        RECT 0.390 8.090 3.890 8.180 ;
        RECT 0.390 7.600 0.610 8.090 ;
        RECT 1.130 7.600 1.330 8.090 ;
        RECT 1.880 7.940 2.220 8.080 ;
        RECT 10.390 8.030 10.560 8.920 ;
        RECT 17.010 8.030 17.180 8.920 ;
        RECT 23.680 8.180 26.990 9.070 ;
        RECT 23.680 8.090 27.180 8.180 ;
        RECT 25.350 7.940 25.690 8.080 ;
        RECT 1.880 7.910 2.320 7.940 ;
        RECT 1.990 7.720 2.320 7.910 ;
        RECT 2.000 7.680 2.320 7.720 ;
        RECT 25.250 7.910 25.690 7.940 ;
        RECT 25.250 7.720 25.580 7.910 ;
        RECT 25.250 7.680 25.570 7.720 ;
        RECT 26.240 7.600 26.440 8.090 ;
        RECT 26.960 7.600 27.180 8.090 ;
        RECT 0.390 7.560 3.890 7.600 ;
        RECT 0.400 7.390 3.890 7.560 ;
        RECT 23.680 7.560 27.180 7.600 ;
        RECT 0.400 7.220 4.100 7.390 ;
        RECT 0.400 7.050 3.890 7.220 ;
        RECT 0.390 6.620 3.890 7.050 ;
        RECT 0.390 6.430 0.610 6.620 ;
        RECT 1.130 6.430 1.330 6.620 ;
        RECT 1.880 6.530 2.220 6.620 ;
        RECT 10.390 6.580 10.560 7.470 ;
        RECT 17.010 6.580 17.180 7.470 ;
        RECT 23.680 7.390 27.170 7.560 ;
        RECT 23.470 7.220 27.170 7.390 ;
        RECT 23.680 7.050 27.170 7.220 ;
        RECT 23.680 6.620 27.180 7.050 ;
        RECT 25.350 6.530 25.690 6.620 ;
        RECT 26.240 6.430 26.440 6.620 ;
        RECT 26.960 6.430 27.180 6.620 ;
        RECT 0.580 5.180 3.890 6.130 ;
        RECT 0.390 5.150 3.890 5.180 ;
        RECT 0.390 4.590 0.610 5.150 ;
        RECT 0.390 4.560 0.600 4.590 ;
        RECT 1.130 4.580 1.330 5.150 ;
        RECT 1.880 4.940 2.220 5.080 ;
        RECT 10.390 5.040 10.560 5.930 ;
        RECT 17.010 5.040 17.180 5.930 ;
        RECT 23.680 5.180 26.990 6.130 ;
        RECT 23.680 5.150 27.180 5.180 ;
        RECT 25.350 4.940 25.690 5.080 ;
        RECT 1.880 4.910 2.320 4.940 ;
        RECT 1.990 4.720 2.320 4.910 ;
        RECT 2.000 4.680 2.320 4.720 ;
        RECT 25.250 4.910 25.690 4.940 ;
        RECT 25.250 4.720 25.580 4.910 ;
        RECT 25.250 4.680 25.570 4.720 ;
        RECT 26.240 4.580 26.440 5.150 ;
        RECT 26.960 4.590 27.180 5.150 ;
        RECT 0.400 4.210 0.600 4.560 ;
        RECT 26.970 4.560 27.180 4.590 ;
        RECT 1.880 4.390 2.220 4.460 ;
        RECT 25.350 4.390 25.690 4.460 ;
        RECT 1.880 4.290 2.320 4.390 ;
        RECT 1.990 4.170 2.320 4.290 ;
        RECT 2.000 4.130 2.320 4.170 ;
        RECT 25.250 4.290 25.690 4.390 ;
        RECT 25.250 4.170 25.580 4.290 ;
        RECT 26.970 4.210 27.170 4.560 ;
        RECT 25.250 4.130 25.570 4.170 ;
      LAYER mcon ;
        RECT 2.150 10.440 2.320 10.480 ;
        RECT 2.090 10.310 2.320 10.440 ;
        RECT 2.090 10.270 2.260 10.310 ;
        RECT 0.420 9.860 0.590 10.030 ;
        RECT 1.150 9.830 1.320 10.000 ;
        RECT 2.090 9.790 2.260 9.890 ;
        RECT 2.090 9.720 2.320 9.790 ;
        RECT 2.150 9.620 2.320 9.720 ;
        RECT 10.390 10.240 10.560 10.410 ;
        RECT 17.010 10.240 17.180 10.410 ;
        RECT 25.250 10.440 25.420 10.480 ;
        RECT 25.250 10.310 25.480 10.440 ;
        RECT 25.310 10.270 25.480 10.310 ;
        RECT 25.310 9.790 25.480 9.890 ;
        RECT 26.250 9.830 26.420 10.000 ;
        RECT 26.980 9.860 27.150 10.030 ;
        RECT 25.250 9.720 25.480 9.790 ;
        RECT 25.250 9.620 25.420 9.720 ;
        RECT 2.150 8.840 2.320 9.010 ;
        RECT 2.150 8.150 2.320 8.320 ;
        RECT 10.390 8.720 10.560 8.890 ;
        RECT 0.420 7.590 0.590 7.760 ;
        RECT 17.010 8.720 17.180 8.890 ;
        RECT 25.250 8.840 25.420 9.010 ;
        RECT 25.250 8.150 25.420 8.320 ;
        RECT 1.150 7.620 1.320 7.790 ;
        RECT 2.090 7.730 2.260 7.900 ;
        RECT 25.310 7.730 25.480 7.900 ;
        RECT 26.250 7.620 26.420 7.790 ;
        RECT 2.150 7.430 2.320 7.540 ;
        RECT 2.090 7.370 2.320 7.430 ;
        RECT 26.980 7.590 27.150 7.760 ;
        RECT 2.090 7.180 2.260 7.370 ;
        RECT 3.660 7.220 3.840 7.390 ;
        RECT 10.390 7.270 10.560 7.440 ;
        RECT 0.420 6.850 0.590 7.020 ;
        RECT 1.150 6.820 1.320 6.990 ;
        RECT 2.090 6.850 2.260 6.880 ;
        RECT 2.090 6.710 2.320 6.850 ;
        RECT 2.150 6.680 2.320 6.710 ;
        RECT 17.010 7.270 17.180 7.440 ;
        RECT 25.250 7.430 25.420 7.540 ;
        RECT 23.730 7.220 23.910 7.390 ;
        RECT 25.250 7.370 25.480 7.430 ;
        RECT 25.310 7.180 25.480 7.370 ;
        RECT 25.310 6.850 25.480 6.880 ;
        RECT 25.250 6.710 25.480 6.850 ;
        RECT 26.250 6.820 26.420 6.990 ;
        RECT 26.980 6.850 27.150 7.020 ;
        RECT 25.250 6.680 25.420 6.710 ;
        RECT 2.150 5.900 2.320 6.070 ;
        RECT 2.150 5.210 2.320 5.380 ;
        RECT 10.390 5.730 10.560 5.900 ;
        RECT 0.420 4.590 0.590 4.760 ;
        RECT 17.010 5.730 17.180 5.900 ;
        RECT 25.250 5.900 25.420 6.070 ;
        RECT 25.250 5.210 25.420 5.380 ;
        RECT 1.150 4.620 1.320 4.790 ;
        RECT 2.090 4.730 2.260 4.900 ;
        RECT 25.310 4.730 25.480 4.900 ;
        RECT 26.250 4.620 26.420 4.790 ;
        RECT 26.980 4.590 27.150 4.760 ;
        RECT 2.090 4.180 2.260 4.350 ;
        RECT 25.310 4.180 25.480 4.350 ;
      LAYER met1 ;
        RECT 0.360 10.090 0.520 10.790 ;
        RECT 0.360 9.540 0.630 10.090 ;
        RECT 0.350 9.490 0.630 9.540 ;
        RECT 0.770 9.750 0.960 10.740 ;
        RECT 1.170 10.060 1.330 10.790 ;
        RECT 2.120 10.520 2.360 10.540 ;
        RECT 2.010 10.200 2.360 10.520 ;
        RECT 1.130 10.040 1.330 10.060 ;
        RECT 1.120 9.800 1.350 10.040 ;
        RECT 2.120 9.970 2.360 10.200 ;
        RECT 2.010 9.900 2.360 9.970 ;
        RECT 1.120 9.750 1.330 9.800 ;
        RECT 0.770 9.630 0.940 9.750 ;
        RECT 0.350 9.400 0.520 9.490 ;
        RECT 0.360 8.890 0.520 9.400 ;
        RECT 0.770 8.890 0.930 9.630 ;
        RECT 1.170 8.890 1.330 9.750 ;
        RECT 2.010 9.650 2.350 9.900 ;
        RECT 2.120 9.640 2.350 9.650 ;
        RECT 2.110 9.420 2.350 9.640 ;
        RECT 10.360 9.340 10.590 10.630 ;
        RECT 0.360 8.220 0.520 8.730 ;
        RECT 0.350 8.130 0.520 8.220 ;
        RECT 0.350 8.080 0.630 8.130 ;
        RECT 0.360 7.530 0.630 8.080 ;
        RECT 0.770 7.990 0.930 8.730 ;
        RECT 0.770 7.870 0.940 7.990 ;
        RECT 1.170 7.870 1.330 8.730 ;
        RECT 2.120 8.430 2.360 9.070 ;
        RECT 2.120 8.170 2.350 8.430 ;
        RECT 2.110 7.970 2.350 8.170 ;
        RECT 0.360 7.080 0.520 7.530 ;
        RECT 0.360 6.530 0.630 7.080 ;
        RECT 0.350 6.480 0.630 6.530 ;
        RECT 0.770 6.740 0.960 7.870 ;
        RECT 1.120 7.820 1.330 7.870 ;
        RECT 2.010 7.950 2.350 7.970 ;
        RECT 1.120 7.580 1.350 7.820 ;
        RECT 2.010 7.650 2.330 7.950 ;
        RECT 10.360 7.820 10.590 9.110 ;
        RECT 1.130 7.560 1.330 7.580 ;
        RECT 1.170 7.050 1.330 7.560 ;
        RECT 2.120 7.510 2.360 7.600 ;
        RECT 2.010 7.100 2.360 7.510 ;
        RECT 3.660 7.420 3.790 7.440 ;
        RECT 3.630 7.190 3.870 7.420 ;
        RECT 3.660 7.150 3.770 7.190 ;
        RECT 1.130 7.030 1.330 7.050 ;
        RECT 1.120 6.790 1.350 7.030 ;
        RECT 2.120 6.960 2.360 7.100 ;
        RECT 1.120 6.740 1.330 6.790 ;
        RECT 0.770 6.620 0.940 6.740 ;
        RECT 0.350 6.390 0.520 6.480 ;
        RECT 0.360 5.880 0.520 6.390 ;
        RECT 0.770 5.880 0.930 6.620 ;
        RECT 1.170 5.880 1.330 6.740 ;
        RECT 2.010 6.640 2.350 6.960 ;
        RECT 2.110 6.480 2.350 6.640 ;
        RECT 10.360 6.370 10.590 7.660 ;
        RECT 0.360 5.220 0.520 5.730 ;
        RECT 0.350 5.130 0.520 5.220 ;
        RECT 0.350 5.080 0.630 5.130 ;
        RECT 0.360 4.530 0.630 5.080 ;
        RECT 0.770 4.990 0.930 5.730 ;
        RECT 0.770 4.870 0.940 4.990 ;
        RECT 1.170 4.870 1.330 5.730 ;
        RECT 2.120 5.490 2.360 6.130 ;
        RECT 2.120 5.230 2.350 5.490 ;
        RECT 2.110 5.010 2.350 5.230 ;
        RECT 0.360 3.830 0.520 4.530 ;
        RECT 0.770 3.880 0.960 4.870 ;
        RECT 1.120 4.820 1.330 4.870 ;
        RECT 1.120 4.580 1.350 4.820 ;
        RECT 2.010 4.650 2.330 4.970 ;
        RECT 10.360 4.830 10.590 6.120 ;
        RECT 1.130 4.560 1.330 4.580 ;
        RECT 1.170 3.830 1.330 4.560 ;
        RECT 2.010 4.100 2.330 4.420 ;
        RECT 10.960 4.280 11.230 10.330 ;
        RECT 16.340 4.280 16.610 10.330 ;
        RECT 16.980 9.340 17.210 10.630 ;
        RECT 25.210 10.520 25.450 10.540 ;
        RECT 25.210 10.200 25.560 10.520 ;
        RECT 25.210 9.970 25.450 10.200 ;
        RECT 26.240 10.060 26.400 10.790 ;
        RECT 26.240 10.040 26.440 10.060 ;
        RECT 25.210 9.900 25.560 9.970 ;
        RECT 25.220 9.650 25.560 9.900 ;
        RECT 26.220 9.800 26.450 10.040 ;
        RECT 26.240 9.750 26.450 9.800 ;
        RECT 26.610 9.750 26.800 10.740 ;
        RECT 27.050 10.090 27.210 10.790 ;
        RECT 25.220 9.640 25.450 9.650 ;
        RECT 25.220 9.420 25.460 9.640 ;
        RECT 16.980 7.820 17.210 9.110 ;
        RECT 25.210 8.430 25.450 9.070 ;
        RECT 26.240 8.890 26.400 9.750 ;
        RECT 26.630 9.630 26.800 9.750 ;
        RECT 26.640 8.890 26.800 9.630 ;
        RECT 26.940 9.540 27.210 10.090 ;
        RECT 26.940 9.490 27.220 9.540 ;
        RECT 27.050 9.400 27.220 9.490 ;
        RECT 27.050 8.890 27.210 9.400 ;
        RECT 25.220 8.170 25.450 8.430 ;
        RECT 25.220 7.970 25.460 8.170 ;
        RECT 25.220 7.950 25.560 7.970 ;
        RECT 16.980 6.370 17.210 7.660 ;
        RECT 25.240 7.650 25.560 7.950 ;
        RECT 26.240 7.870 26.400 8.730 ;
        RECT 26.640 7.990 26.800 8.730 ;
        RECT 27.050 8.220 27.210 8.730 ;
        RECT 27.050 8.130 27.220 8.220 ;
        RECT 26.630 7.870 26.800 7.990 ;
        RECT 26.240 7.820 26.450 7.870 ;
        RECT 25.210 7.510 25.450 7.600 ;
        RECT 26.220 7.580 26.450 7.820 ;
        RECT 26.240 7.560 26.440 7.580 ;
        RECT 23.780 7.420 23.910 7.440 ;
        RECT 23.700 7.190 23.940 7.420 ;
        RECT 23.800 7.150 23.910 7.190 ;
        RECT 25.210 7.100 25.560 7.510 ;
        RECT 25.210 6.960 25.450 7.100 ;
        RECT 26.240 7.050 26.400 7.560 ;
        RECT 26.240 7.030 26.440 7.050 ;
        RECT 25.220 6.640 25.560 6.960 ;
        RECT 26.220 6.790 26.450 7.030 ;
        RECT 26.240 6.740 26.450 6.790 ;
        RECT 26.610 6.740 26.800 7.870 ;
        RECT 26.940 8.080 27.220 8.130 ;
        RECT 26.940 7.530 27.210 8.080 ;
        RECT 27.050 7.080 27.210 7.530 ;
        RECT 25.220 6.480 25.460 6.640 ;
        RECT 16.980 4.830 17.210 6.120 ;
        RECT 25.210 5.490 25.450 6.130 ;
        RECT 26.240 5.880 26.400 6.740 ;
        RECT 26.630 6.620 26.800 6.740 ;
        RECT 26.640 5.880 26.800 6.620 ;
        RECT 26.940 6.530 27.210 7.080 ;
        RECT 26.940 6.480 27.220 6.530 ;
        RECT 27.050 6.390 27.220 6.480 ;
        RECT 27.050 5.880 27.210 6.390 ;
        RECT 25.220 5.230 25.450 5.490 ;
        RECT 25.220 5.010 25.460 5.230 ;
        RECT 25.240 4.650 25.560 4.970 ;
        RECT 26.240 4.870 26.400 5.730 ;
        RECT 26.640 4.990 26.800 5.730 ;
        RECT 27.050 5.220 27.210 5.730 ;
        RECT 27.050 5.130 27.220 5.220 ;
        RECT 26.630 4.870 26.800 4.990 ;
        RECT 26.240 4.820 26.450 4.870 ;
        RECT 26.220 4.580 26.450 4.820 ;
        RECT 26.240 4.560 26.440 4.580 ;
        RECT 25.240 4.100 25.560 4.420 ;
        RECT 26.240 3.830 26.400 4.560 ;
        RECT 26.610 3.880 26.800 4.870 ;
        RECT 26.940 5.080 27.220 5.130 ;
        RECT 26.940 4.530 27.210 5.080 ;
        RECT 27.050 3.830 27.210 4.530 ;
      LAYER via ;
        RECT 2.040 10.230 2.300 10.490 ;
        RECT 2.040 9.680 2.300 9.940 ;
        RECT 2.040 7.680 2.300 7.940 ;
        RECT 2.040 7.130 2.300 7.480 ;
        RECT 2.040 6.670 2.300 6.930 ;
        RECT 2.040 4.680 2.300 4.940 ;
        RECT 2.040 4.130 2.300 4.390 ;
        RECT 25.270 10.230 25.530 10.490 ;
        RECT 25.270 9.680 25.530 9.940 ;
        RECT 25.270 7.680 25.530 7.940 ;
        RECT 25.270 7.130 25.530 7.480 ;
        RECT 25.270 6.670 25.530 6.930 ;
        RECT 25.270 4.680 25.530 4.940 ;
        RECT 25.270 4.130 25.530 4.390 ;
      LAYER met2 ;
        RECT 2.020 10.240 2.330 10.530 ;
        RECT 0.000 10.200 2.330 10.240 ;
        RECT 25.240 10.240 25.550 10.530 ;
        RECT 25.240 10.200 27.570 10.240 ;
        RECT 0.000 10.060 2.180 10.200 ;
        RECT 25.390 10.060 27.570 10.200 ;
        RECT 2.020 9.810 2.330 9.980 ;
        RECT 0.000 9.650 2.330 9.810 ;
        RECT 0.000 9.630 2.170 9.650 ;
        RECT 2.470 9.630 2.560 9.810 ;
        RECT 5.360 9.760 12.240 9.830 ;
        RECT 5.330 9.650 12.240 9.760 ;
        RECT 15.330 9.760 22.210 9.830 ;
        RECT 25.240 9.810 25.550 9.980 ;
        RECT 15.330 9.650 22.240 9.760 ;
        RECT 25.010 9.630 25.100 9.810 ;
        RECT 25.240 9.650 27.570 9.810 ;
        RECT 25.400 9.630 27.570 9.650 ;
        RECT 3.230 9.220 12.240 9.400 ;
        RECT 15.330 9.220 24.340 9.400 ;
        RECT 5.360 8.340 12.240 8.400 ;
        RECT 5.330 8.220 12.240 8.340 ;
        RECT 15.330 8.340 22.210 8.400 ;
        RECT 15.330 8.220 22.240 8.340 ;
        RECT 0.000 7.970 2.170 7.990 ;
        RECT 0.000 7.810 2.330 7.970 ;
        RECT 2.470 7.810 2.560 7.990 ;
        RECT 5.370 7.900 12.240 7.970 ;
        RECT 2.020 7.640 2.330 7.810 ;
        RECT 5.330 7.790 12.240 7.900 ;
        RECT 15.330 7.900 22.200 7.970 ;
        RECT 15.330 7.790 22.240 7.900 ;
        RECT 25.010 7.810 25.100 7.990 ;
        RECT 25.400 7.970 27.570 7.990 ;
        RECT 25.240 7.810 27.570 7.970 ;
        RECT 25.240 7.640 25.550 7.810 ;
        RECT 0.000 7.520 2.180 7.560 ;
        RECT 25.390 7.520 27.570 7.560 ;
        RECT 0.000 7.380 2.330 7.520 ;
        RECT 2.020 7.230 2.330 7.380 ;
        RECT 0.000 7.090 2.330 7.230 ;
        RECT 25.240 7.380 27.570 7.520 ;
        RECT 25.240 7.230 25.550 7.380 ;
        RECT 25.240 7.090 27.570 7.230 ;
        RECT 0.000 7.050 2.180 7.090 ;
        RECT 25.390 7.050 27.570 7.090 ;
        RECT 2.020 6.800 2.330 6.970 ;
        RECT 0.000 6.640 2.330 6.800 ;
        RECT 0.000 6.620 2.170 6.640 ;
        RECT 2.470 6.620 2.560 6.800 ;
        RECT 5.330 6.640 12.240 6.810 ;
        RECT 15.330 6.640 22.240 6.810 ;
        RECT 25.240 6.800 25.550 6.970 ;
        RECT 25.010 6.620 25.100 6.800 ;
        RECT 25.240 6.640 27.570 6.800 ;
        RECT 25.400 6.620 27.570 6.640 ;
        RECT 5.330 6.220 12.240 6.390 ;
        RECT 15.330 6.220 22.240 6.390 ;
        RECT 5.330 5.240 12.240 5.410 ;
        RECT 15.330 5.240 22.240 5.410 ;
        RECT 0.000 4.970 2.170 4.990 ;
        RECT 0.000 4.810 2.330 4.970 ;
        RECT 2.470 4.810 2.560 4.990 ;
        RECT 2.020 4.640 2.330 4.810 ;
        RECT 5.330 4.800 12.240 4.970 ;
        RECT 15.330 4.800 22.240 4.970 ;
        RECT 25.010 4.810 25.100 4.990 ;
        RECT 25.400 4.970 27.570 4.990 ;
        RECT 25.240 4.810 27.570 4.970 ;
        RECT 25.240 4.640 25.550 4.810 ;
        RECT 0.000 4.420 2.180 4.560 ;
        RECT 25.390 4.420 27.570 4.560 ;
        RECT 0.000 4.380 2.330 4.420 ;
        RECT 2.020 4.090 2.330 4.380 ;
        RECT 25.240 4.380 27.570 4.420 ;
        RECT 25.240 4.090 25.550 4.380 ;
        RECT 7.200 3.610 7.320 3.690 ;
        RECT 20.290 3.550 20.410 3.690 ;
  END
END sky130_hilas_swc4x2cellOverlap

MACRO sky130_hilas_FGBias2x1cell
  CLASS CORE ;
  FOREIGN sky130_hilas_FGBias2x1cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.540 BY 10.520 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VTUN
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 0.350 0.470 0.770 6.520 ;
    END
  END VTUN
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2.830 3.660 3.060 6.520 ;
        RECT 2.830 3.370 3.160 3.660 ;
        RECT 2.830 0.470 3.060 3.370 ;
    END
  END VGND
  PIN GATE_CONTROL
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 4.050 0.470 4.280 6.520 ;
    END
  END GATE_CONTROL
  PIN DRAIN1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 5.840 9.120 6.020 ;
    END
  END DRAIN1
  PIN DRAIN4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 9.060 1.140 9.220 1.160 ;
        RECT 0.000 1.090 9.220 1.140 ;
        RECT 0.000 0.990 9.100 1.090 ;
    END
  END DRAIN4
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 11.170 3.660 11.490 3.740 ;
        RECT 10.180 3.480 11.490 3.660 ;
        RECT 10.180 3.310 11.360 3.480 ;
        RECT 10.230 3.160 10.550 3.310 ;
    END
  END VINJ
  PIN OUTPUT1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 9.340 5.000 9.650 5.220 ;
        RECT 9.340 4.890 11.530 5.000 ;
        RECT 9.500 4.780 11.530 4.890 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 9.340 2.240 9.650 2.460 ;
        RECT 9.340 2.130 11.530 2.240 ;
        RECT 9.490 2.030 11.530 2.130 ;
    END
  END OUTPUT2
  PIN GATECOL
    PORT
      LAYER met1 ;
        RECT 10.570 6.480 10.760 6.520 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.570 0.470 10.760 0.520 ;
    END
  END GATECOL
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 11.010 3.770 11.290 6.520 ;
        RECT 11.010 3.450 11.460 3.770 ;
        RECT 11.010 0.470 11.290 3.450 ;
      LAYER via ;
        RECT 11.200 3.480 11.460 3.740 ;
    END
  END VINJ
  OBS
      LAYER nwell ;
        RECT 14.520 10.180 16.250 10.520 ;
        RECT 14.500 8.620 16.250 10.180 ;
        RECT 14.500 6.990 16.230 8.620 ;
        RECT 12.980 6.600 16.290 6.990 ;
        RECT 12.980 6.560 16.530 6.600 ;
        RECT 8.220 6.510 11.530 6.520 ;
        RECT 10.570 6.480 10.760 6.510 ;
        RECT 12.980 4.910 16.540 6.560 ;
        RECT 0.590 1.870 1.150 4.290 ;
        RECT 12.980 3.820 16.290 4.910 ;
        RECT 12.980 1.980 16.290 3.170 ;
        RECT 12.980 0.330 16.540 1.980 ;
        RECT 12.980 0.290 16.530 0.330 ;
        RECT 12.980 0.000 16.290 0.290 ;
      LAYER li1 ;
        RECT 14.920 8.790 15.470 9.220 ;
        RECT 14.920 7.060 15.470 7.490 ;
        RECT 13.880 6.360 14.410 6.530 ;
        RECT 15.690 6.260 15.890 6.610 ;
        RECT 15.690 6.230 15.900 6.260 ;
        RECT 14.120 5.430 14.350 6.120 ;
        RECT 9.350 5.140 9.670 5.180 ;
        RECT 9.350 4.950 9.680 5.140 ;
        RECT 9.350 4.920 9.670 4.950 ;
        RECT 14.130 4.280 14.300 5.430 ;
        RECT 14.960 4.370 15.130 5.980 ;
        RECT 15.680 5.650 15.900 6.230 ;
        RECT 15.690 5.640 15.900 5.650 ;
        RECT 15.330 5.470 15.520 5.480 ;
        RECT 15.330 5.180 15.530 5.470 ;
        RECT 15.320 4.850 15.610 5.180 ;
        RECT 14.960 4.180 15.140 4.370 ;
        RECT 3.040 3.630 3.230 3.950 ;
        RECT 2.950 3.540 3.230 3.630 ;
        RECT 2.950 3.400 6.590 3.540 ;
        RECT 3.040 3.360 6.590 3.400 ;
        RECT 3.040 2.940 3.230 3.360 ;
        RECT 9.350 2.380 9.670 2.420 ;
        RECT 4.070 2.320 4.300 2.360 ;
        RECT 9.350 2.190 9.680 2.380 ;
        RECT 9.350 2.160 9.670 2.190 ;
        RECT 14.130 1.460 14.300 2.710 ;
        RECT 14.960 2.620 15.140 2.810 ;
        RECT 14.120 0.770 14.350 1.460 ;
        RECT 14.960 1.010 15.130 2.620 ;
        RECT 15.320 1.810 15.610 2.140 ;
        RECT 15.330 1.520 15.530 1.810 ;
        RECT 15.330 1.510 15.520 1.520 ;
        RECT 15.690 1.340 15.900 1.350 ;
        RECT 15.680 0.760 15.900 1.340 ;
        RECT 15.690 0.730 15.900 0.760 ;
        RECT 13.880 0.460 14.410 0.630 ;
        RECT 15.690 0.380 15.890 0.730 ;
      LAYER mcon ;
        RECT 14.920 8.870 15.190 9.140 ;
        RECT 14.920 7.140 15.190 7.410 ;
        RECT 14.150 5.910 14.320 6.080 ;
        RECT 15.700 6.060 15.870 6.230 ;
        RECT 14.150 5.460 14.320 5.630 ;
        RECT 9.410 4.960 9.580 5.130 ;
        RECT 15.340 5.220 15.520 5.410 ;
        RECT 2.960 3.430 3.130 3.600 ;
        RECT 9.410 2.200 9.580 2.370 ;
        RECT 14.150 1.260 14.320 1.430 ;
        RECT 15.340 1.580 15.520 1.770 ;
        RECT 14.150 0.810 14.320 0.980 ;
        RECT 15.700 0.760 15.870 0.930 ;
      LAYER met1 ;
        RECT 14.860 6.600 15.250 10.190 ;
        RECT 13.810 6.170 14.120 6.560 ;
        RECT 13.810 6.120 14.360 6.170 ;
        RECT 14.100 5.380 14.360 6.120 ;
        RECT 15.330 5.480 15.520 6.930 ;
        RECT 15.770 6.290 15.930 6.930 ;
        RECT 15.660 5.740 15.930 6.290 ;
        RECT 15.660 5.690 15.940 5.740 ;
        RECT 15.770 5.600 15.940 5.690 ;
        RECT 15.330 5.450 15.550 5.480 ;
        RECT 9.340 4.890 9.660 5.210 ;
        RECT 15.310 5.180 15.560 5.450 ;
        RECT 15.320 5.170 15.560 5.180 ;
        RECT 15.320 4.930 15.550 5.170 ;
        RECT 14.930 4.120 15.170 4.500 ;
        RECT 10.260 3.730 10.520 4.050 ;
        RECT 15.360 3.910 15.520 4.930 ;
        RECT 15.770 3.910 15.930 5.600 ;
        RECT 10.260 3.130 10.520 3.450 ;
        RECT 14.930 2.490 15.170 2.870 ;
        RECT 9.340 2.130 9.660 2.450 ;
        RECT 15.360 2.060 15.520 3.080 ;
        RECT 15.320 1.820 15.550 2.060 ;
        RECT 15.320 1.810 15.560 1.820 ;
        RECT 15.310 1.540 15.560 1.810 ;
        RECT 15.330 1.510 15.550 1.540 ;
        RECT 14.100 0.870 14.360 1.510 ;
        RECT 13.810 0.720 14.360 0.870 ;
        RECT 13.810 0.430 14.120 0.720 ;
        RECT 15.330 0.060 15.520 1.510 ;
        RECT 15.770 1.390 15.930 3.080 ;
        RECT 15.770 1.300 15.940 1.390 ;
        RECT 15.660 1.250 15.940 1.300 ;
        RECT 15.660 0.700 15.930 1.250 ;
        RECT 15.770 0.060 15.930 0.700 ;
      LAYER via ;
        RECT 13.840 6.150 14.100 6.410 ;
        RECT 9.370 4.920 9.630 5.180 ;
        RECT 10.260 3.760 10.520 4.020 ;
        RECT 10.260 3.160 10.520 3.420 ;
        RECT 9.370 2.160 9.630 2.420 ;
        RECT 13.840 0.580 14.100 0.840 ;
      LAYER met2 ;
        RECT 13.810 6.440 14.120 6.450 ;
        RECT 13.810 6.260 16.290 6.440 ;
        RECT 13.810 6.120 14.120 6.260 ;
        RECT 10.230 3.760 10.550 4.020 ;
        RECT 13.810 0.730 14.120 0.870 ;
        RECT 13.810 0.550 16.290 0.730 ;
        RECT 13.810 0.540 14.120 0.550 ;
  END
END sky130_hilas_FGBias2x1cell

MACRO sky130_hilas_drainSelect01
  CLASS CORE ;
  FOREIGN sky130_hilas_drainSelect01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.000 BY 6.110 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DRAIN3
    PORT
      LAYER met2 ;
        RECT 0.000 2.590 0.570 2.600 ;
        RECT 0.000 2.580 1.270 2.590 ;
        RECT 0.000 2.420 2.000 2.580 ;
    END
  END DRAIN3
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.580 6.040 0.830 6.110 ;
    END
  END VINJ
  PIN DRAIN_MUX
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 3.570 6.040 3.800 6.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.570 0.060 3.800 0.140 ;
    END
  END DRAIN_MUX
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 4.920 0.060 5.110 0.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.920 6.060 5.110 6.110 ;
    END
  END VGND
  PIN SELECT2
    ANTENNADIFFAREA 0.322600 ;
    PORT
      LAYER met2 ;
        RECT 4.070 4.000 4.390 4.050 ;
        RECT 5.570 4.000 5.720 4.080 ;
        RECT 6.480 4.000 6.800 4.080 ;
        RECT 4.070 3.810 6.800 4.000 ;
        RECT 4.070 3.790 4.390 3.810 ;
        RECT 6.480 3.760 6.800 3.810 ;
    END
  END SELECT2
  PIN SELECT1
    ANTENNADIFFAREA 0.322600 ;
    PORT
      LAYER met2 ;
        RECT 4.070 5.440 4.390 5.460 ;
        RECT 6.480 5.440 6.800 5.490 ;
        RECT 4.070 5.250 6.800 5.440 ;
        RECT 4.070 5.200 4.390 5.250 ;
        RECT 5.640 5.180 5.720 5.250 ;
        RECT 6.480 5.170 6.800 5.250 ;
    END
  END SELECT1
  PIN SELECT3
    ANTENNADIFFAREA 0.322600 ;
    PORT
      LAYER met2 ;
        RECT 4.070 2.240 4.390 2.260 ;
        RECT 6.480 2.240 6.800 2.290 ;
        RECT 4.070 2.050 6.800 2.240 ;
        RECT 4.070 2.000 4.390 2.050 ;
        RECT 5.640 1.980 5.720 2.050 ;
        RECT 6.480 1.970 6.800 2.050 ;
    END
  END SELECT3
  PIN SELECT4
    ANTENNADIFFAREA 0.322600 ;
    PORT
      LAYER met2 ;
        RECT 4.070 0.800 4.390 0.850 ;
        RECT 5.630 0.800 5.720 0.870 ;
        RECT 6.480 0.800 6.800 0.880 ;
        RECT 4.070 0.610 6.800 0.800 ;
        RECT 4.070 0.590 4.390 0.610 ;
        RECT 6.480 0.560 6.800 0.610 ;
    END
  END SELECT4
  OBS
      LAYER nwell ;
        RECT 2.320 4.630 5.740 5.870 ;
        RECT 0.000 4.620 5.740 4.630 ;
        RECT 2.320 3.380 5.740 4.620 ;
        RECT 2.320 1.430 5.740 2.670 ;
        RECT 0.000 1.410 5.740 1.430 ;
        RECT 2.320 0.180 5.740 1.410 ;
      LAYER li1 ;
        RECT 2.540 4.650 2.710 5.540 ;
        RECT 2.540 3.710 2.710 4.600 ;
        RECT 2.940 3.760 3.110 5.490 ;
        RECT 6.630 5.420 6.870 5.450 ;
        RECT 3.640 5.250 4.600 5.420 ;
        RECT 5.050 5.250 6.390 5.420 ;
        RECT 6.630 5.250 7.200 5.420 ;
        RECT 3.920 5.240 4.090 5.250 ;
        RECT 6.630 5.210 6.870 5.250 ;
        RECT 7.510 5.120 7.680 5.540 ;
        RECT 4.120 4.800 4.460 4.980 ;
        RECT 7.580 4.900 7.750 4.940 ;
        RECT 3.640 4.630 6.390 4.800 ;
        RECT 6.850 4.630 7.220 4.800 ;
        RECT 3.640 4.450 6.390 4.620 ;
        RECT 6.850 4.450 7.220 4.620 ;
        RECT 7.320 4.510 7.510 4.740 ;
        RECT 7.580 4.730 7.810 4.900 ;
        RECT 7.580 4.520 7.750 4.730 ;
        RECT 4.120 4.270 4.460 4.450 ;
        RECT 7.580 4.350 7.810 4.520 ;
        RECT 7.580 4.310 7.750 4.350 ;
        RECT 3.920 4.000 4.090 4.010 ;
        RECT 6.630 4.000 6.870 4.040 ;
        RECT 3.640 3.830 4.600 4.000 ;
        RECT 5.050 3.830 6.390 4.000 ;
        RECT 6.630 3.830 7.200 4.000 ;
        RECT 6.630 3.800 6.870 3.830 ;
        RECT 7.510 3.710 7.680 4.130 ;
        RECT 2.540 1.450 2.710 2.340 ;
        RECT 2.540 0.510 2.710 1.400 ;
        RECT 2.940 0.560 3.110 2.290 ;
        RECT 6.630 2.220 6.870 2.250 ;
        RECT 3.640 2.050 4.600 2.220 ;
        RECT 5.050 2.050 6.390 2.220 ;
        RECT 6.630 2.050 7.200 2.220 ;
        RECT 3.920 2.040 4.090 2.050 ;
        RECT 6.630 2.010 6.870 2.050 ;
        RECT 7.510 1.920 7.680 2.340 ;
        RECT 4.120 1.600 4.460 1.780 ;
        RECT 7.580 1.700 7.750 1.740 ;
        RECT 3.640 1.430 6.390 1.600 ;
        RECT 6.850 1.430 7.220 1.600 ;
        RECT 3.640 1.250 6.390 1.420 ;
        RECT 6.850 1.250 7.220 1.420 ;
        RECT 7.320 1.310 7.510 1.540 ;
        RECT 7.580 1.530 7.810 1.700 ;
        RECT 7.580 1.320 7.750 1.530 ;
        RECT 4.120 1.070 4.460 1.250 ;
        RECT 7.580 1.150 7.810 1.320 ;
        RECT 7.580 1.110 7.750 1.150 ;
        RECT 3.920 0.800 4.090 0.810 ;
        RECT 6.630 0.800 6.870 0.840 ;
        RECT 3.640 0.630 4.600 0.800 ;
        RECT 5.050 0.630 6.390 0.800 ;
        RECT 6.630 0.630 7.200 0.800 ;
        RECT 6.630 0.600 6.870 0.630 ;
        RECT 7.510 0.510 7.680 0.930 ;
      LAYER mcon ;
        RECT 2.540 5.370 2.710 5.540 ;
        RECT 2.540 5.010 2.710 5.180 ;
        RECT 5.920 5.250 6.090 5.420 ;
        RECT 6.670 5.250 6.840 5.420 ;
        RECT 7.510 5.370 7.680 5.540 ;
        RECT 2.940 4.920 3.110 5.090 ;
        RECT 2.540 4.430 2.710 4.600 ;
        RECT 2.540 4.070 2.710 4.240 ;
        RECT 7.330 4.540 7.500 4.710 ;
        RECT 7.640 4.730 7.810 4.900 ;
        RECT 2.940 4.160 3.110 4.330 ;
        RECT 7.640 4.350 7.810 4.520 ;
        RECT 3.920 3.840 4.090 4.010 ;
        RECT 5.920 3.830 6.090 4.000 ;
        RECT 6.670 3.830 6.840 4.000 ;
        RECT 2.540 2.170 2.710 2.340 ;
        RECT 2.540 1.810 2.710 1.980 ;
        RECT 5.920 2.050 6.090 2.220 ;
        RECT 6.670 2.050 6.840 2.220 ;
        RECT 7.510 2.170 7.680 2.340 ;
        RECT 2.940 1.720 3.110 1.890 ;
        RECT 2.540 1.230 2.710 1.400 ;
        RECT 2.540 0.870 2.710 1.040 ;
        RECT 7.330 1.340 7.500 1.510 ;
        RECT 7.640 1.530 7.810 1.700 ;
        RECT 2.940 0.960 3.110 1.130 ;
        RECT 7.640 1.150 7.810 1.320 ;
        RECT 3.920 0.640 4.090 0.810 ;
        RECT 5.920 0.630 6.090 0.800 ;
        RECT 6.670 0.630 6.840 0.800 ;
      LAYER met1 ;
        RECT 2.900 5.600 3.150 5.820 ;
        RECT 0.580 4.620 0.830 4.630 ;
        RECT 2.510 3.650 3.150 5.600 ;
        RECT 4.050 5.440 4.390 5.490 ;
        RECT 3.830 5.420 4.390 5.440 ;
        RECT 3.830 5.250 4.510 5.420 ;
        RECT 3.830 5.210 4.390 5.250 ;
        RECT 4.050 5.170 4.390 5.210 ;
        RECT 4.050 4.040 4.390 4.080 ;
        RECT 3.830 4.000 4.390 4.040 ;
        RECT 3.830 3.830 4.510 4.000 ;
        RECT 3.830 3.810 4.390 3.830 ;
        RECT 4.050 3.760 4.390 3.810 ;
        RECT 2.900 3.430 3.150 3.650 ;
        RECT 5.890 3.430 6.120 5.820 ;
        RECT 7.240 5.600 7.430 5.820 ;
        RECT 6.480 5.460 6.850 5.480 ;
        RECT 6.480 5.200 6.900 5.460 ;
        RECT 6.480 5.190 6.850 5.200 ;
        RECT 7.240 5.110 7.710 5.600 ;
        RECT 7.240 4.770 7.430 5.110 ;
        RECT 7.240 4.480 7.530 4.770 ;
        RECT 7.570 4.670 7.890 4.950 ;
        RECT 7.240 4.140 7.430 4.480 ;
        RECT 7.570 4.300 7.890 4.580 ;
        RECT 6.480 4.050 6.850 4.060 ;
        RECT 6.480 3.790 6.900 4.050 ;
        RECT 6.480 3.770 6.850 3.790 ;
        RECT 7.240 3.650 7.710 4.140 ;
        RECT 7.240 3.430 7.430 3.650 ;
        RECT 2.900 2.400 3.150 2.620 ;
        RECT 0.580 1.420 0.830 1.430 ;
        RECT 2.510 0.450 3.150 2.400 ;
        RECT 4.050 2.240 4.390 2.290 ;
        RECT 3.830 2.220 4.390 2.240 ;
        RECT 3.830 2.050 4.510 2.220 ;
        RECT 3.830 2.010 4.390 2.050 ;
        RECT 4.050 1.970 4.390 2.010 ;
        RECT 4.050 0.840 4.390 0.880 ;
        RECT 3.830 0.800 4.390 0.840 ;
        RECT 3.830 0.630 4.510 0.800 ;
        RECT 3.830 0.610 4.390 0.630 ;
        RECT 4.050 0.560 4.390 0.610 ;
        RECT 2.900 0.230 3.150 0.450 ;
        RECT 5.890 0.230 6.120 2.620 ;
        RECT 7.240 2.400 7.430 2.620 ;
        RECT 6.480 2.260 6.850 2.280 ;
        RECT 6.480 2.000 6.900 2.260 ;
        RECT 6.480 1.990 6.850 2.000 ;
        RECT 7.240 1.910 7.710 2.400 ;
        RECT 7.240 1.570 7.430 1.910 ;
        RECT 7.240 1.280 7.530 1.570 ;
        RECT 7.570 1.470 7.890 1.750 ;
        RECT 7.240 0.940 7.430 1.280 ;
        RECT 7.570 1.100 7.890 1.380 ;
        RECT 6.480 0.850 6.850 0.860 ;
        RECT 6.480 0.590 6.900 0.850 ;
        RECT 6.480 0.570 6.850 0.590 ;
        RECT 7.240 0.450 7.710 0.940 ;
        RECT 7.240 0.230 7.430 0.450 ;
      LAYER via ;
        RECT 4.100 5.200 4.360 5.460 ;
        RECT 4.100 3.790 4.360 4.050 ;
        RECT 6.510 5.200 6.770 5.460 ;
        RECT 7.600 4.680 7.860 4.940 ;
        RECT 7.600 4.310 7.860 4.570 ;
        RECT 6.510 3.790 6.770 4.050 ;
        RECT 4.100 2.000 4.360 2.260 ;
        RECT 4.100 0.590 4.360 0.850 ;
        RECT 6.510 2.000 6.770 2.260 ;
        RECT 7.600 1.480 7.860 1.740 ;
        RECT 7.600 1.110 7.860 1.370 ;
        RECT 6.510 0.590 6.770 0.850 ;
      LAYER met2 ;
        RECT 0.000 5.680 1.780 5.860 ;
        RECT 7.560 4.730 8.000 4.960 ;
        RECT 7.560 4.660 7.900 4.730 ;
        RECT 7.560 4.520 7.900 4.590 ;
        RECT 7.560 4.290 8.000 4.520 ;
        RECT 0.000 3.380 1.780 3.540 ;
        RECT 7.560 1.530 8.000 1.760 ;
        RECT 7.560 1.460 7.900 1.530 ;
        RECT 7.560 1.320 7.900 1.390 ;
        RECT 7.560 1.090 8.000 1.320 ;
        RECT 0.000 0.160 1.780 0.330 ;
  END
END sky130_hilas_drainSelect01

MACRO sky130_hilas_DAC5bit01
  CLASS CORE ;
  FOREIGN sky130_hilas_DAC5bit01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.580 BY 7.990 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 8.350 0.980 8.670 1.110 ;
        RECT 0.000 0.850 8.670 0.980 ;
        RECT 0.000 0.780 8.540 0.850 ;
    END
  END A0
  PIN A1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 11.710 2.100 11.860 5.840 ;
        RECT 0.000 1.900 11.870 2.100 ;
        RECT 0.000 1.890 0.140 1.900 ;
    END
  END A1
  PIN A2
    USE ANALOG ;
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER met2 ;
        RECT 10.110 3.080 10.310 5.680 ;
        RECT 0.000 2.870 10.310 3.080 ;
        RECT 0.320 2.670 0.640 2.870 ;
    END
  END A2
  PIN A3
    USE ANALOG ;
    ANTENNAGATEAREA 0.307500 ;
    PORT
      LAYER met2 ;
        RECT 0.000 4.950 2.060 5.010 ;
        RECT 3.480 4.950 3.700 5.410 ;
        RECT 8.400 4.960 8.650 5.720 ;
        RECT 8.400 4.950 8.680 4.960 ;
        RECT 0.000 4.800 8.680 4.950 ;
        RECT 0.260 4.560 0.620 4.800 ;
        RECT 1.900 4.650 8.680 4.800 ;
    END
  END A3
  PIN A4
    USE ANALOG ;
    ANTENNAGATEAREA 6.324800 ;
    ANTENNADIFFAREA 0.522900 ;
    PORT
      LAYER met2 ;
        RECT 0.320 5.960 0.640 6.190 ;
        RECT 2.030 5.960 2.350 6.230 ;
        RECT 5.230 5.960 5.550 6.230 ;
        RECT 6.840 5.960 7.160 6.240 ;
        RECT 0.000 5.920 7.160 5.960 ;
        RECT 0.000 5.770 7.050 5.920 ;
        RECT 8.460 5.910 8.780 6.230 ;
        RECT 10.070 5.920 10.390 6.240 ;
        RECT 11.680 5.920 12.000 6.240 ;
        RECT 0.000 5.750 0.290 5.770 ;
        RECT 3.750 5.150 4.070 5.470 ;
    END
  END A4
  PIN VPWR
    USE ANALOG ;
    ANTENNADIFFAREA 2.316600 ;
    PORT
      LAYER met2 ;
        RECT 12.970 5.960 13.280 5.980 ;
        RECT 13.640 5.960 13.950 5.980 ;
        RECT 12.710 5.680 13.950 5.960 ;
        RECT 12.970 5.650 13.280 5.680 ;
        RECT 13.460 5.670 13.950 5.680 ;
        RECT 13.640 5.650 13.950 5.670 ;
    END
  END VPWR
  PIN OUT
    USE ANALOG ;
    ANTENNADIFFAREA 0.947700 ;
    PORT
      LAYER met1 ;
        RECT 3.110 0.230 3.340 0.360 ;
        RECT 4.730 0.230 4.960 0.360 ;
        RECT 6.330 0.230 6.560 0.360 ;
        RECT 7.950 0.230 8.180 0.360 ;
        RECT 9.550 0.230 9.780 0.360 ;
        RECT 11.170 0.230 11.400 0.360 ;
        RECT 12.770 0.230 13.000 0.360 ;
        RECT 14.380 0.230 14.610 0.360 ;
        RECT 3.040 0.000 16.580 0.230 ;
    END
  END OUT
  OBS
      LAYER nwell ;
        RECT 0.270 7.030 1.880 7.990 ;
        RECT 1.890 7.030 16.370 7.990 ;
        RECT 0.270 5.820 16.370 7.030 ;
        RECT 0.270 5.110 6.710 5.820 ;
        RECT 6.770 5.360 16.370 5.820 ;
        RECT 8.320 5.110 16.370 5.360 ;
        RECT 0.270 2.940 16.370 5.110 ;
        RECT 0.270 1.980 1.880 2.830 ;
        RECT 1.890 1.980 16.370 2.830 ;
      LAYER li1 ;
        RECT 2.260 6.440 2.430 6.770 ;
        RECT 2.940 6.440 3.110 6.770 ;
        RECT 3.870 6.440 4.040 6.770 ;
        RECT 4.550 6.440 4.720 6.770 ;
        RECT 5.480 6.440 5.650 6.770 ;
        RECT 6.160 6.440 6.330 6.770 ;
        RECT 6.770 6.290 6.980 6.720 ;
        RECT 7.090 6.440 7.260 6.770 ;
        RECT 7.770 6.440 7.940 6.770 ;
        RECT 8.700 6.440 8.870 6.770 ;
        RECT 9.380 6.440 9.550 6.770 ;
        RECT 10.310 6.440 10.480 6.770 ;
        RECT 10.990 6.440 11.160 6.770 ;
        RECT 11.920 6.440 12.090 6.770 ;
        RECT 12.600 6.440 12.770 6.770 ;
        RECT 13.530 6.440 13.700 6.770 ;
        RECT 14.210 6.440 14.380 6.770 ;
        RECT 6.790 6.270 6.960 6.290 ;
        RECT 0.370 5.720 0.580 6.150 ;
        RECT 2.080 5.810 2.290 6.190 ;
        RECT 5.280 5.810 5.490 6.190 ;
        RECT 2.080 5.760 2.430 5.810 ;
        RECT 2.100 5.740 2.430 5.760 ;
        RECT 0.390 5.700 0.560 5.720 ;
        RECT 2.260 5.480 2.430 5.740 ;
        RECT 2.940 5.480 3.110 5.810 ;
        RECT 3.870 5.480 4.040 5.810 ;
        RECT 4.550 5.480 4.720 5.810 ;
        RECT 5.280 5.760 5.650 5.810 ;
        RECT 5.300 5.740 5.470 5.760 ;
        RECT 5.480 5.480 5.650 5.760 ;
        RECT 6.160 5.480 6.330 5.810 ;
        RECT 6.890 5.770 7.100 6.200 ;
        RECT 7.150 5.980 7.320 6.310 ;
        RECT 7.830 5.980 8.000 6.310 ;
        RECT 8.510 5.810 8.720 6.190 ;
        RECT 10.120 5.810 10.330 6.200 ;
        RECT 11.730 5.810 11.940 6.200 ;
        RECT 12.980 5.900 13.300 5.940 ;
        RECT 13.650 5.900 13.970 5.940 ;
        RECT 6.910 5.750 7.080 5.770 ;
        RECT 8.510 5.760 8.870 5.810 ;
        RECT 8.530 5.740 8.870 5.760 ;
        RECT 8.700 5.480 8.870 5.740 ;
        RECT 9.380 5.480 9.550 5.810 ;
        RECT 10.120 5.770 10.480 5.810 ;
        RECT 10.140 5.750 10.480 5.770 ;
        RECT 10.310 5.480 10.480 5.750 ;
        RECT 10.990 5.480 11.160 5.810 ;
        RECT 11.730 5.770 12.090 5.810 ;
        RECT 11.750 5.750 12.090 5.770 ;
        RECT 11.920 5.480 12.090 5.750 ;
        RECT 12.600 5.480 12.770 5.810 ;
        RECT 12.980 5.800 13.310 5.900 ;
        RECT 13.650 5.810 13.980 5.900 ;
        RECT 12.950 5.710 13.310 5.800 ;
        RECT 13.530 5.710 13.980 5.810 ;
        RECT 12.950 5.680 13.300 5.710 ;
        RECT 13.530 5.680 13.970 5.710 ;
        RECT 3.600 5.400 4.030 5.420 ;
        RECT 3.580 5.230 4.030 5.400 ;
        RECT 8.370 5.290 8.540 5.310 ;
        RECT 3.600 5.210 4.030 5.230 ;
        RECT 3.980 5.020 4.150 5.030 ;
        RECT 8.350 5.020 8.560 5.290 ;
        RECT 12.950 5.020 13.160 5.680 ;
        RECT 13.530 5.480 13.790 5.680 ;
        RECT 14.210 5.480 14.380 5.810 ;
        RECT 13.620 5.020 13.790 5.480 ;
        RECT 2.370 4.850 13.800 5.020 ;
        RECT 0.350 4.410 0.560 4.840 ;
        RECT 2.260 4.790 13.800 4.850 ;
        RECT 2.260 4.520 2.540 4.790 ;
        RECT 2.940 4.520 3.110 4.790 ;
        RECT 3.870 4.520 4.150 4.790 ;
        RECT 4.550 4.520 4.720 4.790 ;
        RECT 5.480 4.520 5.740 4.790 ;
        RECT 6.160 4.520 6.330 4.790 ;
        RECT 7.090 4.520 7.360 4.790 ;
        RECT 7.770 4.520 7.940 4.790 ;
        RECT 0.370 4.390 0.540 4.410 ;
        RECT 2.370 3.890 2.540 4.520 ;
        RECT 3.030 3.890 3.200 4.460 ;
        RECT 3.980 3.890 4.150 4.520 ;
        RECT 4.660 3.890 4.830 4.420 ;
        RECT 5.570 3.890 5.740 4.520 ;
        RECT 6.260 3.890 6.430 4.500 ;
        RECT 7.190 3.890 7.360 4.520 ;
        RECT 7.880 3.890 8.050 4.450 ;
        RECT 8.810 3.890 8.980 4.790 ;
        RECT 10.310 4.520 10.580 4.790 ;
        RECT 10.990 4.520 11.160 4.790 ;
        RECT 11.920 4.520 12.190 4.790 ;
        RECT 12.600 4.520 12.770 4.790 ;
        RECT 13.530 4.520 13.800 4.790 ;
        RECT 14.210 4.660 14.380 4.850 ;
        RECT 14.210 4.520 14.480 4.660 ;
        RECT 9.480 3.890 9.650 4.500 ;
        RECT 9.930 4.000 10.140 4.430 ;
        RECT 9.950 3.980 10.120 4.000 ;
        RECT 10.410 3.890 10.580 4.520 ;
        RECT 11.100 3.890 11.270 4.500 ;
        RECT 12.020 3.890 12.190 4.520 ;
        RECT 12.700 3.890 12.870 4.480 ;
        RECT 13.630 3.890 13.800 4.520 ;
        RECT 14.310 3.890 14.480 4.520 ;
        RECT 0.370 3.460 0.580 3.890 ;
        RECT 2.260 3.560 2.540 3.890 ;
        RECT 2.940 3.560 3.200 3.890 ;
        RECT 3.870 3.560 4.150 3.890 ;
        RECT 4.550 3.560 4.830 3.890 ;
        RECT 5.480 3.560 5.740 3.890 ;
        RECT 6.160 3.560 6.430 3.890 ;
        RECT 7.090 3.560 7.360 3.890 ;
        RECT 7.770 3.560 8.050 3.890 ;
        RECT 8.700 3.560 8.980 3.890 ;
        RECT 9.380 3.560 9.650 3.890 ;
        RECT 10.310 3.560 10.580 3.890 ;
        RECT 10.990 3.560 11.270 3.890 ;
        RECT 11.920 3.560 12.190 3.890 ;
        RECT 12.600 3.560 12.870 3.890 ;
        RECT 13.530 3.560 13.800 3.890 ;
        RECT 14.210 3.560 14.480 3.890 ;
        RECT 0.390 3.440 0.560 3.460 ;
        RECT 0.370 2.520 0.580 2.950 ;
        RECT 0.390 2.500 0.560 2.520 ;
        RECT 2.370 1.230 2.540 3.560 ;
        RECT 3.030 0.330 3.200 3.560 ;
        RECT 3.980 1.230 4.150 3.560 ;
        RECT 4.660 0.330 4.830 3.560 ;
        RECT 5.570 1.230 5.740 3.560 ;
        RECT 6.260 0.330 6.430 3.560 ;
        RECT 7.190 1.230 7.360 3.560 ;
        RECT 7.880 0.330 8.050 3.560 ;
        RECT 8.810 1.250 8.980 3.560 ;
        RECT 9.480 0.330 9.650 3.560 ;
        RECT 10.410 1.260 10.580 3.560 ;
        RECT 11.100 0.330 11.270 3.560 ;
        RECT 12.020 1.250 12.190 3.560 ;
        RECT 12.700 0.330 12.870 3.560 ;
        RECT 13.630 1.220 13.800 3.560 ;
        RECT 14.310 0.330 14.480 3.560 ;
        RECT 3.030 0.100 3.320 0.330 ;
        RECT 4.660 0.100 4.940 0.330 ;
        RECT 6.260 0.100 6.540 0.330 ;
        RECT 7.880 0.100 8.160 0.330 ;
        RECT 9.480 0.100 9.760 0.330 ;
        RECT 11.100 0.100 11.380 0.330 ;
        RECT 12.700 0.100 12.980 0.330 ;
        RECT 14.310 0.100 14.590 0.330 ;
        RECT 3.030 0.000 3.200 0.100 ;
        RECT 4.660 0.000 4.830 0.100 ;
        RECT 6.260 0.000 6.430 0.100 ;
        RECT 7.880 0.000 8.050 0.100 ;
        RECT 9.480 0.000 9.650 0.100 ;
        RECT 11.100 0.000 11.270 0.100 ;
        RECT 12.700 0.000 12.870 0.100 ;
        RECT 14.310 0.000 14.480 0.100 ;
      LAYER mcon ;
        RECT 13.040 5.720 13.210 5.890 ;
        RECT 13.710 5.720 13.880 5.890 ;
        RECT 8.370 5.140 8.540 5.310 ;
        RECT 3.140 0.130 3.310 0.300 ;
        RECT 4.760 0.130 4.930 0.300 ;
        RECT 6.360 0.130 6.530 0.300 ;
        RECT 7.980 0.130 8.150 0.300 ;
        RECT 9.580 0.130 9.750 0.300 ;
        RECT 11.200 0.130 11.370 0.300 ;
        RECT 12.800 0.130 12.970 0.300 ;
        RECT 14.410 0.130 14.580 0.300 ;
      LAYER met1 ;
        RECT 6.770 6.500 6.990 6.720 ;
        RECT 6.760 6.240 6.990 6.500 ;
        RECT 0.320 5.870 0.640 6.190 ;
        RECT 2.030 5.910 2.350 6.230 ;
        RECT 5.230 5.910 5.550 6.230 ;
        RECT 6.760 6.210 7.160 6.240 ;
        RECT 6.840 5.920 7.160 6.210 ;
        RECT 0.360 5.640 0.590 5.870 ;
        RECT 2.070 5.680 2.300 5.910 ;
        RECT 5.270 5.680 5.500 5.910 ;
        RECT 6.880 5.690 7.110 5.920 ;
        RECT 8.460 5.910 8.780 6.230 ;
        RECT 10.070 5.920 10.390 6.240 ;
        RECT 11.680 5.920 12.000 6.240 ;
        RECT 8.500 5.680 8.730 5.910 ;
        RECT 10.110 5.690 10.340 5.920 ;
        RECT 11.720 5.690 11.950 5.920 ;
        RECT 12.970 5.650 13.290 5.970 ;
        RECT 13.640 5.650 13.960 5.970 ;
        RECT 3.750 5.430 4.070 5.470 ;
        RECT 3.520 5.200 4.070 5.430 ;
        RECT 3.750 5.150 4.070 5.200 ;
        RECT 8.340 5.080 8.570 5.370 ;
        RECT 0.300 4.560 0.620 4.880 ;
        RECT 8.350 4.860 8.570 5.080 ;
        RECT 0.340 4.330 0.570 4.560 ;
        RECT 9.930 4.210 10.150 4.430 ;
        RECT 0.320 3.610 0.640 3.930 ;
        RECT 9.920 3.920 10.150 4.210 ;
        RECT 0.360 3.380 0.590 3.610 ;
        RECT 6.740 3.550 10.190 3.720 ;
        RECT 0.320 2.670 0.640 2.990 ;
        RECT 0.360 2.440 0.590 2.670 ;
        RECT 8.290 1.140 8.470 2.560 ;
        RECT 9.990 1.710 10.190 3.550 ;
        RECT 8.290 1.020 8.640 1.140 ;
        RECT 8.380 0.820 8.640 1.020 ;
      LAYER via ;
        RECT 0.350 5.900 0.610 6.160 ;
        RECT 2.060 5.940 2.320 6.200 ;
        RECT 5.260 5.940 5.520 6.200 ;
        RECT 6.870 5.950 7.130 6.210 ;
        RECT 8.490 5.940 8.750 6.200 ;
        RECT 10.100 5.950 10.360 6.210 ;
        RECT 11.710 5.950 11.970 6.210 ;
        RECT 13.000 5.680 13.260 5.940 ;
        RECT 13.670 5.680 13.930 5.940 ;
        RECT 3.780 5.180 4.040 5.440 ;
        RECT 0.330 4.590 0.590 4.850 ;
        RECT 0.350 3.640 0.610 3.900 ;
        RECT 0.350 2.700 0.610 2.960 ;
        RECT 8.380 0.850 8.640 1.110 ;
      LAYER met2 ;
        RECT 0.320 3.610 0.640 3.930 ;
  END
END sky130_hilas_DAC5bit01

MACRO sky130_hilas_capacitorSize04
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize04 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.150 BY 7.320 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAP1TERM02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.400 3.900 5.750 4.180 ;
    END
  END CAP1TERM02
  PIN CAP2TERM02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.400 0.900 5.760 1.180 ;
    END
  END CAP2TERM02
  PIN CAP2TERM01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 0.900 0.280 1.180 ;
    END
  END CAP2TERM01
  PIN CAP1TERM01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 3.900 0.270 4.180 ;
    END
  END CAP1TERM01
  OBS
      LAYER met2 ;
        RECT 0.000 4.850 5.750 5.030 ;
        RECT 0.000 4.420 5.800 4.600 ;
        RECT 0.560 4.200 0.930 4.420 ;
        RECT 5.430 4.200 5.800 4.420 ;
        RECT 0.000 3.420 5.750 3.600 ;
        RECT 0.000 2.990 5.750 3.170 ;
        RECT 0.000 1.840 5.750 2.010 ;
        RECT 0.590 1.590 0.960 1.600 ;
        RECT 5.430 1.590 5.800 1.600 ;
        RECT 0.000 1.420 5.800 1.590 ;
        RECT 0.590 1.200 0.960 1.420 ;
        RECT 5.430 1.200 5.800 1.420 ;
        RECT 0.000 0.440 5.750 0.610 ;
        RECT 0.000 0.000 5.750 0.170 ;
      LAYER via2 ;
        RECT 0.610 4.260 0.890 4.540 ;
        RECT 5.480 4.260 5.760 4.540 ;
        RECT 0.640 1.260 0.920 1.540 ;
        RECT 5.480 1.260 5.760 1.540 ;
      LAYER met3 ;
        RECT 5.850 5.040 8.150 7.320 ;
        RECT 0.340 4.000 1.130 4.750 ;
        RECT 3.840 3.640 4.870 4.390 ;
        RECT 5.210 4.310 6.000 4.750 ;
        RECT 5.210 4.000 8.150 4.310 ;
        RECT 5.850 2.030 8.150 4.000 ;
        RECT 0.370 1.000 1.160 1.750 ;
        RECT 3.830 0.650 4.890 1.380 ;
        RECT 5.210 1.000 6.000 1.750 ;
      LAYER via3 ;
        RECT 0.530 4.150 0.960 4.630 ;
        RECT 5.400 4.150 5.830 4.630 ;
        RECT 0.560 1.150 0.990 1.630 ;
        RECT 5.400 1.150 5.830 1.630 ;
      LAYER met4 ;
        RECT 6.700 6.270 7.150 6.280 ;
        RECT 6.680 5.780 7.200 6.270 ;
        RECT 0.430 4.110 1.090 4.720 ;
        RECT 0.240 3.700 3.030 4.110 ;
        RECT 5.300 4.060 5.960 4.720 ;
        RECT 6.700 3.260 7.150 3.270 ;
        RECT 6.680 2.770 7.200 3.260 ;
        RECT 0.460 1.100 1.120 1.720 ;
        RECT 0.460 1.060 2.670 1.100 ;
        RECT 5.300 1.060 5.960 1.720 ;
        RECT 0.550 0.690 2.670 1.060 ;
  END
END sky130_hilas_capacitorSize04

MACRO sky130_hilas_capacitorArray01
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorArray01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.700 BY 14.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM2
    USE ANALOG ;
    PORT
      LAYER met3 ;
        RECT 35.230 2.200 36.380 3.840 ;
        RECT 35.680 2.190 36.380 2.200 ;
    END
  END CAPTERM2
  PIN CAPTERM1
    USE ANALOG ;
    ANTENNADIFFAREA 1.012300 ;
    PORT
      LAYER met3 ;
        RECT 11.250 5.740 11.630 6.030 ;
        RECT 11.170 4.490 11.710 5.740 ;
    END
  END CAPTERM1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 5.390 6.010 5.710 6.020 ;
        RECT 8.760 6.010 9.080 6.100 ;
        RECT 9.320 6.010 9.640 6.070 ;
        RECT 5.390 5.930 9.640 6.010 ;
        RECT 10.740 6.020 11.250 6.050 ;
        RECT 10.740 5.930 11.670 6.020 ;
        RECT 5.390 5.830 11.670 5.930 ;
        RECT 5.390 5.760 5.710 5.830 ;
        RECT 8.880 5.740 11.670 5.830 ;
        RECT 11.170 5.720 11.670 5.740 ;
      LAYER via2 ;
        RECT 11.300 5.720 11.580 6.000 ;
    END
  END VINJ
  PIN GATESELECT
    PORT
      LAYER met1 ;
        RECT 9.120 6.000 9.310 6.050 ;
    END
  END GATESELECT
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 0.360 5.910 0.760 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.360 0.000 0.750 0.120 ;
    END
  END VTUN
  PIN GATE
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 4.420 5.970 4.790 6.050 ;
        RECT 4.410 5.920 4.790 5.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.400 0.130 4.410 0.150 ;
        RECT 4.400 0.010 4.790 0.130 ;
        RECT 4.400 0.000 4.410 0.010 ;
    END
  END GATE
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 0.000 3.510 0.120 3.690 ;
    END
    PORT
      LAYER met2 ;
        RECT 35.690 3.690 36.700 3.700 ;
        RECT 8.940 3.510 36.700 3.690 ;
    END
  END DRAIN2
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 0.010 5.370 0.120 5.550 ;
    END
    PORT
      LAYER met2 ;
        RECT 8.980 5.400 36.700 5.550 ;
        RECT 2.640 5.370 36.700 5.400 ;
        RECT 2.640 5.220 10.260 5.370 ;
    END
  END DRAIN1
  PIN DRAIN4
    PORT
      LAYER met2 ;
        RECT 8.810 0.520 36.700 0.690 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.020 0.520 0.120 0.690 ;
    END
  END DRAIN4
  PIN DRAIN3
    PORT
      LAYER met4 ;
        RECT 10.070 2.300 10.730 2.680 ;
        RECT 13.710 2.300 16.900 2.330 ;
        RECT 19.350 2.300 19.650 2.330 ;
        RECT 10.070 2.020 22.570 2.300 ;
        RECT 10.370 2.000 22.570 2.020 ;
        RECT 13.710 1.630 14.010 2.000 ;
        RECT 16.600 1.660 16.900 2.000 ;
        RECT 19.350 1.660 19.650 2.000 ;
        RECT 16.600 1.630 19.650 1.660 ;
        RECT 22.270 1.630 22.570 2.000 ;
        RECT 13.710 1.330 22.570 1.630 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.020 2.360 0.120 2.530 ;
    END
  END DRAIN3
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2.990 6.050 3.390 10.730 ;
        RECT 2.800 5.990 3.390 6.050 ;
        RECT 2.990 4.230 3.390 5.990 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.730 5.980 6.970 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.800 0.000 3.040 0.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.730 0.000 6.970 0.070 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 17.150 14.670 18.880 14.720 ;
        RECT 2.640 9.390 2.710 9.570 ;
        RECT 13.040 9.230 15.600 11.140 ;
        RECT 3.210 9.040 3.800 9.150 ;
        RECT 6.950 8.980 8.060 9.210 ;
        RECT 11.590 7.550 11.940 7.560 ;
        RECT 11.590 7.390 11.760 7.550 ;
        RECT 11.930 7.390 11.940 7.550 ;
        RECT 13.040 6.050 15.600 8.960 ;
        RECT 15.960 8.230 18.880 14.670 ;
        RECT 21.150 11.140 22.880 12.980 ;
        RECT 15.960 8.180 18.190 8.230 ;
        RECT 10.070 6.040 35.420 6.050 ;
        RECT 3.210 5.760 3.800 5.950 ;
        RECT 6.950 5.740 8.060 6.010 ;
        RECT 10.080 5.970 35.420 6.040 ;
        RECT 0.010 5.370 0.120 5.550 ;
        RECT 0.000 3.510 0.120 3.690 ;
        RECT 0.020 0.520 0.120 0.690 ;
        RECT 10.060 0.060 35.420 5.970 ;
        RECT 10.070 0.010 35.420 0.060 ;
        RECT 12.000 0.000 35.420 0.010 ;
      LAYER li1 ;
        RECT 17.540 11.660 18.090 12.090 ;
        RECT 21.570 11.590 22.120 12.020 ;
        RECT 13.280 10.790 13.600 10.830 ;
        RECT 13.280 10.670 13.610 10.790 ;
        RECT 13.280 10.570 13.720 10.670 ;
        RECT 13.380 10.500 13.720 10.570 ;
        RECT 15.000 10.400 15.200 10.750 ;
        RECT 13.280 10.240 13.600 10.280 ;
        RECT 13.280 10.050 13.610 10.240 ;
        RECT 13.280 10.020 13.720 10.050 ;
        RECT 13.380 9.880 13.720 10.020 ;
        RECT 14.270 9.780 14.470 10.380 ;
        RECT 15.000 10.370 15.210 10.400 ;
        RECT 14.990 9.780 15.210 10.370 ;
        RECT 5.460 8.750 5.630 9.280 ;
        RECT 9.400 8.740 9.570 9.270 ;
        RECT 13.380 8.170 13.720 8.310 ;
        RECT 13.280 8.140 13.720 8.170 ;
        RECT 5.470 7.040 5.640 8.050 ;
        RECT 13.280 7.950 13.610 8.140 ;
        RECT 13.280 7.910 13.600 7.950 ;
        RECT 9.400 6.900 9.570 7.910 ;
        RECT 14.270 7.810 14.470 8.410 ;
        RECT 14.990 7.820 15.210 8.410 ;
        RECT 15.000 7.790 15.210 7.820 ;
        RECT 13.380 7.620 13.720 7.690 ;
        RECT 11.500 7.390 11.940 7.560 ;
        RECT 13.280 7.520 13.720 7.620 ;
        RECT 13.280 7.430 13.610 7.520 ;
        RECT 13.280 7.330 13.720 7.430 ;
        RECT 13.380 7.260 13.720 7.330 ;
        RECT 15.000 7.160 15.200 7.790 ;
        RECT 13.280 7.000 13.600 7.040 ;
        RECT 13.280 6.810 13.610 7.000 ;
        RECT 13.280 6.780 13.720 6.810 ;
        RECT 13.380 6.640 13.720 6.780 ;
        RECT 14.270 6.540 14.470 7.140 ;
        RECT 15.000 7.130 15.210 7.160 ;
        RECT 14.990 6.540 15.210 7.130 ;
        RECT 13.380 4.940 13.720 5.080 ;
        RECT 13.280 4.910 13.720 4.940 ;
        RECT 13.280 4.720 13.610 4.910 ;
        RECT 13.280 4.680 13.600 4.720 ;
        RECT 14.270 4.580 14.470 5.180 ;
        RECT 14.990 4.590 15.210 5.180 ;
        RECT 15.000 4.560 15.210 4.590 ;
        RECT 13.380 4.390 13.720 4.460 ;
        RECT 13.280 4.290 13.720 4.390 ;
        RECT 13.280 4.170 13.610 4.290 ;
        RECT 15.000 4.210 15.200 4.560 ;
        RECT 13.280 4.130 13.600 4.170 ;
      LAYER mcon ;
        RECT 17.540 11.740 17.810 12.010 ;
        RECT 21.570 11.670 21.840 11.940 ;
        RECT 13.340 10.610 13.510 10.780 ;
        RECT 13.340 10.060 13.510 10.230 ;
        RECT 14.280 10.170 14.450 10.340 ;
        RECT 15.010 10.200 15.180 10.370 ;
        RECT 5.460 9.110 5.630 9.280 ;
        RECT 9.400 9.100 9.570 9.270 ;
        RECT 13.340 7.960 13.510 8.130 ;
        RECT 5.470 7.650 5.640 7.820 ;
        RECT 5.470 7.290 5.640 7.460 ;
        RECT 14.280 7.850 14.450 8.020 ;
        RECT 15.010 7.820 15.180 7.990 ;
        RECT 9.400 7.510 9.570 7.680 ;
        RECT 11.760 7.390 11.940 7.560 ;
        RECT 13.340 7.370 13.510 7.580 ;
        RECT 9.400 7.150 9.570 7.320 ;
        RECT 13.340 6.820 13.510 6.990 ;
        RECT 14.280 6.930 14.450 7.100 ;
        RECT 15.010 6.960 15.180 7.130 ;
        RECT 13.340 4.730 13.510 4.900 ;
        RECT 14.280 4.620 14.450 4.790 ;
        RECT 15.010 4.590 15.180 4.760 ;
        RECT 13.340 4.180 13.510 4.350 ;
      LAYER met1 ;
        RECT 5.430 9.320 5.670 10.730 ;
        RECT 7.040 10.400 7.420 10.730 ;
        RECT 9.360 9.340 9.600 10.730 ;
        RECT 13.270 10.540 13.590 10.860 ;
        RECT 11.380 10.460 11.540 10.500 ;
        RECT 11.750 10.450 11.940 10.500 ;
        RECT 12.190 10.450 12.350 10.500 ;
        RECT 14.270 10.400 14.430 11.130 ;
        RECT 14.270 10.380 14.470 10.400 ;
        RECT 13.270 9.990 13.590 10.310 ;
        RECT 14.250 10.140 14.480 10.380 ;
        RECT 14.270 10.090 14.480 10.140 ;
        RECT 14.640 10.090 14.830 11.080 ;
        RECT 15.080 10.430 15.240 11.130 ;
        RECT 5.420 8.660 5.680 9.320 ;
        RECT 9.340 8.680 9.610 9.340 ;
        RECT 14.270 9.230 14.430 10.090 ;
        RECT 14.660 9.970 14.830 10.090 ;
        RECT 14.670 9.230 14.830 9.970 ;
        RECT 14.970 9.880 15.240 10.430 ;
        RECT 14.970 9.830 15.250 9.880 ;
        RECT 15.080 9.740 15.250 9.830 ;
        RECT 15.080 9.230 15.240 9.740 ;
        RECT 5.430 6.050 5.670 8.660 ;
        RECT 5.420 5.730 5.680 6.050 ;
        RECT 8.790 5.810 9.050 6.130 ;
        RECT 9.360 6.090 9.600 8.680 ;
        RECT 13.270 7.880 13.590 8.200 ;
        RECT 14.270 8.100 14.430 8.960 ;
        RECT 14.670 8.220 14.830 8.960 ;
        RECT 15.080 8.450 15.240 8.960 ;
        RECT 15.080 8.360 15.250 8.450 ;
        RECT 14.660 8.100 14.830 8.220 ;
        RECT 14.270 8.050 14.480 8.100 ;
        RECT 14.250 7.810 14.480 8.050 ;
        RECT 14.270 7.790 14.470 7.810 ;
        RECT 11.810 7.590 11.940 7.610 ;
        RECT 11.730 7.570 11.970 7.590 ;
        RECT 11.530 7.380 11.970 7.570 ;
        RECT 11.730 7.360 11.970 7.380 ;
        RECT 11.830 7.320 11.940 7.360 ;
        RECT 13.270 7.300 13.590 7.650 ;
        RECT 14.270 7.160 14.430 7.790 ;
        RECT 14.270 7.140 14.470 7.160 ;
        RECT 13.270 6.750 13.590 7.070 ;
        RECT 14.250 6.900 14.480 7.140 ;
        RECT 14.270 6.850 14.480 6.900 ;
        RECT 14.640 6.850 14.830 8.100 ;
        RECT 14.970 8.310 15.250 8.360 ;
        RECT 14.970 7.760 15.240 8.310 ;
        RECT 16.610 8.180 16.990 14.680 ;
        RECT 17.480 11.200 17.870 13.060 ;
        RECT 21.510 11.130 21.900 12.990 ;
        RECT 15.080 7.190 15.240 7.760 ;
        RECT 9.350 6.050 9.610 6.090 ;
        RECT 9.350 6.000 9.720 6.050 ;
        RECT 9.350 5.770 9.610 6.000 ;
        RECT 14.270 5.990 14.430 6.850 ;
        RECT 14.660 6.730 14.830 6.850 ;
        RECT 14.670 5.990 14.830 6.730 ;
        RECT 14.970 6.640 15.240 7.190 ;
        RECT 14.970 6.590 15.250 6.640 ;
        RECT 15.080 6.500 15.250 6.590 ;
        RECT 15.080 5.990 15.240 6.500 ;
        RECT 5.430 4.230 5.670 5.730 ;
        RECT 7.040 4.230 7.420 4.830 ;
        RECT 9.360 4.230 9.600 5.770 ;
        RECT 13.270 4.650 13.590 4.970 ;
        RECT 14.270 4.870 14.430 5.730 ;
        RECT 14.670 4.990 14.830 5.730 ;
        RECT 15.080 5.220 15.240 5.730 ;
        RECT 15.080 5.130 15.250 5.220 ;
        RECT 14.660 4.870 14.830 4.990 ;
        RECT 14.270 4.820 14.480 4.870 ;
        RECT 14.250 4.580 14.480 4.820 ;
        RECT 14.270 4.560 14.470 4.580 ;
        RECT 13.270 4.100 13.590 4.420 ;
        RECT 14.270 3.830 14.430 4.560 ;
        RECT 14.640 3.880 14.830 4.870 ;
        RECT 14.970 5.080 15.250 5.130 ;
        RECT 14.970 4.530 15.240 5.080 ;
        RECT 15.080 3.830 15.240 4.530 ;
        RECT 8.750 0.010 8.910 0.070 ;
        RECT 9.120 0.010 9.310 0.070 ;
        RECT 9.560 0.010 9.720 0.070 ;
      LAYER via ;
        RECT 13.300 10.570 13.560 10.830 ;
        RECT 13.300 10.020 13.560 10.280 ;
        RECT 5.420 5.760 5.680 6.020 ;
        RECT 8.790 5.840 9.050 6.100 ;
        RECT 13.300 7.910 13.560 8.170 ;
        RECT 13.300 7.330 13.560 7.620 ;
        RECT 13.300 6.780 13.560 7.040 ;
        RECT 9.350 5.800 9.610 6.060 ;
        RECT 13.300 4.680 13.560 4.940 ;
        RECT 13.300 4.130 13.560 4.390 ;
      LAYER met2 ;
        RECT 13.270 10.580 13.580 10.870 ;
        RECT 13.270 10.540 15.600 10.580 ;
        RECT 13.420 10.400 15.600 10.540 ;
        RECT 2.640 9.990 10.270 10.170 ;
        RECT 13.270 10.150 13.580 10.320 ;
        RECT 13.040 9.970 13.130 10.150 ;
        RECT 13.270 9.990 15.600 10.150 ;
        RECT 13.430 9.970 15.600 9.990 ;
        RECT 2.640 9.550 10.270 9.730 ;
        RECT 2.640 8.450 10.270 8.630 ;
        RECT 2.640 8.020 10.270 8.200 ;
        RECT 13.040 8.040 13.130 8.220 ;
        RECT 13.430 8.200 15.600 8.220 ;
        RECT 13.270 8.040 15.600 8.200 ;
        RECT 13.270 7.870 13.580 8.040 ;
        RECT 13.420 7.650 15.600 7.790 ;
        RECT 13.270 7.610 15.600 7.650 ;
        RECT 13.270 7.340 13.580 7.610 ;
        RECT 13.270 7.300 15.600 7.340 ;
        RECT 13.420 7.160 15.600 7.300 ;
        RECT 2.640 6.750 10.260 6.930 ;
        RECT 13.270 6.910 13.580 7.080 ;
        RECT 13.040 6.730 13.130 6.910 ;
        RECT 13.270 6.750 15.600 6.910 ;
        RECT 13.430 6.730 15.600 6.750 ;
        RECT 2.640 6.320 10.270 6.500 ;
        RECT 8.920 4.970 36.700 5.120 ;
        RECT 2.640 4.940 36.700 4.970 ;
        RECT 2.640 4.800 10.240 4.940 ;
        RECT 13.040 4.810 13.130 4.940 ;
        RECT 13.270 4.810 15.600 4.940 ;
        RECT 10.240 4.250 10.610 4.650 ;
        RECT 13.270 4.640 13.580 4.810 ;
        RECT 13.420 4.420 15.600 4.560 ;
        RECT 13.270 4.380 15.600 4.420 ;
        RECT 13.270 4.120 13.580 4.380 ;
        RECT 8.980 3.940 36.700 4.120 ;
        RECT 36.010 2.790 36.700 3.200 ;
        RECT 10.200 2.530 10.570 2.560 ;
        RECT 8.770 2.360 36.700 2.530 ;
        RECT 10.200 2.160 10.570 2.360 ;
        RECT 8.870 1.940 36.700 2.110 ;
        RECT 11.290 1.290 11.660 1.690 ;
        RECT 8.850 0.960 36.700 1.130 ;
      LAYER via2 ;
        RECT 10.290 4.310 10.570 4.590 ;
        RECT 36.080 2.850 36.370 3.130 ;
        RECT 10.250 2.220 10.530 2.500 ;
        RECT 11.340 1.350 11.620 1.630 ;
      LAYER met3 ;
        RECT 10.020 4.050 10.810 4.800 ;
        RECT 9.980 1.960 10.770 2.710 ;
        RECT 11.070 1.090 11.860 1.840 ;
        RECT 11.460 0.790 11.640 1.090 ;
      LAYER via3 ;
        RECT 10.210 4.200 10.640 4.680 ;
        RECT 10.170 2.110 10.600 2.590 ;
        RECT 11.260 1.240 11.690 1.720 ;
      LAYER met4 ;
        RECT 12.790 5.380 16.890 5.680 ;
        RECT 11.100 4.770 13.800 4.880 ;
        RECT 10.110 4.110 10.770 4.770 ;
        RECT 11.100 4.470 14.010 4.770 ;
        RECT 13.500 4.130 14.010 4.470 ;
        RECT 16.510 4.180 16.890 5.380 ;
        RECT 19.350 4.210 22.630 4.510 ;
        RECT 10.410 3.750 11.770 4.050 ;
        RECT 11.470 3.190 11.770 3.750 ;
        RECT 19.350 3.190 19.650 4.210 ;
        RECT 22.330 3.190 22.630 4.210 ;
        RECT 11.470 2.890 22.630 3.190 ;
        RECT 25.030 4.190 33.920 4.490 ;
        RECT 11.160 1.150 11.820 1.810 ;
        RECT 25.030 1.670 25.330 4.190 ;
        RECT 27.860 4.160 30.970 4.190 ;
        RECT 27.860 1.670 28.160 4.160 ;
        RECT 30.670 1.670 30.970 4.160 ;
        RECT 33.620 1.670 33.920 4.190 ;
        RECT 25.030 1.370 33.980 1.670 ;
        RECT 30.670 1.360 33.980 1.370 ;
        RECT 11.340 0.790 11.850 1.090 ;
        RECT 11.550 0.550 11.850 0.790 ;
        RECT 33.680 0.550 33.980 1.360 ;
        RECT 11.550 0.250 33.980 0.550 ;
  END
END sky130_hilas_capacitorArray01

MACRO sky130_hilas_pFETmed
  CLASS CORE ;
  FOREIGN sky130_hilas_pFETmed ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.190 BY 2.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 0.000 0.000 1.190 2.870 ;
      LAYER li1 ;
        RECT 0.240 0.150 0.410 2.640 ;
        RECT 0.790 0.140 0.960 2.640 ;
  END
END sky130_hilas_pFETmed

MACRO sky130_hilas_swc4x1cellOverlap2
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x1cellOverlap2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.240 BY 7.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 8.000 6.980 12.000 7.050 ;
        RECT 8.000 5.070 12.240 6.980 ;
        RECT 8.000 4.910 12.000 5.070 ;
        RECT 8.000 2.060 12.240 4.910 ;
        RECT 8.000 1.910 12.000 2.060 ;
        RECT 8.000 1.000 12.240 1.910 ;
        RECT 9.680 0.000 12.240 1.000 ;
      LAYER li1 ;
        RECT 1.680 5.730 1.850 6.620 ;
        RECT 8.350 6.590 11.660 6.720 ;
        RECT 8.350 6.240 11.840 6.590 ;
        RECT 8.350 5.740 11.850 6.240 ;
        RECT 10.020 5.720 10.360 5.740 ;
        RECT 10.910 5.620 11.110 5.740 ;
        RECT 11.630 5.620 11.850 5.740 ;
        RECT 1.680 4.210 1.850 5.100 ;
        RECT 8.350 4.360 11.660 5.250 ;
        RECT 8.350 4.270 11.850 4.360 ;
        RECT 10.020 4.120 10.360 4.260 ;
        RECT 9.920 4.090 10.360 4.120 ;
        RECT 9.920 3.900 10.250 4.090 ;
        RECT 9.920 3.860 10.240 3.900 ;
        RECT 10.910 3.780 11.110 4.270 ;
        RECT 11.630 3.780 11.850 4.270 ;
        RECT 8.350 3.740 11.850 3.780 ;
        RECT 1.680 2.760 1.850 3.650 ;
        RECT 8.350 3.570 11.840 3.740 ;
        RECT 8.140 3.400 11.840 3.570 ;
        RECT 8.350 3.230 11.840 3.400 ;
        RECT 8.350 2.800 11.850 3.230 ;
        RECT 10.020 2.710 10.360 2.800 ;
        RECT 10.910 2.610 11.110 2.800 ;
        RECT 11.630 2.610 11.850 2.800 ;
        RECT 1.680 1.220 1.850 2.110 ;
        RECT 8.350 1.360 11.660 2.310 ;
        RECT 8.350 1.330 11.850 1.360 ;
        RECT 10.020 1.120 10.360 1.260 ;
        RECT 9.920 1.090 10.360 1.120 ;
        RECT 9.920 0.900 10.250 1.090 ;
        RECT 9.920 0.860 10.240 0.900 ;
        RECT 10.910 0.760 11.110 1.330 ;
        RECT 11.630 0.770 11.850 1.330 ;
        RECT 11.640 0.740 11.850 0.770 ;
        RECT 10.020 0.570 10.360 0.640 ;
        RECT 9.920 0.470 10.360 0.570 ;
        RECT 9.920 0.350 10.250 0.470 ;
        RECT 11.640 0.390 11.840 0.740 ;
        RECT 9.920 0.310 10.240 0.350 ;
      LAYER mcon ;
        RECT 1.680 6.420 1.850 6.590 ;
        RECT 9.920 6.620 10.090 6.660 ;
        RECT 9.920 6.490 10.150 6.620 ;
        RECT 9.980 6.450 10.150 6.490 ;
        RECT 9.980 5.970 10.150 6.070 ;
        RECT 10.920 6.010 11.090 6.180 ;
        RECT 11.650 6.040 11.820 6.210 ;
        RECT 9.920 5.900 10.150 5.970 ;
        RECT 9.920 5.800 10.090 5.900 ;
        RECT 1.680 4.900 1.850 5.070 ;
        RECT 9.920 5.020 10.090 5.190 ;
        RECT 9.920 4.330 10.090 4.500 ;
        RECT 9.980 3.910 10.150 4.080 ;
        RECT 10.920 3.800 11.090 3.970 ;
        RECT 11.650 3.770 11.820 3.940 ;
        RECT 1.680 3.450 1.850 3.620 ;
        RECT 9.920 3.610 10.090 3.720 ;
        RECT 8.400 3.400 8.580 3.570 ;
        RECT 9.920 3.550 10.150 3.610 ;
        RECT 9.980 3.360 10.150 3.550 ;
        RECT 9.980 3.030 10.150 3.060 ;
        RECT 9.920 2.890 10.150 3.030 ;
        RECT 10.920 3.000 11.090 3.170 ;
        RECT 11.650 3.030 11.820 3.200 ;
        RECT 9.920 2.860 10.090 2.890 ;
        RECT 1.680 1.910 1.850 2.080 ;
        RECT 9.920 2.080 10.090 2.250 ;
        RECT 9.920 1.390 10.090 1.560 ;
        RECT 9.980 0.910 10.150 1.080 ;
        RECT 10.920 0.800 11.090 0.970 ;
        RECT 11.650 0.770 11.820 0.940 ;
        RECT 9.980 0.360 10.150 0.530 ;
      LAYER met1 ;
        RECT 1.010 0.460 1.280 6.510 ;
        RECT 1.650 5.520 1.880 6.810 ;
        RECT 9.880 6.700 10.120 6.720 ;
        RECT 9.880 6.380 10.230 6.700 ;
        RECT 9.880 6.150 10.120 6.380 ;
        RECT 10.910 6.240 11.070 6.970 ;
        RECT 10.910 6.220 11.110 6.240 ;
        RECT 9.880 6.080 10.230 6.150 ;
        RECT 9.890 5.830 10.230 6.080 ;
        RECT 10.890 5.980 11.120 6.220 ;
        RECT 10.910 5.930 11.120 5.980 ;
        RECT 11.280 5.930 11.470 6.920 ;
        RECT 11.720 6.270 11.880 6.970 ;
        RECT 9.890 5.820 10.120 5.830 ;
        RECT 9.890 5.600 10.130 5.820 ;
        RECT 1.650 4.000 1.880 5.290 ;
        RECT 9.880 4.610 10.120 5.250 ;
        RECT 10.910 5.070 11.070 5.930 ;
        RECT 11.300 5.810 11.470 5.930 ;
        RECT 11.310 5.070 11.470 5.810 ;
        RECT 11.610 5.720 11.880 6.270 ;
        RECT 11.610 5.670 11.890 5.720 ;
        RECT 11.720 5.580 11.890 5.670 ;
        RECT 11.720 5.070 11.880 5.580 ;
        RECT 9.890 4.350 10.120 4.610 ;
        RECT 9.890 4.150 10.130 4.350 ;
        RECT 9.890 4.130 10.230 4.150 ;
        RECT 1.650 2.550 1.880 3.840 ;
        RECT 9.910 3.830 10.230 4.130 ;
        RECT 10.910 4.050 11.070 4.910 ;
        RECT 11.310 4.170 11.470 4.910 ;
        RECT 11.720 4.400 11.880 4.910 ;
        RECT 11.720 4.310 11.890 4.400 ;
        RECT 11.300 4.050 11.470 4.170 ;
        RECT 10.910 4.000 11.120 4.050 ;
        RECT 9.880 3.690 10.120 3.780 ;
        RECT 10.890 3.760 11.120 4.000 ;
        RECT 10.910 3.740 11.110 3.760 ;
        RECT 8.450 3.600 8.580 3.620 ;
        RECT 8.370 3.370 8.610 3.600 ;
        RECT 8.470 3.330 8.580 3.370 ;
        RECT 9.880 3.280 10.230 3.690 ;
        RECT 9.880 3.140 10.120 3.280 ;
        RECT 10.910 3.230 11.070 3.740 ;
        RECT 10.910 3.210 11.110 3.230 ;
        RECT 9.890 2.820 10.230 3.140 ;
        RECT 10.890 2.970 11.120 3.210 ;
        RECT 10.910 2.920 11.120 2.970 ;
        RECT 11.280 2.920 11.470 4.050 ;
        RECT 11.610 4.260 11.890 4.310 ;
        RECT 11.610 3.710 11.880 4.260 ;
        RECT 11.720 3.260 11.880 3.710 ;
        RECT 9.890 2.660 10.130 2.820 ;
        RECT 1.650 1.010 1.880 2.300 ;
        RECT 9.880 1.670 10.120 2.310 ;
        RECT 10.910 2.060 11.070 2.920 ;
        RECT 11.300 2.800 11.470 2.920 ;
        RECT 11.310 2.060 11.470 2.800 ;
        RECT 11.610 2.710 11.880 3.260 ;
        RECT 11.610 2.660 11.890 2.710 ;
        RECT 11.720 2.570 11.890 2.660 ;
        RECT 11.720 2.060 11.880 2.570 ;
        RECT 9.890 1.410 10.120 1.670 ;
        RECT 9.890 1.190 10.130 1.410 ;
        RECT 9.910 0.830 10.230 1.150 ;
        RECT 10.910 1.050 11.070 1.910 ;
        RECT 11.310 1.170 11.470 1.910 ;
        RECT 11.720 1.400 11.880 1.910 ;
        RECT 11.720 1.310 11.890 1.400 ;
        RECT 11.300 1.050 11.470 1.170 ;
        RECT 10.910 1.000 11.120 1.050 ;
        RECT 10.890 0.760 11.120 1.000 ;
        RECT 10.910 0.740 11.110 0.760 ;
        RECT 9.910 0.280 10.230 0.600 ;
        RECT 10.910 0.010 11.070 0.740 ;
        RECT 11.280 0.060 11.470 1.050 ;
        RECT 11.610 1.260 11.890 1.310 ;
        RECT 11.610 0.710 11.880 1.260 ;
        RECT 11.720 0.010 11.880 0.710 ;
      LAYER via ;
        RECT 9.940 6.410 10.200 6.670 ;
        RECT 9.940 5.860 10.200 6.120 ;
        RECT 9.940 3.860 10.200 4.120 ;
        RECT 9.940 3.310 10.200 3.660 ;
        RECT 9.940 2.850 10.200 3.110 ;
        RECT 9.940 0.860 10.200 1.120 ;
        RECT 9.940 0.310 10.200 0.570 ;
      LAYER met2 ;
        RECT 9.910 6.420 10.220 6.710 ;
        RECT 9.910 6.380 12.240 6.420 ;
        RECT 10.060 6.240 12.240 6.380 ;
        RECT 0.000 5.940 6.880 6.010 ;
        RECT 9.910 5.990 10.220 6.160 ;
        RECT 0.000 5.830 6.910 5.940 ;
        RECT 9.680 5.810 9.770 5.990 ;
        RECT 9.910 5.830 12.240 5.990 ;
        RECT 10.070 5.810 12.240 5.830 ;
        RECT 0.000 5.400 9.010 5.580 ;
        RECT 0.000 4.520 6.880 4.580 ;
        RECT 0.000 4.400 6.910 4.520 ;
        RECT 0.000 4.080 6.870 4.150 ;
        RECT 0.000 3.970 6.910 4.080 ;
        RECT 9.680 3.990 9.770 4.170 ;
        RECT 10.070 4.150 12.240 4.170 ;
        RECT 9.910 3.990 12.240 4.150 ;
        RECT 9.910 3.820 10.220 3.990 ;
        RECT 10.060 3.700 12.240 3.740 ;
        RECT 9.910 3.560 12.240 3.700 ;
        RECT 9.910 3.410 10.220 3.560 ;
        RECT 9.910 3.270 12.240 3.410 ;
        RECT 10.060 3.230 12.240 3.270 ;
        RECT 0.000 2.820 6.910 2.990 ;
        RECT 9.910 2.980 10.220 3.150 ;
        RECT 9.680 2.800 9.770 2.980 ;
        RECT 9.910 2.820 12.240 2.980 ;
        RECT 10.070 2.800 12.240 2.820 ;
        RECT 0.000 2.400 6.910 2.570 ;
        RECT 0.000 1.420 6.910 1.590 ;
        RECT 0.000 0.980 6.910 1.150 ;
        RECT 9.680 0.990 9.770 1.170 ;
        RECT 10.070 1.150 12.240 1.170 ;
        RECT 9.910 0.990 12.240 1.150 ;
        RECT 9.910 0.820 10.220 0.990 ;
        RECT 10.060 0.600 12.240 0.740 ;
        RECT 9.910 0.560 12.240 0.600 ;
        RECT 9.910 0.270 10.220 0.560 ;
  END
END sky130_hilas_swc4x1cellOverlap2

MACRO sky130_hilas_TA2SignalBiasCell
  CLASS CORE ;
  FOREIGN sky130_hilas_TA2SignalBiasCell ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.810 BY 24.010 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VOUT_AMP2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 9.630 12.320 9.780 12.540 ;
    END
  END VOUT_AMP2
  PIN VOUT_AMP1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 9.630 11.500 9.780 11.720 ;
    END
  END VOUT_AMP1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 7.820 8.980 8.160 9.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 7.820 14.890 8.160 15.030 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 8.490 8.980 8.760 9.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.490 14.880 8.760 15.030 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.900 15.020 2.810 15.030 ;
        RECT 0.900 9.420 6.500 15.020 ;
        RECT 10.480 9.470 11.760 12.310 ;
        RECT 0.900 9.240 1.330 9.420 ;
        RECT 0.900 9.010 1.610 9.240 ;
        RECT 0.900 8.990 1.330 9.010 ;
      LAYER met2 ;
        RECT 8.960 15.800 9.270 16.090 ;
        RECT 10.620 15.800 10.930 16.050 ;
        RECT 8.240 15.720 10.930 15.800 ;
        RECT 8.240 15.570 10.780 15.720 ;
        RECT 8.910 15.110 9.220 15.440 ;
        RECT 1.690 15.000 1.930 15.030 ;
        RECT 1.690 14.670 2.100 15.000 ;
        RECT 1.690 14.650 1.930 14.670 ;
        RECT 1.220 14.560 1.930 14.650 ;
        RECT 1.170 14.210 1.930 14.560 ;
        RECT 2.970 14.400 3.520 14.650 ;
        RECT 3.010 14.210 3.320 14.400 ;
        RECT 1.170 13.980 5.710 14.210 ;
        RECT 1.170 13.790 1.930 13.980 ;
        RECT 0.680 13.740 1.930 13.790 ;
        RECT 0.680 13.730 1.620 13.740 ;
        RECT 0.680 13.540 1.560 13.730 ;
        RECT 5.480 13.620 5.710 13.980 ;
        RECT 8.910 13.830 9.220 14.160 ;
        RECT 8.500 13.660 8.830 13.770 ;
        RECT 10.670 13.660 10.980 13.830 ;
        RECT 8.500 13.620 11.150 13.660 ;
        RECT 1.110 13.380 1.420 13.540 ;
        RECT 5.480 13.430 11.150 13.620 ;
        RECT 5.480 13.420 8.830 13.430 ;
        RECT 5.740 13.410 8.830 13.420 ;
        RECT 8.500 12.840 8.830 13.410 ;
        RECT 8.960 13.180 9.270 13.430 ;
        RECT 8.960 12.830 9.270 13.090 ;
        RECT 10.660 12.830 10.970 13.110 ;
        RECT 8.240 12.610 11.150 12.830 ;
        RECT 8.910 12.110 9.220 12.440 ;
        RECT 8.910 10.830 9.220 11.160 ;
        RECT 10.580 10.670 10.890 10.860 ;
        RECT 8.230 10.440 10.940 10.670 ;
        RECT 8.960 10.180 9.270 10.440 ;
    END
  END VPWR
  PIN VIN22
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.290 14.760 5.540 15.020 ;
    END
  END VIN22
  PIN VIN21
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.330 12.090 5.580 12.320 ;
    END
  END VIN21
  PIN VIN11
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 3.770 11.680 4.050 11.920 ;
    END
  END VIN11
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 3.730 9.000 3.990 9.250 ;
    END
  END VIN12
  PIN VBIAS2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.950 9.010 2.600 9.240 ;
    END
  END VBIAS2
  PIN VBIAS1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.910 11.680 2.370 11.920 ;
        RECT 0.910 11.670 1.550 11.680 ;
    END
  END VBIAS1
  OBS
      LAYER nwell ;
        RECT 3.630 21.020 7.240 24.010 ;
        RECT 3.630 17.970 7.240 20.960 ;
        RECT 0.000 16.520 3.610 16.590 ;
        RECT 1.340 16.230 1.790 16.460 ;
        RECT 3.090 16.230 3.540 16.460 ;
        RECT 8.500 14.850 9.780 15.030 ;
        RECT 10.480 13.930 11.760 16.770 ;
        RECT 8.500 8.980 9.780 9.170 ;
        RECT 4.650 7.550 5.100 7.780 ;
        RECT 3.310 7.420 5.170 7.490 ;
        RECT 6.940 3.050 8.800 6.040 ;
        RECT 6.940 0.000 8.800 2.990 ;
      LAYER li1 ;
        RECT 4.040 21.490 4.220 23.540 ;
        RECT 4.850 21.750 5.020 23.530 ;
        RECT 4.770 21.580 5.100 21.750 ;
        RECT 5.790 21.490 5.970 23.540 ;
        RECT 6.600 21.750 6.770 23.530 ;
        RECT 6.520 21.580 6.850 21.750 ;
        RECT 4.040 18.440 4.220 20.490 ;
        RECT 4.850 18.700 5.020 20.480 ;
        RECT 4.770 18.530 5.100 18.700 ;
        RECT 5.790 18.440 5.970 20.490 ;
        RECT 6.600 18.700 6.770 20.480 ;
        RECT 6.520 18.530 6.850 18.700 ;
        RECT 1.600 17.310 1.790 17.330 ;
        RECT 3.350 17.310 3.540 17.330 ;
        RECT 1.460 17.220 1.790 17.310 ;
        RECT 1.460 17.140 1.540 17.220 ;
        RECT 1.600 17.100 1.790 17.220 ;
        RECT 3.210 17.220 3.540 17.310 ;
        RECT 3.210 17.140 3.290 17.220 ;
        RECT 3.350 17.100 3.540 17.220 ;
        RECT 0.410 16.000 0.590 17.060 ;
        RECT 1.060 16.690 1.230 17.020 ;
        RECT 1.140 16.620 1.190 16.690 ;
        RECT 1.140 16.590 1.480 16.620 ;
        RECT 1.020 16.580 1.480 16.590 ;
        RECT 1.020 16.460 1.490 16.580 ;
        RECT 1.160 16.390 1.490 16.460 ;
        RECT 1.160 16.360 1.480 16.390 ;
        RECT 2.160 16.000 2.340 17.060 ;
        RECT 2.810 16.690 2.980 17.020 ;
        RECT 2.890 16.620 2.940 16.690 ;
        RECT 2.890 16.590 3.230 16.620 ;
        RECT 2.770 16.580 3.230 16.590 ;
        RECT 2.770 16.460 3.240 16.580 ;
        RECT 2.910 16.390 3.240 16.460 ;
        RECT 11.040 16.540 11.370 16.710 ;
        RECT 11.480 16.630 11.810 16.800 ;
        RECT 2.910 16.360 3.230 16.390 ;
        RECT 11.040 16.260 11.400 16.540 ;
        RECT 8.970 16.010 9.290 16.050 ;
        RECT 8.970 15.820 9.300 16.010 ;
        RECT 8.970 15.790 9.290 15.820 ;
        RECT 9.370 15.800 9.570 16.130 ;
        RECT 9.960 15.940 10.160 16.130 ;
        RECT 10.690 16.090 11.400 16.260 ;
        RECT 10.630 15.970 10.950 16.010 ;
        RECT 9.650 15.610 9.840 15.620 ;
        RECT 9.850 15.610 10.200 15.940 ;
        RECT 10.630 15.780 10.960 15.970 ;
        RECT 10.630 15.750 10.950 15.780 ;
        RECT 0.430 15.300 0.750 15.340 ;
        RECT 2.180 15.300 2.500 15.340 ;
        RECT 0.430 15.110 0.760 15.300 ;
        RECT 2.180 15.110 2.510 15.300 ;
        RECT 0.430 15.080 0.750 15.110 ;
        RECT 2.180 15.080 2.500 15.110 ;
        RECT 8.740 15.100 8.910 15.430 ;
        RECT 8.920 15.360 9.240 15.400 ;
        RECT 8.920 15.170 9.250 15.360 ;
        RECT 8.920 15.140 9.240 15.170 ;
        RECT 9.370 15.140 9.570 15.470 ;
        RECT 9.650 15.280 10.200 15.610 ;
        RECT 1.800 14.920 2.120 14.960 ;
        RECT 9.850 14.950 10.200 15.280 ;
        RECT 1.800 14.730 2.130 14.920 ;
        RECT 10.690 14.770 11.390 15.650 ;
        RECT 1.800 14.700 2.120 14.730 ;
        RECT 1.570 14.550 1.910 14.560 ;
        RECT 1.320 14.510 1.910 14.550 ;
        RECT 1.240 14.480 1.910 14.510 ;
        RECT 2.990 14.480 3.310 14.510 ;
        RECT 1.230 14.360 1.910 14.480 ;
        RECT 1.150 14.140 1.910 14.360 ;
        RECT 2.980 14.290 3.310 14.480 ;
        RECT 10.030 14.380 10.220 14.610 ;
        RECT 2.990 14.250 3.310 14.290 ;
        RECT 1.150 13.990 1.740 14.140 ;
        RECT 1.080 13.970 1.740 13.990 ;
        RECT 1.080 13.820 1.910 13.970 ;
        RECT 1.080 13.680 1.320 13.820 ;
        RECT 1.740 13.800 1.910 13.820 ;
        RECT 2.830 13.680 3.000 13.990 ;
        RECT 8.740 13.840 8.910 14.170 ;
        RECT 8.920 14.100 9.240 14.130 ;
        RECT 8.920 13.910 9.250 14.100 ;
        RECT 8.920 13.870 9.240 13.910 ;
        RECT 9.370 13.800 9.570 14.130 ;
        RECT 9.850 13.990 10.200 14.320 ;
        RECT 10.680 14.170 11.380 14.350 ;
        RECT 1.080 13.660 1.410 13.680 ;
        RECT 1.090 13.650 1.410 13.660 ;
        RECT 1.080 13.460 1.410 13.650 ;
        RECT 1.090 13.420 1.410 13.460 ;
        RECT 2.640 13.420 3.160 13.680 ;
        RECT 1.150 12.490 1.320 13.420 ;
        RECT 8.550 13.190 8.800 13.730 ;
        RECT 9.650 13.660 10.200 13.990 ;
        RECT 9.650 13.650 9.840 13.660 ;
        RECT 8.970 13.450 9.290 13.480 ;
        RECT 8.970 13.260 9.300 13.450 ;
        RECT 8.970 13.220 9.290 13.260 ;
        RECT 8.550 12.840 8.760 13.190 ;
        RECT 9.370 13.140 9.570 13.470 ;
        RECT 9.850 13.330 10.200 13.660 ;
        RECT 10.680 13.750 11.000 13.790 ;
        RECT 10.680 13.560 11.010 13.750 ;
        RECT 10.680 13.530 11.000 13.560 ;
        RECT 9.960 13.140 10.160 13.330 ;
        RECT 8.970 13.010 9.290 13.050 ;
        RECT 8.970 12.820 9.300 13.010 ;
        RECT 8.970 12.790 9.290 12.820 ;
        RECT 9.370 12.800 9.570 13.130 ;
        RECT 9.960 12.940 10.160 13.130 ;
        RECT 10.670 13.030 10.990 13.070 ;
        RECT 9.650 12.610 9.840 12.620 ;
        RECT 9.850 12.610 10.200 12.940 ;
        RECT 10.670 12.840 11.000 13.030 ;
        RECT 10.670 12.810 10.990 12.840 ;
        RECT 8.740 12.100 8.910 12.430 ;
        RECT 8.920 12.360 9.240 12.400 ;
        RECT 8.920 12.170 9.250 12.360 ;
        RECT 8.920 12.140 9.240 12.170 ;
        RECT 9.370 12.140 9.570 12.470 ;
        RECT 9.650 12.280 10.200 12.610 ;
        RECT 9.850 12.020 10.200 12.280 ;
        RECT 9.850 11.950 10.220 12.020 ;
        RECT 10.030 11.790 10.220 11.950 ;
        RECT 10.680 11.890 11.380 12.070 ;
        RECT 1.160 9.550 1.330 11.330 ;
        RECT 8.740 10.840 8.910 11.170 ;
        RECT 8.920 11.100 9.240 11.130 ;
        RECT 8.920 10.910 9.250 11.100 ;
        RECT 8.920 10.870 9.240 10.910 ;
        RECT 9.370 10.800 9.570 11.130 ;
        RECT 9.850 10.990 10.200 11.320 ;
        RECT 9.650 10.660 10.200 10.990 ;
        RECT 10.690 10.820 11.390 11.470 ;
        RECT 9.650 10.650 9.840 10.660 ;
        RECT 4.400 10.550 4.720 10.590 ;
        RECT 4.390 10.360 4.720 10.550 ;
        RECT 4.400 10.350 4.720 10.360 ;
        RECT 4.390 10.330 4.720 10.350 ;
        RECT 8.970 10.450 9.290 10.480 ;
        RECT 4.390 10.020 4.560 10.330 ;
        RECT 8.970 10.260 9.300 10.450 ;
        RECT 8.970 10.220 9.290 10.260 ;
        RECT 9.370 10.140 9.570 10.470 ;
        RECT 9.850 10.330 10.200 10.660 ;
        RECT 10.590 10.590 11.390 10.820 ;
        RECT 10.590 10.560 10.910 10.590 ;
        RECT 9.960 10.140 10.160 10.330 ;
        RECT 10.690 9.980 11.400 10.150 ;
        RECT 4.550 9.720 4.870 9.760 ;
        RECT 4.540 9.530 4.870 9.720 ;
        RECT 11.040 9.700 11.400 9.980 ;
        RECT 11.040 9.530 11.370 9.700 ;
        RECT 4.550 9.500 4.870 9.530 ;
        RECT 11.480 9.440 11.810 9.610 ;
        RECT 3.740 8.900 4.060 8.930 ;
        RECT 3.740 8.710 4.070 8.900 ;
        RECT 3.740 8.670 4.060 8.710 ;
        RECT 3.720 6.950 3.900 8.010 ;
        RECT 4.470 7.620 4.790 7.650 ;
        RECT 4.470 7.550 4.800 7.620 ;
        RECT 4.330 7.430 4.800 7.550 ;
        RECT 4.330 7.420 4.790 7.430 ;
        RECT 4.450 7.390 4.790 7.420 ;
        RECT 4.450 7.320 4.500 7.390 ;
        RECT 4.370 6.990 4.540 7.320 ;
        RECT 4.770 6.790 4.850 6.870 ;
        RECT 4.910 6.790 5.100 6.910 ;
        RECT 4.770 6.700 5.100 6.790 ;
        RECT 4.910 6.680 5.100 6.700 ;
        RECT 7.350 3.520 7.530 5.570 ;
        RECT 8.080 5.310 8.410 5.480 ;
        RECT 8.160 3.530 8.330 5.310 ;
        RECT 7.350 0.470 7.530 2.520 ;
        RECT 8.080 2.260 8.410 2.430 ;
        RECT 8.160 0.480 8.330 2.260 ;
      LAYER mcon ;
        RECT 1.610 17.130 1.780 17.300 ;
        RECT 3.360 17.130 3.530 17.300 ;
        RECT 1.220 16.400 1.390 16.570 ;
        RECT 2.970 16.400 3.140 16.570 ;
        RECT 9.030 15.830 9.200 16.000 ;
        RECT 10.690 15.790 10.860 15.960 ;
        RECT 0.490 15.120 0.660 15.290 ;
        RECT 2.240 15.120 2.410 15.290 ;
        RECT 8.980 15.180 9.150 15.350 ;
        RECT 9.970 15.440 10.140 15.610 ;
        RECT 1.860 14.740 2.030 14.910 ;
        RECT 1.150 14.190 1.320 14.360 ;
        RECT 1.330 14.300 1.500 14.470 ;
        RECT 1.740 14.140 1.910 14.310 ;
        RECT 3.080 14.300 3.250 14.470 ;
        RECT 10.040 14.410 10.210 14.580 ;
        RECT 1.150 13.850 1.320 14.020 ;
        RECT 8.980 13.920 9.150 14.090 ;
        RECT 1.150 13.640 1.320 13.680 ;
        RECT 1.150 13.510 1.350 13.640 ;
        RECT 1.180 13.470 1.350 13.510 ;
        RECT 2.700 13.460 2.870 13.630 ;
        RECT 2.930 13.470 3.100 13.640 ;
        RECT 8.570 13.560 8.740 13.730 ;
        RECT 9.970 13.660 10.140 13.830 ;
        RECT 1.150 13.170 1.320 13.340 ;
        RECT 1.150 12.830 1.320 13.000 ;
        RECT 9.030 13.270 9.200 13.440 ;
        RECT 10.740 13.570 10.910 13.740 ;
        RECT 8.570 12.860 8.740 13.030 ;
        RECT 9.030 12.830 9.200 13.000 ;
        RECT 10.730 12.850 10.900 13.020 ;
        RECT 8.980 12.180 9.150 12.350 ;
        RECT 9.970 12.440 10.140 12.610 ;
        RECT 10.040 11.820 10.210 11.990 ;
        RECT 1.160 11.160 1.330 11.330 ;
        RECT 1.160 10.820 1.330 10.990 ;
        RECT 8.980 10.920 9.150 11.090 ;
        RECT 9.970 10.660 10.140 10.830 ;
        RECT 1.160 10.480 1.330 10.650 ;
        RECT 4.490 10.370 4.660 10.540 ;
        RECT 1.160 10.140 1.330 10.310 ;
        RECT 9.030 10.270 9.200 10.440 ;
        RECT 10.650 10.600 10.820 10.770 ;
        RECT 1.160 9.800 1.330 9.970 ;
        RECT 4.640 9.540 4.810 9.710 ;
        RECT 3.800 8.720 3.970 8.890 ;
        RECT 4.530 7.440 4.700 7.610 ;
        RECT 4.920 6.710 5.090 6.880 ;
      LAYER met1 ;
        RECT 1.580 17.070 1.810 17.360 ;
        RECT 3.330 17.070 3.560 17.360 ;
        RECT 1.150 16.330 1.470 16.650 ;
        RECT 1.500 15.800 1.710 17.040 ;
        RECT 2.900 16.330 3.220 16.650 ;
        RECT 3.250 15.800 3.460 17.040 ;
        RECT 8.960 16.000 9.280 16.080 ;
        RECT 1.500 15.480 1.830 15.800 ;
        RECT 3.250 15.480 3.580 15.800 ;
        RECT 8.960 15.760 9.530 16.000 ;
        RECT 0.420 15.050 0.740 15.370 ;
        RECT 1.500 15.270 1.710 15.480 ;
        RECT 2.170 15.050 2.490 15.370 ;
        RECT 3.250 15.270 3.460 15.480 ;
        RECT 9.190 15.430 9.530 15.760 ;
        RECT 8.910 15.110 9.530 15.430 ;
        RECT 1.790 14.670 2.110 14.990 ;
        RECT 1.120 14.560 1.650 14.570 ;
        RECT 1.120 14.550 1.910 14.560 ;
        RECT 1.120 14.250 1.940 14.550 ;
        RECT 1.120 13.960 1.970 14.250 ;
        RECT 3.000 14.220 3.320 14.540 ;
        RECT 9.190 14.160 9.530 15.110 ;
        RECT 1.120 13.710 1.940 13.960 ;
        RECT 8.910 13.840 9.530 14.160 ;
        RECT 1.100 13.390 1.760 13.710 ;
        RECT 2.630 13.390 3.170 13.710 ;
        RECT 1.120 9.530 1.760 13.390 ;
        RECT 8.520 12.850 8.840 13.770 ;
        RECT 9.190 13.510 9.530 13.840 ;
        RECT 8.960 13.190 9.530 13.510 ;
        RECT 9.190 13.080 9.530 13.190 ;
        RECT 8.550 12.840 8.840 12.850 ;
        RECT 8.960 12.760 9.530 13.080 ;
        RECT 9.190 12.430 9.530 12.760 ;
        RECT 8.910 12.110 9.530 12.430 ;
        RECT 9.190 11.160 9.530 12.110 ;
        RECT 8.910 10.840 9.530 11.160 ;
        RECT 4.410 10.300 4.730 10.620 ;
        RECT 9.190 10.510 9.530 10.840 ;
        RECT 8.960 10.280 9.530 10.510 ;
        RECT 9.860 15.670 10.130 15.990 ;
        RECT 10.620 15.720 10.940 16.040 ;
        RECT 9.860 15.380 10.170 15.670 ;
        RECT 9.860 14.640 10.130 15.380 ;
        RECT 9.860 14.350 10.240 14.640 ;
        RECT 9.860 13.890 10.130 14.350 ;
        RECT 9.860 13.600 10.170 13.890 ;
        RECT 9.860 12.670 10.130 13.600 ;
        RECT 10.670 13.500 10.990 13.820 ;
        RECT 10.660 12.780 10.980 13.100 ;
        RECT 9.860 12.380 10.170 12.670 ;
        RECT 9.860 12.050 10.130 12.380 ;
        RECT 9.860 11.760 10.240 12.050 ;
        RECT 9.860 10.890 10.130 11.760 ;
        RECT 9.860 10.600 10.170 10.890 ;
        RECT 9.860 10.290 10.130 10.600 ;
        RECT 10.580 10.530 10.900 10.850 ;
        RECT 8.960 10.190 9.280 10.280 ;
        RECT 1.340 9.520 1.760 9.530 ;
        RECT 4.560 9.470 4.880 9.790 ;
        RECT 3.730 8.640 4.050 8.960 ;
        RECT 4.810 8.530 5.020 8.740 ;
        RECT 4.810 8.210 5.140 8.530 ;
        RECT 4.460 7.360 4.780 7.680 ;
        RECT 4.810 6.970 5.020 8.210 ;
        RECT 4.890 6.650 5.120 6.940 ;
      LAYER via ;
        RECT 1.180 16.360 1.440 16.620 ;
        RECT 2.930 16.360 3.190 16.620 ;
        RECT 1.570 15.510 1.830 15.770 ;
        RECT 3.320 15.510 3.580 15.770 ;
        RECT 8.990 15.790 9.250 16.050 ;
        RECT 0.450 15.080 0.710 15.340 ;
        RECT 2.200 15.080 2.460 15.340 ;
        RECT 8.940 15.140 9.200 15.400 ;
        RECT 1.820 14.700 2.080 14.960 ;
        RECT 1.280 14.490 1.540 14.510 ;
        RECT 1.240 13.770 1.830 14.490 ;
        RECT 3.030 14.250 3.290 14.510 ;
        RECT 8.940 13.870 9.200 14.130 ;
        RECT 1.130 13.420 1.390 13.680 ;
        RECT 2.660 13.420 3.140 13.680 ;
        RECT 8.530 12.870 8.790 13.730 ;
        RECT 8.990 13.220 9.250 13.480 ;
        RECT 8.990 12.790 9.250 13.050 ;
        RECT 8.940 12.140 9.200 12.400 ;
        RECT 8.940 10.870 9.200 11.130 ;
        RECT 4.440 10.330 4.700 10.590 ;
        RECT 8.990 10.220 9.250 10.480 ;
        RECT 10.650 15.750 10.910 16.010 ;
        RECT 10.700 13.530 10.960 13.790 ;
        RECT 10.690 12.810 10.950 13.070 ;
        RECT 10.610 10.560 10.870 10.820 ;
        RECT 4.590 9.500 4.850 9.760 ;
        RECT 3.760 8.670 4.020 8.930 ;
        RECT 4.880 8.240 5.140 8.500 ;
        RECT 4.490 7.390 4.750 7.650 ;
      LAYER met2 ;
        RECT 1.150 16.460 1.460 16.660 ;
        RECT 2.900 16.460 3.210 16.660 ;
        RECT 0.920 16.230 1.790 16.460 ;
        RECT 2.670 16.230 3.540 16.460 ;
        RECT 0.920 16.220 1.350 16.230 ;
        RECT 2.670 16.220 3.100 16.230 ;
        RECT 1.540 15.680 1.860 15.770 ;
        RECT 3.290 15.680 3.610 15.770 ;
        RECT 1.400 15.430 1.870 15.680 ;
        RECT 3.150 15.430 3.620 15.680 ;
        RECT 0.420 15.050 0.730 15.380 ;
        RECT 2.170 15.050 2.480 15.380 ;
        RECT 8.470 15.000 8.800 15.210 ;
        RECT 2.430 13.540 3.310 13.790 ;
        RECT 6.350 13.780 6.600 14.150 ;
        RECT 8.470 14.060 8.800 14.270 ;
        RECT 2.630 13.510 3.170 13.540 ;
        RECT 2.630 13.390 4.970 13.510 ;
        RECT 2.780 13.290 4.970 13.390 ;
        RECT 6.380 12.930 6.590 13.220 ;
        RECT 8.470 12.000 8.800 12.210 ;
        RECT 8.470 11.060 8.800 11.270 ;
        RECT 4.820 10.850 6.590 11.050 ;
        RECT 3.250 10.500 3.410 10.680 ;
        RECT 3.230 10.490 3.410 10.500 ;
        RECT 3.010 10.360 3.410 10.490 ;
        RECT 4.420 10.470 4.730 10.630 ;
        RECT 3.010 9.870 3.370 10.360 ;
        RECT 3.990 10.250 4.870 10.470 ;
        RECT 3.990 10.220 6.590 10.250 ;
        RECT 4.530 10.040 6.590 10.220 ;
        RECT 4.570 9.610 4.880 9.800 ;
        RECT 4.530 9.360 5.080 9.610 ;
        RECT 3.730 8.630 4.040 8.960 ;
        RECT 4.710 8.330 5.180 8.580 ;
        RECT 4.850 8.240 5.170 8.330 ;
        RECT 4.230 7.780 4.660 7.790 ;
        RECT 4.230 7.550 5.100 7.780 ;
        RECT 4.460 7.350 4.770 7.550 ;
  END
END sky130_hilas_TA2SignalBiasCell

MACRO sky130_hilas_Tgate4Single01
  CLASS CORE ;
  FOREIGN sky130_hilas_Tgate4Single01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.390 BY 10.470 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPWR
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 0.740 2.260 0.940 2.300 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.740 8.270 0.940 8.310 ;
    END
  END VPWR
  PIN INPUT1_2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 5.390 0.050 5.590 ;
    END
  END INPUT1_2
  PIN SELECT2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 6.370 0.060 6.570 ;
    END
  END SELECT2
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 4.250 8.250 4.440 8.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.250 2.260 4.440 2.320 ;
    END
  END VGND
  PIN OUTPUT2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.690 6.370 4.760 6.570 ;
    END
  END OUTPUT2
  PIN OUTPUT4
    PORT
      LAYER met2 ;
        RECT 4.690 3.170 4.760 3.370 ;
    END
  END OUTPUT4
  PIN OUTPUT3
    PORT
      LAYER met2 ;
        RECT 4.690 3.900 4.760 4.100 ;
    END
  END OUTPUT3
  PIN OUTPUT1
    PORT
      LAYER met2 ;
        RECT 4.690 7.100 4.760 7.300 ;
    END
  END OUTPUT1
  PIN INPUT1_4
    PORT
      LAYER met2 ;
        RECT 0.000 2.190 0.050 2.390 ;
    END
  END INPUT1_4
  PIN SELECT4
    PORT
      LAYER met2 ;
        RECT 0.000 3.170 0.060 3.370 ;
    END
  END SELECT4
  PIN SELECT3
    PORT
      LAYER met2 ;
        RECT 0.000 3.900 0.060 4.100 ;
    END
  END SELECT3
  PIN INPUT1_3
    PORT
      LAYER met2 ;
        RECT 0.000 4.880 0.050 5.080 ;
    END
  END INPUT1_3
  PIN SELECT1
    PORT
      LAYER met2 ;
        RECT 0.000 7.100 0.060 7.300 ;
    END
  END SELECT1
  PIN INPUT1_1
    PORT
      LAYER met2 ;
        RECT 0.000 8.080 0.050 8.280 ;
    END
  END INPUT1_1
  OBS
      LAYER nwell ;
        RECT 5.040 9.790 6.180 10.380 ;
        RECT 4.550 8.950 6.180 9.790 ;
        RECT 2.750 7.930 5.510 8.700 ;
        RECT 0.120 7.520 0.130 7.900 ;
        RECT 2.750 7.760 4.740 7.930 ;
        RECT 2.750 7.140 4.730 7.760 ;
        RECT 5.040 7.140 6.180 7.180 ;
        RECT 2.750 7.090 6.180 7.140 ;
        RECT 5.040 6.590 6.180 7.090 ;
        RECT 4.550 6.580 6.180 6.590 ;
        RECT 2.750 5.750 6.180 6.580 ;
        RECT 2.750 5.740 4.740 5.750 ;
        RECT 2.750 4.730 5.510 5.740 ;
        RECT 2.750 4.720 4.740 4.730 ;
        RECT 2.750 3.890 6.180 4.720 ;
        RECT 4.550 3.880 6.180 3.890 ;
        RECT 5.040 3.380 6.180 3.880 ;
        RECT 2.750 3.330 6.180 3.380 ;
        RECT 2.750 2.710 4.730 3.330 ;
        RECT 5.040 3.290 6.180 3.330 ;
        RECT 2.750 2.540 4.740 2.710 ;
        RECT 2.750 1.770 5.510 2.540 ;
        RECT 4.550 0.680 6.180 1.520 ;
        RECT 5.040 0.090 6.180 0.680 ;
      LAYER li1 ;
        RECT 2.940 9.880 3.580 10.060 ;
        RECT 3.960 9.890 4.310 10.060 ;
        RECT 4.410 10.050 4.600 10.160 ;
        RECT 4.410 9.930 4.740 10.050 ;
        RECT 4.490 9.850 4.740 9.930 ;
        RECT 5.040 9.880 6.180 10.060 ;
        RECT 3.340 9.500 3.510 9.510 ;
        RECT 3.340 9.460 3.740 9.500 ;
        RECT 3.340 9.270 3.750 9.460 ;
        RECT 3.950 9.430 4.140 9.540 ;
        RECT 3.950 9.310 4.290 9.430 ;
        RECT 3.340 9.240 3.740 9.270 ;
        RECT 4.000 9.260 4.290 9.310 ;
        RECT 3.340 9.210 3.510 9.240 ;
        RECT 4.570 9.170 4.740 9.850 ;
        RECT 5.080 9.500 5.250 9.510 ;
        RECT 5.080 9.460 5.410 9.500 ;
        RECT 5.080 9.270 5.420 9.460 ;
        RECT 6.060 9.440 6.250 9.550 ;
        RECT 5.940 9.430 6.250 9.440 ;
        RECT 5.690 9.320 6.250 9.430 ;
        RECT 5.080 9.240 5.410 9.270 ;
        RECT 5.690 9.260 6.070 9.320 ;
        RECT 5.080 9.210 5.250 9.240 ;
        RECT 2.960 8.380 3.170 8.810 ;
        RECT 2.980 8.360 3.150 8.380 ;
        RECT 3.480 8.240 3.670 8.350 ;
        RECT 3.480 8.120 3.900 8.240 ;
        RECT 3.380 8.070 3.900 8.120 ;
        RECT 4.250 8.070 5.510 8.250 ;
        RECT 3.380 7.990 3.570 8.070 ;
        RECT 3.360 7.960 3.570 7.990 ;
        RECT 3.350 7.950 3.570 7.960 ;
        RECT 4.740 7.950 5.070 8.070 ;
        RECT 3.230 7.900 3.570 7.950 ;
        RECT 3.100 7.870 3.570 7.900 ;
        RECT 3.060 7.840 3.570 7.870 ;
        RECT 3.060 7.780 3.550 7.840 ;
        RECT 3.060 7.730 3.400 7.780 ;
        RECT 3.060 7.710 3.320 7.730 ;
        RECT 3.060 7.690 3.290 7.710 ;
        RECT 3.060 7.650 3.270 7.690 ;
        RECT 3.060 7.370 3.230 7.650 ;
        RECT 2.940 6.680 3.580 6.860 ;
        RECT 3.960 6.690 4.310 6.860 ;
        RECT 4.410 6.850 4.600 6.960 ;
        RECT 4.410 6.730 4.740 6.850 ;
        RECT 4.490 6.650 4.740 6.730 ;
        RECT 5.040 6.680 6.180 6.860 ;
        RECT 3.340 6.300 3.510 6.310 ;
        RECT 3.060 6.020 3.230 6.300 ;
        RECT 3.340 6.260 3.740 6.300 ;
        RECT 3.340 6.070 3.750 6.260 ;
        RECT 3.950 6.230 4.140 6.340 ;
        RECT 3.950 6.110 4.290 6.230 ;
        RECT 3.340 6.040 3.740 6.070 ;
        RECT 4.000 6.060 4.290 6.110 ;
        RECT 3.060 5.980 3.270 6.020 ;
        RECT 3.340 6.010 3.510 6.040 ;
        RECT 3.060 5.960 3.290 5.980 ;
        RECT 4.570 5.970 4.740 6.650 ;
        RECT 5.080 6.300 5.250 6.310 ;
        RECT 5.080 6.260 5.410 6.300 ;
        RECT 5.080 6.070 5.420 6.260 ;
        RECT 6.060 6.240 6.250 6.350 ;
        RECT 5.940 6.230 6.250 6.240 ;
        RECT 5.690 6.120 6.250 6.230 ;
        RECT 5.080 6.040 5.410 6.070 ;
        RECT 5.690 6.060 6.070 6.120 ;
        RECT 5.080 6.010 5.250 6.040 ;
        RECT 3.060 5.940 3.320 5.960 ;
        RECT 3.060 5.890 3.400 5.940 ;
        RECT 3.060 5.830 3.550 5.890 ;
        RECT 3.060 5.800 3.570 5.830 ;
        RECT 3.100 5.770 3.570 5.800 ;
        RECT 3.230 5.720 3.570 5.770 ;
        RECT 3.350 5.710 3.570 5.720 ;
        RECT 3.360 5.680 3.570 5.710 ;
        RECT 2.960 4.860 3.170 5.610 ;
        RECT 3.380 5.600 3.570 5.680 ;
        RECT 4.740 5.600 5.070 5.720 ;
        RECT 3.380 5.550 3.900 5.600 ;
        RECT 3.480 5.430 3.900 5.550 ;
        RECT 3.480 5.320 3.670 5.430 ;
        RECT 4.250 5.420 5.510 5.600 ;
        RECT 3.480 5.040 3.670 5.150 ;
        RECT 3.480 4.920 3.900 5.040 ;
        RECT 3.380 4.870 3.900 4.920 ;
        RECT 4.250 4.870 5.510 5.050 ;
        RECT 3.380 4.790 3.570 4.870 ;
        RECT 3.360 4.760 3.570 4.790 ;
        RECT 3.350 4.750 3.570 4.760 ;
        RECT 4.740 4.750 5.070 4.870 ;
        RECT 3.230 4.700 3.570 4.750 ;
        RECT 3.100 4.670 3.570 4.700 ;
        RECT 3.060 4.640 3.570 4.670 ;
        RECT 3.060 4.580 3.550 4.640 ;
        RECT 3.060 4.530 3.400 4.580 ;
        RECT 3.060 4.510 3.320 4.530 ;
        RECT 3.060 4.490 3.290 4.510 ;
        RECT 3.060 4.450 3.270 4.490 ;
        RECT 3.060 4.170 3.230 4.450 ;
        RECT 3.340 4.430 3.510 4.460 ;
        RECT 3.340 4.400 3.740 4.430 ;
        RECT 3.340 4.210 3.750 4.400 ;
        RECT 4.000 4.360 4.290 4.410 ;
        RECT 3.950 4.240 4.290 4.360 ;
        RECT 3.340 4.170 3.740 4.210 ;
        RECT 3.340 4.160 3.510 4.170 ;
        RECT 3.950 4.130 4.140 4.240 ;
        RECT 4.570 3.820 4.740 4.500 ;
        RECT 5.080 4.430 5.250 4.460 ;
        RECT 5.080 4.400 5.410 4.430 ;
        RECT 5.080 4.210 5.420 4.400 ;
        RECT 5.690 4.350 6.070 4.410 ;
        RECT 5.690 4.240 6.250 4.350 ;
        RECT 5.940 4.230 6.250 4.240 ;
        RECT 5.080 4.170 5.410 4.210 ;
        RECT 5.080 4.160 5.250 4.170 ;
        RECT 6.060 4.120 6.250 4.230 ;
        RECT 2.940 3.610 3.580 3.790 ;
        RECT 3.960 3.610 4.310 3.780 ;
        RECT 4.490 3.740 4.740 3.820 ;
        RECT 4.410 3.620 4.740 3.740 ;
        RECT 4.410 3.510 4.600 3.620 ;
        RECT 5.040 3.610 6.180 3.790 ;
        RECT 3.060 2.820 3.230 3.100 ;
        RECT 3.060 2.780 3.270 2.820 ;
        RECT 3.060 2.760 3.290 2.780 ;
        RECT 3.060 2.740 3.320 2.760 ;
        RECT 3.060 2.690 3.400 2.740 ;
        RECT 3.060 2.630 3.550 2.690 ;
        RECT 3.060 2.600 3.570 2.630 ;
        RECT 3.100 2.570 3.570 2.600 ;
        RECT 3.230 2.520 3.570 2.570 ;
        RECT 3.350 2.510 3.570 2.520 ;
        RECT 3.360 2.480 3.570 2.510 ;
        RECT 3.380 2.400 3.570 2.480 ;
        RECT 4.740 2.400 5.070 2.520 ;
        RECT 3.380 2.350 3.900 2.400 ;
        RECT 3.480 2.230 3.900 2.350 ;
        RECT 3.480 2.120 3.670 2.230 ;
        RECT 4.250 2.220 5.510 2.400 ;
        RECT 2.980 2.090 3.150 2.110 ;
        RECT 2.960 1.660 3.170 2.090 ;
        RECT 3.340 1.230 3.510 1.260 ;
        RECT 3.340 1.200 3.740 1.230 ;
        RECT 3.340 1.010 3.750 1.200 ;
        RECT 4.000 1.160 4.290 1.210 ;
        RECT 3.950 1.040 4.290 1.160 ;
        RECT 3.340 0.970 3.740 1.010 ;
        RECT 3.340 0.960 3.510 0.970 ;
        RECT 3.950 0.930 4.140 1.040 ;
        RECT 4.570 0.620 4.740 1.300 ;
        RECT 5.080 1.230 5.250 1.260 ;
        RECT 5.080 1.200 5.410 1.230 ;
        RECT 5.080 1.010 5.420 1.200 ;
        RECT 5.690 1.150 6.070 1.210 ;
        RECT 5.690 1.040 6.250 1.150 ;
        RECT 5.940 1.030 6.250 1.040 ;
        RECT 5.080 0.970 5.410 1.010 ;
        RECT 5.080 0.960 5.250 0.970 ;
        RECT 6.060 0.920 6.250 1.030 ;
        RECT 2.940 0.410 3.580 0.590 ;
        RECT 3.960 0.410 4.310 0.580 ;
        RECT 4.490 0.540 4.740 0.620 ;
        RECT 4.410 0.420 4.740 0.540 ;
        RECT 4.410 0.310 4.600 0.420 ;
        RECT 5.040 0.410 6.180 0.590 ;
      LAYER mcon ;
        RECT 4.420 9.960 4.590 10.130 ;
        RECT 3.480 9.280 3.650 9.450 ;
        RECT 3.960 9.340 4.130 9.510 ;
        RECT 5.150 9.280 5.320 9.450 ;
        RECT 6.070 9.350 6.240 9.520 ;
        RECT 3.490 8.150 3.660 8.320 ;
        RECT 4.420 6.760 4.590 6.930 ;
        RECT 3.480 6.080 3.650 6.250 ;
        RECT 3.960 6.140 4.130 6.310 ;
        RECT 5.150 6.080 5.320 6.250 ;
        RECT 6.070 6.150 6.240 6.320 ;
        RECT 2.980 5.140 3.150 5.330 ;
        RECT 3.490 5.350 3.660 5.520 ;
        RECT 3.490 4.950 3.660 5.120 ;
        RECT 3.480 4.220 3.650 4.390 ;
        RECT 3.960 4.160 4.130 4.330 ;
        RECT 5.150 4.220 5.320 4.390 ;
        RECT 6.070 4.150 6.240 4.320 ;
        RECT 4.420 3.540 4.590 3.710 ;
        RECT 3.490 2.150 3.660 2.320 ;
        RECT 2.980 1.940 3.150 2.110 ;
        RECT 3.480 1.020 3.650 1.190 ;
        RECT 3.960 0.960 4.130 1.130 ;
        RECT 5.150 1.020 5.320 1.190 ;
        RECT 6.070 0.950 6.240 1.120 ;
        RECT 4.420 0.340 4.590 0.510 ;
      LAYER met1 ;
        RECT 3.750 10.300 4.010 10.400 ;
        RECT 3.650 10.230 4.010 10.300 ;
        RECT 3.650 9.980 4.020 10.230 ;
        RECT 3.830 9.570 4.020 9.980 ;
        RECT 4.310 10.190 4.500 10.470 ;
        RECT 4.310 9.900 4.620 10.190 ;
        RECT 5.980 10.090 6.240 10.390 ;
        RECT 5.960 10.070 6.240 10.090 ;
        RECT 3.410 9.210 3.730 9.530 ;
        RECT 3.830 9.480 4.160 9.570 ;
        RECT 3.930 9.280 4.160 9.480 ;
        RECT 4.310 8.950 4.500 9.900 ;
        RECT 5.960 9.580 6.150 10.070 ;
        RECT 5.080 9.210 5.400 9.530 ;
        RECT 5.960 9.500 6.270 9.580 ;
        RECT 5.940 9.290 6.270 9.500 ;
        RECT 5.940 9.210 6.170 9.290 ;
        RECT 2.960 8.650 3.180 8.810 ;
        RECT 2.960 8.590 3.300 8.650 ;
        RECT 2.950 8.330 3.300 8.590 ;
        RECT 3.370 8.380 3.570 8.700 ;
        RECT 6.880 8.660 7.070 8.700 ;
        RECT 2.950 8.300 3.180 8.330 ;
        RECT 3.370 8.090 3.690 8.380 ;
        RECT 3.370 7.090 3.570 8.090 ;
        RECT 3.750 7.100 4.010 7.200 ;
        RECT 3.650 7.030 4.010 7.100 ;
        RECT 3.650 6.780 4.020 7.030 ;
        RECT 3.370 6.330 3.570 6.580 ;
        RECT 3.830 6.370 4.020 6.780 ;
        RECT 4.310 6.990 4.500 7.270 ;
        RECT 4.310 6.700 4.620 6.990 ;
        RECT 5.980 6.890 6.240 7.190 ;
        RECT 6.880 7.090 7.070 7.140 ;
        RECT 5.960 6.870 6.240 6.890 ;
        RECT 3.370 6.010 3.730 6.330 ;
        RECT 3.830 6.280 4.160 6.370 ;
        RECT 3.930 6.080 4.160 6.280 ;
        RECT 2.960 5.450 3.180 5.610 ;
        RECT 3.370 5.580 3.570 6.010 ;
        RECT 4.310 5.750 4.500 6.700 ;
        RECT 5.960 6.380 6.150 6.870 ;
        RECT 6.880 6.530 7.070 6.580 ;
        RECT 5.080 6.010 5.400 6.330 ;
        RECT 5.960 6.300 6.270 6.380 ;
        RECT 5.940 6.090 6.270 6.300 ;
        RECT 5.940 6.010 6.170 6.090 ;
        RECT 2.960 5.390 3.300 5.450 ;
        RECT 2.950 5.080 3.300 5.390 ;
        RECT 2.960 5.020 3.300 5.080 ;
        RECT 3.370 5.290 3.690 5.580 ;
        RECT 6.880 5.460 7.070 5.500 ;
        RECT 3.370 5.180 3.570 5.290 ;
        RECT 2.960 4.860 3.180 5.020 ;
        RECT 3.370 4.890 3.690 5.180 ;
        RECT 6.880 4.970 7.070 5.010 ;
        RECT 3.370 4.460 3.570 4.890 ;
        RECT 3.370 4.140 3.730 4.460 ;
        RECT 3.930 4.190 4.160 4.390 ;
        RECT 3.370 3.890 3.570 4.140 ;
        RECT 3.830 4.100 4.160 4.190 ;
        RECT 3.830 3.690 4.020 4.100 ;
        RECT 3.650 3.440 4.020 3.690 ;
        RECT 4.310 3.770 4.500 4.720 ;
        RECT 5.080 4.140 5.400 4.460 ;
        RECT 5.940 4.380 6.170 4.460 ;
        RECT 5.940 4.170 6.270 4.380 ;
        RECT 5.960 4.090 6.270 4.170 ;
        RECT 4.310 3.480 4.620 3.770 ;
        RECT 5.960 3.600 6.150 4.090 ;
        RECT 6.880 3.890 7.070 3.940 ;
        RECT 5.960 3.580 6.240 3.600 ;
        RECT 3.370 2.380 3.570 3.380 ;
        RECT 3.650 3.370 4.010 3.440 ;
        RECT 3.750 3.270 4.010 3.370 ;
        RECT 4.310 3.200 4.500 3.480 ;
        RECT 5.980 3.280 6.240 3.580 ;
        RECT 6.880 3.330 7.070 3.380 ;
        RECT 2.950 2.140 3.180 2.170 ;
        RECT 2.950 1.880 3.300 2.140 ;
        RECT 2.960 1.820 3.300 1.880 ;
        RECT 3.370 2.090 3.690 2.380 ;
        RECT 2.960 1.660 3.180 1.820 ;
        RECT 3.370 1.770 3.570 2.090 ;
        RECT 6.880 1.770 7.070 1.810 ;
        RECT 3.410 0.940 3.730 1.260 ;
        RECT 3.930 0.990 4.160 1.190 ;
        RECT 3.830 0.900 4.160 0.990 ;
        RECT 3.830 0.490 4.020 0.900 ;
        RECT 3.650 0.240 4.020 0.490 ;
        RECT 4.310 0.570 4.500 1.520 ;
        RECT 5.080 0.940 5.400 1.260 ;
        RECT 5.940 1.180 6.170 1.260 ;
        RECT 5.940 0.970 6.270 1.180 ;
        RECT 5.960 0.890 6.270 0.970 ;
        RECT 4.310 0.280 4.620 0.570 ;
        RECT 5.960 0.400 6.150 0.890 ;
        RECT 5.960 0.380 6.240 0.400 ;
        RECT 3.650 0.170 4.010 0.240 ;
        RECT 3.750 0.070 4.010 0.170 ;
        RECT 4.310 0.000 4.500 0.280 ;
        RECT 5.980 0.080 6.240 0.380 ;
      LAYER via ;
        RECT 3.750 10.110 4.010 10.370 ;
        RECT 5.980 10.100 6.240 10.360 ;
        RECT 3.440 9.240 3.700 9.500 ;
        RECT 5.110 9.240 5.370 9.500 ;
        RECT 3.040 8.360 3.300 8.620 ;
        RECT 3.750 6.910 4.010 7.170 ;
        RECT 5.980 6.900 6.240 7.160 ;
        RECT 3.440 6.040 3.700 6.300 ;
        RECT 5.110 6.040 5.370 6.300 ;
        RECT 3.040 5.050 3.300 5.420 ;
        RECT 3.440 4.170 3.700 4.430 ;
        RECT 3.750 3.300 4.010 3.560 ;
        RECT 5.110 4.170 5.370 4.430 ;
        RECT 5.980 3.310 6.240 3.570 ;
        RECT 3.040 1.850 3.300 2.110 ;
        RECT 3.440 0.970 3.700 1.230 ;
        RECT 3.750 0.100 4.010 0.360 ;
        RECT 5.110 0.970 5.370 1.230 ;
        RECT 5.980 0.110 6.240 0.370 ;
      LAYER met2 ;
        RECT 3.720 10.240 4.040 10.370 ;
        RECT 5.950 10.240 6.270 10.360 ;
        RECT 2.940 10.040 4.820 10.240 ;
        RECT 5.810 10.100 6.270 10.240 ;
        RECT 5.810 10.040 6.180 10.100 ;
        RECT 3.410 9.260 3.720 9.540 ;
        RECT 2.940 9.210 3.720 9.260 ;
        RECT 4.550 9.260 4.770 9.270 ;
        RECT 5.080 9.260 5.390 9.540 ;
        RECT 2.940 9.060 3.510 9.210 ;
        RECT 4.550 9.060 6.180 9.260 ;
        RECT 4.550 9.050 4.770 9.060 ;
        RECT 3.010 8.430 3.330 8.620 ;
        RECT 2.630 8.360 3.330 8.430 ;
        RECT 2.630 8.230 3.240 8.360 ;
        RECT 7.320 8.230 7.390 8.430 ;
        RECT 3.500 7.450 4.620 7.460 ;
        RECT 2.630 7.250 4.620 7.450 ;
        RECT 3.500 7.240 4.620 7.250 ;
        RECT 3.720 7.040 4.040 7.170 ;
        RECT 5.950 7.040 6.270 7.160 ;
        RECT 2.940 6.840 4.820 7.040 ;
        RECT 5.810 6.900 6.270 7.040 ;
        RECT 5.810 6.840 6.180 6.900 ;
        RECT 3.500 6.420 4.620 6.430 ;
        RECT 2.630 6.220 4.620 6.420 ;
        RECT 3.410 6.210 4.620 6.220 ;
        RECT 3.410 6.060 3.720 6.210 ;
        RECT 2.940 6.010 3.720 6.060 ;
        RECT 4.550 6.060 4.770 6.070 ;
        RECT 5.080 6.060 5.390 6.340 ;
        RECT 2.940 5.860 3.510 6.010 ;
        RECT 4.550 5.860 6.180 6.060 ;
        RECT 4.550 5.850 4.770 5.860 ;
        RECT 2.630 5.420 3.240 5.440 ;
        RECT 2.630 5.240 3.330 5.420 ;
        RECT 7.320 5.240 7.390 5.440 ;
        RECT 3.010 5.230 3.330 5.240 ;
        RECT 2.630 5.050 3.330 5.230 ;
        RECT 2.630 5.030 3.240 5.050 ;
        RECT 7.320 5.030 7.390 5.230 ;
        RECT 4.550 4.610 4.770 4.620 ;
        RECT 2.940 4.460 3.510 4.610 ;
        RECT 2.940 4.410 3.720 4.460 ;
        RECT 3.410 4.260 3.720 4.410 ;
        RECT 4.550 4.410 6.180 4.610 ;
        RECT 4.550 4.400 4.770 4.410 ;
        RECT 3.410 4.250 4.620 4.260 ;
        RECT 2.630 4.050 4.620 4.250 ;
        RECT 5.080 4.130 5.390 4.410 ;
        RECT 3.500 4.040 4.620 4.050 ;
        RECT 2.940 3.430 4.820 3.630 ;
        RECT 5.810 3.570 6.180 3.630 ;
        RECT 5.810 3.430 6.270 3.570 ;
        RECT 3.720 3.300 4.040 3.430 ;
        RECT 5.950 3.310 6.270 3.430 ;
        RECT 3.500 3.220 4.620 3.230 ;
        RECT 2.630 3.020 4.620 3.220 ;
        RECT 3.500 3.010 4.620 3.020 ;
        RECT 2.630 2.110 3.240 2.240 ;
        RECT 2.630 2.040 3.330 2.110 ;
        RECT 7.320 2.040 7.390 2.240 ;
        RECT 3.010 1.850 3.330 2.040 ;
        RECT 4.550 1.410 4.770 1.420 ;
        RECT 2.940 1.260 3.510 1.410 ;
        RECT 2.940 1.210 3.720 1.260 ;
        RECT 3.410 0.930 3.720 1.210 ;
        RECT 4.550 1.210 6.180 1.410 ;
        RECT 4.550 1.200 4.770 1.210 ;
        RECT 5.080 0.930 5.390 1.210 ;
        RECT 2.940 0.230 4.820 0.430 ;
        RECT 5.810 0.370 6.180 0.430 ;
        RECT 5.810 0.230 6.270 0.370 ;
        RECT 3.720 0.100 4.040 0.230 ;
        RECT 5.950 0.110 6.270 0.230 ;
  END
END sky130_hilas_Tgate4Single01

MACRO sky130_hilas_VinjDecode2to4
  CLASS CORE ;
  FOREIGN sky130_hilas_VinjDecode2to4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.320 BY 7.560 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN OUTPUT00
    PORT
      LAYER met2 ;
        RECT 12.820 6.270 12.950 6.440 ;
    END
  END OUTPUT00
  PIN OUTPUT01
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 12.940 5.010 13.310 5.090 ;
        RECT 12.940 5.000 13.970 5.010 ;
        RECT 15.850 5.000 16.160 5.160 ;
        RECT 12.940 4.930 16.320 5.000 ;
        RECT 12.820 4.830 16.320 4.930 ;
        RECT 12.820 4.760 12.950 4.830 ;
    END
  END OUTPUT01
  PIN OUTPUT10
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 12.940 3.500 13.310 3.580 ;
        RECT 12.940 3.490 13.970 3.500 ;
        RECT 15.850 3.490 16.160 3.650 ;
        RECT 12.940 3.420 16.320 3.490 ;
        RECT 12.820 3.320 16.320 3.420 ;
        RECT 12.820 3.250 12.950 3.320 ;
    END
  END OUTPUT10
  PIN OUTPUT11
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 12.940 1.990 13.310 2.070 ;
        RECT 12.940 1.980 13.970 1.990 ;
        RECT 15.850 1.980 16.160 2.140 ;
        RECT 12.940 1.920 16.320 1.980 ;
        RECT 12.820 1.810 16.320 1.920 ;
        RECT 12.820 1.750 12.950 1.810 ;
    END
  END OUTPUT11
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 11.660 7.510 11.930 7.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.660 1.540 11.930 1.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.180 7.470 3.410 7.560 ;
    END
  END VGND
  PIN VINJ
    ANTENNADIFFAREA 0.691200 ;
    PORT
      LAYER met1 ;
        RECT 6.540 1.590 6.770 6.120 ;
        RECT 6.690 1.540 6.910 1.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.690 7.490 6.910 7.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.610 7.480 0.830 7.560 ;
    END
  END VINJ
  PIN IN2
    PORT
      LAYER met2 ;
        RECT 0.000 5.480 0.110 5.660 ;
    END
  END IN2
  PIN IN1
    PORT
      LAYER met2 ;
        RECT 0.000 6.990 0.110 7.170 ;
    END
  END IN1
  PIN ENABLE
    PORT
      LAYER met2 ;
        RECT 0.000 3.970 0.110 4.150 ;
    END
  END ENABLE
  OBS
      LAYER nwell ;
        RECT 6.690 7.490 6.910 7.550 ;
        RECT 3.360 1.500 5.340 6.160 ;
        RECT 6.690 1.540 6.910 1.590 ;
        RECT 9.450 0.000 12.890 6.160 ;
      LAYER li1 ;
        RECT 3.980 5.730 4.150 5.870 ;
        RECT 10.070 5.730 10.240 5.870 ;
        RECT 10.800 5.750 10.970 5.830 ;
        RECT 11.610 5.750 11.780 5.830 ;
        RECT 13.150 5.790 13.320 5.910 ;
        RECT 3.980 5.560 4.170 5.730 ;
        RECT 3.980 5.460 4.150 5.560 ;
        RECT 3.550 5.080 3.720 5.180 ;
        RECT 3.530 4.910 3.720 5.080 ;
        RECT 3.550 4.850 3.720 4.910 ;
        RECT 3.970 5.120 4.140 5.180 ;
        RECT 3.970 4.850 4.220 5.120 ;
        RECT 4.710 5.100 4.960 5.180 ;
        RECT 4.710 4.930 6.010 5.100 ;
        RECT 6.570 5.090 6.740 5.720 ;
        RECT 10.070 5.560 10.260 5.730 ;
        RECT 10.070 5.460 10.240 5.560 ;
        RECT 10.800 5.180 11.010 5.750 ;
        RECT 11.570 5.500 11.780 5.750 ;
        RECT 12.170 5.570 12.340 5.670 ;
        RECT 13.110 5.620 13.320 5.790 ;
        RECT 15.040 5.720 15.300 5.790 ;
        RECT 15.840 5.720 16.020 5.850 ;
        RECT 13.150 5.580 13.320 5.620 ;
        RECT 11.570 5.180 11.740 5.500 ;
        RECT 12.140 5.400 12.340 5.570 ;
        RECT 12.170 5.300 12.340 5.400 ;
        RECT 13.710 5.540 14.580 5.710 ;
        RECT 15.040 5.540 16.020 5.720 ;
        RECT 3.980 4.830 4.220 4.850 ;
        RECT 4.790 4.840 4.960 4.930 ;
        RECT 6.490 4.920 6.820 5.090 ;
        RECT 9.640 5.080 9.810 5.180 ;
        RECT 9.620 4.910 9.810 5.080 ;
        RECT 9.640 4.850 9.810 4.910 ;
        RECT 10.060 5.120 10.230 5.180 ;
        RECT 10.060 4.850 10.310 5.120 ;
        RECT 10.800 4.930 11.050 5.180 ;
        RECT 10.070 4.830 10.310 4.850 ;
        RECT 10.880 4.840 11.050 4.930 ;
        RECT 11.530 4.930 11.740 5.180 ;
        RECT 13.710 5.100 13.880 5.540 ;
        RECT 15.040 5.100 15.300 5.540 ;
        RECT 15.840 5.430 16.020 5.540 ;
        RECT 12.250 4.930 13.880 5.100 ;
        RECT 14.330 4.930 15.300 5.100 ;
        RECT 15.750 4.930 16.090 5.100 ;
        RECT 11.530 4.850 11.700 4.930 ;
        RECT 13.020 4.890 13.190 4.930 ;
        RECT 3.980 4.220 4.150 4.360 ;
        RECT 10.070 4.220 10.240 4.360 ;
        RECT 10.800 4.240 10.970 4.320 ;
        RECT 11.610 4.240 11.780 4.320 ;
        RECT 13.150 4.280 13.320 4.400 ;
        RECT 3.980 4.050 4.170 4.220 ;
        RECT 3.980 3.950 4.150 4.050 ;
        RECT 3.550 3.570 3.720 3.670 ;
        RECT 3.530 3.400 3.720 3.570 ;
        RECT 3.550 3.340 3.720 3.400 ;
        RECT 3.970 3.610 4.140 3.670 ;
        RECT 3.970 3.340 4.220 3.610 ;
        RECT 4.710 3.590 4.960 3.670 ;
        RECT 4.710 3.420 6.010 3.590 ;
        RECT 6.570 3.580 6.740 4.210 ;
        RECT 10.070 4.050 10.260 4.220 ;
        RECT 10.070 3.950 10.240 4.050 ;
        RECT 10.800 3.670 11.010 4.240 ;
        RECT 11.570 3.990 11.780 4.240 ;
        RECT 12.170 4.060 12.340 4.160 ;
        RECT 13.110 4.110 13.320 4.280 ;
        RECT 15.040 4.210 15.300 4.280 ;
        RECT 15.840 4.210 16.020 4.340 ;
        RECT 13.150 4.070 13.320 4.110 ;
        RECT 11.570 3.670 11.740 3.990 ;
        RECT 12.140 3.890 12.340 4.060 ;
        RECT 12.170 3.790 12.340 3.890 ;
        RECT 13.710 4.030 14.580 4.200 ;
        RECT 15.040 4.030 16.020 4.210 ;
        RECT 3.980 3.320 4.220 3.340 ;
        RECT 4.790 3.330 4.960 3.420 ;
        RECT 6.490 3.410 6.820 3.580 ;
        RECT 9.640 3.570 9.810 3.670 ;
        RECT 9.620 3.400 9.810 3.570 ;
        RECT 9.640 3.340 9.810 3.400 ;
        RECT 10.060 3.610 10.230 3.670 ;
        RECT 10.060 3.340 10.310 3.610 ;
        RECT 10.800 3.420 11.050 3.670 ;
        RECT 10.070 3.320 10.310 3.340 ;
        RECT 10.880 3.330 11.050 3.420 ;
        RECT 11.530 3.420 11.740 3.670 ;
        RECT 13.710 3.590 13.880 4.030 ;
        RECT 15.040 3.590 15.300 4.030 ;
        RECT 15.840 3.920 16.020 4.030 ;
        RECT 12.250 3.420 13.880 3.590 ;
        RECT 14.330 3.420 15.300 3.590 ;
        RECT 15.750 3.420 16.090 3.590 ;
        RECT 11.530 3.340 11.700 3.420 ;
        RECT 13.020 3.380 13.190 3.420 ;
        RECT 3.980 2.710 4.150 2.850 ;
        RECT 10.070 2.710 10.240 2.850 ;
        RECT 10.800 2.730 10.970 2.810 ;
        RECT 11.610 2.730 11.780 2.810 ;
        RECT 13.150 2.770 13.320 2.890 ;
        RECT 3.980 2.540 4.170 2.710 ;
        RECT 3.980 2.440 4.150 2.540 ;
        RECT 3.550 2.060 3.720 2.160 ;
        RECT 3.530 1.890 3.720 2.060 ;
        RECT 3.550 1.830 3.720 1.890 ;
        RECT 3.970 2.100 4.140 2.160 ;
        RECT 3.970 1.830 4.220 2.100 ;
        RECT 4.710 2.080 4.960 2.160 ;
        RECT 4.710 1.910 6.010 2.080 ;
        RECT 6.570 2.070 6.740 2.700 ;
        RECT 10.070 2.540 10.260 2.710 ;
        RECT 10.070 2.440 10.240 2.540 ;
        RECT 10.800 2.160 11.010 2.730 ;
        RECT 11.570 2.480 11.780 2.730 ;
        RECT 12.170 2.550 12.340 2.650 ;
        RECT 13.110 2.600 13.320 2.770 ;
        RECT 15.040 2.700 15.300 2.770 ;
        RECT 15.840 2.700 16.020 2.830 ;
        RECT 13.150 2.560 13.320 2.600 ;
        RECT 11.570 2.160 11.740 2.480 ;
        RECT 12.140 2.380 12.340 2.550 ;
        RECT 12.170 2.280 12.340 2.380 ;
        RECT 13.710 2.520 14.580 2.690 ;
        RECT 15.040 2.520 16.020 2.700 ;
        RECT 3.980 1.810 4.220 1.830 ;
        RECT 4.790 1.820 4.960 1.910 ;
        RECT 6.490 1.900 6.820 2.070 ;
        RECT 9.640 2.060 9.810 2.160 ;
        RECT 9.620 1.890 9.810 2.060 ;
        RECT 9.640 1.830 9.810 1.890 ;
        RECT 10.060 2.100 10.230 2.160 ;
        RECT 10.060 1.830 10.310 2.100 ;
        RECT 10.800 1.910 11.050 2.160 ;
        RECT 10.070 1.810 10.310 1.830 ;
        RECT 10.880 1.820 11.050 1.910 ;
        RECT 11.530 1.910 11.740 2.160 ;
        RECT 13.710 2.080 13.880 2.520 ;
        RECT 15.040 2.080 15.300 2.520 ;
        RECT 15.840 2.410 16.020 2.520 ;
        RECT 12.250 1.910 13.880 2.080 ;
        RECT 14.330 1.910 15.300 2.080 ;
        RECT 15.750 1.910 16.090 2.080 ;
        RECT 11.530 1.830 11.700 1.910 ;
        RECT 13.020 1.870 13.190 1.910 ;
        RECT 10.070 1.210 10.240 1.350 ;
        RECT 10.800 1.230 10.970 1.310 ;
        RECT 11.610 1.230 11.780 1.310 ;
        RECT 13.150 1.270 13.320 1.390 ;
        RECT 10.070 1.040 10.260 1.210 ;
        RECT 10.070 0.940 10.240 1.040 ;
        RECT 10.800 0.660 11.010 1.230 ;
        RECT 11.570 0.980 11.780 1.230 ;
        RECT 12.170 1.050 12.340 1.150 ;
        RECT 13.110 1.100 13.320 1.270 ;
        RECT 15.040 1.200 15.300 1.270 ;
        RECT 15.840 1.200 16.020 1.330 ;
        RECT 13.150 1.060 13.320 1.100 ;
        RECT 11.570 0.660 11.740 0.980 ;
        RECT 12.140 0.880 12.340 1.050 ;
        RECT 12.170 0.780 12.340 0.880 ;
        RECT 13.710 1.020 14.580 1.190 ;
        RECT 15.040 1.020 16.020 1.200 ;
        RECT 9.640 0.560 9.810 0.660 ;
        RECT 9.620 0.390 9.810 0.560 ;
        RECT 9.640 0.330 9.810 0.390 ;
        RECT 10.060 0.600 10.230 0.660 ;
        RECT 10.060 0.330 10.310 0.600 ;
        RECT 10.800 0.410 11.050 0.660 ;
        RECT 10.070 0.310 10.310 0.330 ;
        RECT 10.880 0.320 11.050 0.410 ;
        RECT 11.530 0.410 11.740 0.660 ;
        RECT 13.710 0.580 13.880 1.020 ;
        RECT 15.040 0.580 15.300 1.020 ;
        RECT 15.840 0.910 16.020 1.020 ;
        RECT 12.250 0.410 13.880 0.580 ;
        RECT 14.330 0.410 15.300 0.580 ;
        RECT 15.750 0.410 16.090 0.580 ;
        RECT 11.530 0.330 11.700 0.410 ;
        RECT 13.020 0.370 13.190 0.410 ;
      LAYER mcon ;
        RECT 4.000 5.560 4.170 5.730 ;
        RECT 10.090 5.560 10.260 5.730 ;
        RECT 6.570 5.200 6.740 5.370 ;
        RECT 4.010 4.880 4.180 5.050 ;
        RECT 5.350 4.930 5.520 5.100 ;
        RECT 10.100 4.880 10.270 5.050 ;
        RECT 15.070 5.220 15.250 5.400 ;
        RECT 4.000 4.050 4.170 4.220 ;
        RECT 10.090 4.050 10.260 4.220 ;
        RECT 6.570 3.690 6.740 3.860 ;
        RECT 4.010 3.370 4.180 3.540 ;
        RECT 5.350 3.420 5.520 3.590 ;
        RECT 10.100 3.370 10.270 3.540 ;
        RECT 15.070 3.710 15.250 3.890 ;
        RECT 4.000 2.540 4.170 2.710 ;
        RECT 10.090 2.540 10.260 2.710 ;
        RECT 6.570 2.180 6.740 2.350 ;
        RECT 4.010 1.860 4.180 2.030 ;
        RECT 5.350 1.910 5.520 2.080 ;
        RECT 10.100 1.860 10.270 2.030 ;
        RECT 15.070 2.200 15.250 2.380 ;
        RECT 10.090 1.040 10.260 1.210 ;
        RECT 10.100 0.360 10.270 0.530 ;
        RECT 15.070 0.700 15.250 0.880 ;
      LAYER met1 ;
        RECT 3.670 7.210 3.940 7.500 ;
        RECT 3.630 6.940 3.960 7.210 ;
        RECT 3.670 6.160 3.940 6.940 ;
        RECT 3.660 5.830 3.940 6.160 ;
        RECT 4.130 6.120 4.400 6.600 ;
        RECT 3.670 5.800 3.940 5.830 ;
        RECT 3.440 4.840 3.750 5.190 ;
        RECT 3.440 3.330 3.750 3.680 ;
        RECT 3.970 2.980 4.400 6.120 ;
        RECT 4.590 5.610 4.860 7.070 ;
        RECT 5.540 6.570 5.830 6.620 ;
        RECT 5.520 6.220 5.830 6.570 ;
        RECT 4.540 5.340 4.870 5.610 ;
        RECT 4.590 4.030 4.860 5.340 ;
        RECT 5.540 5.140 5.830 6.220 ;
        RECT 10.060 5.780 10.280 6.120 ;
        RECT 10.060 5.520 10.290 5.780 ;
        RECT 5.270 5.130 5.830 5.140 ;
        RECT 4.570 3.700 4.860 4.030 ;
        RECT 4.590 3.680 4.860 3.700 ;
        RECT 5.060 4.880 5.830 5.130 ;
        RECT 5.060 4.740 5.340 4.880 ;
        RECT 5.060 3.630 5.330 4.740 ;
        RECT 5.540 3.630 5.830 4.880 ;
        RECT 9.530 4.840 9.840 5.190 ;
        RECT 10.060 5.120 10.280 5.520 ;
        RECT 12.080 5.360 12.410 5.620 ;
        RECT 13.050 5.580 13.480 5.870 ;
        RECT 10.060 4.810 10.310 5.120 ;
        RECT 12.920 4.830 13.310 5.100 ;
        RECT 10.060 4.270 10.280 4.810 ;
        RECT 10.060 4.010 10.290 4.270 ;
        RECT 5.060 3.570 5.830 3.630 ;
        RECT 5.060 3.370 5.840 3.570 ;
        RECT 3.970 2.650 4.430 2.980 ;
        RECT 3.970 2.600 4.400 2.650 ;
        RECT 3.970 2.500 4.200 2.600 ;
        RECT 5.060 2.530 5.330 3.370 ;
        RECT 3.440 1.820 3.750 2.170 ;
        RECT 3.970 2.100 4.190 2.500 ;
        RECT 5.040 2.200 5.330 2.530 ;
        RECT 5.060 2.170 5.330 2.200 ;
        RECT 5.540 3.220 5.840 3.370 ;
        RECT 9.530 3.330 9.840 3.680 ;
        RECT 10.060 3.610 10.280 4.010 ;
        RECT 12.080 3.850 12.410 4.110 ;
        RECT 13.050 4.070 13.480 4.360 ;
        RECT 10.060 3.300 10.310 3.610 ;
        RECT 12.920 3.320 13.310 3.590 ;
        RECT 5.540 2.120 5.830 3.220 ;
        RECT 10.060 2.760 10.280 3.300 ;
        RECT 10.060 2.500 10.290 2.760 ;
        RECT 3.970 1.790 4.220 2.100 ;
        RECT 5.270 1.860 5.830 2.120 ;
        RECT 3.970 1.590 4.190 1.790 ;
        RECT 5.540 1.680 5.830 1.860 ;
        RECT 9.530 1.820 9.840 2.170 ;
        RECT 10.060 2.100 10.280 2.500 ;
        RECT 12.080 2.340 12.410 2.600 ;
        RECT 13.050 2.560 13.480 2.850 ;
        RECT 10.060 1.790 10.310 2.100 ;
        RECT 12.920 1.810 13.310 2.080 ;
        RECT 10.060 1.260 10.280 1.790 ;
        RECT 10.060 1.000 10.290 1.260 ;
        RECT 9.530 0.320 9.840 0.670 ;
        RECT 10.060 0.600 10.280 1.000 ;
        RECT 12.080 0.840 12.410 1.100 ;
        RECT 13.050 1.060 13.480 1.350 ;
        RECT 10.060 0.290 10.310 0.600 ;
        RECT 12.920 0.310 13.310 0.580 ;
        RECT 10.060 0.090 10.280 0.290 ;
        RECT 15.030 0.090 15.300 6.130 ;
        RECT 15.850 4.840 16.160 5.160 ;
        RECT 15.850 3.330 16.160 3.650 ;
        RECT 15.850 1.820 16.160 2.140 ;
        RECT 15.850 0.320 16.160 0.640 ;
      LAYER via ;
        RECT 3.660 6.940 3.930 7.210 ;
        RECT 4.590 6.750 4.860 7.020 ;
        RECT 3.660 5.860 3.930 6.130 ;
        RECT 4.130 6.260 4.400 6.530 ;
        RECT 3.470 4.870 3.730 5.130 ;
        RECT 5.520 6.250 5.810 6.540 ;
        RECT 4.570 5.340 4.840 5.610 ;
        RECT 4.120 4.180 4.390 4.450 ;
        RECT 3.470 3.360 3.730 3.620 ;
        RECT 4.570 3.730 4.840 4.000 ;
        RECT 5.300 5.040 5.560 5.140 ;
        RECT 5.070 5.000 5.560 5.040 ;
        RECT 5.070 4.880 5.820 5.000 ;
        RECT 5.070 4.770 5.340 4.880 ;
        RECT 5.560 4.740 5.820 4.880 ;
        RECT 9.560 4.870 9.820 5.130 ;
        RECT 12.120 5.360 12.380 5.620 ;
        RECT 13.110 5.610 13.370 5.870 ;
        RECT 12.980 4.830 13.240 5.090 ;
        RECT 5.300 3.540 5.560 3.630 ;
        RECT 5.300 3.370 5.840 3.540 ;
        RECT 4.160 2.680 4.430 2.950 ;
        RECT 3.470 1.850 3.730 2.110 ;
        RECT 5.040 2.230 5.310 2.500 ;
        RECT 5.550 3.250 5.840 3.370 ;
        RECT 9.560 3.360 9.820 3.620 ;
        RECT 12.120 3.850 12.380 4.110 ;
        RECT 13.110 4.100 13.370 4.360 ;
        RECT 12.980 3.320 13.240 3.580 ;
        RECT 5.300 2.000 5.560 2.120 ;
        RECT 5.300 1.860 5.830 2.000 ;
        RECT 5.540 1.710 5.830 1.860 ;
        RECT 9.560 1.850 9.820 2.110 ;
        RECT 12.120 2.340 12.380 2.600 ;
        RECT 13.110 2.590 13.370 2.850 ;
        RECT 12.980 1.810 13.240 2.070 ;
        RECT 9.560 0.350 9.820 0.610 ;
        RECT 12.120 0.840 12.380 1.100 ;
        RECT 13.110 1.090 13.370 1.350 ;
        RECT 12.980 0.310 13.240 0.570 ;
        RECT 15.880 4.870 16.140 5.130 ;
        RECT 15.880 3.360 16.140 3.620 ;
        RECT 15.880 1.850 16.140 2.110 ;
        RECT 15.880 0.350 16.140 0.610 ;
      LAYER met2 ;
        RECT 3.710 7.400 6.080 7.410 ;
        RECT 3.690 7.250 6.080 7.400 ;
        RECT 3.690 7.240 3.960 7.250 ;
        RECT 3.660 7.170 3.960 7.240 ;
        RECT 3.430 6.990 3.960 7.170 ;
        RECT 3.660 6.910 3.930 6.990 ;
        RECT 4.560 6.960 4.890 7.020 ;
        RECT 4.560 6.800 6.080 6.960 ;
        RECT 4.560 6.750 4.890 6.800 ;
        RECT 4.100 6.500 4.430 6.530 ;
        RECT 3.430 6.320 4.450 6.500 ;
        RECT 4.100 6.310 4.450 6.320 ;
        RECT 5.490 6.470 5.840 6.540 ;
        RECT 5.490 6.310 6.080 6.470 ;
        RECT 4.100 6.260 4.430 6.310 ;
        RECT 5.490 6.250 5.840 6.310 ;
        RECT 3.630 6.070 3.960 6.130 ;
        RECT 3.630 5.910 5.270 6.070 ;
        RECT 3.630 5.860 3.960 5.910 ;
        RECT 5.110 5.900 5.270 5.910 ;
        RECT 5.110 5.740 6.070 5.900 ;
        RECT 9.440 5.810 13.480 5.970 ;
        RECT 3.360 5.550 6.970 5.730 ;
        RECT 3.430 5.480 4.840 5.550 ;
        RECT 12.080 5.540 12.410 5.620 ;
        RECT 13.060 5.580 13.480 5.810 ;
        RECT 11.810 5.520 12.410 5.540 ;
        RECT 4.570 5.450 4.840 5.480 ;
        RECT 4.570 5.310 4.850 5.450 ;
        RECT 4.620 5.290 4.850 5.310 ;
        RECT 5.120 5.290 6.080 5.450 ;
        RECT 9.450 5.360 12.410 5.520 ;
        RECT 5.120 5.140 5.280 5.290 ;
        RECT 3.440 5.030 3.760 5.130 ;
        RECT 5.120 5.060 5.590 5.140 ;
        RECT 5.120 5.040 6.970 5.060 ;
        RECT 3.430 4.990 3.760 5.030 ;
        RECT 5.040 4.990 6.970 5.040 ;
        RECT 9.530 5.030 9.850 5.130 ;
        RECT 3.430 4.880 6.970 4.990 ;
        RECT 3.430 4.810 5.370 4.880 ;
        RECT 5.040 4.770 5.370 4.810 ;
        RECT 5.530 4.800 6.080 4.880 ;
        RECT 9.450 4.870 9.850 5.030 ;
        RECT 5.530 4.740 5.850 4.800 ;
        RECT 4.090 4.390 4.420 4.450 ;
        RECT 4.090 4.230 6.080 4.390 ;
        RECT 9.440 4.300 13.480 4.460 ;
        RECT 4.090 4.220 4.420 4.230 ;
        RECT 3.360 4.040 6.970 4.220 ;
        RECT 12.080 4.030 12.410 4.110 ;
        RECT 13.060 4.070 13.480 4.300 ;
        RECT 11.810 4.010 12.410 4.030 ;
        RECT 4.540 3.940 4.870 4.000 ;
        RECT 4.540 3.780 6.080 3.940 ;
        RECT 9.450 3.850 12.410 4.010 ;
        RECT 4.540 3.730 4.870 3.780 ;
        RECT 3.440 3.520 3.760 3.620 ;
        RECT 3.430 3.480 3.760 3.520 ;
        RECT 5.270 3.550 5.590 3.630 ;
        RECT 5.270 3.480 6.970 3.550 ;
        RECT 9.530 3.520 9.850 3.620 ;
        RECT 3.430 3.370 6.970 3.480 ;
        RECT 3.430 3.300 6.080 3.370 ;
        RECT 9.450 3.360 9.850 3.520 ;
        RECT 5.520 3.290 6.080 3.300 ;
        RECT 5.520 3.250 5.870 3.290 ;
        RECT 4.130 2.890 4.460 2.950 ;
        RECT 4.130 2.730 6.080 2.890 ;
        RECT 9.440 2.790 13.480 2.950 ;
        RECT 4.130 2.710 4.460 2.730 ;
        RECT 3.360 2.530 6.970 2.710 ;
        RECT 12.080 2.520 12.410 2.600 ;
        RECT 13.060 2.560 13.480 2.790 ;
        RECT 11.810 2.500 12.410 2.520 ;
        RECT 5.010 2.440 5.340 2.500 ;
        RECT 5.010 2.280 6.080 2.440 ;
        RECT 9.450 2.340 12.410 2.500 ;
        RECT 5.010 2.230 5.340 2.280 ;
        RECT 3.440 2.010 3.760 2.110 ;
        RECT 3.430 1.850 3.760 2.010 ;
        RECT 5.270 2.040 5.590 2.120 ;
        RECT 5.270 1.860 6.970 2.040 ;
        RECT 9.530 2.010 9.850 2.110 ;
        RECT 5.510 1.790 6.080 1.860 ;
        RECT 9.450 1.850 9.850 2.010 ;
        RECT 5.510 1.710 5.860 1.790 ;
        RECT 9.440 1.290 13.480 1.450 ;
        RECT 12.080 1.020 12.410 1.100 ;
        RECT 13.060 1.060 13.480 1.290 ;
        RECT 11.810 1.000 12.410 1.020 ;
        RECT 9.450 0.840 12.410 1.000 ;
        RECT 9.530 0.510 9.850 0.610 ;
        RECT 9.450 0.350 9.850 0.510 ;
        RECT 12.940 0.490 13.310 0.570 ;
        RECT 12.940 0.480 13.970 0.490 ;
        RECT 15.850 0.480 16.160 0.640 ;
        RECT 12.940 0.310 16.320 0.480 ;
  END
END sky130_hilas_VinjDecode2to4

MACRO sky130_hilas_TA2Cell_1FG
  CLASS CORE ;
  FOREIGN sky130_hilas_TA2Cell_1FG ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.900 BY 23.320 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 17.820 10.230 18.300 10.240 ;
        RECT 17.820 9.990 18.710 10.230 ;
    END
  END VIN12
  PIN VIN11
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 17.870 13.750 18.710 13.950 ;
    END
  END VIN11
  PIN VIN21
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 32.610 12.090 32.930 12.330 ;
    END
  END VIN21
  PIN VIN22
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 32.530 14.760 32.840 15.000 ;
    END
  END VIN22
  PIN VPWR
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 35.760 14.880 36.040 15.030 ;
    END
    PORT
      LAYER met1 ;
        RECT 35.770 8.980 36.040 9.190 ;
    END
  END VPWR
  PIN VGND
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 35.530 16.460 35.850 16.540 ;
        RECT 34.540 16.280 35.850 16.460 ;
        RECT 34.540 16.110 35.720 16.280 ;
        RECT 34.590 15.960 34.910 16.110 ;
    END
    PORT
      LAYER met2 ;
        RECT 23.150 9.330 23.470 9.340 ;
        RECT 33.590 9.330 33.920 9.470 ;
        RECT 23.150 9.170 33.920 9.330 ;
        RECT 23.150 9.160 23.840 9.170 ;
        RECT 23.150 9.040 23.470 9.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.440 14.940 17.670 15.020 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.230 14.940 23.460 15.030 ;
    END
  END VGND
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 6.890 15.040 7.200 15.260 ;
        RECT 5.010 14.860 16.540 15.040 ;
        RECT 31.410 14.860 31.730 14.980 ;
        RECT 5.010 14.830 31.730 14.860 ;
        RECT 6.320 14.820 31.730 14.830 ;
        RECT 9.210 14.680 31.730 14.820 ;
        RECT 14.180 14.410 14.490 14.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.410 8.980 31.690 9.030 ;
    END
    PORT
      LAYER met1 ;
        RECT 9.210 14.980 9.490 15.030 ;
        RECT 9.210 14.700 9.530 14.980 ;
      LAYER via ;
        RECT 9.240 14.710 9.500 14.970 ;
    END
  END VINJ
  PIN OUTPUT1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 36.950 12.320 37.060 12.550 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 36.950 11.500 37.060 11.720 ;
    END
  END OUTPUT2
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 8.970 14.350 9.040 14.530 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 8.970 9.480 9.050 9.660 ;
    END
  END DRAIN2
  PIN COLSEL2
    PORT
      LAYER met1 ;
        RECT 9.740 14.970 9.930 15.030 ;
    END
  END COLSEL2
  PIN GATE2
    PORT
      LAYER met1 ;
        RECT 16.220 14.940 16.450 15.020 ;
    END
  END GATE2
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT 24.450 14.950 24.680 15.030 ;
    END
  END GATE1
  PIN COLSEL1
    PORT
      LAYER met1 ;
        RECT 30.970 14.950 31.160 15.030 ;
    END
    PORT
      LAYER met1 ;
        RECT 30.970 8.980 31.160 9.030 ;
    END
  END COLSEL1
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 19.730 14.870 21.170 15.030 ;
    END
  END VTUN
  OBS
      LAYER nwell ;
        RECT 0.290 22.980 2.020 23.320 ;
        RECT 38.880 22.980 40.610 23.320 ;
        RECT 0.290 21.420 2.040 22.980 ;
        RECT 0.310 19.790 2.040 21.420 ;
        RECT 38.860 21.420 40.610 22.980 ;
        RECT 38.860 19.790 40.590 21.420 ;
        RECT 0.250 19.400 3.560 19.790 ;
        RECT 0.010 19.360 3.560 19.400 ;
        RECT 0.000 17.710 3.560 19.360 ;
        RECT 37.340 19.400 40.650 19.790 ;
        RECT 37.340 19.360 40.890 19.400 ;
        RECT 32.580 19.310 35.890 19.320 ;
        RECT 34.930 19.280 35.120 19.310 ;
        RECT 0.250 16.620 3.560 17.710 ;
        RECT 37.340 17.710 40.900 19.360 ;
        RECT 0.250 14.780 3.560 15.970 ;
        RECT 8.970 15.020 10.950 15.030 ;
        RECT 0.000 13.130 3.560 14.780 ;
        RECT 15.390 14.670 15.950 17.090 ;
        RECT 24.950 14.670 25.510 17.090 ;
        RECT 37.340 16.620 40.650 17.710 ;
        RECT 37.760 15.970 39.040 16.620 ;
        RECT 31.930 15.020 33.400 15.030 ;
        RECT 35.780 14.850 37.060 15.030 ;
        RECT 37.340 14.780 40.650 15.970 ;
        RECT 8.970 14.350 9.040 14.530 ;
        RECT 0.010 13.090 3.560 13.130 ;
        RECT 0.250 12.800 3.560 13.090 ;
        RECT 37.340 13.130 40.900 14.780 ;
        RECT 37.340 13.090 40.890 13.130 ;
        RECT 37.340 12.800 40.650 13.090 ;
        RECT 8.970 9.480 9.050 9.660 ;
        RECT 37.760 9.470 39.040 12.310 ;
        RECT 35.780 8.980 37.060 9.170 ;
        RECT 31.930 7.550 32.380 7.780 ;
        RECT 30.590 7.420 32.450 7.490 ;
        RECT 34.220 3.050 36.080 6.040 ;
        RECT 34.220 0.000 36.080 2.990 ;
      LAYER li1 ;
        RECT 1.070 21.590 1.620 22.020 ;
        RECT 39.280 21.590 39.830 22.020 ;
        RECT 1.070 19.860 1.620 20.290 ;
        RECT 39.280 19.860 39.830 20.290 ;
        RECT 0.650 19.060 0.850 19.410 ;
        RECT 2.130 19.160 2.660 19.330 ;
        RECT 38.240 19.160 38.770 19.330 ;
        RECT 0.640 19.030 0.850 19.060 ;
        RECT 0.640 18.450 0.860 19.030 ;
        RECT 0.640 18.440 0.850 18.450 ;
        RECT 1.020 18.270 1.210 18.280 ;
        RECT 1.010 17.980 1.210 18.270 ;
        RECT 0.930 17.650 1.220 17.980 ;
        RECT 1.410 17.170 1.580 18.780 ;
        RECT 2.190 18.230 2.420 18.920 ;
        RECT 9.610 18.310 14.670 19.140 ;
        RECT 40.050 19.060 40.250 19.410 ;
        RECT 40.050 19.030 40.260 19.060 ;
        RECT 14.120 18.230 14.600 18.310 ;
        RECT 38.480 18.230 38.710 18.920 ;
        RECT 1.400 16.980 1.580 17.170 ;
        RECT 2.240 17.080 2.410 18.230 ;
        RECT 14.120 18.130 14.450 18.230 ;
        RECT 14.120 17.980 14.270 18.130 ;
        RECT 6.870 17.940 7.190 17.980 ;
        RECT 6.860 17.750 7.190 17.940 ;
        RECT 6.870 17.720 7.190 17.750 ;
        RECT 33.710 17.940 34.030 17.980 ;
        RECT 33.710 17.750 34.040 17.940 ;
        RECT 33.710 17.720 34.030 17.750 ;
        RECT 38.490 17.080 38.660 18.230 ;
        RECT 39.320 17.170 39.490 18.780 ;
        RECT 40.040 18.450 40.260 19.030 ;
        RECT 40.050 18.440 40.260 18.450 ;
        RECT 39.690 18.270 39.880 18.280 ;
        RECT 39.690 17.980 39.890 18.270 ;
        RECT 39.680 17.650 39.970 17.980 ;
        RECT 39.320 16.980 39.500 17.170 ;
        RECT 13.310 16.430 13.500 16.750 ;
        RECT 27.400 16.430 27.590 16.750 ;
        RECT 13.310 16.340 13.590 16.430 ;
        RECT 9.950 16.200 13.590 16.340 ;
        RECT 27.310 16.340 27.590 16.430 ;
        RECT 38.320 16.540 38.650 16.710 ;
        RECT 38.760 16.630 39.090 16.800 ;
        RECT 27.310 16.200 30.950 16.340 ;
        RECT 38.320 16.260 38.680 16.540 ;
        RECT 9.950 16.160 13.500 16.200 ;
        RECT 13.310 15.740 13.500 16.160 ;
        RECT 27.400 16.160 30.950 16.200 ;
        RECT 27.400 15.740 27.590 16.160 ;
        RECT 36.250 16.010 36.570 16.050 ;
        RECT 36.250 15.820 36.580 16.010 ;
        RECT 36.250 15.790 36.570 15.820 ;
        RECT 36.650 15.800 36.850 16.130 ;
        RECT 37.240 15.940 37.440 16.130 ;
        RECT 37.970 16.090 38.680 16.260 ;
        RECT 37.910 15.970 38.230 16.010 ;
        RECT 36.930 15.610 37.120 15.620 ;
        RECT 37.130 15.610 37.480 15.940 ;
        RECT 37.910 15.780 38.240 15.970 ;
        RECT 37.910 15.750 38.230 15.780 ;
        RECT 1.400 15.420 1.580 15.610 ;
        RECT 0.930 14.610 1.220 14.940 ;
        RECT 1.010 14.320 1.210 14.610 ;
        RECT 1.020 14.310 1.210 14.320 ;
        RECT 0.640 14.140 0.850 14.150 ;
        RECT 0.640 13.560 0.860 14.140 ;
        RECT 1.410 13.810 1.580 15.420 ;
        RECT 2.240 14.260 2.410 15.510 ;
        RECT 6.870 15.180 7.190 15.220 ;
        RECT 6.860 14.990 7.190 15.180 ;
        RECT 33.710 15.180 34.030 15.220 ;
        RECT 12.240 15.120 12.470 15.160 ;
        RECT 28.430 15.120 28.660 15.160 ;
        RECT 6.870 14.960 7.190 14.990 ;
        RECT 33.710 14.990 34.040 15.180 ;
        RECT 36.020 15.100 36.190 15.430 ;
        RECT 36.200 15.360 36.520 15.400 ;
        RECT 36.200 15.170 36.530 15.360 ;
        RECT 36.200 15.140 36.520 15.170 ;
        RECT 36.650 15.140 36.850 15.470 ;
        RECT 36.930 15.280 37.480 15.610 ;
        RECT 33.710 14.960 34.030 14.990 ;
        RECT 37.130 14.950 37.480 15.280 ;
        RECT 37.970 14.770 38.670 15.650 ;
        RECT 39.320 15.420 39.500 15.610 ;
        RECT 14.160 14.660 14.480 14.700 ;
        RECT 14.150 14.470 14.480 14.660 ;
        RECT 14.160 14.440 14.480 14.470 ;
        RECT 14.280 14.300 14.300 14.440 ;
        RECT 37.310 14.380 37.500 14.610 ;
        RECT 38.490 14.350 38.660 14.770 ;
        RECT 2.190 13.570 2.420 14.260 ;
        RECT 14.280 14.220 14.630 14.300 ;
        RECT 0.640 13.530 0.850 13.560 ;
        RECT 0.650 13.180 0.850 13.530 ;
        RECT 2.130 13.260 2.660 13.430 ;
        RECT 9.580 13.370 14.630 14.220 ;
        RECT 36.020 13.840 36.190 14.170 ;
        RECT 36.200 14.100 36.520 14.130 ;
        RECT 36.200 13.910 36.530 14.100 ;
        RECT 36.200 13.870 36.520 13.910 ;
        RECT 36.650 13.800 36.850 14.130 ;
        RECT 37.130 13.990 37.480 14.320 ;
        RECT 37.960 14.260 38.660 14.350 ;
        RECT 37.960 14.170 38.710 14.260 ;
        RECT 36.930 13.660 37.480 13.990 ;
        RECT 36.930 13.650 37.120 13.660 ;
        RECT 36.250 13.450 36.570 13.480 ;
        RECT 36.250 13.260 36.580 13.450 ;
        RECT 36.250 13.220 36.570 13.260 ;
        RECT 36.650 13.140 36.850 13.470 ;
        RECT 37.130 13.330 37.480 13.660 ;
        RECT 37.960 13.750 38.280 13.790 ;
        RECT 37.960 13.560 38.290 13.750 ;
        RECT 38.480 13.570 38.710 14.170 ;
        RECT 39.320 13.810 39.490 15.420 ;
        RECT 39.680 14.610 39.970 14.940 ;
        RECT 39.690 14.320 39.890 14.610 ;
        RECT 39.690 14.310 39.880 14.320 ;
        RECT 40.050 14.140 40.260 14.150 ;
        RECT 40.040 13.560 40.260 14.140 ;
        RECT 37.960 13.530 38.280 13.560 ;
        RECT 40.050 13.530 40.260 13.560 ;
        RECT 37.240 13.140 37.440 13.330 ;
        RECT 38.240 13.260 38.770 13.430 ;
        RECT 40.050 13.180 40.250 13.530 ;
        RECT 36.250 13.010 36.570 13.050 ;
        RECT 36.250 12.820 36.580 13.010 ;
        RECT 36.250 12.790 36.570 12.820 ;
        RECT 36.650 12.800 36.850 13.130 ;
        RECT 37.240 12.940 37.440 13.130 ;
        RECT 37.950 13.030 38.270 13.070 ;
        RECT 36.930 12.610 37.120 12.620 ;
        RECT 37.130 12.610 37.480 12.940 ;
        RECT 37.950 12.840 38.280 13.030 ;
        RECT 37.950 12.810 38.270 12.840 ;
        RECT 17.460 11.450 17.660 12.460 ;
        RECT 23.210 11.450 23.500 12.460 ;
        RECT 36.020 12.100 36.190 12.430 ;
        RECT 36.200 12.360 36.520 12.400 ;
        RECT 36.200 12.170 36.530 12.360 ;
        RECT 36.200 12.140 36.520 12.170 ;
        RECT 36.650 12.140 36.850 12.470 ;
        RECT 36.930 12.280 37.480 12.610 ;
        RECT 37.130 12.020 37.480 12.280 ;
        RECT 37.130 11.950 37.500 12.020 ;
        RECT 37.310 11.790 37.500 11.950 ;
        RECT 37.960 11.890 38.660 12.070 ;
        RECT 36.020 10.840 36.190 11.170 ;
        RECT 36.200 11.100 36.520 11.130 ;
        RECT 36.200 10.910 36.530 11.100 ;
        RECT 36.200 10.870 36.520 10.910 ;
        RECT 36.650 10.800 36.850 11.130 ;
        RECT 37.130 10.990 37.480 11.320 ;
        RECT 36.930 10.660 37.480 10.990 ;
        RECT 37.970 10.820 38.670 11.470 ;
        RECT 36.930 10.650 37.120 10.660 ;
        RECT 31.680 10.550 32.000 10.590 ;
        RECT 31.670 10.360 32.000 10.550 ;
        RECT 31.680 10.350 32.000 10.360 ;
        RECT 31.670 10.330 32.000 10.350 ;
        RECT 36.250 10.450 36.570 10.480 ;
        RECT 31.670 10.020 31.840 10.330 ;
        RECT 36.250 10.260 36.580 10.450 ;
        RECT 36.250 10.220 36.570 10.260 ;
        RECT 36.650 10.140 36.850 10.470 ;
        RECT 37.130 10.330 37.480 10.660 ;
        RECT 37.870 10.590 38.670 10.820 ;
        RECT 37.870 10.560 38.190 10.590 ;
        RECT 37.240 10.140 37.440 10.330 ;
        RECT 37.970 9.980 38.680 10.150 ;
        RECT 31.830 9.720 32.150 9.760 ;
        RECT 31.820 9.530 32.150 9.720 ;
        RECT 38.320 9.700 38.680 9.980 ;
        RECT 38.320 9.530 38.650 9.700 ;
        RECT 31.830 9.500 32.150 9.530 ;
        RECT 38.760 9.440 39.090 9.610 ;
        RECT 31.020 8.900 31.340 8.930 ;
        RECT 31.020 8.710 31.350 8.900 ;
        RECT 31.020 8.670 31.340 8.710 ;
        RECT 31.000 6.950 31.180 8.010 ;
        RECT 31.750 7.620 32.070 7.650 ;
        RECT 31.750 7.550 32.080 7.620 ;
        RECT 31.610 7.430 32.080 7.550 ;
        RECT 31.610 7.420 32.070 7.430 ;
        RECT 31.730 7.390 32.070 7.420 ;
        RECT 31.730 7.320 31.780 7.390 ;
        RECT 31.650 6.990 31.820 7.320 ;
        RECT 32.050 6.790 32.130 6.870 ;
        RECT 32.190 6.790 32.380 6.910 ;
        RECT 32.050 6.700 32.380 6.790 ;
        RECT 32.190 6.680 32.380 6.700 ;
        RECT 34.630 3.520 34.810 5.570 ;
        RECT 35.360 5.310 35.690 5.480 ;
        RECT 35.440 3.530 35.610 5.310 ;
        RECT 34.630 0.470 34.810 2.520 ;
        RECT 35.360 2.260 35.690 2.430 ;
        RECT 35.440 0.480 35.610 2.260 ;
      LAYER mcon ;
        RECT 1.350 21.670 1.620 21.940 ;
        RECT 39.280 21.670 39.550 21.940 ;
        RECT 1.350 19.940 1.620 20.210 ;
        RECT 39.280 19.940 39.550 20.210 ;
        RECT 2.480 19.160 2.660 19.330 ;
        RECT 0.670 18.860 0.840 19.030 ;
        RECT 1.020 18.020 1.200 18.210 ;
        RECT 2.220 18.710 2.390 18.880 ;
        RECT 2.220 18.260 2.390 18.430 ;
        RECT 14.220 18.170 14.390 18.340 ;
        RECT 38.510 18.710 38.680 18.880 ;
        RECT 40.060 18.860 40.230 19.030 ;
        RECT 38.510 18.260 38.680 18.430 ;
        RECT 6.960 17.760 7.130 17.930 ;
        RECT 33.770 17.760 33.940 17.930 ;
        RECT 39.700 18.020 39.880 18.210 ;
        RECT 13.410 16.230 13.580 16.400 ;
        RECT 27.320 16.230 27.490 16.400 ;
        RECT 36.310 15.830 36.480 16.000 ;
        RECT 37.970 15.790 38.140 15.960 ;
        RECT 1.020 14.380 1.200 14.570 ;
        RECT 6.960 15.000 7.130 15.170 ;
        RECT 33.770 15.000 33.940 15.170 ;
        RECT 36.260 15.180 36.430 15.350 ;
        RECT 37.250 15.440 37.420 15.610 ;
        RECT 14.250 14.480 14.420 14.650 ;
        RECT 37.320 14.410 37.490 14.580 ;
        RECT 2.220 14.060 2.390 14.230 ;
        RECT 0.670 13.560 0.840 13.730 ;
        RECT 2.220 13.610 2.390 13.780 ;
        RECT 2.480 13.260 2.660 13.430 ;
        RECT 36.260 13.920 36.430 14.090 ;
        RECT 37.250 13.660 37.420 13.830 ;
        RECT 38.510 14.060 38.680 14.230 ;
        RECT 36.310 13.270 36.480 13.440 ;
        RECT 39.700 14.380 39.880 14.570 ;
        RECT 38.020 13.570 38.190 13.740 ;
        RECT 38.510 13.610 38.680 13.780 ;
        RECT 40.060 13.560 40.230 13.730 ;
        RECT 36.310 12.830 36.480 13.000 ;
        RECT 38.010 12.850 38.180 13.020 ;
        RECT 17.470 12.220 17.640 12.390 ;
        RECT 17.480 11.500 17.650 11.670 ;
        RECT 23.260 12.220 23.430 12.390 ;
        RECT 36.260 12.180 36.430 12.350 ;
        RECT 37.250 12.440 37.420 12.610 ;
        RECT 37.320 11.820 37.490 11.990 ;
        RECT 23.260 11.500 23.430 11.670 ;
        RECT 36.260 10.920 36.430 11.090 ;
        RECT 37.250 10.660 37.420 10.830 ;
        RECT 31.770 10.370 31.940 10.540 ;
        RECT 36.310 10.270 36.480 10.440 ;
        RECT 37.930 10.600 38.100 10.770 ;
        RECT 31.920 9.540 32.090 9.710 ;
        RECT 31.080 8.720 31.250 8.890 ;
        RECT 31.810 7.440 31.980 7.610 ;
        RECT 32.200 6.710 32.370 6.880 ;
      LAYER met1 ;
        RECT 0.610 19.090 0.770 19.730 ;
        RECT 0.610 18.540 0.880 19.090 ;
        RECT 0.600 18.490 0.880 18.540 ;
        RECT 0.600 18.400 0.770 18.490 ;
        RECT 0.610 16.710 0.770 18.400 ;
        RECT 1.020 18.280 1.210 19.730 ;
        RECT 1.290 19.400 1.680 22.990 ;
        RECT 39.220 19.400 39.610 22.990 ;
        RECT 2.420 18.970 2.730 19.360 ;
        RECT 0.990 18.250 1.210 18.280 ;
        RECT 2.180 18.920 2.730 18.970 ;
        RECT 0.980 17.980 1.230 18.250 ;
        RECT 2.180 18.180 2.440 18.920 ;
        RECT 0.980 17.970 1.220 17.980 ;
        RECT 0.990 17.730 1.220 17.970 ;
        RECT 1.020 16.710 1.180 17.730 ;
        RECT 1.370 16.920 1.610 17.300 ;
        RECT 0.610 14.190 0.770 15.880 ;
        RECT 1.020 14.860 1.180 15.880 ;
        RECT 1.370 15.290 1.610 15.670 ;
        RECT 0.990 14.620 1.220 14.860 ;
        RECT 0.980 14.610 1.220 14.620 ;
        RECT 0.980 14.340 1.230 14.610 ;
        RECT 0.990 14.310 1.210 14.340 ;
        RECT 0.600 14.100 0.770 14.190 ;
        RECT 0.600 14.050 0.880 14.100 ;
        RECT 0.610 13.500 0.880 14.050 ;
        RECT 0.610 12.860 0.770 13.500 ;
        RECT 1.020 12.860 1.210 14.310 ;
        RECT 2.180 13.670 2.440 14.310 ;
        RECT 2.180 13.520 2.730 13.670 ;
        RECT 2.420 13.230 2.730 13.520 ;
        RECT 5.250 13.270 5.530 19.320 ;
        RECT 5.780 19.260 5.970 19.320 ;
        RECT 6.880 17.690 7.200 18.010 ;
        RECT 6.020 16.530 6.280 16.850 ;
        RECT 6.020 15.930 6.280 16.250 ;
        RECT 6.880 14.930 7.200 15.250 ;
        RECT 5.780 13.270 5.970 13.330 ;
        RECT 12.260 13.270 12.490 19.320 ;
        RECT 13.480 18.350 13.710 19.320 ;
        RECT 13.470 18.100 13.710 18.350 ;
        RECT 14.140 18.100 14.460 18.420 ;
        RECT 13.480 16.460 13.710 18.100 ;
        RECT 13.380 16.170 13.710 16.460 ;
        RECT 13.480 13.270 13.710 16.170 ;
        RECT 14.170 14.410 14.490 14.730 ;
        RECT 15.770 13.280 16.190 19.320 ;
        RECT 24.710 13.270 25.130 19.320 ;
        RECT 27.190 16.460 27.420 19.320 ;
        RECT 27.190 16.170 27.520 16.460 ;
        RECT 27.190 13.270 27.420 16.170 ;
        RECT 28.410 13.270 28.640 19.320 ;
        RECT 34.930 19.280 35.120 19.320 ;
        RECT 33.700 17.690 34.020 18.010 ;
        RECT 34.620 16.530 34.880 16.850 ;
        RECT 35.370 16.570 35.650 19.320 ;
        RECT 38.170 18.970 38.480 19.360 ;
        RECT 38.170 18.920 38.720 18.970 ;
        RECT 38.460 18.180 38.720 18.920 ;
        RECT 39.690 18.280 39.880 19.730 ;
        RECT 40.130 19.090 40.290 19.730 ;
        RECT 40.020 18.540 40.290 19.090 ;
        RECT 40.020 18.490 40.300 18.540 ;
        RECT 40.130 18.400 40.300 18.490 ;
        RECT 39.690 18.250 39.910 18.280 ;
        RECT 39.670 17.980 39.920 18.250 ;
        RECT 39.680 17.970 39.920 17.980 ;
        RECT 39.680 17.730 39.910 17.970 ;
        RECT 39.290 16.920 39.530 17.300 ;
        RECT 39.720 16.710 39.880 17.730 ;
        RECT 40.130 16.710 40.290 18.400 ;
        RECT 35.370 16.250 35.820 16.570 ;
        RECT 34.620 15.930 34.880 16.250 ;
        RECT 31.410 14.980 31.690 15.030 ;
        RECT 31.410 14.680 31.730 14.980 ;
        RECT 33.700 14.930 34.020 15.250 ;
        RECT 35.370 15.030 35.650 16.250 ;
        RECT 36.240 16.000 36.560 16.080 ;
        RECT 36.240 15.760 36.810 16.000 ;
        RECT 36.470 15.430 36.810 15.760 ;
        RECT 36.190 15.110 36.810 15.430 ;
        RECT 35.100 14.890 35.650 15.030 ;
        RECT 34.930 13.270 35.120 13.320 ;
        RECT 35.370 13.270 35.650 14.890 ;
        RECT 36.470 14.160 36.810 15.110 ;
        RECT 36.190 13.840 36.810 14.160 ;
        RECT 36.470 13.510 36.810 13.840 ;
        RECT 36.240 13.190 36.810 13.510 ;
        RECT 36.470 13.080 36.810 13.190 ;
        RECT 36.240 12.760 36.810 13.080 ;
        RECT 36.470 12.430 36.810 12.760 ;
        RECT 17.470 12.210 17.640 12.390 ;
        RECT 23.260 12.210 23.430 12.390 ;
        RECT 36.190 12.110 36.810 12.430 ;
        RECT 17.450 11.620 17.770 11.920 ;
        RECT 17.450 11.510 17.690 11.620 ;
        RECT 23.150 11.550 23.470 11.870 ;
        RECT 17.480 11.500 17.650 11.510 ;
        RECT 17.670 11.450 17.690 11.510 ;
        RECT 23.260 11.500 23.430 11.550 ;
        RECT 36.470 11.160 36.810 12.110 ;
        RECT 36.190 10.840 36.810 11.160 ;
        RECT 31.690 10.300 32.010 10.620 ;
        RECT 36.470 10.510 36.810 10.840 ;
        RECT 36.240 10.280 36.810 10.510 ;
        RECT 37.140 15.670 37.410 15.990 ;
        RECT 37.900 15.720 38.220 16.040 ;
        RECT 37.140 15.380 37.450 15.670 ;
        RECT 37.140 14.640 37.410 15.380 ;
        RECT 39.290 15.290 39.530 15.670 ;
        RECT 39.720 14.860 39.880 15.880 ;
        RECT 37.140 14.350 37.520 14.640 ;
        RECT 39.680 14.620 39.910 14.860 ;
        RECT 39.680 14.610 39.920 14.620 ;
        RECT 37.140 13.890 37.410 14.350 ;
        RECT 39.670 14.340 39.920 14.610 ;
        RECT 39.690 14.310 39.910 14.340 ;
        RECT 37.140 13.600 37.450 13.890 ;
        RECT 37.950 13.670 38.270 13.820 ;
        RECT 38.460 13.670 38.720 14.310 ;
        RECT 37.140 12.670 37.410 13.600 ;
        RECT 37.950 13.520 38.720 13.670 ;
        RECT 37.950 13.500 38.480 13.520 ;
        RECT 38.170 13.230 38.480 13.500 ;
        RECT 37.940 12.780 38.260 13.100 ;
        RECT 39.690 12.860 39.880 14.310 ;
        RECT 40.130 14.190 40.290 15.880 ;
        RECT 40.130 14.100 40.300 14.190 ;
        RECT 40.020 14.050 40.300 14.100 ;
        RECT 40.020 13.500 40.290 14.050 ;
        RECT 40.130 12.860 40.290 13.500 ;
        RECT 37.140 12.380 37.450 12.670 ;
        RECT 37.140 12.050 37.410 12.380 ;
        RECT 37.140 11.760 37.520 12.050 ;
        RECT 37.140 10.890 37.410 11.760 ;
        RECT 37.140 10.600 37.450 10.890 ;
        RECT 37.140 10.290 37.410 10.600 ;
        RECT 37.860 10.530 38.180 10.850 ;
        RECT 36.240 10.190 36.560 10.280 ;
        RECT 31.840 9.470 32.160 9.790 ;
        RECT 23.150 9.040 23.470 9.340 ;
        RECT 33.590 9.180 33.920 9.470 ;
        RECT 33.580 9.150 34.000 9.180 ;
        RECT 34.600 9.170 35.100 9.180 ;
        RECT 34.600 9.150 35.440 9.170 ;
        RECT 33.580 9.040 35.440 9.150 ;
        RECT 33.860 9.010 34.760 9.040 ;
        RECT 35.100 8.980 35.440 9.040 ;
        RECT 31.010 8.640 31.330 8.960 ;
        RECT 32.090 8.530 32.300 8.740 ;
        RECT 32.090 8.210 32.420 8.530 ;
        RECT 31.740 7.360 32.060 7.680 ;
        RECT 32.090 6.970 32.300 8.210 ;
        RECT 32.170 6.650 32.400 6.940 ;
      LAYER via ;
        RECT 2.440 18.950 2.700 19.210 ;
        RECT 2.440 13.380 2.700 13.640 ;
        RECT 6.910 17.720 7.170 17.980 ;
        RECT 6.020 16.560 6.280 16.820 ;
        RECT 6.020 15.960 6.280 16.220 ;
        RECT 6.910 14.960 7.170 15.220 ;
        RECT 14.170 18.130 14.430 18.390 ;
        RECT 14.200 14.440 14.460 14.700 ;
        RECT 33.730 17.720 33.990 17.980 ;
        RECT 34.620 16.560 34.880 16.820 ;
        RECT 38.200 18.950 38.460 19.210 ;
        RECT 35.560 16.280 35.820 16.540 ;
        RECT 34.620 15.960 34.880 16.220 ;
        RECT 31.440 14.700 31.700 14.960 ;
        RECT 33.730 14.960 33.990 15.220 ;
        RECT 36.270 15.790 36.530 16.050 ;
        RECT 36.220 15.140 36.480 15.400 ;
        RECT 36.220 13.870 36.480 14.130 ;
        RECT 36.270 13.220 36.530 13.480 ;
        RECT 36.270 12.790 36.530 13.050 ;
        RECT 36.220 12.140 36.480 12.400 ;
        RECT 17.480 11.640 17.740 11.900 ;
        RECT 23.180 11.580 23.440 11.840 ;
        RECT 36.220 10.870 36.480 11.130 ;
        RECT 31.720 10.330 31.980 10.590 ;
        RECT 36.270 10.220 36.530 10.480 ;
        RECT 37.930 15.750 38.190 16.010 ;
        RECT 37.980 13.640 38.240 13.790 ;
        RECT 37.980 13.530 38.460 13.640 ;
        RECT 38.200 13.380 38.460 13.530 ;
        RECT 37.970 12.810 38.230 13.070 ;
        RECT 37.890 10.560 38.150 10.820 ;
        RECT 31.870 9.500 32.130 9.760 ;
        RECT 23.180 9.060 23.440 9.320 ;
        RECT 33.620 9.190 33.890 9.450 ;
        RECT 31.040 8.670 31.300 8.930 ;
        RECT 32.160 8.240 32.420 8.500 ;
        RECT 31.770 7.390 32.030 7.650 ;
      LAYER met2 ;
        RECT 2.420 19.240 2.730 19.250 ;
        RECT 0.250 19.060 2.730 19.240 ;
        RECT 2.420 18.920 2.730 19.060 ;
        RECT 38.170 19.240 38.480 19.250 ;
        RECT 38.170 19.060 40.650 19.240 ;
        RECT 38.170 18.920 38.480 19.060 ;
        RECT 7.420 18.640 16.540 18.820 ;
        RECT 24.360 18.640 33.480 18.820 ;
        RECT 14.150 18.230 14.460 18.430 ;
        RECT 14.150 18.220 14.750 18.230 ;
        RECT 14.150 18.100 16.540 18.220 ;
        RECT 14.290 18.060 16.540 18.100 ;
        RECT 14.600 18.040 16.540 18.060 ;
        RECT 6.890 17.800 7.200 18.020 ;
        RECT 5.010 17.790 7.200 17.800 ;
        RECT 33.700 17.800 34.010 18.020 ;
        RECT 5.010 17.580 16.540 17.790 ;
        RECT 33.700 17.690 35.890 17.800 ;
        RECT 33.860 17.580 35.890 17.690 ;
        RECT 6.320 17.570 16.540 17.580 ;
        RECT 5.990 16.600 16.540 16.820 ;
        RECT 5.990 16.560 6.310 16.600 ;
        RECT 34.590 16.560 34.910 16.820 ;
        RECT 6.100 16.220 6.360 16.460 ;
        RECT 5.990 16.110 6.360 16.220 ;
        RECT 5.990 15.960 6.310 16.110 ;
        RECT 36.240 15.800 36.550 16.090 ;
        RECT 37.900 15.800 38.210 16.050 ;
        RECT 35.520 15.720 38.210 15.800 ;
        RECT 35.520 15.570 38.060 15.720 ;
        RECT 33.700 15.040 34.010 15.260 ;
        RECT 35.750 15.040 36.080 15.210 ;
        RECT 36.190 15.110 36.500 15.440 ;
        RECT 33.700 15.000 36.080 15.040 ;
        RECT 33.700 14.930 35.890 15.000 ;
        RECT 33.850 14.830 35.890 14.930 ;
        RECT 14.590 14.300 16.540 14.510 ;
        RECT 33.640 14.130 33.860 14.150 ;
        RECT 7.320 13.940 7.480 13.960 ;
        RECT 33.420 13.940 33.580 13.960 ;
        RECT 7.320 13.890 16.540 13.940 ;
        RECT 7.440 13.790 16.540 13.890 ;
        RECT 24.360 13.890 33.580 13.940 ;
        RECT 24.360 13.790 33.460 13.890 ;
        RECT 33.590 13.790 33.860 14.130 ;
        RECT 35.750 14.060 36.080 14.270 ;
        RECT 36.190 13.830 36.500 14.160 ;
        RECT 37.950 13.670 38.260 13.830 ;
        RECT 2.420 13.530 2.730 13.670 ;
        RECT 37.950 13.660 38.480 13.670 ;
        RECT 0.250 13.350 2.730 13.530 ;
        RECT 35.780 13.530 38.480 13.660 ;
        RECT 2.420 13.340 2.730 13.350 ;
        RECT 18.320 13.280 28.460 13.500 ;
        RECT 31.850 13.290 32.200 13.510 ;
        RECT 35.780 13.430 40.650 13.530 ;
        RECT 18.270 12.310 27.280 12.530 ;
        RECT 17.450 11.870 17.770 11.920 ;
        RECT 17.450 11.620 23.470 11.870 ;
        RECT 23.150 11.550 23.470 11.620 ;
        RECT 18.320 10.530 23.980 10.750 ;
        RECT 23.760 10.200 23.980 10.530 ;
        RECT 27.060 10.700 27.280 12.310 ;
        RECT 28.240 12.080 28.460 13.280 ;
        RECT 33.660 13.220 33.860 13.230 ;
        RECT 33.660 12.890 33.880 13.220 ;
        RECT 36.240 13.180 36.550 13.430 ;
        RECT 38.170 13.350 40.650 13.430 ;
        RECT 38.170 13.340 38.480 13.350 ;
        RECT 33.680 12.880 33.880 12.890 ;
        RECT 36.240 12.830 36.550 13.090 ;
        RECT 37.940 12.830 38.250 13.110 ;
        RECT 35.520 12.610 38.430 12.830 ;
        RECT 28.210 12.040 28.460 12.080 ;
        RECT 28.210 11.400 28.470 12.040 ;
        RECT 35.750 12.000 36.080 12.210 ;
        RECT 36.190 12.110 36.500 12.440 ;
        RECT 28.210 11.190 32.340 11.400 ;
        RECT 32.130 11.050 32.340 11.190 ;
        RECT 35.750 11.060 36.080 11.270 ;
        RECT 32.130 10.840 34.150 11.050 ;
        RECT 36.190 10.830 36.500 11.160 ;
        RECT 27.060 10.480 29.910 10.700 ;
        RECT 37.860 10.670 38.170 10.860 ;
        RECT 31.700 10.470 32.010 10.630 ;
        RECT 31.270 10.250 32.150 10.470 ;
        RECT 35.510 10.440 38.220 10.670 ;
        RECT 28.130 10.200 34.150 10.250 ;
        RECT 23.760 10.040 34.150 10.200 ;
        RECT 36.240 10.180 36.550 10.440 ;
        RECT 23.760 9.980 28.520 10.040 ;
        RECT 31.850 9.610 32.160 9.800 ;
        RECT 31.810 9.360 32.360 9.610 ;
        RECT 31.010 8.630 31.320 8.960 ;
        RECT 31.990 8.330 32.460 8.580 ;
        RECT 32.130 8.240 32.450 8.330 ;
        RECT 31.510 7.780 31.940 7.790 ;
        RECT 31.510 7.550 32.380 7.780 ;
        RECT 31.740 7.350 32.050 7.550 ;
  END
END sky130_hilas_TA2Cell_1FG

MACRO sky130_hilas_swc4x1cellOverlap
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x1cellOverlap ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 10.510 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 14.520 9.060 16.250 10.510 ;
        RECT 7.740 6.980 10.460 7.510 ;
        RECT 14.490 7.220 16.250 9.060 ;
        RECT 7.740 5.070 12.970 6.980 ;
        RECT 7.740 4.910 10.460 5.070 ;
        RECT 7.740 4.420 12.970 4.910 ;
        RECT 14.520 4.460 16.250 7.220 ;
        RECT 7.730 2.060 12.970 4.420 ;
        RECT 7.730 1.910 10.450 2.060 ;
        RECT 7.730 0.920 12.970 1.910 ;
        RECT 10.410 0.000 12.970 0.920 ;
      LAYER li1 ;
        RECT 14.910 7.670 15.460 8.100 ;
        RECT 8.140 5.940 10.090 7.110 ;
        RECT 10.650 6.630 10.970 6.670 ;
        RECT 10.650 6.510 10.980 6.630 ;
        RECT 10.650 6.410 11.090 6.510 ;
        RECT 10.750 6.340 11.090 6.410 ;
        RECT 12.370 6.240 12.570 6.590 ;
        RECT 10.650 6.080 10.970 6.120 ;
        RECT 10.650 5.890 10.980 6.080 ;
        RECT 10.650 5.860 11.090 5.890 ;
        RECT 10.750 5.720 11.090 5.860 ;
        RECT 11.640 5.620 11.840 6.220 ;
        RECT 12.370 6.210 12.580 6.240 ;
        RECT 12.360 5.620 12.580 6.210 ;
        RECT 8.140 4.410 10.090 5.580 ;
        RECT 10.750 4.120 11.090 4.260 ;
        RECT 10.650 4.090 11.090 4.120 ;
        RECT 8.130 2.850 10.080 4.020 ;
        RECT 10.650 3.900 10.980 4.090 ;
        RECT 10.650 3.860 10.970 3.900 ;
        RECT 11.640 3.760 11.840 4.360 ;
        RECT 12.360 3.770 12.580 4.360 ;
        RECT 12.370 3.740 12.580 3.770 ;
        RECT 10.650 3.640 10.970 3.660 ;
        RECT 10.650 3.330 11.090 3.640 ;
        RECT 10.650 3.310 10.970 3.330 ;
        RECT 12.370 3.230 12.570 3.740 ;
        RECT 10.650 3.070 10.970 3.110 ;
        RECT 10.650 2.880 10.980 3.070 ;
        RECT 10.650 2.850 11.090 2.880 ;
        RECT 10.750 2.710 11.090 2.850 ;
        RECT 11.640 2.610 11.840 3.210 ;
        RECT 12.370 3.200 12.580 3.230 ;
        RECT 12.360 2.610 12.580 3.200 ;
        RECT 8.130 1.310 10.080 2.480 ;
        RECT 10.750 1.120 11.090 1.260 ;
        RECT 10.650 1.090 11.090 1.120 ;
        RECT 10.650 0.900 10.980 1.090 ;
        RECT 10.650 0.860 10.970 0.900 ;
        RECT 11.640 0.760 11.840 1.360 ;
        RECT 12.360 0.770 12.580 1.360 ;
        RECT 12.370 0.740 12.580 0.770 ;
        RECT 10.750 0.570 11.090 0.640 ;
        RECT 10.650 0.470 11.090 0.570 ;
        RECT 10.650 0.350 10.980 0.470 ;
        RECT 12.370 0.390 12.570 0.740 ;
        RECT 10.650 0.310 10.970 0.350 ;
      LAYER mcon ;
        RECT 14.910 7.750 15.180 8.020 ;
        RECT 8.620 6.770 8.790 6.940 ;
        RECT 8.620 6.430 8.790 6.600 ;
        RECT 10.710 6.450 10.880 6.620 ;
        RECT 8.620 6.090 8.790 6.260 ;
        RECT 10.710 5.900 10.880 6.070 ;
        RECT 11.650 6.010 11.820 6.180 ;
        RECT 12.380 6.040 12.550 6.210 ;
        RECT 8.620 5.240 8.790 5.410 ;
        RECT 8.620 4.900 8.790 5.070 ;
        RECT 8.620 4.560 8.790 4.730 ;
        RECT 10.710 3.910 10.880 4.080 ;
        RECT 8.610 3.680 8.780 3.850 ;
        RECT 11.650 3.800 11.820 3.970 ;
        RECT 12.380 3.770 12.550 3.940 ;
        RECT 8.610 3.340 8.780 3.510 ;
        RECT 9.130 3.400 9.310 3.570 ;
        RECT 10.710 3.360 10.880 3.610 ;
        RECT 8.610 3.000 8.780 3.170 ;
        RECT 10.710 2.890 10.880 3.060 ;
        RECT 11.650 3.000 11.820 3.170 ;
        RECT 12.380 3.030 12.550 3.200 ;
        RECT 8.610 2.140 8.780 2.310 ;
        RECT 8.610 1.800 8.780 1.970 ;
        RECT 8.610 1.460 8.780 1.630 ;
        RECT 10.710 0.910 10.880 1.080 ;
        RECT 11.650 0.800 11.820 0.970 ;
        RECT 12.380 0.770 12.550 0.940 ;
        RECT 10.710 0.360 10.880 0.530 ;
      LAYER met1 ;
        RECT 14.850 7.210 15.240 9.070 ;
        RECT 8.580 6.520 8.840 7.000 ;
        RECT 0.360 0.460 0.760 6.450 ;
        RECT 8.570 6.000 8.840 6.520 ;
        RECT 10.640 6.380 10.960 6.700 ;
        RECT 11.640 6.240 11.800 6.970 ;
        RECT 11.640 6.220 11.840 6.240 ;
        RECT 8.570 5.550 8.830 6.000 ;
        RECT 10.640 5.830 10.960 6.150 ;
        RECT 11.620 5.980 11.850 6.220 ;
        RECT 11.640 5.930 11.850 5.980 ;
        RECT 12.010 5.930 12.200 6.920 ;
        RECT 12.450 6.270 12.610 6.970 ;
        RECT 8.580 4.990 8.840 5.470 ;
        RECT 11.640 5.070 11.800 5.930 ;
        RECT 12.030 5.810 12.200 5.930 ;
        RECT 12.040 5.070 12.200 5.810 ;
        RECT 12.340 5.720 12.610 6.270 ;
        RECT 12.340 5.670 12.620 5.720 ;
        RECT 12.450 5.580 12.620 5.670 ;
        RECT 12.450 5.070 12.610 5.580 ;
        RECT 8.570 4.470 8.840 4.990 ;
        RECT 8.570 4.020 8.830 4.470 ;
        RECT 8.570 3.430 8.830 3.910 ;
        RECT 10.640 3.830 10.960 4.150 ;
        RECT 11.640 4.050 11.800 4.910 ;
        RECT 12.040 4.170 12.200 4.910 ;
        RECT 12.450 4.400 12.610 4.910 ;
        RECT 12.450 4.310 12.620 4.400 ;
        RECT 12.030 4.050 12.200 4.170 ;
        RECT 11.640 4.000 11.850 4.050 ;
        RECT 11.620 3.760 11.850 4.000 ;
        RECT 11.640 3.740 11.840 3.760 ;
        RECT 9.180 3.600 9.310 3.620 ;
        RECT 8.560 2.910 8.830 3.430 ;
        RECT 9.100 3.370 9.340 3.600 ;
        RECT 9.200 3.330 9.310 3.370 ;
        RECT 10.640 3.280 10.960 3.690 ;
        RECT 11.640 3.230 11.800 3.740 ;
        RECT 11.640 3.210 11.840 3.230 ;
        RECT 8.560 2.460 8.820 2.910 ;
        RECT 10.640 2.820 10.960 3.140 ;
        RECT 11.620 2.970 11.850 3.210 ;
        RECT 11.640 2.920 11.850 2.970 ;
        RECT 12.010 2.920 12.200 4.050 ;
        RECT 12.340 4.260 12.620 4.310 ;
        RECT 12.340 3.710 12.610 4.260 ;
        RECT 12.450 3.260 12.610 3.710 ;
        RECT 8.570 1.890 8.830 2.370 ;
        RECT 11.640 2.060 11.800 2.920 ;
        RECT 12.030 2.800 12.200 2.920 ;
        RECT 12.040 2.060 12.200 2.800 ;
        RECT 12.340 2.710 12.610 3.260 ;
        RECT 12.340 2.660 12.620 2.710 ;
        RECT 12.450 2.570 12.620 2.660 ;
        RECT 12.450 2.060 12.610 2.570 ;
        RECT 8.560 1.370 8.830 1.890 ;
        RECT 8.560 0.920 8.820 1.370 ;
        RECT 10.640 0.830 10.960 1.150 ;
        RECT 11.640 1.050 11.800 1.910 ;
        RECT 12.040 1.170 12.200 1.910 ;
        RECT 12.450 1.400 12.610 1.910 ;
        RECT 12.450 1.310 12.620 1.400 ;
        RECT 12.030 1.050 12.200 1.170 ;
        RECT 11.640 1.000 11.850 1.050 ;
        RECT 11.620 0.760 11.850 1.000 ;
        RECT 11.640 0.740 11.840 0.760 ;
        RECT 10.640 0.280 10.960 0.600 ;
        RECT 11.640 0.010 11.800 0.740 ;
        RECT 12.010 0.060 12.200 1.050 ;
        RECT 12.340 1.260 12.620 1.310 ;
        RECT 12.340 0.710 12.610 1.260 ;
        RECT 12.450 0.010 12.610 0.710 ;
      LAYER via ;
        RECT 10.670 6.410 10.930 6.670 ;
        RECT 10.670 5.860 10.930 6.120 ;
        RECT 10.670 3.860 10.930 4.120 ;
        RECT 10.670 3.310 10.930 3.660 ;
        RECT 10.670 2.850 10.930 3.110 ;
        RECT 10.670 0.860 10.930 1.120 ;
        RECT 10.670 0.310 10.930 0.570 ;
      LAYER met2 ;
        RECT 10.640 6.420 10.950 6.710 ;
        RECT 10.640 6.380 12.970 6.420 ;
        RECT 10.790 6.240 12.970 6.380 ;
        RECT 0.000 5.940 7.610 6.010 ;
        RECT 10.640 5.990 10.950 6.160 ;
        RECT 0.000 5.830 7.640 5.940 ;
        RECT 10.410 5.810 10.500 5.990 ;
        RECT 10.640 5.830 12.970 5.990 ;
        RECT 10.800 5.810 12.970 5.830 ;
        RECT 0.000 5.400 9.740 5.580 ;
        RECT 0.000 4.520 7.610 4.580 ;
        RECT 0.000 4.400 7.640 4.520 ;
        RECT 0.000 4.080 7.600 4.150 ;
        RECT 0.000 3.970 7.640 4.080 ;
        RECT 10.410 3.990 10.500 4.170 ;
        RECT 10.800 4.150 12.970 4.170 ;
        RECT 10.640 3.990 12.970 4.150 ;
        RECT 10.640 3.820 10.950 3.990 ;
        RECT 10.790 3.700 12.970 3.740 ;
        RECT 10.640 3.560 12.970 3.700 ;
        RECT 10.640 3.410 10.950 3.560 ;
        RECT 10.640 3.270 12.970 3.410 ;
        RECT 10.790 3.230 12.970 3.270 ;
        RECT 0.020 2.820 7.640 2.990 ;
        RECT 10.640 2.980 10.950 3.150 ;
        RECT 10.410 2.800 10.500 2.980 ;
        RECT 10.640 2.820 12.970 2.980 ;
        RECT 10.800 2.800 12.970 2.820 ;
        RECT 0.020 2.400 7.640 2.570 ;
        RECT 0.020 1.420 7.640 1.590 ;
        RECT 0.800 1.330 2.340 1.420 ;
        RECT 0.020 0.980 7.640 1.150 ;
        RECT 10.410 0.990 10.500 1.170 ;
        RECT 10.800 1.150 12.970 1.170 ;
        RECT 10.640 0.990 12.970 1.150 ;
        RECT 10.640 0.820 10.950 0.990 ;
        RECT 10.790 0.600 12.970 0.740 ;
        RECT 10.640 0.560 12.970 0.600 ;
        RECT 10.640 0.270 10.950 0.560 ;
  END
END sky130_hilas_swc4x1cellOverlap

MACRO sky130_hilas_capacitorSize02
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize02 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.610 BY 7.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 7.660 2.390 7.970 2.670 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.020 2.370 0.290 2.650 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 0.000 4.850 7.970 5.030 ;
        RECT 0.000 4.420 7.970 4.600 ;
        RECT 0.030 3.420 7.970 3.600 ;
        RECT 0.030 3.090 7.970 3.170 ;
        RECT 0.030 2.990 8.090 3.090 ;
        RECT 0.600 2.670 0.970 2.990 ;
        RECT 7.720 2.690 8.090 2.990 ;
        RECT 0.030 1.840 7.970 2.010 ;
        RECT 0.030 1.420 7.970 1.590 ;
        RECT 0.030 0.440 7.970 0.610 ;
        RECT 0.030 0.000 7.970 0.170 ;
      LAYER via2 ;
        RECT 0.650 2.730 0.930 3.010 ;
        RECT 7.770 2.750 8.050 3.030 ;
      LAYER met3 ;
        RECT 5.380 7.840 7.690 7.870 ;
        RECT 0.380 2.470 1.170 3.220 ;
        RECT 5.380 2.060 9.610 7.840 ;
        RECT 7.660 2.040 9.610 2.060 ;
      LAYER via3 ;
        RECT 0.570 2.620 1.000 3.100 ;
        RECT 7.690 2.640 8.120 3.120 ;
      LAYER met4 ;
        RECT 0.470 2.770 1.130 3.190 ;
        RECT 5.760 3.140 8.770 3.610 ;
        RECT 1.160 2.770 2.170 2.780 ;
        RECT 0.450 2.270 3.800 2.770 ;
        RECT 7.590 2.550 8.250 3.140 ;
        RECT 0.450 2.260 1.520 2.270 ;
        RECT 3.160 1.150 3.790 2.270 ;
        RECT 3.160 0.850 5.310 1.150 ;
        RECT 3.490 0.840 5.310 0.850 ;
  END
END sky130_hilas_capacitorSize02

MACRO sky130_hilas_TopProtectStructure
  CLASS CORE ;
  FOREIGN sky130_hilas_TopProtectStructure ;
  ORIGIN 0.000 0.000 ;
  SIZE 393.720 BY 458.320 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN IO07
    PORT
      LAYER met1 ;
        RECT 371.600 180.790 372.850 184.680 ;
    END
  END IO07
  PIN IO08
    PORT
      LAYER met1 ;
        RECT 371.600 209.400 372.850 213.290 ;
    END
  END IO08
  PIN IO09
    PORT
      LAYER met1 ;
        RECT 371.580 237.980 372.830 241.870 ;
    END
  END IO09
  PIN IO10
    PORT
      LAYER met1 ;
        RECT 371.600 266.590 372.850 270.480 ;
    END
  END IO10
  PIN IO11
    PORT
      LAYER met1 ;
        RECT 371.590 295.150 372.840 299.040 ;
    END
  END IO11
  PIN IO12
    PORT
      LAYER met1 ;
        RECT 371.590 323.750 372.840 327.640 ;
    END
  END IO12
  PIN IO13
    PORT
      LAYER met1 ;
        RECT 371.600 352.350 372.850 356.240 ;
    END
  END IO13
  PIN IO25
    PORT
      LAYER met1 ;
        RECT 0.000 353.050 1.250 356.940 ;
    END
  END IO25
  PIN IO26
    PORT
      LAYER met1 ;
        RECT 0.010 324.470 1.260 328.360 ;
    END
  END IO26
  PIN IO27
    PORT
      LAYER met1 ;
        RECT 0.000 295.870 1.250 299.760 ;
    END
  END IO27
  PIN IO28
    PORT
      LAYER met1 ;
        RECT 0.020 267.280 1.270 271.170 ;
    END
  END IO28
  PIN IO29
    PORT
      LAYER met1 ;
        RECT 0.010 238.700 1.260 242.590 ;
    END
  END IO29
  PIN IO30
    PORT
      LAYER met1 ;
        RECT 0.000 210.100 1.250 213.990 ;
    END
  END IO30
  PIN IO31
    PORT
      LAYER met1 ;
        RECT 0.010 181.520 1.260 185.410 ;
    END
  END IO31
  PIN IO32
    PORT
      LAYER met1 ;
        RECT 0.040 152.940 1.290 156.830 ;
    END
  END IO32
  PIN IO33
    PORT
      LAYER met1 ;
        RECT 0.020 124.330 1.270 128.220 ;
    END
  END IO33
  PIN IO34
    PORT
      LAYER met1 ;
        RECT 0.010 95.740 1.260 99.630 ;
    END
  END IO34
  PIN IO35
    PORT
      LAYER met1 ;
        RECT 0.010 67.150 1.260 71.040 ;
    END
  END IO35
  PIN IO36
    PORT
      LAYER met1 ;
        RECT 0.020 38.560 1.270 42.450 ;
    END
  END IO36
  PIN IO37
    PORT
      LAYER met1 ;
        RECT 0.020 9.980 1.270 13.870 ;
    END
  END IO37
  PIN VSSA1
    PORT
      LAYER met2 ;
        RECT 3.420 385.010 16.350 385.020 ;
        RECT 3.290 383.620 16.350 385.010 ;
        RECT 3.290 382.100 5.580 383.620 ;
        RECT 3.740 382.060 5.580 382.100 ;
        RECT 4.180 373.540 5.580 382.060 ;
    END
  END VSSA1
  PIN ANALOG10
    ANTENNAGATEAREA 0.136700 ;
    ANTENNADIFFAREA 1261.030029 ;
    PORT
      LAYER nwell ;
        RECT 24.920 444.600 30.860 456.650 ;
        RECT 24.920 416.010 30.860 428.060 ;
        RECT 24.920 387.420 30.860 399.470 ;
        RECT 30.800 381.200 42.850 387.140 ;
        RECT 59.390 381.200 71.440 387.140 ;
        RECT 87.980 381.200 100.030 387.140 ;
        RECT 24.920 358.830 30.860 370.880 ;
        RECT 24.920 330.240 30.860 342.290 ;
        RECT 24.920 301.650 30.860 313.700 ;
        RECT 24.920 273.060 30.860 285.110 ;
        RECT 24.920 244.470 30.860 256.520 ;
        RECT 24.920 215.880 30.860 227.930 ;
        RECT 24.920 187.290 30.860 199.340 ;
        RECT 24.920 158.700 30.860 170.750 ;
        RECT 24.920 130.110 30.860 142.160 ;
        RECT 24.920 101.520 30.860 113.570 ;
      LAYER met2 ;
        RECT 23.990 431.130 25.390 458.320 ;
        RECT 30.290 457.800 31.690 458.320 ;
        RECT 30.290 457.720 31.820 457.800 ;
        RECT 30.290 456.710 32.330 457.720 ;
        RECT 27.280 456.070 32.330 456.710 ;
        RECT 30.290 455.790 32.330 456.070 ;
        RECT 30.290 455.170 32.400 455.790 ;
        RECT 23.990 430.620 25.400 431.130 ;
        RECT 23.990 430.450 26.510 430.620 ;
        RECT 23.990 430.200 25.400 430.450 ;
        RECT 23.990 402.540 25.390 430.200 ;
        RECT 30.290 429.210 31.690 455.170 ;
        RECT 30.290 429.130 31.820 429.210 ;
        RECT 30.290 428.120 32.330 429.130 ;
        RECT 27.280 427.480 32.330 428.120 ;
        RECT 30.290 427.200 32.330 427.480 ;
        RECT 30.290 426.580 32.400 427.200 ;
        RECT 23.990 402.030 25.400 402.540 ;
        RECT 23.990 401.860 26.510 402.030 ;
        RECT 23.990 401.610 25.400 401.860 ;
        RECT 23.990 388.070 25.390 401.610 ;
        RECT 30.290 400.620 31.690 426.580 ;
        RECT 30.290 400.540 31.820 400.620 ;
        RECT 30.290 399.530 32.330 400.540 ;
        RECT 27.280 398.890 32.330 399.530 ;
        RECT 30.290 398.610 32.330 398.890 ;
        RECT 30.290 397.990 32.400 398.610 ;
        RECT 30.290 388.070 31.690 397.990 ;
        RECT 15.930 386.670 101.700 388.070 ;
        RECT 16.400 386.660 17.330 386.670 ;
        RECT 16.650 385.550 16.820 386.660 ;
        RECT 23.990 381.770 25.390 386.670 ;
        RECT 30.290 381.770 31.690 386.670 ;
        RECT 44.990 386.660 45.920 386.670 ;
        RECT 73.580 386.660 74.510 386.670 ;
        RECT 45.240 385.550 45.410 386.660 ;
        RECT 73.830 385.550 74.000 386.660 ;
        RECT 42.270 381.770 42.910 384.780 ;
        RECT 70.860 381.770 71.500 384.780 ;
        RECT 99.450 381.770 100.090 384.780 ;
        RECT 15.930 380.370 101.700 381.770 ;
        RECT 23.990 373.950 25.390 380.370 ;
        RECT 23.990 373.440 25.400 373.950 ;
        RECT 23.990 373.270 26.510 373.440 ;
        RECT 23.990 373.020 25.400 373.270 ;
        RECT 14.870 359.920 17.760 361.880 ;
        RECT 23.990 359.920 25.390 373.020 ;
        RECT 30.290 372.030 31.690 380.370 ;
        RECT 41.370 380.240 44.000 380.370 ;
        RECT 69.960 380.240 72.590 380.370 ;
        RECT 98.550 380.240 101.180 380.370 ;
        RECT 41.370 379.730 43.920 380.240 ;
        RECT 69.960 379.730 72.510 380.240 ;
        RECT 98.550 379.730 101.100 380.240 ;
        RECT 41.370 379.660 41.990 379.730 ;
        RECT 69.960 379.660 70.580 379.730 ;
        RECT 98.550 379.660 99.170 379.730 ;
        RECT 30.290 371.950 31.820 372.030 ;
        RECT 30.290 370.940 32.330 371.950 ;
        RECT 27.280 370.300 32.330 370.940 ;
        RECT 30.290 370.020 32.330 370.300 ;
        RECT 30.290 369.400 32.400 370.020 ;
        RECT 27.100 364.260 29.740 365.440 ;
        RECT 30.290 364.260 31.690 369.400 ;
        RECT 27.020 362.010 127.330 364.260 ;
        RECT 27.100 361.840 29.740 362.010 ;
        RECT 30.290 359.920 31.690 362.010 ;
        RECT 14.840 358.060 126.960 359.920 ;
        RECT 23.990 355.480 25.390 358.060 ;
        RECT 30.290 355.480 31.690 358.060 ;
        RECT 23.730 353.400 127.250 355.480 ;
        RECT 23.730 344.850 25.810 353.400 ;
        RECT 30.290 350.600 31.690 353.400 ;
        RECT 27.890 348.520 127.730 350.600 ;
        RECT 23.730 344.680 26.510 344.850 ;
        RECT 23.730 333.290 25.810 344.680 ;
        RECT 27.890 342.350 29.970 348.520 ;
        RECT 30.290 343.440 31.690 348.520 ;
        RECT 32.230 343.700 127.730 345.780 ;
        RECT 30.290 343.360 31.820 343.440 ;
        RECT 32.230 343.360 34.310 343.700 ;
        RECT 30.290 342.350 34.310 343.360 ;
        RECT 27.280 341.710 34.310 342.350 ;
        RECT 23.660 329.920 26.000 333.290 ;
        RECT 23.730 329.050 25.810 329.920 ;
        RECT 23.990 316.770 25.390 329.050 ;
        RECT 23.990 316.260 25.400 316.770 ;
        RECT 23.990 316.090 26.510 316.260 ;
        RECT 23.990 315.840 25.400 316.090 ;
        RECT 23.990 288.180 25.390 315.840 ;
        RECT 27.890 313.760 29.970 341.710 ;
        RECT 30.290 340.810 34.310 341.710 ;
        RECT 30.290 314.850 31.690 340.810 ;
        RECT 30.290 314.770 31.820 314.850 ;
        RECT 32.230 314.770 34.310 340.810 ;
        RECT 30.290 313.760 34.310 314.770 ;
        RECT 27.280 313.120 34.310 313.760 ;
        RECT 27.890 304.690 29.970 313.120 ;
        RECT 27.670 301.280 29.970 304.690 ;
        RECT 27.890 300.950 29.970 301.280 ;
        RECT 30.290 312.220 34.310 313.120 ;
        RECT 23.990 287.670 25.400 288.180 ;
        RECT 23.990 287.500 26.510 287.670 ;
        RECT 23.990 287.250 25.400 287.500 ;
        RECT 23.990 259.590 25.390 287.250 ;
        RECT 30.290 286.260 31.690 312.220 ;
        RECT 30.290 286.180 31.820 286.260 ;
        RECT 32.230 286.180 34.310 312.220 ;
        RECT 30.290 285.170 34.310 286.180 ;
        RECT 27.280 284.530 34.310 285.170 ;
        RECT 30.290 283.630 34.310 284.530 ;
        RECT 23.990 259.080 25.400 259.590 ;
        RECT 23.990 258.910 26.510 259.080 ;
        RECT 23.990 258.660 25.400 258.910 ;
        RECT 23.990 231.000 25.390 258.660 ;
        RECT 30.290 257.670 31.690 283.630 ;
        RECT 32.230 276.210 34.310 283.630 ;
        RECT 32.020 272.610 34.590 276.210 ;
        RECT 32.230 272.570 34.310 272.610 ;
        RECT 30.290 257.590 31.820 257.670 ;
        RECT 30.290 256.580 32.330 257.590 ;
        RECT 27.280 255.940 32.330 256.580 ;
        RECT 30.290 255.660 32.330 255.940 ;
        RECT 30.290 255.040 32.400 255.660 ;
        RECT 23.990 230.490 25.400 231.000 ;
        RECT 23.990 230.320 26.510 230.490 ;
        RECT 23.990 230.070 25.400 230.320 ;
        RECT 23.990 202.410 25.390 230.070 ;
        RECT 30.290 229.080 31.690 255.040 ;
        RECT 30.290 229.000 31.820 229.080 ;
        RECT 30.290 227.990 32.330 229.000 ;
        RECT 27.280 227.350 32.330 227.990 ;
        RECT 30.290 227.070 32.330 227.350 ;
        RECT 30.290 226.450 32.400 227.070 ;
        RECT 23.990 201.900 25.400 202.410 ;
        RECT 23.990 201.730 26.510 201.900 ;
        RECT 23.990 201.480 25.400 201.730 ;
        RECT 23.990 173.820 25.390 201.480 ;
        RECT 30.290 200.490 31.690 226.450 ;
        RECT 30.290 200.410 31.820 200.490 ;
        RECT 30.290 199.400 32.330 200.410 ;
        RECT 27.280 198.760 32.330 199.400 ;
        RECT 30.290 198.480 32.330 198.760 ;
        RECT 30.290 197.860 32.400 198.480 ;
        RECT 23.990 173.310 25.400 173.820 ;
        RECT 23.990 173.140 26.510 173.310 ;
        RECT 23.990 172.890 25.400 173.140 ;
        RECT 23.990 145.230 25.390 172.890 ;
        RECT 30.290 171.900 31.690 197.860 ;
        RECT 30.290 171.820 31.820 171.900 ;
        RECT 30.290 170.810 32.330 171.820 ;
        RECT 27.280 170.170 32.330 170.810 ;
        RECT 30.290 169.890 32.330 170.170 ;
        RECT 30.290 169.270 32.400 169.890 ;
        RECT 23.990 144.720 25.400 145.230 ;
        RECT 23.990 144.550 26.510 144.720 ;
        RECT 23.990 144.300 25.400 144.550 ;
        RECT 23.990 116.640 25.390 144.300 ;
        RECT 30.290 143.310 31.690 169.270 ;
        RECT 30.290 143.230 31.820 143.310 ;
        RECT 30.290 142.220 32.330 143.230 ;
        RECT 27.280 141.580 32.330 142.220 ;
        RECT 30.290 141.300 32.330 141.580 ;
        RECT 30.290 140.680 32.400 141.300 ;
        RECT 23.990 116.130 25.400 116.640 ;
        RECT 23.990 115.960 26.510 116.130 ;
        RECT 23.990 115.710 25.400 115.960 ;
        RECT 23.990 88.050 25.390 115.710 ;
        RECT 30.290 114.720 31.690 140.680 ;
        RECT 30.290 114.640 31.820 114.720 ;
        RECT 30.290 113.630 32.330 114.640 ;
        RECT 27.280 112.990 32.330 113.630 ;
        RECT 30.290 112.710 32.330 112.990 ;
        RECT 30.290 112.090 32.400 112.710 ;
        RECT 23.990 87.540 25.400 88.050 ;
        RECT 23.990 87.370 26.510 87.540 ;
        RECT 23.990 87.120 25.400 87.370 ;
        RECT 23.990 86.650 25.390 87.120 ;
        RECT 30.290 86.650 31.690 112.090 ;
    END
  END ANALOG10
  PIN ANALOG09
    PORT
      LAYER met1 ;
        RECT 52.230 389.570 56.130 390.160 ;
        RECT 52.230 389.070 52.520 389.570 ;
        RECT 52.210 387.900 56.100 389.070 ;
    END
  END ANALOG09
  PIN ANALOG08
    PORT
      LAYER met1 ;
        RECT 80.820 389.570 84.720 390.160 ;
        RECT 80.820 389.070 81.110 389.570 ;
        RECT 80.800 387.900 84.690 389.070 ;
    END
  END ANALOG08
  PIN ANALOG07
    PORT
      LAYER met1 ;
        RECT 122.700 387.930 126.590 389.100 ;
    END
  END ANALOG07
  PIN ANALOG06
    PORT
      LAYER met1 ;
        RECT 164.840 389.570 168.740 390.160 ;
        RECT 164.840 389.080 165.130 389.570 ;
        RECT 164.820 387.910 168.710 389.080 ;
    END
  END ANALOG06
  PIN ANALOG05
    PORT
      LAYER met1 ;
        RECT 193.430 389.570 197.330 390.160 ;
        RECT 193.430 389.080 193.720 389.570 ;
        RECT 193.410 387.910 197.300 389.080 ;
    END
  END ANALOG05
  PIN ANALOG04
    PORT
      LAYER met1 ;
        RECT 222.020 389.570 225.920 390.160 ;
        RECT 222.020 389.080 222.310 389.570 ;
        RECT 222.010 387.910 225.900 389.080 ;
    END
  END ANALOG04
  PIN ANALOG03
    PORT
      LAYER met1 ;
        RECT 250.610 389.570 254.510 390.160 ;
        RECT 250.610 389.080 250.900 389.570 ;
        RECT 250.600 387.910 254.490 389.080 ;
    END
  END ANALOG03
  PIN ANALOG02
    PORT
      LAYER met1 ;
        RECT 279.200 389.570 283.100 390.160 ;
        RECT 279.200 389.080 279.490 389.570 ;
        RECT 279.190 387.910 283.080 389.080 ;
    END
  END ANALOG02
  PIN ANALOG01
    PORT
      LAYER met1 ;
        RECT 307.790 389.570 311.690 390.160 ;
        RECT 307.790 389.070 308.080 389.570 ;
        RECT 307.780 387.900 311.670 389.070 ;
    END
  END ANALOG01
  PIN ANALOG00
    PORT
      LAYER met1 ;
        RECT 336.380 389.570 340.280 390.160 ;
        RECT 336.380 389.070 336.670 389.570 ;
        RECT 336.370 387.900 340.260 389.070 ;
    END
  END ANALOG00
  PIN VSSA1
    PORT
      LAYER met2 ;
        RECT 368.490 385.020 369.680 385.030 ;
        RECT 356.690 384.500 369.680 385.020 ;
        RECT 356.480 383.740 369.680 384.500 ;
        RECT 367.520 382.420 369.680 383.740 ;
        RECT 367.520 373.190 368.800 382.420 ;
        RECT 368.040 372.450 368.800 373.190 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.150 0.330 5.550 2.300 ;
    END
    PORT
      LAYER met2 ;
        RECT 368.060 173.390 368.800 173.730 ;
        RECT 367.400 172.990 368.810 173.390 ;
        RECT 367.420 172.300 368.800 172.990 ;
        RECT 367.410 171.130 368.810 172.300 ;
    END
  END VSSA1
  PIN VDDA1
    PORT
      LAYER met2 ;
        RECT 10.450 0.000 11.850 3.660 ;
    END
    PORT
      LAYER met2 ;
        RECT 361.080 172.360 362.480 173.140 ;
        RECT 361.070 172.240 362.480 172.360 ;
        RECT 361.060 172.090 362.480 172.240 ;
        RECT 361.060 171.190 362.470 172.090 ;
    END
  END VDDA1
  PIN LADATAOUT01
    PORT
      LAYER met2 ;
        RECT 146.050 6.780 148.070 301.800 ;
        RECT 146.050 5.220 148.080 6.780 ;
        RECT 146.050 5.210 148.070 5.220 ;
    END
  END LADATAOUT01
  PIN LADATAOUT00
    PORT
      LAYER met2 ;
        RECT 141.990 5.210 144.010 301.800 ;
    END
  END LADATAOUT00
  PIN LADATAOUT02
    PORT
      LAYER met2 ;
        RECT 150.020 6.770 152.040 301.800 ;
        RECT 150.010 5.210 152.040 6.770 ;
    END
  END LADATAOUT02
  PIN LADATAOUT03
    PORT
      LAYER met2 ;
        RECT 154.020 6.770 156.040 301.800 ;
        RECT 154.010 5.210 156.040 6.770 ;
    END
  END LADATAOUT03
  PIN LADATAOUT04
    PORT
      LAYER met2 ;
        RECT 158.070 5.210 160.090 301.800 ;
    END
  END LADATAOUT04
  PIN LADATAOUT05
    PORT
      LAYER met2 ;
        RECT 162.080 6.780 164.100 301.800 ;
        RECT 162.070 5.220 164.100 6.780 ;
        RECT 162.080 5.210 164.100 5.220 ;
    END
  END LADATAOUT05
  PIN LADATAOUT06
    PORT
      LAYER met2 ;
        RECT 166.080 5.210 168.100 301.800 ;
    END
  END LADATAOUT06
  PIN LADATAOUT07
    PORT
      LAYER met2 ;
        RECT 170.170 5.210 172.190 301.800 ;
    END
  END LADATAOUT07
  PIN LADATAOUT08
    PORT
      LAYER met2 ;
        RECT 174.300 6.770 176.320 301.800 ;
        RECT 174.290 5.210 176.320 6.770 ;
    END
  END LADATAOUT08
  PIN LADATAOUT09
    PORT
      LAYER met2 ;
        RECT 178.300 6.770 180.320 301.800 ;
        RECT 178.290 5.210 180.320 6.770 ;
    END
  END LADATAOUT09
  PIN LADATAOUT10
    PORT
      LAYER met2 ;
        RECT 182.260 6.770 184.280 301.800 ;
        RECT 182.250 5.210 184.280 6.770 ;
    END
  END LADATAOUT10
  PIN LADATAOUT11
    PORT
      LAYER met2 ;
        RECT 186.310 6.780 188.330 301.800 ;
        RECT 186.310 5.220 188.340 6.780 ;
        RECT 186.310 5.210 188.330 5.220 ;
    END
  END LADATAOUT11
  PIN LADATAOUT12
    PORT
      LAYER met2 ;
        RECT 190.400 5.210 192.420 301.800 ;
    END
  END LADATAOUT12
  PIN LADATAOUT13
    PORT
      LAYER met2 ;
        RECT 194.410 6.760 196.430 301.800 ;
        RECT 194.410 5.210 196.440 6.760 ;
        RECT 194.420 5.200 196.440 5.210 ;
    END
  END LADATAOUT13
  PIN LADATAOUT14
    PORT
      LAYER met2 ;
        RECT 198.450 6.770 200.470 301.800 ;
        RECT 198.450 5.210 200.480 6.770 ;
    END
  END LADATAOUT14
  PIN LADATAOUT15
    PORT
      LAYER met2 ;
        RECT 202.540 6.750 204.560 301.800 ;
        RECT 202.540 5.210 204.570 6.750 ;
        RECT 202.550 5.190 204.570 5.210 ;
    END
  END LADATAOUT15
  PIN LADATA16
    PORT
      LAYER met2 ;
        RECT 206.590 5.210 208.610 301.800 ;
    END
  END LADATA16
  PIN LADATAOUT17
    PORT
      LAYER met2 ;
        RECT 210.560 5.210 212.580 301.800 ;
    END
  END LADATAOUT17
  PIN LADATAOUT18
    PORT
      LAYER met2 ;
        RECT 214.680 5.210 216.700 301.800 ;
    END
  END LADATAOUT18
  PIN LADATAOUT19
    PORT
      LAYER met2 ;
        RECT 218.810 5.200 220.830 301.800 ;
    END
  END LADATAOUT19
  PIN LADATAOUT20
    PORT
      LAYER met2 ;
        RECT 222.820 5.210 224.840 301.800 ;
    END
  END LADATAOUT20
  PIN LADATAOUT21
    PORT
      LAYER met2 ;
        RECT 226.830 6.890 228.850 301.800 ;
        RECT 226.830 5.230 228.870 6.890 ;
    END
  END LADATAOUT21
  PIN LADATAOUT22
    PORT
      LAYER met2 ;
        RECT 230.920 6.870 232.940 301.800 ;
        RECT 230.920 5.210 232.950 6.870 ;
    END
  END LADATAOUT22
  PIN LADATAOUT23
    PORT
      LAYER met2 ;
        RECT 235.090 5.210 237.110 301.800 ;
    END
  END LADATAOUT23
  PIN LADATAOUT24
    PORT
      LAYER met2 ;
        RECT 239.090 6.870 241.110 301.800 ;
        RECT 239.090 5.210 241.120 6.870 ;
    END
  END LADATAOUT24
  PIN LADATAIN00
    PORT
      LAYER met2 ;
        RECT 243.100 6.870 245.120 301.800 ;
        RECT 243.070 5.210 245.120 6.870 ;
    END
  END LADATAIN00
  PIN LADATAIN01
    PORT
      LAYER met2 ;
        RECT 247.060 6.870 249.080 301.800 ;
        RECT 247.050 5.210 249.080 6.870 ;
    END
  END LADATAIN01
  PIN LADATAIN02
    PORT
      LAYER met2 ;
        RECT 251.110 6.870 253.130 301.800 ;
        RECT 251.110 5.210 253.150 6.870 ;
    END
  END LADATAIN02
  PIN LADATAIN03
    PORT
      LAYER met2 ;
        RECT 255.170 6.870 257.190 301.800 ;
        RECT 255.170 5.210 257.210 6.870 ;
    END
  END LADATAIN03
  PIN VCCA
    ANTENNADIFFAREA 0.272000 ;
    PORT
      LAYER nwell ;
        RECT 203.610 341.920 206.170 343.830 ;
      LAYER met2 ;
        RECT 243.440 356.810 266.770 357.240 ;
        RECT 203.990 342.370 204.310 342.420 ;
        RECT 199.210 342.210 204.310 342.370 ;
        RECT 203.990 342.160 204.310 342.210 ;
        RECT 203.470 341.440 203.790 341.490 ;
        RECT 199.210 341.280 203.790 341.440 ;
        RECT 203.470 341.230 203.790 341.280 ;
        RECT 203.000 339.600 203.320 339.650 ;
        RECT 199.210 339.440 203.320 339.600 ;
        RECT 203.000 339.390 203.320 339.440 ;
        RECT 202.500 338.670 202.820 338.720 ;
        RECT 199.210 338.510 202.820 338.670 ;
        RECT 202.500 338.460 202.820 338.510 ;
        RECT 203.970 332.750 260.510 333.250 ;
        RECT 254.410 332.350 256.420 332.370 ;
        RECT 203.430 331.850 256.420 332.350 ;
        RECT 202.960 331.430 252.230 331.450 ;
        RECT 202.960 330.950 252.340 331.430 ;
        RECT 250.330 330.890 252.340 330.950 ;
        RECT 254.410 330.890 256.420 331.850 ;
        RECT 258.500 330.890 260.510 332.750 ;
        RECT 243.260 330.550 333.310 330.890 ;
        RECT 202.480 330.050 333.310 330.550 ;
        RECT 243.260 328.800 333.310 330.050 ;
        RECT 246.470 327.580 248.480 328.800 ;
        RECT 250.330 327.580 252.340 328.800 ;
        RECT 254.410 327.580 256.420 328.800 ;
        RECT 258.500 327.580 260.510 328.800 ;
        RECT 264.230 327.580 268.760 327.660 ;
        RECT 243.540 326.430 268.830 327.580 ;
        RECT 246.470 325.380 248.480 326.430 ;
        RECT 250.330 325.380 252.340 326.430 ;
        RECT 254.410 325.380 256.420 326.430 ;
        RECT 258.500 325.380 260.510 326.430 ;
        RECT 264.230 326.410 268.760 326.430 ;
        RECT 243.580 323.290 329.070 325.380 ;
        RECT 246.470 312.750 248.480 323.290 ;
        RECT 246.410 312.230 248.480 312.750 ;
        RECT 250.330 312.750 252.340 323.290 ;
        RECT 246.410 312.100 248.440 312.230 ;
        RECT 250.330 312.100 252.400 312.750 ;
        RECT 254.410 312.730 256.420 323.290 ;
        RECT 258.500 312.750 260.510 323.290 ;
        RECT 250.330 312.060 252.340 312.100 ;
        RECT 254.410 312.080 256.450 312.730 ;
        RECT 258.470 312.170 260.510 312.750 ;
        RECT 258.470 312.100 260.500 312.170 ;
        RECT 254.410 312.000 256.420 312.080 ;
        RECT 326.980 191.860 329.070 323.290 ;
        RECT 331.220 218.330 333.310 328.800 ;
        RECT 331.050 214.620 333.480 218.330 ;
        RECT 326.990 189.960 329.070 191.860 ;
        RECT 326.990 189.840 329.080 189.960 ;
        RECT 326.880 189.780 329.080 189.840 ;
        RECT 326.620 186.100 329.150 189.780 ;
        RECT 326.880 186.080 328.970 186.100 ;
        RECT 263.390 164.230 267.990 165.010 ;
        RECT 263.390 162.550 362.540 164.230 ;
        RECT 263.390 161.260 362.670 162.550 ;
        RECT 263.390 160.440 267.990 161.260 ;
    END
  END VCCA
  OBS
      LAYER nwell ;
        RECT 125.380 382.570 135.070 387.170 ;
        RECT 137.720 382.790 140.430 382.830 ;
        RECT 124.780 381.180 135.070 382.570 ;
        RECT 137.710 381.140 140.430 382.790 ;
        RECT 142.910 381.090 145.130 382.780 ;
        RECT 172.000 381.200 184.050 387.140 ;
        RECT 200.590 381.200 212.640 387.140 ;
        RECT 229.180 381.200 241.230 387.140 ;
        RECT 255.360 382.260 257.090 382.600 ;
        RECT 210.480 380.700 212.230 381.200 ;
        RECT 137.720 379.800 140.430 379.840 ;
        RECT 137.710 379.530 140.430 379.800 ;
        RECT 125.330 375.500 128.070 379.000 ;
        RECT 137.000 377.890 141.000 379.530 ;
        RECT 210.500 379.070 212.230 380.700 ;
        RECT 255.340 380.700 257.090 382.260 ;
        RECT 257.770 381.200 269.820 387.140 ;
        RECT 286.360 381.200 298.410 387.140 ;
        RECT 314.950 381.200 327.000 387.140 ;
        RECT 343.540 381.200 355.590 387.140 ;
        RECT 255.340 379.070 257.070 380.700 ;
        RECT 137.710 377.140 140.430 377.890 ;
        RECT 142.210 377.380 143.820 378.170 ;
        RECT 144.320 377.380 144.830 377.550 ;
        RECT 144.870 377.380 146.020 377.550 ;
        RECT 137.000 373.540 141.000 376.730 ;
        RECT 142.210 376.200 146.210 377.380 ;
        RECT 142.210 376.190 143.000 376.200 ;
        RECT 144.320 376.190 146.210 376.200 ;
        RECT 143.000 376.000 143.270 376.180 ;
        RECT 144.320 375.990 144.830 376.190 ;
        RECT 144.870 376.000 146.020 376.190 ;
        RECT 210.440 375.900 213.750 379.070 ;
        RECT 253.820 378.680 257.130 379.070 ;
        RECT 230.290 378.640 233.000 378.680 ;
        RECT 253.820 378.640 257.370 378.680 ;
        RECT 230.290 376.990 233.010 378.640 ;
        RECT 249.060 378.590 252.370 378.600 ;
        RECT 251.410 378.560 251.600 378.590 ;
        RECT 253.820 376.990 257.380 378.640 ;
        RECT 210.730 375.250 212.480 375.900 ;
        RECT 149.930 374.680 150.150 374.790 ;
        RECT 210.440 373.040 213.750 375.250 ;
        RECT 225.580 374.310 226.140 376.370 ;
        RECT 225.440 374.300 228.750 374.310 ;
        RECT 225.580 373.950 226.140 374.300 ;
        RECT 168.990 372.050 170.760 372.120 ;
        RECT 171.770 370.950 173.540 372.540 ;
        RECT 168.990 370.300 170.760 370.460 ;
        RECT 171.770 369.200 173.540 370.790 ;
        RECT 174.630 370.640 177.130 372.120 ;
        RECT 210.440 370.960 214.000 373.040 ;
        RECT 225.960 372.560 226.380 372.630 ;
        RECT 230.290 372.410 233.010 374.060 ;
        RECT 241.430 373.950 241.990 376.370 ;
        RECT 249.320 376.230 251.050 376.570 ;
        RECT 249.300 374.670 251.050 376.230 ;
        RECT 253.820 375.900 257.130 376.990 ;
        RECT 254.240 375.250 255.520 375.900 ;
        RECT 249.300 374.310 251.030 374.670 ;
        RECT 248.410 374.300 251.030 374.310 ;
        RECT 247.910 373.990 248.230 374.290 ;
        RECT 249.300 373.040 251.030 374.300 ;
        RECT 252.260 374.130 253.540 374.310 ;
        RECT 253.820 374.060 257.130 375.250 ;
        RECT 247.780 372.650 251.090 373.040 ;
        RECT 247.780 372.610 251.330 372.650 ;
        RECT 243.020 372.560 246.330 372.570 ;
        RECT 245.370 372.530 245.560 372.560 ;
        RECT 230.290 372.370 233.000 372.410 ;
        RECT 174.630 370.440 177.160 370.640 ;
        RECT 168.990 368.550 170.760 368.710 ;
        RECT 171.770 367.450 173.540 369.040 ;
        RECT 168.990 366.800 170.760 366.960 ;
        RECT 146.740 363.250 148.770 366.220 ;
        RECT 171.770 365.700 173.540 367.290 ;
        RECT 168.990 365.120 170.760 365.210 ;
        RECT 174.630 365.120 177.130 370.440 ;
        RECT 210.690 369.870 214.000 370.960 ;
        RECT 247.780 370.960 251.340 372.610 ;
        RECT 253.820 372.410 257.380 374.060 ;
        RECT 253.820 372.370 257.370 372.410 ;
        RECT 253.820 372.080 257.130 372.370 ;
        RECT 210.690 368.030 214.000 369.220 ;
        RECT 219.410 368.270 221.390 368.280 ;
        RECT 210.440 366.380 214.000 368.030 ;
        RECT 225.830 367.920 226.390 370.340 ;
        RECT 235.390 367.920 235.950 370.340 ;
        RECT 247.780 369.870 251.090 370.960 ;
        RECT 240.920 369.180 242.060 369.770 ;
        RECT 248.200 369.220 249.480 369.870 ;
        RECT 240.430 368.340 242.060 369.180 ;
        RECT 242.370 368.270 243.840 368.280 ;
        RECT 246.220 368.100 247.500 368.280 ;
        RECT 219.410 367.600 219.480 367.780 ;
        RECT 238.630 367.320 241.390 368.090 ;
        RECT 247.780 368.030 251.090 369.220 ;
        RECT 254.240 368.750 255.520 371.590 ;
        RECT 252.260 368.260 253.540 368.450 ;
        RECT 236.000 366.910 236.010 367.290 ;
        RECT 238.630 367.150 240.620 367.320 ;
        RECT 238.630 366.530 240.610 367.150 ;
        RECT 247.780 366.770 251.340 368.030 ;
        RECT 247.070 366.700 251.340 366.770 ;
        RECT 240.920 366.530 242.060 366.570 ;
        RECT 238.630 366.480 242.060 366.530 ;
        RECT 210.450 366.340 214.000 366.380 ;
        RECT 210.690 366.050 214.000 366.340 ;
        RECT 240.920 365.980 242.060 366.480 ;
        RECT 247.780 366.380 251.340 366.700 ;
        RECT 247.780 366.340 251.330 366.380 ;
        RECT 247.780 366.050 251.090 366.340 ;
        RECT 240.430 365.970 242.060 365.980 ;
        RECT 238.630 365.140 242.060 365.970 ;
        RECT 238.630 365.130 240.620 365.140 ;
        RECT 238.630 364.120 241.390 365.130 ;
        RECT 238.630 364.110 240.620 364.120 ;
        RECT 184.270 363.650 184.300 363.660 ;
        RECT 169.510 363.510 171.280 363.620 ;
        RECT 175.150 363.510 177.650 363.620 ;
        RECT 183.590 363.350 184.300 363.650 ;
        RECT 183.590 363.310 184.270 363.350 ;
        RECT 147.560 363.140 148.100 363.250 ;
        RECT 147.380 362.690 148.100 363.140 ;
        RECT 145.530 362.510 148.100 362.690 ;
        RECT 168.990 361.920 170.760 362.010 ;
        RECT 168.990 360.170 170.760 360.330 ;
        RECT 171.770 359.840 173.540 361.430 ;
        RECT 168.990 358.420 170.760 358.580 ;
        RECT 171.770 358.090 173.540 359.680 ;
        RECT 168.990 356.670 170.760 356.830 ;
        RECT 171.770 356.340 173.540 357.930 ;
        RECT 174.630 356.690 177.130 362.010 ;
        RECT 183.580 357.260 184.280 363.310 ;
        RECT 238.630 363.280 242.060 364.110 ;
        RECT 240.430 363.270 242.060 363.280 ;
        RECT 188.350 361.960 191.770 363.190 ;
        RECT 219.410 362.730 219.490 362.910 ;
        RECT 240.920 362.770 242.060 363.270 ;
        RECT 238.630 362.720 242.060 362.770 ;
        RECT 248.200 362.720 249.480 365.560 ;
        RECT 194.050 361.960 194.060 362.410 ;
        RECT 238.630 362.100 240.610 362.720 ;
        RECT 240.920 362.680 242.060 362.720 ;
        RECT 246.220 362.230 247.500 362.420 ;
        RECT 250.700 362.330 252.560 365.320 ;
        RECT 188.350 361.940 194.090 361.960 ;
        RECT 188.350 360.700 191.770 361.940 ;
        RECT 194.050 361.220 194.060 361.940 ;
        RECT 238.630 361.930 240.620 362.100 ;
        RECT 199.730 361.610 201.460 361.660 ;
        RECT 235.720 361.610 237.450 361.660 ;
        RECT 194.050 361.170 194.100 361.220 ;
        RECT 194.050 361.070 194.110 361.170 ;
        RECT 188.350 358.750 191.770 359.990 ;
        RECT 194.060 359.950 194.110 361.070 ;
        RECT 188.350 358.740 194.090 358.750 ;
        RECT 188.350 357.500 191.770 358.740 ;
        RECT 195.730 358.080 197.460 359.920 ;
        RECT 183.590 357.060 184.280 357.260 ;
        RECT 174.630 356.490 177.160 356.690 ;
        RECT 168.990 355.010 170.760 355.080 ;
        RECT 171.770 354.590 173.540 356.180 ;
        RECT 174.630 355.010 177.130 356.490 ;
        RECT 199.730 355.170 202.650 361.610 ;
        RECT 207.480 360.160 208.040 360.700 ;
        RECT 203.010 356.170 205.570 358.080 ;
        RECT 215.900 356.330 215.970 356.510 ;
        RECT 221.210 356.330 221.280 356.510 ;
        RECT 231.610 356.170 234.170 358.080 ;
        RECT 210.550 355.920 211.660 356.150 ;
        RECT 214.810 355.980 215.400 356.090 ;
        RECT 221.780 355.980 222.370 356.090 ;
        RECT 225.520 355.920 226.630 356.150 ;
        RECT 200.420 355.120 202.650 355.170 ;
        RECT 203.010 352.930 205.570 355.900 ;
        RECT 206.670 354.490 207.020 354.500 ;
        RECT 206.670 354.330 206.680 354.490 ;
        RECT 206.850 354.330 207.020 354.490 ;
        RECT 230.160 354.490 230.510 354.500 ;
        RECT 230.160 354.330 230.330 354.490 ;
        RECT 230.500 354.330 230.510 354.490 ;
        RECT 200.330 352.770 202.060 352.830 ;
        RECT 168.990 351.790 170.760 351.880 ;
        RECT 168.990 350.040 170.760 350.200 ;
        RECT 171.770 349.710 173.540 351.300 ;
        RECT 168.990 348.290 170.760 348.450 ;
        RECT 171.770 347.960 173.540 349.550 ;
        RECT 168.990 346.540 170.760 346.700 ;
        RECT 171.770 346.210 173.540 347.800 ;
        RECT 174.630 346.560 177.130 351.880 ;
        RECT 188.330 351.490 191.750 352.720 ;
        RECT 200.330 352.670 203.250 352.770 ;
        RECT 210.550 352.680 211.660 352.950 ;
        RECT 214.810 352.700 215.400 352.890 ;
        RECT 221.780 352.700 222.370 352.890 ;
        RECT 225.520 352.680 226.630 352.950 ;
        RECT 228.370 352.810 228.460 353.110 ;
        RECT 231.610 352.930 234.170 355.900 ;
        RECT 234.530 355.170 237.450 361.610 ;
        RECT 238.630 361.160 241.390 361.930 ;
        RECT 240.430 360.740 242.060 360.910 ;
        RECT 242.370 360.800 242.820 361.030 ;
        RECT 240.430 360.670 242.890 360.740 ;
        RECT 240.430 360.070 242.060 360.670 ;
        RECT 240.920 359.920 242.060 360.070 ;
        RECT 239.720 359.480 242.060 359.920 ;
        RECT 239.720 358.080 241.450 359.480 ;
        RECT 244.660 356.300 246.520 359.290 ;
        RECT 250.700 359.280 252.560 362.270 ;
        RECT 234.530 355.120 236.760 355.170 ;
        RECT 244.660 353.250 246.520 356.240 ;
        RECT 188.330 351.470 194.070 351.490 ;
        RECT 188.330 350.230 191.750 351.470 ;
        RECT 188.330 348.280 191.750 349.520 ;
        RECT 196.330 349.200 198.060 351.040 ;
        RECT 200.330 350.760 205.570 352.670 ;
        RECT 231.610 350.760 234.170 352.670 ;
        RECT 188.330 348.270 194.070 348.280 ;
        RECT 188.330 347.030 191.750 348.270 ;
        RECT 174.630 346.360 177.160 346.560 ;
        RECT 168.990 344.880 170.760 344.950 ;
        RECT 171.770 344.460 173.540 346.050 ;
        RECT 174.630 344.880 177.130 346.360 ;
        RECT 200.330 346.330 203.250 350.760 ;
        RECT 208.530 350.630 208.660 350.690 ;
        RECT 208.530 350.510 208.600 350.630 ;
        RECT 203.610 347.330 206.170 349.240 ;
        RECT 201.020 346.280 203.250 346.330 ;
        RECT 203.610 344.090 206.170 347.080 ;
        RECT 211.150 347.040 212.260 347.310 ;
        RECT 215.410 347.100 216.000 347.260 ;
        RECT 208.970 346.120 209.060 346.200 ;
        RECT 207.450 345.620 207.620 345.680 ;
        RECT 207.270 345.610 207.620 345.620 ;
        RECT 207.270 345.510 207.280 345.610 ;
        RECT 207.450 345.510 207.620 345.610 ;
        RECT 208.740 344.140 211.700 344.150 ;
        RECT 208.740 343.990 209.150 344.140 ;
        RECT 214.430 344.050 214.810 344.150 ;
        RECT 208.740 343.980 209.330 343.990 ;
        RECT 168.950 342.730 170.720 342.820 ;
        RECT 168.950 340.980 170.720 341.140 ;
        RECT 171.730 340.650 173.500 342.240 ;
        RECT 148.810 337.100 151.180 339.970 ;
        RECT 152.650 338.020 153.210 339.990 ;
        RECT 168.950 339.230 170.720 339.390 ;
        RECT 171.730 338.900 173.500 340.490 ;
        RECT 168.950 337.480 170.720 337.640 ;
        RECT 171.730 337.150 173.500 338.740 ;
        RECT 174.590 337.500 177.090 342.820 ;
        RECT 183.580 337.540 185.330 343.510 ;
        RECT 188.360 342.220 191.780 343.450 ;
        RECT 208.740 342.220 209.150 343.980 ;
        RECT 211.150 343.840 212.260 344.030 ;
        RECT 218.460 344.010 218.860 344.150 ;
        RECT 215.410 343.860 216.000 344.010 ;
        RECT 188.360 342.200 194.100 342.220 ;
        RECT 188.360 340.960 191.780 342.200 ;
        RECT 208.630 341.800 209.150 342.220 ;
        RECT 208.630 341.600 209.140 341.800 ;
        RECT 208.630 341.070 209.150 341.600 ;
        RECT 188.360 339.010 191.780 340.250 ;
        RECT 188.360 339.000 194.100 339.010 ;
        RECT 188.360 337.760 191.780 339.000 ;
        RECT 208.740 338.110 209.150 341.070 ;
        RECT 183.580 337.510 186.600 337.540 ;
        RECT 174.590 337.300 177.120 337.500 ;
        RECT 185.720 337.350 186.600 337.510 ;
        RECT 168.950 335.820 170.720 335.890 ;
        RECT 171.730 335.400 173.500 336.990 ;
        RECT 174.590 335.820 177.090 337.300 ;
        RECT 185.480 331.980 187.500 336.070 ;
        RECT 185.480 331.950 190.300 331.980 ;
        RECT 177.100 331.860 180.490 331.950 ;
        RECT 182.710 331.890 190.300 331.950 ;
        RECT 192.520 331.890 195.910 331.980 ;
        RECT 182.710 331.860 190.770 331.890 ;
        RECT 143.560 330.460 144.180 330.550 ;
        RECT 143.560 324.850 147.420 330.460 ;
        RECT 177.100 326.250 180.960 331.860 ;
        RECT 180.340 326.160 180.960 326.250 ;
        RECT 182.240 330.380 190.770 331.860 ;
        RECT 182.240 326.250 186.100 330.380 ;
        RECT 186.910 326.280 190.770 330.380 ;
        RECT 182.240 326.160 182.860 326.250 ;
        RECT 190.150 326.190 190.770 326.280 ;
        RECT 192.050 326.280 195.910 331.890 ;
        RECT 192.050 326.190 192.670 326.280 ;
        RECT 144.030 324.760 147.420 324.850 ;
        RECT 229.180 311.500 230.030 325.980 ;
        RECT 230.140 317.930 235.190 325.980 ;
        RECT 230.140 316.320 232.310 317.930 ;
        RECT 232.560 316.380 235.190 317.930 ;
        RECT 233.020 316.320 235.190 316.380 ;
        RECT 230.140 311.500 235.190 316.320 ;
        RECT 238.120 314.260 239.470 329.730 ;
        RECT 238.110 313.790 239.470 314.260 ;
        RECT 230.140 311.490 234.230 311.500 ;
        RECT 229.180 309.880 230.030 311.490 ;
        RECT 230.140 309.880 235.190 311.490 ;
        RECT 384.760 272.340 390.700 284.390 ;
        RECT 384.760 243.750 390.700 255.800 ;
        RECT 384.760 215.160 390.700 227.210 ;
        RECT 384.760 186.570 390.700 198.620 ;
        RECT 384.760 157.980 390.700 170.030 ;
        RECT 384.760 129.390 390.700 141.440 ;
        RECT 384.760 100.800 390.700 112.850 ;
      LAYER li1 ;
        RECT 24.080 457.110 31.610 457.660 ;
        RECT 22.390 444.140 23.870 444.390 ;
        RECT 24.080 444.200 24.590 457.110 ;
        RECT 30.940 457.100 31.610 457.110 ;
        RECT 27.240 456.210 30.700 456.650 ;
        RECT 25.310 456.110 30.700 456.210 ;
        RECT 25.310 456.040 30.590 456.110 ;
        RECT 25.310 445.130 25.480 456.040 ;
        RECT 25.810 455.630 30.040 455.650 ;
        RECT 25.790 445.520 30.120 455.630 ;
        RECT 25.850 445.470 26.020 445.520 ;
        RECT 30.420 445.130 30.590 456.040 ;
        RECT 25.310 444.960 30.590 445.130 ;
        RECT 30.350 444.950 30.590 444.960 ;
        RECT 31.100 444.200 31.610 457.100 ;
        RECT 24.080 443.690 31.610 444.200 ;
        RECT 22.380 437.670 23.840 437.710 ;
        RECT 22.380 437.500 23.850 437.670 ;
        RECT 22.380 437.460 23.840 437.500 ;
        RECT 24.080 431.080 24.590 443.690 ;
        RECT 24.950 442.900 30.930 443.130 ;
        RECT 25.040 431.840 30.690 442.900 ;
        RECT 31.100 433.330 31.610 443.690 ;
        RECT 31.090 433.310 31.610 433.330 ;
        RECT 25.040 431.830 30.750 431.840 ;
        RECT 24.960 431.660 30.750 431.830 ;
        RECT 25.050 431.650 30.750 431.660 ;
        RECT 30.520 431.580 30.690 431.650 ;
        RECT 31.090 431.530 31.620 433.310 ;
        RECT 31.100 431.510 31.620 431.530 ;
        RECT 24.080 430.790 26.520 431.080 ;
        RECT 31.100 431.000 31.610 431.510 ;
        RECT 31.100 430.790 31.630 431.000 ;
        RECT 24.080 430.310 31.630 430.790 ;
        RECT 24.080 430.280 31.440 430.310 ;
        RECT 24.080 428.520 31.610 429.070 ;
        RECT 22.390 415.550 23.870 415.800 ;
        RECT 24.080 415.610 24.590 428.520 ;
        RECT 30.940 428.510 31.610 428.520 ;
        RECT 27.240 427.620 30.700 428.060 ;
        RECT 25.310 427.520 30.700 427.620 ;
        RECT 25.310 427.450 30.590 427.520 ;
        RECT 25.310 416.540 25.480 427.450 ;
        RECT 25.810 427.040 30.040 427.060 ;
        RECT 25.790 416.930 30.120 427.040 ;
        RECT 25.850 416.880 26.020 416.930 ;
        RECT 30.420 416.540 30.590 427.450 ;
        RECT 25.310 416.370 30.590 416.540 ;
        RECT 30.350 416.360 30.590 416.370 ;
        RECT 31.100 415.610 31.610 428.510 ;
        RECT 24.080 415.100 31.610 415.610 ;
        RECT 22.380 409.080 23.840 409.120 ;
        RECT 22.380 408.910 23.850 409.080 ;
        RECT 22.380 408.870 23.840 408.910 ;
        RECT 24.080 402.490 24.590 415.100 ;
        RECT 24.950 414.310 30.930 414.540 ;
        RECT 25.040 403.250 30.690 414.310 ;
        RECT 31.100 404.740 31.610 415.100 ;
        RECT 31.090 404.720 31.610 404.740 ;
        RECT 25.040 403.240 30.750 403.250 ;
        RECT 24.960 403.070 30.750 403.240 ;
        RECT 25.050 403.060 30.750 403.070 ;
        RECT 30.520 402.990 30.690 403.060 ;
        RECT 31.090 402.940 31.620 404.720 ;
        RECT 31.100 402.920 31.620 402.940 ;
        RECT 24.080 402.200 26.520 402.490 ;
        RECT 31.100 402.410 31.610 402.920 ;
        RECT 31.100 402.200 31.630 402.410 ;
        RECT 24.080 401.720 31.630 402.200 ;
        RECT 24.080 401.690 31.440 401.720 ;
        RECT 24.080 399.930 31.610 400.480 ;
        RECT 23.660 388.220 23.910 389.680 ;
        RECT 23.700 388.210 23.870 388.220 ;
        RECT 24.080 387.980 24.590 399.930 ;
        RECT 30.940 399.920 31.610 399.930 ;
        RECT 27.240 399.030 30.700 399.470 ;
        RECT 25.310 398.930 30.700 399.030 ;
        RECT 25.310 398.860 30.590 398.930 ;
        RECT 25.310 387.980 25.480 398.860 ;
        RECT 25.810 398.450 30.040 398.470 ;
        RECT 25.790 388.340 30.120 398.450 ;
        RECT 30.420 389.670 30.590 398.860 ;
        RECT 25.850 388.290 26.020 388.340 ;
        RECT 30.340 388.190 30.590 389.670 ;
        RECT 30.420 387.980 30.590 388.190 ;
        RECT 31.100 387.980 31.610 399.920 ;
        RECT 52.250 388.220 52.500 389.680 ;
        RECT 52.290 388.210 52.460 388.220 ;
        RECT 58.930 388.190 59.180 389.670 ;
        RECT 80.840 388.220 81.090 389.680 ;
        RECT 80.880 388.210 81.050 388.220 ;
        RECT 87.520 388.190 87.770 389.670 ;
        RECT 164.860 388.220 165.110 389.680 ;
        RECT 164.900 388.210 165.070 388.220 ;
        RECT 171.540 388.190 171.790 389.670 ;
        RECT 193.450 388.220 193.700 389.680 ;
        RECT 193.490 388.210 193.660 388.220 ;
        RECT 200.130 388.190 200.380 389.670 ;
        RECT 222.040 388.220 222.290 389.680 ;
        RECT 222.080 388.210 222.250 388.220 ;
        RECT 228.720 388.190 228.970 389.670 ;
        RECT 250.630 388.220 250.880 389.680 ;
        RECT 250.670 388.210 250.840 388.220 ;
        RECT 257.310 388.190 257.560 389.670 ;
        RECT 279.220 388.220 279.470 389.680 ;
        RECT 279.260 388.210 279.430 388.220 ;
        RECT 285.900 388.190 286.150 389.670 ;
        RECT 307.810 388.220 308.060 389.680 ;
        RECT 307.850 388.210 308.020 388.220 ;
        RECT 314.490 388.190 314.740 389.670 ;
        RECT 336.400 388.220 336.650 389.680 ;
        RECT 336.440 388.210 336.610 388.220 ;
        RECT 343.080 388.190 343.330 389.670 ;
        RECT 16.480 387.470 43.860 387.980 ;
        RECT 16.480 385.540 17.280 387.470 ;
        RECT 17.860 387.020 18.030 387.100 ;
        RECT 22.390 387.020 23.870 387.210 ;
        RECT 24.080 387.020 24.590 387.470 ;
        RECT 29.100 387.020 29.330 387.110 ;
        RECT 29.890 387.020 30.400 387.470 ;
        RECT 31.100 387.020 31.610 387.470 ;
        RECT 17.860 387.010 31.610 387.020 ;
        RECT 17.850 386.750 31.610 387.010 ;
        RECT 17.850 386.580 42.410 386.750 ;
        RECT 17.850 386.510 31.610 386.580 ;
        RECT 17.850 385.950 29.330 386.510 ;
        RECT 29.890 385.950 30.400 386.510 ;
        RECT 17.850 385.720 30.930 385.950 ;
        RECT 16.480 380.960 16.990 385.540 ;
        RECT 17.850 381.540 30.690 385.720 ;
        RECT 17.780 381.370 30.690 381.540 ;
        RECT 17.850 381.310 18.040 381.370 ;
        RECT 17.730 380.960 19.530 380.970 ;
        RECT 24.080 380.960 24.590 381.370 ;
        RECT 25.040 380.960 30.690 381.370 ;
        RECT 31.100 381.640 31.610 386.510 ;
        RECT 31.720 386.250 41.830 386.270 ;
        RECT 31.720 386.210 41.850 386.250 ;
        RECT 31.670 386.040 41.850 386.210 ;
        RECT 31.720 382.020 41.850 386.040 ;
        RECT 42.240 384.820 42.410 386.580 ;
        RECT 31.720 381.940 41.830 382.020 ;
        RECT 42.240 381.640 42.850 384.820 ;
        RECT 31.100 381.470 42.850 381.640 ;
        RECT 31.100 380.960 31.610 381.470 ;
        RECT 42.310 381.360 42.850 381.470 ;
        RECT 43.310 381.120 43.860 387.470 ;
        RECT 43.300 380.960 43.860 381.120 ;
        RECT 16.480 380.620 43.860 380.960 ;
        RECT 45.070 387.470 72.450 387.980 ;
        RECT 45.070 385.540 45.870 387.470 ;
        RECT 46.450 387.020 46.620 387.100 ;
        RECT 57.690 387.020 57.920 387.110 ;
        RECT 46.450 387.010 57.920 387.020 ;
        RECT 45.070 380.960 45.580 385.540 ;
        RECT 46.440 381.540 57.920 387.010 ;
        RECT 46.370 381.370 57.920 381.540 ;
        RECT 46.440 381.310 46.630 381.370 ;
        RECT 57.690 381.130 57.920 381.370 ;
        RECT 46.320 380.960 48.120 380.970 ;
        RECT 58.480 380.960 58.990 387.470 ;
        RECT 59.750 386.580 71.000 386.750 ;
        RECT 59.750 381.710 59.920 386.580 ;
        RECT 60.310 386.250 70.420 386.270 ;
        RECT 60.310 386.210 70.440 386.250 ;
        RECT 60.260 386.040 70.440 386.210 ;
        RECT 60.310 382.020 70.440 386.040 ;
        RECT 70.830 384.820 71.000 386.580 ;
        RECT 60.310 381.940 70.420 382.020 ;
        RECT 59.740 381.640 59.920 381.710 ;
        RECT 70.830 381.640 71.440 384.820 ;
        RECT 59.740 381.470 71.440 381.640 ;
        RECT 70.900 381.360 71.440 381.470 ;
        RECT 71.900 381.120 72.450 387.470 ;
        RECT 71.890 380.960 72.450 381.120 ;
        RECT 45.070 380.620 72.450 380.960 ;
        RECT 73.660 387.470 101.040 387.980 ;
        RECT 73.660 385.540 74.460 387.470 ;
        RECT 75.040 387.020 75.210 387.100 ;
        RECT 86.280 387.020 86.510 387.110 ;
        RECT 75.040 387.010 86.510 387.020 ;
        RECT 73.660 380.960 74.170 385.540 ;
        RECT 75.030 381.540 86.510 387.010 ;
        RECT 74.960 381.370 86.510 381.540 ;
        RECT 75.030 381.310 75.220 381.370 ;
        RECT 86.280 381.130 86.510 381.370 ;
        RECT 74.910 380.960 76.710 380.970 ;
        RECT 87.070 380.960 87.580 387.470 ;
        RECT 88.340 386.580 99.590 386.750 ;
        RECT 88.340 381.710 88.510 386.580 ;
        RECT 88.900 386.250 99.010 386.270 ;
        RECT 88.900 386.210 99.030 386.250 ;
        RECT 88.850 386.040 99.030 386.210 ;
        RECT 88.900 382.020 99.030 386.040 ;
        RECT 99.420 384.820 99.590 386.580 ;
        RECT 88.900 381.940 99.010 382.020 ;
        RECT 88.330 381.640 88.510 381.710 ;
        RECT 99.420 381.640 100.030 384.820 ;
        RECT 88.330 381.470 100.030 381.640 ;
        RECT 99.490 381.360 100.030 381.470 ;
        RECT 100.490 381.120 101.040 387.470 ;
        RECT 142.840 386.690 143.060 387.810 ;
        RECT 142.790 386.500 143.120 386.690 ;
        RECT 149.580 386.500 149.820 387.850 ;
        RECT 157.680 387.470 185.060 387.980 ;
        RECT 157.680 386.300 158.480 387.470 ;
        RECT 159.060 387.020 159.230 387.100 ;
        RECT 170.300 387.020 170.530 387.110 ;
        RECT 159.060 387.010 170.530 387.020 ;
        RECT 159.050 386.300 170.530 387.010 ;
        RECT 171.090 386.300 171.600 387.470 ;
        RECT 172.360 386.580 183.610 386.750 ;
        RECT 172.360 386.300 172.530 386.580 ;
        RECT 100.480 380.960 101.040 381.120 ;
        RECT 73.660 380.620 101.040 380.960 ;
        RECT 16.510 380.450 43.860 380.620 ;
        RECT 45.100 380.450 72.450 380.620 ;
        RECT 73.690 380.450 101.040 380.620 ;
        RECT 122.080 386.270 176.820 386.300 ;
        RECT 122.080 386.250 183.030 386.270 ;
        RECT 122.080 386.030 183.050 386.250 ;
        RECT 122.080 385.900 146.420 386.030 ;
        RECT 155.110 385.900 183.050 386.030 ;
        RECT 16.510 380.430 17.200 380.450 ;
        RECT 17.710 380.440 19.510 380.450 ;
        RECT 22.380 380.320 23.850 380.450 ;
        RECT 22.380 380.280 23.840 380.320 ;
        RECT 24.080 373.900 24.590 380.450 ;
        RECT 25.040 374.660 30.690 380.450 ;
        RECT 31.100 376.150 31.610 380.450 ;
        RECT 45.100 380.430 45.790 380.450 ;
        RECT 46.300 380.440 48.100 380.450 ;
        RECT 73.690 380.430 74.380 380.450 ;
        RECT 74.890 380.440 76.690 380.450 ;
        RECT 122.080 378.300 122.250 385.900 ;
        RECT 157.680 385.540 158.480 385.900 ;
        RECT 125.240 381.480 125.410 382.150 ;
        RECT 139.900 381.660 140.130 382.350 ;
        RECT 144.600 381.610 144.830 382.300 ;
        RECT 157.680 380.960 158.190 385.540 ;
        RECT 159.050 381.540 170.530 385.900 ;
        RECT 158.980 381.370 170.530 381.540 ;
        RECT 159.050 381.310 159.240 381.370 ;
        RECT 170.300 381.130 170.530 381.370 ;
        RECT 158.930 380.960 160.730 380.970 ;
        RECT 171.090 380.960 171.600 385.900 ;
        RECT 172.360 381.710 172.530 385.900 ;
        RECT 172.920 382.020 183.050 385.900 ;
        RECT 183.440 384.820 183.610 386.580 ;
        RECT 172.920 381.940 183.030 382.020 ;
        RECT 172.350 381.640 172.530 381.710 ;
        RECT 176.650 381.640 176.820 381.940 ;
        RECT 183.440 381.640 184.050 384.820 ;
        RECT 172.350 381.470 184.050 381.640 ;
        RECT 176.650 380.960 176.820 381.470 ;
        RECT 183.510 381.360 184.050 381.470 ;
        RECT 184.510 381.120 185.060 387.470 ;
        RECT 184.500 380.960 185.060 381.120 ;
        RECT 157.680 380.620 185.060 380.960 ;
        RECT 186.270 387.470 213.650 387.980 ;
        RECT 186.270 385.540 187.070 387.470 ;
        RECT 187.650 387.020 187.820 387.100 ;
        RECT 198.890 387.020 199.120 387.110 ;
        RECT 187.650 387.010 199.120 387.020 ;
        RECT 186.270 380.960 186.780 385.540 ;
        RECT 187.640 381.540 199.120 387.010 ;
        RECT 187.570 381.370 199.120 381.540 ;
        RECT 187.640 381.310 187.830 381.370 ;
        RECT 198.890 381.130 199.120 381.370 ;
        RECT 187.520 380.960 189.320 380.970 ;
        RECT 199.680 380.960 200.190 387.470 ;
        RECT 200.950 386.580 212.200 386.750 ;
        RECT 200.950 381.710 201.120 386.580 ;
        RECT 201.510 386.250 211.620 386.270 ;
        RECT 201.510 386.210 211.640 386.250 ;
        RECT 201.460 386.040 211.640 386.210 ;
        RECT 201.510 382.020 211.640 386.040 ;
        RECT 212.030 384.820 212.200 386.580 ;
        RECT 201.510 381.940 211.620 382.020 ;
        RECT 200.940 381.640 201.120 381.710 ;
        RECT 212.030 381.640 212.640 384.820 ;
        RECT 200.940 381.470 212.640 381.640 ;
        RECT 212.100 381.360 212.640 381.470 ;
        RECT 211.260 380.960 211.810 381.300 ;
        RECT 213.100 381.120 213.650 387.470 ;
        RECT 213.090 380.960 213.650 381.120 ;
        RECT 186.270 380.620 213.650 380.960 ;
        RECT 214.860 387.470 242.240 387.980 ;
        RECT 214.860 385.540 215.660 387.470 ;
        RECT 216.240 387.020 216.410 387.100 ;
        RECT 227.480 387.020 227.710 387.110 ;
        RECT 216.240 387.010 227.710 387.020 ;
        RECT 214.860 380.960 215.370 385.540 ;
        RECT 216.230 381.540 227.710 387.010 ;
        RECT 216.160 381.370 227.710 381.540 ;
        RECT 216.230 381.310 216.420 381.370 ;
        RECT 227.480 381.130 227.710 381.370 ;
        RECT 216.110 380.960 217.910 380.970 ;
        RECT 228.270 380.960 228.780 387.470 ;
        RECT 229.540 386.580 240.790 386.750 ;
        RECT 229.540 381.710 229.710 386.580 ;
        RECT 230.100 386.250 240.210 386.270 ;
        RECT 230.100 386.210 240.230 386.250 ;
        RECT 230.050 386.040 240.230 386.210 ;
        RECT 230.100 382.020 240.230 386.040 ;
        RECT 240.620 384.820 240.790 386.580 ;
        RECT 230.100 381.940 240.210 382.020 ;
        RECT 229.530 381.640 229.710 381.710 ;
        RECT 240.620 381.640 241.230 384.820 ;
        RECT 229.530 381.470 241.230 381.640 ;
        RECT 240.690 381.360 241.230 381.470 ;
        RECT 241.690 381.120 242.240 387.470 ;
        RECT 241.680 380.960 242.240 381.120 ;
        RECT 214.860 380.620 242.240 380.960 ;
        RECT 243.450 387.470 270.830 387.980 ;
        RECT 243.450 385.540 244.250 387.470 ;
        RECT 244.830 387.020 245.000 387.100 ;
        RECT 256.070 387.020 256.300 387.110 ;
        RECT 244.830 387.010 256.300 387.020 ;
        RECT 243.450 380.960 243.960 385.540 ;
        RECT 244.820 381.540 256.300 387.010 ;
        RECT 244.750 381.370 256.300 381.540 ;
        RECT 244.820 381.310 245.010 381.370 ;
        RECT 256.070 381.300 256.300 381.370 ;
        RECT 244.700 380.960 246.500 380.970 ;
        RECT 255.760 380.960 256.310 381.300 ;
        RECT 256.860 380.960 257.370 387.470 ;
        RECT 258.130 386.580 269.380 386.750 ;
        RECT 258.130 381.710 258.300 386.580 ;
        RECT 258.690 386.250 268.800 386.270 ;
        RECT 258.690 386.210 268.820 386.250 ;
        RECT 258.640 386.040 268.820 386.210 ;
        RECT 258.690 382.020 268.820 386.040 ;
        RECT 269.210 384.820 269.380 386.580 ;
        RECT 258.690 381.940 268.800 382.020 ;
        RECT 258.120 381.640 258.300 381.710 ;
        RECT 269.210 381.640 269.820 384.820 ;
        RECT 258.120 381.470 269.820 381.640 ;
        RECT 269.280 381.360 269.820 381.470 ;
        RECT 270.280 381.120 270.830 387.470 ;
        RECT 270.270 380.960 270.830 381.120 ;
        RECT 243.450 380.620 270.830 380.960 ;
        RECT 272.040 387.470 299.420 387.980 ;
        RECT 272.040 385.540 272.840 387.470 ;
        RECT 273.420 387.020 273.590 387.100 ;
        RECT 284.660 387.020 284.890 387.110 ;
        RECT 273.420 387.010 284.890 387.020 ;
        RECT 272.040 380.960 272.550 385.540 ;
        RECT 273.410 381.540 284.890 387.010 ;
        RECT 273.340 381.370 284.890 381.540 ;
        RECT 273.410 381.310 273.600 381.370 ;
        RECT 284.660 381.130 284.890 381.370 ;
        RECT 273.290 380.960 275.090 380.970 ;
        RECT 285.450 380.960 285.960 387.470 ;
        RECT 286.720 386.580 297.970 386.750 ;
        RECT 286.720 381.710 286.890 386.580 ;
        RECT 287.280 386.250 297.390 386.270 ;
        RECT 287.280 386.210 297.410 386.250 ;
        RECT 287.230 386.040 297.410 386.210 ;
        RECT 287.280 382.020 297.410 386.040 ;
        RECT 297.800 384.820 297.970 386.580 ;
        RECT 287.280 381.940 297.390 382.020 ;
        RECT 286.710 381.640 286.890 381.710 ;
        RECT 297.800 381.640 298.410 384.820 ;
        RECT 286.710 381.470 298.410 381.640 ;
        RECT 297.870 381.360 298.410 381.470 ;
        RECT 298.870 381.120 299.420 387.470 ;
        RECT 298.860 380.960 299.420 381.120 ;
        RECT 272.040 380.620 299.420 380.960 ;
        RECT 300.630 387.470 328.010 387.980 ;
        RECT 300.630 385.540 301.430 387.470 ;
        RECT 302.010 387.020 302.180 387.100 ;
        RECT 313.250 387.020 313.480 387.110 ;
        RECT 302.010 387.010 313.480 387.020 ;
        RECT 300.630 380.960 301.140 385.540 ;
        RECT 302.000 381.540 313.480 387.010 ;
        RECT 301.930 381.370 313.480 381.540 ;
        RECT 302.000 381.310 302.190 381.370 ;
        RECT 313.250 381.130 313.480 381.370 ;
        RECT 301.880 380.960 303.680 380.970 ;
        RECT 314.040 380.960 314.550 387.470 ;
        RECT 315.310 386.580 326.560 386.750 ;
        RECT 315.310 381.710 315.480 386.580 ;
        RECT 315.870 386.250 325.980 386.270 ;
        RECT 315.870 386.210 326.000 386.250 ;
        RECT 315.820 386.040 326.000 386.210 ;
        RECT 315.870 382.020 326.000 386.040 ;
        RECT 326.390 384.820 326.560 386.580 ;
        RECT 315.870 381.940 325.980 382.020 ;
        RECT 315.300 381.640 315.480 381.710 ;
        RECT 326.390 381.640 327.000 384.820 ;
        RECT 315.300 381.470 327.000 381.640 ;
        RECT 326.460 381.360 327.000 381.470 ;
        RECT 327.460 381.120 328.010 387.470 ;
        RECT 327.450 380.960 328.010 381.120 ;
        RECT 300.630 380.620 328.010 380.960 ;
        RECT 329.220 387.470 356.600 387.980 ;
        RECT 329.220 385.540 330.020 387.470 ;
        RECT 330.600 387.020 330.770 387.100 ;
        RECT 341.840 387.020 342.070 387.110 ;
        RECT 330.600 387.010 342.070 387.020 ;
        RECT 329.220 380.960 329.730 385.540 ;
        RECT 330.590 381.540 342.070 387.010 ;
        RECT 330.520 381.370 342.070 381.540 ;
        RECT 330.590 381.310 330.780 381.370 ;
        RECT 341.840 381.130 342.070 381.370 ;
        RECT 330.470 380.960 332.270 380.970 ;
        RECT 342.630 380.960 343.140 387.470 ;
        RECT 343.900 386.580 355.150 386.750 ;
        RECT 343.900 381.710 344.070 386.580 ;
        RECT 344.460 386.250 354.570 386.270 ;
        RECT 344.460 386.210 354.590 386.250 ;
        RECT 344.410 386.040 354.590 386.210 ;
        RECT 344.460 382.020 354.590 386.040 ;
        RECT 354.980 384.820 355.150 386.580 ;
        RECT 344.460 381.940 354.570 382.020 ;
        RECT 343.890 381.640 344.070 381.710 ;
        RECT 354.980 381.640 355.590 384.820 ;
        RECT 343.890 381.470 355.590 381.640 ;
        RECT 355.050 381.360 355.590 381.470 ;
        RECT 356.050 381.120 356.600 387.470 ;
        RECT 356.040 380.960 356.600 381.120 ;
        RECT 329.220 380.620 356.600 380.960 ;
        RECT 157.710 380.450 185.060 380.620 ;
        RECT 186.300 380.450 213.650 380.620 ;
        RECT 214.890 380.450 242.240 380.620 ;
        RECT 243.480 380.450 270.830 380.620 ;
        RECT 272.070 380.450 299.420 380.620 ;
        RECT 300.660 380.450 328.010 380.620 ;
        RECT 329.250 380.450 356.600 380.620 ;
        RECT 157.710 380.430 158.400 380.450 ;
        RECT 158.910 380.440 160.710 380.450 ;
        RECT 139.900 379.200 140.130 379.360 ;
        RECT 125.200 378.690 125.370 379.020 ;
        RECT 125.440 378.580 125.530 378.720 ;
        RECT 126.600 378.690 126.770 379.020 ;
        RECT 125.330 378.400 126.330 378.580 ;
        RECT 126.820 378.570 126.900 378.720 ;
        RECT 128.530 378.610 129.200 378.780 ;
        RECT 126.730 378.400 127.740 378.570 ;
        RECT 137.340 378.220 140.650 379.200 ;
        RECT 176.650 378.820 176.820 380.450 ;
        RECT 186.300 380.430 186.990 380.450 ;
        RECT 187.500 380.440 189.300 380.450 ;
        RECT 214.890 380.430 215.580 380.450 ;
        RECT 216.090 380.440 217.890 380.450 ;
        RECT 243.480 380.430 244.170 380.450 ;
        RECT 244.680 380.440 246.480 380.450 ;
        RECT 272.070 380.430 272.760 380.450 ;
        RECT 273.270 380.440 275.070 380.450 ;
        RECT 300.660 380.430 301.350 380.450 ;
        RECT 301.860 380.440 303.660 380.450 ;
        RECT 329.250 380.430 329.940 380.450 ;
        RECT 330.450 380.440 332.250 380.450 ;
        RECT 211.260 379.140 211.810 379.570 ;
        RECT 255.760 379.140 256.310 379.570 ;
        RECT 210.840 378.340 211.040 378.690 ;
        RECT 212.320 378.440 212.850 378.610 ;
        RECT 254.720 378.440 255.250 378.610 ;
        RECT 210.830 378.310 211.040 378.340 ;
        RECT 256.530 378.340 256.730 378.690 ;
        RECT 256.530 378.310 256.740 378.340 ;
        RECT 126.400 377.870 126.720 377.910 ;
        RECT 126.390 377.720 126.720 377.870 ;
        RECT 125.660 377.550 127.740 377.720 ;
        RECT 128.270 377.690 128.940 377.860 ;
        RECT 139.900 377.660 140.130 378.220 ;
        RECT 148.520 377.960 150.880 378.130 ;
        RECT 142.590 377.580 142.760 377.910 ;
        RECT 143.270 377.580 143.440 377.910 ;
        RECT 210.830 377.730 211.050 378.310 ;
        RECT 210.830 377.720 211.040 377.730 ;
        RECT 125.840 377.140 127.660 377.310 ;
        RECT 128.360 377.150 128.570 377.580 ;
        RECT 211.210 377.550 211.400 377.560 ;
        RECT 128.380 377.130 128.550 377.150 ;
        RECT 141.790 377.130 142.110 377.170 ;
        RECT 126.400 377.030 126.720 377.070 ;
        RECT 126.390 376.900 126.720 377.030 ;
        RECT 141.780 376.940 142.110 377.130 ;
        RECT 142.660 377.020 142.830 377.370 ;
        RECT 211.200 377.260 211.400 377.550 ;
        RECT 143.150 377.210 143.470 377.250 ;
        RECT 143.140 377.020 143.470 377.210 ;
        RECT 143.840 377.200 144.160 377.240 ;
        RECT 141.790 376.910 142.110 376.940 ;
        RECT 125.660 376.730 127.740 376.900 ;
        RECT 142.230 376.760 142.830 377.020 ;
        RECT 143.150 376.990 143.470 377.020 ;
        RECT 143.830 377.010 144.160 377.200 ;
        RECT 143.840 376.980 144.160 377.010 ;
        RECT 211.140 376.930 211.410 377.260 ;
        RECT 151.160 376.780 151.330 376.800 ;
        RECT 128.270 376.260 128.940 376.430 ;
        RECT 31.090 376.130 31.610 376.150 ;
        RECT 25.040 374.650 30.750 374.660 ;
        RECT 24.960 374.480 30.750 374.650 ;
        RECT 25.050 374.470 30.750 374.480 ;
        RECT 30.520 374.400 30.690 374.470 ;
        RECT 31.090 374.350 31.620 376.130 ;
        RECT 125.660 375.890 126.330 376.060 ;
        RECT 127.060 375.890 127.740 376.060 ;
        RECT 127.940 375.770 128.130 375.910 ;
        RECT 127.940 375.680 129.210 375.770 ;
        RECT 128.070 375.600 129.210 375.680 ;
        RECT 137.340 375.420 140.650 376.400 ;
        RECT 128.060 375.170 128.230 375.210 ;
        RECT 128.060 375.140 128.440 375.170 ;
        RECT 125.660 374.770 126.330 374.940 ;
        RECT 126.630 374.810 126.800 375.140 ;
        RECT 128.060 374.950 128.450 375.140 ;
        RECT 128.540 374.990 129.210 375.160 ;
        RECT 126.860 374.770 127.740 374.940 ;
        RECT 128.060 374.910 128.440 374.950 ;
        RECT 128.060 374.880 128.230 374.910 ;
        RECT 31.100 374.330 31.620 374.350 ;
        RECT 24.080 373.610 26.520 373.900 ;
        RECT 31.100 373.820 31.610 374.330 ;
        RECT 126.380 374.230 126.700 374.270 ;
        RECT 127.810 374.250 128.130 374.290 ;
        RECT 126.370 374.100 126.700 374.230 ;
        RECT 127.800 374.100 128.130 374.250 ;
        RECT 125.650 373.930 129.230 374.100 ;
        RECT 137.340 373.870 140.650 374.850 ;
        RECT 141.290 373.900 141.460 376.550 ;
        RECT 142.660 376.360 142.830 376.760 ;
        RECT 148.270 376.610 151.330 376.780 ;
        RECT 151.160 375.960 151.330 376.610 ;
        RECT 211.600 376.450 211.770 378.060 ;
        RECT 217.750 378.050 217.940 378.280 ;
        RECT 211.590 376.260 211.770 376.450 ;
        RECT 212.430 376.360 212.600 378.050 ;
        RECT 213.020 377.860 213.350 378.030 ;
        RECT 214.370 377.860 214.720 378.030 ;
        RECT 218.030 378.000 218.910 378.170 ;
        RECT 218.220 377.610 218.410 377.720 ;
        RECT 218.110 377.490 218.410 377.610 ;
        RECT 218.740 377.610 218.910 378.000 ;
        RECT 218.110 377.440 218.330 377.490 ;
        RECT 218.740 377.440 219.130 377.610 ;
        RECT 230.590 377.510 230.820 378.200 ;
        RECT 254.960 377.510 255.190 378.200 ;
        RECT 213.020 377.070 213.350 377.240 ;
        RECT 214.370 377.070 214.720 377.240 ;
        RECT 250.190 377.220 250.510 377.260 ;
        RECT 250.190 377.030 250.520 377.220 ;
        RECT 250.190 377.000 250.510 377.030 ;
        RECT 216.820 376.650 217.140 376.690 ;
        RECT 218.070 376.650 219.150 376.820 ;
        RECT 219.480 376.650 220.560 376.820 ;
        RECT 216.810 376.460 217.140 376.650 ;
        RECT 213.020 376.280 213.350 376.450 ;
        RECT 214.370 376.280 214.710 376.450 ;
        RECT 216.820 376.430 217.140 376.460 ;
        RECT 254.970 376.360 255.140 377.510 ;
        RECT 255.800 376.450 255.970 378.060 ;
        RECT 256.520 377.730 256.740 378.310 ;
        RECT 256.530 377.720 256.740 377.730 ;
        RECT 256.170 377.550 256.360 377.560 ;
        RECT 256.170 377.260 256.370 377.550 ;
        RECT 256.160 376.930 256.450 377.260 ;
        RECT 217.750 376.060 217.940 376.290 ;
        RECT 255.800 376.260 255.980 376.450 ;
        RECT 151.160 375.790 152.430 375.960 ;
        RECT 218.050 375.860 218.130 376.030 ;
        RECT 31.100 373.610 31.630 373.820 ;
        RECT 125.590 373.650 125.910 373.690 ;
        RECT 126.520 373.650 126.840 373.690 ;
        RECT 127.220 373.650 127.540 373.690 ;
        RECT 127.960 373.650 128.280 373.690 ;
        RECT 24.080 373.130 31.630 373.610 ;
        RECT 125.580 373.460 125.910 373.650 ;
        RECT 126.510 373.460 126.840 373.650 ;
        RECT 127.210 373.460 127.540 373.650 ;
        RECT 127.950 373.480 128.280 373.650 ;
        RECT 128.670 373.640 128.990 373.680 ;
        RECT 128.660 373.480 128.990 373.640 ;
        RECT 141.290 373.510 141.470 373.900 ;
        RECT 151.160 373.530 151.330 375.790 ;
        RECT 218.610 375.710 218.820 376.140 ;
        RECT 218.630 375.690 218.800 375.710 ;
        RECT 153.280 374.570 153.450 375.460 ;
        RECT 211.510 374.840 212.060 375.270 ;
        RECT 216.810 374.960 217.130 375.000 ;
        RECT 217.760 374.990 217.950 375.220 ;
        RECT 218.080 375.120 218.130 375.290 ;
        RECT 218.220 375.170 218.410 375.400 ;
        RECT 219.220 375.290 219.390 375.860 ;
        RECT 223.500 375.710 223.690 376.030 ;
        RECT 243.880 375.710 244.070 376.030 ;
        RECT 223.500 375.620 223.780 375.710 ;
        RECT 220.140 375.480 223.780 375.620 ;
        RECT 243.790 375.620 244.070 375.710 ;
        RECT 254.800 375.820 255.130 375.990 ;
        RECT 255.240 375.910 255.570 376.080 ;
        RECT 243.790 375.480 247.430 375.620 ;
        RECT 254.800 375.540 255.160 375.820 ;
        RECT 220.140 375.440 223.690 375.480 ;
        RECT 218.500 375.260 218.550 375.270 ;
        RECT 219.130 375.260 219.210 375.270 ;
        RECT 218.500 375.220 219.210 375.260 ;
        RECT 218.500 375.180 219.230 375.220 ;
        RECT 218.460 375.060 219.300 375.180 ;
        RECT 223.500 375.020 223.690 375.440 ;
        RECT 243.880 375.440 247.430 375.480 ;
        RECT 243.880 375.020 244.070 375.440 ;
        RECT 252.730 375.290 253.050 375.330 ;
        RECT 211.590 374.700 211.770 374.840 ;
        RECT 211.140 373.890 211.410 374.220 ;
        RECT 211.200 373.600 211.400 373.890 ;
        RECT 211.210 373.590 211.400 373.600 ;
        RECT 211.600 373.540 211.770 374.700 ;
        RECT 127.950 373.460 128.990 373.480 ;
        RECT 141.070 373.470 141.470 373.510 ;
        RECT 150.930 373.490 151.330 373.530 ;
        RECT 125.590 373.430 125.910 373.460 ;
        RECT 126.520 373.430 126.840 373.460 ;
        RECT 127.220 373.430 127.540 373.460 ;
        RECT 127.960 373.430 128.990 373.460 ;
        RECT 125.700 373.420 128.990 373.430 ;
        RECT 125.700 373.260 129.130 373.420 ;
        RECT 141.060 373.280 141.470 373.470 ;
        RECT 150.920 373.380 151.330 373.490 ;
        RECT 210.830 373.420 211.040 373.430 ;
        RECT 150.920 373.300 151.250 373.380 ;
        RECT 128.280 373.250 129.130 373.260 ;
        RECT 141.070 373.250 141.470 373.280 ;
        RECT 150.930 373.270 151.250 373.300 ;
        RECT 141.290 373.170 141.470 373.250 ;
        RECT 24.080 373.100 31.440 373.130 ;
        RECT 210.830 372.840 211.050 373.420 ;
        RECT 211.510 373.110 212.060 373.540 ;
        RECT 211.600 373.090 211.770 373.110 ;
        RECT 212.430 373.100 212.600 374.790 ;
        RECT 213.020 374.700 213.350 374.870 ;
        RECT 214.370 374.700 214.710 374.870 ;
        RECT 216.800 374.770 217.130 374.960 ;
        RECT 249.720 374.840 250.270 375.270 ;
        RECT 252.730 375.100 253.060 375.290 ;
        RECT 252.730 375.070 253.050 375.100 ;
        RECT 253.130 375.080 253.330 375.410 ;
        RECT 253.720 375.220 253.920 375.410 ;
        RECT 254.450 375.370 255.160 375.540 ;
        RECT 254.390 375.250 254.710 375.290 ;
        RECT 253.410 374.890 253.600 374.900 ;
        RECT 253.610 374.890 253.960 375.220 ;
        RECT 254.390 375.060 254.720 375.250 ;
        RECT 254.390 375.030 254.710 375.060 ;
        RECT 216.810 374.740 217.130 374.770 ;
        RECT 218.070 374.330 219.150 374.500 ;
        RECT 219.470 374.330 220.710 374.500 ;
        RECT 250.190 374.460 250.510 374.500 ;
        RECT 244.910 374.400 245.140 374.440 ;
        RECT 250.190 374.270 250.520 374.460 ;
        RECT 252.500 374.380 252.670 374.710 ;
        RECT 252.680 374.640 253.000 374.680 ;
        RECT 252.680 374.450 253.010 374.640 ;
        RECT 252.680 374.420 253.000 374.450 ;
        RECT 253.130 374.420 253.330 374.750 ;
        RECT 253.410 374.560 253.960 374.890 ;
        RECT 250.190 374.240 250.510 374.270 ;
        RECT 253.610 374.230 253.960 374.560 ;
        RECT 213.020 373.910 213.350 374.080 ;
        RECT 214.370 373.910 214.720 374.080 ;
        RECT 219.800 374.010 219.970 374.070 ;
        RECT 254.450 374.050 255.150 374.930 ;
        RECT 255.800 374.700 255.980 374.890 ;
        RECT 218.210 373.710 218.400 373.820 ;
        RECT 219.780 373.800 219.990 374.010 ;
        RECT 219.800 373.730 219.970 373.800 ;
        RECT 218.110 373.590 218.400 373.710 ;
        RECT 218.670 373.700 219.130 373.710 ;
        RECT 218.110 373.540 218.320 373.590 ;
        RECT 218.670 373.550 219.140 373.700 ;
        RECT 253.790 373.660 253.980 373.890 ;
        RECT 254.970 373.630 255.140 374.050 ;
        RECT 218.670 373.540 219.130 373.550 ;
        RECT 213.020 373.120 213.350 373.290 ;
        RECT 214.370 373.120 214.720 373.290 ;
        RECT 217.780 373.200 217.970 373.310 ;
        RECT 218.670 373.200 218.860 373.540 ;
        RECT 217.780 373.080 218.860 373.200 ;
        RECT 217.900 373.020 218.860 373.080 ;
        RECT 230.590 372.850 230.820 373.540 ;
        RECT 249.720 373.110 250.270 373.540 ;
        RECT 252.500 373.120 252.670 373.450 ;
        RECT 252.680 373.380 253.000 373.410 ;
        RECT 252.680 373.190 253.010 373.380 ;
        RECT 252.680 373.150 253.000 373.190 ;
        RECT 253.130 373.080 253.330 373.410 ;
        RECT 253.610 373.270 253.960 373.600 ;
        RECT 254.440 373.540 255.140 373.630 ;
        RECT 254.440 373.450 255.190 373.540 ;
        RECT 253.410 372.940 253.960 373.270 ;
        RECT 253.410 372.930 253.600 372.940 ;
        RECT 210.830 372.810 211.040 372.840 ;
        RECT 210.840 372.460 211.040 372.810 ;
        RECT 252.730 372.730 253.050 372.760 ;
        RECT 211.090 372.310 211.290 372.660 ;
        RECT 212.320 372.580 212.850 372.710 ;
        RECT 212.320 372.540 213.100 372.580 ;
        RECT 212.570 372.410 213.100 372.540 ;
        RECT 248.680 372.410 249.210 372.580 ;
        RECT 211.080 372.280 211.290 372.310 ;
        RECT 150.080 372.130 151.600 372.140 ;
        RECT 24.080 371.340 31.610 371.890 ;
        RECT 150.080 371.340 151.630 372.130 ;
        RECT 173.430 372.070 173.780 372.170 ;
        RECT 177.020 372.120 177.190 372.160 ;
        RECT 176.040 372.100 177.190 372.120 ;
        RECT 175.090 372.070 175.550 372.100 ;
        RECT 172.020 371.900 172.780 372.070 ;
        RECT 173.030 371.900 174.200 372.070 ;
        RECT 174.440 371.930 175.550 372.070 ;
        RECT 176.000 371.930 177.190 372.100 ;
        RECT 174.440 371.900 175.260 371.930 ;
        RECT 172.020 371.890 172.250 371.900 ;
        RECT 171.980 371.450 172.250 371.890 ;
        RECT 175.000 371.760 175.260 371.900 ;
        RECT 173.460 371.450 173.790 371.710 ;
        RECT 174.410 371.660 174.700 371.690 ;
        RECT 174.370 371.490 174.700 371.660 ;
        RECT 174.410 371.450 174.700 371.490 ;
        RECT 175.000 371.590 176.180 371.760 ;
        RECT 211.080 371.700 211.300 372.280 ;
        RECT 211.080 371.690 211.290 371.700 ;
        RECT 175.000 371.450 175.260 371.590 ;
        RECT 22.390 358.370 23.870 358.620 ;
        RECT 24.080 358.430 24.590 371.340 ;
        RECT 30.940 371.330 31.610 371.340 ;
        RECT 27.240 370.440 30.700 370.880 ;
        RECT 25.310 370.340 30.700 370.440 ;
        RECT 25.310 370.270 30.590 370.340 ;
        RECT 25.310 359.360 25.480 370.270 ;
        RECT 25.810 369.860 30.040 369.880 ;
        RECT 25.790 359.750 30.120 369.860 ;
        RECT 25.850 359.700 26.020 359.750 ;
        RECT 30.420 359.360 30.590 370.270 ;
        RECT 25.310 359.190 30.590 359.360 ;
        RECT 30.350 359.180 30.590 359.190 ;
        RECT 31.100 358.430 31.610 371.330 ;
        RECT 171.430 371.310 171.600 371.370 ;
        RECT 171.400 371.090 171.620 371.310 ;
        RECT 171.950 371.270 172.280 371.450 ;
        RECT 172.530 371.280 174.690 371.450 ;
        RECT 174.930 371.280 175.260 371.450 ;
        RECT 175.400 371.440 176.180 371.590 ;
        RECT 175.030 371.230 175.260 371.280 ;
        RECT 171.430 371.040 171.600 371.090 ;
        RECT 175.030 371.000 175.200 371.230 ;
        RECT 175.550 371.090 175.760 371.420 ;
        RECT 176.000 371.150 176.180 371.440 ;
        RECT 176.460 371.430 176.790 371.600 ;
        RECT 211.460 371.520 211.650 371.530 ;
        RECT 174.820 370.990 175.200 371.000 ;
        RECT 174.820 370.930 175.290 370.990 ;
        RECT 176.540 370.970 176.720 371.430 ;
        RECT 176.730 371.250 177.350 371.420 ;
        RECT 211.450 371.230 211.650 371.520 ;
        RECT 174.480 370.880 175.290 370.930 ;
        RECT 174.470 370.820 175.290 370.880 ;
        RECT 174.470 370.760 175.210 370.820 ;
        RECT 175.760 370.800 176.720 370.970 ;
        RECT 211.370 370.900 211.660 371.230 ;
        RECT 174.820 370.710 175.210 370.760 ;
        RECT 211.850 370.420 212.020 372.030 ;
        RECT 212.630 371.480 212.860 372.170 ;
        RECT 220.050 371.560 225.110 372.390 ;
        RECT 250.490 372.310 250.690 372.660 ;
        RECT 252.730 372.540 253.060 372.730 ;
        RECT 252.730 372.500 253.050 372.540 ;
        RECT 253.130 372.420 253.330 372.750 ;
        RECT 253.610 372.610 253.960 372.940 ;
        RECT 254.440 373.030 254.760 373.070 ;
        RECT 254.440 372.840 254.770 373.030 ;
        RECT 254.960 372.850 255.190 373.450 ;
        RECT 255.800 373.090 255.970 374.700 ;
        RECT 256.160 373.890 256.450 374.220 ;
        RECT 256.170 373.600 256.370 373.890 ;
        RECT 256.170 373.590 256.360 373.600 ;
        RECT 256.530 373.420 256.740 373.430 ;
        RECT 256.520 372.840 256.740 373.420 ;
        RECT 254.440 372.810 254.760 372.840 ;
        RECT 256.530 372.810 256.740 372.840 ;
        RECT 253.720 372.420 253.920 372.610 ;
        RECT 254.720 372.540 255.250 372.710 ;
        RECT 256.530 372.460 256.730 372.810 ;
        RECT 250.490 372.280 250.700 372.310 ;
        RECT 224.560 371.480 225.040 371.560 ;
        RECT 248.920 371.480 249.150 372.170 ;
        RECT 173.430 370.320 173.780 370.420 ;
        RECT 177.020 370.370 177.190 370.410 ;
        RECT 176.040 370.350 177.190 370.370 ;
        RECT 175.090 370.320 175.550 370.350 ;
        RECT 172.020 370.150 172.780 370.320 ;
        RECT 173.030 370.150 174.200 370.320 ;
        RECT 174.440 370.180 175.550 370.320 ;
        RECT 176.000 370.180 177.190 370.350 ;
        RECT 211.840 370.230 212.020 370.420 ;
        RECT 212.680 370.330 212.850 371.480 ;
        RECT 224.560 371.380 224.890 371.480 ;
        RECT 224.560 371.230 224.710 371.380 ;
        RECT 217.310 371.190 217.630 371.230 ;
        RECT 217.300 371.000 217.630 371.190 ;
        RECT 217.310 370.970 217.630 371.000 ;
        RECT 244.150 371.190 244.470 371.230 ;
        RECT 244.150 371.000 244.480 371.190 ;
        RECT 244.150 370.970 244.470 371.000 ;
        RECT 248.930 370.330 249.100 371.480 ;
        RECT 249.760 370.420 249.930 372.030 ;
        RECT 250.480 371.700 250.700 372.280 ;
        RECT 252.730 372.290 253.050 372.330 ;
        RECT 252.730 372.100 253.060 372.290 ;
        RECT 252.730 372.070 253.050 372.100 ;
        RECT 253.130 372.080 253.330 372.410 ;
        RECT 253.720 372.220 253.920 372.410 ;
        RECT 254.430 372.310 254.750 372.350 ;
        RECT 253.410 371.890 253.600 371.900 ;
        RECT 253.610 371.890 253.960 372.220 ;
        RECT 254.430 372.120 254.760 372.310 ;
        RECT 254.430 372.090 254.750 372.120 ;
        RECT 250.490 371.690 250.700 371.700 ;
        RECT 250.130 371.520 250.320 371.530 ;
        RECT 250.130 371.230 250.330 371.520 ;
        RECT 252.500 371.380 252.670 371.710 ;
        RECT 252.680 371.640 253.000 371.680 ;
        RECT 252.680 371.450 253.010 371.640 ;
        RECT 252.680 371.420 253.000 371.450 ;
        RECT 253.130 371.420 253.330 371.750 ;
        RECT 253.410 371.560 253.960 371.890 ;
        RECT 253.610 371.300 253.960 371.560 ;
        RECT 253.610 371.230 253.980 371.300 ;
        RECT 250.120 370.900 250.410 371.230 ;
        RECT 253.790 371.070 253.980 371.230 ;
        RECT 254.440 371.170 255.140 371.350 ;
        RECT 249.760 370.230 249.940 370.420 ;
        RECT 174.440 370.150 175.260 370.180 ;
        RECT 172.020 370.140 172.250 370.150 ;
        RECT 171.980 369.700 172.250 370.140 ;
        RECT 175.000 370.010 175.260 370.150 ;
        RECT 252.500 370.120 252.670 370.450 ;
        RECT 252.680 370.380 253.000 370.410 ;
        RECT 252.680 370.190 253.010 370.380 ;
        RECT 252.680 370.150 253.000 370.190 ;
        RECT 253.130 370.080 253.330 370.410 ;
        RECT 253.610 370.270 253.960 370.600 ;
        RECT 173.460 369.700 173.790 369.960 ;
        RECT 174.410 369.910 174.700 369.940 ;
        RECT 174.370 369.740 174.700 369.910 ;
        RECT 174.410 369.700 174.700 369.740 ;
        RECT 175.000 369.840 176.180 370.010 ;
        RECT 175.000 369.700 175.260 369.840 ;
        RECT 171.430 369.560 171.600 369.620 ;
        RECT 171.400 369.340 171.620 369.560 ;
        RECT 171.950 369.520 172.280 369.700 ;
        RECT 172.530 369.530 174.690 369.700 ;
        RECT 174.930 369.530 175.260 369.700 ;
        RECT 175.400 369.690 176.180 369.840 ;
        RECT 175.030 369.480 175.260 369.530 ;
        RECT 171.430 369.290 171.600 369.340 ;
        RECT 175.030 369.250 175.200 369.480 ;
        RECT 175.550 369.340 175.760 369.670 ;
        RECT 176.000 369.400 176.180 369.690 ;
        RECT 176.460 369.680 176.790 369.850 ;
        RECT 223.750 369.680 223.940 370.000 ;
        RECT 237.840 369.680 238.030 370.000 ;
        RECT 248.160 369.830 248.480 369.870 ;
        RECT 174.820 369.240 175.200 369.250 ;
        RECT 174.820 369.180 175.290 369.240 ;
        RECT 176.540 369.220 176.720 369.680 ;
        RECT 176.730 369.500 177.350 369.670 ;
        RECT 223.750 369.590 224.030 369.680 ;
        RECT 220.390 369.450 224.030 369.590 ;
        RECT 237.750 369.590 238.030 369.680 ;
        RECT 248.150 369.640 248.480 369.830 ;
        RECT 248.160 369.630 248.480 369.640 ;
        RECT 248.150 369.610 248.480 369.630 ;
        RECT 248.760 369.790 249.090 369.960 ;
        RECT 249.200 369.880 249.530 370.050 ;
        RECT 253.410 369.940 253.960 370.270 ;
        RECT 254.450 370.100 255.150 370.750 ;
        RECT 253.410 369.930 253.600 369.940 ;
        RECT 237.750 369.450 241.390 369.590 ;
        RECT 220.390 369.410 223.940 369.450 ;
        RECT 174.480 369.130 175.290 369.180 ;
        RECT 174.470 369.070 175.290 369.130 ;
        RECT 174.470 369.010 175.210 369.070 ;
        RECT 175.760 369.050 176.720 369.220 ;
        RECT 174.820 368.960 175.210 369.010 ;
        RECT 147.310 368.830 147.630 368.870 ;
        RECT 148.400 368.840 148.720 368.880 ;
        RECT 147.310 368.760 147.640 368.830 ;
        RECT 147.310 368.610 147.680 368.760 ;
        RECT 147.480 368.430 147.680 368.610 ;
        RECT 148.070 368.430 148.270 368.760 ;
        RECT 148.400 368.650 148.730 368.840 ;
        RECT 148.400 368.620 148.720 368.650 ;
        RECT 173.430 368.570 173.780 368.670 ;
        RECT 177.020 368.620 177.190 368.660 ;
        RECT 176.040 368.600 177.190 368.620 ;
        RECT 175.090 368.570 175.550 368.600 ;
        RECT 172.020 368.400 172.780 368.570 ;
        RECT 173.030 368.400 174.200 368.570 ;
        RECT 174.440 368.430 175.550 368.570 ;
        RECT 176.000 368.430 177.190 368.600 ;
        RECT 174.440 368.400 175.260 368.430 ;
        RECT 172.020 368.390 172.250 368.400 ;
        RECT 146.930 368.120 147.260 368.290 ;
        RECT 145.770 367.920 146.090 367.960 ;
        RECT 171.980 367.950 172.250 368.390 ;
        RECT 175.000 368.260 175.260 368.400 ;
        RECT 173.460 367.950 173.790 368.210 ;
        RECT 174.410 368.160 174.700 368.190 ;
        RECT 174.370 367.990 174.700 368.160 ;
        RECT 174.410 367.950 174.700 367.990 ;
        RECT 175.000 368.090 176.180 368.260 ;
        RECT 198.050 368.180 198.720 369.050 ;
        RECT 210.330 368.200 212.430 369.050 ;
        RECT 223.750 368.990 223.940 369.410 ;
        RECT 237.840 369.410 242.060 369.450 ;
        RECT 237.840 368.990 238.030 369.410 ;
        RECT 238.820 369.270 239.460 369.410 ;
        RECT 239.840 369.280 240.190 369.410 ;
        RECT 240.290 369.320 240.620 369.410 ;
        RECT 240.370 369.240 240.620 369.320 ;
        RECT 240.920 369.270 242.060 369.410 ;
        RECT 239.220 368.890 239.390 368.900 ;
        RECT 239.220 368.850 239.620 368.890 ;
        RECT 175.000 367.950 175.260 368.090 ;
        RECT 145.770 367.730 146.100 367.920 ;
        RECT 147.320 367.840 147.640 367.880 ;
        RECT 148.410 367.850 148.730 367.890 ;
        RECT 147.320 367.770 147.650 367.840 ;
        RECT 147.660 367.770 147.830 367.820 ;
        RECT 148.150 367.770 148.340 367.810 ;
        RECT 147.320 367.740 147.830 367.770 ;
        RECT 148.080 367.740 148.340 367.770 ;
        RECT 145.770 367.700 146.090 367.730 ;
        RECT 145.790 367.630 146.000 367.700 ;
        RECT 147.320 367.620 148.340 367.740 ;
        RECT 148.410 367.660 148.740 367.850 ;
        RECT 171.430 367.810 171.600 367.870 ;
        RECT 148.410 367.630 148.730 367.660 ;
        RECT 147.490 367.580 148.340 367.620 ;
        RECT 171.400 367.590 171.620 367.810 ;
        RECT 171.950 367.770 172.280 367.950 ;
        RECT 172.530 367.780 174.690 367.950 ;
        RECT 174.930 367.780 175.260 367.950 ;
        RECT 175.400 367.940 176.180 368.090 ;
        RECT 175.030 367.730 175.260 367.780 ;
        RECT 147.490 367.490 148.280 367.580 ;
        RECT 171.430 367.540 171.600 367.590 ;
        RECT 175.030 367.500 175.200 367.730 ;
        RECT 175.550 367.590 175.760 367.920 ;
        RECT 176.000 367.650 176.180 367.940 ;
        RECT 176.460 367.930 176.790 368.100 ;
        RECT 147.490 367.440 147.840 367.490 ;
        RECT 148.080 367.440 148.280 367.490 ;
        RECT 174.820 367.490 175.200 367.500 ;
        RECT 147.660 367.430 147.840 367.440 ;
        RECT 174.820 367.430 175.290 367.490 ;
        RECT 176.540 367.470 176.720 367.930 ;
        RECT 176.730 367.750 177.350 367.920 ;
        RECT 211.370 367.860 211.660 368.190 ;
        RECT 211.450 367.570 211.650 367.860 ;
        RECT 211.460 367.560 211.650 367.570 ;
        RECT 174.480 367.380 175.290 367.430 ;
        RECT 174.470 367.320 175.290 367.380 ;
        RECT 146.940 367.130 147.270 367.300 ;
        RECT 174.470 367.260 175.210 367.320 ;
        RECT 175.760 367.300 176.720 367.470 ;
        RECT 211.080 367.390 211.290 367.400 ;
        RECT 174.820 367.210 175.210 367.260 ;
        RECT 145.750 367.000 146.070 367.040 ;
        RECT 145.750 366.810 146.080 367.000 ;
        RECT 147.320 366.850 147.640 366.890 ;
        RECT 148.410 366.860 148.730 366.900 ;
        RECT 145.750 366.780 146.070 366.810 ;
        RECT 147.320 366.780 147.650 366.850 ;
        RECT 147.320 366.630 147.690 366.780 ;
        RECT 147.490 366.450 147.690 366.630 ;
        RECT 148.080 366.450 148.280 366.780 ;
        RECT 148.410 366.670 148.740 366.860 ;
        RECT 173.430 366.820 173.780 366.920 ;
        RECT 177.020 366.870 177.190 366.910 ;
        RECT 176.040 366.850 177.190 366.870 ;
        RECT 175.090 366.820 175.550 366.850 ;
        RECT 148.410 366.640 148.730 366.670 ;
        RECT 172.020 366.650 172.780 366.820 ;
        RECT 173.030 366.650 174.200 366.820 ;
        RECT 174.440 366.680 175.550 366.820 ;
        RECT 176.000 366.680 177.190 366.850 ;
        RECT 211.080 366.810 211.300 367.390 ;
        RECT 211.850 367.060 212.020 368.200 ;
        RECT 212.680 367.510 212.850 368.760 ;
        RECT 239.220 368.660 239.630 368.850 ;
        RECT 239.830 368.820 240.020 368.930 ;
        RECT 239.830 368.700 240.170 368.820 ;
        RECT 239.220 368.630 239.620 368.660 ;
        RECT 239.880 368.650 240.170 368.700 ;
        RECT 239.220 368.600 239.390 368.630 ;
        RECT 240.450 368.560 240.620 369.240 ;
        RECT 246.690 369.260 247.010 369.300 ;
        RECT 246.690 369.070 247.020 369.260 ;
        RECT 246.690 369.040 247.010 369.070 ;
        RECT 247.090 369.050 247.290 369.380 ;
        RECT 247.680 369.190 247.880 369.380 ;
        RECT 248.150 369.300 248.320 369.610 ;
        RECT 248.760 369.510 249.120 369.790 ;
        RECT 248.410 369.340 249.120 369.510 ;
        RECT 252.730 369.730 253.050 369.760 ;
        RECT 252.730 369.540 253.060 369.730 ;
        RECT 252.730 369.500 253.050 369.540 ;
        RECT 253.130 369.420 253.330 369.750 ;
        RECT 253.610 369.610 253.960 369.940 ;
        RECT 254.350 369.870 255.150 370.100 ;
        RECT 254.350 369.840 254.670 369.870 ;
        RECT 253.720 369.420 253.920 369.610 ;
        RECT 254.450 369.260 255.160 369.430 ;
        RECT 248.350 369.220 248.670 369.260 ;
        RECT 240.960 368.890 241.130 368.900 ;
        RECT 240.960 368.850 241.290 368.890 ;
        RECT 240.960 368.660 241.300 368.850 ;
        RECT 241.940 368.830 242.130 368.940 ;
        RECT 241.820 368.820 242.130 368.830 ;
        RECT 241.570 368.710 242.130 368.820 ;
        RECT 247.370 368.860 247.560 368.870 ;
        RECT 247.570 368.860 247.920 369.190 ;
        RECT 248.350 369.040 248.680 369.220 ;
        RECT 248.310 369.030 248.680 369.040 ;
        RECT 248.310 369.000 248.670 369.030 ;
        RECT 240.960 368.630 241.290 368.660 ;
        RECT 241.570 368.650 241.950 368.710 ;
        RECT 240.960 368.600 241.130 368.630 ;
        RECT 217.310 368.430 217.630 368.470 ;
        RECT 217.300 368.240 217.630 368.430 ;
        RECT 244.150 368.430 244.470 368.470 ;
        RECT 222.680 368.370 222.910 368.410 ;
        RECT 238.870 368.370 239.100 368.410 ;
        RECT 217.310 368.210 217.630 368.240 ;
        RECT 244.150 368.240 244.480 368.430 ;
        RECT 246.460 368.350 246.630 368.680 ;
        RECT 246.640 368.610 246.960 368.650 ;
        RECT 246.640 368.420 246.970 368.610 ;
        RECT 246.640 368.390 246.960 368.420 ;
        RECT 247.090 368.390 247.290 368.720 ;
        RECT 247.370 368.530 247.920 368.860 ;
        RECT 248.300 368.900 248.630 369.000 ;
        RECT 254.800 368.980 255.160 369.260 ;
        RECT 248.300 368.810 249.110 368.900 ;
        RECT 248.310 368.780 249.110 368.810 ;
        RECT 244.150 368.210 244.470 368.240 ;
        RECT 247.570 368.210 247.920 368.530 ;
        RECT 247.500 368.200 247.920 368.210 ;
        RECT 224.600 367.910 224.920 367.950 ;
        RECT 224.590 367.720 224.920 367.910 ;
        RECT 238.840 367.770 239.050 368.200 ;
        RECT 247.500 368.180 247.820 368.200 ;
        RECT 247.500 367.990 247.830 368.180 ;
        RECT 248.410 368.020 249.110 368.780 ;
        RECT 249.760 368.670 249.940 368.860 ;
        RECT 254.800 368.810 255.130 368.980 ;
        RECT 255.240 368.720 255.570 368.890 ;
        RECT 247.500 367.950 247.820 367.990 ;
        RECT 238.860 367.750 239.030 367.770 ;
        RECT 224.600 367.690 224.920 367.720 ;
        RECT 224.720 367.550 224.740 367.690 ;
        RECT 239.360 367.630 239.550 367.740 ;
        RECT 212.630 366.820 212.860 367.510 ;
        RECT 224.720 367.470 225.070 367.550 ;
        RECT 239.360 367.510 239.780 367.630 ;
        RECT 211.080 366.780 211.290 366.810 ;
        RECT 174.440 366.650 175.260 366.680 ;
        RECT 172.020 366.640 172.250 366.650 ;
        RECT 146.940 366.160 147.270 366.310 ;
        RECT 171.980 366.200 172.250 366.640 ;
        RECT 175.000 366.510 175.260 366.650 ;
        RECT 173.460 366.200 173.790 366.460 ;
        RECT 174.410 366.410 174.700 366.440 ;
        RECT 174.370 366.240 174.700 366.410 ;
        RECT 174.410 366.200 174.700 366.240 ;
        RECT 175.000 366.340 176.180 366.510 ;
        RECT 211.090 366.430 211.290 366.780 ;
        RECT 212.570 366.510 213.100 366.680 ;
        RECT 220.020 366.620 225.070 367.470 ;
        RECT 239.260 367.460 239.780 367.510 ;
        RECT 240.130 367.460 241.390 367.640 ;
        RECT 247.750 367.630 247.940 367.860 ;
        RECT 248.930 367.600 249.100 368.020 ;
        RECT 239.260 367.380 239.450 367.460 ;
        RECT 239.240 367.350 239.450 367.380 ;
        RECT 239.230 367.340 239.450 367.350 ;
        RECT 240.620 367.340 240.950 367.460 ;
        RECT 239.110 367.290 239.450 367.340 ;
        RECT 238.980 367.260 239.450 367.290 ;
        RECT 238.940 367.230 239.450 367.260 ;
        RECT 238.940 367.170 239.430 367.230 ;
        RECT 238.940 367.120 239.280 367.170 ;
        RECT 238.940 367.100 239.200 367.120 ;
        RECT 238.940 367.080 239.170 367.100 ;
        RECT 246.460 367.090 246.630 367.420 ;
        RECT 246.640 367.350 246.960 367.380 ;
        RECT 246.640 367.160 246.970 367.350 ;
        RECT 246.640 367.120 246.960 367.160 ;
        RECT 238.940 367.040 239.150 367.080 ;
        RECT 247.090 367.050 247.290 367.380 ;
        RECT 247.570 367.290 247.920 367.570 ;
        RECT 248.400 367.510 249.100 367.600 ;
        RECT 248.400 367.420 249.150 367.510 ;
        RECT 247.480 367.240 247.920 367.290 ;
        RECT 238.940 366.760 239.110 367.040 ;
        RECT 247.370 366.900 247.920 367.240 ;
        RECT 248.400 367.000 248.720 367.040 ;
        RECT 248.400 366.930 248.730 367.000 ;
        RECT 246.690 366.700 247.010 366.730 ;
        RECT 246.690 366.510 247.020 366.700 ;
        RECT 246.690 366.470 247.010 366.510 ;
        RECT 247.090 366.390 247.290 366.720 ;
        RECT 247.480 366.580 247.920 366.900 ;
        RECT 248.230 366.830 248.730 366.930 ;
        RECT 248.090 366.810 248.730 366.830 ;
        RECT 248.920 366.820 249.150 367.420 ;
        RECT 249.760 367.060 249.930 368.670 ;
        RECT 250.120 367.860 250.410 368.190 ;
        RECT 250.130 367.570 250.330 367.860 ;
        RECT 250.130 367.560 250.320 367.570 ;
        RECT 250.490 367.390 250.700 367.400 ;
        RECT 250.480 366.810 250.700 367.390 ;
        RECT 248.090 366.780 248.720 366.810 ;
        RECT 250.490 366.780 250.700 366.810 ;
        RECT 248.090 366.710 248.560 366.780 ;
        RECT 248.090 366.700 248.550 366.710 ;
        RECT 248.210 366.670 248.550 366.700 ;
        RECT 248.210 366.600 248.260 366.670 ;
        RECT 175.000 366.200 175.260 366.340 ;
        RECT 146.940 366.140 147.550 366.160 ;
        RECT 147.230 366.120 147.550 366.140 ;
        RECT 145.730 366.010 146.050 366.050 ;
        RECT 145.730 365.820 146.060 366.010 ;
        RECT 147.230 365.950 147.560 366.120 ;
        RECT 171.430 366.060 171.600 366.120 ;
        RECT 148.530 366.020 148.850 366.060 ;
        RECT 147.230 365.900 147.710 365.950 ;
        RECT 145.730 365.790 146.050 365.820 ;
        RECT 147.400 365.770 147.710 365.900 ;
        RECT 147.380 365.750 147.710 365.770 ;
        RECT 147.540 365.620 147.710 365.750 ;
        RECT 148.220 365.620 148.390 365.950 ;
        RECT 148.530 365.830 148.860 366.020 ;
        RECT 171.400 365.840 171.620 366.060 ;
        RECT 171.950 366.020 172.280 366.200 ;
        RECT 172.530 366.030 174.690 366.200 ;
        RECT 174.930 366.030 175.260 366.200 ;
        RECT 175.400 366.190 176.180 366.340 ;
        RECT 175.030 365.980 175.260 366.030 ;
        RECT 148.530 365.800 148.850 365.830 ;
        RECT 171.430 365.790 171.600 365.840 ;
        RECT 175.030 365.750 175.200 365.980 ;
        RECT 175.550 365.840 175.760 366.170 ;
        RECT 176.000 365.900 176.180 366.190 ;
        RECT 176.460 366.180 176.790 366.350 ;
        RECT 174.820 365.740 175.200 365.750 ;
        RECT 174.820 365.680 175.290 365.740 ;
        RECT 176.540 365.720 176.720 366.180 ;
        RECT 176.730 366.000 177.350 366.170 ;
        RECT 238.820 366.070 239.460 366.250 ;
        RECT 239.840 366.080 240.190 366.250 ;
        RECT 240.290 366.240 240.480 366.350 ;
        RECT 246.690 366.260 247.010 366.300 ;
        RECT 240.290 366.120 240.620 366.240 ;
        RECT 240.370 366.040 240.620 366.120 ;
        RECT 240.920 366.070 242.060 366.250 ;
        RECT 246.690 366.070 247.020 366.260 ;
        RECT 246.690 366.040 247.010 366.070 ;
        RECT 247.090 366.050 247.290 366.380 ;
        RECT 247.480 366.230 247.660 366.580 ;
        RECT 247.680 366.390 247.880 366.580 ;
        RECT 247.680 366.190 247.880 366.380 ;
        RECT 248.130 366.270 248.300 366.600 ;
        RECT 248.680 366.510 249.210 366.680 ;
        RECT 250.490 366.430 250.690 366.780 ;
        RECT 248.390 366.280 248.710 366.320 ;
        RECT 248.390 366.190 248.720 366.280 ;
        RECT 174.480 365.630 175.290 365.680 ;
        RECT 174.470 365.570 175.290 365.630 ;
        RECT 174.470 365.510 175.210 365.570 ;
        RECT 175.760 365.550 176.720 365.720 ;
        RECT 174.820 365.460 175.210 365.510 ;
        RECT 147.160 365.420 147.590 365.440 ;
        RECT 147.140 365.250 147.590 365.420 ;
        RECT 147.160 365.230 147.590 365.250 ;
        RECT 147.230 365.130 147.550 365.170 ;
        RECT 147.230 364.960 147.560 365.130 ;
        RECT 148.530 365.030 148.850 365.070 ;
        RECT 147.230 364.910 147.710 364.960 ;
        RECT 147.400 364.780 147.710 364.910 ;
        RECT 147.380 364.760 147.710 364.780 ;
        RECT 147.540 364.630 147.710 364.760 ;
        RECT 148.220 364.630 148.390 364.960 ;
        RECT 148.530 364.840 148.860 365.030 ;
        RECT 148.530 364.810 148.850 364.840 ;
        RECT 227.900 364.700 228.100 365.710 ;
        RECT 233.650 364.700 233.940 365.710 ;
        RECT 239.220 365.690 239.390 365.700 ;
        RECT 238.940 365.410 239.110 365.690 ;
        RECT 239.220 365.650 239.620 365.690 ;
        RECT 239.220 365.460 239.630 365.650 ;
        RECT 239.830 365.620 240.020 365.730 ;
        RECT 239.830 365.500 240.170 365.620 ;
        RECT 239.220 365.430 239.620 365.460 ;
        RECT 239.880 365.450 240.170 365.500 ;
        RECT 238.940 365.370 239.150 365.410 ;
        RECT 239.220 365.400 239.390 365.430 ;
        RECT 238.940 365.350 239.170 365.370 ;
        RECT 240.450 365.360 240.620 366.040 ;
        RECT 247.370 365.860 247.560 365.870 ;
        RECT 247.570 365.860 247.920 366.190 ;
        RECT 248.390 366.060 248.860 366.190 ;
        RECT 248.530 365.980 248.860 366.060 ;
        RECT 248.670 365.960 248.860 365.980 ;
        RECT 240.960 365.690 241.130 365.700 ;
        RECT 240.960 365.650 241.290 365.690 ;
        RECT 240.960 365.460 241.300 365.650 ;
        RECT 241.940 365.630 242.130 365.740 ;
        RECT 241.820 365.620 242.130 365.630 ;
        RECT 241.570 365.510 242.130 365.620 ;
        RECT 240.960 365.430 241.290 365.460 ;
        RECT 241.570 365.450 241.950 365.510 ;
        RECT 240.960 365.400 241.130 365.430 ;
        RECT 246.460 365.350 246.630 365.680 ;
        RECT 246.640 365.610 246.960 365.650 ;
        RECT 246.640 365.420 246.970 365.610 ;
        RECT 246.640 365.390 246.960 365.420 ;
        RECT 247.090 365.390 247.290 365.720 ;
        RECT 247.370 365.530 247.920 365.860 ;
        RECT 238.940 365.330 239.200 365.350 ;
        RECT 238.940 365.280 239.280 365.330 ;
        RECT 238.940 365.220 239.430 365.280 ;
        RECT 247.570 365.270 247.920 365.530 ;
        RECT 238.940 365.190 239.450 365.220 ;
        RECT 247.570 365.200 247.940 365.270 ;
        RECT 238.980 365.160 239.450 365.190 ;
        RECT 239.110 365.110 239.450 365.160 ;
        RECT 239.230 365.100 239.450 365.110 ;
        RECT 239.240 365.070 239.450 365.100 ;
        RECT 147.160 364.430 147.590 364.450 ;
        RECT 147.140 364.260 147.590 364.430 ;
        RECT 147.160 364.240 147.590 364.260 ;
        RECT 238.840 364.250 239.050 365.000 ;
        RECT 239.260 364.990 239.450 365.070 ;
        RECT 240.620 364.990 240.950 365.110 ;
        RECT 247.750 365.040 247.940 365.200 ;
        RECT 248.400 365.140 249.100 365.320 ;
        RECT 239.260 364.940 239.780 364.990 ;
        RECT 239.360 364.820 239.780 364.940 ;
        RECT 239.360 364.710 239.550 364.820 ;
        RECT 240.130 364.810 241.390 364.990 ;
        RECT 239.360 364.430 239.550 364.540 ;
        RECT 239.360 364.310 239.780 364.430 ;
        RECT 239.260 364.260 239.780 364.310 ;
        RECT 240.130 364.260 241.390 364.440 ;
        RECT 239.260 364.180 239.450 364.260 ;
        RECT 147.230 364.140 147.550 364.180 ;
        RECT 239.240 364.150 239.450 364.180 ;
        RECT 239.230 364.140 239.450 364.150 ;
        RECT 240.620 364.140 240.950 364.260 ;
        RECT 147.230 363.970 147.560 364.140 ;
        RECT 239.110 364.090 239.450 364.140 ;
        RECT 246.460 364.090 246.630 364.420 ;
        RECT 246.640 364.350 246.960 364.380 ;
        RECT 246.640 364.160 246.970 364.350 ;
        RECT 246.640 364.120 246.960 364.160 ;
        RECT 148.530 364.040 148.850 364.080 ;
        RECT 238.980 364.060 239.450 364.090 ;
        RECT 147.230 363.920 147.710 363.970 ;
        RECT 147.400 363.790 147.710 363.920 ;
        RECT 147.380 363.780 147.710 363.790 ;
        RECT 147.380 363.770 147.870 363.780 ;
        RECT 147.540 363.690 147.870 363.770 ;
        RECT 147.540 363.610 147.930 363.690 ;
        RECT 148.220 363.640 148.390 363.970 ;
        RECT 148.530 363.850 148.860 364.040 ;
        RECT 238.940 364.030 239.450 364.060 ;
        RECT 247.090 364.050 247.290 364.380 ;
        RECT 247.570 364.240 247.920 364.570 ;
        RECT 238.940 363.970 239.430 364.030 ;
        RECT 238.940 363.920 239.280 363.970 ;
        RECT 238.940 363.900 239.200 363.920 ;
        RECT 247.370 363.910 247.920 364.240 ;
        RECT 248.410 364.070 249.110 364.720 ;
        RECT 247.370 363.900 247.560 363.910 ;
        RECT 238.940 363.880 239.170 363.900 ;
        RECT 148.530 363.820 148.850 363.850 ;
        RECT 238.940 363.840 239.150 363.880 ;
        RECT 147.700 363.500 147.930 363.610 ;
        RECT 238.940 363.560 239.110 363.840 ;
        RECT 239.220 363.820 239.390 363.850 ;
        RECT 239.220 363.790 239.620 363.820 ;
        RECT 239.220 363.600 239.630 363.790 ;
        RECT 239.880 363.750 240.170 363.800 ;
        RECT 239.830 363.630 240.170 363.750 ;
        RECT 239.220 363.560 239.620 363.600 ;
        RECT 239.220 363.550 239.390 363.560 ;
        RECT 239.830 363.520 240.020 363.630 ;
        RECT 147.160 363.440 147.590 363.460 ;
        RECT 147.140 363.270 147.590 363.440 ;
        RECT 147.160 363.250 147.590 363.270 ;
        RECT 240.450 363.210 240.620 363.890 ;
        RECT 240.960 363.820 241.130 363.850 ;
        RECT 240.960 363.790 241.290 363.820 ;
        RECT 242.120 363.800 242.440 363.840 ;
        RECT 240.960 363.600 241.300 363.790 ;
        RECT 241.570 363.740 241.950 363.800 ;
        RECT 242.110 363.740 242.440 363.800 ;
        RECT 241.570 363.630 242.440 363.740 ;
        RECT 241.820 363.620 242.440 363.630 ;
        RECT 240.960 363.560 241.290 363.600 ;
        RECT 241.940 363.580 242.440 363.620 ;
        RECT 246.690 363.700 247.010 363.730 ;
        RECT 240.960 363.550 241.130 363.560 ;
        RECT 241.940 363.510 242.280 363.580 ;
        RECT 242.110 363.270 242.280 363.510 ;
        RECT 246.690 363.510 247.020 363.700 ;
        RECT 246.690 363.470 247.010 363.510 ;
        RECT 247.090 363.390 247.290 363.720 ;
        RECT 247.570 363.580 247.920 363.910 ;
        RECT 248.310 363.840 249.110 364.070 ;
        RECT 248.310 363.810 248.630 363.840 ;
        RECT 247.680 363.390 247.880 363.580 ;
        RECT 248.410 363.230 249.120 363.400 ;
        RECT 238.820 363.000 239.460 363.180 ;
        RECT 239.840 363.000 240.190 363.170 ;
        RECT 240.370 363.130 240.620 363.210 ;
        RECT 240.290 363.010 240.620 363.130 ;
        RECT 240.290 362.900 240.480 363.010 ;
        RECT 240.920 363.000 242.060 363.180 ;
        RECT 242.270 362.970 242.590 363.010 ;
        RECT 186.410 362.440 186.580 362.860 ;
        RECT 187.220 362.740 187.460 362.770 ;
        RECT 186.890 362.570 187.460 362.740 ;
        RECT 187.700 362.570 189.040 362.740 ;
        RECT 189.490 362.570 190.450 362.740 ;
        RECT 187.220 362.530 187.460 362.570 ;
        RECT 190.000 362.560 190.170 362.570 ;
        RECT 186.340 362.220 186.510 362.260 ;
        RECT 186.280 362.050 186.510 362.220 ;
        RECT 189.630 362.120 189.970 362.300 ;
        RECT 186.340 361.840 186.510 362.050 ;
        RECT 186.280 361.670 186.510 361.840 ;
        RECT 186.580 361.830 186.770 362.060 ;
        RECT 186.870 361.950 187.240 362.120 ;
        RECT 187.700 361.950 190.450 362.120 ;
        RECT 186.870 361.770 187.240 361.940 ;
        RECT 187.700 361.770 190.450 361.940 ;
        RECT 174.820 361.620 175.210 361.670 ;
        RECT 186.340 361.630 186.510 361.670 ;
        RECT 174.470 361.560 175.210 361.620 ;
        RECT 189.630 361.590 189.970 361.770 ;
        RECT 174.470 361.500 175.290 361.560 ;
        RECT 174.480 361.450 175.290 361.500 ;
        RECT 174.820 361.390 175.290 361.450 ;
        RECT 175.760 361.410 176.720 361.580 ;
        RECT 174.820 361.380 175.200 361.390 ;
        RECT 171.430 361.290 171.600 361.340 ;
        RECT 171.400 361.070 171.620 361.290 ;
        RECT 175.030 361.150 175.200 361.380 ;
        RECT 171.430 361.010 171.600 361.070 ;
        RECT 171.950 360.930 172.280 361.110 ;
        RECT 175.030 361.100 175.260 361.150 ;
        RECT 172.530 360.930 174.690 361.100 ;
        RECT 174.930 360.930 175.260 361.100 ;
        RECT 175.550 360.960 175.760 361.290 ;
        RECT 176.000 360.940 176.180 361.230 ;
        RECT 176.540 360.950 176.720 361.410 ;
        RECT 176.730 360.960 177.350 361.130 ;
        RECT 186.410 361.030 186.580 361.450 ;
        RECT 187.220 361.320 187.460 361.360 ;
        RECT 190.000 361.320 190.170 361.330 ;
        RECT 186.890 361.150 187.460 361.320 ;
        RECT 187.700 361.150 189.040 361.320 ;
        RECT 189.490 361.150 190.450 361.320 ;
        RECT 187.220 361.120 187.460 361.150 ;
        RECT 190.980 361.080 191.150 362.810 ;
        RECT 191.380 361.970 191.550 362.860 ;
        RECT 242.260 362.780 242.590 362.970 ;
        RECT 248.760 362.950 249.120 363.230 ;
        RECT 248.760 362.780 249.090 362.950 ;
        RECT 242.270 362.750 242.590 362.780 ;
        RECT 249.200 362.690 249.530 362.860 ;
        RECT 251.110 362.800 251.290 364.850 ;
        RECT 251.840 364.590 252.170 364.760 ;
        RECT 251.920 362.810 252.090 364.590 ;
        RECT 238.940 362.210 239.110 362.490 ;
        RECT 238.940 362.170 239.150 362.210 ;
        RECT 238.940 362.150 239.170 362.170 ;
        RECT 241.460 362.150 241.780 362.180 ;
        RECT 238.940 362.130 239.200 362.150 ;
        RECT 238.940 362.080 239.280 362.130 ;
        RECT 238.940 362.020 239.430 362.080 ;
        RECT 238.940 361.990 239.450 362.020 ;
        RECT 238.980 361.960 239.450 361.990 ;
        RECT 191.380 361.030 191.550 361.920 ;
        RECT 239.110 361.910 239.450 361.960 ;
        RECT 241.460 361.960 241.790 362.150 ;
        RECT 241.460 361.920 241.780 361.960 ;
        RECT 239.230 361.900 239.450 361.910 ;
        RECT 239.240 361.870 239.450 361.900 ;
        RECT 239.260 361.790 239.450 361.870 ;
        RECT 240.620 361.790 240.950 361.910 ;
        RECT 239.260 361.740 239.780 361.790 ;
        RECT 239.360 361.620 239.780 361.740 ;
        RECT 239.360 361.510 239.550 361.620 ;
        RECT 240.130 361.610 241.390 361.790 ;
        RECT 238.860 361.480 239.030 361.500 ;
        RECT 238.840 361.050 239.050 361.480 ;
        RECT 171.980 360.490 172.250 360.930 ;
        RECT 173.460 360.670 173.790 360.930 ;
        RECT 174.410 360.890 174.700 360.930 ;
        RECT 174.370 360.720 174.700 360.890 ;
        RECT 174.410 360.690 174.700 360.720 ;
        RECT 175.000 360.790 175.260 360.930 ;
        RECT 175.400 360.790 176.180 360.940 ;
        RECT 172.020 360.480 172.250 360.490 ;
        RECT 175.000 360.620 176.180 360.790 ;
        RECT 176.460 360.780 176.790 360.950 ;
        RECT 239.220 360.620 239.390 360.650 ;
        RECT 175.000 360.480 175.260 360.620 ;
        RECT 172.020 360.310 172.780 360.480 ;
        RECT 173.030 360.310 174.200 360.480 ;
        RECT 174.440 360.450 175.260 360.480 ;
        RECT 239.220 360.590 239.620 360.620 ;
        RECT 174.440 360.310 175.550 360.450 ;
        RECT 173.430 360.210 173.780 360.310 ;
        RECT 175.090 360.280 175.550 360.310 ;
        RECT 176.000 360.280 177.190 360.450 ;
        RECT 239.220 360.400 239.630 360.590 ;
        RECT 239.880 360.550 240.170 360.600 ;
        RECT 239.830 360.430 240.170 360.550 ;
        RECT 239.220 360.360 239.620 360.400 ;
        RECT 239.220 360.350 239.390 360.360 ;
        RECT 239.830 360.320 240.020 360.430 ;
        RECT 176.040 360.260 177.190 360.280 ;
        RECT 177.020 360.220 177.190 360.260 ;
        RECT 240.450 360.010 240.620 360.690 ;
        RECT 240.960 360.620 241.130 360.650 ;
        RECT 240.960 360.590 241.290 360.620 ;
        RECT 241.440 360.600 241.620 361.260 ;
        RECT 242.190 360.870 242.510 360.900 ;
        RECT 242.190 360.800 242.520 360.870 ;
        RECT 242.050 360.680 242.520 360.800 ;
        RECT 242.050 360.670 242.510 360.680 ;
        RECT 242.170 360.640 242.510 360.670 ;
        RECT 240.960 360.400 241.300 360.590 ;
        RECT 241.440 360.540 241.950 360.600 ;
        RECT 242.170 360.570 242.220 360.640 ;
        RECT 242.090 360.540 242.260 360.570 ;
        RECT 241.440 360.430 242.260 360.540 ;
        RECT 240.960 360.360 241.290 360.400 ;
        RECT 240.960 360.350 241.130 360.360 ;
        RECT 241.440 360.200 241.620 360.430 ;
        RECT 241.820 360.420 242.260 360.430 ;
        RECT 241.940 360.310 242.260 360.420 ;
        RECT 242.090 360.240 242.260 360.310 ;
        RECT 174.820 359.870 175.210 359.920 ;
        RECT 174.470 359.810 175.210 359.870 ;
        RECT 174.470 359.750 175.290 359.810 ;
        RECT 174.480 359.700 175.290 359.750 ;
        RECT 174.820 359.640 175.290 359.700 ;
        RECT 175.760 359.660 176.720 359.830 ;
        RECT 238.820 359.800 239.460 359.980 ;
        RECT 239.840 359.800 240.190 359.970 ;
        RECT 240.370 359.930 240.620 360.010 ;
        RECT 242.490 360.040 242.570 360.120 ;
        RECT 242.630 360.040 242.820 360.160 ;
        RECT 240.290 359.810 240.620 359.930 ;
        RECT 240.290 359.700 240.480 359.810 ;
        RECT 240.920 359.800 242.060 359.980 ;
        RECT 242.490 359.950 242.820 360.040 ;
        RECT 242.630 359.930 242.820 359.950 ;
        RECT 251.110 359.750 251.290 361.800 ;
        RECT 251.840 361.540 252.170 361.710 ;
        RECT 251.920 359.760 252.090 361.540 ;
        RECT 174.820 359.630 175.200 359.640 ;
        RECT 171.430 359.540 171.600 359.590 ;
        RECT 171.400 359.320 171.620 359.540 ;
        RECT 175.030 359.400 175.200 359.630 ;
        RECT 171.430 359.260 171.600 359.320 ;
        RECT 171.950 359.180 172.280 359.360 ;
        RECT 175.030 359.350 175.260 359.400 ;
        RECT 172.530 359.180 174.690 359.350 ;
        RECT 174.930 359.180 175.260 359.350 ;
        RECT 175.550 359.210 175.760 359.540 ;
        RECT 176.000 359.190 176.180 359.480 ;
        RECT 176.540 359.200 176.720 359.660 ;
        RECT 176.730 359.210 177.350 359.380 ;
        RECT 186.410 359.240 186.580 359.660 ;
        RECT 187.220 359.540 187.460 359.570 ;
        RECT 186.890 359.370 187.460 359.540 ;
        RECT 187.700 359.370 189.040 359.540 ;
        RECT 189.490 359.370 190.450 359.540 ;
        RECT 187.220 359.330 187.460 359.370 ;
        RECT 190.000 359.360 190.170 359.370 ;
        RECT 171.980 358.740 172.250 359.180 ;
        RECT 173.460 358.920 173.790 359.180 ;
        RECT 174.410 359.140 174.700 359.180 ;
        RECT 174.370 358.970 174.700 359.140 ;
        RECT 174.410 358.940 174.700 358.970 ;
        RECT 175.000 359.040 175.260 359.180 ;
        RECT 175.400 359.040 176.180 359.190 ;
        RECT 172.020 358.730 172.250 358.740 ;
        RECT 175.000 358.870 176.180 359.040 ;
        RECT 176.460 359.030 176.790 359.200 ;
        RECT 186.340 359.020 186.510 359.060 ;
        RECT 175.000 358.730 175.260 358.870 ;
        RECT 186.280 358.850 186.510 359.020 ;
        RECT 189.630 358.920 189.970 359.100 ;
        RECT 172.020 358.560 172.780 358.730 ;
        RECT 173.030 358.560 174.200 358.730 ;
        RECT 174.440 358.700 175.260 358.730 ;
        RECT 174.440 358.560 175.550 358.700 ;
        RECT 173.430 358.460 173.780 358.560 ;
        RECT 175.090 358.530 175.550 358.560 ;
        RECT 176.000 358.530 177.190 358.700 ;
        RECT 186.340 358.640 186.510 358.850 ;
        RECT 176.040 358.510 177.190 358.530 ;
        RECT 177.020 358.470 177.190 358.510 ;
        RECT 186.280 358.470 186.510 358.640 ;
        RECT 186.580 358.630 186.770 358.860 ;
        RECT 186.870 358.750 187.240 358.920 ;
        RECT 187.700 358.750 190.450 358.920 ;
        RECT 186.870 358.570 187.240 358.740 ;
        RECT 187.700 358.570 190.450 358.740 ;
        RECT 186.340 358.430 186.510 358.470 ;
        RECT 24.080 357.920 31.610 358.430 ;
        RECT 189.630 358.390 189.970 358.570 ;
        RECT 174.820 358.120 175.210 358.170 ;
        RECT 174.470 358.060 175.210 358.120 ;
        RECT 174.470 358.000 175.290 358.060 ;
        RECT 174.480 357.950 175.290 358.000 ;
        RECT 22.380 351.900 23.840 351.940 ;
        RECT 22.380 351.730 23.850 351.900 ;
        RECT 22.380 351.690 23.840 351.730 ;
        RECT 24.080 345.310 24.590 357.920 ;
        RECT 24.950 357.130 30.930 357.360 ;
        RECT 25.040 346.070 30.690 357.130 ;
        RECT 31.100 347.560 31.610 357.920 ;
        RECT 174.820 357.890 175.290 357.950 ;
        RECT 175.760 357.910 176.720 358.080 ;
        RECT 174.820 357.880 175.200 357.890 ;
        RECT 171.430 357.790 171.600 357.840 ;
        RECT 171.400 357.570 171.620 357.790 ;
        RECT 175.030 357.650 175.200 357.880 ;
        RECT 171.430 357.510 171.600 357.570 ;
        RECT 171.950 357.430 172.280 357.610 ;
        RECT 175.030 357.600 175.260 357.650 ;
        RECT 172.530 357.430 174.690 357.600 ;
        RECT 174.930 357.430 175.260 357.600 ;
        RECT 175.550 357.460 175.760 357.790 ;
        RECT 176.000 357.440 176.180 357.730 ;
        RECT 176.540 357.450 176.720 357.910 ;
        RECT 186.410 357.830 186.580 358.250 ;
        RECT 187.220 358.120 187.460 358.160 ;
        RECT 190.000 358.120 190.170 358.130 ;
        RECT 186.890 357.950 187.460 358.120 ;
        RECT 187.700 357.950 189.040 358.120 ;
        RECT 189.490 357.950 190.450 358.120 ;
        RECT 187.220 357.920 187.460 357.950 ;
        RECT 190.980 357.880 191.150 359.610 ;
        RECT 191.380 358.770 191.550 359.660 ;
        RECT 191.380 357.830 191.550 358.720 ;
        RECT 196.490 358.530 197.040 358.960 ;
        RECT 200.520 358.600 201.070 359.030 ;
        RECT 236.110 358.600 236.660 359.030 ;
        RECT 240.140 358.530 240.690 358.960 ;
        RECT 205.010 357.730 205.330 357.770 ;
        RECT 176.730 357.460 177.350 357.630 ;
        RECT 171.980 356.990 172.250 357.430 ;
        RECT 173.460 357.170 173.790 357.430 ;
        RECT 174.410 357.390 174.700 357.430 ;
        RECT 174.370 357.220 174.700 357.390 ;
        RECT 174.410 357.190 174.700 357.220 ;
        RECT 175.000 357.290 175.260 357.430 ;
        RECT 175.400 357.290 176.180 357.440 ;
        RECT 172.020 356.980 172.250 356.990 ;
        RECT 175.000 357.120 176.180 357.290 ;
        RECT 176.460 357.280 176.790 357.450 ;
        RECT 203.410 357.340 203.610 357.690 ;
        RECT 205.000 357.610 205.330 357.730 ;
        RECT 204.890 357.510 205.330 357.610 ;
        RECT 231.850 357.730 232.170 357.770 ;
        RECT 231.850 357.610 232.180 357.730 ;
        RECT 231.850 357.510 232.290 357.610 ;
        RECT 204.890 357.440 205.230 357.510 ;
        RECT 231.950 357.440 232.290 357.510 ;
        RECT 203.400 357.310 203.610 357.340 ;
        RECT 233.570 357.340 233.770 357.690 ;
        RECT 175.000 356.980 175.260 357.120 ;
        RECT 172.020 356.810 172.780 356.980 ;
        RECT 173.030 356.810 174.200 356.980 ;
        RECT 174.440 356.950 175.260 356.980 ;
        RECT 174.440 356.810 175.550 356.950 ;
        RECT 173.430 356.710 173.780 356.810 ;
        RECT 175.090 356.780 175.550 356.810 ;
        RECT 176.000 356.780 177.190 356.950 ;
        RECT 176.040 356.760 177.190 356.780 ;
        RECT 177.020 356.720 177.190 356.760 ;
        RECT 203.400 356.720 203.620 357.310 ;
        RECT 204.140 356.720 204.340 357.320 ;
        RECT 205.010 357.180 205.330 357.220 ;
        RECT 205.000 356.990 205.330 357.180 ;
        RECT 204.890 356.960 205.330 356.990 ;
        RECT 231.850 357.180 232.170 357.220 ;
        RECT 231.850 356.990 232.180 357.180 ;
        RECT 231.850 356.960 232.290 356.990 ;
        RECT 204.890 356.820 205.230 356.960 ;
        RECT 231.950 356.820 232.290 356.960 ;
        RECT 232.840 356.720 233.040 357.320 ;
        RECT 233.570 357.310 233.780 357.340 ;
        RECT 233.560 356.720 233.780 357.310 ;
        RECT 245.070 356.770 245.250 358.820 ;
        RECT 245.800 358.560 246.130 358.730 ;
        RECT 245.880 356.780 246.050 358.560 ;
        RECT 174.820 356.370 175.210 356.420 ;
        RECT 174.470 356.310 175.210 356.370 ;
        RECT 174.470 356.250 175.290 356.310 ;
        RECT 174.480 356.200 175.290 356.250 ;
        RECT 174.820 356.140 175.290 356.200 ;
        RECT 175.760 356.160 176.720 356.330 ;
        RECT 174.820 356.130 175.200 356.140 ;
        RECT 171.430 356.040 171.600 356.090 ;
        RECT 171.400 355.820 171.620 356.040 ;
        RECT 175.030 355.900 175.200 356.130 ;
        RECT 171.430 355.760 171.600 355.820 ;
        RECT 171.950 355.680 172.280 355.860 ;
        RECT 175.030 355.850 175.260 355.900 ;
        RECT 172.530 355.680 174.690 355.850 ;
        RECT 174.930 355.680 175.260 355.850 ;
        RECT 175.550 355.710 175.760 356.040 ;
        RECT 176.000 355.690 176.180 355.980 ;
        RECT 176.540 355.700 176.720 356.160 ;
        RECT 176.730 355.710 177.350 355.880 ;
        RECT 171.980 355.240 172.250 355.680 ;
        RECT 173.460 355.420 173.790 355.680 ;
        RECT 174.410 355.640 174.700 355.680 ;
        RECT 174.370 355.470 174.700 355.640 ;
        RECT 174.410 355.440 174.700 355.470 ;
        RECT 175.000 355.540 175.260 355.680 ;
        RECT 175.400 355.540 176.180 355.690 ;
        RECT 172.020 355.230 172.250 355.240 ;
        RECT 175.000 355.370 176.180 355.540 ;
        RECT 176.460 355.530 176.790 355.700 ;
        RECT 209.040 355.680 209.210 356.210 ;
        RECT 212.980 355.690 213.150 356.220 ;
        RECT 224.030 355.690 224.200 356.220 ;
        RECT 227.970 355.680 228.140 356.210 ;
        RECT 175.000 355.230 175.260 355.370 ;
        RECT 172.020 355.060 172.780 355.230 ;
        RECT 173.030 355.060 174.200 355.230 ;
        RECT 174.440 355.200 175.260 355.230 ;
        RECT 174.440 355.060 175.550 355.200 ;
        RECT 173.430 354.960 173.780 355.060 ;
        RECT 175.090 355.030 175.550 355.060 ;
        RECT 176.000 355.030 177.190 355.200 ;
        RECT 176.040 355.010 177.190 355.030 ;
        RECT 177.020 354.970 177.190 355.010 ;
        RECT 203.400 354.760 203.620 355.350 ;
        RECT 203.400 354.730 203.610 354.760 ;
        RECT 204.140 354.750 204.340 355.350 ;
        RECT 204.890 355.110 205.230 355.250 ;
        RECT 231.950 355.110 232.290 355.250 ;
        RECT 204.890 355.080 205.330 355.110 ;
        RECT 205.000 354.890 205.330 355.080 ;
        RECT 231.850 355.080 232.290 355.110 ;
        RECT 205.010 354.850 205.330 354.890 ;
        RECT 203.410 354.100 203.610 354.730 ;
        RECT 204.890 354.560 205.230 354.630 ;
        RECT 204.890 354.460 205.330 354.560 ;
        RECT 205.000 354.370 205.330 354.460 ;
        RECT 204.890 354.270 205.330 354.370 ;
        RECT 206.670 354.330 207.110 354.500 ;
        RECT 204.890 354.200 205.230 354.270 ;
        RECT 203.400 354.070 203.610 354.100 ;
        RECT 203.400 353.480 203.620 354.070 ;
        RECT 204.140 353.480 204.340 354.080 ;
        RECT 205.010 353.940 205.330 353.980 ;
        RECT 205.000 353.750 205.330 353.940 ;
        RECT 209.040 353.840 209.210 354.850 ;
        RECT 212.970 353.980 213.140 354.990 ;
        RECT 224.040 353.980 224.210 354.990 ;
        RECT 231.850 354.890 232.180 355.080 ;
        RECT 231.850 354.850 232.170 354.890 ;
        RECT 227.970 353.840 228.140 354.850 ;
        RECT 232.840 354.750 233.040 355.350 ;
        RECT 233.560 354.760 233.780 355.350 ;
        RECT 233.570 354.730 233.780 354.760 ;
        RECT 231.950 354.560 232.290 354.630 ;
        RECT 230.070 354.330 230.510 354.500 ;
        RECT 231.850 354.460 232.290 354.560 ;
        RECT 231.850 354.370 232.180 354.460 ;
        RECT 231.850 354.270 232.290 354.370 ;
        RECT 231.950 354.200 232.290 354.270 ;
        RECT 233.570 354.100 233.770 354.730 ;
        RECT 231.850 353.940 232.170 353.980 ;
        RECT 204.890 353.720 205.330 353.750 ;
        RECT 231.850 353.750 232.180 353.940 ;
        RECT 231.850 353.720 232.290 353.750 ;
        RECT 204.890 353.580 205.230 353.720 ;
        RECT 231.950 353.580 232.290 353.720 ;
        RECT 232.840 353.480 233.040 354.080 ;
        RECT 233.570 354.070 233.780 354.100 ;
        RECT 233.560 353.480 233.780 354.070 ;
        RECT 245.070 353.720 245.250 355.770 ;
        RECT 245.800 355.510 246.130 355.680 ;
        RECT 245.880 353.730 246.050 355.510 ;
        RECT 186.390 351.970 186.560 352.390 ;
        RECT 187.200 352.270 187.440 352.300 ;
        RECT 186.870 352.100 187.440 352.270 ;
        RECT 187.680 352.100 189.020 352.270 ;
        RECT 189.470 352.100 190.430 352.270 ;
        RECT 187.200 352.060 187.440 352.100 ;
        RECT 189.980 352.090 190.150 352.100 ;
        RECT 186.320 351.750 186.490 351.790 ;
        RECT 186.260 351.580 186.490 351.750 ;
        RECT 189.610 351.650 189.950 351.830 ;
        RECT 174.820 351.490 175.210 351.540 ;
        RECT 174.470 351.430 175.210 351.490 ;
        RECT 174.470 351.370 175.290 351.430 ;
        RECT 174.480 351.320 175.290 351.370 ;
        RECT 174.820 351.260 175.290 351.320 ;
        RECT 175.760 351.280 176.720 351.450 ;
        RECT 186.320 351.370 186.490 351.580 ;
        RECT 174.820 351.250 175.200 351.260 ;
        RECT 171.430 351.160 171.600 351.210 ;
        RECT 171.400 350.940 171.620 351.160 ;
        RECT 175.030 351.020 175.200 351.250 ;
        RECT 171.430 350.880 171.600 350.940 ;
        RECT 171.950 350.800 172.280 350.980 ;
        RECT 175.030 350.970 175.260 351.020 ;
        RECT 172.530 350.800 174.690 350.970 ;
        RECT 174.930 350.800 175.260 350.970 ;
        RECT 175.550 350.830 175.760 351.160 ;
        RECT 176.000 350.810 176.180 351.100 ;
        RECT 176.540 350.820 176.720 351.280 ;
        RECT 186.260 351.200 186.490 351.370 ;
        RECT 186.560 351.360 186.750 351.590 ;
        RECT 186.850 351.480 187.220 351.650 ;
        RECT 187.680 351.480 190.430 351.650 ;
        RECT 186.850 351.300 187.220 351.470 ;
        RECT 187.680 351.300 190.430 351.470 ;
        RECT 186.320 351.160 186.490 351.200 ;
        RECT 189.610 351.120 189.950 351.300 ;
        RECT 176.730 350.830 177.350 351.000 ;
        RECT 171.980 350.360 172.250 350.800 ;
        RECT 173.460 350.540 173.790 350.800 ;
        RECT 174.410 350.760 174.700 350.800 ;
        RECT 174.370 350.590 174.700 350.760 ;
        RECT 174.410 350.560 174.700 350.590 ;
        RECT 175.000 350.660 175.260 350.800 ;
        RECT 175.400 350.660 176.180 350.810 ;
        RECT 172.020 350.350 172.250 350.360 ;
        RECT 175.000 350.490 176.180 350.660 ;
        RECT 176.460 350.650 176.790 350.820 ;
        RECT 186.390 350.560 186.560 350.980 ;
        RECT 187.200 350.850 187.440 350.890 ;
        RECT 189.980 350.850 190.150 350.860 ;
        RECT 186.870 350.680 187.440 350.850 ;
        RECT 187.680 350.680 189.020 350.850 ;
        RECT 189.470 350.680 190.430 350.850 ;
        RECT 187.200 350.650 187.440 350.680 ;
        RECT 190.960 350.610 191.130 352.340 ;
        RECT 191.360 351.500 191.530 352.390 ;
        RECT 203.400 351.530 203.620 352.120 ;
        RECT 203.400 351.500 203.610 351.530 ;
        RECT 204.140 351.520 204.340 352.120 ;
        RECT 204.890 351.880 205.230 352.020 ;
        RECT 231.950 351.880 232.290 352.020 ;
        RECT 204.890 351.850 205.330 351.880 ;
        RECT 205.000 351.660 205.330 351.850 ;
        RECT 205.010 351.620 205.330 351.660 ;
        RECT 231.850 351.850 232.290 351.880 ;
        RECT 231.850 351.660 232.180 351.850 ;
        RECT 231.850 351.620 232.170 351.660 ;
        RECT 232.840 351.520 233.040 352.120 ;
        RECT 233.560 351.530 233.780 352.120 ;
        RECT 191.360 350.560 191.530 351.450 ;
        RECT 203.410 351.150 203.610 351.500 ;
        RECT 233.570 351.500 233.780 351.530 ;
        RECT 204.890 351.330 205.230 351.400 ;
        RECT 231.950 351.330 232.290 351.400 ;
        RECT 204.890 351.230 205.330 351.330 ;
        RECT 205.000 351.110 205.330 351.230 ;
        RECT 205.010 351.070 205.330 351.110 ;
        RECT 231.850 351.230 232.290 351.330 ;
        RECT 231.850 351.110 232.180 351.230 ;
        RECT 233.570 351.150 233.770 351.500 ;
        RECT 231.850 351.070 232.170 351.110 ;
        RECT 175.000 350.350 175.260 350.490 ;
        RECT 172.020 350.180 172.780 350.350 ;
        RECT 173.030 350.180 174.200 350.350 ;
        RECT 174.440 350.320 175.260 350.350 ;
        RECT 174.440 350.180 175.550 350.320 ;
        RECT 173.430 350.080 173.780 350.180 ;
        RECT 175.090 350.150 175.550 350.180 ;
        RECT 176.000 350.150 177.190 350.320 ;
        RECT 176.040 350.130 177.190 350.150 ;
        RECT 177.020 350.090 177.190 350.130 ;
        RECT 174.820 349.740 175.210 349.790 ;
        RECT 174.470 349.680 175.210 349.740 ;
        RECT 174.470 349.620 175.290 349.680 ;
        RECT 174.480 349.570 175.290 349.620 ;
        RECT 174.820 349.510 175.290 349.570 ;
        RECT 175.760 349.530 176.720 349.700 ;
        RECT 197.090 349.650 197.640 350.080 ;
        RECT 201.120 349.720 201.670 350.150 ;
        RECT 174.820 349.500 175.200 349.510 ;
        RECT 171.430 349.410 171.600 349.460 ;
        RECT 171.400 349.190 171.620 349.410 ;
        RECT 175.030 349.270 175.200 349.500 ;
        RECT 171.430 349.130 171.600 349.190 ;
        RECT 171.950 349.050 172.280 349.230 ;
        RECT 175.030 349.220 175.260 349.270 ;
        RECT 172.530 349.050 174.690 349.220 ;
        RECT 174.930 349.050 175.260 349.220 ;
        RECT 175.550 349.080 175.760 349.410 ;
        RECT 176.000 349.060 176.180 349.350 ;
        RECT 176.540 349.070 176.720 349.530 ;
        RECT 176.730 349.080 177.350 349.250 ;
        RECT 171.980 348.610 172.250 349.050 ;
        RECT 173.460 348.790 173.790 349.050 ;
        RECT 174.410 349.010 174.700 349.050 ;
        RECT 174.370 348.840 174.700 349.010 ;
        RECT 174.410 348.810 174.700 348.840 ;
        RECT 175.000 348.910 175.260 349.050 ;
        RECT 175.400 348.910 176.180 349.060 ;
        RECT 172.020 348.600 172.250 348.610 ;
        RECT 175.000 348.740 176.180 348.910 ;
        RECT 176.460 348.900 176.790 349.070 ;
        RECT 186.390 348.770 186.560 349.190 ;
        RECT 187.200 349.070 187.440 349.100 ;
        RECT 186.870 348.900 187.440 349.070 ;
        RECT 187.680 348.900 189.020 349.070 ;
        RECT 189.470 348.900 190.430 349.070 ;
        RECT 187.200 348.860 187.440 348.900 ;
        RECT 189.980 348.890 190.150 348.900 ;
        RECT 175.000 348.600 175.260 348.740 ;
        RECT 172.020 348.430 172.780 348.600 ;
        RECT 173.030 348.430 174.200 348.600 ;
        RECT 174.440 348.570 175.260 348.600 ;
        RECT 174.440 348.430 175.550 348.570 ;
        RECT 173.430 348.330 173.780 348.430 ;
        RECT 175.090 348.400 175.550 348.430 ;
        RECT 176.000 348.400 177.190 348.570 ;
        RECT 186.320 348.550 186.490 348.590 ;
        RECT 176.040 348.380 177.190 348.400 ;
        RECT 186.260 348.380 186.490 348.550 ;
        RECT 189.610 348.450 189.950 348.630 ;
        RECT 177.020 348.340 177.190 348.380 ;
        RECT 186.320 348.170 186.490 348.380 ;
        RECT 174.820 347.990 175.210 348.040 ;
        RECT 186.260 348.000 186.490 348.170 ;
        RECT 186.560 348.160 186.750 348.390 ;
        RECT 186.850 348.280 187.220 348.450 ;
        RECT 187.680 348.280 190.430 348.450 ;
        RECT 186.850 348.100 187.220 348.270 ;
        RECT 187.680 348.100 190.430 348.270 ;
        RECT 174.470 347.930 175.210 347.990 ;
        RECT 186.320 347.960 186.490 348.000 ;
        RECT 174.470 347.870 175.290 347.930 ;
        RECT 174.480 347.820 175.290 347.870 ;
        RECT 174.820 347.760 175.290 347.820 ;
        RECT 175.760 347.780 176.720 347.950 ;
        RECT 189.610 347.920 189.950 348.100 ;
        RECT 174.820 347.750 175.200 347.760 ;
        RECT 171.430 347.660 171.600 347.710 ;
        RECT 31.090 347.540 31.610 347.560 ;
        RECT 25.040 346.060 30.750 346.070 ;
        RECT 24.960 345.890 30.750 346.060 ;
        RECT 25.050 345.880 30.750 345.890 ;
        RECT 30.520 345.810 30.690 345.880 ;
        RECT 31.090 345.760 31.620 347.540 ;
        RECT 171.400 347.440 171.620 347.660 ;
        RECT 175.030 347.520 175.200 347.750 ;
        RECT 171.430 347.380 171.600 347.440 ;
        RECT 171.950 347.300 172.280 347.480 ;
        RECT 175.030 347.470 175.260 347.520 ;
        RECT 172.530 347.300 174.690 347.470 ;
        RECT 174.930 347.300 175.260 347.470 ;
        RECT 175.550 347.330 175.760 347.660 ;
        RECT 176.000 347.310 176.180 347.600 ;
        RECT 176.540 347.320 176.720 347.780 ;
        RECT 176.730 347.330 177.350 347.500 ;
        RECT 186.390 347.360 186.560 347.780 ;
        RECT 187.200 347.650 187.440 347.690 ;
        RECT 189.980 347.650 190.150 347.660 ;
        RECT 186.870 347.480 187.440 347.650 ;
        RECT 187.680 347.480 189.020 347.650 ;
        RECT 189.470 347.480 190.430 347.650 ;
        RECT 187.200 347.450 187.440 347.480 ;
        RECT 190.960 347.410 191.130 349.140 ;
        RECT 191.360 348.300 191.530 349.190 ;
        RECT 205.610 348.890 205.930 348.930 ;
        RECT 204.010 348.500 204.210 348.850 ;
        RECT 205.600 348.770 205.930 348.890 ;
        RECT 205.490 348.670 205.930 348.770 ;
        RECT 205.490 348.600 205.830 348.670 ;
        RECT 204.000 348.470 204.210 348.500 ;
        RECT 191.360 347.360 191.530 348.250 ;
        RECT 204.000 347.880 204.220 348.470 ;
        RECT 204.740 347.880 204.940 348.480 ;
        RECT 205.610 348.340 205.930 348.380 ;
        RECT 205.600 348.150 205.930 348.340 ;
        RECT 205.490 348.120 205.930 348.150 ;
        RECT 205.490 347.980 205.830 348.120 ;
        RECT 171.980 346.860 172.250 347.300 ;
        RECT 173.460 347.040 173.790 347.300 ;
        RECT 174.410 347.260 174.700 347.300 ;
        RECT 174.370 347.090 174.700 347.260 ;
        RECT 174.410 347.060 174.700 347.090 ;
        RECT 175.000 347.160 175.260 347.300 ;
        RECT 175.400 347.160 176.180 347.310 ;
        RECT 172.020 346.850 172.250 346.860 ;
        RECT 175.000 346.990 176.180 347.160 ;
        RECT 176.460 347.150 176.790 347.320 ;
        RECT 175.000 346.850 175.260 346.990 ;
        RECT 172.020 346.680 172.780 346.850 ;
        RECT 173.030 346.680 174.200 346.850 ;
        RECT 174.440 346.820 175.260 346.850 ;
        RECT 174.440 346.680 175.550 346.820 ;
        RECT 173.430 346.580 173.780 346.680 ;
        RECT 175.090 346.650 175.550 346.680 ;
        RECT 176.000 346.650 177.190 346.820 ;
        RECT 209.770 346.780 209.940 347.310 ;
        RECT 213.790 346.810 213.960 347.340 ;
        RECT 176.040 346.630 177.190 346.650 ;
        RECT 177.020 346.590 177.190 346.630 ;
        RECT 174.820 346.240 175.210 346.290 ;
        RECT 174.470 346.180 175.210 346.240 ;
        RECT 174.470 346.120 175.290 346.180 ;
        RECT 174.480 346.070 175.290 346.120 ;
        RECT 174.820 346.010 175.290 346.070 ;
        RECT 175.760 346.030 176.720 346.200 ;
        RECT 174.820 346.000 175.200 346.010 ;
        RECT 171.430 345.910 171.600 345.960 ;
        RECT 31.100 345.740 31.620 345.760 ;
        RECT 24.080 345.020 26.520 345.310 ;
        RECT 31.100 345.230 31.610 345.740 ;
        RECT 171.400 345.690 171.620 345.910 ;
        RECT 175.030 345.770 175.200 346.000 ;
        RECT 171.430 345.630 171.600 345.690 ;
        RECT 171.950 345.550 172.280 345.730 ;
        RECT 175.030 345.720 175.260 345.770 ;
        RECT 172.530 345.550 174.690 345.720 ;
        RECT 174.930 345.550 175.260 345.720 ;
        RECT 175.550 345.580 175.760 345.910 ;
        RECT 176.000 345.560 176.180 345.850 ;
        RECT 176.540 345.570 176.720 346.030 ;
        RECT 204.000 345.940 204.220 346.530 ;
        RECT 204.000 345.910 204.210 345.940 ;
        RECT 204.740 345.930 204.940 346.530 ;
        RECT 205.490 346.290 205.830 346.430 ;
        RECT 205.490 346.260 205.930 346.290 ;
        RECT 205.600 346.070 205.930 346.260 ;
        RECT 205.610 346.030 205.930 346.070 ;
        RECT 176.730 345.580 177.350 345.750 ;
        RECT 31.100 345.020 31.630 345.230 ;
        RECT 171.980 345.110 172.250 345.550 ;
        RECT 173.460 345.290 173.790 345.550 ;
        RECT 174.410 345.510 174.700 345.550 ;
        RECT 174.370 345.340 174.700 345.510 ;
        RECT 174.410 345.310 174.700 345.340 ;
        RECT 175.000 345.410 175.260 345.550 ;
        RECT 175.400 345.410 176.180 345.560 ;
        RECT 24.080 344.540 31.630 345.020 ;
        RECT 172.020 345.100 172.250 345.110 ;
        RECT 175.000 345.240 176.180 345.410 ;
        RECT 176.460 345.400 176.790 345.570 ;
        RECT 204.010 345.260 204.210 345.910 ;
        RECT 205.490 345.740 205.830 345.810 ;
        RECT 205.490 345.640 205.930 345.740 ;
        RECT 205.600 345.530 205.930 345.640 ;
        RECT 205.490 345.430 205.930 345.530 ;
        RECT 207.270 345.510 207.710 345.680 ;
        RECT 205.490 345.360 205.830 345.430 ;
        RECT 175.000 345.100 175.260 345.240 ;
        RECT 172.020 344.930 172.780 345.100 ;
        RECT 173.030 344.930 174.200 345.100 ;
        RECT 174.440 345.070 175.260 345.100 ;
        RECT 204.000 345.230 204.210 345.260 ;
        RECT 174.440 344.930 175.550 345.070 ;
        RECT 173.430 344.830 173.780 344.930 ;
        RECT 175.090 344.900 175.550 344.930 ;
        RECT 176.000 344.900 177.190 345.070 ;
        RECT 176.040 344.880 177.190 344.900 ;
        RECT 177.020 344.840 177.190 344.880 ;
        RECT 204.000 344.640 204.220 345.230 ;
        RECT 204.740 344.640 204.940 345.240 ;
        RECT 205.610 345.100 205.930 345.140 ;
        RECT 205.600 344.910 205.930 345.100 ;
        RECT 209.760 344.920 209.930 346.110 ;
        RECT 205.490 344.880 205.930 344.910 ;
        RECT 213.780 344.880 213.950 346.050 ;
        RECT 205.490 344.740 205.830 344.880 ;
        RECT 24.080 344.510 31.440 344.540 ;
        RECT 24.080 342.750 31.610 343.300 ;
        RECT 22.390 329.780 23.870 330.030 ;
        RECT 24.080 329.840 24.590 342.750 ;
        RECT 30.940 342.740 31.610 342.750 ;
        RECT 27.240 341.850 30.700 342.290 ;
        RECT 25.310 341.750 30.700 341.850 ;
        RECT 25.310 341.680 30.590 341.750 ;
        RECT 25.310 330.770 25.480 341.680 ;
        RECT 25.810 341.270 30.040 341.290 ;
        RECT 25.790 331.160 30.120 341.270 ;
        RECT 25.850 331.110 26.020 331.160 ;
        RECT 30.420 330.770 30.590 341.680 ;
        RECT 25.310 330.600 30.590 330.770 ;
        RECT 30.350 330.590 30.590 330.600 ;
        RECT 31.100 329.840 31.610 342.740 ;
        RECT 151.720 342.860 152.040 342.890 ;
        RECT 152.370 342.860 152.690 342.890 ;
        RECT 151.720 342.670 152.050 342.860 ;
        RECT 152.370 342.670 152.700 342.860 ;
        RECT 186.420 342.700 186.590 343.120 ;
        RECT 187.230 343.000 187.470 343.030 ;
        RECT 186.900 342.830 187.470 343.000 ;
        RECT 187.710 342.830 189.050 343.000 ;
        RECT 189.500 342.830 190.460 343.000 ;
        RECT 187.230 342.790 187.470 342.830 ;
        RECT 190.010 342.820 190.180 342.830 ;
        RECT 150.630 342.450 150.800 342.650 ;
        RECT 151.180 342.450 151.350 342.650 ;
        RECT 151.720 342.630 152.040 342.670 ;
        RECT 152.370 342.630 152.690 342.670 ;
        RECT 150.500 342.420 150.820 342.450 ;
        RECT 151.180 342.420 151.520 342.450 ;
        RECT 150.500 342.230 150.830 342.420 ;
        RECT 151.180 342.230 151.530 342.420 ;
        RECT 150.500 342.190 150.820 342.230 ;
        RECT 151.180 342.190 151.520 342.230 ;
        RECT 149.880 340.620 150.050 340.640 ;
        RECT 149.860 340.500 150.070 340.620 ;
        RECT 149.860 340.190 150.260 340.500 ;
        RECT 150.630 340.250 150.800 342.190 ;
        RECT 151.180 340.250 151.350 342.190 ;
        RECT 151.820 340.250 151.990 342.630 ;
        RECT 152.370 340.630 152.540 342.630 ;
        RECT 186.350 342.480 186.520 342.520 ;
        RECT 174.780 342.430 175.170 342.480 ;
        RECT 174.430 342.370 175.170 342.430 ;
        RECT 174.430 342.310 175.250 342.370 ;
        RECT 174.440 342.260 175.250 342.310 ;
        RECT 174.780 342.200 175.250 342.260 ;
        RECT 175.720 342.220 176.680 342.390 ;
        RECT 186.290 342.310 186.520 342.480 ;
        RECT 189.640 342.380 189.980 342.560 ;
        RECT 174.780 342.190 175.160 342.200 ;
        RECT 152.800 341.330 152.970 342.180 ;
        RECT 171.390 342.100 171.560 342.150 ;
        RECT 171.360 341.880 171.580 342.100 ;
        RECT 174.990 341.960 175.160 342.190 ;
        RECT 171.390 341.820 171.560 341.880 ;
        RECT 171.910 341.740 172.240 341.920 ;
        RECT 174.990 341.910 175.220 341.960 ;
        RECT 172.490 341.740 174.650 341.910 ;
        RECT 174.890 341.740 175.220 341.910 ;
        RECT 175.510 341.770 175.720 342.100 ;
        RECT 175.960 341.750 176.140 342.040 ;
        RECT 176.500 341.760 176.680 342.220 ;
        RECT 186.350 342.100 186.520 342.310 ;
        RECT 176.690 341.770 177.310 341.940 ;
        RECT 186.290 341.930 186.520 342.100 ;
        RECT 186.590 342.090 186.780 342.320 ;
        RECT 186.880 342.210 187.250 342.380 ;
        RECT 187.710 342.210 190.460 342.380 ;
        RECT 186.880 342.030 187.250 342.200 ;
        RECT 187.710 342.030 190.460 342.200 ;
        RECT 186.350 341.890 186.520 341.930 ;
        RECT 189.640 341.850 189.980 342.030 ;
        RECT 171.940 341.300 172.210 341.740 ;
        RECT 173.420 341.480 173.750 341.740 ;
        RECT 174.370 341.700 174.660 341.740 ;
        RECT 174.330 341.530 174.660 341.700 ;
        RECT 174.370 341.500 174.660 341.530 ;
        RECT 174.960 341.600 175.220 341.740 ;
        RECT 175.360 341.600 176.140 341.750 ;
        RECT 171.980 341.290 172.210 341.300 ;
        RECT 174.960 341.430 176.140 341.600 ;
        RECT 176.420 341.590 176.750 341.760 ;
        RECT 174.960 341.290 175.220 341.430 ;
        RECT 186.420 341.290 186.590 341.710 ;
        RECT 187.230 341.580 187.470 341.620 ;
        RECT 190.010 341.580 190.180 341.590 ;
        RECT 186.900 341.410 187.470 341.580 ;
        RECT 187.710 341.410 189.050 341.580 ;
        RECT 189.500 341.410 190.460 341.580 ;
        RECT 187.230 341.380 187.470 341.410 ;
        RECT 190.990 341.340 191.160 343.070 ;
        RECT 191.390 342.230 191.560 343.120 ;
        RECT 204.000 342.690 204.220 343.280 ;
        RECT 204.000 342.660 204.210 342.690 ;
        RECT 204.740 342.680 204.940 343.280 ;
        RECT 221.610 343.240 221.820 343.260 ;
        RECT 205.490 343.040 205.830 343.180 ;
        RECT 221.590 343.070 222.260 343.240 ;
        RECT 205.490 343.010 205.930 343.040 ;
        RECT 205.600 342.820 205.930 343.010 ;
        RECT 205.610 342.780 205.930 342.820 ;
        RECT 220.820 342.950 221.140 342.990 ;
        RECT 220.820 342.860 221.150 342.950 ;
        RECT 221.590 342.860 221.840 343.070 ;
        RECT 220.820 342.840 222.320 342.860 ;
        RECT 220.820 342.740 222.400 342.840 ;
        RECT 220.670 342.690 222.400 342.740 ;
        RECT 204.010 342.310 204.210 342.660 ;
        RECT 205.490 342.490 205.830 342.560 ;
        RECT 220.670 342.520 221.340 342.690 ;
        RECT 221.510 342.670 221.840 342.690 ;
        RECT 222.060 342.670 222.400 342.690 ;
        RECT 205.490 342.390 205.930 342.490 ;
        RECT 220.670 342.480 220.990 342.520 ;
        RECT 205.600 342.270 205.930 342.390 ;
        RECT 205.610 342.230 205.930 342.270 ;
        RECT 220.670 342.270 220.990 342.310 ;
        RECT 221.000 342.270 221.340 342.520 ;
        RECT 221.590 342.500 221.760 342.670 ;
        RECT 222.150 342.500 222.320 342.670 ;
        RECT 221.510 342.290 221.840 342.500 ;
        RECT 222.060 342.290 222.400 342.500 ;
        RECT 191.390 341.290 191.560 342.180 ;
        RECT 220.670 342.100 221.340 342.270 ;
        RECT 221.590 342.120 221.760 342.290 ;
        RECT 222.150 342.120 222.320 342.290 ;
        RECT 221.510 342.100 221.840 342.120 ;
        RECT 222.060 342.100 222.400 342.120 ;
        RECT 220.670 342.050 222.400 342.100 ;
        RECT 220.820 341.950 222.400 342.050 ;
        RECT 220.820 341.930 222.320 341.950 ;
        RECT 220.820 341.840 221.150 341.930 ;
        RECT 220.820 341.800 221.140 341.840 ;
        RECT 221.590 341.720 221.840 341.930 ;
        RECT 222.720 341.870 223.230 342.920 ;
        RECT 221.590 341.550 222.260 341.720 ;
        RECT 221.610 341.530 221.820 341.550 ;
        RECT 171.980 341.120 172.740 341.290 ;
        RECT 172.990 341.120 174.160 341.290 ;
        RECT 174.400 341.260 175.220 341.290 ;
        RECT 174.400 341.120 175.510 341.260 ;
        RECT 173.390 341.020 173.740 341.120 ;
        RECT 175.050 341.090 175.510 341.120 ;
        RECT 175.960 341.090 177.150 341.260 ;
        RECT 176.000 341.070 177.150 341.090 ;
        RECT 176.980 341.030 177.150 341.070 ;
        RECT 174.780 340.680 175.170 340.730 ;
        RECT 152.370 340.610 152.860 340.630 ;
        RECT 174.430 340.620 175.170 340.680 ;
        RECT 152.370 340.440 152.880 340.610 ;
        RECT 174.430 340.560 175.250 340.620 ;
        RECT 174.440 340.510 175.250 340.560 ;
        RECT 174.780 340.450 175.250 340.510 ;
        RECT 175.720 340.470 176.680 340.640 ;
        RECT 221.610 340.470 221.820 340.490 ;
        RECT 174.780 340.440 175.160 340.450 ;
        RECT 152.370 340.420 152.860 340.440 ;
        RECT 152.370 340.250 152.540 340.420 ;
        RECT 171.390 340.350 171.560 340.400 ;
        RECT 150.050 340.070 150.260 340.190 ;
        RECT 171.360 340.130 171.580 340.350 ;
        RECT 174.990 340.210 175.160 340.440 ;
        RECT 152.440 340.070 152.870 340.090 ;
        RECT 171.390 340.070 171.560 340.130 ;
        RECT 150.070 340.050 150.240 340.070 ;
        RECT 152.440 339.900 152.890 340.070 ;
        RECT 171.910 339.990 172.240 340.170 ;
        RECT 174.990 340.160 175.220 340.210 ;
        RECT 172.490 339.990 174.650 340.160 ;
        RECT 174.890 339.990 175.220 340.160 ;
        RECT 175.510 340.020 175.720 340.350 ;
        RECT 175.960 340.000 176.140 340.290 ;
        RECT 176.500 340.010 176.680 340.470 ;
        RECT 221.590 340.300 222.260 340.470 ;
        RECT 176.690 340.020 177.310 340.190 ;
        RECT 220.820 340.180 221.140 340.220 ;
        RECT 220.820 340.090 221.150 340.180 ;
        RECT 221.590 340.090 221.840 340.300 ;
        RECT 220.820 340.070 222.320 340.090 ;
        RECT 152.440 339.880 152.870 339.900 ;
        RECT 147.450 338.100 147.960 338.280 ;
        RECT 147.390 338.070 147.960 338.100 ;
        RECT 147.380 337.880 147.960 338.070 ;
        RECT 147.390 337.840 147.960 337.880 ;
        RECT 144.080 337.630 144.400 337.660 ;
        RECT 145.180 337.640 145.500 337.670 ;
        RECT 146.270 337.640 146.590 337.670 ;
        RECT 144.070 337.570 144.400 337.630 ;
        RECT 145.170 337.570 145.500 337.640 ;
        RECT 142.640 335.170 142.810 337.570 ;
        RECT 143.190 335.170 143.360 337.570 ;
        RECT 143.740 335.170 143.910 337.570 ;
        RECT 144.070 337.440 144.460 337.570 ;
        RECT 144.080 337.400 144.460 337.440 ;
        RECT 144.290 335.100 144.460 337.400 ;
        RECT 144.840 336.990 145.010 337.570 ;
        RECT 145.170 337.450 145.560 337.570 ;
        RECT 146.260 337.450 146.590 337.640 ;
        RECT 147.450 337.630 147.960 337.840 ;
        RECT 147.400 337.600 147.960 337.630 ;
        RECT 145.180 337.410 145.560 337.450 ;
        RECT 146.270 337.410 146.590 337.450 ;
        RECT 147.390 337.410 147.970 337.600 ;
        RECT 144.630 336.960 145.010 336.990 ;
        RECT 144.620 336.770 145.010 336.960 ;
        RECT 144.630 336.730 145.010 336.770 ;
        RECT 144.840 335.620 145.010 336.730 ;
        RECT 144.630 335.590 145.010 335.620 ;
        RECT 144.620 335.400 145.010 335.590 ;
        RECT 144.630 335.360 145.010 335.400 ;
        RECT 144.840 335.100 145.010 335.360 ;
        RECT 145.390 335.100 145.560 337.410 ;
        RECT 147.400 337.370 147.970 337.410 ;
        RECT 147.460 337.270 147.970 337.370 ;
        RECT 149.050 337.330 149.220 339.820 ;
        RECT 149.600 337.330 149.770 339.830 ;
        RECT 150.230 337.330 150.400 339.820 ;
        RECT 150.780 338.570 150.950 339.830 ;
        RECT 171.940 339.550 172.210 339.990 ;
        RECT 173.420 339.730 173.750 339.990 ;
        RECT 174.370 339.950 174.660 339.990 ;
        RECT 174.330 339.780 174.660 339.950 ;
        RECT 174.370 339.750 174.660 339.780 ;
        RECT 174.960 339.850 175.220 339.990 ;
        RECT 175.360 339.850 176.140 340.000 ;
        RECT 171.980 339.540 172.210 339.550 ;
        RECT 174.960 339.680 176.140 339.850 ;
        RECT 176.420 339.840 176.750 340.010 ;
        RECT 220.820 339.970 222.400 340.070 ;
        RECT 220.670 339.920 222.400 339.970 ;
        RECT 174.960 339.540 175.220 339.680 ;
        RECT 152.790 338.780 152.960 339.450 ;
        RECT 171.980 339.370 172.740 339.540 ;
        RECT 172.990 339.370 174.160 339.540 ;
        RECT 174.400 339.510 175.220 339.540 ;
        RECT 174.400 339.370 175.510 339.510 ;
        RECT 173.390 339.270 173.740 339.370 ;
        RECT 175.050 339.340 175.510 339.370 ;
        RECT 175.960 339.340 177.150 339.510 ;
        RECT 186.420 339.500 186.590 339.920 ;
        RECT 187.230 339.800 187.470 339.830 ;
        RECT 186.900 339.630 187.470 339.800 ;
        RECT 187.710 339.630 189.050 339.800 ;
        RECT 189.500 339.630 190.460 339.800 ;
        RECT 187.230 339.590 187.470 339.630 ;
        RECT 190.010 339.620 190.180 339.630 ;
        RECT 176.000 339.320 177.150 339.340 ;
        RECT 176.980 339.280 177.150 339.320 ;
        RECT 186.350 339.280 186.520 339.320 ;
        RECT 186.290 339.110 186.520 339.280 ;
        RECT 189.640 339.180 189.980 339.360 ;
        RECT 174.780 338.930 175.170 338.980 ;
        RECT 174.430 338.870 175.170 338.930 ;
        RECT 186.350 338.900 186.520 339.110 ;
        RECT 174.430 338.810 175.250 338.870 ;
        RECT 174.440 338.760 175.250 338.810 ;
        RECT 174.780 338.700 175.250 338.760 ;
        RECT 175.720 338.720 176.680 338.890 ;
        RECT 186.290 338.730 186.520 338.900 ;
        RECT 186.590 338.890 186.780 339.120 ;
        RECT 186.880 339.010 187.250 339.180 ;
        RECT 187.710 339.010 190.460 339.180 ;
        RECT 186.880 338.830 187.250 339.000 ;
        RECT 187.710 338.830 190.460 339.000 ;
        RECT 174.780 338.690 175.160 338.700 ;
        RECT 171.390 338.600 171.560 338.650 ;
        RECT 150.530 338.310 150.950 338.570 ;
        RECT 150.780 337.330 150.950 338.310 ;
        RECT 151.220 338.530 151.540 338.560 ;
        RECT 151.220 338.340 151.550 338.530 ;
        RECT 171.360 338.380 171.580 338.600 ;
        RECT 174.990 338.460 175.160 338.690 ;
        RECT 151.220 338.300 151.540 338.340 ;
        RECT 171.390 338.320 171.560 338.380 ;
        RECT 171.910 338.240 172.240 338.420 ;
        RECT 174.990 338.410 175.220 338.460 ;
        RECT 172.490 338.240 174.650 338.410 ;
        RECT 174.890 338.240 175.220 338.410 ;
        RECT 175.510 338.270 175.720 338.600 ;
        RECT 175.960 338.250 176.140 338.540 ;
        RECT 176.500 338.260 176.680 338.720 ;
        RECT 186.350 338.690 186.520 338.730 ;
        RECT 189.640 338.650 189.980 338.830 ;
        RECT 176.690 338.270 177.310 338.440 ;
        RECT 171.940 337.800 172.210 338.240 ;
        RECT 173.420 337.980 173.750 338.240 ;
        RECT 174.370 338.200 174.660 338.240 ;
        RECT 174.330 338.030 174.660 338.200 ;
        RECT 174.370 338.000 174.660 338.030 ;
        RECT 174.960 338.100 175.220 338.240 ;
        RECT 175.360 338.100 176.140 338.250 ;
        RECT 171.980 337.790 172.210 337.800 ;
        RECT 174.960 337.930 176.140 338.100 ;
        RECT 176.420 338.090 176.750 338.260 ;
        RECT 186.420 338.090 186.590 338.510 ;
        RECT 187.230 338.380 187.470 338.420 ;
        RECT 190.010 338.380 190.180 338.390 ;
        RECT 186.900 338.210 187.470 338.380 ;
        RECT 187.710 338.210 189.050 338.380 ;
        RECT 189.500 338.210 190.460 338.380 ;
        RECT 187.230 338.180 187.470 338.210 ;
        RECT 190.990 338.140 191.160 339.870 ;
        RECT 191.390 339.030 191.560 339.920 ;
        RECT 220.670 339.750 221.340 339.920 ;
        RECT 221.510 339.900 221.840 339.920 ;
        RECT 222.060 339.900 222.400 339.920 ;
        RECT 220.670 339.710 220.990 339.750 ;
        RECT 220.670 339.500 220.990 339.540 ;
        RECT 221.000 339.500 221.340 339.750 ;
        RECT 221.590 339.730 221.760 339.900 ;
        RECT 222.150 339.730 222.320 339.900 ;
        RECT 221.510 339.520 221.840 339.730 ;
        RECT 222.060 339.520 222.400 339.730 ;
        RECT 208.690 339.370 209.010 339.410 ;
        RECT 208.690 339.200 209.020 339.370 ;
        RECT 220.670 339.330 221.340 339.500 ;
        RECT 221.590 339.350 221.760 339.520 ;
        RECT 222.150 339.350 222.320 339.520 ;
        RECT 221.510 339.330 221.840 339.350 ;
        RECT 222.060 339.330 222.400 339.350 ;
        RECT 220.670 339.280 222.400 339.330 ;
        RECT 208.600 339.180 209.020 339.200 ;
        RECT 220.820 339.180 222.400 339.280 ;
        RECT 208.600 339.150 209.010 339.180 ;
        RECT 220.820 339.160 222.320 339.180 ;
        RECT 191.390 338.090 191.560 338.980 ;
        RECT 208.600 338.450 208.780 339.150 ;
        RECT 220.820 339.070 221.150 339.160 ;
        RECT 220.820 339.030 221.140 339.070 ;
        RECT 221.590 338.950 221.840 339.160 ;
        RECT 222.720 339.100 223.230 340.150 ;
        RECT 221.590 338.780 222.260 338.950 ;
        RECT 221.610 338.760 221.820 338.780 ;
        RECT 208.600 338.410 209.060 338.450 ;
        RECT 208.600 338.280 209.070 338.410 ;
        RECT 208.740 338.220 209.070 338.280 ;
        RECT 208.740 338.190 209.060 338.220 ;
        RECT 174.960 337.790 175.220 337.930 ;
        RECT 151.700 337.760 152.020 337.790 ;
        RECT 151.700 337.570 152.030 337.760 ;
        RECT 152.410 337.700 152.730 337.730 ;
        RECT 151.700 337.530 152.020 337.570 ;
        RECT 152.410 337.510 152.740 337.700 ;
        RECT 171.980 337.620 172.740 337.790 ;
        RECT 172.990 337.620 174.160 337.790 ;
        RECT 174.400 337.760 175.220 337.790 ;
        RECT 174.400 337.620 175.510 337.760 ;
        RECT 173.390 337.520 173.740 337.620 ;
        RECT 175.050 337.590 175.510 337.620 ;
        RECT 175.960 337.590 177.150 337.760 ;
        RECT 176.000 337.570 177.150 337.590 ;
        RECT 176.980 337.530 177.150 337.570 ;
        RECT 152.410 337.470 152.730 337.510 ;
        RECT 174.780 337.180 175.170 337.230 ;
        RECT 174.430 337.120 175.170 337.180 ;
        RECT 145.730 336.960 146.050 336.990 ;
        RECT 146.830 336.960 147.150 336.990 ;
        RECT 145.720 336.770 146.050 336.960 ;
        RECT 146.820 336.770 147.150 336.960 ;
        RECT 145.730 336.730 146.050 336.770 ;
        RECT 146.830 336.730 147.150 336.770 ;
        RECT 147.750 335.860 147.920 337.080 ;
        RECT 174.430 337.060 175.250 337.120 ;
        RECT 174.440 337.010 175.250 337.060 ;
        RECT 174.780 336.950 175.250 337.010 ;
        RECT 175.720 336.970 176.680 337.140 ;
        RECT 174.780 336.940 175.160 336.950 ;
        RECT 171.390 336.850 171.560 336.900 ;
        RECT 171.360 336.630 171.580 336.850 ;
        RECT 174.990 336.710 175.160 336.940 ;
        RECT 171.390 336.570 171.560 336.630 ;
        RECT 171.910 336.490 172.240 336.670 ;
        RECT 174.990 336.660 175.220 336.710 ;
        RECT 172.490 336.490 174.650 336.660 ;
        RECT 174.890 336.490 175.220 336.660 ;
        RECT 175.510 336.520 175.720 336.850 ;
        RECT 175.960 336.500 176.140 336.790 ;
        RECT 176.500 336.510 176.680 336.970 ;
        RECT 176.690 336.520 177.310 336.690 ;
        RECT 171.940 336.050 172.210 336.490 ;
        RECT 173.420 336.230 173.750 336.490 ;
        RECT 174.370 336.450 174.660 336.490 ;
        RECT 174.330 336.280 174.660 336.450 ;
        RECT 174.370 336.250 174.660 336.280 ;
        RECT 174.960 336.350 175.220 336.490 ;
        RECT 175.360 336.350 176.140 336.500 ;
        RECT 171.980 336.040 172.210 336.050 ;
        RECT 174.960 336.180 176.140 336.350 ;
        RECT 176.420 336.340 176.750 336.510 ;
        RECT 174.960 336.040 175.220 336.180 ;
        RECT 171.980 335.870 172.740 336.040 ;
        RECT 172.990 335.870 174.160 336.040 ;
        RECT 174.400 336.010 175.220 336.040 ;
        RECT 174.400 335.870 175.510 336.010 ;
        RECT 173.390 335.770 173.740 335.870 ;
        RECT 175.050 335.840 175.510 335.870 ;
        RECT 175.960 335.840 177.150 336.010 ;
        RECT 176.000 335.820 177.150 335.840 ;
        RECT 176.980 335.780 177.150 335.820 ;
        RECT 145.730 335.590 146.050 335.620 ;
        RECT 146.830 335.590 147.150 335.620 ;
        RECT 145.720 335.480 146.050 335.590 ;
        RECT 146.820 335.480 147.150 335.590 ;
        RECT 145.720 335.400 146.110 335.480 ;
        RECT 145.730 335.360 146.110 335.400 ;
        RECT 145.940 335.100 146.110 335.360 ;
        RECT 146.490 335.100 146.660 335.480 ;
        RECT 146.820 335.400 147.210 335.480 ;
        RECT 146.830 335.360 147.210 335.400 ;
        RECT 147.040 335.100 147.210 335.360 ;
        RECT 144.080 334.860 144.400 334.890 ;
        RECT 145.180 334.860 145.500 334.890 ;
        RECT 146.270 334.860 146.590 334.890 ;
        RECT 144.070 334.790 144.400 334.860 ;
        RECT 145.170 334.790 145.500 334.860 ;
        RECT 142.640 332.390 142.810 334.790 ;
        RECT 143.190 332.390 143.360 334.790 ;
        RECT 143.740 332.390 143.910 334.790 ;
        RECT 144.070 334.670 144.460 334.790 ;
        RECT 144.080 334.630 144.460 334.670 ;
        RECT 144.290 333.550 144.460 334.630 ;
        RECT 144.070 333.520 144.460 333.550 ;
        RECT 144.060 333.330 144.460 333.520 ;
        RECT 144.070 333.290 144.460 333.330 ;
        RECT 144.290 332.390 144.460 333.290 ;
        RECT 144.840 332.850 145.010 334.790 ;
        RECT 145.170 334.670 145.560 334.790 ;
        RECT 146.260 334.670 146.590 334.860 ;
        RECT 145.180 334.630 145.560 334.670 ;
        RECT 146.270 334.630 146.590 334.670 ;
        RECT 145.390 333.540 145.560 334.630 ;
        RECT 154.080 333.580 154.840 334.000 ;
        RECT 145.180 333.510 145.560 333.540 ;
        RECT 145.170 333.320 145.560 333.510 ;
        RECT 146.270 333.490 146.590 333.520 ;
        RECT 145.180 333.280 145.560 333.320 ;
        RECT 146.260 333.300 146.590 333.490 ;
        RECT 144.630 332.820 145.010 332.850 ;
        RECT 144.620 332.630 145.010 332.820 ;
        RECT 144.630 332.590 145.010 332.630 ;
        RECT 144.840 332.390 145.010 332.590 ;
        RECT 145.390 332.390 145.560 333.280 ;
        RECT 146.270 333.260 146.590 333.300 ;
        RECT 145.730 332.810 146.050 332.840 ;
        RECT 146.820 332.810 147.140 332.840 ;
        RECT 145.720 332.620 146.050 332.810 ;
        RECT 146.810 332.620 147.140 332.810 ;
        RECT 154.100 332.790 154.840 333.580 ;
        RECT 145.730 332.580 146.050 332.620 ;
        RECT 146.820 332.580 147.140 332.620 ;
        RECT 187.150 331.720 187.320 331.750 ;
        RECT 177.340 331.690 177.510 331.720 ;
        RECT 177.340 331.650 177.660 331.690 ;
        RECT 177.340 331.460 177.670 331.650 ;
        RECT 177.340 331.430 177.660 331.460 ;
        RECT 147.490 330.540 148.000 330.720 ;
        RECT 147.430 330.510 148.000 330.540 ;
        RECT 147.420 330.320 148.000 330.510 ;
        RECT 144.260 330.100 144.430 330.320 ;
        RECT 144.120 330.070 144.440 330.100 ;
        RECT 144.110 329.880 144.440 330.070 ;
        RECT 144.120 329.840 144.440 329.880 ;
        RECT 24.080 329.330 31.610 329.840 ;
        RECT 22.380 323.310 23.840 323.350 ;
        RECT 22.380 323.140 23.850 323.310 ;
        RECT 22.380 323.100 23.840 323.140 ;
        RECT 24.080 316.720 24.590 329.330 ;
        RECT 24.950 328.540 30.930 328.770 ;
        RECT 25.040 317.480 30.690 328.540 ;
        RECT 31.100 318.970 31.610 329.330 ;
        RECT 144.260 327.920 144.430 329.840 ;
        RECT 144.810 329.430 144.980 330.320 ;
        RECT 145.360 330.110 145.530 330.320 ;
        RECT 145.220 330.080 145.540 330.110 ;
        RECT 145.210 329.890 145.540 330.080 ;
        RECT 145.220 329.850 145.540 329.890 ;
        RECT 144.670 329.400 144.990 329.430 ;
        RECT 144.660 329.210 144.990 329.400 ;
        RECT 144.670 329.170 144.990 329.210 ;
        RECT 144.810 328.060 144.980 329.170 ;
        RECT 144.670 328.030 144.990 328.060 ;
        RECT 144.660 327.920 144.990 328.030 ;
        RECT 145.360 327.920 145.530 329.850 ;
        RECT 145.910 329.430 146.080 330.320 ;
        RECT 146.460 330.110 146.630 330.320 ;
        RECT 146.310 330.080 146.630 330.110 ;
        RECT 146.300 329.890 146.630 330.080 ;
        RECT 146.310 329.850 146.630 329.890 ;
        RECT 145.770 329.400 146.090 329.430 ;
        RECT 145.760 329.210 146.090 329.400 ;
        RECT 145.770 329.170 146.090 329.210 ;
        RECT 145.910 328.060 146.080 329.170 ;
        RECT 145.770 328.030 146.090 328.060 ;
        RECT 145.760 327.920 146.090 328.030 ;
        RECT 146.460 327.920 146.630 329.850 ;
        RECT 147.010 329.430 147.180 330.310 ;
        RECT 147.430 330.280 148.000 330.320 ;
        RECT 147.490 330.070 148.000 330.280 ;
        RECT 147.440 330.040 148.000 330.070 ;
        RECT 147.430 329.850 148.010 330.040 ;
        RECT 147.440 329.810 148.010 329.850 ;
        RECT 147.490 329.790 148.010 329.810 ;
        RECT 147.500 329.710 148.010 329.790 ;
        RECT 146.870 329.400 147.190 329.430 ;
        RECT 146.860 329.210 147.190 329.400 ;
        RECT 177.340 329.230 177.510 331.430 ;
        RECT 177.890 331.010 178.060 331.720 ;
        RECT 178.440 331.690 178.610 331.720 ;
        RECT 178.430 331.650 178.750 331.690 ;
        RECT 178.430 331.460 178.760 331.650 ;
        RECT 178.430 331.430 178.750 331.460 ;
        RECT 177.890 330.970 178.210 331.010 ;
        RECT 177.890 330.780 178.220 330.970 ;
        RECT 177.890 330.750 178.210 330.780 ;
        RECT 177.890 329.640 178.060 330.750 ;
        RECT 177.890 329.600 178.210 329.640 ;
        RECT 177.890 329.410 178.220 329.600 ;
        RECT 177.890 329.380 178.210 329.410 ;
        RECT 177.890 329.220 178.060 329.380 ;
        RECT 178.440 329.220 178.610 331.430 ;
        RECT 178.990 330.990 179.160 331.720 ;
        RECT 179.540 331.680 179.710 331.720 ;
        RECT 179.530 331.640 179.850 331.680 ;
        RECT 179.530 331.450 179.860 331.640 ;
        RECT 179.530 331.420 179.850 331.450 ;
        RECT 178.980 330.950 179.300 330.990 ;
        RECT 178.980 330.760 179.310 330.950 ;
        RECT 178.980 330.730 179.300 330.760 ;
        RECT 178.990 329.640 179.160 330.730 ;
        RECT 178.980 329.600 179.300 329.640 ;
        RECT 178.980 329.410 179.310 329.600 ;
        RECT 178.980 329.380 179.300 329.410 ;
        RECT 178.990 329.220 179.160 329.380 ;
        RECT 179.540 329.220 179.710 331.420 ;
        RECT 180.090 330.980 180.260 331.720 ;
        RECT 180.090 330.940 180.410 330.980 ;
        RECT 180.090 330.750 180.420 330.940 ;
        RECT 180.570 330.900 180.740 331.660 ;
        RECT 182.460 330.900 182.630 331.660 ;
        RECT 182.940 330.980 183.110 331.720 ;
        RECT 183.490 331.680 183.660 331.720 ;
        RECT 183.350 331.640 183.670 331.680 ;
        RECT 183.340 331.450 183.670 331.640 ;
        RECT 183.350 331.420 183.670 331.450 ;
        RECT 182.790 330.940 183.110 330.980 ;
        RECT 182.780 330.750 183.110 330.940 ;
        RECT 180.090 330.720 180.410 330.750 ;
        RECT 182.790 330.720 183.110 330.750 ;
        RECT 180.090 329.640 180.260 330.720 ;
        RECT 182.940 329.640 183.110 330.720 ;
        RECT 180.080 329.600 180.400 329.640 ;
        RECT 182.800 329.600 183.120 329.640 ;
        RECT 180.080 329.410 180.410 329.600 ;
        RECT 182.790 329.410 183.120 329.600 ;
        RECT 180.080 329.380 180.400 329.410 ;
        RECT 182.800 329.380 183.120 329.410 ;
        RECT 180.090 329.220 180.260 329.380 ;
        RECT 182.940 329.220 183.110 329.380 ;
        RECT 183.490 329.220 183.660 331.420 ;
        RECT 184.040 330.990 184.210 331.720 ;
        RECT 184.590 331.690 184.760 331.720 ;
        RECT 184.450 331.650 184.770 331.690 ;
        RECT 184.440 331.460 184.770 331.650 ;
        RECT 184.450 331.430 184.770 331.460 ;
        RECT 183.900 330.950 184.220 330.990 ;
        RECT 183.890 330.760 184.220 330.950 ;
        RECT 183.900 330.730 184.220 330.760 ;
        RECT 184.040 329.640 184.210 330.730 ;
        RECT 183.900 329.600 184.220 329.640 ;
        RECT 183.890 329.410 184.220 329.600 ;
        RECT 183.900 329.380 184.220 329.410 ;
        RECT 184.040 329.220 184.210 329.380 ;
        RECT 184.590 329.220 184.760 331.430 ;
        RECT 185.140 331.010 185.310 331.720 ;
        RECT 185.690 331.690 185.860 331.720 ;
        RECT 185.540 331.650 185.860 331.690 ;
        RECT 185.530 331.460 185.860 331.650 ;
        RECT 185.540 331.430 185.860 331.460 ;
        RECT 184.990 330.970 185.310 331.010 ;
        RECT 184.980 330.780 185.310 330.970 ;
        RECT 184.990 330.750 185.310 330.780 ;
        RECT 185.140 329.640 185.310 330.750 ;
        RECT 184.990 329.600 185.310 329.640 ;
        RECT 184.980 329.410 185.310 329.600 ;
        RECT 184.990 329.380 185.310 329.410 ;
        RECT 185.140 329.220 185.310 329.380 ;
        RECT 185.690 329.230 185.860 331.430 ;
        RECT 187.150 331.680 187.470 331.720 ;
        RECT 187.150 331.490 187.480 331.680 ;
        RECT 187.150 331.460 187.470 331.490 ;
        RECT 187.150 329.260 187.320 331.460 ;
        RECT 187.700 331.040 187.870 331.750 ;
        RECT 188.250 331.720 188.420 331.750 ;
        RECT 188.240 331.680 188.560 331.720 ;
        RECT 188.240 331.490 188.570 331.680 ;
        RECT 188.240 331.460 188.560 331.490 ;
        RECT 187.700 331.000 188.020 331.040 ;
        RECT 187.700 330.810 188.030 331.000 ;
        RECT 187.700 330.780 188.020 330.810 ;
        RECT 187.700 329.670 187.870 330.780 ;
        RECT 187.700 329.630 188.020 329.670 ;
        RECT 187.700 329.440 188.030 329.630 ;
        RECT 187.700 329.410 188.020 329.440 ;
        RECT 187.700 329.250 187.870 329.410 ;
        RECT 188.250 329.250 188.420 331.460 ;
        RECT 188.800 331.020 188.970 331.750 ;
        RECT 189.350 331.710 189.520 331.750 ;
        RECT 189.340 331.670 189.660 331.710 ;
        RECT 189.340 331.480 189.670 331.670 ;
        RECT 189.340 331.450 189.660 331.480 ;
        RECT 188.790 330.980 189.110 331.020 ;
        RECT 188.790 330.790 189.120 330.980 ;
        RECT 188.790 330.760 189.110 330.790 ;
        RECT 188.800 329.670 188.970 330.760 ;
        RECT 188.790 329.630 189.110 329.670 ;
        RECT 188.790 329.440 189.120 329.630 ;
        RECT 188.790 329.410 189.110 329.440 ;
        RECT 188.800 329.250 188.970 329.410 ;
        RECT 189.350 329.250 189.520 331.450 ;
        RECT 189.900 331.010 190.070 331.750 ;
        RECT 189.900 330.970 190.220 331.010 ;
        RECT 189.900 330.780 190.230 330.970 ;
        RECT 190.380 330.930 190.550 331.690 ;
        RECT 192.270 330.930 192.440 331.690 ;
        RECT 192.750 331.010 192.920 331.750 ;
        RECT 193.300 331.710 193.470 331.750 ;
        RECT 193.160 331.670 193.480 331.710 ;
        RECT 193.150 331.480 193.480 331.670 ;
        RECT 193.160 331.450 193.480 331.480 ;
        RECT 192.600 330.970 192.920 331.010 ;
        RECT 192.590 330.780 192.920 330.970 ;
        RECT 189.900 330.750 190.220 330.780 ;
        RECT 192.600 330.750 192.920 330.780 ;
        RECT 189.900 329.670 190.070 330.750 ;
        RECT 192.750 329.670 192.920 330.750 ;
        RECT 189.890 329.630 190.210 329.670 ;
        RECT 192.610 329.630 192.930 329.670 ;
        RECT 189.890 329.440 190.220 329.630 ;
        RECT 192.600 329.440 192.930 329.630 ;
        RECT 189.890 329.410 190.210 329.440 ;
        RECT 192.610 329.410 192.930 329.440 ;
        RECT 189.900 329.250 190.070 329.410 ;
        RECT 192.750 329.250 192.920 329.410 ;
        RECT 193.300 329.250 193.470 331.450 ;
        RECT 193.850 331.020 194.020 331.750 ;
        RECT 194.400 331.720 194.570 331.750 ;
        RECT 194.260 331.680 194.580 331.720 ;
        RECT 194.250 331.490 194.580 331.680 ;
        RECT 194.260 331.460 194.580 331.490 ;
        RECT 193.710 330.980 194.030 331.020 ;
        RECT 193.700 330.790 194.030 330.980 ;
        RECT 193.710 330.760 194.030 330.790 ;
        RECT 193.850 329.670 194.020 330.760 ;
        RECT 193.710 329.630 194.030 329.670 ;
        RECT 193.700 329.440 194.030 329.630 ;
        RECT 193.710 329.410 194.030 329.440 ;
        RECT 193.850 329.250 194.020 329.410 ;
        RECT 194.400 329.250 194.570 331.460 ;
        RECT 194.950 331.040 195.120 331.750 ;
        RECT 195.500 331.720 195.670 331.750 ;
        RECT 195.350 331.680 195.670 331.720 ;
        RECT 195.340 331.490 195.670 331.680 ;
        RECT 195.350 331.460 195.670 331.490 ;
        RECT 194.800 331.000 195.120 331.040 ;
        RECT 194.790 330.810 195.120 331.000 ;
        RECT 194.800 330.780 195.120 330.810 ;
        RECT 194.950 329.670 195.120 330.780 ;
        RECT 194.800 329.630 195.120 329.670 ;
        RECT 194.790 329.440 195.120 329.630 ;
        RECT 194.800 329.410 195.120 329.440 ;
        RECT 194.950 329.250 195.120 329.410 ;
        RECT 195.500 329.260 195.670 331.460 ;
        RECT 196.910 329.490 197.080 331.890 ;
        RECT 197.460 329.490 197.630 331.890 ;
        RECT 198.010 329.490 198.180 331.890 ;
        RECT 198.560 330.990 198.730 331.890 ;
        RECT 199.110 331.690 199.280 331.890 ;
        RECT 198.900 331.650 199.280 331.690 ;
        RECT 198.890 331.460 199.280 331.650 ;
        RECT 198.900 331.430 199.280 331.460 ;
        RECT 198.340 330.950 198.730 330.990 ;
        RECT 198.330 330.760 198.730 330.950 ;
        RECT 198.340 330.730 198.730 330.760 ;
        RECT 198.560 329.650 198.730 330.730 ;
        RECT 198.350 329.610 198.730 329.650 ;
        RECT 198.340 329.490 198.730 329.610 ;
        RECT 199.110 329.490 199.280 331.430 ;
        RECT 199.660 331.000 199.830 331.890 ;
        RECT 200.000 331.660 200.320 331.700 ;
        RECT 201.090 331.660 201.410 331.700 ;
        RECT 199.990 331.470 200.320 331.660 ;
        RECT 201.080 331.470 201.410 331.660 ;
        RECT 200.000 331.440 200.320 331.470 ;
        RECT 201.090 331.440 201.410 331.470 ;
        RECT 199.450 330.960 199.830 331.000 ;
        RECT 200.540 330.980 200.860 331.020 ;
        RECT 199.440 330.770 199.830 330.960 ;
        RECT 200.530 330.790 200.860 330.980 ;
        RECT 199.450 330.740 199.830 330.770 ;
        RECT 200.540 330.760 200.860 330.790 ;
        RECT 199.660 329.650 199.830 330.740 ;
        RECT 199.450 329.610 199.830 329.650 ;
        RECT 200.540 329.610 200.860 329.650 ;
        RECT 199.440 329.490 199.830 329.610 ;
        RECT 198.340 329.420 198.670 329.490 ;
        RECT 199.440 329.420 199.770 329.490 ;
        RECT 200.530 329.420 200.860 329.610 ;
        RECT 198.350 329.390 198.670 329.420 ;
        RECT 199.450 329.390 199.770 329.420 ;
        RECT 200.540 329.390 200.860 329.420 ;
        RECT 146.870 329.170 147.190 329.210 ;
        RECT 147.010 328.060 147.180 329.170 ;
        RECT 177.280 329.140 177.440 329.170 ;
        RECT 177.280 328.910 177.450 329.140 ;
        RECT 177.830 329.130 177.990 329.170 ;
        RECT 177.280 328.870 177.650 328.910 ;
        RECT 177.830 328.890 178.000 329.130 ;
        RECT 178.380 328.910 178.550 329.200 ;
        RECT 178.930 329.130 179.090 329.170 ;
        RECT 179.480 329.130 179.640 329.170 ;
        RECT 180.030 329.150 180.190 329.170 ;
        RECT 183.010 329.150 183.170 329.170 ;
        RECT 177.280 328.790 177.660 328.870 ;
        RECT 177.830 328.790 178.060 328.890 ;
        RECT 178.380 328.870 178.750 328.910 ;
        RECT 178.930 328.890 179.100 329.130 ;
        RECT 179.480 328.910 179.650 329.130 ;
        RECT 178.380 328.790 178.760 328.870 ;
        RECT 178.930 328.790 179.160 328.890 ;
        RECT 179.480 328.870 179.850 328.910 ;
        RECT 180.030 328.890 180.200 329.150 ;
        RECT 183.000 328.890 183.170 329.150 ;
        RECT 183.560 329.130 183.720 329.170 ;
        RECT 184.110 329.130 184.270 329.170 ;
        RECT 183.550 328.910 183.720 329.130 ;
        RECT 179.480 328.790 179.860 328.870 ;
        RECT 180.030 328.790 180.260 328.890 ;
        RECT 177.330 328.680 177.660 328.790 ;
        RECT 177.330 328.650 177.650 328.680 ;
        RECT 146.870 328.030 147.190 328.060 ;
        RECT 146.860 327.920 147.190 328.030 ;
        RECT 144.260 327.820 144.490 327.920 ;
        RECT 144.660 327.840 145.040 327.920 ;
        RECT 144.320 327.560 144.490 327.820 ;
        RECT 144.670 327.800 145.040 327.840 ;
        RECT 145.360 327.820 145.590 327.920 ;
        RECT 145.760 327.840 146.140 327.920 ;
        RECT 144.870 327.580 145.040 327.800 ;
        RECT 145.420 327.580 145.590 327.820 ;
        RECT 145.770 327.800 146.140 327.840 ;
        RECT 146.460 327.820 146.690 327.920 ;
        RECT 146.860 327.840 147.240 327.920 ;
        RECT 144.330 327.540 144.490 327.560 ;
        RECT 144.880 327.540 145.040 327.580 ;
        RECT 145.430 327.540 145.590 327.580 ;
        RECT 145.970 327.510 146.140 327.800 ;
        RECT 146.520 327.580 146.690 327.820 ;
        RECT 146.870 327.800 147.240 327.840 ;
        RECT 146.530 327.540 146.690 327.580 ;
        RECT 147.070 327.570 147.240 327.800 ;
        RECT 147.080 327.540 147.240 327.570 ;
        RECT 177.340 327.540 177.510 328.650 ;
        RECT 177.330 327.500 177.650 327.540 ;
        RECT 144.260 327.330 144.430 327.490 ;
        RECT 144.120 327.300 144.440 327.330 ;
        RECT 144.110 327.110 144.440 327.300 ;
        RECT 144.120 327.070 144.440 327.110 ;
        RECT 144.260 325.990 144.430 327.070 ;
        RECT 144.110 325.960 144.430 325.990 ;
        RECT 143.780 325.050 143.950 325.810 ;
        RECT 144.100 325.770 144.430 325.960 ;
        RECT 144.110 325.730 144.430 325.770 ;
        RECT 144.260 324.990 144.430 325.730 ;
        RECT 144.810 325.290 144.980 327.490 ;
        RECT 145.360 327.330 145.530 327.490 ;
        RECT 145.220 327.300 145.540 327.330 ;
        RECT 145.210 327.110 145.540 327.300 ;
        RECT 145.220 327.070 145.540 327.110 ;
        RECT 145.360 325.980 145.530 327.070 ;
        RECT 145.220 325.950 145.540 325.980 ;
        RECT 145.210 325.760 145.540 325.950 ;
        RECT 145.220 325.720 145.540 325.760 ;
        RECT 144.670 325.260 144.990 325.290 ;
        RECT 144.660 325.070 144.990 325.260 ;
        RECT 144.670 325.030 144.990 325.070 ;
        RECT 144.810 324.990 144.980 325.030 ;
        RECT 145.360 324.990 145.530 325.720 ;
        RECT 145.910 325.280 146.080 327.490 ;
        RECT 146.460 327.330 146.630 327.490 ;
        RECT 146.310 327.300 146.630 327.330 ;
        RECT 146.300 327.110 146.630 327.300 ;
        RECT 146.310 327.070 146.630 327.110 ;
        RECT 146.460 325.960 146.630 327.070 ;
        RECT 146.310 325.930 146.630 325.960 ;
        RECT 146.300 325.740 146.630 325.930 ;
        RECT 146.310 325.700 146.630 325.740 ;
        RECT 145.770 325.250 146.090 325.280 ;
        RECT 145.760 325.060 146.090 325.250 ;
        RECT 145.770 325.020 146.090 325.060 ;
        RECT 145.910 324.990 146.080 325.020 ;
        RECT 146.460 324.990 146.630 325.700 ;
        RECT 147.010 325.280 147.180 327.480 ;
        RECT 177.330 327.310 177.660 327.500 ;
        RECT 177.330 327.280 177.650 327.310 ;
        RECT 176.510 326.920 177.020 327.000 ;
        RECT 176.510 326.900 177.030 326.920 ;
        RECT 176.510 326.860 177.080 326.900 ;
        RECT 176.510 326.670 177.090 326.860 ;
        RECT 176.520 326.640 177.080 326.670 ;
        RECT 176.520 326.430 177.030 326.640 ;
        RECT 176.520 326.390 177.090 326.430 ;
        RECT 177.340 326.400 177.510 327.280 ;
        RECT 177.890 326.860 178.060 328.790 ;
        RECT 178.430 328.680 178.760 328.790 ;
        RECT 178.430 328.650 178.750 328.680 ;
        RECT 178.440 327.540 178.610 328.650 ;
        RECT 178.430 327.500 178.750 327.540 ;
        RECT 178.430 327.310 178.760 327.500 ;
        RECT 178.430 327.280 178.750 327.310 ;
        RECT 177.890 326.820 178.210 326.860 ;
        RECT 177.890 326.630 178.220 326.820 ;
        RECT 177.890 326.600 178.210 326.630 ;
        RECT 177.890 326.390 178.060 326.600 ;
        RECT 178.440 326.390 178.610 327.280 ;
        RECT 178.990 326.860 179.160 328.790 ;
        RECT 179.530 328.680 179.860 328.790 ;
        RECT 179.530 328.650 179.850 328.680 ;
        RECT 179.540 327.540 179.710 328.650 ;
        RECT 179.530 327.500 179.850 327.540 ;
        RECT 179.530 327.310 179.860 327.500 ;
        RECT 179.530 327.280 179.850 327.310 ;
        RECT 178.980 326.820 179.300 326.860 ;
        RECT 178.980 326.630 179.310 326.820 ;
        RECT 178.980 326.600 179.300 326.630 ;
        RECT 178.990 326.390 179.160 326.600 ;
        RECT 179.540 326.390 179.710 327.280 ;
        RECT 180.090 326.870 180.260 328.790 ;
        RECT 182.940 328.790 183.170 328.890 ;
        RECT 183.350 328.870 183.720 328.910 ;
        RECT 184.100 328.890 184.270 329.130 ;
        RECT 184.650 328.910 184.820 329.200 ;
        RECT 187.090 329.170 187.250 329.200 ;
        RECT 185.210 329.130 185.370 329.170 ;
        RECT 185.760 329.140 185.920 329.170 ;
        RECT 183.340 328.790 183.720 328.870 ;
        RECT 184.040 328.790 184.270 328.890 ;
        RECT 184.450 328.870 184.820 328.910 ;
        RECT 185.200 328.890 185.370 329.130 ;
        RECT 185.750 328.910 185.920 329.140 ;
        RECT 184.440 328.790 184.820 328.870 ;
        RECT 185.140 328.790 185.370 328.890 ;
        RECT 185.550 328.870 185.920 328.910 ;
        RECT 185.540 328.790 185.920 328.870 ;
        RECT 187.090 328.940 187.260 329.170 ;
        RECT 187.640 329.160 187.800 329.200 ;
        RECT 187.090 328.900 187.460 328.940 ;
        RECT 187.640 328.920 187.810 329.160 ;
        RECT 188.190 328.940 188.360 329.230 ;
        RECT 188.740 329.160 188.900 329.200 ;
        RECT 189.290 329.160 189.450 329.200 ;
        RECT 189.840 329.180 190.000 329.200 ;
        RECT 192.820 329.180 192.980 329.200 ;
        RECT 187.090 328.820 187.470 328.900 ;
        RECT 187.640 328.820 187.870 328.920 ;
        RECT 188.190 328.900 188.560 328.940 ;
        RECT 188.740 328.920 188.910 329.160 ;
        RECT 189.290 328.940 189.460 329.160 ;
        RECT 188.190 328.820 188.570 328.900 ;
        RECT 188.740 328.820 188.970 328.920 ;
        RECT 189.290 328.900 189.660 328.940 ;
        RECT 189.840 328.920 190.010 329.180 ;
        RECT 192.810 328.920 192.980 329.180 ;
        RECT 193.370 329.160 193.530 329.200 ;
        RECT 193.920 329.160 194.080 329.200 ;
        RECT 193.360 328.940 193.530 329.160 ;
        RECT 189.290 328.820 189.670 328.900 ;
        RECT 189.840 328.820 190.070 328.920 ;
        RECT 182.940 326.870 183.110 328.790 ;
        RECT 183.340 328.680 183.670 328.790 ;
        RECT 183.350 328.650 183.670 328.680 ;
        RECT 183.490 327.540 183.660 328.650 ;
        RECT 183.350 327.500 183.670 327.540 ;
        RECT 183.340 327.310 183.670 327.500 ;
        RECT 183.350 327.280 183.670 327.310 ;
        RECT 180.080 326.830 180.400 326.870 ;
        RECT 182.800 326.830 183.120 326.870 ;
        RECT 180.080 326.640 180.410 326.830 ;
        RECT 182.790 326.640 183.120 326.830 ;
        RECT 180.080 326.610 180.400 326.640 ;
        RECT 182.800 326.610 183.120 326.640 ;
        RECT 180.090 326.390 180.260 326.610 ;
        RECT 182.940 326.390 183.110 326.610 ;
        RECT 183.490 326.390 183.660 327.280 ;
        RECT 184.040 326.860 184.210 328.790 ;
        RECT 184.440 328.680 184.770 328.790 ;
        RECT 184.450 328.650 184.770 328.680 ;
        RECT 184.590 327.540 184.760 328.650 ;
        RECT 184.450 327.500 184.770 327.540 ;
        RECT 184.440 327.310 184.770 327.500 ;
        RECT 184.450 327.280 184.770 327.310 ;
        RECT 183.900 326.820 184.220 326.860 ;
        RECT 183.890 326.630 184.220 326.820 ;
        RECT 183.900 326.600 184.220 326.630 ;
        RECT 184.040 326.390 184.210 326.600 ;
        RECT 184.590 326.390 184.760 327.280 ;
        RECT 185.140 326.860 185.310 328.790 ;
        RECT 185.540 328.680 185.870 328.790 ;
        RECT 187.140 328.710 187.470 328.820 ;
        RECT 187.140 328.680 187.460 328.710 ;
        RECT 185.550 328.650 185.870 328.680 ;
        RECT 185.690 327.540 185.860 328.650 ;
        RECT 187.150 327.570 187.320 328.680 ;
        RECT 185.550 327.500 185.870 327.540 ;
        RECT 185.540 327.310 185.870 327.500 ;
        RECT 187.140 327.530 187.460 327.570 ;
        RECT 187.140 327.340 187.470 327.530 ;
        RECT 187.140 327.310 187.460 327.340 ;
        RECT 185.550 327.280 185.870 327.310 ;
        RECT 184.990 326.820 185.310 326.860 ;
        RECT 184.980 326.630 185.310 326.820 ;
        RECT 184.990 326.600 185.310 326.630 ;
        RECT 185.140 326.390 185.310 326.600 ;
        RECT 185.690 326.400 185.860 327.280 ;
        RECT 186.320 327.000 186.830 327.030 ;
        RECT 186.180 326.950 186.830 327.000 ;
        RECT 186.180 326.930 186.840 326.950 ;
        RECT 186.180 326.920 186.890 326.930 ;
        RECT 186.170 326.900 186.890 326.920 ;
        RECT 186.120 326.890 186.890 326.900 ;
        RECT 186.120 326.860 186.900 326.890 ;
        RECT 186.110 326.700 186.900 326.860 ;
        RECT 186.110 326.670 186.890 326.700 ;
        RECT 186.120 326.640 186.840 326.670 ;
        RECT 186.170 326.460 186.840 326.640 ;
        RECT 186.170 326.430 186.900 326.460 ;
        RECT 187.150 326.430 187.320 327.310 ;
        RECT 187.700 326.890 187.870 328.820 ;
        RECT 188.240 328.710 188.570 328.820 ;
        RECT 188.240 328.680 188.560 328.710 ;
        RECT 188.250 327.570 188.420 328.680 ;
        RECT 188.240 327.530 188.560 327.570 ;
        RECT 188.240 327.340 188.570 327.530 ;
        RECT 188.240 327.310 188.560 327.340 ;
        RECT 187.700 326.850 188.020 326.890 ;
        RECT 187.700 326.660 188.030 326.850 ;
        RECT 187.700 326.630 188.020 326.660 ;
        RECT 186.110 326.420 186.900 326.430 ;
        RECT 187.700 326.420 187.870 326.630 ;
        RECT 188.250 326.420 188.420 327.310 ;
        RECT 188.800 326.890 188.970 328.820 ;
        RECT 189.340 328.710 189.670 328.820 ;
        RECT 189.340 328.680 189.660 328.710 ;
        RECT 189.350 327.570 189.520 328.680 ;
        RECT 189.340 327.530 189.660 327.570 ;
        RECT 189.340 327.340 189.670 327.530 ;
        RECT 189.340 327.310 189.660 327.340 ;
        RECT 188.790 326.850 189.110 326.890 ;
        RECT 188.790 326.660 189.120 326.850 ;
        RECT 188.790 326.630 189.110 326.660 ;
        RECT 188.800 326.420 188.970 326.630 ;
        RECT 189.350 326.420 189.520 327.310 ;
        RECT 189.900 326.900 190.070 328.820 ;
        RECT 192.750 328.820 192.980 328.920 ;
        RECT 193.160 328.900 193.530 328.940 ;
        RECT 193.910 328.920 194.080 329.160 ;
        RECT 194.460 328.940 194.630 329.230 ;
        RECT 195.020 329.160 195.180 329.200 ;
        RECT 195.570 329.170 195.730 329.200 ;
        RECT 193.150 328.820 193.530 328.900 ;
        RECT 193.850 328.820 194.080 328.920 ;
        RECT 194.260 328.900 194.630 328.940 ;
        RECT 195.010 328.920 195.180 329.160 ;
        RECT 195.560 328.940 195.730 329.170 ;
        RECT 194.250 328.820 194.630 328.900 ;
        RECT 194.950 328.820 195.180 328.920 ;
        RECT 195.360 328.900 195.730 328.940 ;
        RECT 195.350 328.820 195.730 328.900 ;
        RECT 192.750 326.900 192.920 328.820 ;
        RECT 193.150 328.710 193.480 328.820 ;
        RECT 193.160 328.680 193.480 328.710 ;
        RECT 193.300 327.570 193.470 328.680 ;
        RECT 193.160 327.530 193.480 327.570 ;
        RECT 193.150 327.340 193.480 327.530 ;
        RECT 193.160 327.310 193.480 327.340 ;
        RECT 189.890 326.860 190.210 326.900 ;
        RECT 192.610 326.860 192.930 326.900 ;
        RECT 189.890 326.670 190.220 326.860 ;
        RECT 192.600 326.670 192.930 326.860 ;
        RECT 189.890 326.640 190.210 326.670 ;
        RECT 192.610 326.640 192.930 326.670 ;
        RECT 189.900 326.420 190.070 326.640 ;
        RECT 192.750 326.420 192.920 326.640 ;
        RECT 193.300 326.420 193.470 327.310 ;
        RECT 193.850 326.890 194.020 328.820 ;
        RECT 194.250 328.710 194.580 328.820 ;
        RECT 194.260 328.680 194.580 328.710 ;
        RECT 194.400 327.570 194.570 328.680 ;
        RECT 194.260 327.530 194.580 327.570 ;
        RECT 194.250 327.340 194.580 327.530 ;
        RECT 194.260 327.310 194.580 327.340 ;
        RECT 193.710 326.850 194.030 326.890 ;
        RECT 193.700 326.660 194.030 326.850 ;
        RECT 193.710 326.630 194.030 326.660 ;
        RECT 193.850 326.420 194.020 326.630 ;
        RECT 194.400 326.420 194.570 327.310 ;
        RECT 194.950 326.890 195.120 328.820 ;
        RECT 195.350 328.710 195.680 328.820 ;
        RECT 195.360 328.680 195.680 328.710 ;
        RECT 195.500 327.570 195.670 328.680 ;
        RECT 195.360 327.530 195.680 327.570 ;
        RECT 195.350 327.340 195.680 327.530 ;
        RECT 195.360 327.310 195.680 327.340 ;
        RECT 194.800 326.850 195.120 326.890 ;
        RECT 194.790 326.660 195.120 326.850 ;
        RECT 194.800 326.630 195.120 326.660 ;
        RECT 194.950 326.420 195.120 326.630 ;
        RECT 195.500 326.430 195.670 327.310 ;
        RECT 195.990 326.950 196.500 327.030 ;
        RECT 195.980 326.930 196.500 326.950 ;
        RECT 195.930 326.890 196.500 326.930 ;
        RECT 195.920 326.700 196.500 326.890 ;
        RECT 196.910 326.710 197.080 329.110 ;
        RECT 197.460 326.710 197.630 329.110 ;
        RECT 198.010 326.710 198.180 329.110 ;
        RECT 198.560 326.880 198.730 329.180 ;
        RECT 199.110 328.920 199.280 329.180 ;
        RECT 198.900 328.880 199.280 328.920 ;
        RECT 198.890 328.690 199.280 328.880 ;
        RECT 198.900 328.660 199.280 328.690 ;
        RECT 199.110 327.550 199.280 328.660 ;
        RECT 198.900 327.510 199.280 327.550 ;
        RECT 198.890 327.320 199.280 327.510 ;
        RECT 198.900 327.290 199.280 327.320 ;
        RECT 198.350 326.840 198.730 326.880 ;
        RECT 198.340 326.710 198.730 326.840 ;
        RECT 199.110 326.710 199.280 327.290 ;
        RECT 199.660 326.870 199.830 329.180 ;
        RECT 200.210 328.920 200.380 329.180 ;
        RECT 200.000 328.880 200.380 328.920 ;
        RECT 199.990 328.800 200.380 328.880 ;
        RECT 200.760 328.800 200.930 329.180 ;
        RECT 201.310 328.920 201.480 329.180 ;
        RECT 201.100 328.880 201.480 328.920 ;
        RECT 201.090 328.800 201.480 328.880 ;
        RECT 199.990 328.690 200.320 328.800 ;
        RECT 201.090 328.690 201.420 328.800 ;
        RECT 200.000 328.660 200.320 328.690 ;
        RECT 201.100 328.660 201.420 328.690 ;
        RECT 200.000 327.510 200.320 327.550 ;
        RECT 201.100 327.510 201.420 327.550 ;
        RECT 199.990 327.320 200.320 327.510 ;
        RECT 201.090 327.320 201.420 327.510 ;
        RECT 200.000 327.290 200.320 327.320 ;
        RECT 201.100 327.290 201.420 327.320 ;
        RECT 202.020 327.200 202.190 328.420 ;
        RECT 201.730 326.910 202.240 327.010 ;
        RECT 201.670 326.870 202.240 326.910 ;
        RECT 199.450 326.830 199.830 326.870 ;
        RECT 200.540 326.830 200.860 326.870 ;
        RECT 199.440 326.710 199.830 326.830 ;
        RECT 195.930 326.670 196.490 326.700 ;
        RECT 195.980 326.460 196.490 326.670 ;
        RECT 198.340 326.650 198.670 326.710 ;
        RECT 198.350 326.620 198.670 326.650 ;
        RECT 199.440 326.640 199.770 326.710 ;
        RECT 200.530 326.640 200.860 326.830 ;
        RECT 201.660 326.680 202.240 326.870 ;
        RECT 201.670 326.650 202.230 326.680 ;
        RECT 199.450 326.610 199.770 326.640 ;
        RECT 200.540 326.610 200.860 326.640 ;
        RECT 195.920 326.420 196.490 326.460 ;
        RECT 201.720 326.440 202.230 326.650 ;
        RECT 186.110 326.390 186.910 326.420 ;
        RECT 176.520 326.200 177.100 326.390 ;
        RECT 186.100 326.230 186.910 326.390 ;
        RECT 195.910 326.230 196.490 326.420 ;
        RECT 201.660 326.400 202.230 326.440 ;
        RECT 186.100 326.200 186.900 326.230 ;
        RECT 195.920 326.200 196.490 326.230 ;
        RECT 201.650 326.210 202.230 326.400 ;
        RECT 176.520 326.170 177.090 326.200 ;
        RECT 186.110 326.170 186.840 326.200 ;
        RECT 176.520 325.990 177.030 326.170 ;
        RECT 186.170 326.020 186.840 326.170 ;
        RECT 195.980 326.020 196.490 326.200 ;
        RECT 201.660 326.180 202.230 326.210 ;
        RECT 186.170 325.990 186.680 326.020 ;
        RECT 201.720 326.000 202.230 326.180 ;
        RECT 146.860 325.250 147.180 325.280 ;
        RECT 146.850 325.060 147.180 325.250 ;
        RECT 146.860 325.020 147.180 325.060 ;
        RECT 147.010 324.990 147.180 325.020 ;
        RECT 148.430 324.890 150.820 325.260 ;
        RECT 148.480 321.630 150.820 324.890 ;
        RECT 227.300 324.090 227.530 324.200 ;
        RECT 227.200 323.990 231.860 324.090 ;
        RECT 227.200 323.920 232.050 323.990 ;
        RECT 230.760 323.820 231.090 323.920 ;
        RECT 231.720 323.820 232.050 323.920 ;
        RECT 232.680 323.820 233.010 323.990 ;
        RECT 233.640 323.820 233.970 323.990 ;
        RECT 232.910 323.580 233.100 323.590 ;
        RECT 228.420 323.400 232.220 323.410 ;
        RECT 232.880 323.400 233.140 323.580 ;
        RECT 228.420 323.260 233.140 323.400 ;
        RECT 228.420 323.240 233.010 323.260 ;
        RECT 230.760 323.140 231.090 323.240 ;
        RECT 231.720 323.230 233.010 323.240 ;
        RECT 231.720 323.140 232.220 323.230 ;
        RECT 232.680 323.140 233.010 323.230 ;
        RECT 233.640 323.140 233.970 323.310 ;
        RECT 231.990 322.770 232.220 323.140 ;
        RECT 232.910 322.910 233.100 322.920 ;
        RECT 232.880 322.770 233.140 322.910 ;
        RECT 231.990 322.590 233.140 322.770 ;
        RECT 227.300 322.480 227.530 322.590 ;
        RECT 231.990 322.560 233.000 322.590 ;
        RECT 227.200 322.310 231.680 322.480 ;
        RECT 231.990 322.380 232.220 322.560 ;
        RECT 230.760 322.210 231.090 322.310 ;
        RECT 231.720 322.210 232.220 322.380 ;
        RECT 232.680 322.210 233.010 322.380 ;
        RECT 233.640 322.210 233.970 322.380 ;
        RECT 231.990 321.800 232.220 322.210 ;
        RECT 228.450 321.630 232.220 321.800 ;
        RECT 148.480 321.620 150.810 321.630 ;
        RECT 230.760 321.530 231.090 321.630 ;
        RECT 231.720 321.530 232.220 321.630 ;
        RECT 232.680 321.550 233.010 321.700 ;
        RECT 232.680 321.530 233.400 321.550 ;
        RECT 233.640 321.530 233.970 321.700 ;
        RECT 227.300 320.880 227.530 320.990 ;
        RECT 227.200 320.710 231.700 320.880 ;
        RECT 231.990 320.770 232.220 321.530 ;
        RECT 232.950 321.360 233.400 321.530 ;
        RECT 232.970 321.340 233.400 321.360 ;
        RECT 230.760 320.600 231.090 320.710 ;
        RECT 231.720 320.600 232.220 320.770 ;
        RECT 232.680 320.600 233.010 320.770 ;
        RECT 233.640 320.600 233.970 320.770 ;
        RECT 231.990 320.190 232.220 320.600 ;
        RECT 228.460 320.020 232.220 320.190 ;
        RECT 230.760 319.920 231.090 320.020 ;
        RECT 231.720 319.920 232.220 320.020 ;
        RECT 232.680 319.940 233.010 320.090 ;
        RECT 232.680 319.920 233.400 319.940 ;
        RECT 233.640 319.920 233.970 320.090 ;
        RECT 231.200 319.730 231.630 319.750 ;
        RECT 231.180 319.560 231.630 319.730 ;
        RECT 231.200 319.540 231.630 319.560 ;
        RECT 227.300 319.260 227.530 319.370 ;
        RECT 227.200 319.090 231.700 319.260 ;
        RECT 230.760 318.990 231.090 319.090 ;
        RECT 31.090 318.950 31.610 318.970 ;
        RECT 25.040 317.470 30.750 317.480 ;
        RECT 24.960 317.300 30.750 317.470 ;
        RECT 25.050 317.290 30.750 317.300 ;
        RECT 30.520 317.220 30.690 317.290 ;
        RECT 31.090 317.170 31.620 318.950 ;
        RECT 231.990 318.590 232.220 319.920 ;
        RECT 232.950 319.750 233.400 319.920 ;
        RECT 232.970 319.730 233.400 319.750 ;
        RECT 232.680 318.990 233.010 319.160 ;
        RECT 233.640 318.990 233.970 319.160 ;
        RECT 228.450 318.420 232.220 318.590 ;
        RECT 230.760 318.310 231.090 318.420 ;
        RECT 231.990 318.170 232.220 318.420 ;
        RECT 232.680 318.330 233.010 318.480 ;
        RECT 232.680 318.310 233.390 318.330 ;
        RECT 233.640 318.310 233.970 318.480 ;
        RECT 231.990 318.150 232.490 318.170 ;
        RECT 231.990 317.980 232.510 318.150 ;
        RECT 232.940 318.140 233.390 318.310 ;
        RECT 232.960 318.120 233.390 318.140 ;
        RECT 231.990 317.960 232.490 317.980 ;
        RECT 227.300 317.660 227.530 317.770 ;
        RECT 227.200 317.490 231.650 317.660 ;
        RECT 231.990 317.550 232.220 317.960 ;
        RECT 230.760 317.380 231.090 317.490 ;
        RECT 231.720 317.380 232.220 317.550 ;
        RECT 233.180 317.440 233.510 317.610 ;
        RECT 233.640 317.380 233.970 317.550 ;
        RECT 31.100 317.150 31.620 317.170 ;
        RECT 24.080 316.430 26.520 316.720 ;
        RECT 31.100 316.640 31.610 317.150 ;
        RECT 231.990 316.970 232.220 317.380 ;
        RECT 228.430 316.800 232.220 316.970 ;
        RECT 230.760 316.700 231.090 316.800 ;
        RECT 231.720 316.700 232.220 316.800 ;
        RECT 233.180 316.760 233.510 316.930 ;
        RECT 31.100 316.430 31.630 316.640 ;
        RECT 24.080 315.950 31.630 316.430 ;
        RECT 227.300 316.040 227.530 316.150 ;
        RECT 24.080 315.920 31.440 315.950 ;
        RECT 227.200 315.870 231.700 316.040 ;
        RECT 231.990 315.940 232.220 316.700 ;
        RECT 232.970 316.690 233.400 316.710 ;
        RECT 233.640 316.700 233.970 316.870 ;
        RECT 232.950 316.520 233.400 316.690 ;
        RECT 233.490 316.570 233.920 316.590 ;
        RECT 232.970 316.500 233.400 316.520 ;
        RECT 233.470 316.400 233.920 316.570 ;
        RECT 233.490 316.380 233.920 316.400 ;
        RECT 230.760 315.770 231.090 315.870 ;
        RECT 231.720 315.770 232.220 315.940 ;
        RECT 232.680 315.770 233.010 315.940 ;
        RECT 233.640 315.770 233.970 315.940 ;
        RECT 231.990 315.350 232.220 315.770 ;
        RECT 228.430 315.180 232.220 315.350 ;
        RECT 230.760 315.090 231.090 315.180 ;
        RECT 231.720 315.090 232.220 315.180 ;
        RECT 232.680 315.100 233.010 315.260 ;
        RECT 232.680 315.090 233.390 315.100 ;
        RECT 233.640 315.090 233.970 315.260 ;
        RECT 24.080 314.160 31.610 314.710 ;
        RECT 227.300 314.440 227.530 314.550 ;
        RECT 227.200 314.270 231.620 314.440 ;
        RECT 231.990 314.330 232.220 315.090 ;
        RECT 232.960 315.080 233.390 315.090 ;
        RECT 232.940 314.910 233.390 315.080 ;
        RECT 232.960 314.890 233.390 314.910 ;
        RECT 238.660 314.630 239.030 329.500 ;
        RECT 238.660 314.380 239.040 314.630 ;
        RECT 230.760 314.160 231.090 314.270 ;
        RECT 231.720 314.160 232.220 314.330 ;
        RECT 232.680 314.160 233.010 314.330 ;
        RECT 233.640 314.160 233.970 314.330 ;
        RECT 22.390 301.190 23.870 301.440 ;
        RECT 24.080 301.250 24.590 314.160 ;
        RECT 30.940 314.150 31.610 314.160 ;
        RECT 27.240 313.260 30.700 313.700 ;
        RECT 25.310 313.160 30.700 313.260 ;
        RECT 25.310 313.090 30.590 313.160 ;
        RECT 25.310 302.180 25.480 313.090 ;
        RECT 25.810 312.680 30.040 312.700 ;
        RECT 25.790 302.570 30.120 312.680 ;
        RECT 25.850 302.520 26.020 302.570 ;
        RECT 30.420 302.180 30.590 313.090 ;
        RECT 25.310 302.010 30.590 302.180 ;
        RECT 30.350 302.000 30.590 302.010 ;
        RECT 31.100 301.250 31.610 314.150 ;
        RECT 231.990 313.760 232.220 314.160 ;
        RECT 228.430 313.590 232.230 313.760 ;
        RECT 230.760 313.480 231.090 313.590 ;
        RECT 231.720 313.480 232.220 313.590 ;
        RECT 227.300 312.810 227.530 312.930 ;
        RECT 227.200 312.640 231.660 312.810 ;
        RECT 231.990 312.720 232.220 313.480 ;
        RECT 232.410 313.210 232.620 313.640 ;
        RECT 232.680 313.480 233.010 313.650 ;
        RECT 233.640 313.480 233.970 313.650 ;
        RECT 232.430 313.190 232.600 313.210 ;
        RECT 230.760 312.550 231.090 312.640 ;
        RECT 231.720 312.550 232.220 312.720 ;
        RECT 232.680 312.550 233.010 312.720 ;
        RECT 233.640 312.550 233.970 312.720 ;
        RECT 231.990 312.150 232.220 312.550 ;
        RECT 228.430 311.980 232.220 312.150 ;
        RECT 230.760 311.870 231.090 311.980 ;
        RECT 231.720 311.870 232.050 311.980 ;
        RECT 232.680 311.900 233.010 312.040 ;
        RECT 232.680 311.870 233.390 311.900 ;
        RECT 233.640 311.870 233.970 312.040 ;
        RECT 232.940 311.710 233.390 311.870 ;
        RECT 232.960 311.690 233.390 311.710 ;
        RECT 229.720 310.170 230.150 310.190 ;
        RECT 230.660 310.170 231.090 310.190 ;
        RECT 232.920 310.170 233.350 310.190 ;
        RECT 229.700 310.000 230.150 310.170 ;
        RECT 230.640 310.000 231.090 310.170 ;
        RECT 231.610 310.150 232.040 310.170 ;
        RECT 229.720 309.980 230.150 310.000 ;
        RECT 230.660 309.980 231.090 310.000 ;
        RECT 231.590 309.980 232.040 310.150 ;
        RECT 232.900 310.000 233.350 310.170 ;
        RECT 232.920 309.980 233.350 310.000 ;
        RECT 231.610 309.960 232.040 309.980 ;
        RECT 24.080 300.740 31.610 301.250 ;
        RECT 22.380 294.720 23.840 294.760 ;
        RECT 22.380 294.550 23.850 294.720 ;
        RECT 22.380 294.510 23.840 294.550 ;
        RECT 24.080 288.130 24.590 300.740 ;
        RECT 24.950 299.950 30.930 300.180 ;
        RECT 25.040 288.890 30.690 299.950 ;
        RECT 31.100 290.380 31.610 300.740 ;
        RECT 31.090 290.360 31.610 290.380 ;
        RECT 25.040 288.880 30.750 288.890 ;
        RECT 24.960 288.710 30.750 288.880 ;
        RECT 25.050 288.700 30.750 288.710 ;
        RECT 30.520 288.630 30.690 288.700 ;
        RECT 31.090 288.580 31.620 290.360 ;
        RECT 31.100 288.560 31.620 288.580 ;
        RECT 24.080 287.840 26.520 288.130 ;
        RECT 31.100 288.050 31.610 288.560 ;
        RECT 31.100 287.840 31.630 288.050 ;
        RECT 24.080 287.360 31.630 287.840 ;
        RECT 24.080 287.330 31.440 287.360 ;
        RECT 24.080 285.570 31.610 286.120 ;
        RECT 22.390 272.600 23.870 272.850 ;
        RECT 24.080 272.660 24.590 285.570 ;
        RECT 30.940 285.560 31.610 285.570 ;
        RECT 27.240 284.670 30.700 285.110 ;
        RECT 25.310 284.570 30.700 284.670 ;
        RECT 25.310 284.500 30.590 284.570 ;
        RECT 25.310 273.590 25.480 284.500 ;
        RECT 25.810 284.090 30.040 284.110 ;
        RECT 25.790 273.980 30.120 284.090 ;
        RECT 25.850 273.930 26.020 273.980 ;
        RECT 30.420 273.590 30.590 284.500 ;
        RECT 25.310 273.420 30.590 273.590 ;
        RECT 30.350 273.410 30.590 273.420 ;
        RECT 31.100 272.660 31.610 285.560 ;
        RECT 24.080 272.150 31.610 272.660 ;
        RECT 22.380 266.130 23.840 266.170 ;
        RECT 22.380 265.960 23.850 266.130 ;
        RECT 22.380 265.920 23.840 265.960 ;
        RECT 24.080 259.540 24.590 272.150 ;
        RECT 24.950 271.360 30.930 271.590 ;
        RECT 25.040 260.300 30.690 271.360 ;
        RECT 31.100 261.790 31.610 272.150 ;
        RECT 31.090 261.770 31.610 261.790 ;
        RECT 384.010 284.850 391.540 285.400 ;
        RECT 384.010 284.840 384.680 284.850 ;
        RECT 384.010 271.940 384.520 284.840 ;
        RECT 384.920 283.950 388.380 284.390 ;
        RECT 384.920 283.850 390.310 283.950 ;
        RECT 385.030 283.780 390.310 283.850 ;
        RECT 385.030 272.870 385.200 283.780 ;
        RECT 385.580 283.370 389.810 283.390 ;
        RECT 385.500 273.260 389.830 283.370 ;
        RECT 389.600 273.210 389.770 273.260 ;
        RECT 390.140 272.870 390.310 283.780 ;
        RECT 385.030 272.700 390.310 272.870 ;
        RECT 385.030 272.690 385.270 272.700 ;
        RECT 391.030 271.940 391.540 284.850 ;
        RECT 384.010 271.430 391.540 271.940 ;
        RECT 391.750 271.880 393.230 272.130 ;
        RECT 25.040 260.290 30.750 260.300 ;
        RECT 24.960 260.120 30.750 260.290 ;
        RECT 25.050 260.110 30.750 260.120 ;
        RECT 30.520 260.040 30.690 260.110 ;
        RECT 31.090 259.990 31.620 261.770 ;
        RECT 384.010 261.070 384.520 271.430 ;
        RECT 384.690 270.640 390.670 270.870 ;
        RECT 384.010 261.050 384.530 261.070 ;
        RECT 31.100 259.970 31.620 259.990 ;
        RECT 24.080 259.250 26.520 259.540 ;
        RECT 31.100 259.460 31.610 259.970 ;
        RECT 31.100 259.250 31.630 259.460 ;
        RECT 384.000 259.270 384.530 261.050 ;
        RECT 384.930 259.580 390.580 270.640 ;
        RECT 384.870 259.570 390.580 259.580 ;
        RECT 384.870 259.400 390.660 259.570 ;
        RECT 384.870 259.390 390.570 259.400 ;
        RECT 384.930 259.320 385.100 259.390 ;
        RECT 384.000 259.250 384.520 259.270 ;
        RECT 24.080 258.770 31.630 259.250 ;
        RECT 24.080 258.740 31.440 258.770 ;
        RECT 384.010 258.740 384.520 259.250 ;
        RECT 391.030 258.820 391.540 271.430 ;
        RECT 391.780 265.410 393.240 265.450 ;
        RECT 391.770 265.240 393.240 265.410 ;
        RECT 391.780 265.200 393.240 265.240 ;
        RECT 383.990 258.530 384.520 258.740 ;
        RECT 389.100 258.530 391.540 258.820 ;
        RECT 383.990 258.050 391.540 258.530 ;
        RECT 384.180 258.020 391.540 258.050 ;
        RECT 24.080 256.980 31.610 257.530 ;
        RECT 22.390 244.010 23.870 244.260 ;
        RECT 24.080 244.070 24.590 256.980 ;
        RECT 30.940 256.970 31.610 256.980 ;
        RECT 27.240 256.080 30.700 256.520 ;
        RECT 25.310 255.980 30.700 256.080 ;
        RECT 25.310 255.910 30.590 255.980 ;
        RECT 25.310 245.000 25.480 255.910 ;
        RECT 25.810 255.500 30.040 255.520 ;
        RECT 25.790 245.390 30.120 255.500 ;
        RECT 25.850 245.340 26.020 245.390 ;
        RECT 30.420 245.000 30.590 255.910 ;
        RECT 25.310 244.830 30.590 245.000 ;
        RECT 30.350 244.820 30.590 244.830 ;
        RECT 31.100 244.070 31.610 256.970 ;
        RECT 24.080 243.560 31.610 244.070 ;
        RECT 22.380 237.540 23.840 237.580 ;
        RECT 22.380 237.370 23.850 237.540 ;
        RECT 22.380 237.330 23.840 237.370 ;
        RECT 24.080 230.950 24.590 243.560 ;
        RECT 24.950 242.770 30.930 243.000 ;
        RECT 25.040 231.710 30.690 242.770 ;
        RECT 31.100 233.200 31.610 243.560 ;
        RECT 31.090 233.180 31.610 233.200 ;
        RECT 384.010 256.260 391.540 256.810 ;
        RECT 384.010 256.250 384.680 256.260 ;
        RECT 384.010 243.350 384.520 256.250 ;
        RECT 384.920 255.360 388.380 255.800 ;
        RECT 384.920 255.260 390.310 255.360 ;
        RECT 385.030 255.190 390.310 255.260 ;
        RECT 385.030 244.280 385.200 255.190 ;
        RECT 385.580 254.780 389.810 254.800 ;
        RECT 385.500 244.670 389.830 254.780 ;
        RECT 389.600 244.620 389.770 244.670 ;
        RECT 390.140 244.280 390.310 255.190 ;
        RECT 385.030 244.110 390.310 244.280 ;
        RECT 385.030 244.100 385.270 244.110 ;
        RECT 391.030 243.350 391.540 256.260 ;
        RECT 384.010 242.840 391.540 243.350 ;
        RECT 391.750 243.290 393.230 243.540 ;
        RECT 25.040 231.700 30.750 231.710 ;
        RECT 24.960 231.530 30.750 231.700 ;
        RECT 25.050 231.520 30.750 231.530 ;
        RECT 30.520 231.450 30.690 231.520 ;
        RECT 31.090 231.400 31.620 233.180 ;
        RECT 384.010 232.480 384.520 242.840 ;
        RECT 384.690 242.050 390.670 242.280 ;
        RECT 384.010 232.460 384.530 232.480 ;
        RECT 31.100 231.380 31.620 231.400 ;
        RECT 24.080 230.660 26.520 230.950 ;
        RECT 31.100 230.870 31.610 231.380 ;
        RECT 31.100 230.660 31.630 230.870 ;
        RECT 384.000 230.680 384.530 232.460 ;
        RECT 384.930 230.990 390.580 242.050 ;
        RECT 384.870 230.980 390.580 230.990 ;
        RECT 384.870 230.810 390.660 230.980 ;
        RECT 384.870 230.800 390.570 230.810 ;
        RECT 384.930 230.730 385.100 230.800 ;
        RECT 384.000 230.660 384.520 230.680 ;
        RECT 24.080 230.180 31.630 230.660 ;
        RECT 24.080 230.150 31.440 230.180 ;
        RECT 384.010 230.150 384.520 230.660 ;
        RECT 391.030 230.230 391.540 242.840 ;
        RECT 391.780 236.820 393.240 236.860 ;
        RECT 391.770 236.650 393.240 236.820 ;
        RECT 391.780 236.610 393.240 236.650 ;
        RECT 383.990 229.940 384.520 230.150 ;
        RECT 389.100 229.940 391.540 230.230 ;
        RECT 383.990 229.460 391.540 229.940 ;
        RECT 384.180 229.430 391.540 229.460 ;
        RECT 24.080 228.390 31.610 228.940 ;
        RECT 22.390 215.420 23.870 215.670 ;
        RECT 24.080 215.480 24.590 228.390 ;
        RECT 30.940 228.380 31.610 228.390 ;
        RECT 27.240 227.490 30.700 227.930 ;
        RECT 25.310 227.390 30.700 227.490 ;
        RECT 25.310 227.320 30.590 227.390 ;
        RECT 25.310 216.410 25.480 227.320 ;
        RECT 25.810 226.910 30.040 226.930 ;
        RECT 25.790 216.800 30.120 226.910 ;
        RECT 25.850 216.750 26.020 216.800 ;
        RECT 30.420 216.410 30.590 227.320 ;
        RECT 25.310 216.240 30.590 216.410 ;
        RECT 30.350 216.230 30.590 216.240 ;
        RECT 31.100 215.480 31.610 228.380 ;
        RECT 24.080 214.970 31.610 215.480 ;
        RECT 22.380 208.950 23.840 208.990 ;
        RECT 22.380 208.780 23.850 208.950 ;
        RECT 22.380 208.740 23.840 208.780 ;
        RECT 24.080 202.360 24.590 214.970 ;
        RECT 24.950 214.180 30.930 214.410 ;
        RECT 25.040 203.120 30.690 214.180 ;
        RECT 31.100 204.610 31.610 214.970 ;
        RECT 31.090 204.590 31.610 204.610 ;
        RECT 384.010 227.670 391.540 228.220 ;
        RECT 384.010 227.660 384.680 227.670 ;
        RECT 384.010 214.760 384.520 227.660 ;
        RECT 384.920 226.770 388.380 227.210 ;
        RECT 384.920 226.670 390.310 226.770 ;
        RECT 385.030 226.600 390.310 226.670 ;
        RECT 385.030 215.690 385.200 226.600 ;
        RECT 385.580 226.190 389.810 226.210 ;
        RECT 385.500 216.080 389.830 226.190 ;
        RECT 389.600 216.030 389.770 216.080 ;
        RECT 390.140 215.690 390.310 226.600 ;
        RECT 385.030 215.520 390.310 215.690 ;
        RECT 385.030 215.510 385.270 215.520 ;
        RECT 391.030 214.760 391.540 227.670 ;
        RECT 384.010 214.250 391.540 214.760 ;
        RECT 391.750 214.700 393.230 214.950 ;
        RECT 25.040 203.110 30.750 203.120 ;
        RECT 24.960 202.940 30.750 203.110 ;
        RECT 25.050 202.930 30.750 202.940 ;
        RECT 30.520 202.860 30.690 202.930 ;
        RECT 31.090 202.810 31.620 204.590 ;
        RECT 384.010 203.890 384.520 214.250 ;
        RECT 384.690 213.460 390.670 213.690 ;
        RECT 384.010 203.870 384.530 203.890 ;
        RECT 31.100 202.790 31.620 202.810 ;
        RECT 24.080 202.070 26.520 202.360 ;
        RECT 31.100 202.280 31.610 202.790 ;
        RECT 31.100 202.070 31.630 202.280 ;
        RECT 384.000 202.090 384.530 203.870 ;
        RECT 384.930 202.400 390.580 213.460 ;
        RECT 384.870 202.390 390.580 202.400 ;
        RECT 384.870 202.220 390.660 202.390 ;
        RECT 384.870 202.210 390.570 202.220 ;
        RECT 384.930 202.140 385.100 202.210 ;
        RECT 384.000 202.070 384.520 202.090 ;
        RECT 24.080 201.590 31.630 202.070 ;
        RECT 24.080 201.560 31.440 201.590 ;
        RECT 384.010 201.560 384.520 202.070 ;
        RECT 391.030 201.640 391.540 214.250 ;
        RECT 391.780 208.230 393.240 208.270 ;
        RECT 391.770 208.060 393.240 208.230 ;
        RECT 391.780 208.020 393.240 208.060 ;
        RECT 383.990 201.350 384.520 201.560 ;
        RECT 389.100 201.350 391.540 201.640 ;
        RECT 383.990 200.870 391.540 201.350 ;
        RECT 384.180 200.840 391.540 200.870 ;
        RECT 24.080 199.800 31.610 200.350 ;
        RECT 22.390 186.830 23.870 187.080 ;
        RECT 24.080 186.890 24.590 199.800 ;
        RECT 30.940 199.790 31.610 199.800 ;
        RECT 27.240 198.900 30.700 199.340 ;
        RECT 25.310 198.800 30.700 198.900 ;
        RECT 25.310 198.730 30.590 198.800 ;
        RECT 25.310 187.820 25.480 198.730 ;
        RECT 25.810 198.320 30.040 198.340 ;
        RECT 25.790 188.210 30.120 198.320 ;
        RECT 25.850 188.160 26.020 188.210 ;
        RECT 30.420 187.820 30.590 198.730 ;
        RECT 25.310 187.650 30.590 187.820 ;
        RECT 30.350 187.640 30.590 187.650 ;
        RECT 31.100 186.890 31.610 199.790 ;
        RECT 24.080 186.380 31.610 186.890 ;
        RECT 22.380 180.360 23.840 180.400 ;
        RECT 22.380 180.190 23.850 180.360 ;
        RECT 22.380 180.150 23.840 180.190 ;
        RECT 24.080 173.770 24.590 186.380 ;
        RECT 24.950 185.590 30.930 185.820 ;
        RECT 25.040 174.530 30.690 185.590 ;
        RECT 31.100 176.020 31.610 186.380 ;
        RECT 31.090 176.000 31.610 176.020 ;
        RECT 384.010 199.080 391.540 199.630 ;
        RECT 384.010 199.070 384.680 199.080 ;
        RECT 384.010 186.170 384.520 199.070 ;
        RECT 384.920 198.180 388.380 198.620 ;
        RECT 384.920 198.080 390.310 198.180 ;
        RECT 385.030 198.010 390.310 198.080 ;
        RECT 385.030 187.100 385.200 198.010 ;
        RECT 385.580 197.600 389.810 197.620 ;
        RECT 385.500 187.490 389.830 197.600 ;
        RECT 389.600 187.440 389.770 187.490 ;
        RECT 390.140 187.100 390.310 198.010 ;
        RECT 385.030 186.930 390.310 187.100 ;
        RECT 385.030 186.920 385.270 186.930 ;
        RECT 391.030 186.170 391.540 199.080 ;
        RECT 384.010 185.660 391.540 186.170 ;
        RECT 391.750 186.110 393.230 186.360 ;
        RECT 25.040 174.520 30.750 174.530 ;
        RECT 24.960 174.350 30.750 174.520 ;
        RECT 25.050 174.340 30.750 174.350 ;
        RECT 30.520 174.270 30.690 174.340 ;
        RECT 31.090 174.220 31.620 176.000 ;
        RECT 384.010 175.300 384.520 185.660 ;
        RECT 384.690 184.870 390.670 185.100 ;
        RECT 384.010 175.280 384.530 175.300 ;
        RECT 31.100 174.200 31.620 174.220 ;
        RECT 24.080 173.480 26.520 173.770 ;
        RECT 31.100 173.690 31.610 174.200 ;
        RECT 31.100 173.480 31.630 173.690 ;
        RECT 384.000 173.500 384.530 175.280 ;
        RECT 384.930 173.810 390.580 184.870 ;
        RECT 384.870 173.800 390.580 173.810 ;
        RECT 384.870 173.630 390.660 173.800 ;
        RECT 384.870 173.620 390.570 173.630 ;
        RECT 384.930 173.550 385.100 173.620 ;
        RECT 384.000 173.480 384.520 173.500 ;
        RECT 24.080 173.000 31.630 173.480 ;
        RECT 24.080 172.970 31.440 173.000 ;
        RECT 384.010 172.970 384.520 173.480 ;
        RECT 391.030 173.050 391.540 185.660 ;
        RECT 391.780 179.640 393.240 179.680 ;
        RECT 391.770 179.470 393.240 179.640 ;
        RECT 391.780 179.430 393.240 179.470 ;
        RECT 383.990 172.760 384.520 172.970 ;
        RECT 389.100 172.760 391.540 173.050 ;
        RECT 383.990 172.280 391.540 172.760 ;
        RECT 384.180 172.250 391.540 172.280 ;
        RECT 24.080 171.210 31.610 171.760 ;
        RECT 22.390 158.240 23.870 158.490 ;
        RECT 24.080 158.300 24.590 171.210 ;
        RECT 30.940 171.200 31.610 171.210 ;
        RECT 27.240 170.310 30.700 170.750 ;
        RECT 25.310 170.210 30.700 170.310 ;
        RECT 25.310 170.140 30.590 170.210 ;
        RECT 25.310 159.230 25.480 170.140 ;
        RECT 25.810 169.730 30.040 169.750 ;
        RECT 25.790 159.620 30.120 169.730 ;
        RECT 25.850 159.570 26.020 159.620 ;
        RECT 30.420 159.230 30.590 170.140 ;
        RECT 25.310 159.060 30.590 159.230 ;
        RECT 30.350 159.050 30.590 159.060 ;
        RECT 31.100 158.300 31.610 171.200 ;
        RECT 24.080 157.790 31.610 158.300 ;
        RECT 22.380 151.770 23.840 151.810 ;
        RECT 22.380 151.600 23.850 151.770 ;
        RECT 22.380 151.560 23.840 151.600 ;
        RECT 24.080 145.180 24.590 157.790 ;
        RECT 24.950 157.000 30.930 157.230 ;
        RECT 25.040 145.940 30.690 157.000 ;
        RECT 31.100 147.430 31.610 157.790 ;
        RECT 31.090 147.410 31.610 147.430 ;
        RECT 384.010 170.490 391.540 171.040 ;
        RECT 384.010 170.480 384.680 170.490 ;
        RECT 384.010 157.580 384.520 170.480 ;
        RECT 384.920 169.590 388.380 170.030 ;
        RECT 384.920 169.490 390.310 169.590 ;
        RECT 385.030 169.420 390.310 169.490 ;
        RECT 385.030 158.510 385.200 169.420 ;
        RECT 385.580 169.010 389.810 169.030 ;
        RECT 385.500 158.900 389.830 169.010 ;
        RECT 389.600 158.850 389.770 158.900 ;
        RECT 390.140 158.510 390.310 169.420 ;
        RECT 385.030 158.340 390.310 158.510 ;
        RECT 385.030 158.330 385.270 158.340 ;
        RECT 391.030 157.580 391.540 170.490 ;
        RECT 384.010 157.070 391.540 157.580 ;
        RECT 391.750 157.520 393.230 157.770 ;
        RECT 25.040 145.930 30.750 145.940 ;
        RECT 24.960 145.760 30.750 145.930 ;
        RECT 25.050 145.750 30.750 145.760 ;
        RECT 30.520 145.680 30.690 145.750 ;
        RECT 31.090 145.630 31.620 147.410 ;
        RECT 384.010 146.710 384.520 157.070 ;
        RECT 384.690 156.280 390.670 156.510 ;
        RECT 384.010 146.690 384.530 146.710 ;
        RECT 31.100 145.610 31.620 145.630 ;
        RECT 24.080 144.890 26.520 145.180 ;
        RECT 31.100 145.100 31.610 145.610 ;
        RECT 31.100 144.890 31.630 145.100 ;
        RECT 384.000 144.910 384.530 146.690 ;
        RECT 384.930 145.220 390.580 156.280 ;
        RECT 384.870 145.210 390.580 145.220 ;
        RECT 384.870 145.040 390.660 145.210 ;
        RECT 384.870 145.030 390.570 145.040 ;
        RECT 384.930 144.960 385.100 145.030 ;
        RECT 384.000 144.890 384.520 144.910 ;
        RECT 24.080 144.410 31.630 144.890 ;
        RECT 24.080 144.380 31.440 144.410 ;
        RECT 384.010 144.380 384.520 144.890 ;
        RECT 391.030 144.460 391.540 157.070 ;
        RECT 391.780 151.050 393.240 151.090 ;
        RECT 391.770 150.880 393.240 151.050 ;
        RECT 391.780 150.840 393.240 150.880 ;
        RECT 383.990 144.170 384.520 144.380 ;
        RECT 389.100 144.170 391.540 144.460 ;
        RECT 383.990 143.690 391.540 144.170 ;
        RECT 384.180 143.660 391.540 143.690 ;
        RECT 24.080 142.620 31.610 143.170 ;
        RECT 22.390 129.650 23.870 129.900 ;
        RECT 24.080 129.710 24.590 142.620 ;
        RECT 30.940 142.610 31.610 142.620 ;
        RECT 27.240 141.720 30.700 142.160 ;
        RECT 25.310 141.620 30.700 141.720 ;
        RECT 25.310 141.550 30.590 141.620 ;
        RECT 25.310 130.640 25.480 141.550 ;
        RECT 25.810 141.140 30.040 141.160 ;
        RECT 25.790 131.030 30.120 141.140 ;
        RECT 25.850 130.980 26.020 131.030 ;
        RECT 30.420 130.640 30.590 141.550 ;
        RECT 25.310 130.470 30.590 130.640 ;
        RECT 30.350 130.460 30.590 130.470 ;
        RECT 31.100 129.710 31.610 142.610 ;
        RECT 24.080 129.200 31.610 129.710 ;
        RECT 22.380 123.180 23.840 123.220 ;
        RECT 22.380 123.010 23.850 123.180 ;
        RECT 22.380 122.970 23.840 123.010 ;
        RECT 24.080 116.590 24.590 129.200 ;
        RECT 24.950 128.410 30.930 128.640 ;
        RECT 25.040 117.350 30.690 128.410 ;
        RECT 31.100 118.840 31.610 129.200 ;
        RECT 31.090 118.820 31.610 118.840 ;
        RECT 384.010 141.900 391.540 142.450 ;
        RECT 384.010 141.890 384.680 141.900 ;
        RECT 384.010 128.990 384.520 141.890 ;
        RECT 384.920 141.000 388.380 141.440 ;
        RECT 384.920 140.900 390.310 141.000 ;
        RECT 385.030 140.830 390.310 140.900 ;
        RECT 385.030 129.920 385.200 140.830 ;
        RECT 385.580 140.420 389.810 140.440 ;
        RECT 385.500 130.310 389.830 140.420 ;
        RECT 389.600 130.260 389.770 130.310 ;
        RECT 390.140 129.920 390.310 140.830 ;
        RECT 385.030 129.750 390.310 129.920 ;
        RECT 385.030 129.740 385.270 129.750 ;
        RECT 391.030 128.990 391.540 141.900 ;
        RECT 384.010 128.480 391.540 128.990 ;
        RECT 391.750 128.930 393.230 129.180 ;
        RECT 25.040 117.340 30.750 117.350 ;
        RECT 24.960 117.170 30.750 117.340 ;
        RECT 25.050 117.160 30.750 117.170 ;
        RECT 30.520 117.090 30.690 117.160 ;
        RECT 31.090 117.040 31.620 118.820 ;
        RECT 384.010 118.120 384.520 128.480 ;
        RECT 384.690 127.690 390.670 127.920 ;
        RECT 384.010 118.100 384.530 118.120 ;
        RECT 31.100 117.020 31.620 117.040 ;
        RECT 24.080 116.300 26.520 116.590 ;
        RECT 31.100 116.510 31.610 117.020 ;
        RECT 31.100 116.300 31.630 116.510 ;
        RECT 384.000 116.320 384.530 118.100 ;
        RECT 384.930 116.630 390.580 127.690 ;
        RECT 384.870 116.620 390.580 116.630 ;
        RECT 384.870 116.450 390.660 116.620 ;
        RECT 384.870 116.440 390.570 116.450 ;
        RECT 384.930 116.370 385.100 116.440 ;
        RECT 384.000 116.300 384.520 116.320 ;
        RECT 24.080 115.820 31.630 116.300 ;
        RECT 24.080 115.790 31.440 115.820 ;
        RECT 384.010 115.790 384.520 116.300 ;
        RECT 391.030 115.870 391.540 128.480 ;
        RECT 391.780 122.460 393.240 122.500 ;
        RECT 391.770 122.290 393.240 122.460 ;
        RECT 391.780 122.250 393.240 122.290 ;
        RECT 383.990 115.580 384.520 115.790 ;
        RECT 389.100 115.580 391.540 115.870 ;
        RECT 383.990 115.100 391.540 115.580 ;
        RECT 384.180 115.070 391.540 115.100 ;
        RECT 24.080 114.030 31.610 114.580 ;
        RECT 22.390 101.060 23.870 101.310 ;
        RECT 24.080 101.120 24.590 114.030 ;
        RECT 30.940 114.020 31.610 114.030 ;
        RECT 27.240 113.130 30.700 113.570 ;
        RECT 25.310 113.030 30.700 113.130 ;
        RECT 25.310 112.960 30.590 113.030 ;
        RECT 25.310 102.050 25.480 112.960 ;
        RECT 25.810 112.550 30.040 112.570 ;
        RECT 25.790 102.440 30.120 112.550 ;
        RECT 25.850 102.390 26.020 102.440 ;
        RECT 30.420 102.050 30.590 112.960 ;
        RECT 25.310 101.880 30.590 102.050 ;
        RECT 30.350 101.870 30.590 101.880 ;
        RECT 31.100 101.120 31.610 114.020 ;
        RECT 24.080 100.610 31.610 101.120 ;
        RECT 22.380 94.590 23.840 94.630 ;
        RECT 22.380 94.420 23.850 94.590 ;
        RECT 22.380 94.380 23.840 94.420 ;
        RECT 24.080 88.000 24.590 100.610 ;
        RECT 24.950 99.820 30.930 100.050 ;
        RECT 25.040 88.760 30.690 99.820 ;
        RECT 31.100 90.250 31.610 100.610 ;
        RECT 31.090 90.230 31.610 90.250 ;
        RECT 384.010 113.310 391.540 113.860 ;
        RECT 384.010 113.300 384.680 113.310 ;
        RECT 384.010 100.400 384.520 113.300 ;
        RECT 384.920 112.410 388.380 112.850 ;
        RECT 384.920 112.310 390.310 112.410 ;
        RECT 385.030 112.240 390.310 112.310 ;
        RECT 385.030 101.330 385.200 112.240 ;
        RECT 385.580 111.830 389.810 111.850 ;
        RECT 385.500 101.720 389.830 111.830 ;
        RECT 389.600 101.670 389.770 101.720 ;
        RECT 390.140 101.330 390.310 112.240 ;
        RECT 385.030 101.160 390.310 101.330 ;
        RECT 385.030 101.150 385.270 101.160 ;
        RECT 391.030 100.400 391.540 113.310 ;
        RECT 384.010 99.890 391.540 100.400 ;
        RECT 391.750 100.340 393.230 100.590 ;
        RECT 25.040 88.750 30.750 88.760 ;
        RECT 24.960 88.580 30.750 88.750 ;
        RECT 25.050 88.570 30.750 88.580 ;
        RECT 30.520 88.500 30.690 88.570 ;
        RECT 31.090 88.450 31.620 90.230 ;
        RECT 384.010 89.530 384.520 99.890 ;
        RECT 384.690 99.100 390.670 99.330 ;
        RECT 384.010 89.510 384.530 89.530 ;
        RECT 31.100 88.430 31.620 88.450 ;
        RECT 24.080 87.710 26.520 88.000 ;
        RECT 31.100 87.920 31.610 88.430 ;
        RECT 31.100 87.710 31.630 87.920 ;
        RECT 384.000 87.730 384.530 89.510 ;
        RECT 384.930 88.040 390.580 99.100 ;
        RECT 384.870 88.030 390.580 88.040 ;
        RECT 384.870 87.860 390.660 88.030 ;
        RECT 384.870 87.850 390.570 87.860 ;
        RECT 384.930 87.780 385.100 87.850 ;
        RECT 384.000 87.710 384.520 87.730 ;
        RECT 24.080 87.230 31.630 87.710 ;
        RECT 24.080 87.200 31.440 87.230 ;
        RECT 384.010 87.200 384.520 87.710 ;
        RECT 391.030 87.280 391.540 99.890 ;
        RECT 391.780 93.870 393.240 93.910 ;
        RECT 391.770 93.700 393.240 93.870 ;
        RECT 391.780 93.660 393.240 93.700 ;
        RECT 383.990 86.990 384.520 87.200 ;
        RECT 389.100 86.990 391.540 87.280 ;
        RECT 383.990 86.510 391.540 86.990 ;
        RECT 384.180 86.480 391.540 86.510 ;
      LAYER mcon ;
        RECT 24.480 457.290 25.410 457.490 ;
        RECT 24.250 453.720 24.430 456.880 ;
        RECT 27.350 456.220 30.650 456.570 ;
        RECT 22.410 444.180 22.580 444.350 ;
        RECT 22.770 444.180 22.940 444.350 ;
        RECT 23.130 444.180 23.300 444.350 ;
        RECT 23.490 444.180 23.660 444.350 ;
        RECT 26.140 445.720 26.310 455.170 ;
        RECT 26.890 445.710 27.060 455.100 ;
        RECT 27.610 445.740 27.780 455.140 ;
        RECT 28.270 445.750 28.440 455.120 ;
        RECT 28.920 445.740 29.090 455.190 ;
        RECT 29.560 445.750 29.730 455.140 ;
        RECT 22.730 437.500 22.900 437.670 ;
        RECT 23.090 437.500 23.260 437.670 ;
        RECT 23.460 437.500 23.630 437.670 ;
        RECT 24.250 432.220 24.420 432.230 ;
        RECT 24.240 430.360 24.420 432.220 ;
        RECT 25.380 431.990 25.550 442.970 ;
        RECT 26.000 431.990 26.170 442.970 ;
        RECT 26.620 432.000 26.790 442.980 ;
        RECT 27.200 432.020 27.370 443.000 ;
        RECT 27.790 432.030 27.960 443.010 ;
        RECT 28.390 432.030 28.560 443.010 ;
        RECT 28.990 431.980 29.160 442.960 ;
        RECT 29.600 431.990 29.770 442.970 ;
        RECT 30.200 431.980 30.370 442.960 ;
        RECT 24.610 430.800 26.520 430.980 ;
        RECT 24.610 430.400 26.510 430.580 ;
        RECT 24.480 428.700 25.410 428.900 ;
        RECT 24.250 425.130 24.430 428.290 ;
        RECT 27.350 427.630 30.650 427.980 ;
        RECT 22.410 415.590 22.580 415.760 ;
        RECT 22.770 415.590 22.940 415.760 ;
        RECT 23.130 415.590 23.300 415.760 ;
        RECT 23.490 415.590 23.660 415.760 ;
        RECT 26.140 417.130 26.310 426.580 ;
        RECT 26.890 417.120 27.060 426.510 ;
        RECT 27.610 417.150 27.780 426.550 ;
        RECT 28.270 417.160 28.440 426.530 ;
        RECT 28.920 417.150 29.090 426.600 ;
        RECT 29.560 417.160 29.730 426.550 ;
        RECT 22.730 408.910 22.900 409.080 ;
        RECT 23.090 408.910 23.260 409.080 ;
        RECT 23.460 408.910 23.630 409.080 ;
        RECT 24.250 403.630 24.420 403.640 ;
        RECT 24.240 401.770 24.420 403.630 ;
        RECT 25.380 403.400 25.550 414.380 ;
        RECT 26.000 403.400 26.170 414.380 ;
        RECT 26.620 403.410 26.790 414.390 ;
        RECT 27.200 403.430 27.370 414.410 ;
        RECT 27.790 403.440 27.960 414.420 ;
        RECT 28.390 403.440 28.560 414.420 ;
        RECT 28.990 403.390 29.160 414.370 ;
        RECT 29.600 403.400 29.770 414.380 ;
        RECT 30.200 403.390 30.370 414.370 ;
        RECT 24.610 402.210 26.520 402.390 ;
        RECT 24.610 401.810 26.510 401.990 ;
        RECT 24.480 400.110 25.410 400.310 ;
        RECT 24.250 396.540 24.430 399.700 ;
        RECT 27.350 399.040 30.650 399.390 ;
        RECT 23.700 389.160 23.870 389.330 ;
        RECT 23.700 388.800 23.870 388.970 ;
        RECT 23.700 388.430 23.870 388.600 ;
        RECT 26.140 388.540 26.310 397.990 ;
        RECT 26.890 388.530 27.060 397.920 ;
        RECT 27.610 388.560 27.780 397.960 ;
        RECT 28.270 388.570 28.440 397.940 ;
        RECT 28.920 388.560 29.090 398.010 ;
        RECT 29.560 388.570 29.730 397.960 ;
        RECT 30.380 389.480 30.550 389.650 ;
        RECT 30.380 389.120 30.550 389.290 ;
        RECT 30.380 388.760 30.550 388.930 ;
        RECT 30.380 388.400 30.550 388.570 ;
        RECT 52.290 389.160 52.460 389.330 ;
        RECT 52.290 388.800 52.460 388.970 ;
        RECT 52.290 388.430 52.460 388.600 ;
        RECT 58.970 389.480 59.140 389.650 ;
        RECT 58.970 389.120 59.140 389.290 ;
        RECT 58.970 388.760 59.140 388.930 ;
        RECT 58.970 388.400 59.140 388.570 ;
        RECT 80.880 389.160 81.050 389.330 ;
        RECT 80.880 388.800 81.050 388.970 ;
        RECT 80.880 388.430 81.050 388.600 ;
        RECT 87.560 389.480 87.730 389.650 ;
        RECT 87.560 389.120 87.730 389.290 ;
        RECT 87.560 388.760 87.730 388.930 ;
        RECT 87.560 388.400 87.730 388.570 ;
        RECT 164.900 389.160 165.070 389.330 ;
        RECT 164.900 388.800 165.070 388.970 ;
        RECT 164.900 388.430 165.070 388.600 ;
        RECT 171.580 389.480 171.750 389.650 ;
        RECT 171.580 389.120 171.750 389.290 ;
        RECT 171.580 388.760 171.750 388.930 ;
        RECT 171.580 388.400 171.750 388.570 ;
        RECT 193.490 389.160 193.660 389.330 ;
        RECT 193.490 388.800 193.660 388.970 ;
        RECT 193.490 388.430 193.660 388.600 ;
        RECT 200.170 389.480 200.340 389.650 ;
        RECT 200.170 389.120 200.340 389.290 ;
        RECT 200.170 388.760 200.340 388.930 ;
        RECT 200.170 388.400 200.340 388.570 ;
        RECT 222.080 389.160 222.250 389.330 ;
        RECT 222.080 388.800 222.250 388.970 ;
        RECT 222.080 388.430 222.250 388.600 ;
        RECT 228.760 389.480 228.930 389.650 ;
        RECT 228.760 389.120 228.930 389.290 ;
        RECT 228.760 388.760 228.930 388.930 ;
        RECT 228.760 388.400 228.930 388.570 ;
        RECT 250.670 389.160 250.840 389.330 ;
        RECT 250.670 388.800 250.840 388.970 ;
        RECT 250.670 388.430 250.840 388.600 ;
        RECT 257.350 389.480 257.520 389.650 ;
        RECT 257.350 389.120 257.520 389.290 ;
        RECT 257.350 388.760 257.520 388.930 ;
        RECT 257.350 388.400 257.520 388.570 ;
        RECT 279.260 389.160 279.430 389.330 ;
        RECT 279.260 388.800 279.430 388.970 ;
        RECT 279.260 388.430 279.430 388.600 ;
        RECT 285.940 389.480 286.110 389.650 ;
        RECT 285.940 389.120 286.110 389.290 ;
        RECT 285.940 388.760 286.110 388.930 ;
        RECT 285.940 388.400 286.110 388.570 ;
        RECT 307.850 389.160 308.020 389.330 ;
        RECT 307.850 388.800 308.020 388.970 ;
        RECT 307.850 388.430 308.020 388.600 ;
        RECT 314.530 389.480 314.700 389.650 ;
        RECT 314.530 389.120 314.700 389.290 ;
        RECT 314.530 388.760 314.700 388.930 ;
        RECT 314.530 388.400 314.700 388.570 ;
        RECT 336.440 389.160 336.610 389.330 ;
        RECT 336.440 388.800 336.610 388.970 ;
        RECT 336.440 388.430 336.610 388.600 ;
        RECT 343.120 389.480 343.290 389.650 ;
        RECT 343.120 389.120 343.290 389.290 ;
        RECT 343.120 388.760 343.290 388.930 ;
        RECT 343.120 388.400 343.290 388.570 ;
        RECT 16.560 387.810 18.420 387.820 ;
        RECT 16.560 387.640 18.430 387.810 ;
        RECT 39.920 387.630 43.080 387.810 ;
        RECT 16.600 385.550 16.780 387.450 ;
        RECT 17.000 385.540 17.180 387.450 ;
        RECT 22.410 387.000 22.580 387.170 ;
        RECT 22.770 387.000 22.940 387.170 ;
        RECT 23.130 387.000 23.300 387.170 ;
        RECT 23.490 387.000 23.660 387.170 ;
        RECT 18.190 386.510 29.170 386.680 ;
        RECT 18.190 385.890 29.170 386.060 ;
        RECT 25.380 385.440 25.550 385.790 ;
        RECT 26.000 385.440 26.170 385.790 ;
        RECT 26.620 385.440 26.790 385.800 ;
        RECT 27.200 385.440 27.370 385.820 ;
        RECT 27.790 385.440 27.960 385.830 ;
        RECT 28.390 385.440 28.560 385.830 ;
        RECT 28.990 385.440 29.160 385.780 ;
        RECT 18.200 385.270 29.180 385.440 ;
        RECT 25.380 384.860 25.550 385.270 ;
        RECT 26.000 384.860 26.170 385.270 ;
        RECT 26.620 384.860 26.790 385.270 ;
        RECT 27.200 384.860 27.370 385.270 ;
        RECT 27.790 384.860 27.960 385.270 ;
        RECT 28.390 384.860 28.560 385.270 ;
        RECT 28.990 384.860 29.160 385.270 ;
        RECT 18.220 384.690 29.200 384.860 ;
        RECT 25.380 384.270 25.550 384.690 ;
        RECT 26.000 384.270 26.170 384.690 ;
        RECT 26.620 384.270 26.790 384.690 ;
        RECT 27.200 384.270 27.370 384.690 ;
        RECT 27.790 384.270 27.960 384.690 ;
        RECT 28.390 384.270 28.560 384.690 ;
        RECT 28.990 384.270 29.160 384.690 ;
        RECT 18.230 384.100 29.210 384.270 ;
        RECT 25.380 383.670 25.550 384.100 ;
        RECT 26.000 383.670 26.170 384.100 ;
        RECT 26.620 383.670 26.790 384.100 ;
        RECT 27.200 383.670 27.370 384.100 ;
        RECT 27.790 383.670 27.960 384.100 ;
        RECT 28.390 383.670 28.560 384.100 ;
        RECT 28.990 383.670 29.160 384.100 ;
        RECT 18.230 383.500 29.210 383.670 ;
        RECT 25.380 383.070 25.550 383.500 ;
        RECT 26.000 383.070 26.170 383.500 ;
        RECT 26.620 383.070 26.790 383.500 ;
        RECT 27.200 383.070 27.370 383.500 ;
        RECT 27.790 383.070 27.960 383.500 ;
        RECT 28.390 383.070 28.560 383.500 ;
        RECT 28.990 383.070 29.160 383.500 ;
        RECT 18.180 382.900 29.160 383.070 ;
        RECT 25.380 382.460 25.550 382.900 ;
        RECT 26.000 382.460 26.170 382.900 ;
        RECT 26.620 382.460 26.790 382.900 ;
        RECT 27.200 382.460 27.370 382.900 ;
        RECT 27.790 382.460 27.960 382.900 ;
        RECT 28.390 382.460 28.560 382.900 ;
        RECT 28.990 382.460 29.160 382.900 ;
        RECT 18.190 382.290 29.170 382.460 ;
        RECT 25.380 381.860 25.550 382.290 ;
        RECT 26.000 381.860 26.170 382.290 ;
        RECT 26.620 381.860 26.790 382.290 ;
        RECT 27.200 381.860 27.370 382.290 ;
        RECT 27.790 381.860 27.960 382.290 ;
        RECT 28.390 381.860 28.560 382.290 ;
        RECT 28.990 381.860 29.160 382.290 ;
        RECT 18.180 381.690 29.160 381.860 ;
        RECT 22.730 380.320 22.900 380.490 ;
        RECT 23.090 380.320 23.260 380.490 ;
        RECT 23.460 380.320 23.630 380.490 ;
        RECT 24.250 375.040 24.420 375.050 ;
        RECT 24.240 373.180 24.420 375.040 ;
        RECT 25.380 374.810 25.550 381.690 ;
        RECT 26.000 374.810 26.170 381.690 ;
        RECT 26.620 374.820 26.790 381.690 ;
        RECT 27.200 374.840 27.370 381.690 ;
        RECT 27.790 374.850 27.960 381.690 ;
        RECT 28.390 374.850 28.560 381.690 ;
        RECT 28.990 374.800 29.160 381.690 ;
        RECT 29.600 374.810 29.770 385.790 ;
        RECT 30.200 374.800 30.370 385.780 ;
        RECT 31.920 385.750 41.370 385.920 ;
        RECT 31.910 385.000 41.300 385.170 ;
        RECT 31.940 384.280 41.340 384.450 ;
        RECT 31.950 383.620 41.320 383.790 ;
        RECT 31.940 382.970 41.390 383.140 ;
        RECT 31.950 382.330 41.340 382.500 ;
        RECT 43.490 386.650 43.690 387.580 ;
        RECT 42.420 381.410 42.770 384.710 ;
        RECT 45.150 387.810 47.010 387.820 ;
        RECT 45.150 387.640 47.020 387.810 ;
        RECT 68.510 387.630 71.670 387.810 ;
        RECT 45.190 385.550 45.370 387.450 ;
        RECT 45.590 385.540 45.770 387.450 ;
        RECT 46.780 386.510 57.760 386.680 ;
        RECT 46.780 385.890 57.760 386.060 ;
        RECT 46.790 385.270 57.770 385.440 ;
        RECT 46.810 384.690 57.790 384.860 ;
        RECT 46.820 384.100 57.800 384.270 ;
        RECT 46.820 383.500 57.800 383.670 ;
        RECT 46.770 382.900 57.750 383.070 ;
        RECT 46.780 382.290 57.760 382.460 ;
        RECT 46.770 381.690 57.750 381.860 ;
        RECT 60.510 385.750 69.960 385.920 ;
        RECT 60.500 385.000 69.890 385.170 ;
        RECT 60.530 384.280 69.930 384.450 ;
        RECT 60.540 383.620 69.910 383.790 ;
        RECT 60.530 382.970 69.980 383.140 ;
        RECT 60.540 382.330 69.930 382.500 ;
        RECT 72.080 386.650 72.280 387.580 ;
        RECT 71.010 381.410 71.360 384.710 ;
        RECT 73.740 387.810 75.600 387.820 ;
        RECT 73.740 387.640 75.610 387.810 ;
        RECT 97.100 387.630 100.260 387.810 ;
        RECT 73.780 385.550 73.960 387.450 ;
        RECT 74.180 385.540 74.360 387.450 ;
        RECT 75.370 386.510 86.350 386.680 ;
        RECT 75.370 385.890 86.350 386.060 ;
        RECT 75.380 385.270 86.360 385.440 ;
        RECT 75.400 384.690 86.380 384.860 ;
        RECT 75.410 384.100 86.390 384.270 ;
        RECT 75.410 383.500 86.390 383.670 ;
        RECT 75.360 382.900 86.340 383.070 ;
        RECT 75.370 382.290 86.350 382.460 ;
        RECT 75.360 381.690 86.340 381.860 ;
        RECT 89.100 385.750 98.550 385.920 ;
        RECT 89.090 385.000 98.480 385.170 ;
        RECT 89.120 384.280 98.520 384.450 ;
        RECT 89.130 383.620 98.500 383.790 ;
        RECT 89.120 382.970 98.570 383.140 ;
        RECT 89.130 382.330 98.520 382.500 ;
        RECT 100.670 386.650 100.870 387.580 ;
        RECT 142.870 387.610 143.040 387.780 ;
        RECT 142.870 387.250 143.040 387.420 ;
        RECT 142.870 386.890 143.040 387.060 ;
        RECT 99.600 381.410 99.950 384.710 ;
        RECT 142.870 386.530 143.040 386.700 ;
        RECT 149.620 387.440 149.790 387.610 ;
        RECT 149.620 387.080 149.790 387.250 ;
        RECT 149.620 386.720 149.790 386.890 ;
        RECT 157.760 387.810 159.620 387.820 ;
        RECT 157.760 387.640 159.630 387.810 ;
        RECT 181.120 387.630 184.280 387.810 ;
        RECT 157.800 386.090 157.980 387.450 ;
        RECT 158.200 386.090 158.380 387.450 ;
        RECT 159.390 386.510 170.370 386.680 ;
        RECT 122.420 385.920 146.320 386.090 ;
        RECT 155.200 385.920 176.370 386.090 ;
        RECT 157.800 385.550 157.980 385.920 ;
        RECT 158.200 385.540 158.380 385.920 ;
        RECT 159.390 385.890 170.370 385.920 ;
        RECT 125.240 381.730 125.410 381.900 ;
        RECT 139.930 382.140 140.100 382.310 ;
        RECT 139.930 381.690 140.100 381.860 ;
        RECT 144.630 382.090 144.800 382.260 ;
        RECT 144.630 381.640 144.800 381.810 ;
        RECT 159.400 385.270 170.380 385.440 ;
        RECT 159.420 384.690 170.400 384.860 ;
        RECT 159.430 384.100 170.410 384.270 ;
        RECT 159.430 383.500 170.410 383.670 ;
        RECT 159.380 382.900 170.360 383.070 ;
        RECT 159.390 382.290 170.370 382.460 ;
        RECT 159.380 381.690 170.360 381.860 ;
        RECT 173.120 385.750 182.570 385.920 ;
        RECT 173.110 385.000 182.500 385.170 ;
        RECT 173.140 384.280 182.540 384.450 ;
        RECT 173.150 383.620 182.520 383.790 ;
        RECT 173.140 382.970 182.590 383.140 ;
        RECT 173.150 382.330 182.540 382.500 ;
        RECT 184.690 386.650 184.890 387.580 ;
        RECT 183.620 381.410 183.970 384.710 ;
        RECT 186.350 387.810 188.210 387.820 ;
        RECT 186.350 387.640 188.220 387.810 ;
        RECT 209.710 387.630 212.870 387.810 ;
        RECT 186.390 385.550 186.570 387.450 ;
        RECT 186.790 385.540 186.970 387.450 ;
        RECT 187.980 386.510 198.960 386.680 ;
        RECT 187.980 385.890 198.960 386.060 ;
        RECT 187.990 385.270 198.970 385.440 ;
        RECT 188.010 384.690 198.990 384.860 ;
        RECT 188.020 384.100 199.000 384.270 ;
        RECT 188.020 383.500 199.000 383.670 ;
        RECT 187.970 382.900 198.950 383.070 ;
        RECT 187.980 382.290 198.960 382.460 ;
        RECT 187.970 381.690 198.950 381.860 ;
        RECT 201.710 385.750 211.160 385.920 ;
        RECT 201.700 385.000 211.090 385.170 ;
        RECT 201.730 384.280 211.130 384.450 ;
        RECT 201.740 383.620 211.110 383.790 ;
        RECT 201.730 382.970 211.180 383.140 ;
        RECT 201.740 382.330 211.130 382.500 ;
        RECT 213.280 386.650 213.480 387.580 ;
        RECT 212.210 381.410 212.560 384.710 ;
        RECT 211.540 380.950 211.810 381.220 ;
        RECT 214.940 387.810 216.800 387.820 ;
        RECT 214.940 387.640 216.810 387.810 ;
        RECT 238.300 387.630 241.460 387.810 ;
        RECT 214.980 385.550 215.160 387.450 ;
        RECT 215.380 385.540 215.560 387.450 ;
        RECT 216.570 386.510 227.550 386.680 ;
        RECT 216.570 385.890 227.550 386.060 ;
        RECT 216.580 385.270 227.560 385.440 ;
        RECT 216.600 384.690 227.580 384.860 ;
        RECT 216.610 384.100 227.590 384.270 ;
        RECT 216.610 383.500 227.590 383.670 ;
        RECT 216.560 382.900 227.540 383.070 ;
        RECT 216.570 382.290 227.550 382.460 ;
        RECT 216.560 381.690 227.540 381.860 ;
        RECT 230.300 385.750 239.750 385.920 ;
        RECT 230.290 385.000 239.680 385.170 ;
        RECT 230.320 384.280 239.720 384.450 ;
        RECT 230.330 383.620 239.700 383.790 ;
        RECT 230.320 382.970 239.770 383.140 ;
        RECT 230.330 382.330 239.720 382.500 ;
        RECT 241.870 386.650 242.070 387.580 ;
        RECT 240.800 381.410 241.150 384.710 ;
        RECT 243.530 387.810 245.390 387.820 ;
        RECT 243.530 387.640 245.400 387.810 ;
        RECT 266.890 387.630 270.050 387.810 ;
        RECT 243.570 385.550 243.750 387.450 ;
        RECT 243.970 385.540 244.150 387.450 ;
        RECT 245.160 386.510 256.140 386.680 ;
        RECT 245.160 385.890 256.140 386.060 ;
        RECT 245.170 385.270 256.150 385.440 ;
        RECT 245.190 384.690 256.170 384.860 ;
        RECT 245.200 384.100 256.180 384.270 ;
        RECT 245.200 383.500 256.180 383.670 ;
        RECT 245.150 382.900 256.130 383.070 ;
        RECT 245.160 382.290 256.140 382.460 ;
        RECT 245.150 381.690 256.130 381.860 ;
        RECT 255.760 380.950 256.030 381.220 ;
        RECT 258.890 385.750 268.340 385.920 ;
        RECT 258.880 385.000 268.270 385.170 ;
        RECT 258.910 384.280 268.310 384.450 ;
        RECT 258.920 383.620 268.290 383.790 ;
        RECT 258.910 382.970 268.360 383.140 ;
        RECT 258.920 382.330 268.310 382.500 ;
        RECT 270.460 386.650 270.660 387.580 ;
        RECT 269.390 381.410 269.740 384.710 ;
        RECT 272.120 387.810 273.980 387.820 ;
        RECT 272.120 387.640 273.990 387.810 ;
        RECT 295.480 387.630 298.640 387.810 ;
        RECT 272.160 385.550 272.340 387.450 ;
        RECT 272.560 385.540 272.740 387.450 ;
        RECT 273.750 386.510 284.730 386.680 ;
        RECT 273.750 385.890 284.730 386.060 ;
        RECT 273.760 385.270 284.740 385.440 ;
        RECT 273.780 384.690 284.760 384.860 ;
        RECT 273.790 384.100 284.770 384.270 ;
        RECT 273.790 383.500 284.770 383.670 ;
        RECT 273.740 382.900 284.720 383.070 ;
        RECT 273.750 382.290 284.730 382.460 ;
        RECT 273.740 381.690 284.720 381.860 ;
        RECT 287.480 385.750 296.930 385.920 ;
        RECT 287.470 385.000 296.860 385.170 ;
        RECT 287.500 384.280 296.900 384.450 ;
        RECT 287.510 383.620 296.880 383.790 ;
        RECT 287.500 382.970 296.950 383.140 ;
        RECT 287.510 382.330 296.900 382.500 ;
        RECT 299.050 386.650 299.250 387.580 ;
        RECT 297.980 381.410 298.330 384.710 ;
        RECT 300.710 387.810 302.570 387.820 ;
        RECT 300.710 387.640 302.580 387.810 ;
        RECT 324.070 387.630 327.230 387.810 ;
        RECT 300.750 385.550 300.930 387.450 ;
        RECT 301.150 385.540 301.330 387.450 ;
        RECT 302.340 386.510 313.320 386.680 ;
        RECT 302.340 385.890 313.320 386.060 ;
        RECT 302.350 385.270 313.330 385.440 ;
        RECT 302.370 384.690 313.350 384.860 ;
        RECT 302.380 384.100 313.360 384.270 ;
        RECT 302.380 383.500 313.360 383.670 ;
        RECT 302.330 382.900 313.310 383.070 ;
        RECT 302.340 382.290 313.320 382.460 ;
        RECT 302.330 381.690 313.310 381.860 ;
        RECT 316.070 385.750 325.520 385.920 ;
        RECT 316.060 385.000 325.450 385.170 ;
        RECT 316.090 384.280 325.490 384.450 ;
        RECT 316.100 383.620 325.470 383.790 ;
        RECT 316.090 382.970 325.540 383.140 ;
        RECT 316.100 382.330 325.490 382.500 ;
        RECT 327.640 386.650 327.840 387.580 ;
        RECT 326.570 381.410 326.920 384.710 ;
        RECT 329.300 387.810 331.160 387.820 ;
        RECT 329.300 387.640 331.170 387.810 ;
        RECT 352.660 387.630 355.820 387.810 ;
        RECT 329.340 385.550 329.520 387.450 ;
        RECT 329.740 385.540 329.920 387.450 ;
        RECT 330.930 386.510 341.910 386.680 ;
        RECT 330.930 385.890 341.910 386.060 ;
        RECT 330.940 385.270 341.920 385.440 ;
        RECT 330.960 384.690 341.940 384.860 ;
        RECT 330.970 384.100 341.950 384.270 ;
        RECT 330.970 383.500 341.950 383.670 ;
        RECT 330.920 382.900 341.900 383.070 ;
        RECT 330.930 382.290 341.910 382.460 ;
        RECT 330.920 381.690 341.900 381.860 ;
        RECT 344.660 385.750 354.110 385.920 ;
        RECT 344.650 385.000 354.040 385.170 ;
        RECT 344.680 384.280 354.080 384.450 ;
        RECT 344.690 383.620 354.060 383.790 ;
        RECT 344.680 382.970 354.130 383.140 ;
        RECT 344.690 382.330 354.080 382.500 ;
        RECT 356.230 386.650 356.430 387.580 ;
        RECT 355.160 381.410 355.510 384.710 ;
        RECT 139.930 379.150 140.100 379.320 ;
        RECT 138.910 378.970 139.080 379.140 ;
        RECT 128.780 378.610 128.950 378.780 ;
        RECT 139.930 378.700 140.100 378.870 ;
        RECT 211.540 379.220 211.810 379.490 ;
        RECT 255.760 379.220 256.030 379.490 ;
        RECT 125.910 378.400 126.080 378.570 ;
        RECT 127.320 378.400 127.490 378.570 ;
        RECT 138.910 378.280 139.080 378.450 ;
        RECT 212.670 378.440 212.850 378.610 ;
        RECT 139.930 378.140 140.100 378.310 ;
        RECT 210.860 378.140 211.030 378.310 ;
        RECT 148.890 377.960 149.060 378.130 ;
        RECT 149.260 377.960 149.430 378.130 ;
        RECT 149.620 377.960 149.790 378.130 ;
        RECT 149.980 377.960 150.150 378.130 ;
        RECT 150.340 377.960 150.520 378.130 ;
        RECT 150.710 377.960 150.880 378.130 ;
        RECT 125.910 377.550 126.080 377.720 ;
        RECT 126.490 377.690 126.660 377.860 ;
        RECT 127.320 377.550 127.490 377.720 ;
        RECT 128.520 377.690 128.690 377.860 ;
        RECT 139.930 377.690 140.100 377.860 ;
        RECT 217.760 378.080 217.930 378.250 ;
        RECT 126.090 377.140 126.260 377.310 ;
        RECT 127.150 377.140 127.320 377.310 ;
        RECT 125.910 376.730 126.080 376.900 ;
        RECT 126.490 376.850 126.660 377.020 ;
        RECT 141.880 376.950 142.050 377.120 ;
        RECT 211.210 377.300 211.390 377.490 ;
        RECT 143.240 377.030 143.410 377.200 ;
        RECT 127.320 376.730 127.490 376.900 ;
        RECT 143.930 377.020 144.100 377.190 ;
        RECT 128.520 376.260 128.690 376.430 ;
        RECT 138.910 376.170 139.080 376.340 ;
        RECT 125.910 375.890 126.080 376.060 ;
        RECT 127.320 375.890 127.490 376.060 ;
        RECT 127.950 375.710 128.120 375.880 ;
        RECT 138.910 375.480 139.080 375.650 ;
        RECT 125.910 374.770 126.080 374.940 ;
        RECT 128.180 374.960 128.350 375.130 ;
        RECT 128.790 374.990 128.960 375.160 ;
        RECT 127.320 374.770 127.490 374.940 ;
        RECT 138.910 374.620 139.080 374.790 ;
        RECT 24.610 373.620 26.520 373.800 ;
        RECT 126.470 374.050 126.640 374.220 ;
        RECT 127.900 374.070 128.070 374.240 ;
        RECT 138.910 373.930 139.080 374.100 ;
        RECT 218.230 377.520 218.400 377.690 ;
        RECT 230.620 377.990 230.790 378.160 ;
        RECT 230.620 377.540 230.790 377.710 ;
        RECT 254.990 377.990 255.160 378.160 ;
        RECT 256.540 378.140 256.710 378.310 ;
        RECT 254.990 377.540 255.160 377.710 ;
        RECT 250.250 377.040 250.420 377.210 ;
        RECT 216.910 376.470 217.080 376.640 ;
        RECT 256.180 377.300 256.360 377.490 ;
        RECT 217.760 376.090 217.930 376.260 ;
        RECT 125.680 373.470 125.850 373.640 ;
        RECT 126.610 373.470 126.780 373.640 ;
        RECT 127.310 373.470 127.480 373.640 ;
        RECT 128.050 373.470 128.220 373.640 ;
        RECT 128.760 373.460 128.930 373.630 ;
        RECT 153.280 375.260 153.450 375.430 ;
        RECT 211.790 374.920 212.060 375.190 ;
        RECT 217.770 375.020 217.940 375.190 ;
        RECT 218.230 375.200 218.400 375.370 ;
        RECT 223.600 375.510 223.770 375.680 ;
        RECT 243.800 375.510 243.970 375.680 ;
        RECT 211.210 373.660 211.390 373.850 ;
        RECT 24.610 373.220 26.510 373.400 ;
        RECT 141.160 373.290 141.330 373.460 ;
        RECT 151.020 373.310 151.190 373.480 ;
        RECT 211.790 373.190 212.060 373.460 ;
        RECT 216.900 374.780 217.070 374.950 ;
        RECT 249.720 374.920 249.990 375.190 ;
        RECT 252.790 375.110 252.960 375.280 ;
        RECT 254.450 375.070 254.620 375.240 ;
        RECT 250.250 374.280 250.420 374.450 ;
        RECT 252.740 374.460 252.910 374.630 ;
        RECT 253.730 374.720 253.900 374.890 ;
        RECT 218.220 373.620 218.390 373.790 ;
        RECT 253.800 373.690 253.970 373.860 ;
        RECT 217.790 373.110 217.960 373.280 ;
        RECT 230.620 373.340 230.790 373.510 ;
        RECT 249.720 373.190 249.990 373.460 ;
        RECT 252.740 373.200 252.910 373.370 ;
        RECT 210.860 372.840 211.030 373.010 ;
        RECT 230.620 372.890 230.790 373.060 ;
        RECT 253.730 372.940 253.900 373.110 ;
        RECT 254.990 373.340 255.160 373.510 ;
        RECT 212.670 372.540 212.850 372.710 ;
        RECT 212.920 372.410 213.100 372.580 ;
        RECT 24.480 371.520 25.410 371.720 ;
        RECT 150.150 371.370 150.580 372.110 ;
        RECT 173.510 371.940 173.720 372.150 ;
        RECT 211.110 372.110 211.280 372.280 ;
        RECT 172.040 371.570 172.210 371.740 ;
        RECT 174.470 371.470 174.640 371.640 ;
        RECT 24.250 367.950 24.430 371.110 ;
        RECT 27.350 370.450 30.650 370.800 ;
        RECT 22.410 358.410 22.580 358.580 ;
        RECT 22.770 358.410 22.940 358.580 ;
        RECT 23.130 358.410 23.300 358.580 ;
        RECT 23.490 358.410 23.660 358.580 ;
        RECT 26.140 359.950 26.310 369.400 ;
        RECT 26.890 359.940 27.060 369.330 ;
        RECT 27.610 359.970 27.780 369.370 ;
        RECT 28.270 359.980 28.440 369.350 ;
        RECT 28.920 359.970 29.090 369.420 ;
        RECT 29.560 359.980 29.730 369.370 ;
        RECT 175.510 371.510 175.680 371.680 ;
        RECT 176.550 371.170 176.720 371.340 ;
        RECT 211.460 371.270 211.640 371.460 ;
        RECT 176.550 370.810 176.720 370.980 ;
        RECT 212.660 371.960 212.830 372.130 ;
        RECT 212.660 371.510 212.830 371.680 ;
        RECT 252.790 372.550 252.960 372.720 ;
        RECT 256.180 373.660 256.360 373.850 ;
        RECT 254.500 372.850 254.670 373.020 ;
        RECT 254.990 372.890 255.160 373.060 ;
        RECT 256.540 372.840 256.710 373.010 ;
        RECT 173.510 370.190 173.720 370.400 ;
        RECT 224.660 371.420 224.830 371.590 ;
        RECT 248.950 371.960 249.120 372.130 ;
        RECT 250.500 372.110 250.670 372.280 ;
        RECT 248.950 371.510 249.120 371.680 ;
        RECT 217.400 371.010 217.570 371.180 ;
        RECT 244.210 371.010 244.380 371.180 ;
        RECT 252.790 372.110 252.960 372.280 ;
        RECT 254.490 372.130 254.660 372.300 ;
        RECT 250.140 371.270 250.320 371.460 ;
        RECT 252.740 371.460 252.910 371.630 ;
        RECT 253.730 371.720 253.900 371.890 ;
        RECT 253.800 371.100 253.970 371.270 ;
        RECT 172.040 369.820 172.210 369.990 ;
        RECT 252.740 370.200 252.910 370.370 ;
        RECT 174.470 369.720 174.640 369.890 ;
        RECT 175.510 369.760 175.680 369.930 ;
        RECT 176.550 369.420 176.720 369.590 ;
        RECT 223.850 369.480 224.020 369.650 ;
        RECT 237.760 369.480 237.930 369.650 ;
        RECT 248.250 369.650 248.420 369.820 ;
        RECT 253.730 369.940 253.900 370.110 ;
        RECT 176.550 369.060 176.720 369.230 ;
        RECT 147.370 368.650 147.540 368.820 ;
        RECT 148.460 368.660 148.630 368.830 ;
        RECT 173.510 368.440 173.720 368.650 ;
        RECT 172.040 368.070 172.210 368.240 ;
        RECT 174.470 367.970 174.640 368.140 ;
        RECT 198.440 368.210 198.700 369.030 ;
        RECT 210.390 368.240 210.710 369.030 ;
        RECT 240.300 369.350 240.470 369.520 ;
        RECT 211.840 368.670 212.020 368.860 ;
        RECT 145.830 367.740 146.000 367.910 ;
        RECT 147.380 367.660 147.550 367.830 ;
        RECT 148.160 367.610 148.330 367.780 ;
        RECT 148.470 367.670 148.640 367.840 ;
        RECT 175.510 368.010 175.680 368.180 ;
        RECT 176.550 367.670 176.720 367.840 ;
        RECT 211.460 367.630 211.640 367.820 ;
        RECT 176.550 367.310 176.720 367.480 ;
        RECT 145.810 366.820 145.980 366.990 ;
        RECT 239.360 368.670 239.530 368.840 ;
        RECT 239.840 368.730 240.010 368.900 ;
        RECT 246.750 369.080 246.920 369.250 ;
        RECT 252.790 369.550 252.960 369.720 ;
        RECT 254.410 369.880 254.580 370.050 ;
        RECT 241.030 368.670 241.200 368.840 ;
        RECT 241.950 368.740 242.120 368.910 ;
        RECT 248.410 369.040 248.580 369.210 ;
        RECT 217.400 368.250 217.570 368.420 ;
        RECT 244.210 368.250 244.380 368.420 ;
        RECT 246.700 368.430 246.870 368.600 ;
        RECT 247.690 368.690 247.860 368.860 ;
        RECT 248.400 368.820 248.570 368.990 ;
        RECT 224.690 367.730 224.860 367.900 ;
        RECT 247.560 368.000 247.730 368.170 ;
        RECT 212.660 367.310 212.830 367.480 ;
        RECT 239.370 367.540 239.540 367.710 ;
        RECT 247.760 367.660 247.930 367.830 ;
        RECT 147.380 366.670 147.550 366.840 ;
        RECT 148.470 366.680 148.640 366.850 ;
        RECT 173.510 366.690 173.720 366.900 ;
        RECT 211.110 366.810 211.280 366.980 ;
        RECT 212.660 366.860 212.830 367.030 ;
        RECT 172.040 366.320 172.210 366.490 ;
        RECT 174.470 366.220 174.640 366.390 ;
        RECT 212.920 366.510 213.100 366.680 ;
        RECT 246.700 367.170 246.870 367.340 ;
        RECT 247.690 366.910 247.860 367.080 ;
        RECT 248.950 367.310 249.120 367.480 ;
        RECT 250.140 367.630 250.320 367.820 ;
        RECT 246.750 366.520 246.920 366.690 ;
        RECT 145.790 365.830 145.960 366.000 ;
        RECT 147.290 365.940 147.460 366.110 ;
        RECT 148.590 365.840 148.760 366.010 ;
        RECT 175.510 366.260 175.680 366.430 ;
        RECT 248.460 366.890 248.630 366.990 ;
        RECT 248.290 366.820 248.630 366.890 ;
        RECT 248.950 366.860 249.120 367.030 ;
        RECT 248.290 366.720 248.460 366.820 ;
        RECT 250.500 366.810 250.670 366.980 ;
        RECT 176.550 365.920 176.720 366.090 ;
        RECT 240.300 366.150 240.470 366.320 ;
        RECT 246.750 366.080 246.920 366.250 ;
        RECT 176.550 365.560 176.720 365.730 ;
        RECT 227.910 365.470 228.080 365.640 ;
        RECT 147.290 364.950 147.460 365.120 ;
        RECT 148.590 364.850 148.760 365.020 ;
        RECT 227.920 364.750 228.090 364.920 ;
        RECT 233.700 365.470 233.870 365.640 ;
        RECT 239.360 365.470 239.530 365.640 ;
        RECT 239.840 365.530 240.010 365.700 ;
        RECT 248.450 366.100 248.620 366.270 ;
        RECT 248.680 365.990 248.850 366.160 ;
        RECT 241.030 365.470 241.200 365.640 ;
        RECT 241.950 365.540 242.120 365.710 ;
        RECT 246.700 365.430 246.870 365.600 ;
        RECT 247.690 365.690 247.860 365.860 ;
        RECT 233.700 364.750 233.870 364.920 ;
        RECT 247.760 365.070 247.930 365.240 ;
        RECT 238.860 364.530 239.030 364.720 ;
        RECT 239.370 364.740 239.540 364.910 ;
        RECT 239.370 364.340 239.540 364.510 ;
        RECT 147.290 363.960 147.460 364.130 ;
        RECT 246.700 364.170 246.870 364.340 ;
        RECT 147.730 363.510 147.900 363.680 ;
        RECT 148.590 363.860 148.760 364.030 ;
        RECT 247.690 363.910 247.860 364.080 ;
        RECT 239.360 363.610 239.530 363.780 ;
        RECT 239.840 363.550 240.010 363.720 ;
        RECT 241.030 363.610 241.200 363.780 ;
        RECT 241.950 363.540 242.120 363.710 ;
        RECT 242.210 363.620 242.380 363.790 ;
        RECT 246.750 363.520 246.920 363.690 ;
        RECT 248.370 363.850 248.540 364.020 ;
        RECT 240.300 362.930 240.470 363.100 ;
        RECT 186.410 362.690 186.580 362.860 ;
        RECT 187.250 362.570 187.420 362.740 ;
        RECT 188.000 362.570 188.170 362.740 ;
        RECT 186.280 362.050 186.450 362.220 ;
        RECT 190.980 362.240 191.150 362.410 ;
        RECT 186.590 361.860 186.760 362.030 ;
        RECT 191.380 362.690 191.550 362.860 ;
        RECT 242.360 362.790 242.530 362.960 ;
        RECT 191.380 362.330 191.550 362.500 ;
        RECT 176.550 361.400 176.720 361.570 ;
        RECT 190.980 361.480 191.150 361.650 ;
        RECT 176.550 361.040 176.720 361.210 ;
        RECT 187.250 361.150 187.420 361.320 ;
        RECT 188.000 361.150 188.170 361.320 ;
        RECT 190.000 361.160 190.170 361.330 ;
        RECT 191.380 361.750 191.550 361.920 ;
        RECT 241.520 361.970 241.690 362.140 ;
        RECT 191.380 361.390 191.550 361.560 ;
        RECT 239.370 361.540 239.540 361.710 ;
        RECT 238.860 361.330 239.030 361.500 ;
        RECT 172.040 360.640 172.210 360.810 ;
        RECT 174.470 360.740 174.640 360.910 ;
        RECT 175.510 360.700 175.680 360.870 ;
        RECT 173.510 360.230 173.720 360.440 ;
        RECT 239.360 360.410 239.530 360.580 ;
        RECT 239.840 360.350 240.010 360.520 ;
        RECT 242.250 360.690 242.420 360.860 ;
        RECT 241.030 360.410 241.200 360.580 ;
        RECT 241.950 360.340 242.120 360.510 ;
        RECT 176.550 359.650 176.720 359.820 ;
        RECT 240.300 359.730 240.470 359.900 ;
        RECT 242.640 359.960 242.810 360.130 ;
        RECT 176.550 359.290 176.720 359.460 ;
        RECT 186.410 359.490 186.580 359.660 ;
        RECT 187.250 359.370 187.420 359.540 ;
        RECT 188.000 359.370 188.170 359.540 ;
        RECT 172.040 358.890 172.210 359.060 ;
        RECT 174.470 358.990 174.640 359.160 ;
        RECT 175.510 358.950 175.680 359.120 ;
        RECT 186.280 358.850 186.450 359.020 ;
        RECT 190.980 359.040 191.150 359.210 ;
        RECT 173.510 358.480 173.720 358.690 ;
        RECT 186.590 358.660 186.760 358.830 ;
        RECT 191.380 359.490 191.550 359.660 ;
        RECT 191.380 359.130 191.550 359.300 ;
        RECT 190.980 358.280 191.150 358.450 ;
        RECT 22.730 351.730 22.900 351.900 ;
        RECT 23.090 351.730 23.260 351.900 ;
        RECT 23.460 351.730 23.630 351.900 ;
        RECT 24.250 346.450 24.420 346.460 ;
        RECT 24.240 344.590 24.420 346.450 ;
        RECT 25.380 346.220 25.550 357.200 ;
        RECT 26.000 346.220 26.170 357.200 ;
        RECT 26.620 346.230 26.790 357.210 ;
        RECT 27.200 346.250 27.370 357.230 ;
        RECT 27.790 346.260 27.960 357.240 ;
        RECT 28.390 346.260 28.560 357.240 ;
        RECT 28.990 346.210 29.160 357.190 ;
        RECT 29.600 346.220 29.770 357.200 ;
        RECT 30.200 346.210 30.370 357.190 ;
        RECT 176.550 357.900 176.720 358.070 ;
        RECT 187.250 357.950 187.420 358.120 ;
        RECT 188.000 357.950 188.170 358.120 ;
        RECT 190.000 357.960 190.170 358.130 ;
        RECT 191.380 358.550 191.550 358.720 ;
        RECT 196.770 358.610 197.040 358.880 ;
        RECT 200.800 358.680 201.070 358.950 ;
        RECT 236.110 358.680 236.380 358.950 ;
        RECT 240.140 358.610 240.410 358.880 ;
        RECT 191.380 358.190 191.550 358.360 ;
        RECT 176.550 357.540 176.720 357.710 ;
        RECT 172.040 357.140 172.210 357.310 ;
        RECT 174.470 357.240 174.640 357.410 ;
        RECT 175.510 357.200 175.680 357.370 ;
        RECT 205.100 357.550 205.270 357.720 ;
        RECT 231.910 357.550 232.080 357.720 ;
        RECT 203.430 357.140 203.600 357.310 ;
        RECT 173.510 356.730 173.720 356.940 ;
        RECT 204.160 357.110 204.330 357.280 ;
        RECT 205.100 357.000 205.270 357.170 ;
        RECT 231.910 357.000 232.080 357.170 ;
        RECT 232.850 357.110 233.020 357.280 ;
        RECT 233.580 357.140 233.750 357.310 ;
        RECT 176.550 356.150 176.720 356.320 ;
        RECT 176.550 355.790 176.720 355.960 ;
        RECT 209.040 356.040 209.210 356.210 ;
        RECT 172.040 355.390 172.210 355.560 ;
        RECT 174.470 355.490 174.640 355.660 ;
        RECT 175.510 355.450 175.680 355.620 ;
        RECT 212.980 356.050 213.150 356.220 ;
        RECT 224.030 356.050 224.200 356.220 ;
        RECT 227.970 356.040 228.140 356.210 ;
        RECT 173.510 354.980 173.720 355.190 ;
        RECT 203.430 354.760 203.600 354.930 ;
        RECT 204.160 354.790 204.330 354.960 ;
        RECT 205.100 354.900 205.270 355.070 ;
        RECT 205.100 354.310 205.270 354.520 ;
        RECT 209.040 354.450 209.210 354.620 ;
        RECT 209.040 354.090 209.210 354.260 ;
        RECT 203.430 353.900 203.600 354.070 ;
        RECT 204.160 353.870 204.330 354.040 ;
        RECT 205.100 353.760 205.270 353.930 ;
        RECT 212.970 354.590 213.140 354.760 ;
        RECT 212.970 354.230 213.140 354.400 ;
        RECT 231.910 354.900 232.080 355.070 ;
        RECT 224.040 354.590 224.210 354.760 ;
        RECT 224.040 354.230 224.210 354.400 ;
        RECT 232.850 354.790 233.020 354.960 ;
        RECT 233.580 354.760 233.750 354.930 ;
        RECT 227.970 354.450 228.140 354.620 ;
        RECT 230.330 354.330 230.510 354.500 ;
        RECT 231.910 354.310 232.080 354.520 ;
        RECT 227.970 354.090 228.140 354.260 ;
        RECT 231.910 353.760 232.080 353.930 ;
        RECT 232.850 353.870 233.020 354.040 ;
        RECT 233.580 353.900 233.750 354.070 ;
        RECT 186.390 352.220 186.560 352.390 ;
        RECT 187.230 352.100 187.400 352.270 ;
        RECT 187.980 352.100 188.150 352.270 ;
        RECT 186.260 351.580 186.430 351.750 ;
        RECT 190.960 351.770 191.130 351.940 ;
        RECT 176.550 351.270 176.720 351.440 ;
        RECT 186.570 351.390 186.740 351.560 ;
        RECT 191.360 352.220 191.530 352.390 ;
        RECT 191.360 351.860 191.530 352.030 ;
        RECT 203.430 351.530 203.600 351.700 ;
        RECT 204.160 351.560 204.330 351.730 ;
        RECT 205.100 351.670 205.270 351.840 ;
        RECT 231.910 351.670 232.080 351.840 ;
        RECT 232.850 351.560 233.020 351.730 ;
        RECT 233.580 351.530 233.750 351.700 ;
        RECT 176.550 350.910 176.720 351.080 ;
        RECT 190.960 351.010 191.130 351.180 ;
        RECT 172.040 350.510 172.210 350.680 ;
        RECT 174.470 350.610 174.640 350.780 ;
        RECT 175.510 350.570 175.680 350.740 ;
        RECT 187.230 350.680 187.400 350.850 ;
        RECT 187.980 350.680 188.150 350.850 ;
        RECT 189.980 350.690 190.150 350.860 ;
        RECT 191.360 351.280 191.530 351.450 ;
        RECT 205.100 351.120 205.270 351.290 ;
        RECT 191.360 350.920 191.530 351.090 ;
        RECT 231.910 351.120 232.080 351.290 ;
        RECT 173.510 350.100 173.720 350.310 ;
        RECT 197.370 349.730 197.640 350.000 ;
        RECT 176.550 349.520 176.720 349.690 ;
        RECT 201.400 349.800 201.670 350.070 ;
        RECT 176.550 349.160 176.720 349.330 ;
        RECT 172.040 348.760 172.210 348.930 ;
        RECT 174.470 348.860 174.640 349.030 ;
        RECT 175.510 348.820 175.680 348.990 ;
        RECT 186.390 349.020 186.560 349.190 ;
        RECT 187.230 348.900 187.400 349.070 ;
        RECT 187.980 348.900 188.150 349.070 ;
        RECT 173.510 348.350 173.720 348.560 ;
        RECT 186.260 348.380 186.430 348.550 ;
        RECT 190.960 348.570 191.130 348.740 ;
        RECT 186.570 348.190 186.740 348.360 ;
        RECT 176.550 347.770 176.720 347.940 ;
        RECT 191.360 349.020 191.530 349.190 ;
        RECT 191.360 348.660 191.530 348.830 ;
        RECT 205.700 348.710 205.870 348.880 ;
        RECT 204.030 348.300 204.200 348.470 ;
        RECT 190.960 347.810 191.130 347.980 ;
        RECT 176.550 347.410 176.720 347.580 ;
        RECT 187.230 347.480 187.400 347.650 ;
        RECT 187.980 347.480 188.150 347.650 ;
        RECT 189.980 347.490 190.150 347.660 ;
        RECT 191.360 348.080 191.530 348.250 ;
        RECT 191.360 347.720 191.530 347.890 ;
        RECT 204.760 348.270 204.930 348.440 ;
        RECT 205.700 348.160 205.870 348.330 ;
        RECT 172.040 347.010 172.210 347.180 ;
        RECT 174.470 347.110 174.640 347.280 ;
        RECT 175.510 347.070 175.680 347.240 ;
        RECT 209.770 347.140 209.940 347.310 ;
        RECT 173.510 346.600 173.720 346.810 ;
        RECT 213.790 347.170 213.960 347.340 ;
        RECT 176.550 346.020 176.720 346.190 ;
        RECT 24.610 345.030 26.520 345.210 ;
        RECT 204.030 345.940 204.200 346.110 ;
        RECT 204.760 345.970 204.930 346.140 ;
        RECT 205.700 346.080 205.870 346.250 ;
        RECT 209.760 345.940 209.930 346.110 ;
        RECT 176.550 345.660 176.720 345.830 ;
        RECT 172.040 345.260 172.210 345.430 ;
        RECT 174.470 345.360 174.640 345.530 ;
        RECT 175.510 345.320 175.680 345.490 ;
        RECT 205.700 345.470 205.870 345.700 ;
        RECT 173.510 344.850 173.720 345.060 ;
        RECT 209.760 345.280 209.930 345.450 ;
        RECT 204.030 345.060 204.200 345.230 ;
        RECT 24.610 344.630 26.510 344.810 ;
        RECT 204.760 345.030 204.930 345.200 ;
        RECT 205.700 344.920 205.870 345.090 ;
        RECT 213.780 345.880 213.950 346.050 ;
        RECT 213.780 345.240 213.950 345.410 ;
        RECT 24.480 342.930 25.410 343.130 ;
        RECT 186.420 342.950 186.590 343.120 ;
        RECT 24.250 339.360 24.430 342.520 ;
        RECT 27.350 341.860 30.650 342.210 ;
        RECT 22.410 329.820 22.580 329.990 ;
        RECT 22.770 329.820 22.940 329.990 ;
        RECT 23.130 329.820 23.300 329.990 ;
        RECT 23.490 329.820 23.660 329.990 ;
        RECT 26.140 331.360 26.310 340.810 ;
        RECT 26.890 331.350 27.060 340.740 ;
        RECT 27.610 331.380 27.780 340.780 ;
        RECT 28.270 331.390 28.440 340.760 ;
        RECT 28.920 331.380 29.090 340.830 ;
        RECT 29.560 331.390 29.730 340.780 ;
        RECT 151.780 342.680 151.950 342.850 ;
        RECT 152.430 342.680 152.600 342.850 ;
        RECT 187.260 342.830 187.430 343.000 ;
        RECT 188.010 342.830 188.180 343.000 ;
        RECT 150.560 342.240 150.730 342.410 ;
        RECT 151.260 342.240 151.430 342.410 ;
        RECT 149.880 340.470 150.050 340.640 ;
        RECT 176.510 342.210 176.680 342.380 ;
        RECT 186.290 342.310 186.460 342.480 ;
        RECT 190.990 342.500 191.160 342.670 ;
        RECT 152.800 342.010 152.970 342.180 ;
        RECT 176.510 341.850 176.680 342.020 ;
        RECT 186.600 342.120 186.770 342.290 ;
        RECT 191.390 342.950 191.560 343.120 ;
        RECT 191.390 342.590 191.560 342.760 ;
        RECT 204.030 342.690 204.200 342.860 ;
        RECT 221.630 343.070 221.800 343.240 ;
        RECT 204.760 342.720 204.930 342.890 ;
        RECT 205.700 342.830 205.870 343.000 ;
        RECT 220.880 342.770 221.050 342.940 ;
        RECT 220.730 342.530 220.900 342.700 ;
        RECT 205.700 342.280 205.870 342.450 ;
        RECT 222.890 342.500 223.060 342.670 ;
        RECT 172.000 341.450 172.170 341.620 ;
        RECT 174.430 341.550 174.600 341.720 ;
        RECT 175.470 341.510 175.640 341.680 ;
        RECT 190.990 341.740 191.160 341.910 ;
        RECT 187.260 341.410 187.430 341.580 ;
        RECT 188.010 341.410 188.180 341.580 ;
        RECT 190.010 341.420 190.180 341.590 ;
        RECT 191.390 342.010 191.560 342.180 ;
        RECT 220.730 342.090 220.900 342.260 ;
        RECT 222.890 342.120 223.060 342.290 ;
        RECT 191.390 341.650 191.560 341.820 ;
        RECT 220.880 341.850 221.050 342.020 ;
        RECT 221.630 341.550 221.800 341.720 ;
        RECT 173.470 341.040 173.680 341.250 ;
        RECT 152.710 340.440 152.880 340.610 ;
        RECT 176.510 340.460 176.680 340.630 ;
        RECT 152.720 339.900 152.890 340.070 ;
        RECT 176.510 340.100 176.680 340.270 ;
        RECT 221.630 340.300 221.800 340.470 ;
        RECT 147.480 337.890 147.650 338.060 ;
        RECT 144.170 337.450 144.340 337.620 ;
        RECT 145.270 337.460 145.440 337.630 ;
        RECT 146.360 337.460 146.530 337.630 ;
        RECT 147.490 337.420 147.660 337.590 ;
        RECT 144.720 336.780 144.890 336.950 ;
        RECT 144.720 335.410 144.890 335.580 ;
        RECT 172.000 339.700 172.170 339.870 ;
        RECT 174.430 339.800 174.600 339.970 ;
        RECT 175.470 339.760 175.640 339.930 ;
        RECT 220.880 340.000 221.050 340.170 ;
        RECT 186.420 339.750 186.590 339.920 ;
        RECT 173.470 339.290 173.680 339.500 ;
        RECT 187.260 339.630 187.430 339.800 ;
        RECT 188.010 339.630 188.180 339.800 ;
        RECT 152.790 339.030 152.960 339.200 ;
        RECT 186.290 339.110 186.460 339.280 ;
        RECT 190.990 339.300 191.160 339.470 ;
        RECT 176.510 338.710 176.680 338.880 ;
        RECT 186.600 338.920 186.770 339.090 ;
        RECT 150.590 338.360 150.760 338.530 ;
        RECT 151.280 338.350 151.450 338.520 ;
        RECT 191.390 339.750 191.560 339.920 ;
        RECT 220.730 339.760 220.900 339.930 ;
        RECT 191.390 339.390 191.560 339.560 ;
        RECT 222.890 339.730 223.060 339.900 ;
        RECT 208.750 339.190 208.920 339.360 ;
        RECT 220.730 339.320 220.900 339.490 ;
        RECT 222.890 339.350 223.060 339.520 ;
        RECT 176.510 338.350 176.680 338.520 ;
        RECT 190.990 338.540 191.160 338.710 ;
        RECT 172.000 337.950 172.170 338.120 ;
        RECT 174.430 338.050 174.600 338.220 ;
        RECT 175.470 338.010 175.640 338.180 ;
        RECT 187.260 338.210 187.430 338.380 ;
        RECT 188.010 338.210 188.180 338.380 ;
        RECT 190.010 338.220 190.180 338.390 ;
        RECT 191.390 338.810 191.560 338.980 ;
        RECT 191.390 338.450 191.560 338.620 ;
        RECT 220.880 339.080 221.050 339.250 ;
        RECT 221.630 338.780 221.800 338.950 ;
        RECT 208.800 338.230 208.970 338.400 ;
        RECT 151.760 337.580 151.930 337.750 ;
        RECT 152.470 337.520 152.640 337.690 ;
        RECT 173.470 337.540 173.680 337.750 ;
        RECT 145.820 336.780 145.990 336.950 ;
        RECT 146.920 336.780 147.090 336.950 ;
        RECT 147.750 336.910 147.920 337.080 ;
        RECT 176.510 336.960 176.680 337.130 ;
        RECT 176.510 336.600 176.680 336.770 ;
        RECT 147.750 336.220 147.920 336.390 ;
        RECT 172.000 336.200 172.170 336.370 ;
        RECT 174.430 336.300 174.600 336.470 ;
        RECT 175.470 336.260 175.640 336.430 ;
        RECT 173.470 335.790 173.680 336.000 ;
        RECT 145.820 335.410 145.990 335.580 ;
        RECT 146.920 335.410 147.090 335.580 ;
        RECT 144.170 334.680 144.340 334.850 ;
        RECT 144.160 333.340 144.330 333.510 ;
        RECT 145.270 334.680 145.440 334.850 ;
        RECT 146.360 334.680 146.530 334.850 ;
        RECT 154.300 333.660 154.470 334.000 ;
        RECT 154.670 333.660 154.840 334.000 ;
        RECT 145.270 333.330 145.440 333.500 ;
        RECT 146.360 333.310 146.530 333.480 ;
        RECT 144.720 332.640 144.890 332.810 ;
        RECT 145.820 332.630 145.990 332.800 ;
        RECT 146.910 332.630 147.080 332.800 ;
        RECT 177.400 331.470 177.570 331.640 ;
        RECT 147.520 330.330 147.690 330.500 ;
        RECT 144.210 329.890 144.380 330.060 ;
        RECT 22.730 323.140 22.900 323.310 ;
        RECT 23.090 323.140 23.260 323.310 ;
        RECT 23.460 323.140 23.630 323.310 ;
        RECT 24.250 317.860 24.420 317.870 ;
        RECT 24.240 316.000 24.420 317.860 ;
        RECT 25.380 317.630 25.550 328.610 ;
        RECT 26.000 317.630 26.170 328.610 ;
        RECT 26.620 317.640 26.790 328.620 ;
        RECT 27.200 317.660 27.370 328.640 ;
        RECT 27.790 317.670 27.960 328.650 ;
        RECT 28.390 317.670 28.560 328.650 ;
        RECT 28.990 317.620 29.160 328.600 ;
        RECT 29.600 317.630 29.770 328.610 ;
        RECT 30.200 317.620 30.370 328.600 ;
        RECT 145.310 329.900 145.480 330.070 ;
        RECT 144.760 329.220 144.930 329.390 ;
        RECT 144.760 327.850 144.930 328.020 ;
        RECT 146.400 329.900 146.570 330.070 ;
        RECT 145.860 329.220 146.030 329.390 ;
        RECT 145.860 327.850 146.030 328.020 ;
        RECT 147.530 329.860 147.700 330.030 ;
        RECT 146.960 329.220 147.130 329.390 ;
        RECT 178.490 331.470 178.660 331.640 ;
        RECT 177.950 330.790 178.120 330.960 ;
        RECT 177.950 329.420 178.120 329.590 ;
        RECT 179.590 331.460 179.760 331.630 ;
        RECT 179.040 330.770 179.210 330.940 ;
        RECT 179.040 329.420 179.210 329.590 ;
        RECT 180.570 331.490 180.740 331.660 ;
        RECT 180.570 331.130 180.740 331.300 ;
        RECT 180.150 330.760 180.320 330.930 ;
        RECT 182.460 331.490 182.630 331.660 ;
        RECT 182.460 331.130 182.630 331.300 ;
        RECT 183.440 331.460 183.610 331.630 ;
        RECT 182.880 330.760 183.050 330.930 ;
        RECT 180.140 329.420 180.310 329.590 ;
        RECT 182.890 329.420 183.060 329.590 ;
        RECT 184.540 331.470 184.710 331.640 ;
        RECT 183.990 330.770 184.160 330.940 ;
        RECT 183.990 329.420 184.160 329.590 ;
        RECT 185.630 331.470 185.800 331.640 ;
        RECT 185.080 330.790 185.250 330.960 ;
        RECT 185.080 329.420 185.250 329.590 ;
        RECT 187.210 331.500 187.380 331.670 ;
        RECT 188.300 331.500 188.470 331.670 ;
        RECT 187.760 330.820 187.930 330.990 ;
        RECT 187.760 329.450 187.930 329.620 ;
        RECT 189.400 331.490 189.570 331.660 ;
        RECT 188.850 330.800 189.020 330.970 ;
        RECT 188.850 329.450 189.020 329.620 ;
        RECT 190.380 331.520 190.550 331.690 ;
        RECT 190.380 331.160 190.550 331.330 ;
        RECT 189.960 330.790 190.130 330.960 ;
        RECT 192.270 331.520 192.440 331.690 ;
        RECT 192.270 331.160 192.440 331.330 ;
        RECT 193.250 331.490 193.420 331.660 ;
        RECT 192.690 330.790 192.860 330.960 ;
        RECT 189.950 329.450 190.120 329.620 ;
        RECT 192.700 329.450 192.870 329.620 ;
        RECT 194.350 331.500 194.520 331.670 ;
        RECT 193.800 330.800 193.970 330.970 ;
        RECT 193.800 329.450 193.970 329.620 ;
        RECT 195.440 331.500 195.610 331.670 ;
        RECT 194.890 330.820 195.060 330.990 ;
        RECT 194.890 329.450 195.060 329.620 ;
        RECT 198.990 331.470 199.160 331.640 ;
        RECT 198.430 330.770 198.600 330.940 ;
        RECT 198.440 329.430 198.610 329.600 ;
        RECT 200.090 331.480 200.260 331.650 ;
        RECT 201.180 331.480 201.350 331.650 ;
        RECT 199.540 330.780 199.710 330.950 ;
        RECT 200.630 330.800 200.800 330.970 ;
        RECT 199.540 329.430 199.710 329.600 ;
        RECT 200.630 329.430 200.800 329.600 ;
        RECT 177.390 328.690 177.560 328.860 ;
        RECT 146.960 327.850 147.130 328.020 ;
        RECT 144.210 327.120 144.380 327.290 ;
        RECT 144.200 325.780 144.370 325.950 ;
        RECT 143.780 325.410 143.950 325.580 ;
        RECT 145.310 327.120 145.480 327.290 ;
        RECT 145.310 325.770 145.480 325.940 ;
        RECT 144.760 325.080 144.930 325.250 ;
        RECT 146.400 327.120 146.570 327.290 ;
        RECT 146.400 325.750 146.570 325.920 ;
        RECT 145.860 325.070 146.030 325.240 ;
        RECT 177.390 327.320 177.560 327.490 ;
        RECT 176.820 326.680 176.990 326.850 ;
        RECT 178.490 328.690 178.660 328.860 ;
        RECT 178.490 327.320 178.660 327.490 ;
        RECT 177.950 326.640 178.120 326.810 ;
        RECT 179.590 328.690 179.760 328.860 ;
        RECT 179.590 327.320 179.760 327.490 ;
        RECT 179.040 326.640 179.210 326.810 ;
        RECT 183.440 328.690 183.610 328.860 ;
        RECT 183.440 327.320 183.610 327.490 ;
        RECT 180.140 326.650 180.310 326.820 ;
        RECT 182.890 326.650 183.060 326.820 ;
        RECT 184.540 328.690 184.710 328.860 ;
        RECT 184.540 327.320 184.710 327.490 ;
        RECT 183.990 326.640 184.160 326.810 ;
        RECT 185.640 328.690 185.810 328.860 ;
        RECT 187.200 328.720 187.370 328.890 ;
        RECT 185.640 327.320 185.810 327.490 ;
        RECT 187.200 327.350 187.370 327.520 ;
        RECT 185.080 326.640 185.250 326.810 ;
        RECT 186.210 326.680 186.380 326.850 ;
        RECT 186.630 326.710 186.800 326.880 ;
        RECT 188.300 328.720 188.470 328.890 ;
        RECT 188.300 327.350 188.470 327.520 ;
        RECT 187.760 326.670 187.930 326.840 ;
        RECT 189.400 328.720 189.570 328.890 ;
        RECT 189.400 327.350 189.570 327.520 ;
        RECT 188.850 326.670 189.020 326.840 ;
        RECT 193.250 328.720 193.420 328.890 ;
        RECT 193.250 327.350 193.420 327.520 ;
        RECT 189.950 326.680 190.120 326.850 ;
        RECT 192.700 326.680 192.870 326.850 ;
        RECT 194.350 328.720 194.520 328.890 ;
        RECT 194.350 327.350 194.520 327.520 ;
        RECT 193.800 326.670 193.970 326.840 ;
        RECT 195.450 328.720 195.620 328.890 ;
        RECT 195.450 327.350 195.620 327.520 ;
        RECT 194.890 326.670 195.060 326.840 ;
        RECT 196.020 326.710 196.190 326.880 ;
        RECT 198.990 328.700 199.160 328.870 ;
        RECT 198.990 327.330 199.160 327.500 ;
        RECT 198.440 326.660 198.610 326.830 ;
        RECT 200.090 328.700 200.260 328.870 ;
        RECT 201.190 328.700 201.360 328.870 ;
        RECT 202.020 328.250 202.190 328.420 ;
        RECT 202.020 327.890 202.190 328.060 ;
        RECT 200.090 327.330 200.260 327.500 ;
        RECT 201.190 327.330 201.360 327.500 ;
        RECT 199.540 326.650 199.710 326.820 ;
        RECT 200.630 326.650 200.800 326.820 ;
        RECT 201.760 326.690 201.930 326.860 ;
        RECT 176.830 326.210 177.000 326.380 ;
        RECT 186.200 326.210 186.370 326.380 ;
        RECT 186.640 326.240 186.810 326.410 ;
        RECT 196.010 326.240 196.180 326.410 ;
        RECT 201.750 326.220 201.920 326.390 ;
        RECT 146.950 325.070 147.120 325.240 ;
        RECT 148.490 321.690 148.660 325.210 ;
        RECT 148.850 321.690 149.020 325.210 ;
        RECT 149.210 321.690 149.380 325.210 ;
        RECT 149.900 321.690 150.070 325.210 ;
        RECT 150.260 321.690 150.430 325.210 ;
        RECT 150.620 321.690 150.790 325.210 ;
        RECT 227.330 324.020 227.500 324.190 ;
        RECT 232.920 323.320 233.090 323.490 ;
        RECT 232.920 322.650 233.090 322.820 ;
        RECT 227.330 322.410 227.500 322.580 ;
        RECT 227.330 320.810 227.500 320.980 ;
        RECT 227.330 319.190 227.500 319.360 ;
        RECT 232.340 317.980 232.510 318.150 ;
        RECT 227.330 317.590 227.500 317.760 ;
        RECT 24.610 316.440 26.520 316.620 ;
        RECT 24.610 316.040 26.510 316.220 ;
        RECT 227.330 315.970 227.500 316.140 ;
        RECT 24.480 314.340 25.410 314.540 ;
        RECT 227.330 314.370 227.500 314.540 ;
        RECT 238.860 314.480 239.030 329.430 ;
        RECT 24.250 310.770 24.430 313.930 ;
        RECT 27.350 313.270 30.650 313.620 ;
        RECT 22.410 301.230 22.580 301.400 ;
        RECT 22.770 301.230 22.940 301.400 ;
        RECT 23.130 301.230 23.300 301.400 ;
        RECT 23.490 301.230 23.660 301.400 ;
        RECT 26.140 302.770 26.310 312.220 ;
        RECT 26.890 302.760 27.060 312.150 ;
        RECT 27.610 302.790 27.780 312.190 ;
        RECT 28.270 302.800 28.440 312.170 ;
        RECT 28.920 302.790 29.090 312.240 ;
        RECT 29.560 302.800 29.730 312.190 ;
        RECT 227.330 312.750 227.500 312.920 ;
        RECT 22.730 294.550 22.900 294.720 ;
        RECT 23.090 294.550 23.260 294.720 ;
        RECT 23.460 294.550 23.630 294.720 ;
        RECT 24.250 289.270 24.420 289.280 ;
        RECT 24.240 287.410 24.420 289.270 ;
        RECT 25.380 289.040 25.550 300.020 ;
        RECT 26.000 289.040 26.170 300.020 ;
        RECT 26.620 289.050 26.790 300.030 ;
        RECT 27.200 289.070 27.370 300.050 ;
        RECT 27.790 289.080 27.960 300.060 ;
        RECT 28.390 289.080 28.560 300.060 ;
        RECT 28.990 289.030 29.160 300.010 ;
        RECT 29.600 289.040 29.770 300.020 ;
        RECT 30.200 289.030 30.370 300.010 ;
        RECT 24.610 287.850 26.520 288.030 ;
        RECT 24.610 287.450 26.510 287.630 ;
        RECT 24.480 285.750 25.410 285.950 ;
        RECT 24.250 282.180 24.430 285.340 ;
        RECT 27.350 284.680 30.650 285.030 ;
        RECT 22.410 272.640 22.580 272.810 ;
        RECT 22.770 272.640 22.940 272.810 ;
        RECT 23.130 272.640 23.300 272.810 ;
        RECT 23.490 272.640 23.660 272.810 ;
        RECT 26.140 274.180 26.310 283.630 ;
        RECT 26.890 274.170 27.060 283.560 ;
        RECT 27.610 274.200 27.780 283.600 ;
        RECT 28.270 274.210 28.440 283.580 ;
        RECT 28.920 274.200 29.090 283.650 ;
        RECT 29.560 274.210 29.730 283.600 ;
        RECT 22.730 265.960 22.900 266.130 ;
        RECT 23.090 265.960 23.260 266.130 ;
        RECT 23.460 265.960 23.630 266.130 ;
        RECT 24.250 260.680 24.420 260.690 ;
        RECT 24.240 258.820 24.420 260.680 ;
        RECT 25.380 260.450 25.550 271.430 ;
        RECT 26.000 260.450 26.170 271.430 ;
        RECT 26.620 260.460 26.790 271.440 ;
        RECT 27.200 260.480 27.370 271.460 ;
        RECT 27.790 260.490 27.960 271.470 ;
        RECT 28.390 260.490 28.560 271.470 ;
        RECT 28.990 260.440 29.160 271.420 ;
        RECT 29.600 260.450 29.770 271.430 ;
        RECT 30.200 260.440 30.370 271.420 ;
        RECT 390.210 285.030 391.140 285.230 ;
        RECT 384.970 283.960 388.270 284.310 ;
        RECT 385.890 273.490 386.060 282.880 ;
        RECT 386.530 273.480 386.700 282.930 ;
        RECT 387.180 273.490 387.350 282.860 ;
        RECT 387.840 273.480 388.010 282.880 ;
        RECT 388.560 273.450 388.730 282.840 ;
        RECT 389.310 273.460 389.480 282.910 ;
        RECT 391.190 281.460 391.370 284.620 ;
        RECT 391.960 271.920 392.130 272.090 ;
        RECT 392.320 271.920 392.490 272.090 ;
        RECT 392.680 271.920 392.850 272.090 ;
        RECT 393.040 271.920 393.210 272.090 ;
        RECT 24.610 259.260 26.520 259.440 ;
        RECT 385.250 259.720 385.420 270.700 ;
        RECT 385.850 259.730 386.020 270.710 ;
        RECT 386.460 259.720 386.630 270.700 ;
        RECT 387.060 259.770 387.230 270.750 ;
        RECT 387.660 259.770 387.830 270.750 ;
        RECT 388.250 259.760 388.420 270.740 ;
        RECT 388.830 259.740 389.000 270.720 ;
        RECT 389.450 259.730 389.620 270.710 ;
        RECT 390.070 259.730 390.240 270.710 ;
        RECT 391.990 265.240 392.160 265.410 ;
        RECT 392.360 265.240 392.530 265.410 ;
        RECT 392.720 265.240 392.890 265.410 ;
        RECT 24.610 258.860 26.510 259.040 ;
        RECT 391.200 259.960 391.370 259.970 ;
        RECT 389.100 258.540 391.010 258.720 ;
        RECT 389.110 258.140 391.010 258.320 ;
        RECT 391.200 258.100 391.380 259.960 ;
        RECT 24.480 257.160 25.410 257.360 ;
        RECT 24.250 253.590 24.430 256.750 ;
        RECT 27.350 256.090 30.650 256.440 ;
        RECT 22.410 244.050 22.580 244.220 ;
        RECT 22.770 244.050 22.940 244.220 ;
        RECT 23.130 244.050 23.300 244.220 ;
        RECT 23.490 244.050 23.660 244.220 ;
        RECT 26.140 245.590 26.310 255.040 ;
        RECT 26.890 245.580 27.060 254.970 ;
        RECT 27.610 245.610 27.780 255.010 ;
        RECT 28.270 245.620 28.440 254.990 ;
        RECT 28.920 245.610 29.090 255.060 ;
        RECT 29.560 245.620 29.730 255.010 ;
        RECT 22.730 237.370 22.900 237.540 ;
        RECT 23.090 237.370 23.260 237.540 ;
        RECT 23.460 237.370 23.630 237.540 ;
        RECT 24.250 232.090 24.420 232.100 ;
        RECT 24.240 230.230 24.420 232.090 ;
        RECT 25.380 231.860 25.550 242.840 ;
        RECT 26.000 231.860 26.170 242.840 ;
        RECT 26.620 231.870 26.790 242.850 ;
        RECT 27.200 231.890 27.370 242.870 ;
        RECT 27.790 231.900 27.960 242.880 ;
        RECT 28.390 231.900 28.560 242.880 ;
        RECT 28.990 231.850 29.160 242.830 ;
        RECT 29.600 231.860 29.770 242.840 ;
        RECT 30.200 231.850 30.370 242.830 ;
        RECT 390.210 256.440 391.140 256.640 ;
        RECT 384.970 255.370 388.270 255.720 ;
        RECT 385.890 244.900 386.060 254.290 ;
        RECT 386.530 244.890 386.700 254.340 ;
        RECT 387.180 244.900 387.350 254.270 ;
        RECT 387.840 244.890 388.010 254.290 ;
        RECT 388.560 244.860 388.730 254.250 ;
        RECT 389.310 244.870 389.480 254.320 ;
        RECT 391.190 252.870 391.370 256.030 ;
        RECT 391.960 243.330 392.130 243.500 ;
        RECT 392.320 243.330 392.490 243.500 ;
        RECT 392.680 243.330 392.850 243.500 ;
        RECT 393.040 243.330 393.210 243.500 ;
        RECT 24.610 230.670 26.520 230.850 ;
        RECT 385.250 231.130 385.420 242.110 ;
        RECT 385.850 231.140 386.020 242.120 ;
        RECT 386.460 231.130 386.630 242.110 ;
        RECT 387.060 231.180 387.230 242.160 ;
        RECT 387.660 231.180 387.830 242.160 ;
        RECT 388.250 231.170 388.420 242.150 ;
        RECT 388.830 231.150 389.000 242.130 ;
        RECT 389.450 231.140 389.620 242.120 ;
        RECT 390.070 231.140 390.240 242.120 ;
        RECT 391.990 236.650 392.160 236.820 ;
        RECT 392.360 236.650 392.530 236.820 ;
        RECT 392.720 236.650 392.890 236.820 ;
        RECT 24.610 230.270 26.510 230.450 ;
        RECT 391.200 231.370 391.370 231.380 ;
        RECT 389.100 229.950 391.010 230.130 ;
        RECT 389.110 229.550 391.010 229.730 ;
        RECT 391.200 229.510 391.380 231.370 ;
        RECT 24.480 228.570 25.410 228.770 ;
        RECT 24.250 225.000 24.430 228.160 ;
        RECT 27.350 227.500 30.650 227.850 ;
        RECT 22.410 215.460 22.580 215.630 ;
        RECT 22.770 215.460 22.940 215.630 ;
        RECT 23.130 215.460 23.300 215.630 ;
        RECT 23.490 215.460 23.660 215.630 ;
        RECT 26.140 217.000 26.310 226.450 ;
        RECT 26.890 216.990 27.060 226.380 ;
        RECT 27.610 217.020 27.780 226.420 ;
        RECT 28.270 217.030 28.440 226.400 ;
        RECT 28.920 217.020 29.090 226.470 ;
        RECT 29.560 217.030 29.730 226.420 ;
        RECT 22.730 208.780 22.900 208.950 ;
        RECT 23.090 208.780 23.260 208.950 ;
        RECT 23.460 208.780 23.630 208.950 ;
        RECT 24.250 203.500 24.420 203.510 ;
        RECT 24.240 201.640 24.420 203.500 ;
        RECT 25.380 203.270 25.550 214.250 ;
        RECT 26.000 203.270 26.170 214.250 ;
        RECT 26.620 203.280 26.790 214.260 ;
        RECT 27.200 203.300 27.370 214.280 ;
        RECT 27.790 203.310 27.960 214.290 ;
        RECT 28.390 203.310 28.560 214.290 ;
        RECT 28.990 203.260 29.160 214.240 ;
        RECT 29.600 203.270 29.770 214.250 ;
        RECT 30.200 203.260 30.370 214.240 ;
        RECT 390.210 227.850 391.140 228.050 ;
        RECT 384.970 226.780 388.270 227.130 ;
        RECT 385.890 216.310 386.060 225.700 ;
        RECT 386.530 216.300 386.700 225.750 ;
        RECT 387.180 216.310 387.350 225.680 ;
        RECT 387.840 216.300 388.010 225.700 ;
        RECT 388.560 216.270 388.730 225.660 ;
        RECT 389.310 216.280 389.480 225.730 ;
        RECT 391.190 224.280 391.370 227.440 ;
        RECT 391.960 214.740 392.130 214.910 ;
        RECT 392.320 214.740 392.490 214.910 ;
        RECT 392.680 214.740 392.850 214.910 ;
        RECT 393.040 214.740 393.210 214.910 ;
        RECT 24.610 202.080 26.520 202.260 ;
        RECT 385.250 202.540 385.420 213.520 ;
        RECT 385.850 202.550 386.020 213.530 ;
        RECT 386.460 202.540 386.630 213.520 ;
        RECT 387.060 202.590 387.230 213.570 ;
        RECT 387.660 202.590 387.830 213.570 ;
        RECT 388.250 202.580 388.420 213.560 ;
        RECT 388.830 202.560 389.000 213.540 ;
        RECT 389.450 202.550 389.620 213.530 ;
        RECT 390.070 202.550 390.240 213.530 ;
        RECT 391.990 208.060 392.160 208.230 ;
        RECT 392.360 208.060 392.530 208.230 ;
        RECT 392.720 208.060 392.890 208.230 ;
        RECT 24.610 201.680 26.510 201.860 ;
        RECT 391.200 202.780 391.370 202.790 ;
        RECT 389.100 201.360 391.010 201.540 ;
        RECT 389.110 200.960 391.010 201.140 ;
        RECT 391.200 200.920 391.380 202.780 ;
        RECT 24.480 199.980 25.410 200.180 ;
        RECT 24.250 196.410 24.430 199.570 ;
        RECT 27.350 198.910 30.650 199.260 ;
        RECT 22.410 186.870 22.580 187.040 ;
        RECT 22.770 186.870 22.940 187.040 ;
        RECT 23.130 186.870 23.300 187.040 ;
        RECT 23.490 186.870 23.660 187.040 ;
        RECT 26.140 188.410 26.310 197.860 ;
        RECT 26.890 188.400 27.060 197.790 ;
        RECT 27.610 188.430 27.780 197.830 ;
        RECT 28.270 188.440 28.440 197.810 ;
        RECT 28.920 188.430 29.090 197.880 ;
        RECT 29.560 188.440 29.730 197.830 ;
        RECT 22.730 180.190 22.900 180.360 ;
        RECT 23.090 180.190 23.260 180.360 ;
        RECT 23.460 180.190 23.630 180.360 ;
        RECT 24.250 174.910 24.420 174.920 ;
        RECT 24.240 173.050 24.420 174.910 ;
        RECT 25.380 174.680 25.550 185.660 ;
        RECT 26.000 174.680 26.170 185.660 ;
        RECT 26.620 174.690 26.790 185.670 ;
        RECT 27.200 174.710 27.370 185.690 ;
        RECT 27.790 174.720 27.960 185.700 ;
        RECT 28.390 174.720 28.560 185.700 ;
        RECT 28.990 174.670 29.160 185.650 ;
        RECT 29.600 174.680 29.770 185.660 ;
        RECT 30.200 174.670 30.370 185.650 ;
        RECT 390.210 199.260 391.140 199.460 ;
        RECT 384.970 198.190 388.270 198.540 ;
        RECT 385.890 187.720 386.060 197.110 ;
        RECT 386.530 187.710 386.700 197.160 ;
        RECT 387.180 187.720 387.350 197.090 ;
        RECT 387.840 187.710 388.010 197.110 ;
        RECT 388.560 187.680 388.730 197.070 ;
        RECT 389.310 187.690 389.480 197.140 ;
        RECT 391.190 195.690 391.370 198.850 ;
        RECT 391.960 186.150 392.130 186.320 ;
        RECT 392.320 186.150 392.490 186.320 ;
        RECT 392.680 186.150 392.850 186.320 ;
        RECT 393.040 186.150 393.210 186.320 ;
        RECT 24.610 173.490 26.520 173.670 ;
        RECT 385.250 173.950 385.420 184.930 ;
        RECT 385.850 173.960 386.020 184.940 ;
        RECT 386.460 173.950 386.630 184.930 ;
        RECT 387.060 174.000 387.230 184.980 ;
        RECT 387.660 174.000 387.830 184.980 ;
        RECT 388.250 173.990 388.420 184.970 ;
        RECT 388.830 173.970 389.000 184.950 ;
        RECT 389.450 173.960 389.620 184.940 ;
        RECT 390.070 173.960 390.240 184.940 ;
        RECT 391.990 179.470 392.160 179.640 ;
        RECT 392.360 179.470 392.530 179.640 ;
        RECT 392.720 179.470 392.890 179.640 ;
        RECT 24.610 173.090 26.510 173.270 ;
        RECT 391.200 174.190 391.370 174.200 ;
        RECT 389.100 172.770 391.010 172.950 ;
        RECT 389.110 172.370 391.010 172.550 ;
        RECT 391.200 172.330 391.380 174.190 ;
        RECT 24.480 171.390 25.410 171.590 ;
        RECT 24.250 167.820 24.430 170.980 ;
        RECT 27.350 170.320 30.650 170.670 ;
        RECT 22.410 158.280 22.580 158.450 ;
        RECT 22.770 158.280 22.940 158.450 ;
        RECT 23.130 158.280 23.300 158.450 ;
        RECT 23.490 158.280 23.660 158.450 ;
        RECT 26.140 159.820 26.310 169.270 ;
        RECT 26.890 159.810 27.060 169.200 ;
        RECT 27.610 159.840 27.780 169.240 ;
        RECT 28.270 159.850 28.440 169.220 ;
        RECT 28.920 159.840 29.090 169.290 ;
        RECT 29.560 159.850 29.730 169.240 ;
        RECT 22.730 151.600 22.900 151.770 ;
        RECT 23.090 151.600 23.260 151.770 ;
        RECT 23.460 151.600 23.630 151.770 ;
        RECT 24.250 146.320 24.420 146.330 ;
        RECT 24.240 144.460 24.420 146.320 ;
        RECT 25.380 146.090 25.550 157.070 ;
        RECT 26.000 146.090 26.170 157.070 ;
        RECT 26.620 146.100 26.790 157.080 ;
        RECT 27.200 146.120 27.370 157.100 ;
        RECT 27.790 146.130 27.960 157.110 ;
        RECT 28.390 146.130 28.560 157.110 ;
        RECT 28.990 146.080 29.160 157.060 ;
        RECT 29.600 146.090 29.770 157.070 ;
        RECT 30.200 146.080 30.370 157.060 ;
        RECT 390.210 170.670 391.140 170.870 ;
        RECT 384.970 169.600 388.270 169.950 ;
        RECT 385.890 159.130 386.060 168.520 ;
        RECT 386.530 159.120 386.700 168.570 ;
        RECT 387.180 159.130 387.350 168.500 ;
        RECT 387.840 159.120 388.010 168.520 ;
        RECT 388.560 159.090 388.730 168.480 ;
        RECT 389.310 159.100 389.480 168.550 ;
        RECT 391.190 167.100 391.370 170.260 ;
        RECT 391.960 157.560 392.130 157.730 ;
        RECT 392.320 157.560 392.490 157.730 ;
        RECT 392.680 157.560 392.850 157.730 ;
        RECT 393.040 157.560 393.210 157.730 ;
        RECT 24.610 144.900 26.520 145.080 ;
        RECT 385.250 145.360 385.420 156.340 ;
        RECT 385.850 145.370 386.020 156.350 ;
        RECT 386.460 145.360 386.630 156.340 ;
        RECT 387.060 145.410 387.230 156.390 ;
        RECT 387.660 145.410 387.830 156.390 ;
        RECT 388.250 145.400 388.420 156.380 ;
        RECT 388.830 145.380 389.000 156.360 ;
        RECT 389.450 145.370 389.620 156.350 ;
        RECT 390.070 145.370 390.240 156.350 ;
        RECT 391.990 150.880 392.160 151.050 ;
        RECT 392.360 150.880 392.530 151.050 ;
        RECT 392.720 150.880 392.890 151.050 ;
        RECT 24.610 144.500 26.510 144.680 ;
        RECT 391.200 145.600 391.370 145.610 ;
        RECT 389.100 144.180 391.010 144.360 ;
        RECT 389.110 143.780 391.010 143.960 ;
        RECT 391.200 143.740 391.380 145.600 ;
        RECT 24.480 142.800 25.410 143.000 ;
        RECT 24.250 139.230 24.430 142.390 ;
        RECT 27.350 141.730 30.650 142.080 ;
        RECT 22.410 129.690 22.580 129.860 ;
        RECT 22.770 129.690 22.940 129.860 ;
        RECT 23.130 129.690 23.300 129.860 ;
        RECT 23.490 129.690 23.660 129.860 ;
        RECT 26.140 131.230 26.310 140.680 ;
        RECT 26.890 131.220 27.060 140.610 ;
        RECT 27.610 131.250 27.780 140.650 ;
        RECT 28.270 131.260 28.440 140.630 ;
        RECT 28.920 131.250 29.090 140.700 ;
        RECT 29.560 131.260 29.730 140.650 ;
        RECT 22.730 123.010 22.900 123.180 ;
        RECT 23.090 123.010 23.260 123.180 ;
        RECT 23.460 123.010 23.630 123.180 ;
        RECT 24.250 117.730 24.420 117.740 ;
        RECT 24.240 115.870 24.420 117.730 ;
        RECT 25.380 117.500 25.550 128.480 ;
        RECT 26.000 117.500 26.170 128.480 ;
        RECT 26.620 117.510 26.790 128.490 ;
        RECT 27.200 117.530 27.370 128.510 ;
        RECT 27.790 117.540 27.960 128.520 ;
        RECT 28.390 117.540 28.560 128.520 ;
        RECT 28.990 117.490 29.160 128.470 ;
        RECT 29.600 117.500 29.770 128.480 ;
        RECT 30.200 117.490 30.370 128.470 ;
        RECT 390.210 142.080 391.140 142.280 ;
        RECT 384.970 141.010 388.270 141.360 ;
        RECT 385.890 130.540 386.060 139.930 ;
        RECT 386.530 130.530 386.700 139.980 ;
        RECT 387.180 130.540 387.350 139.910 ;
        RECT 387.840 130.530 388.010 139.930 ;
        RECT 388.560 130.500 388.730 139.890 ;
        RECT 389.310 130.510 389.480 139.960 ;
        RECT 391.190 138.510 391.370 141.670 ;
        RECT 391.960 128.970 392.130 129.140 ;
        RECT 392.320 128.970 392.490 129.140 ;
        RECT 392.680 128.970 392.850 129.140 ;
        RECT 393.040 128.970 393.210 129.140 ;
        RECT 24.610 116.310 26.520 116.490 ;
        RECT 385.250 116.770 385.420 127.750 ;
        RECT 385.850 116.780 386.020 127.760 ;
        RECT 386.460 116.770 386.630 127.750 ;
        RECT 387.060 116.820 387.230 127.800 ;
        RECT 387.660 116.820 387.830 127.800 ;
        RECT 388.250 116.810 388.420 127.790 ;
        RECT 388.830 116.790 389.000 127.770 ;
        RECT 389.450 116.780 389.620 127.760 ;
        RECT 390.070 116.780 390.240 127.760 ;
        RECT 391.990 122.290 392.160 122.460 ;
        RECT 392.360 122.290 392.530 122.460 ;
        RECT 392.720 122.290 392.890 122.460 ;
        RECT 24.610 115.910 26.510 116.090 ;
        RECT 391.200 117.010 391.370 117.020 ;
        RECT 389.100 115.590 391.010 115.770 ;
        RECT 389.110 115.190 391.010 115.370 ;
        RECT 391.200 115.150 391.380 117.010 ;
        RECT 24.480 114.210 25.410 114.410 ;
        RECT 24.250 110.640 24.430 113.800 ;
        RECT 27.350 113.140 30.650 113.490 ;
        RECT 22.410 101.100 22.580 101.270 ;
        RECT 22.770 101.100 22.940 101.270 ;
        RECT 23.130 101.100 23.300 101.270 ;
        RECT 23.490 101.100 23.660 101.270 ;
        RECT 26.140 102.640 26.310 112.090 ;
        RECT 26.890 102.630 27.060 112.020 ;
        RECT 27.610 102.660 27.780 112.060 ;
        RECT 28.270 102.670 28.440 112.040 ;
        RECT 28.920 102.660 29.090 112.110 ;
        RECT 29.560 102.670 29.730 112.060 ;
        RECT 22.730 94.420 22.900 94.590 ;
        RECT 23.090 94.420 23.260 94.590 ;
        RECT 23.460 94.420 23.630 94.590 ;
        RECT 24.250 89.140 24.420 89.150 ;
        RECT 24.240 87.280 24.420 89.140 ;
        RECT 25.380 88.910 25.550 99.890 ;
        RECT 26.000 88.910 26.170 99.890 ;
        RECT 26.620 88.920 26.790 99.900 ;
        RECT 27.200 88.940 27.370 99.920 ;
        RECT 27.790 88.950 27.960 99.930 ;
        RECT 28.390 88.950 28.560 99.930 ;
        RECT 28.990 88.900 29.160 99.880 ;
        RECT 29.600 88.910 29.770 99.890 ;
        RECT 30.200 88.900 30.370 99.880 ;
        RECT 390.210 113.490 391.140 113.690 ;
        RECT 384.970 112.420 388.270 112.770 ;
        RECT 385.890 101.950 386.060 111.340 ;
        RECT 386.530 101.940 386.700 111.390 ;
        RECT 387.180 101.950 387.350 111.320 ;
        RECT 387.840 101.940 388.010 111.340 ;
        RECT 388.560 101.910 388.730 111.300 ;
        RECT 389.310 101.920 389.480 111.370 ;
        RECT 391.190 109.920 391.370 113.080 ;
        RECT 391.960 100.380 392.130 100.550 ;
        RECT 392.320 100.380 392.490 100.550 ;
        RECT 392.680 100.380 392.850 100.550 ;
        RECT 393.040 100.380 393.210 100.550 ;
        RECT 24.610 87.720 26.520 87.900 ;
        RECT 385.250 88.180 385.420 99.160 ;
        RECT 385.850 88.190 386.020 99.170 ;
        RECT 386.460 88.180 386.630 99.160 ;
        RECT 387.060 88.230 387.230 99.210 ;
        RECT 387.660 88.230 387.830 99.210 ;
        RECT 388.250 88.220 388.420 99.200 ;
        RECT 388.830 88.200 389.000 99.180 ;
        RECT 389.450 88.190 389.620 99.170 ;
        RECT 390.070 88.190 390.240 99.170 ;
        RECT 391.990 93.700 392.160 93.870 ;
        RECT 392.360 93.700 392.530 93.870 ;
        RECT 392.720 93.700 392.890 93.870 ;
        RECT 24.610 87.320 26.510 87.500 ;
        RECT 391.200 88.420 391.370 88.430 ;
        RECT 389.100 87.000 391.010 87.180 ;
        RECT 389.110 86.600 391.010 86.780 ;
        RECT 391.200 86.560 391.380 88.420 ;
      LAYER met1 ;
        RECT 24.490 457.640 25.480 457.650 ;
        RECT 24.090 457.120 25.480 457.640 ;
        RECT 24.090 453.510 24.580 457.120 ;
        RECT 27.290 456.590 30.710 456.640 ;
        RECT 27.280 456.020 30.720 456.590 ;
        RECT 25.870 446.190 30.170 455.250 ;
        RECT 31.850 455.200 32.570 455.750 ;
        RECT 31.850 455.190 32.350 455.200 ;
        RECT 32.000 446.190 32.770 446.210 ;
        RECT 23.470 444.440 32.770 446.190 ;
        RECT 22.520 444.430 32.770 444.440 ;
        RECT 22.360 444.080 32.770 444.430 ;
        RECT 22.520 444.070 32.770 444.080 ;
        RECT 23.470 443.720 32.770 444.070 ;
        RECT 23.840 442.280 32.770 443.720 ;
        RECT 21.900 437.730 22.490 441.340 ;
        RECT 21.900 437.440 23.840 437.730 ;
        RECT 23.380 432.540 24.190 433.890 ;
        RECT 25.300 432.570 30.450 442.280 ;
        RECT 32.000 442.260 32.770 442.280 ;
        RECT 35.050 434.810 35.690 438.750 ;
        RECT 23.380 432.480 24.640 432.540 ;
        RECT 23.380 431.900 24.660 432.480 ;
        RECT 25.310 431.900 30.450 432.570 ;
        RECT 23.380 431.150 24.640 431.900 ;
        RECT 23.380 430.430 32.270 431.150 ;
        RECT 23.380 430.200 26.600 430.430 ;
        RECT 23.380 430.170 24.640 430.200 ;
        RECT 23.380 429.990 24.190 430.170 ;
        RECT 24.490 429.050 25.480 429.060 ;
        RECT 24.090 428.530 25.480 429.050 ;
        RECT 24.090 424.920 24.580 428.530 ;
        RECT 27.290 428.000 30.710 428.050 ;
        RECT 27.280 427.430 30.720 428.000 ;
        RECT 25.870 417.600 30.170 426.660 ;
        RECT 31.850 426.610 32.570 427.160 ;
        RECT 31.850 426.600 32.350 426.610 ;
        RECT 32.000 417.600 32.770 417.620 ;
        RECT 23.470 415.850 32.770 417.600 ;
        RECT 22.520 415.840 32.770 415.850 ;
        RECT 22.360 415.490 32.770 415.840 ;
        RECT 22.520 415.480 32.770 415.490 ;
        RECT 23.470 415.130 32.770 415.480 ;
        RECT 23.840 413.690 32.770 415.130 ;
        RECT 21.900 409.140 22.490 412.750 ;
        RECT 21.900 408.850 23.840 409.140 ;
        RECT 23.380 403.950 24.190 405.300 ;
        RECT 25.300 403.980 30.450 413.690 ;
        RECT 32.000 413.670 32.770 413.690 ;
        RECT 35.050 406.230 35.690 410.170 ;
        RECT 23.380 403.890 24.640 403.950 ;
        RECT 23.380 403.310 24.660 403.890 ;
        RECT 25.310 403.310 30.450 403.980 ;
        RECT 23.380 402.560 24.640 403.310 ;
        RECT 23.380 401.840 32.270 402.560 ;
        RECT 23.380 401.610 26.600 401.840 ;
        RECT 23.380 401.580 24.640 401.610 ;
        RECT 23.380 401.400 24.190 401.580 ;
        RECT 24.490 400.460 25.480 400.470 ;
        RECT 24.090 399.940 25.480 400.460 ;
        RECT 24.090 396.330 24.580 399.940 ;
        RECT 27.290 399.410 30.710 399.460 ;
        RECT 27.280 398.840 30.720 399.410 ;
        RECT 25.870 390.160 30.170 398.070 ;
        RECT 31.850 398.020 32.570 398.570 ;
        RECT 31.850 398.010 32.350 398.020 ;
        RECT 23.640 389.570 30.170 390.160 ;
        RECT 23.640 389.080 23.930 389.570 ;
        RECT 25.870 389.080 30.170 389.570 ;
        RECT 30.280 389.540 30.630 389.700 ;
        RECT 58.870 389.540 59.220 389.700 ;
        RECT 87.460 389.540 87.810 389.700 ;
        RECT 171.480 389.540 171.830 389.700 ;
        RECT 200.070 389.540 200.420 389.700 ;
        RECT 228.660 389.540 229.010 389.700 ;
        RECT 257.250 389.540 257.600 389.700 ;
        RECT 285.840 389.540 286.190 389.700 ;
        RECT 314.430 389.540 314.780 389.700 ;
        RECT 343.020 389.540 343.370 389.700 ;
        RECT 23.620 389.010 30.170 389.080 ;
        RECT 30.270 389.010 30.640 389.540 ;
        RECT 32.000 389.010 32.770 389.030 ;
        RECT 16.190 387.870 20.080 388.670 ;
        RECT 16.370 387.420 18.740 387.870 ;
        RECT 16.400 385.460 17.350 387.420 ;
        RECT 18.100 387.400 18.680 387.420 ;
        RECT 23.470 387.260 32.770 389.010 ;
        RECT 39.710 387.570 43.840 387.970 ;
        RECT 44.780 387.870 48.670 388.670 ;
        RECT 58.860 388.590 59.230 389.540 ;
        RECT 58.510 388.220 60.980 388.590 ;
        RECT 39.710 387.480 43.850 387.570 ;
        RECT 22.520 387.250 32.770 387.260 ;
        RECT 22.360 386.900 32.770 387.250 ;
        RECT 22.520 386.890 32.770 386.900 ;
        RECT 23.470 386.760 32.770 386.890 ;
        RECT 18.770 386.750 32.770 386.760 ;
        RECT 16.630 379.790 17.350 385.460 ;
        RECT 18.100 386.190 32.770 386.750 ;
        RECT 43.320 386.580 43.850 387.480 ;
        RECT 44.960 387.420 47.330 387.870 ;
        RECT 18.100 381.890 41.450 386.190 ;
        RECT 44.990 385.460 45.940 387.420 ;
        RECT 46.690 387.400 47.270 387.420 ;
        RECT 57.070 386.760 60.980 388.220 ;
        RECT 68.300 387.570 72.430 387.970 ;
        RECT 73.370 387.870 77.260 388.670 ;
        RECT 87.450 388.590 87.820 389.540 ;
        RECT 87.100 388.220 89.570 388.590 ;
        RECT 68.300 387.480 72.440 387.570 ;
        RECT 47.360 386.750 60.980 386.760 ;
        RECT 42.220 384.770 42.790 384.780 ;
        RECT 18.100 381.610 32.390 381.890 ;
        RECT 21.900 380.550 22.490 381.610 ;
        RECT 21.900 380.260 23.840 380.550 ;
        RECT 25.300 380.060 32.390 381.610 ;
        RECT 25.300 379.290 32.410 380.060 ;
        RECT 25.300 378.700 30.450 379.290 ;
        RECT 21.010 376.230 24.960 377.000 ;
        RECT 23.380 375.360 24.190 376.230 ;
        RECT 25.300 375.390 32.370 378.700 ;
        RECT 35.060 377.620 35.700 381.560 ;
        RECT 42.220 381.350 42.840 384.770 ;
        RECT 42.220 381.340 42.790 381.350 ;
        RECT 41.390 379.710 41.950 380.210 ;
        RECT 45.220 379.790 45.940 385.460 ;
        RECT 46.690 386.190 60.980 386.750 ;
        RECT 71.910 386.580 72.440 387.480 ;
        RECT 73.550 387.420 75.920 387.870 ;
        RECT 46.690 381.890 70.040 386.190 ;
        RECT 73.580 385.460 74.530 387.420 ;
        RECT 75.280 387.400 75.860 387.420 ;
        RECT 85.660 386.760 89.570 388.220 ;
        RECT 96.890 387.570 101.020 387.970 ;
        RECT 115.270 387.890 119.160 388.690 ;
        RECT 142.760 387.820 145.170 388.460 ;
        RECT 96.890 387.480 101.030 387.570 ;
        RECT 75.950 386.750 89.570 386.760 ;
        RECT 70.810 384.770 71.380 384.780 ;
        RECT 46.690 381.610 60.980 381.890 ;
        RECT 57.070 380.060 60.980 381.610 ;
        RECT 70.810 381.350 71.430 384.770 ;
        RECT 70.810 381.340 71.380 381.350 ;
        RECT 41.400 379.490 41.950 379.710 ;
        RECT 57.050 379.290 61.000 380.060 ;
        RECT 69.980 379.710 70.540 380.210 ;
        RECT 73.810 379.790 74.530 385.460 ;
        RECT 75.280 386.190 89.570 386.750 ;
        RECT 100.500 386.580 101.030 387.480 ;
        RECT 142.780 386.470 143.190 387.820 ;
        RECT 149.510 387.160 149.920 387.930 ;
        RECT 157.390 387.870 161.280 388.670 ;
        RECT 171.470 388.590 171.840 389.540 ;
        RECT 171.120 388.220 173.590 388.590 ;
        RECT 157.570 387.420 159.940 387.870 ;
        RECT 149.240 386.890 149.920 387.160 ;
        RECT 149.240 386.460 150.930 386.890 ;
        RECT 122.030 386.280 146.400 386.300 ;
        RECT 75.280 381.890 98.630 386.190 ;
        RECT 121.970 385.890 146.400 386.280 ;
        RECT 99.400 384.770 99.970 384.780 ;
        RECT 75.280 381.610 89.570 381.890 ;
        RECT 85.660 380.060 89.570 381.610 ;
        RECT 99.400 381.350 100.020 384.770 ;
        RECT 99.400 381.340 99.970 381.350 ;
        RECT 69.990 379.490 70.540 379.710 ;
        RECT 85.640 379.290 89.590 380.060 ;
        RECT 98.570 379.710 99.130 380.210 ;
        RECT 98.580 379.490 99.130 379.710 ;
        RECT 49.610 376.230 53.560 377.000 ;
        RECT 23.380 375.300 24.640 375.360 ;
        RECT 23.380 374.720 24.660 375.300 ;
        RECT 25.310 374.720 32.370 375.390 ;
        RECT 23.380 373.970 24.640 374.720 ;
        RECT 29.140 373.970 32.370 374.720 ;
        RECT 23.380 373.250 32.370 373.970 ;
        RECT 23.380 373.020 26.600 373.250 ;
        RECT 23.380 372.990 24.640 373.020 ;
        RECT 23.380 372.810 24.190 372.990 ;
        RECT 24.490 371.870 25.480 371.880 ;
        RECT 24.090 371.350 25.480 371.870 ;
        RECT 24.090 367.740 24.580 371.350 ;
        RECT 29.140 370.870 32.370 373.250 ;
        RECT 27.290 370.820 32.370 370.870 ;
        RECT 27.280 370.250 32.370 370.820 ;
        RECT 29.140 369.980 32.370 370.250 ;
        RECT 29.140 369.480 32.570 369.980 ;
        RECT 25.870 369.430 32.570 369.480 ;
        RECT 25.870 361.970 32.370 369.430 ;
        RECT 57.730 369.000 60.960 378.700 ;
        RECT 78.190 376.230 82.140 377.000 ;
        RECT 86.320 373.290 89.550 378.700 ;
        RECT 121.970 377.640 122.380 385.890 ;
        RECT 132.240 382.020 132.740 382.500 ;
        RECT 125.200 381.640 125.440 382.000 ;
        RECT 132.340 379.060 132.730 382.020 ;
        RECT 139.890 381.610 140.150 382.400 ;
        RECT 144.590 381.560 144.850 382.350 ;
        RECT 125.780 378.650 126.040 378.950 ;
        RECT 128.640 378.810 128.900 379.000 ;
        RECT 128.640 378.680 129.010 378.810 ;
        RECT 125.780 378.630 126.190 378.650 ;
        RECT 125.810 378.340 126.190 378.630 ;
        RECT 127.220 378.340 128.250 378.650 ;
        RECT 128.720 378.580 129.010 378.680 ;
        RECT 125.770 377.780 126.030 377.920 ;
        RECT 125.770 377.600 126.120 377.780 ;
        RECT 126.410 377.620 126.730 377.940 ;
        RECT 127.180 377.780 127.440 377.930 ;
        RECT 127.180 377.610 127.520 377.780 ;
        RECT 125.880 377.550 126.120 377.600 ;
        RECT 127.290 377.550 127.520 377.610 ;
        RECT 125.820 377.470 127.570 377.550 ;
        RECT 125.770 377.150 127.570 377.470 ;
        RECT 125.820 377.050 127.570 377.150 ;
        RECT 98.860 376.490 99.030 376.610 ;
        RECT 85.890 370.550 89.720 373.290 ;
        RECT 98.510 369.930 99.030 376.490 ;
        RECT 98.450 369.420 99.100 369.930 ;
        RECT 57.570 366.110 61.070 369.000 ;
        RECT 14.530 361.890 17.920 361.960 ;
        RECT 13.560 361.800 17.920 361.890 ;
        RECT 10.330 358.570 17.920 361.800 ;
        RECT 25.870 360.420 30.170 361.970 ;
        RECT 98.510 361.740 99.030 369.420 ;
        RECT 101.910 365.510 102.320 376.720 ;
        RECT 120.960 376.230 123.440 377.000 ;
        RECT 125.770 376.890 127.570 377.050 ;
        RECT 125.770 376.730 126.120 376.890 ;
        RECT 126.410 376.780 126.730 376.890 ;
        RECT 127.200 376.750 127.520 376.890 ;
        RECT 125.880 376.670 126.120 376.730 ;
        RECT 127.290 376.670 127.520 376.750 ;
        RECT 125.880 375.700 126.110 376.120 ;
        RECT 125.770 375.380 126.110 375.700 ;
        RECT 125.880 374.710 126.110 375.380 ;
        RECT 127.290 374.710 127.520 376.120 ;
        RECT 128.010 375.940 128.250 378.340 ;
        RECT 132.340 378.570 132.810 379.060 ;
        RECT 132.340 378.560 132.790 378.570 ;
        RECT 138.880 378.560 139.120 379.200 ;
        RECT 139.890 378.620 140.150 379.410 ;
        RECT 144.090 378.640 144.330 379.050 ;
        RECT 128.730 377.890 129.000 378.020 ;
        RECT 128.410 377.660 129.090 377.890 ;
        RECT 128.300 377.300 128.620 377.620 ;
        RECT 128.670 377.600 129.090 377.660 ;
        RECT 128.350 377.070 128.580 377.300 ;
        RECT 128.860 376.660 129.090 377.600 ;
        RECT 128.730 376.630 129.090 376.660 ;
        RECT 128.730 376.480 130.180 376.630 ;
        RECT 128.730 376.460 129.000 376.480 ;
        RECT 128.410 376.230 129.000 376.460 ;
        RECT 127.920 375.650 128.250 375.940 ;
        RECT 128.010 375.570 128.250 375.650 ;
        RECT 128.110 374.880 128.430 375.200 ;
        RECT 128.730 375.190 129.000 376.230 ;
        RECT 129.020 375.190 130.180 376.480 ;
        RECT 128.730 374.960 130.180 375.190 ;
        RECT 129.020 374.720 130.180 374.960 ;
        RECT 132.340 374.720 132.730 378.560 ;
        RECT 138.880 378.300 139.110 378.560 ;
        RECT 138.870 378.080 139.110 378.300 ;
        RECT 133.750 377.420 134.010 377.740 ;
        RECT 139.890 377.610 140.150 378.400 ;
        RECT 148.570 378.390 150.930 386.460 ;
        RECT 157.600 386.300 158.550 387.420 ;
        RECT 159.300 387.400 159.880 387.420 ;
        RECT 169.680 386.760 173.590 388.220 ;
        RECT 180.910 387.570 185.040 387.970 ;
        RECT 185.980 387.870 189.870 388.670 ;
        RECT 200.060 388.590 200.430 389.540 ;
        RECT 199.710 388.220 202.180 388.590 ;
        RECT 180.910 387.480 185.050 387.570 ;
        RECT 159.970 386.750 173.590 386.760 ;
        RECT 159.300 386.300 173.590 386.750 ;
        RECT 184.520 386.580 185.050 387.480 ;
        RECT 186.160 387.420 188.530 387.870 ;
        RECT 155.200 386.290 176.560 386.300 ;
        RECT 155.140 386.190 176.560 386.290 ;
        RECT 155.140 385.890 182.650 386.190 ;
        RECT 157.600 385.460 158.550 385.890 ;
        RECT 157.830 383.310 158.550 385.460 ;
        RECT 159.300 383.310 182.650 385.890 ;
        RECT 186.190 385.460 187.140 387.420 ;
        RECT 187.890 387.400 188.470 387.420 ;
        RECT 198.270 386.760 202.180 388.220 ;
        RECT 209.500 387.570 213.630 387.970 ;
        RECT 214.580 387.870 218.470 388.670 ;
        RECT 228.650 388.590 229.020 389.540 ;
        RECT 228.300 388.220 230.770 388.590 ;
        RECT 209.500 387.480 213.640 387.570 ;
        RECT 188.560 386.750 202.180 386.760 ;
        RECT 157.830 382.300 182.650 383.310 ;
        RECT 152.930 381.700 155.700 381.940 ;
        RECT 152.930 381.290 153.170 381.700 ;
        RECT 148.450 377.570 150.930 378.390 ;
        RECT 154.640 378.160 154.900 379.050 ;
        RECT 133.760 375.200 134.000 377.420 ;
        RECT 141.800 376.880 142.120 377.200 ;
        RECT 143.160 376.960 143.480 377.280 ;
        RECT 143.850 376.950 144.170 377.270 ;
        RECT 138.880 375.760 139.120 376.400 ;
        RECT 138.880 375.500 139.110 375.760 ;
        RECT 138.870 375.280 139.110 375.500 ;
        RECT 133.670 374.720 134.090 375.200 ;
        RECT 138.880 374.720 139.120 374.850 ;
        RECT 139.560 374.720 139.850 375.880 ;
        RECT 144.080 374.720 144.320 374.880 ;
        RECT 149.900 374.720 150.210 375.590 ;
        RECT 152.920 374.720 153.160 375.830 ;
        RECT 153.250 374.720 153.480 375.650 ;
        RECT 153.860 374.720 154.110 375.050 ;
        RECT 155.460 374.720 155.700 381.700 ;
        RECT 157.830 379.790 158.550 382.300 ;
        RECT 159.300 381.890 182.650 382.300 ;
        RECT 183.420 384.770 183.990 384.780 ;
        RECT 159.300 381.640 173.590 381.890 ;
        RECT 158.770 381.610 173.590 381.640 ;
        RECT 158.770 381.370 161.800 381.610 ;
        RECT 163.480 381.380 163.740 381.610 ;
        RECT 126.390 373.980 126.710 374.300 ;
        RECT 127.820 374.000 128.140 374.320 ;
        RECT 125.600 373.400 125.920 373.720 ;
        RECT 126.530 373.400 126.850 373.720 ;
        RECT 127.230 373.400 127.550 373.720 ;
        RECT 127.970 373.400 128.290 373.720 ;
        RECT 128.680 373.390 129.000 373.710 ;
        RECT 129.020 373.590 156.380 374.720 ;
        RECT 129.020 373.390 156.570 373.590 ;
        RECT 130.720 373.000 131.010 373.390 ;
        RECT 101.790 365.040 102.320 365.510 ;
        RECT 98.310 361.010 99.030 361.740 ;
        RECT 32.000 360.420 32.770 360.440 ;
        RECT 23.470 358.670 32.770 360.420 ;
        RECT 22.520 358.660 32.770 358.670 ;
        RECT 13.560 357.890 17.920 358.570 ;
        RECT 22.360 358.310 32.770 358.660 ;
        RECT 22.520 358.300 32.770 358.310 ;
        RECT 23.470 357.950 32.770 358.300 ;
        RECT 23.840 356.510 32.770 357.950 ;
        RECT 21.900 351.960 22.490 355.570 ;
        RECT 21.900 351.670 23.840 351.960 ;
        RECT 23.390 346.770 24.200 348.120 ;
        RECT 25.300 346.800 30.450 356.510 ;
        RECT 32.000 356.490 32.770 356.510 ;
        RECT 35.050 349.040 35.690 352.980 ;
        RECT 23.390 346.710 24.640 346.770 ;
        RECT 23.390 346.130 24.660 346.710 ;
        RECT 25.310 346.130 30.450 346.800 ;
        RECT 23.390 345.380 24.640 346.130 ;
        RECT 23.390 344.660 32.270 345.380 ;
        RECT 23.390 344.430 26.600 344.660 ;
        RECT 23.390 344.400 24.640 344.430 ;
        RECT 23.390 344.220 24.200 344.400 ;
        RECT 24.490 343.280 25.480 343.290 ;
        RECT 24.090 342.760 25.480 343.280 ;
        RECT 24.090 339.150 24.580 342.760 ;
        RECT 27.290 342.230 30.710 342.280 ;
        RECT 27.280 341.660 30.720 342.230 ;
        RECT 25.870 333.250 30.170 340.890 ;
        RECT 31.850 340.840 32.570 341.390 ;
        RECT 31.850 340.830 32.350 340.840 ;
        RECT 23.700 333.210 30.170 333.250 ;
        RECT 10.330 331.830 30.170 333.210 ;
        RECT 32.000 331.830 32.770 331.850 ;
        RECT 10.330 329.980 32.770 331.830 ;
        RECT 22.360 329.720 32.770 329.980 ;
        RECT 22.520 329.710 32.770 329.720 ;
        RECT 23.470 329.360 32.770 329.710 ;
        RECT 23.840 327.920 32.770 329.360 ;
        RECT 21.900 323.370 22.490 326.980 ;
        RECT 21.900 323.080 23.840 323.370 ;
        RECT 23.380 318.180 24.190 319.530 ;
        RECT 25.300 318.210 30.450 327.920 ;
        RECT 32.000 327.900 32.770 327.920 ;
        RECT 98.510 325.660 99.030 361.010 ;
        RECT 101.910 360.790 102.320 365.040 ;
        RECT 101.770 360.200 102.390 360.790 ;
        RECT 98.430 325.060 99.060 325.660 ;
        RECT 101.910 324.640 102.320 360.200 ;
        RECT 35.060 320.460 35.700 324.400 ;
        RECT 101.860 324.140 102.340 324.640 ;
        RECT 132.340 320.450 132.730 373.390 ;
        RECT 139.540 373.290 139.950 373.390 ;
        RECT 141.080 373.220 141.400 373.390 ;
        RECT 144.080 373.000 144.320 373.390 ;
        RECT 149.900 373.000 150.210 373.390 ;
        RECT 150.940 373.240 151.260 373.390 ;
        RECT 152.920 372.600 153.160 373.390 ;
        RECT 153.860 373.180 154.110 373.390 ;
        RECT 153.860 373.000 154.120 373.180 ;
        RECT 152.870 372.260 153.210 372.600 ;
        RECT 150.120 372.160 150.610 372.170 ;
        RECT 147.300 368.580 147.620 368.900 ;
        RECT 148.390 368.590 148.710 368.910 ;
        RECT 145.760 367.670 146.080 367.990 ;
        RECT 147.310 367.590 147.630 367.910 ;
        RECT 145.740 366.750 146.060 367.070 ;
        RECT 145.720 365.760 146.040 366.080 ;
        RECT 146.190 363.470 146.420 366.950 ;
        RECT 146.860 366.330 147.080 366.950 ;
        RECT 147.310 366.600 147.630 366.920 ;
        RECT 146.830 366.010 147.090 366.330 ;
        RECT 146.860 365.450 147.080 366.010 ;
        RECT 147.220 365.870 147.540 366.190 ;
        RECT 147.310 365.450 147.630 365.490 ;
        RECT 146.860 365.410 147.630 365.450 ;
        RECT 146.800 365.220 147.630 365.410 ;
        RECT 146.800 365.090 147.080 365.220 ;
        RECT 147.310 365.200 147.630 365.220 ;
        RECT 146.860 364.490 147.080 365.090 ;
        RECT 147.220 365.170 147.630 365.200 ;
        RECT 147.220 364.880 147.540 365.170 ;
        RECT 146.810 364.460 147.080 364.490 ;
        RECT 147.310 364.460 147.630 364.500 ;
        RECT 146.810 364.230 147.630 364.460 ;
        RECT 146.810 364.170 147.080 364.230 ;
        RECT 147.310 364.210 147.630 364.230 ;
        RECT 146.160 363.150 146.420 363.470 ;
        RECT 146.190 362.510 146.420 363.150 ;
        RECT 146.120 362.190 146.420 362.510 ;
        RECT 146.190 361.550 146.420 362.190 ;
        RECT 146.160 361.230 146.420 361.550 ;
        RECT 146.190 346.480 146.420 361.230 ;
        RECT 146.860 363.470 147.080 364.170 ;
        RECT 147.220 364.180 147.630 364.210 ;
        RECT 147.220 363.890 147.540 364.180 ;
        RECT 147.640 363.780 147.860 368.390 ;
        RECT 147.620 363.710 147.860 363.780 ;
        RECT 148.040 367.840 148.260 368.390 ;
        RECT 148.040 367.550 148.360 367.840 ;
        RECT 148.400 367.600 148.720 367.920 ;
        RECT 147.620 363.610 147.960 363.710 ;
        RECT 147.310 363.470 147.630 363.510 ;
        RECT 146.860 363.240 147.630 363.470 ;
        RECT 146.860 346.480 147.080 363.240 ;
        RECT 147.310 363.190 147.630 363.240 ;
        RECT 147.640 363.480 147.960 363.610 ;
        RECT 147.640 362.510 147.860 363.480 ;
        RECT 148.040 362.510 148.260 367.550 ;
        RECT 148.400 366.610 148.720 366.930 ;
        RECT 149.550 366.670 149.770 371.220 ;
        RECT 150.110 371.010 150.620 372.160 ;
        RECT 155.050 371.990 156.380 373.390 ;
        RECT 158.740 372.200 159.050 375.900 ;
        RECT 155.460 371.230 155.700 371.990 ;
        RECT 158.660 371.830 159.050 372.200 ;
        RECT 161.530 371.690 161.800 381.370 ;
        RECT 169.680 380.060 173.590 381.610 ;
        RECT 169.660 379.290 173.610 380.060 ;
        RECT 175.250 379.950 175.670 381.890 ;
        RECT 183.420 381.350 184.040 384.770 ;
        RECT 183.420 381.340 183.990 381.350 ;
        RECT 175.250 379.470 175.720 379.950 ;
        RECT 182.590 379.710 183.150 380.210 ;
        RECT 182.600 379.490 183.150 379.710 ;
        RECT 171.440 379.190 171.860 379.290 ;
        RECT 171.400 378.710 171.880 379.190 ;
        RECT 162.210 376.240 166.160 377.010 ;
        RECT 162.700 372.690 162.950 375.840 ;
        RECT 169.740 373.340 170.060 373.390 ;
        RECT 169.650 373.050 170.060 373.340 ;
        RECT 162.660 372.330 162.990 372.690 ;
        RECT 169.230 372.050 169.470 372.120 ;
        RECT 161.490 371.380 161.830 371.690 ;
        RECT 169.260 371.630 169.500 371.680 ;
        RECT 150.060 370.910 150.620 371.010 ;
        RECT 155.410 370.910 155.750 371.230 ;
        RECT 149.950 370.510 150.620 370.910 ;
        RECT 149.950 370.480 150.610 370.510 ;
        RECT 149.950 366.670 150.170 370.480 ;
        RECT 169.230 370.300 169.470 370.370 ;
        RECT 169.650 369.550 169.890 373.050 ;
        RECT 170.340 372.480 173.570 378.710 ;
        RECT 176.950 377.100 177.390 377.600 ;
        RECT 182.670 377.100 183.110 377.600 ;
        RECT 172.010 372.120 172.250 372.480 ;
        RECT 172.010 372.060 172.480 372.120 ;
        RECT 172.010 371.680 172.250 372.060 ;
        RECT 172.010 371.620 172.510 371.680 ;
        RECT 171.270 371.040 171.680 371.370 ;
        RECT 172.010 370.860 172.250 371.620 ;
        RECT 172.010 370.370 172.250 370.790 ;
        RECT 172.010 370.310 172.480 370.370 ;
        RECT 171.270 369.290 171.680 369.620 ;
        RECT 172.010 369.110 172.250 370.310 ;
        RECT 172.590 369.480 172.900 372.480 ;
        RECT 173.430 371.900 173.780 372.190 ;
        RECT 173.430 371.880 173.630 371.900 ;
        RECT 174.390 371.690 174.700 371.700 ;
        RECT 174.390 371.420 174.710 371.690 ;
        RECT 174.410 371.410 174.700 371.420 ;
        RECT 174.950 370.860 175.260 372.550 ;
        RECT 175.430 371.480 175.750 371.760 ;
        RECT 176.500 371.680 176.790 372.120 ;
        RECT 176.500 371.590 176.820 371.680 ;
        RECT 175.430 371.460 175.790 371.480 ;
        RECT 175.510 371.150 175.790 371.460 ;
        RECT 173.430 370.150 173.780 370.440 ;
        RECT 173.430 370.130 173.630 370.150 ;
        RECT 174.390 369.940 174.700 369.950 ;
        RECT 174.390 369.670 174.710 369.940 ;
        RECT 174.410 369.660 174.700 369.670 ;
        RECT 174.950 369.110 175.260 370.800 ;
        RECT 175.430 369.730 175.750 370.010 ;
        RECT 175.430 369.710 175.790 369.730 ;
        RECT 175.510 369.400 175.790 369.710 ;
        RECT 151.170 368.360 151.520 368.820 ;
        RECT 167.600 368.380 167.970 368.690 ;
        RECT 172.010 368.620 172.250 369.040 ;
        RECT 169.230 368.550 169.470 368.620 ;
        RECT 172.010 368.560 172.480 368.620 ;
        RECT 150.570 368.000 150.820 368.120 ;
        RECT 150.540 367.540 150.860 368.000 ;
        RECT 150.570 366.750 150.820 367.540 ;
        RECT 150.570 366.430 150.860 366.750 ;
        RECT 148.520 365.770 148.840 366.090 ;
        RECT 150.570 365.830 150.820 366.430 ;
        RECT 150.570 365.510 150.860 365.830 ;
        RECT 148.520 364.780 148.840 365.100 ;
        RECT 150.570 364.910 150.820 365.510 ;
        RECT 150.570 364.590 150.830 364.910 ;
        RECT 148.520 363.790 148.840 364.110 ;
        RECT 146.080 345.950 146.420 346.480 ;
        RECT 146.740 345.950 147.080 346.480 ;
        RECT 144.770 345.210 145.000 345.280 ;
        RECT 144.730 344.950 145.050 345.210 ;
        RECT 144.280 344.840 144.510 344.880 ;
        RECT 144.240 344.520 144.510 344.840 ;
        RECT 134.930 343.280 135.650 343.980 ;
        RECT 134.940 338.130 135.600 343.280 ;
        RECT 144.280 341.000 144.510 344.520 ;
        RECT 144.770 342.480 145.000 344.950 ;
        RECT 146.190 344.860 146.420 345.950 ;
        RECT 146.860 345.220 147.080 345.950 ;
        RECT 148.620 345.240 148.890 345.280 ;
        RECT 146.840 344.900 147.100 345.220 ;
        RECT 148.600 344.910 148.890 345.240 ;
        RECT 146.180 344.540 146.440 344.860 ;
        RECT 148.070 343.370 148.360 343.400 ;
        RECT 144.770 342.110 145.500 342.480 ;
        RECT 144.280 340.930 144.540 341.000 ;
        RECT 144.260 340.920 144.540 340.930 ;
        RECT 144.230 340.610 144.550 340.920 ;
        RECT 140.130 338.750 140.560 339.180 ;
        RECT 134.940 337.410 135.680 338.130 ;
        RECT 140.180 332.940 140.550 338.750 ;
        RECT 144.090 337.370 144.410 337.690 ;
        RECT 144.770 337.020 145.000 342.110 ;
        RECT 148.620 341.940 148.890 344.910 ;
        RECT 148.500 341.690 148.890 341.940 ;
        RECT 149.100 344.840 149.340 344.880 ;
        RECT 149.100 344.520 149.360 344.840 ;
        RECT 149.100 341.380 149.340 344.520 ;
        RECT 148.500 341.150 149.340 341.380 ;
        RECT 147.400 337.810 147.720 338.130 ;
        RECT 145.190 337.380 145.510 337.700 ;
        RECT 146.280 337.380 146.600 337.700 ;
        RECT 147.410 337.340 147.730 337.660 ;
        RECT 144.640 336.700 145.000 337.020 ;
        RECT 145.740 336.700 146.060 337.020 ;
        RECT 146.840 336.700 147.160 337.020 ;
        RECT 144.770 335.650 145.000 336.700 ;
        RECT 147.690 336.680 147.980 337.110 ;
        RECT 147.690 336.660 148.160 336.680 ;
        RECT 147.700 336.360 148.160 336.660 ;
        RECT 147.700 335.830 147.980 336.360 ;
        RECT 147.710 335.800 147.980 335.830 ;
        RECT 144.640 335.330 145.000 335.650 ;
        RECT 145.740 335.330 146.060 335.650 ;
        RECT 146.840 335.330 147.160 335.650 ;
        RECT 144.090 334.600 144.410 334.920 ;
        RECT 144.770 334.610 145.000 335.330 ;
        RECT 145.190 334.610 145.510 334.920 ;
        RECT 146.280 334.610 146.600 334.920 ;
        RECT 144.770 334.380 147.220 334.610 ;
        RECT 146.900 334.050 147.220 334.380 ;
        RECT 144.080 333.260 144.400 333.580 ;
        RECT 145.190 333.250 145.510 333.570 ;
        RECT 146.280 333.230 146.600 333.550 ;
        RECT 140.140 332.510 140.570 332.940 ;
        RECT 144.640 332.560 144.960 332.880 ;
        RECT 145.740 332.550 146.060 332.870 ;
        RECT 146.830 332.550 147.150 332.870 ;
        RECT 147.660 332.480 147.990 332.510 ;
        RECT 147.520 332.400 147.990 332.480 ;
        RECT 147.280 332.160 147.990 332.400 ;
        RECT 147.660 332.090 147.990 332.160 ;
        RECT 143.150 326.850 143.440 327.200 ;
        RECT 143.160 326.280 143.420 326.850 ;
        RECT 143.800 325.750 144.060 330.730 ;
        RECT 147.440 330.250 147.760 330.570 ;
        RECT 144.130 329.810 144.450 330.130 ;
        RECT 145.230 329.820 145.550 330.140 ;
        RECT 146.320 329.820 146.640 330.140 ;
        RECT 147.450 329.780 147.770 330.100 ;
        RECT 144.680 329.140 145.000 329.460 ;
        RECT 145.780 329.140 146.100 329.460 ;
        RECT 146.880 329.140 147.200 329.460 ;
        RECT 144.680 327.770 145.000 328.090 ;
        RECT 145.780 327.770 146.100 328.090 ;
        RECT 146.880 327.770 147.200 328.090 ;
        RECT 144.130 327.040 144.450 327.360 ;
        RECT 145.230 327.040 145.550 327.360 ;
        RECT 146.320 327.040 146.640 327.360 ;
        RECT 149.100 326.490 149.340 341.150 ;
        RECT 149.550 340.480 149.770 361.230 ;
        RECT 149.950 343.090 150.170 361.230 ;
        RECT 150.570 344.240 150.820 364.590 ;
        RECT 151.190 363.820 151.450 368.360 ;
        RECT 166.960 366.660 167.350 367.030 ;
        RECT 166.380 365.170 166.770 365.560 ;
        RECT 151.190 363.500 151.470 363.820 ;
        RECT 165.740 363.580 166.130 363.960 ;
        RECT 165.770 363.570 166.110 363.580 ;
        RECT 151.190 362.860 151.450 363.500 ;
        RECT 165.130 363.380 165.470 363.390 ;
        RECT 165.120 362.990 165.480 363.380 ;
        RECT 151.190 362.540 151.480 362.860 ;
        RECT 151.190 361.900 151.450 362.540 ;
        RECT 151.190 361.580 151.470 361.900 ;
        RECT 150.570 344.220 150.830 344.240 ;
        RECT 150.560 343.940 150.840 344.220 ;
        RECT 150.570 343.920 150.830 343.940 ;
        RECT 149.910 342.770 150.230 343.090 ;
        RECT 149.950 341.180 150.170 342.770 ;
        RECT 150.570 342.480 150.820 343.920 ;
        RECT 150.490 342.160 150.820 342.480 ;
        RECT 149.950 340.860 150.280 341.180 ;
        RECT 149.950 340.700 150.170 340.860 ;
        RECT 149.850 340.500 150.170 340.700 ;
        RECT 149.510 340.160 149.790 340.480 ;
        RECT 149.850 340.190 150.270 340.500 ;
        RECT 149.550 327.190 149.770 340.160 ;
        RECT 149.950 339.990 150.270 340.190 ;
        RECT 149.950 339.630 150.170 339.990 ;
        RECT 149.950 339.310 150.280 339.630 ;
        RECT 149.950 334.950 150.170 339.310 ;
        RECT 150.570 338.600 150.820 342.160 ;
        RECT 151.190 342.480 151.450 361.580 ;
        RECT 164.510 361.430 164.870 361.820 ;
        RECT 163.860 359.890 164.270 360.290 ;
        RECT 163.330 358.330 163.690 358.720 ;
        RECT 162.750 353.270 163.080 353.290 ;
        RECT 162.690 352.850 163.080 353.270 ;
        RECT 162.120 351.660 162.450 351.680 ;
        RECT 162.070 351.270 162.460 351.660 ;
        RECT 161.500 350.110 161.830 350.120 ;
        RECT 161.470 349.720 161.830 350.110 ;
        RECT 160.850 348.240 161.240 348.640 ;
        RECT 160.180 343.070 160.610 343.470 ;
        RECT 151.710 342.600 152.030 342.920 ;
        RECT 152.360 342.600 152.680 342.920 ;
        RECT 151.190 342.160 151.510 342.480 ;
        RECT 151.190 339.910 151.450 342.160 ;
        RECT 152.740 341.300 153.030 342.210 ;
        RECT 159.520 341.500 159.930 341.900 ;
        RECT 152.390 340.640 152.710 340.680 ;
        RECT 152.390 340.410 152.940 340.640 ;
        RECT 153.200 340.500 153.210 340.730 ;
        RECT 152.390 340.360 152.710 340.410 ;
        RECT 152.400 340.100 152.720 340.140 ;
        RECT 151.180 339.590 151.490 339.910 ;
        RECT 152.400 339.870 152.950 340.100 ;
        RECT 152.400 339.820 152.720 339.870 ;
        RECT 158.910 339.860 159.300 340.260 ;
        RECT 150.520 338.280 150.840 338.600 ;
        RECT 151.190 338.590 151.450 339.590 ;
        RECT 152.730 339.280 153.000 339.460 ;
        RECT 152.710 338.960 153.030 339.280 ;
        RECT 152.730 338.790 153.000 338.960 ;
        RECT 149.950 334.470 150.240 334.950 ;
        RECT 149.950 332.510 150.170 334.470 ;
        RECT 149.930 332.090 150.190 332.510 ;
        RECT 149.950 327.470 150.170 332.090 ;
        RECT 150.570 328.850 150.820 338.280 ;
        RECT 151.190 338.270 151.530 338.590 ;
        RECT 158.220 338.420 158.630 338.810 ;
        RECT 150.530 328.450 150.830 328.850 ;
        RECT 149.950 327.330 150.190 327.470 ;
        RECT 149.510 326.840 149.820 327.190 ;
        RECT 149.960 326.700 150.190 327.330 ;
        RECT 143.750 324.940 144.060 325.750 ;
        RECT 144.120 325.700 144.440 326.020 ;
        RECT 145.230 325.690 145.550 326.010 ;
        RECT 146.320 325.670 146.640 325.990 ;
        RECT 148.310 325.930 149.340 326.490 ;
        RECT 149.950 326.670 150.190 326.700 ;
        RECT 148.310 325.820 149.100 325.930 ;
        RECT 144.680 325.000 145.000 325.320 ;
        RECT 145.780 324.990 146.100 325.310 ;
        RECT 146.870 324.990 147.190 325.310 ;
        RECT 149.950 325.280 150.170 326.670 ;
        RECT 143.800 324.740 144.060 324.940 ;
        RECT 148.420 321.600 150.840 325.280 ;
        RECT 151.190 321.310 151.450 338.270 ;
        RECT 151.690 337.500 152.010 337.820 ;
        RECT 152.400 337.440 152.720 337.760 ;
        RECT 154.010 333.270 154.940 334.920 ;
        RECT 154.100 332.790 154.840 333.270 ;
        RECT 151.100 320.900 151.450 321.310 ;
        RECT 132.170 319.930 132.730 320.450 ;
        RECT 23.380 318.120 24.640 318.180 ;
        RECT 23.380 317.540 24.660 318.120 ;
        RECT 25.310 317.540 30.450 318.210 ;
        RECT 23.380 316.790 24.640 317.540 ;
        RECT 23.380 316.070 32.270 316.790 ;
        RECT 23.380 315.840 26.600 316.070 ;
        RECT 23.380 315.810 24.640 315.840 ;
        RECT 23.380 315.630 24.190 315.810 ;
        RECT 158.280 315.080 158.610 338.420 ;
        RECT 158.230 315.070 158.660 315.080 ;
        RECT 24.490 314.690 25.480 314.700 ;
        RECT 24.090 314.170 25.480 314.690 ;
        RECT 158.200 314.610 158.690 315.070 ;
        RECT 158.230 314.590 158.660 314.610 ;
        RECT 158.930 314.290 159.260 339.860 ;
        RECT 24.090 310.560 24.580 314.170 ;
        RECT 158.840 313.800 159.330 314.290 ;
        RECT 27.290 313.640 30.710 313.690 ;
        RECT 27.280 313.070 30.720 313.640 ;
        RECT 159.580 313.580 159.910 341.500 ;
        RECT 159.550 313.120 159.950 313.580 ;
        RECT 25.870 304.620 30.170 312.300 ;
        RECT 31.850 312.250 32.570 312.800 ;
        RECT 159.340 312.630 159.920 312.740 ;
        RECT 160.250 312.630 160.580 343.070 ;
        RECT 160.890 317.210 161.220 348.240 ;
        RECT 160.890 312.750 161.210 317.210 ;
        RECT 161.500 313.360 161.830 349.720 ;
        RECT 162.120 313.610 162.450 351.270 ;
        RECT 162.750 314.640 163.080 352.850 ;
        RECT 163.350 314.940 163.680 358.330 ;
        RECT 163.930 315.510 164.260 359.890 ;
        RECT 164.540 316.540 164.870 361.430 ;
        RECT 165.130 317.150 165.460 362.990 ;
        RECT 165.770 317.820 166.100 363.570 ;
        RECT 166.390 318.470 166.720 365.170 ;
        RECT 166.990 319.100 167.320 366.660 ;
        RECT 167.620 319.710 167.950 368.380 ;
        RECT 171.270 367.540 171.680 367.870 ;
        RECT 172.010 367.360 172.250 368.560 ;
        RECT 173.430 368.400 173.780 368.690 ;
        RECT 173.430 368.380 173.630 368.400 ;
        RECT 174.390 368.190 174.700 368.200 ;
        RECT 174.390 367.920 174.710 368.190 ;
        RECT 174.410 367.910 174.700 367.920 ;
        RECT 174.950 367.360 175.260 369.050 ;
        RECT 175.430 367.980 175.750 368.260 ;
        RECT 175.430 367.960 175.790 367.980 ;
        RECT 175.510 367.650 175.790 367.960 ;
        RECT 172.010 366.870 172.250 367.290 ;
        RECT 169.230 366.800 169.470 366.870 ;
        RECT 172.010 366.810 172.480 366.870 ;
        RECT 171.270 365.790 171.680 366.120 ;
        RECT 172.010 365.610 172.250 366.810 ;
        RECT 173.430 366.650 173.780 366.940 ;
        RECT 173.430 366.630 173.630 366.650 ;
        RECT 174.390 366.440 174.700 366.450 ;
        RECT 174.390 366.170 174.710 366.440 ;
        RECT 174.410 366.160 174.700 366.170 ;
        RECT 174.950 365.610 175.260 367.300 ;
        RECT 175.430 366.230 175.750 366.510 ;
        RECT 175.430 366.210 175.790 366.230 ;
        RECT 175.510 365.900 175.790 366.210 ;
        RECT 176.500 365.120 176.790 371.590 ;
        RECT 177.020 369.500 177.310 377.100 ;
        RECT 181.980 376.630 182.590 376.770 ;
        RECT 182.760 376.630 183.010 377.100 ;
        RECT 184.460 377.060 185.190 383.930 ;
        RECT 186.420 379.790 187.140 385.460 ;
        RECT 187.890 386.190 202.180 386.750 ;
        RECT 213.110 386.580 213.640 387.480 ;
        RECT 214.750 387.420 217.120 387.870 ;
        RECT 187.890 386.030 211.240 386.190 ;
        RECT 214.780 386.030 215.730 387.420 ;
        RECT 216.480 387.400 217.060 387.420 ;
        RECT 218.290 386.760 219.010 387.770 ;
        RECT 226.860 386.760 230.770 388.220 ;
        RECT 238.090 387.570 242.220 387.970 ;
        RECT 243.170 387.870 247.060 388.670 ;
        RECT 257.240 388.590 257.610 389.540 ;
        RECT 256.890 388.220 259.360 388.590 ;
        RECT 238.090 387.480 242.230 387.570 ;
        RECT 217.150 386.750 230.770 386.760 ;
        RECT 216.480 386.190 230.770 386.750 ;
        RECT 241.700 386.580 242.230 387.480 ;
        RECT 243.340 387.420 245.710 387.870 ;
        RECT 216.480 386.030 239.830 386.190 ;
        RECT 187.890 385.310 239.830 386.030 ;
        RECT 243.370 385.460 244.320 387.420 ;
        RECT 245.070 387.400 245.650 387.420 ;
        RECT 255.450 386.760 259.360 388.220 ;
        RECT 266.680 387.570 270.810 387.970 ;
        RECT 271.750 387.870 275.640 388.670 ;
        RECT 285.830 388.590 286.200 389.540 ;
        RECT 285.480 388.220 287.950 388.590 ;
        RECT 266.680 387.480 270.820 387.570 ;
        RECT 245.740 386.750 259.360 386.760 ;
        RECT 187.890 381.890 211.240 385.310 ;
        RECT 212.010 384.770 212.580 384.780 ;
        RECT 187.890 381.610 202.180 381.890 ;
        RECT 178.210 376.110 178.710 376.550 ;
        RECT 169.260 364.680 169.500 364.730 ;
        RECT 172.200 364.680 172.510 364.740 ;
        RECT 176.530 364.680 176.820 364.800 ;
        RECT 169.750 363.510 169.990 363.620 ;
        RECT 172.690 363.510 173.000 363.620 ;
        RECT 177.020 363.470 177.310 363.630 ;
        RECT 178.480 363.110 178.670 376.110 ;
        RECT 181.960 374.670 183.140 376.630 ;
        RECT 181.160 373.760 183.140 374.670 ;
        RECT 181.160 373.580 183.010 373.760 ;
        RECT 181.160 372.890 181.890 373.580 ;
        RECT 182.760 363.070 183.010 373.580 ;
        RECT 184.620 366.670 184.790 377.060 ;
        RECT 186.400 373.600 187.120 377.460 ;
        RECT 189.620 376.530 190.590 381.610 ;
        RECT 198.270 380.060 202.180 381.610 ;
        RECT 198.250 379.290 202.200 380.060 ;
        RECT 195.010 378.690 196.480 379.220 ;
        RECT 189.600 376.060 190.610 376.530 ;
        RECT 190.800 376.230 194.750 377.000 ;
        RECT 192.640 376.080 193.080 376.230 ;
        RECT 186.840 372.330 187.180 372.620 ;
        RECT 186.890 372.300 187.150 372.330 ;
        RECT 185.010 368.770 185.270 369.090 ;
        RECT 185.040 366.540 185.230 368.770 ;
        RECT 186.910 366.520 187.120 372.300 ;
        RECT 190.480 371.700 190.740 371.710 ;
        RECT 190.460 371.400 190.760 371.700 ;
        RECT 190.480 371.390 190.740 371.400 ;
        RECT 187.310 370.370 187.650 370.690 ;
        RECT 187.380 366.540 187.570 370.370 ;
        RECT 187.750 368.280 188.040 368.600 ;
        RECT 187.790 366.520 188.000 368.280 ;
        RECT 188.790 367.800 189.130 368.120 ;
        RECT 188.870 366.550 189.050 367.800 ;
        RECT 190.510 363.310 190.710 371.390 ;
        RECT 192.740 366.500 192.970 376.080 ;
        RECT 193.640 372.310 193.920 372.630 ;
        RECT 193.200 371.400 193.480 371.720 ;
        RECT 188.980 363.240 189.170 363.310 ;
        RECT 190.290 363.230 190.710 363.310 ;
        RECT 186.660 362.920 186.850 363.140 ;
        RECT 169.260 362.400 169.500 362.450 ;
        RECT 172.200 362.390 172.510 362.450 ;
        RECT 176.530 362.330 176.820 362.450 ;
        RECT 186.380 362.430 186.850 362.920 ;
        RECT 187.240 362.780 187.610 362.800 ;
        RECT 187.190 362.520 187.610 362.780 ;
        RECT 187.240 362.510 187.610 362.520 ;
        RECT 171.270 361.010 171.680 361.340 ;
        RECT 169.230 360.260 169.470 360.330 ;
        RECT 172.010 360.320 172.250 361.520 ;
        RECT 174.410 360.960 174.700 360.970 ;
        RECT 174.390 360.690 174.710 360.960 ;
        RECT 174.390 360.680 174.700 360.690 ;
        RECT 173.430 360.480 173.630 360.500 ;
        RECT 172.010 360.260 172.480 360.320 ;
        RECT 172.010 359.840 172.250 360.260 ;
        RECT 173.430 360.190 173.780 360.480 ;
        RECT 174.950 359.830 175.260 361.520 ;
        RECT 175.510 360.920 175.790 361.230 ;
        RECT 175.430 360.900 175.790 360.920 ;
        RECT 175.430 360.620 175.750 360.900 ;
        RECT 171.270 359.260 171.680 359.590 ;
        RECT 169.230 358.510 169.470 358.580 ;
        RECT 172.010 358.570 172.250 359.770 ;
        RECT 174.410 359.210 174.700 359.220 ;
        RECT 174.390 358.940 174.710 359.210 ;
        RECT 174.390 358.930 174.700 358.940 ;
        RECT 173.430 358.730 173.630 358.750 ;
        RECT 172.010 358.510 172.480 358.570 ;
        RECT 172.010 358.090 172.250 358.510 ;
        RECT 173.430 358.440 173.780 358.730 ;
        RECT 174.950 358.080 175.260 359.770 ;
        RECT 175.510 359.170 175.790 359.480 ;
        RECT 175.430 359.150 175.790 359.170 ;
        RECT 175.430 358.870 175.750 359.150 ;
        RECT 171.270 357.510 171.680 357.840 ;
        RECT 169.230 356.760 169.470 356.830 ;
        RECT 169.260 355.450 169.500 355.500 ;
        RECT 169.230 355.010 169.470 355.080 ;
        RECT 169.650 353.100 169.890 357.470 ;
        RECT 172.010 356.820 172.250 358.020 ;
        RECT 172.010 356.760 172.480 356.820 ;
        RECT 172.010 356.340 172.250 356.760 ;
        RECT 171.270 355.760 171.680 356.090 ;
        RECT 172.010 355.510 172.250 356.270 ;
        RECT 172.010 355.450 172.510 355.510 ;
        RECT 172.010 355.070 172.250 355.450 ;
        RECT 172.010 355.010 172.480 355.070 ;
        RECT 172.010 354.590 172.250 355.010 ;
        RECT 172.590 353.030 172.900 357.540 ;
        RECT 174.410 357.460 174.700 357.470 ;
        RECT 174.390 357.190 174.710 357.460 ;
        RECT 174.390 357.180 174.700 357.190 ;
        RECT 173.430 356.980 173.630 357.000 ;
        RECT 173.430 356.690 173.780 356.980 ;
        RECT 174.950 356.330 175.260 358.020 ;
        RECT 175.510 357.420 175.790 357.730 ;
        RECT 175.430 357.400 175.790 357.420 ;
        RECT 175.430 357.120 175.750 357.400 ;
        RECT 174.410 355.710 174.700 355.720 ;
        RECT 174.390 355.440 174.710 355.710 ;
        RECT 174.390 355.430 174.700 355.440 ;
        RECT 173.430 355.230 173.630 355.250 ;
        RECT 173.430 354.940 173.780 355.230 ;
        RECT 174.950 354.580 175.260 356.270 ;
        RECT 175.510 355.670 175.790 355.980 ;
        RECT 175.430 355.650 175.790 355.670 ;
        RECT 175.430 355.370 175.750 355.650 ;
        RECT 176.500 355.540 176.790 362.010 ;
        RECT 186.200 361.990 186.520 362.270 ;
        RECT 186.660 362.090 186.850 362.430 ;
        RECT 186.200 361.620 186.520 361.900 ;
        RECT 186.560 361.800 186.850 362.090 ;
        RECT 186.660 361.460 186.850 361.800 ;
        RECT 186.380 360.970 186.850 361.460 ;
        RECT 187.240 361.370 187.610 361.380 ;
        RECT 187.190 361.110 187.610 361.370 ;
        RECT 187.240 361.090 187.610 361.110 ;
        RECT 186.660 360.750 186.850 360.970 ;
        RECT 187.970 360.750 188.200 363.140 ;
        RECT 189.700 362.760 190.040 362.810 ;
        RECT 189.700 362.740 190.260 362.760 ;
        RECT 189.580 362.570 190.260 362.740 ;
        RECT 189.700 362.530 190.260 362.570 ;
        RECT 189.700 362.490 190.040 362.530 ;
        RECT 189.700 361.360 190.040 361.400 ;
        RECT 189.700 361.320 190.260 361.360 ;
        RECT 189.580 361.150 190.260 361.320 ;
        RECT 190.510 361.160 190.710 363.230 ;
        RECT 189.700 361.130 190.260 361.150 ;
        RECT 189.700 361.080 190.040 361.130 ;
        RECT 190.490 361.030 190.710 361.160 ;
        RECT 190.940 362.920 191.190 363.140 ;
        RECT 190.440 360.700 190.770 361.030 ;
        RECT 190.940 360.970 191.580 362.920 ;
        RECT 193.230 361.950 193.450 371.400 ;
        RECT 193.230 361.940 193.510 361.950 ;
        RECT 190.940 360.750 191.190 360.970 ;
        RECT 192.970 360.590 192.980 360.750 ;
        RECT 186.660 359.720 186.850 359.940 ;
        RECT 186.380 359.230 186.850 359.720 ;
        RECT 187.240 359.580 187.610 359.600 ;
        RECT 187.190 359.320 187.610 359.580 ;
        RECT 187.240 359.310 187.610 359.320 ;
        RECT 186.200 358.790 186.520 359.070 ;
        RECT 186.660 358.890 186.850 359.230 ;
        RECT 186.200 358.420 186.520 358.700 ;
        RECT 186.560 358.600 186.850 358.890 ;
        RECT 186.660 358.260 186.850 358.600 ;
        RECT 186.380 357.770 186.850 358.260 ;
        RECT 187.240 358.170 187.610 358.180 ;
        RECT 187.190 357.910 187.610 358.170 ;
        RECT 187.240 357.890 187.610 357.910 ;
        RECT 186.660 357.550 186.850 357.770 ;
        RECT 187.970 357.550 188.200 359.940 ;
        RECT 190.940 359.720 191.190 359.940 ;
        RECT 193.230 359.860 193.450 361.940 ;
        RECT 193.220 359.790 193.450 359.860 ;
        RECT 189.700 359.560 190.040 359.610 ;
        RECT 189.700 359.540 190.260 359.560 ;
        RECT 189.580 359.370 190.260 359.540 ;
        RECT 189.700 359.330 190.260 359.370 ;
        RECT 189.700 359.290 190.040 359.330 ;
        RECT 189.700 358.160 190.040 358.200 ;
        RECT 189.700 358.120 190.260 358.160 ;
        RECT 189.580 357.950 190.260 358.120 ;
        RECT 189.700 357.930 190.260 357.950 ;
        RECT 189.700 357.880 190.040 357.930 ;
        RECT 190.940 357.770 191.580 359.720 ;
        RECT 193.210 359.190 193.410 359.790 ;
        RECT 193.660 359.340 193.890 372.310 ;
        RECT 195.030 366.310 195.450 378.690 ;
        RECT 196.060 366.310 196.480 378.690 ;
        RECT 198.440 376.040 198.880 376.540 ;
        RECT 198.540 369.060 198.770 376.040 ;
        RECT 198.930 372.480 202.160 378.700 ;
        RECT 202.960 370.790 204.240 381.890 ;
        RECT 206.720 377.570 207.000 377.690 ;
        RECT 206.720 377.070 207.050 377.570 ;
        RECT 202.960 370.710 204.260 370.790 ;
        RECT 202.950 370.410 204.260 370.710 ;
        RECT 199.730 369.760 200.030 370.080 ;
        RECT 198.410 369.050 198.770 369.060 ;
        RECT 198.380 368.160 198.770 369.050 ;
        RECT 198.540 366.500 198.770 368.160 ;
        RECT 199.760 366.500 199.990 369.760 ;
        RECT 206.040 369.210 206.470 369.550 ;
        RECT 206.280 366.540 206.470 369.210 ;
        RECT 206.720 366.450 207.000 377.070 ;
        RECT 208.420 372.310 208.680 372.630 ;
        RECT 207.530 371.440 207.790 371.760 ;
        RECT 207.560 367.720 207.750 371.440 ;
        RECT 208.440 367.720 208.660 372.310 ;
        RECT 210.410 369.090 210.750 381.890 ;
        RECT 211.480 380.210 211.870 382.270 ;
        RECT 212.010 381.350 212.630 384.770 ;
        RECT 215.010 381.860 215.730 385.310 ;
        RECT 214.910 381.850 215.730 381.860 ;
        RECT 214.860 381.400 215.730 381.850 ;
        RECT 216.480 384.110 239.830 385.310 ;
        RECT 240.600 384.770 241.170 384.780 ;
        RECT 216.480 381.890 239.960 384.110 ;
        RECT 216.480 381.610 230.770 381.890 ;
        RECT 212.010 381.340 212.580 381.350 ;
        RECT 211.180 379.710 211.870 380.210 ;
        RECT 211.190 379.490 211.870 379.710 ;
        RECT 210.800 378.370 210.960 379.010 ;
        RECT 210.800 377.820 211.070 378.370 ;
        RECT 210.790 377.770 211.070 377.820 ;
        RECT 210.790 377.680 210.960 377.770 ;
        RECT 210.800 375.990 210.960 377.680 ;
        RECT 211.210 377.560 211.400 379.010 ;
        RECT 211.480 378.680 211.870 379.490 ;
        RECT 214.910 379.790 215.730 381.400 ;
        RECT 226.860 380.060 230.770 381.610 ;
        RECT 212.610 378.200 212.920 378.640 ;
        RECT 211.180 377.530 211.400 377.560 ;
        RECT 211.170 377.260 211.420 377.530 ;
        RECT 211.170 377.250 211.410 377.260 ;
        RECT 211.180 377.010 211.410 377.250 ;
        RECT 211.210 375.990 211.370 377.010 ;
        RECT 211.560 376.240 211.800 376.580 ;
        RECT 211.560 376.200 212.120 376.240 ;
        RECT 210.800 373.470 210.960 375.160 ;
        RECT 211.210 374.140 211.370 375.160 ;
        RECT 211.730 374.950 212.120 376.200 ;
        RECT 211.560 374.570 212.120 374.950 ;
        RECT 211.180 373.900 211.410 374.140 ;
        RECT 211.170 373.890 211.410 373.900 ;
        RECT 211.170 373.620 211.420 373.890 ;
        RECT 211.180 373.590 211.400 373.620 ;
        RECT 210.790 373.380 210.960 373.470 ;
        RECT 210.790 373.360 211.070 373.380 ;
        RECT 211.210 373.360 211.400 373.590 ;
        RECT 210.790 373.330 211.400 373.360 ;
        RECT 210.800 372.990 211.400 373.330 ;
        RECT 210.800 372.980 211.070 372.990 ;
        RECT 211.080 372.980 211.400 372.990 ;
        RECT 210.800 372.780 211.400 372.980 ;
        RECT 210.800 372.140 210.960 372.780 ;
        RECT 211.050 372.140 211.400 372.780 ;
        RECT 211.050 371.790 211.350 372.140 ;
        RECT 211.040 371.650 211.350 371.790 ;
        RECT 211.050 369.960 211.350 371.650 ;
        RECT 211.460 371.530 211.650 372.980 ;
        RECT 211.730 372.650 212.120 374.570 ;
        RECT 212.610 372.610 212.920 372.950 ;
        RECT 212.610 372.510 213.170 372.610 ;
        RECT 212.860 372.220 213.170 372.510 ;
        RECT 211.430 371.500 211.650 371.530 ;
        RECT 212.620 372.170 213.170 372.220 ;
        RECT 211.420 371.230 211.670 371.500 ;
        RECT 212.620 371.430 212.880 372.170 ;
        RECT 211.420 371.220 211.660 371.230 ;
        RECT 211.430 370.980 211.660 371.220 ;
        RECT 211.460 369.960 211.620 370.980 ;
        RECT 211.810 370.170 212.050 370.550 ;
        RECT 211.080 369.130 211.350 369.960 ;
        RECT 210.360 369.010 210.750 369.090 ;
        RECT 210.350 368.240 210.750 369.010 ;
        RECT 210.360 368.170 210.750 368.240 ;
        RECT 207.390 367.030 208.070 367.720 ;
        RECT 208.430 367.030 209.110 367.720 ;
        RECT 210.410 366.390 210.750 368.170 ;
        RECT 211.050 367.610 211.350 369.130 ;
        RECT 211.460 368.110 211.620 369.130 ;
        RECT 211.810 368.540 212.050 368.920 ;
        RECT 211.430 367.870 211.660 368.110 ;
        RECT 211.420 367.860 211.660 367.870 ;
        RECT 211.420 367.610 211.670 367.860 ;
        RECT 211.050 367.440 211.760 367.610 ;
        RECT 211.040 367.300 211.760 367.440 ;
        RECT 211.050 367.110 211.760 367.300 ;
        RECT 211.050 366.460 211.350 367.110 ;
        RECT 211.050 366.110 211.210 366.460 ;
        RECT 211.460 366.110 211.650 367.110 ;
        RECT 212.620 366.920 212.880 367.560 ;
        RECT 212.620 366.770 213.170 366.920 ;
        RECT 212.860 366.480 213.170 366.770 ;
        RECT 193.220 359.160 193.450 359.190 ;
        RECT 193.230 358.750 193.450 359.160 ;
        RECT 193.230 358.740 193.510 358.750 ;
        RECT 190.940 357.550 191.190 357.770 ;
        RECT 176.500 355.450 176.820 355.540 ;
        RECT 176.500 355.010 176.790 355.450 ;
        RECT 177.020 353.050 177.310 357.520 ;
        RECT 178.480 353.560 178.670 357.460 ;
        RECT 179.790 353.660 180.020 357.500 ;
        RECT 182.760 353.670 183.010 357.520 ;
        RECT 193.230 357.330 193.450 358.740 ;
        RECT 196.710 358.070 197.100 359.930 ;
        RECT 200.740 358.140 201.130 360.000 ;
        RECT 188.980 357.260 189.170 357.310 ;
        RECT 190.290 357.260 190.520 357.330 ;
        RECT 193.230 357.260 193.510 357.330 ;
        RECT 193.230 355.960 193.450 357.260 ;
        RECT 193.230 355.870 193.580 355.960 ;
        RECT 193.230 355.650 193.740 355.870 ;
        RECT 201.620 355.120 202.000 361.620 ;
        RECT 203.370 357.370 203.530 358.070 ;
        RECT 203.370 356.820 203.640 357.370 ;
        RECT 203.360 356.770 203.640 356.820 ;
        RECT 203.780 357.030 203.970 358.020 ;
        RECT 204.180 357.340 204.340 358.070 ;
        RECT 205.020 357.480 205.340 357.800 ;
        RECT 214.910 357.670 215.280 379.790 ;
        RECT 226.840 379.290 230.790 380.060 ;
        RECT 215.560 378.550 215.720 378.600 ;
        RECT 215.970 378.540 216.160 378.600 ;
        RECT 215.700 377.950 216.160 378.380 ;
        RECT 217.840 378.310 218.050 378.600 ;
        RECT 217.730 378.020 218.050 378.310 ;
        RECT 215.720 372.600 216.090 377.950 ;
        RECT 216.830 376.400 217.150 376.720 ;
        RECT 217.840 376.320 218.050 378.020 ;
        RECT 218.310 377.750 218.500 378.600 ;
        RECT 218.200 377.460 218.500 377.750 ;
        RECT 217.730 376.030 218.050 376.320 ;
        RECT 216.200 375.780 216.460 375.840 ;
        RECT 217.840 375.810 218.050 376.030 ;
        RECT 216.200 375.520 216.560 375.780 ;
        RECT 216.320 375.360 216.560 375.520 ;
        RECT 218.310 375.430 218.500 377.460 ;
        RECT 218.720 376.140 218.930 378.600 ;
        RECT 219.800 377.000 219.980 378.600 ;
        RECT 219.390 376.230 223.340 377.000 ;
        RECT 218.600 375.630 218.930 376.140 ;
        RECT 217.860 375.250 218.050 375.300 ;
        RECT 216.820 374.710 217.140 375.030 ;
        RECT 217.740 374.960 218.050 375.250 ;
        RECT 218.200 375.140 218.500 375.430 ;
        RECT 216.470 373.240 216.920 373.670 ;
        RECT 217.860 373.340 218.050 374.960 ;
        RECT 218.310 373.850 218.500 375.140 ;
        RECT 218.190 373.560 218.500 373.850 ;
        RECT 215.560 372.550 216.160 372.600 ;
        RECT 215.690 366.520 216.090 372.550 ;
        RECT 216.220 372.510 216.410 372.570 ;
        RECT 216.490 370.100 216.860 373.240 ;
        RECT 217.540 373.050 217.550 373.060 ;
        RECT 217.760 373.050 218.050 373.340 ;
        RECT 217.850 372.550 218.080 373.050 ;
        RECT 218.310 372.550 218.500 373.560 ;
        RECT 218.720 372.550 218.930 375.630 ;
        RECT 219.800 374.070 219.980 376.230 ;
        RECT 223.670 375.740 223.900 378.600 ;
        RECT 223.570 375.450 223.900 375.740 ;
        RECT 219.740 373.730 220.030 374.070 ;
        RECT 219.800 372.550 219.980 373.730 ;
        RECT 217.320 370.940 217.640 371.260 ;
        RECT 219.830 370.620 220.390 371.270 ;
        RECT 220.780 371.110 221.340 371.690 ;
        RECT 221.860 371.570 222.420 372.160 ;
        RECT 216.460 369.780 216.860 370.100 ;
        RECT 216.490 369.500 216.860 369.780 ;
        RECT 216.460 369.180 216.860 369.500 ;
        RECT 216.220 366.520 216.410 366.580 ;
        RECT 206.260 357.390 206.420 357.440 ;
        RECT 206.670 357.390 206.860 357.440 ;
        RECT 207.070 357.400 207.230 357.440 ;
        RECT 204.140 357.320 204.340 357.340 ;
        RECT 204.130 357.080 204.360 357.320 ;
        RECT 204.130 357.030 204.340 357.080 ;
        RECT 203.780 356.910 203.950 357.030 ;
        RECT 203.360 356.680 203.530 356.770 ;
        RECT 203.370 356.170 203.530 356.680 ;
        RECT 203.780 356.170 203.940 356.910 ;
        RECT 204.180 356.170 204.340 357.030 ;
        RECT 205.020 356.930 205.340 357.250 ;
        RECT 209.010 356.280 209.250 357.670 ;
        RECT 211.190 357.340 211.570 357.670 ;
        RECT 203.370 355.390 203.530 355.900 ;
        RECT 203.360 355.300 203.530 355.390 ;
        RECT 203.360 355.250 203.640 355.300 ;
        RECT 178.460 353.060 178.670 353.560 ;
        RECT 179.770 353.250 180.020 353.660 ;
        RECT 182.740 353.250 183.010 353.670 ;
        RECT 184.520 353.820 184.800 354.930 ;
        RECT 185.050 354.240 185.240 354.840 ;
        RECT 187.050 354.400 187.440 354.420 ;
        RECT 187.040 354.310 187.440 354.400 ;
        RECT 186.890 354.300 187.440 354.310 ;
        RECT 185.050 354.050 186.650 354.240 ;
        RECT 184.520 353.540 186.240 353.820 ;
        RECT 186.040 353.310 186.240 353.540 ;
        RECT 178.460 352.930 178.650 353.060 ;
        RECT 179.770 352.820 180.000 353.250 ;
        RECT 182.740 352.880 182.990 353.250 ;
        RECT 186.050 353.010 186.210 353.310 ;
        RECT 186.460 352.930 186.650 354.050 ;
        RECT 186.860 354.060 187.440 354.300 ;
        RECT 186.860 354.040 187.430 354.060 ;
        RECT 186.860 354.030 187.050 354.040 ;
        RECT 186.860 353.190 187.030 354.030 ;
        RECT 191.530 353.970 191.760 354.880 ;
        RECT 192.750 354.000 192.980 354.880 ;
        RECT 191.010 353.900 191.760 353.970 ;
        RECT 190.980 353.740 191.760 353.900 ;
        RECT 192.730 353.940 192.980 354.000 ;
        RECT 196.060 354.070 196.480 355.070 ;
        RECT 190.980 353.290 191.390 353.740 ;
        RECT 186.860 352.920 187.020 353.190 ;
        RECT 188.960 352.770 189.150 352.840 ;
        RECT 190.270 352.760 190.500 352.840 ;
        RECT 190.980 352.800 191.360 353.290 ;
        RECT 192.730 352.940 192.970 353.940 ;
        RECT 196.060 353.890 196.490 354.070 ;
        RECT 196.060 353.500 196.500 353.890 ;
        RECT 198.540 353.680 198.770 354.880 ;
        RECT 196.090 353.290 196.500 353.500 ;
        RECT 196.090 352.780 196.490 353.290 ;
        RECT 198.530 352.940 198.770 353.680 ;
        RECT 199.760 353.990 199.990 354.880 ;
        RECT 203.370 354.700 203.640 355.250 ;
        RECT 203.780 355.160 203.940 355.900 ;
        RECT 203.780 355.040 203.950 355.160 ;
        RECT 204.180 355.040 204.340 355.900 ;
        RECT 209.000 355.620 209.270 356.280 ;
        RECT 212.940 356.260 213.180 357.670 ;
        RECT 203.370 354.130 203.530 354.700 ;
        RECT 199.760 353.610 200.520 353.990 ;
        RECT 200.140 353.150 200.520 353.610 ;
        RECT 203.370 353.580 203.640 354.130 ;
        RECT 203.360 353.530 203.640 353.580 ;
        RECT 203.780 353.790 203.970 355.040 ;
        RECT 204.130 354.990 204.340 355.040 ;
        RECT 204.130 354.750 204.360 354.990 ;
        RECT 205.020 354.820 205.340 355.140 ;
        RECT 204.140 354.730 204.340 354.750 ;
        RECT 204.180 354.100 204.340 354.730 ;
        RECT 205.020 354.240 205.340 354.590 ;
        RECT 204.140 354.080 204.340 354.100 ;
        RECT 204.130 353.840 204.360 354.080 ;
        RECT 205.020 353.860 205.340 354.010 ;
        RECT 206.280 353.860 206.470 354.840 ;
        RECT 206.720 354.550 207.000 354.930 ;
        RECT 206.670 354.530 207.000 354.550 ;
        RECT 206.640 354.510 207.000 354.530 ;
        RECT 206.640 354.320 207.080 354.510 ;
        RECT 206.640 354.300 207.000 354.320 ;
        RECT 206.670 354.260 207.000 354.300 ;
        RECT 204.130 353.790 204.340 353.840 ;
        RECT 203.780 353.670 203.950 353.790 ;
        RECT 203.360 353.440 203.530 353.530 ;
        RECT 203.370 352.930 203.530 353.440 ;
        RECT 203.780 352.930 203.940 353.670 ;
        RECT 204.180 352.930 204.340 353.790 ;
        RECT 204.450 353.490 204.730 353.810 ;
        RECT 204.880 353.670 206.470 353.860 ;
        RECT 204.480 353.010 204.640 353.490 ;
        RECT 204.880 353.340 205.070 353.670 ;
        RECT 206.720 353.480 207.000 354.260 ;
        RECT 205.330 353.470 207.000 353.480 ;
        RECT 204.850 353.230 205.070 353.340 ;
        RECT 204.850 352.930 205.040 353.230 ;
        RECT 205.290 353.200 207.000 353.470 ;
        RECT 205.290 353.010 205.450 353.200 ;
        RECT 209.010 353.090 209.250 355.620 ;
        RECT 212.930 355.600 213.190 356.260 ;
        RECT 208.740 353.030 209.250 353.090 ;
        RECT 208.740 352.950 209.260 353.030 ;
        RECT 212.940 352.990 213.180 355.600 ;
        RECT 214.910 354.490 215.620 357.670 ;
        RECT 214.880 354.030 215.620 354.490 ;
        RECT 214.910 353.990 215.620 354.030 ;
        RECT 215.220 352.990 215.620 353.990 ;
        RECT 215.720 353.900 216.090 366.520 ;
        RECT 215.690 353.440 216.130 353.900 ;
        RECT 215.720 353.390 216.090 353.440 ;
        RECT 208.730 352.800 209.260 352.950 ;
        RECT 209.300 352.940 209.490 352.990 ;
        RECT 209.700 352.940 209.860 352.990 ;
        RECT 211.640 352.900 211.880 352.990 ;
        RECT 186.640 352.450 186.830 352.670 ;
        RECT 169.260 352.270 169.500 352.320 ;
        RECT 172.200 352.260 172.510 352.320 ;
        RECT 176.530 352.200 176.820 352.320 ;
        RECT 186.360 351.960 186.830 352.450 ;
        RECT 187.220 352.310 187.590 352.330 ;
        RECT 187.170 352.050 187.590 352.310 ;
        RECT 187.220 352.040 187.590 352.050 ;
        RECT 171.270 350.880 171.680 351.210 ;
        RECT 169.230 350.130 169.470 350.200 ;
        RECT 172.010 350.190 172.250 351.390 ;
        RECT 174.410 350.830 174.700 350.840 ;
        RECT 174.390 350.560 174.710 350.830 ;
        RECT 174.390 350.550 174.700 350.560 ;
        RECT 173.430 350.350 173.630 350.370 ;
        RECT 172.010 350.130 172.480 350.190 ;
        RECT 172.010 349.710 172.250 350.130 ;
        RECT 173.430 350.060 173.780 350.350 ;
        RECT 174.950 349.700 175.260 351.390 ;
        RECT 175.510 350.790 175.790 351.100 ;
        RECT 175.430 350.770 175.790 350.790 ;
        RECT 175.430 350.490 175.750 350.770 ;
        RECT 171.270 349.130 171.680 349.460 ;
        RECT 169.230 348.380 169.470 348.450 ;
        RECT 172.010 348.440 172.250 349.640 ;
        RECT 174.410 349.080 174.700 349.090 ;
        RECT 174.390 348.810 174.710 349.080 ;
        RECT 174.390 348.800 174.700 348.810 ;
        RECT 173.430 348.600 173.630 348.620 ;
        RECT 172.010 348.380 172.480 348.440 ;
        RECT 172.010 347.960 172.250 348.380 ;
        RECT 173.430 348.310 173.780 348.600 ;
        RECT 174.950 347.950 175.260 349.640 ;
        RECT 175.510 349.040 175.790 349.350 ;
        RECT 175.430 349.020 175.790 349.040 ;
        RECT 175.430 348.740 175.750 349.020 ;
        RECT 171.270 347.380 171.680 347.710 ;
        RECT 169.230 346.630 169.470 346.700 ;
        RECT 169.650 346.480 169.890 347.340 ;
        RECT 172.010 346.690 172.250 347.890 ;
        RECT 172.010 346.630 172.480 346.690 ;
        RECT 169.260 345.320 169.500 345.370 ;
        RECT 169.230 344.880 169.470 344.950 ;
        RECT 169.650 343.570 169.990 346.480 ;
        RECT 172.010 346.210 172.250 346.630 ;
        RECT 172.590 346.480 172.900 347.410 ;
        RECT 174.410 347.330 174.700 347.340 ;
        RECT 174.390 347.060 174.710 347.330 ;
        RECT 174.390 347.050 174.700 347.060 ;
        RECT 173.430 346.850 173.630 346.870 ;
        RECT 173.430 346.560 173.780 346.850 ;
        RECT 171.270 345.630 171.680 345.960 ;
        RECT 172.010 345.380 172.250 346.140 ;
        RECT 172.010 345.320 172.510 345.380 ;
        RECT 172.010 344.940 172.250 345.320 ;
        RECT 172.010 344.880 172.480 344.940 ;
        RECT 172.010 344.460 172.250 344.880 ;
        RECT 172.590 343.570 173.000 346.480 ;
        RECT 174.950 346.200 175.260 347.890 ;
        RECT 175.510 347.290 175.790 347.600 ;
        RECT 175.430 347.270 175.790 347.290 ;
        RECT 175.430 346.990 175.750 347.270 ;
        RECT 174.410 345.580 174.700 345.590 ;
        RECT 174.390 345.310 174.710 345.580 ;
        RECT 174.390 345.300 174.700 345.310 ;
        RECT 173.430 345.100 173.630 345.120 ;
        RECT 173.430 344.810 173.780 345.100 ;
        RECT 174.950 344.450 175.260 346.140 ;
        RECT 175.510 345.540 175.790 345.850 ;
        RECT 175.430 345.520 175.790 345.540 ;
        RECT 175.430 345.240 175.750 345.520 ;
        RECT 176.500 345.410 176.790 351.880 ;
        RECT 186.180 351.520 186.500 351.800 ;
        RECT 186.640 351.620 186.830 351.960 ;
        RECT 186.180 351.150 186.500 351.430 ;
        RECT 186.540 351.330 186.830 351.620 ;
        RECT 186.640 350.990 186.830 351.330 ;
        RECT 186.360 350.500 186.830 350.990 ;
        RECT 187.220 350.900 187.590 350.910 ;
        RECT 187.170 350.640 187.590 350.900 ;
        RECT 187.220 350.620 187.590 350.640 ;
        RECT 186.640 350.280 186.830 350.500 ;
        RECT 187.950 350.280 188.180 352.670 ;
        RECT 190.920 352.450 191.170 352.670 ;
        RECT 189.680 352.290 190.020 352.340 ;
        RECT 189.680 352.270 190.240 352.290 ;
        RECT 189.560 352.100 190.240 352.270 ;
        RECT 189.680 352.060 190.240 352.100 ;
        RECT 189.680 352.020 190.020 352.060 ;
        RECT 189.680 350.890 190.020 350.930 ;
        RECT 189.680 350.850 190.240 350.890 ;
        RECT 189.560 350.680 190.240 350.850 ;
        RECT 189.680 350.660 190.240 350.680 ;
        RECT 189.680 350.610 190.020 350.660 ;
        RECT 190.920 350.500 191.560 352.450 ;
        RECT 193.240 351.470 193.490 351.480 ;
        RECT 190.920 350.280 191.170 350.500 ;
        RECT 186.640 349.250 186.830 349.470 ;
        RECT 186.360 348.760 186.830 349.250 ;
        RECT 187.220 349.110 187.590 349.130 ;
        RECT 187.170 348.850 187.590 349.110 ;
        RECT 187.220 348.840 187.590 348.850 ;
        RECT 186.180 348.320 186.500 348.600 ;
        RECT 186.640 348.420 186.830 348.760 ;
        RECT 186.180 347.950 186.500 348.230 ;
        RECT 186.540 348.130 186.830 348.420 ;
        RECT 186.640 347.790 186.830 348.130 ;
        RECT 176.500 345.320 176.820 345.410 ;
        RECT 176.500 344.880 176.790 345.320 ;
        RECT 177.020 343.570 177.310 347.390 ;
        RECT 169.750 343.330 169.990 343.570 ;
        RECT 172.690 343.300 173.000 343.570 ;
        RECT 178.480 343.300 178.670 347.390 ;
        RECT 179.790 346.350 180.020 347.430 ;
        RECT 179.700 345.870 180.030 346.350 ;
        RECT 179.790 343.260 180.020 345.870 ;
        RECT 182.760 343.470 183.010 347.450 ;
        RECT 186.080 343.410 186.240 347.460 ;
        RECT 186.360 347.300 186.830 347.790 ;
        RECT 187.220 347.700 187.590 347.710 ;
        RECT 187.170 347.440 187.590 347.700 ;
        RECT 187.220 347.420 187.590 347.440 ;
        RECT 186.640 347.080 186.830 347.300 ;
        RECT 187.950 347.080 188.180 349.470 ;
        RECT 190.920 349.250 191.170 349.470 ;
        RECT 189.680 349.090 190.020 349.140 ;
        RECT 189.680 349.070 190.240 349.090 ;
        RECT 189.560 348.900 190.240 349.070 ;
        RECT 189.680 348.860 190.240 348.900 ;
        RECT 189.680 348.820 190.020 348.860 ;
        RECT 189.680 347.690 190.020 347.730 ;
        RECT 189.680 347.650 190.240 347.690 ;
        RECT 188.830 346.840 189.070 347.540 ;
        RECT 189.560 347.480 190.240 347.650 ;
        RECT 189.680 347.460 190.240 347.480 ;
        RECT 189.680 347.410 190.020 347.460 ;
        RECT 190.920 347.300 191.560 349.250 ;
        RECT 197.310 349.190 197.700 351.050 ;
        RECT 201.340 349.260 201.730 351.120 ;
        RECT 193.240 348.270 193.490 348.280 ;
        RECT 190.920 347.080 191.390 347.300 ;
        RECT 188.830 346.790 189.150 346.840 ;
        RECT 190.270 346.790 190.500 346.860 ;
        RECT 188.830 343.820 189.070 346.790 ;
        RECT 188.810 343.570 189.200 343.820 ;
        RECT 169.220 343.210 169.460 343.260 ;
        RECT 172.160 343.200 172.470 343.260 ;
        RECT 176.490 343.140 176.780 343.260 ;
        RECT 186.670 343.180 186.860 343.400 ;
        RECT 171.230 341.820 171.640 342.150 ;
        RECT 169.190 341.070 169.430 341.140 ;
        RECT 171.970 341.130 172.210 342.330 ;
        RECT 174.370 341.770 174.660 341.780 ;
        RECT 174.350 341.500 174.670 341.770 ;
        RECT 174.350 341.490 174.660 341.500 ;
        RECT 173.390 341.290 173.590 341.310 ;
        RECT 171.970 341.070 172.440 341.130 ;
        RECT 171.970 340.650 172.210 341.070 ;
        RECT 173.390 341.000 173.740 341.290 ;
        RECT 174.910 340.640 175.220 342.330 ;
        RECT 175.470 341.730 175.750 342.040 ;
        RECT 175.390 341.710 175.750 341.730 ;
        RECT 175.390 341.430 175.710 341.710 ;
        RECT 171.230 340.070 171.640 340.400 ;
        RECT 169.190 339.320 169.430 339.390 ;
        RECT 171.970 339.380 172.210 340.580 ;
        RECT 174.370 340.020 174.660 340.030 ;
        RECT 174.350 339.750 174.670 340.020 ;
        RECT 174.350 339.740 174.660 339.750 ;
        RECT 173.390 339.540 173.590 339.560 ;
        RECT 171.970 339.320 172.440 339.380 ;
        RECT 171.970 338.900 172.210 339.320 ;
        RECT 173.390 339.250 173.740 339.540 ;
        RECT 174.910 338.890 175.220 340.580 ;
        RECT 175.470 339.980 175.750 340.290 ;
        RECT 175.390 339.960 175.750 339.980 ;
        RECT 175.390 339.680 175.710 339.960 ;
        RECT 171.230 338.320 171.640 338.650 ;
        RECT 169.190 337.570 169.430 337.640 ;
        RECT 171.970 337.630 172.210 338.830 ;
        RECT 174.370 338.270 174.660 338.280 ;
        RECT 174.350 338.000 174.670 338.270 ;
        RECT 174.350 337.990 174.660 338.000 ;
        RECT 173.390 337.790 173.590 337.810 ;
        RECT 171.970 337.570 172.440 337.630 ;
        RECT 169.220 336.260 169.460 336.310 ;
        RECT 169.190 335.820 169.430 335.890 ;
        RECT 169.650 324.940 169.890 337.570 ;
        RECT 171.970 337.150 172.210 337.570 ;
        RECT 171.230 336.570 171.640 336.900 ;
        RECT 171.970 336.320 172.210 337.080 ;
        RECT 172.590 336.490 172.900 337.640 ;
        RECT 173.390 337.500 173.740 337.790 ;
        RECT 174.910 337.140 175.220 338.830 ;
        RECT 175.470 338.230 175.750 338.540 ;
        RECT 175.390 338.210 175.750 338.230 ;
        RECT 175.390 337.930 175.710 338.210 ;
        RECT 174.370 336.520 174.660 336.530 ;
        RECT 171.970 336.260 172.470 336.320 ;
        RECT 171.970 335.880 172.210 336.260 ;
        RECT 172.550 336.160 172.920 336.490 ;
        RECT 174.350 336.250 174.670 336.520 ;
        RECT 174.350 336.240 174.660 336.250 ;
        RECT 171.970 335.820 172.440 335.880 ;
        RECT 171.970 335.400 172.210 335.820 ;
        RECT 172.590 334.950 172.900 336.160 ;
        RECT 173.390 336.040 173.590 336.060 ;
        RECT 173.390 335.750 173.740 336.040 ;
        RECT 174.910 335.390 175.220 337.080 ;
        RECT 175.470 336.480 175.750 336.790 ;
        RECT 175.390 336.460 175.750 336.480 ;
        RECT 175.390 336.180 175.710 336.460 ;
        RECT 176.460 336.350 176.750 342.820 ;
        RECT 186.390 342.690 186.860 343.180 ;
        RECT 187.250 343.040 187.620 343.060 ;
        RECT 187.200 342.780 187.620 343.040 ;
        RECT 187.250 342.770 187.620 342.780 ;
        RECT 184.110 342.140 184.430 342.480 ;
        RECT 186.210 342.250 186.530 342.530 ;
        RECT 186.670 342.350 186.860 342.690 ;
        RECT 177.020 337.000 177.310 337.620 ;
        RECT 177.520 337.020 177.860 337.340 ;
        RECT 176.990 336.650 177.340 337.000 ;
        RECT 176.460 336.260 176.780 336.350 ;
        RECT 176.460 336.190 176.750 336.260 ;
        RECT 177.020 336.190 177.310 336.650 ;
        RECT 177.520 336.410 177.770 337.020 ;
        RECT 178.480 336.430 178.670 337.630 ;
        RECT 182.760 336.960 183.010 337.690 ;
        RECT 184.190 337.380 184.400 342.140 ;
        RECT 186.210 341.880 186.530 342.160 ;
        RECT 186.570 342.060 186.860 342.350 ;
        RECT 186.670 341.720 186.860 342.060 ;
        RECT 186.390 341.230 186.860 341.720 ;
        RECT 187.250 341.630 187.620 341.640 ;
        RECT 187.200 341.370 187.620 341.630 ;
        RECT 187.250 341.350 187.620 341.370 ;
        RECT 186.670 341.010 186.860 341.230 ;
        RECT 187.980 341.010 188.210 343.400 ;
        RECT 188.950 343.320 189.200 343.570 ;
        RECT 190.300 343.490 190.530 343.570 ;
        RECT 191.010 343.400 191.390 347.080 ;
        RECT 192.760 343.800 193.000 347.540 ;
        RECT 193.240 346.790 193.490 346.860 ;
        RECT 192.760 343.530 193.230 343.800 ;
        RECT 190.950 343.190 191.390 343.400 ;
        RECT 192.960 343.300 193.230 343.530 ;
        RECT 190.950 343.180 191.200 343.190 ;
        RECT 189.710 343.020 190.050 343.070 ;
        RECT 189.710 343.000 190.270 343.020 ;
        RECT 189.590 342.830 190.270 343.000 ;
        RECT 189.710 342.790 190.270 342.830 ;
        RECT 189.710 342.750 190.050 342.790 ;
        RECT 189.710 341.620 190.050 341.660 ;
        RECT 189.710 341.580 190.270 341.620 ;
        RECT 189.590 341.410 190.270 341.580 ;
        RECT 189.710 341.390 190.270 341.410 ;
        RECT 189.710 341.340 190.050 341.390 ;
        RECT 190.950 341.230 191.590 343.180 ;
        RECT 195.040 343.170 195.440 347.700 ;
        RECT 198.560 345.030 198.800 347.540 ;
        RECT 202.220 346.280 202.600 352.780 ;
        RECT 208.890 352.710 209.260 352.800 ;
        RECT 203.370 352.160 203.530 352.670 ;
        RECT 203.360 352.070 203.530 352.160 ;
        RECT 203.360 352.020 203.640 352.070 ;
        RECT 203.370 351.470 203.640 352.020 ;
        RECT 203.780 351.930 203.940 352.670 ;
        RECT 203.780 351.810 203.950 351.930 ;
        RECT 204.180 351.810 204.340 352.670 ;
        RECT 208.890 352.650 209.250 352.710 ;
        RECT 212.930 352.670 213.190 352.990 ;
        RECT 213.820 352.890 214.200 352.990 ;
        RECT 215.220 352.930 215.810 352.990 ;
        RECT 203.370 350.770 203.530 351.470 ;
        RECT 203.780 350.820 203.970 351.810 ;
        RECT 204.130 351.760 204.340 351.810 ;
        RECT 204.130 351.520 204.360 351.760 ;
        RECT 205.020 351.590 205.340 351.910 ;
        RECT 204.140 351.500 204.340 351.520 ;
        RECT 204.180 350.770 204.340 351.500 ;
        RECT 205.020 351.040 205.340 351.360 ;
        RECT 209.010 351.170 209.250 352.650 ;
        RECT 211.190 351.170 211.570 351.770 ;
        RECT 212.940 351.170 213.180 352.670 ;
        RECT 215.220 351.170 215.620 352.930 ;
        RECT 216.490 351.550 216.860 369.180 ;
        RECT 217.360 368.500 217.790 368.600 ;
        RECT 217.320 368.180 217.790 368.500 ;
        RECT 219.850 368.280 220.350 370.620 ;
        RECT 217.360 368.160 217.790 368.180 ;
        RECT 219.650 368.220 220.370 368.280 ;
        RECT 216.460 351.540 216.860 351.550 ;
        RECT 216.450 351.120 216.870 351.540 ;
        RECT 216.490 351.110 216.860 351.120 ;
        RECT 203.970 348.530 204.130 349.230 ;
        RECT 203.970 347.980 204.240 348.530 ;
        RECT 203.960 347.930 204.240 347.980 ;
        RECT 204.380 348.190 204.570 349.180 ;
        RECT 204.780 348.500 204.940 349.230 ;
        RECT 205.620 348.640 205.940 348.960 ;
        RECT 204.740 348.480 204.940 348.500 ;
        RECT 206.860 348.490 207.020 348.560 ;
        RECT 207.270 348.490 207.460 348.560 ;
        RECT 207.670 348.490 207.830 348.560 ;
        RECT 204.730 348.240 204.960 348.480 ;
        RECT 204.730 348.190 204.940 348.240 ;
        RECT 204.380 348.070 204.550 348.190 ;
        RECT 203.960 347.840 204.130 347.930 ;
        RECT 203.970 347.330 204.130 347.840 ;
        RECT 204.380 347.330 204.540 348.070 ;
        RECT 204.780 347.330 204.940 348.190 ;
        RECT 205.620 348.090 205.940 348.410 ;
        RECT 203.970 346.570 204.130 347.080 ;
        RECT 203.960 346.480 204.130 346.570 ;
        RECT 203.960 346.430 204.240 346.480 ;
        RECT 203.970 345.880 204.240 346.430 ;
        RECT 204.380 346.340 204.540 347.080 ;
        RECT 204.380 346.220 204.550 346.340 ;
        RECT 204.780 346.220 204.940 347.080 ;
        RECT 209.730 347.010 209.980 348.830 ;
        RECT 211.790 348.460 212.170 348.830 ;
        RECT 213.740 347.030 214.010 348.830 ;
        RECT 208.890 346.940 209.050 347.000 ;
        RECT 209.300 346.950 209.490 347.010 ;
        RECT 209.700 346.950 209.980 347.010 ;
        RECT 203.970 345.290 204.130 345.880 ;
        RECT 198.560 344.790 199.140 345.030 ;
        RECT 198.900 343.450 199.140 344.790 ;
        RECT 203.970 344.740 204.240 345.290 ;
        RECT 203.960 344.690 204.240 344.740 ;
        RECT 204.380 344.950 204.570 346.220 ;
        RECT 204.730 346.170 204.940 346.220 ;
        RECT 204.730 345.930 204.960 346.170 ;
        RECT 205.620 346.000 205.940 346.320 ;
        RECT 204.740 345.910 204.940 345.930 ;
        RECT 204.780 345.260 204.940 345.910 ;
        RECT 205.620 345.400 205.940 345.770 ;
        RECT 207.240 345.680 207.480 345.710 ;
        RECT 207.240 345.590 207.670 345.680 ;
        RECT 206.860 345.580 207.020 345.590 ;
        RECT 207.240 345.580 207.830 345.590 ;
        RECT 207.240 345.510 207.670 345.580 ;
        RECT 207.240 345.480 207.480 345.510 ;
        RECT 207.270 345.380 207.380 345.480 ;
        RECT 204.740 345.240 204.940 345.260 ;
        RECT 204.730 345.000 204.960 345.240 ;
        RECT 204.730 344.950 204.940 345.000 ;
        RECT 204.380 344.830 204.550 344.950 ;
        RECT 203.960 344.600 204.130 344.690 ;
        RECT 203.970 344.090 204.130 344.600 ;
        RECT 204.380 344.090 204.540 344.830 ;
        RECT 204.780 344.090 204.940 344.950 ;
        RECT 205.620 344.850 205.940 345.170 ;
        RECT 209.730 344.150 209.980 346.950 ;
        RECT 211.640 346.940 211.880 347.020 ;
        RECT 213.740 346.940 214.200 347.030 ;
        RECT 215.570 346.940 215.810 347.010 ;
        RECT 209.500 344.080 209.660 344.150 ;
        RECT 209.730 344.120 210.100 344.150 ;
        RECT 209.710 344.090 210.100 344.120 ;
        RECT 209.700 344.080 210.100 344.090 ;
        RECT 210.310 344.080 210.470 344.150 ;
        RECT 213.740 344.090 214.010 346.940 ;
        RECT 203.970 343.320 204.130 343.830 ;
        RECT 203.960 343.230 204.130 343.320 ;
        RECT 203.960 343.180 204.240 343.230 ;
        RECT 203.970 342.630 204.240 343.180 ;
        RECT 204.380 343.090 204.540 343.830 ;
        RECT 204.380 342.970 204.550 343.090 ;
        RECT 204.780 342.970 204.940 343.830 ;
        RECT 209.700 343.810 210.000 344.080 ;
        RECT 209.710 343.790 209.990 343.810 ;
        RECT 203.970 342.450 204.130 342.630 ;
        RECT 193.270 342.200 193.520 342.210 ;
        RECT 203.970 342.130 204.280 342.450 ;
        RECT 203.970 341.930 204.260 342.130 ;
        RECT 204.380 341.980 204.570 342.970 ;
        RECT 204.730 342.920 204.940 342.970 ;
        RECT 204.730 342.680 204.960 342.920 ;
        RECT 205.620 342.750 205.940 343.070 ;
        RECT 204.740 342.660 204.940 342.680 ;
        RECT 204.780 341.930 204.940 342.660 ;
        RECT 206.860 342.520 207.020 342.590 ;
        RECT 207.270 342.520 207.460 342.590 ;
        RECT 207.670 342.520 207.830 342.590 ;
        RECT 205.620 342.200 205.940 342.520 ;
        RECT 208.730 342.220 208.990 342.440 ;
        RECT 209.730 342.330 209.980 343.790 ;
        RECT 212.020 343.670 212.280 343.990 ;
        RECT 213.720 343.780 214.030 344.090 ;
        RECT 214.430 344.050 214.810 344.150 ;
        RECT 211.930 342.940 212.140 343.570 ;
        RECT 211.930 342.830 212.260 342.940 ;
        RECT 212.000 342.620 212.260 342.830 ;
        RECT 211.790 342.330 212.170 342.610 ;
        RECT 213.740 342.330 214.010 343.780 ;
        RECT 215.820 342.330 216.220 348.830 ;
        RECT 217.370 346.370 217.740 368.160 ;
        RECT 219.650 367.950 220.350 368.220 ;
        RECT 217.850 352.860 218.250 352.990 ;
        RECT 218.930 352.890 219.330 352.990 ;
        RECT 218.250 352.630 218.930 352.850 ;
        RECT 217.850 346.940 218.250 347.060 ;
        RECT 218.930 346.940 219.330 347.060 ;
        RECT 217.330 345.860 217.820 346.370 ;
        RECT 217.370 345.830 217.740 345.860 ;
        RECT 218.460 343.870 218.860 344.150 ;
        RECT 208.630 342.120 208.990 342.220 ;
        RECT 190.950 341.010 191.200 341.230 ;
        RECT 203.500 341.200 203.760 341.520 ;
        RECT 185.450 340.450 185.840 340.700 ;
        RECT 184.730 339.350 185.070 339.690 ;
        RECT 184.770 339.330 184.990 339.350 ;
        RECT 184.160 337.060 184.440 337.380 ;
        RECT 184.770 337.050 184.970 339.330 ;
        RECT 185.230 337.510 185.420 337.870 ;
        RECT 182.730 336.670 183.070 336.960 ;
        RECT 184.730 336.730 185.010 337.050 ;
        RECT 185.190 337.040 185.470 337.510 ;
        RECT 176.450 335.910 177.310 336.190 ;
        RECT 176.370 335.900 177.310 335.910 ;
        RECT 177.470 336.300 177.770 336.410 ;
        RECT 176.370 335.430 176.830 335.900 ;
        RECT 172.540 334.470 172.960 334.950 ;
        RECT 177.470 334.790 177.660 336.300 ;
        RECT 178.420 336.110 178.740 336.430 ;
        RECT 181.100 335.900 181.850 336.090 ;
        RECT 181.350 335.060 181.850 335.900 ;
        RECT 185.660 335.820 185.840 340.450 ;
        RECT 186.670 339.980 186.860 340.200 ;
        RECT 186.390 339.490 186.860 339.980 ;
        RECT 187.250 339.840 187.620 339.860 ;
        RECT 187.200 339.580 187.620 339.840 ;
        RECT 187.250 339.570 187.620 339.580 ;
        RECT 186.210 339.050 186.530 339.330 ;
        RECT 186.670 339.150 186.860 339.490 ;
        RECT 186.210 338.680 186.530 338.960 ;
        RECT 186.570 338.860 186.860 339.150 ;
        RECT 186.670 338.520 186.860 338.860 ;
        RECT 186.390 338.030 186.860 338.520 ;
        RECT 187.250 338.430 187.620 338.440 ;
        RECT 187.200 338.170 187.620 338.430 ;
        RECT 187.250 338.150 187.620 338.170 ;
        RECT 186.670 337.810 186.860 338.030 ;
        RECT 187.980 337.810 188.210 340.200 ;
        RECT 190.950 339.980 191.200 340.200 ;
        RECT 189.710 339.820 190.050 339.870 ;
        RECT 189.710 339.800 190.270 339.820 ;
        RECT 189.590 339.630 190.270 339.800 ;
        RECT 189.710 339.590 190.270 339.630 ;
        RECT 189.710 339.550 190.050 339.590 ;
        RECT 189.710 338.420 190.050 338.460 ;
        RECT 189.710 338.380 190.270 338.420 ;
        RECT 189.590 338.210 190.270 338.380 ;
        RECT 189.710 338.190 190.270 338.210 ;
        RECT 189.710 338.140 190.050 338.190 ;
        RECT 190.950 338.030 191.590 339.980 ;
        RECT 203.030 339.360 203.290 339.680 ;
        RECT 193.270 339.000 193.520 339.010 ;
        RECT 202.530 338.430 202.790 338.750 ;
        RECT 190.950 337.810 191.200 338.030 ;
        RECT 186.980 336.980 187.240 337.010 ;
        RECT 186.960 336.680 187.260 336.980 ;
        RECT 186.980 336.670 187.240 336.680 ;
        RECT 185.660 335.520 186.140 335.820 ;
        RECT 186.990 335.750 187.210 336.670 ;
        RECT 188.950 336.540 189.200 337.770 ;
        RECT 190.300 337.520 190.530 337.590 ;
        RECT 192.960 336.560 193.230 337.790 ;
        RECT 193.270 337.520 193.520 337.590 ;
        RECT 195.780 336.990 196.210 337.390 ;
        RECT 188.940 336.280 189.260 336.540 ;
        RECT 192.960 336.250 193.310 336.560 ;
        RECT 185.740 335.410 186.140 335.520 ;
        RECT 186.930 335.350 187.270 335.750 ;
        RECT 186.990 335.270 187.210 335.350 ;
        RECT 190.940 335.080 191.880 336.010 ;
        RECT 195.820 335.200 196.170 336.990 ;
        RECT 197.640 336.430 197.860 337.750 ;
        RECT 198.900 337.030 199.130 337.750 ;
        RECT 198.900 336.800 202.110 337.030 ;
        RECT 198.900 336.790 199.130 336.800 ;
        RECT 197.350 336.190 197.860 336.430 ;
        RECT 177.030 334.470 177.660 334.790 ;
        RECT 180.860 334.740 181.100 335.060 ;
        RECT 182.100 334.740 182.340 335.060 ;
        RECT 190.670 334.760 190.910 335.080 ;
        RECT 191.910 334.760 192.150 335.080 ;
        RECT 197.350 334.940 197.580 336.190 ;
        RECT 201.880 335.830 202.110 336.800 ;
        RECT 201.830 335.430 202.140 335.830 ;
        RECT 197.240 334.500 197.700 334.940 ;
        RECT 177.030 334.370 177.470 334.470 ;
        RECT 180.860 333.400 181.100 333.720 ;
        RECT 182.100 333.390 182.340 333.710 ;
        RECT 190.670 333.420 190.910 333.740 ;
        RECT 191.910 333.410 192.150 333.730 ;
        RECT 201.880 332.260 202.110 335.430 ;
        RECT 201.750 332.040 202.110 332.260 ;
        RECT 180.460 331.770 180.720 331.970 ;
        RECT 182.480 331.770 182.740 331.970 ;
        RECT 177.330 331.400 177.650 331.720 ;
        RECT 178.420 331.400 178.740 331.720 ;
        RECT 179.520 331.390 179.840 331.710 ;
        RECT 177.240 329.190 177.560 330.940 ;
        RECT 177.880 330.720 178.200 331.040 ;
        RECT 178.970 330.700 179.290 331.020 ;
        RECT 180.080 330.690 180.400 331.010 ;
        RECT 180.460 330.960 180.770 331.770 ;
        RECT 182.430 330.960 182.740 331.770 ;
        RECT 190.270 331.800 190.530 332.000 ;
        RECT 192.290 331.800 192.550 332.000 ;
        RECT 201.550 331.810 202.110 332.040 ;
        RECT 201.550 331.800 202.090 331.810 ;
        RECT 183.360 331.390 183.680 331.710 ;
        RECT 184.460 331.400 184.780 331.720 ;
        RECT 185.550 331.400 185.870 331.720 ;
        RECT 187.140 331.430 187.460 331.750 ;
        RECT 188.230 331.430 188.550 331.750 ;
        RECT 189.330 331.420 189.650 331.740 ;
        RECT 177.880 329.350 178.200 329.670 ;
        RECT 178.970 329.350 179.290 329.670 ;
        RECT 180.070 329.350 180.390 329.670 ;
        RECT 177.120 328.590 177.660 329.190 ;
        RECT 178.420 328.620 178.740 328.940 ;
        RECT 179.520 328.620 179.840 328.940 ;
        RECT 177.320 327.250 177.640 327.570 ;
        RECT 178.420 327.250 178.740 327.570 ;
        RECT 179.520 327.250 179.840 327.570 ;
        RECT 176.750 326.610 177.070 326.930 ;
        RECT 177.880 326.570 178.200 326.890 ;
        RECT 178.970 326.570 179.290 326.890 ;
        RECT 180.070 326.580 180.390 326.900 ;
        RECT 176.760 326.140 177.080 326.460 ;
        RECT 180.460 325.980 180.720 330.960 ;
        RECT 180.860 330.630 181.100 330.950 ;
        RECT 182.100 330.620 182.340 330.940 ;
        RECT 181.100 329.970 181.360 330.430 ;
        RECT 181.840 329.990 182.100 330.430 ;
        RECT 181.090 329.630 181.370 329.970 ;
        RECT 181.830 329.650 182.110 329.990 ;
        RECT 181.100 328.220 181.360 329.630 ;
        RECT 181.840 328.220 182.100 329.650 ;
        RECT 169.250 323.620 169.900 324.940 ;
        RECT 181.100 324.790 182.100 328.220 ;
        RECT 182.480 325.980 182.740 330.960 ;
        RECT 182.800 330.690 183.120 331.010 ;
        RECT 183.910 330.700 184.230 331.020 ;
        RECT 185.000 330.720 185.320 331.040 ;
        RECT 182.810 329.350 183.130 329.670 ;
        RECT 183.910 329.350 184.230 329.670 ;
        RECT 185.000 329.350 185.320 329.670 ;
        RECT 185.610 328.940 185.950 330.960 ;
        RECT 183.360 328.620 183.680 328.940 ;
        RECT 184.460 328.620 184.780 328.940 ;
        RECT 185.560 328.620 185.950 328.940 ;
        RECT 185.610 328.170 185.950 328.620 ;
        RECT 187.040 328.970 187.380 330.950 ;
        RECT 187.690 330.750 188.010 331.070 ;
        RECT 188.780 330.730 189.100 331.050 ;
        RECT 189.890 330.720 190.210 331.040 ;
        RECT 190.270 330.990 190.580 331.800 ;
        RECT 192.240 330.990 192.550 331.800 ;
        RECT 193.170 331.420 193.490 331.740 ;
        RECT 194.270 331.430 194.590 331.750 ;
        RECT 195.360 331.430 195.680 331.750 ;
        RECT 198.910 331.400 199.230 331.720 ;
        RECT 200.010 331.410 200.330 331.730 ;
        RECT 201.100 331.410 201.420 331.730 ;
        RECT 187.690 329.380 188.010 329.700 ;
        RECT 188.780 329.380 189.100 329.700 ;
        RECT 189.880 329.380 190.200 329.700 ;
        RECT 187.040 328.650 187.450 328.970 ;
        RECT 188.230 328.650 188.550 328.970 ;
        RECT 189.330 328.650 189.650 328.970 ;
        RECT 185.550 327.650 186.010 328.170 ;
        RECT 187.040 327.600 187.380 328.650 ;
        RECT 183.360 327.250 183.680 327.570 ;
        RECT 184.460 327.250 184.780 327.570 ;
        RECT 185.560 327.250 185.880 327.570 ;
        RECT 187.040 327.280 187.450 327.600 ;
        RECT 188.230 327.280 188.550 327.600 ;
        RECT 189.330 327.280 189.650 327.600 ;
        RECT 182.810 326.580 183.130 326.900 ;
        RECT 183.910 326.570 184.230 326.890 ;
        RECT 185.000 326.570 185.320 326.890 ;
        RECT 186.130 326.610 186.450 326.930 ;
        RECT 186.560 326.640 186.880 326.960 ;
        RECT 186.950 326.760 187.470 327.280 ;
        RECT 187.690 326.600 188.010 326.920 ;
        RECT 188.780 326.600 189.100 326.920 ;
        RECT 189.880 326.610 190.200 326.930 ;
        RECT 186.120 326.140 186.440 326.460 ;
        RECT 186.570 326.170 186.890 326.490 ;
        RECT 190.270 326.010 190.530 330.990 ;
        RECT 190.670 330.650 190.910 330.970 ;
        RECT 191.910 330.650 192.150 330.970 ;
        RECT 190.910 329.970 191.170 330.460 ;
        RECT 190.900 329.630 191.180 329.970 ;
        RECT 190.910 328.450 191.170 329.630 ;
        RECT 191.650 328.450 191.910 330.460 ;
        RECT 190.910 324.850 191.910 328.450 ;
        RECT 192.290 326.010 192.550 330.990 ;
        RECT 192.610 330.720 192.930 331.040 ;
        RECT 193.720 330.730 194.040 331.050 ;
        RECT 194.810 330.750 195.130 331.070 ;
        RECT 192.620 329.380 192.940 329.700 ;
        RECT 193.720 329.380 194.040 329.700 ;
        RECT 194.810 329.380 195.130 329.700 ;
        RECT 195.460 328.970 195.730 330.990 ;
        RECT 198.350 330.700 198.670 331.020 ;
        RECT 199.460 330.710 199.780 331.030 ;
        RECT 200.550 330.730 200.870 331.050 ;
        RECT 202.530 330.590 202.780 338.430 ;
        RECT 203.030 331.490 203.280 339.360 ;
        RECT 203.510 332.400 203.760 341.200 ;
        RECT 204.010 333.290 204.260 341.930 ;
        RECT 208.630 341.430 208.840 342.120 ;
        RECT 208.630 341.110 208.970 341.430 ;
        RECT 208.630 341.070 208.840 341.110 ;
        RECT 212.000 340.960 212.260 341.060 ;
        RECT 211.910 340.740 212.260 340.960 ;
        RECT 211.910 339.880 212.070 340.740 ;
        RECT 211.870 339.560 212.130 339.880 ;
        RECT 211.910 339.460 212.070 339.560 ;
        RECT 208.680 339.120 209.000 339.440 ;
        RECT 208.730 338.160 209.050 338.480 ;
        RECT 214.430 338.100 214.810 338.200 ;
        RECT 219.850 334.790 220.350 367.950 ;
        RECT 220.780 344.150 221.280 371.110 ;
        RECT 221.910 357.670 222.410 371.570 ;
        RECT 222.700 366.520 222.930 372.570 ;
        RECT 223.040 372.190 223.620 372.750 ;
        RECT 223.670 372.550 223.900 375.450 ;
        RECT 225.960 374.310 226.380 378.600 ;
        RECT 227.520 378.250 230.750 378.700 ;
        RECT 227.520 377.460 230.830 378.250 ;
        RECT 225.800 374.290 226.400 374.310 ;
        RECT 225.640 374.250 226.400 374.290 ;
        RECT 225.640 373.990 226.380 374.250 ;
        RECT 225.960 372.570 226.380 373.990 ;
        RECT 227.520 373.590 230.750 377.460 ;
        RECT 227.520 372.800 230.830 373.590 ;
        RECT 221.560 352.990 222.410 357.670 ;
        RECT 223.040 352.990 223.540 372.190 ;
        RECT 223.920 371.600 224.150 372.570 ;
        RECT 225.960 372.550 226.630 372.570 ;
        RECT 223.910 371.350 224.150 371.600 ;
        RECT 224.580 371.350 224.900 371.670 ;
        RECT 223.920 369.710 224.150 371.350 ;
        RECT 223.820 369.420 224.150 369.710 ;
        RECT 223.920 366.520 224.150 369.420 ;
        RECT 224.610 367.660 224.930 367.980 ;
        RECT 226.210 366.530 226.630 372.550 ;
        RECT 227.520 372.480 230.750 372.800 ;
        RECT 231.900 370.590 233.180 381.890 ;
        RECT 239.770 380.210 239.960 381.890 ;
        RECT 240.600 381.350 241.220 384.770 ;
        RECT 240.600 381.340 241.170 381.350 ;
        RECT 239.770 379.490 240.330 380.210 ;
        RECT 243.600 379.790 244.320 385.460 ;
        RECT 245.070 386.190 259.360 386.750 ;
        RECT 270.290 386.580 270.820 387.480 ;
        RECT 271.930 387.420 274.300 387.870 ;
        RECT 245.070 381.890 268.420 386.190 ;
        RECT 271.960 385.460 272.910 387.420 ;
        RECT 273.660 387.400 274.240 387.420 ;
        RECT 284.040 386.760 287.950 388.220 ;
        RECT 295.270 387.570 299.400 387.970 ;
        RECT 300.340 387.870 304.230 388.670 ;
        RECT 314.420 388.590 314.790 389.540 ;
        RECT 314.070 388.220 316.540 388.590 ;
        RECT 295.270 387.480 299.410 387.570 ;
        RECT 274.330 386.750 287.950 386.760 ;
        RECT 269.190 384.770 269.760 384.780 ;
        RECT 245.070 381.610 259.360 381.890 ;
        RECT 255.450 380.060 259.360 381.610 ;
        RECT 269.190 381.350 269.810 384.770 ;
        RECT 269.190 381.340 269.760 381.350 ;
        RECT 236.450 376.090 236.640 376.100 ;
        RECT 239.770 376.090 239.960 379.490 ;
        RECT 255.430 379.290 259.380 380.060 ;
        RECT 268.360 379.710 268.920 380.210 ;
        RECT 272.190 379.790 272.910 385.460 ;
        RECT 273.660 386.190 287.950 386.750 ;
        RECT 298.880 386.580 299.410 387.480 ;
        RECT 300.520 387.420 302.890 387.870 ;
        RECT 273.660 381.890 297.010 386.190 ;
        RECT 300.550 385.460 301.500 387.420 ;
        RECT 302.250 387.400 302.830 387.420 ;
        RECT 312.630 386.760 316.540 388.220 ;
        RECT 323.860 387.570 327.990 387.970 ;
        RECT 328.940 387.870 332.830 388.670 ;
        RECT 343.010 388.590 343.380 389.540 ;
        RECT 342.660 388.220 345.130 388.590 ;
        RECT 323.860 387.480 328.000 387.570 ;
        RECT 302.920 386.750 316.540 386.760 ;
        RECT 297.780 384.770 298.350 384.780 ;
        RECT 273.660 381.610 287.950 381.890 ;
        RECT 284.040 380.060 287.950 381.610 ;
        RECT 297.780 381.350 298.400 384.770 ;
        RECT 297.780 381.340 298.350 381.350 ;
        RECT 268.370 379.490 268.920 379.710 ;
        RECT 284.020 379.290 287.970 380.060 ;
        RECT 296.950 379.710 297.510 380.210 ;
        RECT 300.780 379.790 301.500 385.460 ;
        RECT 302.250 386.190 316.540 386.750 ;
        RECT 327.470 386.580 328.000 387.480 ;
        RECT 329.110 387.420 331.480 387.870 ;
        RECT 302.250 381.890 325.600 386.190 ;
        RECT 329.140 385.460 330.090 387.420 ;
        RECT 330.840 387.400 331.420 387.420 ;
        RECT 341.220 386.760 345.130 388.220 ;
        RECT 352.450 387.570 356.580 387.970 ;
        RECT 352.450 387.480 356.590 387.570 ;
        RECT 331.510 386.750 345.130 386.760 ;
        RECT 326.370 384.770 326.940 384.780 ;
        RECT 302.250 381.610 316.540 381.890 ;
        RECT 312.630 380.060 316.540 381.610 ;
        RECT 326.370 381.350 326.990 384.770 ;
        RECT 326.370 381.340 326.940 381.350 ;
        RECT 296.960 379.490 297.510 379.710 ;
        RECT 312.610 379.290 316.560 380.060 ;
        RECT 325.540 379.710 326.100 380.210 ;
        RECT 329.370 379.790 330.090 385.460 ;
        RECT 330.840 386.190 345.130 386.750 ;
        RECT 356.060 386.580 356.590 387.480 ;
        RECT 330.840 381.890 354.190 386.190 ;
        RECT 354.960 384.770 355.530 384.780 ;
        RECT 330.840 381.610 345.130 381.890 ;
        RECT 341.220 380.060 345.130 381.610 ;
        RECT 354.960 381.350 355.580 384.770 ;
        RECT 354.960 381.340 355.530 381.350 ;
        RECT 325.550 379.490 326.100 379.710 ;
        RECT 341.200 379.290 345.150 380.060 ;
        RECT 354.130 379.710 354.690 380.210 ;
        RECT 354.140 379.490 354.690 379.710 ;
        RECT 255.700 378.680 256.090 379.290 ;
        RECT 256.170 378.700 256.360 379.010 ;
        RECT 256.610 378.700 256.770 379.010 ;
        RECT 241.190 376.090 241.610 378.600 ;
        RECT 243.670 377.460 243.900 378.600 ;
        RECT 243.580 376.090 244.300 377.460 ;
        RECT 236.450 375.740 244.300 376.090 ;
        RECT 236.450 374.310 236.640 375.740 ;
        RECT 236.200 374.160 236.640 374.310 ;
        RECT 237.230 374.160 237.650 374.310 ;
        RECT 236.200 374.020 237.650 374.160 ;
        RECT 236.450 373.610 236.640 374.020 ;
        RECT 231.890 369.250 233.180 370.590 ;
        RECT 231.900 368.760 233.180 369.250 ;
        RECT 228.090 368.270 228.320 368.390 ;
        RECT 233.860 368.310 234.180 368.610 ;
        RECT 226.660 368.190 226.890 368.270 ;
        RECT 227.880 368.190 228.110 368.270 ;
        RECT 230.170 368.120 231.610 368.280 ;
        RECT 233.670 368.190 233.900 368.280 ;
        RECT 234.890 368.200 235.120 368.280 ;
        RECT 235.150 366.520 235.570 372.570 ;
        RECT 237.630 369.710 237.860 372.570 ;
        RECT 237.630 369.420 237.960 369.710 ;
        RECT 236.620 367.660 236.820 367.700 ;
        RECT 236.260 367.580 236.460 367.610 ;
        RECT 236.170 367.080 236.480 367.580 ;
        RECT 232.350 365.810 232.700 366.290 ;
        RECT 227.910 365.460 228.080 365.640 ;
        RECT 227.890 364.870 228.210 365.170 ;
        RECT 227.890 364.760 228.130 364.870 ;
        RECT 227.920 364.750 228.090 364.760 ;
        RECT 228.110 364.700 228.130 364.760 ;
        RECT 228.360 362.610 228.830 363.100 ;
        RECT 224.000 356.260 224.240 357.670 ;
        RECT 225.610 357.340 225.990 357.670 ;
        RECT 227.930 356.280 228.170 357.670 ;
        RECT 223.990 355.600 224.250 356.260 ;
        RECT 227.910 355.620 228.180 356.280 ;
        RECT 224.000 352.990 224.240 355.600 ;
        RECT 227.930 353.100 228.170 355.620 ;
        RECT 228.410 353.100 228.810 362.610 ;
        RECT 229.330 362.000 229.750 362.360 ;
        RECT 227.930 353.030 228.810 353.100 ;
        RECT 221.370 352.940 222.410 352.990 ;
        RECT 221.560 351.170 222.410 352.940 ;
        RECT 222.980 352.890 223.540 352.990 ;
        RECT 221.370 346.940 221.610 347.010 ;
        RECT 221.910 345.300 222.410 351.170 ;
        RECT 223.040 350.470 223.540 352.890 ;
        RECT 223.990 352.670 224.250 352.990 ;
        RECT 225.300 352.920 225.540 352.990 ;
        RECT 227.320 352.940 227.480 352.990 ;
        RECT 227.690 352.940 227.880 352.990 ;
        RECT 227.920 352.820 228.810 353.030 ;
        RECT 227.920 352.710 228.290 352.820 ;
        RECT 224.000 351.170 224.240 352.670 ;
        RECT 227.930 352.650 228.290 352.710 ;
        RECT 225.610 351.170 225.990 351.770 ;
        RECT 227.930 351.170 228.170 352.650 ;
        RECT 222.990 349.910 223.540 350.470 ;
        RECT 223.040 347.090 223.540 349.910 ;
        RECT 222.980 346.940 223.540 347.090 ;
        RECT 225.300 346.940 225.540 347.000 ;
        RECT 227.320 346.950 227.480 347.010 ;
        RECT 227.690 346.950 227.880 347.010 ;
        RECT 228.130 346.950 228.290 347.010 ;
        RECT 221.900 344.740 222.420 345.300 ;
        RECT 221.910 344.150 222.410 344.740 ;
        RECT 220.780 343.690 221.290 344.150 ;
        RECT 221.910 343.690 222.550 344.150 ;
        RECT 220.780 342.770 221.280 343.690 ;
        RECT 220.660 342.450 221.280 342.770 ;
        RECT 220.780 342.340 221.280 342.450 ;
        RECT 220.660 342.020 221.280 342.340 ;
        RECT 220.520 340.910 220.750 341.110 ;
        RECT 220.780 340.070 221.280 342.020 ;
        RECT 221.600 341.490 221.830 343.300 ;
        RECT 221.910 341.120 222.410 343.690 ;
        RECT 223.040 343.160 223.540 346.940 ;
        RECT 222.860 341.630 223.540 343.160 ;
        RECT 221.780 340.910 222.410 341.120 ;
        RECT 220.770 340.000 221.290 340.070 ;
        RECT 220.660 339.680 221.290 340.000 ;
        RECT 220.770 339.570 221.290 339.680 ;
        RECT 220.660 339.550 221.290 339.570 ;
        RECT 220.660 339.250 221.280 339.550 ;
        RECT 219.690 334.220 220.350 334.790 ;
        RECT 203.960 332.710 204.330 333.290 ;
        RECT 203.430 331.820 203.800 332.400 ;
        RECT 202.940 330.910 203.310 331.490 ;
        RECT 198.360 329.360 198.680 329.680 ;
        RECT 199.460 329.360 199.780 329.680 ;
        RECT 200.550 329.360 200.870 329.680 ;
        RECT 193.170 328.650 193.490 328.970 ;
        RECT 194.270 328.650 194.590 328.970 ;
        RECT 195.370 328.650 195.730 328.970 ;
        RECT 201.200 328.950 201.530 330.370 ;
        RECT 202.470 330.020 202.820 330.590 ;
        RECT 195.460 327.600 195.730 328.650 ;
        RECT 198.910 328.630 199.230 328.950 ;
        RECT 200.010 328.630 200.330 328.950 ;
        RECT 201.110 328.630 201.530 328.950 ;
        RECT 193.170 327.280 193.490 327.600 ;
        RECT 194.270 327.280 194.590 327.600 ;
        RECT 195.370 327.280 195.730 327.600 ;
        RECT 201.200 327.580 201.530 328.630 ;
        RECT 201.980 328.450 202.250 328.480 ;
        RECT 201.970 327.920 202.250 328.450 ;
        RECT 201.970 327.620 202.430 327.920 ;
        RECT 192.620 326.610 192.940 326.930 ;
        RECT 193.720 326.600 194.040 326.920 ;
        RECT 194.810 326.600 195.130 326.920 ;
        RECT 195.460 326.400 195.730 327.280 ;
        RECT 198.910 327.260 199.230 327.580 ;
        RECT 200.010 327.260 200.330 327.580 ;
        RECT 201.110 327.260 201.530 327.580 ;
        RECT 195.940 326.640 196.260 326.960 ;
        RECT 198.360 326.590 198.680 326.910 ;
        RECT 199.460 326.580 199.780 326.900 ;
        RECT 200.550 326.580 200.870 326.900 ;
        RECT 195.350 325.840 195.840 326.400 ;
        RECT 195.930 326.170 196.250 326.490 ;
        RECT 190.910 324.810 192.930 324.850 ;
        RECT 180.620 324.750 182.550 324.790 ;
        RECT 180.080 323.560 182.550 324.750 ;
        RECT 167.600 319.330 167.970 319.710 ;
        RECT 166.950 318.710 167.340 319.100 ;
        RECT 166.350 318.080 166.730 318.470 ;
        RECT 165.760 317.450 166.110 317.820 ;
        RECT 165.120 316.770 165.480 317.150 ;
        RECT 164.530 316.530 164.870 316.540 ;
        RECT 164.510 316.160 164.890 316.530 ;
        RECT 164.530 316.150 164.860 316.160 ;
        RECT 162.750 314.310 163.100 314.640 ;
        RECT 162.770 314.250 163.100 314.310 ;
        RECT 161.480 313.030 161.830 313.360 ;
        RECT 161.480 312.960 161.810 313.030 ;
        RECT 159.340 312.300 160.580 312.630 ;
        RECT 160.870 312.330 161.310 312.750 ;
        RECT 31.850 312.240 32.350 312.250 ;
        RECT 159.340 312.190 159.920 312.300 ;
        RECT 180.080 312.070 181.020 323.560 ;
        RECT 190.430 323.530 192.930 324.810 ;
        RECT 192.040 313.530 192.930 323.530 ;
        RECT 201.200 320.380 201.530 327.260 ;
        RECT 201.960 327.600 202.430 327.620 ;
        RECT 201.960 327.170 202.250 327.600 ;
        RECT 201.680 326.620 202.000 326.940 ;
        RECT 201.670 326.150 201.990 326.470 ;
        RECT 219.850 325.910 220.350 334.220 ;
        RECT 220.780 338.350 221.280 339.250 ;
        RECT 221.600 338.720 221.830 340.530 ;
        RECT 221.910 339.850 222.410 340.910 ;
        RECT 223.040 340.390 223.540 341.630 ;
        RECT 221.910 339.800 222.550 339.850 ;
        RECT 221.910 339.790 222.560 339.800 ;
        RECT 221.910 339.470 222.580 339.790 ;
        RECT 221.910 338.350 222.410 339.470 ;
        RECT 222.860 338.860 223.540 340.390 ;
        RECT 220.780 338.100 221.290 338.350 ;
        RECT 221.910 338.100 222.550 338.350 ;
        RECT 220.780 326.820 221.280 338.100 ;
        RECT 221.910 327.690 222.410 338.100 ;
        RECT 223.040 329.200 223.540 338.860 ;
        RECT 225.930 336.760 226.510 337.320 ;
        RECT 225.960 336.750 226.470 336.760 ;
        RECT 223.040 328.640 223.600 329.200 ;
        RECT 223.040 328.510 223.540 328.640 ;
        RECT 225.960 324.880 226.460 336.750 ;
        RECT 225.330 323.600 226.460 324.880 ;
        RECT 227.200 324.220 227.430 326.190 ;
        RECT 227.200 323.990 227.560 324.220 ;
        RECT 227.200 322.610 227.430 323.990 ;
        RECT 227.200 322.380 227.560 322.610 ;
        RECT 227.200 321.010 227.430 322.380 ;
        RECT 227.200 320.780 227.560 321.010 ;
        RECT 201.140 319.990 201.570 320.380 ;
        RECT 227.200 319.390 227.430 320.780 ;
        RECT 227.200 319.160 227.560 319.390 ;
        RECT 228.410 319.260 228.810 352.820 ;
        RECT 229.340 319.800 229.730 362.000 ;
        RECT 230.250 359.610 230.700 360.040 ;
        RECT 229.950 357.400 230.110 357.440 ;
        RECT 230.270 354.510 230.660 359.610 ;
        RECT 231.110 359.350 231.490 359.360 ;
        RECT 231.090 359.050 231.510 359.350 ;
        RECT 230.760 357.390 230.920 357.440 ;
        RECT 230.100 354.320 230.660 354.510 ;
        RECT 230.270 319.800 230.660 354.320 ;
        RECT 228.910 319.600 230.920 319.800 ;
        RECT 227.200 317.790 227.430 319.160 ;
        RECT 228.400 318.800 228.870 319.260 ;
        RECT 229.340 318.460 229.730 319.600 ;
        RECT 228.020 318.080 228.340 318.250 ;
        RECT 229.310 318.080 229.770 318.460 ;
        RECT 228.020 317.990 229.770 318.080 ;
        RECT 228.220 317.900 229.760 317.990 ;
        RECT 227.200 317.560 227.560 317.790 ;
        RECT 230.270 317.640 230.660 319.600 ;
        RECT 227.200 316.170 227.430 317.560 ;
        RECT 230.250 317.180 230.720 317.640 ;
        RECT 230.750 316.350 230.920 319.600 ;
        RECT 231.110 319.760 231.490 359.050 ;
        RECT 231.840 357.480 232.160 357.800 ;
        RECT 231.840 356.930 232.160 357.250 ;
        RECT 231.840 354.820 232.160 355.140 ;
        RECT 231.840 354.240 232.160 354.590 ;
        RECT 231.840 353.690 232.160 354.010 ;
        RECT 231.840 351.590 232.160 351.910 ;
        RECT 231.840 351.040 232.160 351.360 ;
        RECT 232.450 335.820 232.680 365.810 ;
        RECT 233.700 365.460 233.870 365.640 ;
        RECT 233.590 364.800 233.910 365.120 ;
        RECT 233.700 364.750 233.870 364.800 ;
        RECT 236.260 363.830 236.460 367.080 ;
        RECT 237.630 366.520 237.860 369.420 ;
        RECT 238.850 368.200 239.080 372.570 ;
        RECT 239.770 369.790 239.960 375.740 ;
        RECT 240.930 374.230 241.160 374.310 ;
        RECT 241.190 372.550 241.610 375.740 ;
        RECT 243.670 375.450 244.000 375.740 ;
        RECT 243.670 375.350 243.900 375.450 ;
        RECT 243.110 375.260 243.930 375.350 ;
        RECT 243.050 374.570 243.930 375.260 ;
        RECT 243.050 372.550 243.900 374.570 ;
        RECT 244.890 372.550 245.120 378.600 ;
        RECT 251.410 378.560 251.600 378.600 ;
        RECT 250.180 377.000 250.500 377.290 ;
        RECT 251.850 377.000 252.130 378.600 ;
        RECT 254.650 378.250 254.960 378.640 ;
        RECT 254.650 378.200 255.200 378.250 ;
        RECT 254.940 377.460 255.200 378.200 ;
        RECT 247.980 376.230 252.130 377.000 ;
        RECT 247.450 374.230 247.640 374.310 ;
        RECT 247.890 374.290 248.170 374.310 ;
        RECT 247.890 374.230 248.230 374.290 ;
        RECT 247.910 373.990 248.230 374.230 ;
        RECT 249.660 372.650 250.050 376.230 ;
        RECT 251.100 375.810 251.360 376.130 ;
        RECT 251.850 375.850 252.130 376.230 ;
        RECT 255.770 376.200 256.010 376.580 ;
        RECT 251.850 375.530 252.300 375.850 ;
        RECT 256.110 375.550 259.340 378.700 ;
        RECT 276.580 376.230 280.530 377.000 ;
        RECT 251.100 375.210 251.360 375.530 ;
        RECT 250.180 374.210 250.500 374.530 ;
        RECT 251.850 374.310 252.130 375.530 ;
        RECT 252.720 375.280 253.040 375.360 ;
        RECT 252.720 375.040 253.290 375.280 ;
        RECT 252.950 374.710 253.290 375.040 ;
        RECT 252.670 374.390 253.290 374.710 ;
        RECT 251.580 374.170 252.130 374.310 ;
        RECT 239.630 369.690 239.960 369.790 ;
        RECT 239.530 369.370 239.960 369.690 ;
        RECT 239.710 368.960 239.960 369.370 ;
        RECT 240.190 369.580 240.380 369.860 ;
        RECT 240.190 369.290 240.500 369.580 ;
        RECT 241.860 369.480 242.120 369.780 ;
        RECT 241.840 369.460 242.120 369.480 ;
        RECT 239.290 368.600 239.610 368.920 ;
        RECT 239.710 368.870 240.040 368.960 ;
        RECT 239.770 368.670 240.040 368.870 ;
        RECT 239.770 368.610 239.960 368.670 ;
        RECT 239.660 368.310 239.980 368.610 ;
        RECT 240.190 368.340 240.380 369.290 ;
        RECT 241.840 368.970 242.030 369.460 ;
        RECT 240.960 368.600 241.280 368.920 ;
        RECT 241.840 368.890 242.150 368.970 ;
        RECT 241.820 368.680 242.150 368.890 ;
        RECT 241.820 368.600 242.050 368.680 ;
        RECT 238.840 368.040 239.080 368.200 ;
        RECT 238.840 367.980 239.180 368.040 ;
        RECT 238.830 367.720 239.180 367.980 ;
        RECT 239.250 367.770 239.450 368.090 ;
        RECT 238.830 367.690 239.080 367.720 ;
        RECT 238.850 366.520 239.080 367.690 ;
        RECT 239.250 367.480 239.570 367.770 ;
        RECT 239.250 366.480 239.450 367.480 ;
        RECT 239.770 366.590 239.960 368.310 ;
        RECT 241.410 368.200 241.600 368.280 ;
        RECT 241.850 368.230 242.130 368.280 ;
        RECT 241.850 367.930 242.170 368.230 ;
        RECT 242.760 368.050 242.950 368.090 ;
        RECT 240.130 367.640 240.320 367.700 ;
        RECT 239.630 366.490 239.960 366.590 ;
        RECT 239.530 366.170 239.960 366.490 ;
        RECT 239.250 365.720 239.450 365.970 ;
        RECT 239.710 365.760 239.960 366.170 ;
        RECT 240.190 366.380 240.380 366.660 ;
        RECT 240.190 366.090 240.500 366.380 ;
        RECT 241.860 366.280 242.120 366.580 ;
        RECT 242.760 366.480 242.950 366.530 ;
        RECT 241.840 366.260 242.120 366.280 ;
        RECT 239.250 365.400 239.610 365.720 ;
        RECT 239.710 365.670 240.040 365.760 ;
        RECT 239.770 365.470 240.040 365.670 ;
        RECT 238.840 364.840 239.060 365.000 ;
        RECT 239.250 364.970 239.450 365.400 ;
        RECT 238.840 364.780 239.180 364.840 ;
        RECT 238.830 364.470 239.180 364.780 ;
        RECT 238.840 364.410 239.180 364.470 ;
        RECT 239.250 364.680 239.570 364.970 ;
        RECT 239.250 364.570 239.450 364.680 ;
        RECT 238.840 364.250 239.060 364.410 ;
        RECT 239.250 364.280 239.570 364.570 ;
        RECT 239.250 363.850 239.450 364.280 ;
        RECT 239.250 363.530 239.610 363.850 ;
        RECT 239.770 363.840 239.960 365.470 ;
        RECT 240.190 365.140 240.380 366.090 ;
        RECT 241.840 365.770 242.030 366.260 ;
        RECT 242.760 365.920 242.950 365.970 ;
        RECT 240.960 365.400 241.280 365.720 ;
        RECT 241.840 365.690 242.150 365.770 ;
        RECT 241.820 365.480 242.150 365.690 ;
        RECT 241.820 365.400 242.050 365.480 ;
        RECT 242.760 364.850 242.950 364.890 ;
        RECT 242.760 364.360 242.950 364.400 ;
        RECT 239.810 363.580 240.040 363.780 ;
        RECT 239.250 363.280 239.450 363.530 ;
        RECT 239.710 363.490 240.040 363.580 ;
        RECT 239.710 363.080 239.900 363.490 ;
        RECT 239.530 362.830 239.900 363.080 ;
        RECT 240.190 363.160 240.380 364.110 ;
        RECT 240.960 363.530 241.280 363.850 ;
        RECT 241.820 363.770 242.050 363.850 ;
        RECT 242.130 363.770 242.450 363.870 ;
        RECT 241.820 363.560 242.450 363.770 ;
        RECT 241.840 363.550 242.450 363.560 ;
        RECT 241.840 363.480 242.150 363.550 ;
        RECT 240.190 362.870 240.500 363.160 ;
        RECT 241.840 362.990 242.030 363.480 ;
        RECT 242.760 363.280 242.950 363.330 ;
        RECT 241.840 362.970 242.120 362.990 ;
        RECT 233.590 362.290 233.910 362.590 ;
        RECT 239.250 361.770 239.450 362.770 ;
        RECT 239.530 362.760 239.890 362.830 ;
        RECT 239.630 362.660 239.890 362.760 ;
        RECT 240.190 362.590 240.380 362.870 ;
        RECT 241.860 362.670 242.120 362.970 ;
        RECT 242.280 362.720 242.600 363.040 ;
        RECT 242.760 362.720 242.950 362.770 ;
        RECT 241.410 362.230 241.600 362.280 ;
        RECT 241.850 362.230 242.130 362.280 ;
        RECT 241.450 361.890 241.770 362.210 ;
        RECT 242.530 361.780 242.740 361.990 ;
        RECT 236.620 361.650 236.820 361.690 ;
        RECT 232.840 357.340 233.000 358.070 ;
        RECT 232.840 357.320 233.040 357.340 ;
        RECT 232.820 357.080 233.050 357.320 ;
        RECT 232.840 357.030 233.050 357.080 ;
        RECT 233.210 357.030 233.400 358.020 ;
        RECT 233.650 357.370 233.810 358.070 ;
        RECT 232.840 356.170 233.000 357.030 ;
        RECT 233.230 356.910 233.400 357.030 ;
        RECT 233.240 356.170 233.400 356.910 ;
        RECT 233.540 356.820 233.810 357.370 ;
        RECT 233.540 356.770 233.820 356.820 ;
        RECT 233.650 356.680 233.820 356.770 ;
        RECT 233.650 356.170 233.810 356.680 ;
        RECT 232.840 355.040 233.000 355.900 ;
        RECT 233.240 355.160 233.400 355.900 ;
        RECT 233.650 355.390 233.810 355.900 ;
        RECT 233.650 355.300 233.820 355.390 ;
        RECT 233.230 355.040 233.400 355.160 ;
        RECT 232.840 354.990 233.050 355.040 ;
        RECT 232.820 354.750 233.050 354.990 ;
        RECT 232.840 354.730 233.040 354.750 ;
        RECT 232.840 354.100 233.000 354.730 ;
        RECT 232.840 354.080 233.040 354.100 ;
        RECT 232.820 353.840 233.050 354.080 ;
        RECT 232.840 353.790 233.050 353.840 ;
        RECT 233.210 353.790 233.400 355.040 ;
        RECT 233.540 355.250 233.820 355.300 ;
        RECT 233.540 354.700 233.810 355.250 ;
        RECT 235.180 355.120 235.560 361.620 ;
        RECT 238.830 361.530 239.060 361.560 ;
        RECT 238.830 361.270 239.180 361.530 ;
        RECT 238.840 361.210 239.180 361.270 ;
        RECT 239.250 361.480 239.570 361.770 ;
        RECT 240.130 361.650 240.320 361.710 ;
        RECT 238.840 361.050 239.060 361.210 ;
        RECT 239.250 361.160 239.450 361.480 ;
        RECT 242.530 361.460 242.860 361.780 ;
        RECT 239.290 360.330 239.610 360.650 ;
        RECT 239.810 360.380 240.040 360.580 ;
        RECT 239.710 360.290 240.040 360.380 ;
        RECT 236.050 358.140 236.440 360.000 ;
        RECT 239.710 359.880 239.900 360.290 ;
        RECT 240.190 359.960 240.380 360.910 ;
        RECT 240.960 360.330 241.280 360.650 ;
        RECT 241.820 360.570 242.050 360.650 ;
        RECT 242.180 360.610 242.500 360.930 ;
        RECT 241.820 360.360 242.150 360.570 ;
        RECT 241.840 360.280 242.150 360.360 ;
        RECT 240.190 359.930 240.500 359.960 ;
        RECT 239.530 359.630 239.900 359.880 ;
        RECT 240.080 359.670 240.500 359.930 ;
        RECT 241.840 359.790 242.030 360.280 ;
        RECT 242.530 360.220 242.740 361.460 ;
        RECT 242.760 361.160 242.950 361.200 ;
        RECT 242.610 359.900 242.840 360.190 ;
        RECT 241.840 359.770 242.120 359.790 ;
        RECT 239.530 359.560 239.890 359.630 ;
        RECT 239.630 359.460 239.890 359.560 ;
        RECT 240.080 358.070 240.470 359.670 ;
        RECT 241.860 359.470 242.120 359.770 ;
        RECT 243.050 355.570 243.760 372.550 ;
        RECT 245.370 372.530 245.560 372.570 ;
        RECT 244.140 370.940 244.460 371.260 ;
        RECT 245.060 369.780 245.320 370.100 ;
        RECT 245.810 369.820 246.090 372.570 ;
        RECT 248.610 372.220 248.920 372.610 ;
        RECT 248.610 372.170 249.160 372.220 ;
        RECT 248.900 371.430 249.160 372.170 ;
        RECT 250.130 371.530 250.320 372.980 ;
        RECT 250.570 372.340 250.730 372.980 ;
        RECT 251.410 372.550 251.600 372.600 ;
        RECT 251.850 372.550 252.130 374.170 ;
        RECT 252.240 374.160 252.520 374.310 ;
        RECT 252.950 373.440 253.290 374.390 ;
        RECT 252.670 373.120 253.290 373.440 ;
        RECT 252.950 372.790 253.290 373.120 ;
        RECT 252.720 372.470 253.290 372.790 ;
        RECT 252.950 372.360 253.290 372.470 ;
        RECT 250.460 371.790 250.730 372.340 ;
        RECT 252.720 372.040 253.290 372.360 ;
        RECT 250.460 371.740 250.740 371.790 ;
        RECT 250.570 371.650 250.740 371.740 ;
        RECT 252.950 371.710 253.290 372.040 ;
        RECT 250.130 371.500 250.350 371.530 ;
        RECT 250.110 371.230 250.360 371.500 ;
        RECT 250.120 371.220 250.360 371.230 ;
        RECT 250.120 370.980 250.350 371.220 ;
        RECT 249.730 370.170 249.970 370.550 ;
        RECT 250.160 369.960 250.320 370.980 ;
        RECT 250.570 369.960 250.730 371.650 ;
        RECT 252.670 371.390 253.290 371.710 ;
        RECT 252.950 370.440 253.290 371.390 ;
        RECT 252.670 370.120 253.290 370.440 ;
        RECT 245.810 369.500 246.260 369.820 ;
        RECT 248.170 369.580 248.490 369.900 ;
        RECT 252.950 369.790 253.290 370.120 ;
        RECT 252.720 369.560 253.290 369.790 ;
        RECT 253.620 374.950 253.890 375.270 ;
        RECT 254.380 375.000 254.700 375.320 ;
        RECT 255.350 375.270 259.340 375.550 ;
        RECT 255.330 375.070 259.340 375.270 ;
        RECT 253.620 374.660 253.930 374.950 ;
        RECT 253.620 373.920 253.890 374.660 ;
        RECT 253.620 373.630 254.000 373.920 ;
        RECT 253.620 373.170 253.890 373.630 ;
        RECT 255.150 373.590 259.500 375.070 ;
        RECT 253.620 372.880 253.930 373.170 ;
        RECT 254.430 372.950 254.750 373.100 ;
        RECT 254.940 372.950 259.500 373.590 ;
        RECT 253.620 371.950 253.890 372.880 ;
        RECT 254.430 372.800 259.500 372.950 ;
        RECT 254.430 372.780 254.960 372.800 ;
        RECT 254.650 372.510 254.960 372.780 ;
        RECT 254.420 372.060 254.740 372.380 ;
        RECT 253.620 371.660 253.930 371.950 ;
        RECT 253.620 371.330 253.890 371.660 ;
        RECT 255.150 371.370 259.500 372.800 ;
        RECT 253.620 371.040 254.000 371.330 ;
        RECT 253.620 370.170 253.890 371.040 ;
        RECT 284.700 370.890 287.930 378.700 ;
        RECT 305.160 376.230 309.110 377.000 ;
        RECT 253.620 369.880 253.930 370.170 ;
        RECT 253.620 369.570 253.890 369.880 ;
        RECT 254.340 369.810 254.660 370.130 ;
        RECT 245.060 369.180 245.320 369.500 ;
        RECT 244.140 368.180 244.460 368.500 ;
        RECT 245.810 368.280 246.090 369.500 ;
        RECT 252.720 369.470 253.040 369.560 ;
        RECT 246.680 369.250 247.000 369.330 ;
        RECT 246.680 369.010 247.250 369.250 ;
        RECT 246.910 368.680 247.250 369.010 ;
        RECT 246.630 368.360 247.250 368.680 ;
        RECT 245.540 368.140 246.090 368.280 ;
        RECT 245.370 366.520 245.560 366.570 ;
        RECT 245.810 366.520 246.090 368.140 ;
        RECT 246.200 368.130 246.480 368.280 ;
        RECT 246.910 367.410 247.250 368.360 ;
        RECT 247.580 368.920 247.850 369.240 ;
        RECT 248.340 369.070 248.660 369.290 ;
        RECT 248.320 368.970 248.660 369.070 ;
        RECT 247.580 368.630 247.890 368.920 ;
        RECT 248.320 368.750 248.640 368.970 ;
        RECT 247.580 368.310 247.850 368.630 ;
        RECT 249.730 368.540 249.970 368.920 ;
        RECT 250.160 368.760 250.320 369.130 ;
        RECT 250.050 368.460 250.370 368.760 ;
        RECT 250.050 368.430 250.480 368.460 ;
        RECT 250.570 368.430 250.730 369.130 ;
        RECT 251.080 368.450 251.590 368.460 ;
        RECT 251.080 368.430 251.920 368.450 ;
        RECT 250.050 368.400 251.920 368.430 ;
        RECT 247.450 368.260 247.850 368.310 ;
        RECT 247.890 368.260 248.170 368.310 ;
        RECT 250.160 368.300 251.920 368.400 ;
        RECT 247.580 368.240 247.850 368.260 ;
        RECT 247.490 367.920 247.850 368.240 ;
        RECT 250.160 368.110 250.320 368.300 ;
        RECT 250.330 368.290 251.290 368.300 ;
        RECT 246.630 367.090 247.250 367.410 ;
        RECT 246.910 366.760 247.250 367.090 ;
        RECT 246.680 366.440 247.250 366.760 ;
        RECT 246.910 366.330 247.250 366.440 ;
        RECT 246.680 366.010 247.250 366.330 ;
        RECT 246.910 365.680 247.250 366.010 ;
        RECT 246.630 365.360 247.250 365.680 ;
        RECT 246.910 364.410 247.250 365.360 ;
        RECT 246.630 364.090 247.250 364.410 ;
        RECT 246.910 363.760 247.250 364.090 ;
        RECT 246.680 363.530 247.250 363.760 ;
        RECT 247.580 367.890 247.850 367.920 ;
        RECT 247.580 367.600 247.960 367.890 ;
        RECT 248.570 367.810 248.780 368.020 ;
        RECT 250.120 367.870 250.350 368.110 ;
        RECT 250.120 367.860 250.360 367.870 ;
        RECT 247.580 367.140 247.850 367.600 ;
        RECT 248.570 367.560 248.900 367.810 ;
        RECT 250.110 367.590 250.360 367.860 ;
        RECT 250.130 367.560 250.350 367.590 ;
        RECT 248.570 367.490 249.160 367.560 ;
        RECT 247.580 366.850 247.890 367.140 ;
        RECT 248.570 367.070 248.780 367.490 ;
        RECT 248.390 366.960 248.780 367.070 ;
        RECT 248.220 366.920 248.780 366.960 ;
        RECT 248.900 366.920 249.160 367.490 ;
        RECT 247.580 365.920 247.850 366.850 ;
        RECT 248.220 366.770 249.160 366.920 ;
        RECT 248.220 366.750 248.920 366.770 ;
        RECT 248.220 366.640 248.540 366.750 ;
        RECT 248.570 366.480 248.920 366.750 ;
        RECT 248.570 366.350 248.780 366.480 ;
        RECT 248.380 366.250 248.780 366.350 ;
        RECT 248.380 366.220 248.700 366.250 ;
        RECT 248.380 366.030 248.880 366.220 ;
        RECT 250.130 366.110 250.320 367.560 ;
        RECT 250.570 367.440 250.730 368.290 ;
        RECT 251.580 368.260 251.920 368.300 ;
        RECT 252.250 368.260 252.520 368.470 ;
        RECT 250.570 367.350 250.740 367.440 ;
        RECT 250.460 367.300 250.740 367.350 ;
        RECT 250.460 366.750 250.730 367.300 ;
        RECT 284.400 366.840 287.950 370.890 ;
        RECT 250.570 366.110 250.730 366.750 ;
        RECT 248.650 365.930 248.880 366.030 ;
        RECT 247.580 365.630 247.890 365.920 ;
        RECT 247.580 365.300 247.850 365.630 ;
        RECT 247.580 365.010 247.960 365.300 ;
        RECT 313.290 365.260 316.520 378.700 ;
        RECT 333.750 376.230 337.700 377.000 ;
        RECT 247.580 364.140 247.850 365.010 ;
        RECT 247.580 363.850 247.890 364.140 ;
        RECT 247.580 363.540 247.850 363.850 ;
        RECT 248.300 363.780 248.620 364.100 ;
        RECT 246.680 363.440 247.000 363.530 ;
        RECT 313.090 362.730 316.680 365.260 ;
        RECT 244.030 362.430 244.360 362.720 ;
        RECT 244.020 362.400 244.440 362.430 ;
        RECT 245.040 362.420 245.540 362.430 ;
        RECT 245.040 362.400 245.880 362.420 ;
        RECT 244.020 362.290 245.880 362.400 ;
        RECT 244.300 362.260 245.200 362.290 ;
        RECT 245.540 362.230 245.880 362.290 ;
        RECT 246.210 362.230 246.480 362.440 ;
        RECT 341.880 361.770 345.110 378.700 ;
        RECT 341.570 358.150 345.330 361.770 ;
        RECT 355.920 361.080 359.330 361.400 ;
        RECT 355.920 357.850 362.560 361.080 ;
        RECT 242.920 354.780 243.760 355.570 ;
        RECT 233.650 354.130 233.810 354.700 ;
        RECT 232.840 352.930 233.000 353.790 ;
        RECT 233.230 353.670 233.400 353.790 ;
        RECT 233.240 352.930 233.400 353.670 ;
        RECT 233.540 353.580 233.810 354.130 ;
        RECT 233.540 353.530 233.820 353.580 ;
        RECT 233.650 353.440 233.820 353.530 ;
        RECT 233.650 352.930 233.810 353.440 ;
        RECT 232.840 351.810 233.000 352.670 ;
        RECT 233.240 351.930 233.400 352.670 ;
        RECT 233.650 352.160 233.810 352.670 ;
        RECT 233.650 352.070 233.820 352.160 ;
        RECT 233.230 351.810 233.400 351.930 ;
        RECT 232.840 351.760 233.050 351.810 ;
        RECT 232.820 351.520 233.050 351.760 ;
        RECT 232.840 351.500 233.040 351.520 ;
        RECT 232.840 350.770 233.000 351.500 ;
        RECT 233.210 350.820 233.400 351.810 ;
        RECT 233.540 352.020 233.820 352.070 ;
        RECT 233.540 351.470 233.810 352.020 ;
        RECT 233.650 350.770 233.810 351.470 ;
        RECT 238.640 336.740 239.360 337.310 ;
        RECT 232.450 335.590 232.690 335.820 ;
        RECT 232.450 329.780 232.680 335.590 ;
        RECT 238.700 329.730 239.210 336.740 ;
        RECT 238.560 329.680 239.210 329.730 ;
        RECT 238.550 329.500 239.210 329.680 ;
        RECT 238.520 329.490 239.210 329.500 ;
        RECT 238.520 329.120 239.120 329.490 ;
        RECT 238.520 327.250 239.100 329.120 ;
        RECT 264.240 327.690 268.660 357.800 ;
        RECT 355.920 357.360 359.330 357.850 ;
        RECT 347.510 332.490 349.830 332.570 ;
        RECT 347.510 329.260 362.550 332.490 ;
        RECT 347.510 329.200 349.830 329.260 ;
        RECT 238.170 326.260 239.100 327.250 ;
        RECT 264.210 326.370 268.680 327.690 ;
        RECT 238.520 325.480 239.100 326.260 ;
        RECT 238.570 324.880 239.100 325.480 ;
        RECT 238.530 324.870 239.100 324.880 ;
        RECT 238.520 323.870 239.100 324.870 ;
        RECT 232.850 323.250 233.170 323.570 ;
        RECT 238.570 323.270 239.100 323.870 ;
        RECT 232.850 322.580 233.170 322.900 ;
        RECT 238.520 322.260 239.100 323.270 ;
        RECT 238.560 321.660 239.100 322.260 ;
        RECT 233.120 321.560 233.440 321.610 ;
        RECT 232.890 321.330 233.440 321.560 ;
        RECT 233.120 321.290 233.440 321.330 ;
        RECT 238.520 320.640 239.100 321.660 ;
        RECT 238.570 320.040 239.100 320.640 ;
        RECT 233.120 319.950 233.440 320.000 ;
        RECT 231.110 319.540 231.630 319.760 ;
        RECT 232.890 319.720 233.440 319.950 ;
        RECT 233.120 319.680 233.440 319.720 ;
        RECT 231.110 316.840 231.490 319.540 ;
        RECT 238.520 319.030 239.100 320.040 ;
        RECT 238.560 318.430 239.100 319.030 ;
        RECT 233.110 318.340 233.430 318.390 ;
        RECT 232.060 317.960 232.570 318.180 ;
        RECT 232.880 318.110 233.430 318.340 ;
        RECT 233.110 318.070 233.430 318.110 ;
        RECT 232.280 317.950 232.570 317.960 ;
        RECT 231.080 316.380 231.520 316.840 ;
        RECT 233.120 316.720 233.440 316.770 ;
        RECT 232.890 316.600 233.440 316.720 ;
        RECT 232.890 316.490 233.920 316.600 ;
        RECT 238.520 316.560 239.100 318.430 ;
        RECT 233.120 316.450 233.920 316.490 ;
        RECT 233.410 316.380 233.920 316.450 ;
        RECT 233.410 316.370 233.700 316.380 ;
        RECT 227.200 315.940 227.560 316.170 ;
        RECT 227.200 314.570 227.430 315.940 ;
        RECT 233.110 315.110 233.430 315.160 ;
        RECT 232.880 314.880 233.430 315.110 ;
        RECT 233.110 314.840 233.430 314.880 ;
        RECT 227.200 314.340 227.560 314.570 ;
        RECT 238.560 314.350 239.100 316.560 ;
        RECT 192.040 312.800 192.960 313.530 ;
        RECT 227.200 312.950 227.430 314.340 ;
        RECT 232.350 313.360 232.670 313.680 ;
        RECT 232.400 313.130 232.630 313.360 ;
        RECT 192.010 312.070 192.930 312.800 ;
        RECT 227.200 312.720 227.560 312.950 ;
        RECT 227.200 312.650 227.430 312.720 ;
        RECT 233.110 311.910 233.430 311.960 ;
        RECT 232.880 311.680 233.430 311.910 ;
        RECT 233.110 311.640 233.430 311.680 ;
        RECT 229.870 310.200 230.190 310.250 ;
        RECT 230.810 310.200 231.130 310.250 ;
        RECT 229.640 309.970 230.190 310.200 ;
        RECT 230.580 309.970 231.130 310.200 ;
        RECT 231.760 310.180 232.080 310.230 ;
        RECT 233.070 310.200 233.390 310.250 ;
        RECT 229.870 309.930 230.190 309.970 ;
        RECT 230.810 309.930 231.130 309.970 ;
        RECT 231.530 309.950 232.080 310.180 ;
        RECT 232.840 309.970 233.390 310.200 ;
        RECT 231.760 309.910 232.080 309.950 ;
        RECT 233.070 309.930 233.390 309.970 ;
        RECT 10.340 303.240 30.170 304.620 ;
        RECT 32.000 303.240 32.770 303.260 ;
        RECT 10.340 301.390 32.770 303.240 ;
        RECT 22.360 301.130 32.770 301.390 ;
        RECT 22.520 301.120 32.770 301.130 ;
        RECT 23.470 300.770 32.770 301.120 ;
        RECT 23.840 299.330 32.770 300.770 ;
        RECT 21.900 294.780 22.490 298.390 ;
        RECT 21.900 294.490 23.840 294.780 ;
        RECT 23.380 289.590 24.190 290.940 ;
        RECT 25.300 289.620 30.450 299.330 ;
        RECT 32.000 299.310 32.770 299.330 ;
        RECT 35.050 291.870 35.690 295.810 ;
        RECT 23.380 289.530 24.640 289.590 ;
        RECT 23.380 288.950 24.660 289.530 ;
        RECT 25.310 288.950 30.450 289.620 ;
        RECT 23.380 288.200 24.640 288.950 ;
        RECT 23.380 287.480 32.270 288.200 ;
        RECT 23.380 287.250 26.600 287.480 ;
        RECT 23.380 287.220 24.640 287.250 ;
        RECT 23.380 287.040 24.190 287.220 ;
        RECT 24.490 286.100 25.480 286.110 ;
        RECT 24.090 285.580 25.480 286.100 ;
        RECT 24.090 281.970 24.580 285.580 ;
        RECT 27.290 285.050 30.710 285.100 ;
        RECT 27.280 284.480 30.720 285.050 ;
        RECT 25.870 276.030 30.170 283.710 ;
        RECT 31.850 283.660 32.570 284.210 ;
        RECT 31.850 283.650 32.350 283.660 ;
        RECT 32.120 276.030 34.530 276.130 ;
        RECT 10.330 272.800 34.530 276.030 ;
        RECT 22.360 272.700 34.530 272.800 ;
        RECT 22.360 272.540 32.770 272.700 ;
        RECT 22.520 272.530 32.770 272.540 ;
        RECT 23.470 272.180 32.770 272.530 ;
        RECT 23.840 270.740 32.770 272.180 ;
        RECT 21.900 266.190 22.490 269.800 ;
        RECT 21.900 265.900 23.840 266.190 ;
        RECT 23.380 261.000 24.190 262.360 ;
        RECT 25.300 261.030 30.450 270.740 ;
        RECT 32.000 270.720 32.770 270.740 ;
        RECT 35.050 263.280 35.690 267.220 ;
        RECT 23.380 260.940 24.640 261.000 ;
        RECT 23.380 260.360 24.660 260.940 ;
        RECT 25.310 260.360 30.450 261.030 ;
        RECT 23.380 259.610 24.640 260.360 ;
        RECT 23.380 258.890 32.270 259.610 ;
        RECT 23.380 258.660 26.600 258.890 ;
        RECT 23.380 258.630 24.640 258.660 ;
        RECT 23.380 258.460 24.190 258.630 ;
        RECT 24.490 257.510 25.480 257.520 ;
        RECT 24.090 256.990 25.480 257.510 ;
        RECT 24.090 253.380 24.580 256.990 ;
        RECT 27.290 256.460 30.710 256.510 ;
        RECT 27.280 255.890 30.720 256.460 ;
        RECT 25.870 247.440 30.170 255.120 ;
        RECT 31.850 255.070 32.570 255.620 ;
        RECT 31.850 255.060 32.350 255.070 ;
        RECT 36.680 247.440 38.950 247.510 ;
        RECT 10.340 244.210 38.950 247.440 ;
        RECT 22.360 243.950 32.770 244.210 ;
        RECT 36.680 244.110 38.950 244.210 ;
        RECT 22.520 243.940 32.770 243.950 ;
        RECT 23.470 243.590 32.770 243.940 ;
        RECT 23.840 242.150 32.770 243.590 ;
        RECT 21.900 237.600 22.490 241.210 ;
        RECT 21.900 237.310 23.840 237.600 ;
        RECT 23.400 232.410 24.210 233.770 ;
        RECT 25.300 232.440 30.450 242.150 ;
        RECT 32.000 242.130 32.770 242.150 ;
        RECT 35.050 234.680 35.690 238.620 ;
        RECT 23.400 232.350 24.640 232.410 ;
        RECT 23.400 231.770 24.660 232.350 ;
        RECT 25.310 231.770 30.450 232.440 ;
        RECT 23.400 231.020 24.640 231.770 ;
        RECT 23.400 230.300 32.270 231.020 ;
        RECT 23.400 230.070 26.600 230.300 ;
        RECT 23.400 230.040 24.640 230.070 ;
        RECT 23.400 229.870 24.210 230.040 ;
        RECT 24.490 228.920 25.480 228.930 ;
        RECT 24.090 228.400 25.480 228.920 ;
        RECT 24.090 224.790 24.580 228.400 ;
        RECT 27.290 227.870 30.710 227.920 ;
        RECT 27.280 227.300 30.720 227.870 ;
        RECT 25.870 218.850 30.170 226.530 ;
        RECT 31.850 226.480 32.570 227.030 ;
        RECT 31.850 226.470 32.350 226.480 ;
        RECT 41.040 218.850 43.290 218.910 ;
        RECT 10.330 215.620 43.290 218.850 ;
        RECT 22.360 215.360 32.770 215.620 ;
        RECT 41.040 215.540 43.290 215.620 ;
        RECT 22.520 215.350 32.770 215.360 ;
        RECT 23.470 215.000 32.770 215.350 ;
        RECT 23.840 213.560 32.770 215.000 ;
        RECT 21.900 209.010 22.490 212.620 ;
        RECT 21.900 208.720 23.840 209.010 ;
        RECT 23.390 203.820 24.200 205.170 ;
        RECT 25.300 203.850 30.450 213.560 ;
        RECT 32.000 213.540 32.770 213.560 ;
        RECT 35.050 206.090 35.690 210.030 ;
        RECT 23.390 203.760 24.640 203.820 ;
        RECT 23.390 203.180 24.660 203.760 ;
        RECT 25.310 203.180 30.450 203.850 ;
        RECT 23.390 202.430 24.640 203.180 ;
        RECT 23.390 201.710 32.270 202.430 ;
        RECT 23.390 201.480 26.600 201.710 ;
        RECT 23.390 201.450 24.640 201.480 ;
        RECT 23.390 201.270 24.200 201.450 ;
        RECT 24.490 200.330 25.480 200.340 ;
        RECT 24.090 199.810 25.480 200.330 ;
        RECT 24.090 196.200 24.580 199.810 ;
        RECT 27.290 199.280 30.710 199.330 ;
        RECT 27.280 198.710 30.720 199.280 ;
        RECT 25.870 190.260 30.170 197.940 ;
        RECT 31.850 197.890 32.570 198.440 ;
        RECT 31.850 197.880 32.350 197.890 ;
        RECT 45.360 190.260 47.610 190.370 ;
        RECT 10.330 187.030 47.760 190.260 ;
        RECT 22.360 186.770 32.770 187.030 ;
        RECT 45.360 186.920 47.610 187.030 ;
        RECT 22.520 186.760 32.770 186.770 ;
        RECT 23.470 186.410 32.770 186.760 ;
        RECT 23.840 184.970 32.770 186.410 ;
        RECT 21.900 180.420 22.490 184.030 ;
        RECT 21.900 180.130 23.840 180.420 ;
        RECT 23.390 175.230 24.200 176.580 ;
        RECT 25.300 175.260 30.450 184.970 ;
        RECT 32.000 184.950 32.770 184.970 ;
        RECT 35.040 177.520 35.680 181.460 ;
        RECT 23.390 175.170 24.640 175.230 ;
        RECT 23.390 174.590 24.660 175.170 ;
        RECT 25.310 174.590 30.450 175.260 ;
        RECT 23.390 173.840 24.640 174.590 ;
        RECT 23.390 173.120 32.270 173.840 ;
        RECT 23.390 172.890 26.600 173.120 ;
        RECT 23.390 172.860 24.640 172.890 ;
        RECT 23.390 172.680 24.200 172.860 ;
        RECT 24.490 171.740 25.480 171.750 ;
        RECT 24.090 171.220 25.480 171.740 ;
        RECT 24.090 167.610 24.580 171.220 ;
        RECT 27.290 170.690 30.710 170.740 ;
        RECT 27.280 170.120 30.720 170.690 ;
        RECT 25.870 161.670 30.170 169.350 ;
        RECT 31.850 169.300 32.570 169.850 ;
        RECT 31.850 169.290 32.350 169.300 ;
        RECT 264.240 165.070 268.660 326.370 ;
        RECT 343.340 303.900 345.700 304.030 ;
        RECT 343.340 300.670 362.570 303.900 ;
        RECT 343.340 300.570 345.700 300.670 ;
        RECT 390.140 285.380 391.130 285.390 ;
        RECT 390.140 284.860 391.530 285.380 ;
        RECT 384.910 284.330 388.330 284.380 ;
        RECT 384.900 283.760 388.340 284.330 ;
        RECT 383.050 282.940 383.770 283.490 ;
        RECT 383.270 282.930 383.770 282.940 ;
        RECT 339.330 275.310 341.610 275.470 ;
        RECT 339.330 272.080 362.550 275.310 ;
        RECT 382.850 273.930 383.620 273.950 ;
        RECT 385.450 273.930 389.750 282.990 ;
        RECT 391.040 281.250 391.530 284.860 ;
        RECT 382.850 272.180 392.150 273.930 ;
        RECT 382.850 272.170 393.100 272.180 ;
        RECT 339.330 271.970 341.610 272.080 ;
        RECT 382.850 271.820 393.260 272.170 ;
        RECT 382.850 271.810 393.100 271.820 ;
        RECT 382.850 271.460 392.150 271.810 ;
        RECT 382.850 270.020 391.780 271.460 ;
        RECT 382.850 270.000 383.620 270.020 ;
        RECT 379.870 262.560 380.580 266.520 ;
        RECT 385.170 260.310 390.320 270.020 ;
        RECT 393.130 265.470 393.720 269.080 ;
        RECT 391.780 265.180 393.720 265.470 ;
        RECT 385.170 259.640 390.310 260.310 ;
        RECT 391.420 260.280 392.140 261.630 ;
        RECT 390.980 260.220 392.140 260.280 ;
        RECT 390.960 259.640 392.140 260.220 ;
        RECT 390.980 258.890 392.140 259.640 ;
        RECT 383.350 258.170 392.140 258.890 ;
        RECT 389.020 257.940 392.140 258.170 ;
        RECT 390.980 257.910 392.140 257.940 ;
        RECT 391.420 257.740 392.140 257.910 ;
        RECT 390.140 256.790 391.130 256.800 ;
        RECT 390.140 256.270 391.530 256.790 ;
        RECT 384.910 255.740 388.330 255.790 ;
        RECT 384.900 255.170 388.340 255.740 ;
        RECT 383.050 254.350 383.770 254.900 ;
        RECT 383.270 254.340 383.770 254.350 ;
        RECT 335.030 246.720 337.450 246.840 ;
        RECT 335.030 243.490 362.550 246.720 ;
        RECT 382.850 245.340 383.620 245.360 ;
        RECT 385.450 245.340 389.750 254.400 ;
        RECT 391.040 252.660 391.530 256.270 ;
        RECT 382.850 243.590 392.150 245.340 ;
        RECT 382.850 243.580 393.100 243.590 ;
        RECT 335.030 243.330 337.450 243.490 ;
        RECT 382.850 243.230 393.260 243.580 ;
        RECT 382.850 243.220 393.100 243.230 ;
        RECT 382.850 242.870 392.150 243.220 ;
        RECT 382.850 241.430 391.780 242.870 ;
        RECT 382.850 241.410 383.620 241.430 ;
        RECT 379.860 233.960 380.560 237.920 ;
        RECT 385.170 231.720 390.320 241.430 ;
        RECT 393.130 236.880 393.720 240.490 ;
        RECT 391.780 236.590 393.720 236.880 ;
        RECT 385.170 231.050 390.310 231.720 ;
        RECT 391.420 231.690 392.140 233.040 ;
        RECT 390.980 231.630 392.140 231.690 ;
        RECT 390.960 231.050 392.140 231.630 ;
        RECT 390.980 230.300 392.140 231.050 ;
        RECT 383.350 229.580 392.140 230.300 ;
        RECT 389.020 229.350 392.140 229.580 ;
        RECT 390.980 229.320 392.140 229.350 ;
        RECT 391.420 229.150 392.140 229.320 ;
        RECT 390.140 228.200 391.130 228.210 ;
        RECT 390.140 227.680 391.530 228.200 ;
        RECT 384.910 227.150 388.330 227.200 ;
        RECT 384.900 226.580 388.340 227.150 ;
        RECT 383.050 225.760 383.770 226.310 ;
        RECT 383.270 225.750 383.770 225.760 ;
        RECT 331.140 218.130 333.410 218.240 ;
        RECT 331.140 214.900 362.560 218.130 ;
        RECT 382.850 216.750 383.620 216.770 ;
        RECT 385.450 216.750 389.750 225.810 ;
        RECT 391.040 224.070 391.530 227.680 ;
        RECT 382.850 215.000 392.150 216.750 ;
        RECT 382.850 214.990 393.100 215.000 ;
        RECT 331.140 214.770 333.410 214.900 ;
        RECT 382.850 214.640 393.260 214.990 ;
        RECT 382.850 214.630 393.100 214.640 ;
        RECT 382.850 214.280 392.150 214.630 ;
        RECT 382.850 212.840 391.780 214.280 ;
        RECT 382.850 212.820 383.620 212.840 ;
        RECT 379.880 205.370 380.580 209.330 ;
        RECT 385.170 203.130 390.320 212.840 ;
        RECT 393.130 208.290 393.720 211.900 ;
        RECT 391.780 208.000 393.720 208.290 ;
        RECT 385.170 202.460 390.310 203.130 ;
        RECT 391.420 203.100 392.140 204.440 ;
        RECT 390.980 203.040 392.140 203.100 ;
        RECT 390.960 202.460 392.140 203.040 ;
        RECT 390.980 201.710 392.140 202.460 ;
        RECT 383.350 200.990 392.140 201.710 ;
        RECT 389.020 200.760 392.140 200.990 ;
        RECT 390.980 200.730 392.140 200.760 ;
        RECT 391.420 200.550 392.140 200.730 ;
        RECT 390.140 199.610 391.130 199.620 ;
        RECT 390.140 199.090 391.530 199.610 ;
        RECT 384.910 198.560 388.330 198.610 ;
        RECT 384.900 197.990 388.340 198.560 ;
        RECT 383.050 197.170 383.770 197.720 ;
        RECT 383.270 197.160 383.770 197.170 ;
        RECT 326.740 189.540 329.040 189.620 ;
        RECT 326.740 186.310 362.560 189.540 ;
        RECT 382.850 188.160 383.620 188.180 ;
        RECT 385.450 188.160 389.750 197.220 ;
        RECT 391.040 195.480 391.530 199.090 ;
        RECT 382.850 186.410 392.150 188.160 ;
        RECT 382.850 186.400 393.100 186.410 ;
        RECT 326.740 186.210 329.040 186.310 ;
        RECT 382.850 186.050 393.260 186.400 ;
        RECT 382.850 186.040 393.100 186.050 ;
        RECT 382.850 185.690 392.150 186.040 ;
        RECT 382.850 184.250 391.780 185.690 ;
        RECT 382.850 184.230 383.620 184.250 ;
        RECT 379.860 176.780 380.560 180.740 ;
        RECT 385.170 174.540 390.320 184.250 ;
        RECT 393.130 179.700 393.720 183.310 ;
        RECT 391.780 179.410 393.720 179.700 ;
        RECT 385.170 173.870 390.310 174.540 ;
        RECT 391.420 174.510 392.140 175.870 ;
        RECT 390.980 174.450 392.140 174.510 ;
        RECT 390.960 173.870 392.140 174.450 ;
        RECT 390.980 173.120 392.140 173.870 ;
        RECT 383.350 172.400 392.140 173.120 ;
        RECT 389.020 172.170 392.140 172.400 ;
        RECT 390.980 172.140 392.140 172.170 ;
        RECT 391.420 171.980 392.140 172.140 ;
        RECT 390.140 171.020 391.130 171.030 ;
        RECT 390.140 170.500 391.530 171.020 ;
        RECT 384.910 169.970 388.330 170.020 ;
        RECT 384.900 169.400 388.340 169.970 ;
        RECT 383.050 168.580 383.770 169.130 ;
        RECT 383.270 168.570 383.770 168.580 ;
        RECT 49.420 161.670 51.830 161.770 ;
        RECT 10.330 158.440 51.830 161.670 ;
        RECT 263.320 161.330 268.660 165.070 ;
        RECT 263.320 160.370 268.080 161.330 ;
        RECT 22.360 158.180 32.770 158.440 ;
        RECT 49.420 158.260 51.830 158.440 ;
        RECT 382.850 159.570 383.620 159.590 ;
        RECT 385.450 159.570 389.750 168.630 ;
        RECT 391.040 166.890 391.530 170.500 ;
        RECT 22.520 158.170 32.770 158.180 ;
        RECT 23.470 157.820 32.770 158.170 ;
        RECT 23.840 156.380 32.770 157.820 ;
        RECT 21.900 151.830 22.490 155.440 ;
        RECT 21.900 151.540 23.840 151.830 ;
        RECT 23.390 146.640 24.200 147.990 ;
        RECT 25.300 146.670 30.450 156.380 ;
        RECT 32.000 156.360 32.770 156.380 ;
        RECT 382.850 157.820 392.150 159.570 ;
        RECT 382.850 157.810 393.100 157.820 ;
        RECT 382.850 157.460 393.260 157.810 ;
        RECT 382.850 157.450 393.100 157.460 ;
        RECT 382.850 157.100 392.150 157.450 ;
        RECT 382.850 155.660 391.780 157.100 ;
        RECT 382.850 155.640 383.620 155.660 ;
        RECT 35.040 148.920 35.680 152.860 ;
        RECT 379.860 148.180 380.560 152.140 ;
        RECT 23.390 146.580 24.640 146.640 ;
        RECT 23.390 146.000 24.660 146.580 ;
        RECT 25.310 146.000 30.450 146.670 ;
        RECT 23.390 145.250 24.640 146.000 ;
        RECT 385.170 145.950 390.320 155.660 ;
        RECT 393.130 151.110 393.720 154.720 ;
        RECT 391.780 150.820 393.720 151.110 ;
        RECT 385.170 145.280 390.310 145.950 ;
        RECT 391.410 145.920 392.130 147.270 ;
        RECT 390.980 145.860 392.130 145.920 ;
        RECT 390.960 145.280 392.130 145.860 ;
        RECT 23.390 144.530 32.270 145.250 ;
        RECT 390.980 144.530 392.130 145.280 ;
        RECT 23.390 144.300 26.600 144.530 ;
        RECT 23.390 144.270 24.640 144.300 ;
        RECT 23.390 144.090 24.200 144.270 ;
        RECT 383.350 143.810 392.130 144.530 ;
        RECT 389.020 143.580 392.130 143.810 ;
        RECT 390.980 143.550 392.130 143.580 ;
        RECT 391.410 143.380 392.130 143.550 ;
        RECT 24.490 143.150 25.480 143.160 ;
        RECT 24.090 142.630 25.480 143.150 ;
        RECT 24.090 139.020 24.580 142.630 ;
        RECT 390.140 142.430 391.130 142.440 ;
        RECT 27.290 142.100 30.710 142.150 ;
        RECT 27.280 141.530 30.720 142.100 ;
        RECT 390.140 141.910 391.530 142.430 ;
        RECT 384.910 141.380 388.330 141.430 ;
        RECT 25.870 133.080 30.170 140.760 ;
        RECT 31.850 140.710 32.570 141.260 ;
        RECT 384.900 140.810 388.340 141.380 ;
        RECT 31.850 140.700 32.350 140.710 ;
        RECT 383.050 139.990 383.770 140.540 ;
        RECT 383.270 139.980 383.770 139.990 ;
        RECT 53.700 133.080 56.160 133.150 ;
        RECT 10.330 129.850 56.160 133.080 ;
        RECT 22.360 129.590 32.770 129.850 ;
        RECT 53.700 129.800 56.160 129.850 ;
        RECT 382.850 130.980 383.620 131.000 ;
        RECT 385.450 130.980 389.750 140.040 ;
        RECT 391.040 138.300 391.530 141.910 ;
        RECT 22.520 129.580 32.770 129.590 ;
        RECT 23.470 129.230 32.770 129.580 ;
        RECT 23.840 127.790 32.770 129.230 ;
        RECT 21.900 123.240 22.490 126.850 ;
        RECT 21.900 122.950 23.840 123.240 ;
        RECT 23.400 118.050 24.210 119.400 ;
        RECT 25.300 118.080 30.450 127.790 ;
        RECT 32.000 127.770 32.770 127.790 ;
        RECT 382.850 129.230 392.150 130.980 ;
        RECT 382.850 129.220 393.100 129.230 ;
        RECT 382.850 128.870 393.260 129.220 ;
        RECT 382.850 128.860 393.100 128.870 ;
        RECT 382.850 128.510 392.150 128.860 ;
        RECT 382.850 127.070 391.780 128.510 ;
        RECT 382.850 127.050 383.620 127.070 ;
        RECT 35.060 120.320 35.700 124.260 ;
        RECT 379.870 119.600 380.570 123.560 ;
        RECT 23.400 117.990 24.640 118.050 ;
        RECT 23.400 117.410 24.660 117.990 ;
        RECT 25.310 117.410 30.450 118.080 ;
        RECT 23.400 116.660 24.640 117.410 ;
        RECT 385.170 117.360 390.320 127.070 ;
        RECT 393.130 122.520 393.720 126.130 ;
        RECT 391.780 122.230 393.720 122.520 ;
        RECT 385.170 116.690 390.310 117.360 ;
        RECT 391.420 117.330 392.140 118.680 ;
        RECT 390.980 117.270 392.140 117.330 ;
        RECT 390.960 116.690 392.140 117.270 ;
        RECT 23.400 115.940 32.270 116.660 ;
        RECT 390.980 115.940 392.140 116.690 ;
        RECT 23.400 115.710 26.600 115.940 ;
        RECT 23.400 115.680 24.640 115.710 ;
        RECT 23.400 115.500 24.210 115.680 ;
        RECT 383.350 115.220 392.140 115.940 ;
        RECT 389.020 114.990 392.140 115.220 ;
        RECT 390.980 114.960 392.140 114.990 ;
        RECT 391.420 114.790 392.140 114.960 ;
        RECT 24.490 114.560 25.480 114.570 ;
        RECT 24.090 114.040 25.480 114.560 ;
        RECT 24.090 110.430 24.580 114.040 ;
        RECT 390.140 113.840 391.130 113.850 ;
        RECT 27.290 113.510 30.710 113.560 ;
        RECT 27.280 112.940 30.720 113.510 ;
        RECT 390.140 113.320 391.530 113.840 ;
        RECT 384.910 112.790 388.330 112.840 ;
        RECT 25.870 104.490 30.170 112.170 ;
        RECT 31.850 112.120 32.570 112.670 ;
        RECT 384.900 112.220 388.340 112.790 ;
        RECT 31.850 112.110 32.350 112.120 ;
        RECT 383.050 111.400 383.770 111.950 ;
        RECT 383.270 111.390 383.770 111.400 ;
        RECT 58.070 104.490 60.470 104.630 ;
        RECT 10.320 101.260 60.470 104.490 ;
        RECT 22.360 101.000 32.770 101.260 ;
        RECT 58.070 101.160 60.470 101.260 ;
        RECT 382.850 102.390 383.620 102.410 ;
        RECT 385.450 102.390 389.750 111.450 ;
        RECT 391.040 109.710 391.530 113.320 ;
        RECT 22.520 100.990 32.770 101.000 ;
        RECT 23.470 100.640 32.770 100.990 ;
        RECT 23.840 99.200 32.770 100.640 ;
        RECT 21.900 94.650 22.490 98.260 ;
        RECT 21.900 94.360 23.840 94.650 ;
        RECT 23.380 89.460 24.190 90.810 ;
        RECT 25.300 89.490 30.450 99.200 ;
        RECT 32.000 99.180 32.770 99.200 ;
        RECT 382.850 100.640 392.150 102.390 ;
        RECT 382.850 100.630 393.100 100.640 ;
        RECT 382.850 100.280 393.260 100.630 ;
        RECT 382.850 100.270 393.100 100.280 ;
        RECT 382.850 99.920 392.150 100.270 ;
        RECT 382.850 98.480 391.780 99.920 ;
        RECT 382.850 98.460 383.620 98.480 ;
        RECT 35.060 91.750 35.700 95.690 ;
        RECT 379.870 91.000 380.570 94.960 ;
        RECT 23.380 89.400 24.640 89.460 ;
        RECT 23.380 88.820 24.660 89.400 ;
        RECT 25.310 88.820 30.450 89.490 ;
        RECT 23.380 88.070 24.640 88.820 ;
        RECT 385.170 88.770 390.320 98.480 ;
        RECT 393.130 93.930 393.720 97.540 ;
        RECT 391.780 93.640 393.720 93.930 ;
        RECT 385.170 88.100 390.310 88.770 ;
        RECT 391.420 88.740 392.140 90.080 ;
        RECT 390.980 88.680 392.140 88.740 ;
        RECT 390.960 88.100 392.140 88.680 ;
        RECT 23.380 87.350 32.270 88.070 ;
        RECT 390.980 87.350 392.140 88.100 ;
        RECT 23.380 87.120 26.600 87.350 ;
        RECT 23.380 87.090 24.640 87.120 ;
        RECT 23.380 86.910 24.190 87.090 ;
        RECT 383.350 86.630 392.140 87.350 ;
        RECT 389.020 86.400 392.140 86.630 ;
        RECT 390.980 86.370 392.140 86.400 ;
        RECT 391.420 86.190 392.140 86.370 ;
        RECT 62.010 75.900 64.500 75.980 ;
        RECT 10.320 72.670 64.500 75.900 ;
        RECT 62.010 72.480 64.500 72.670 ;
        RECT 66.480 47.310 68.830 47.410 ;
        RECT 10.340 44.080 68.830 47.310 ;
        RECT 66.480 43.950 68.830 44.080 ;
        RECT 70.480 18.720 73.190 18.780 ;
        RECT 10.340 15.490 73.190 18.720 ;
        RECT 70.480 15.370 73.190 15.490 ;
      LAYER via ;
        RECT 24.530 457.210 25.290 457.560 ;
        RECT 24.140 453.780 24.490 456.770 ;
        RECT 27.410 456.180 30.580 456.600 ;
        RECT 31.880 455.210 32.400 455.730 ;
        RECT 24.160 430.390 24.490 432.420 ;
        RECT 24.730 430.330 25.350 431.030 ;
        RECT 24.530 428.620 25.290 428.970 ;
        RECT 24.140 425.190 24.490 428.180 ;
        RECT 27.410 427.590 30.580 428.010 ;
        RECT 31.880 426.620 32.400 427.140 ;
        RECT 24.160 401.800 24.490 403.830 ;
        RECT 24.730 401.740 25.350 402.440 ;
        RECT 24.530 400.030 25.290 400.380 ;
        RECT 24.140 396.600 24.490 399.590 ;
        RECT 27.410 399.000 30.580 399.420 ;
        RECT 31.880 398.030 32.400 398.550 ;
        RECT 16.590 387.570 18.620 387.900 ;
        RECT 16.530 386.710 17.230 387.330 ;
        RECT 39.980 387.570 42.970 387.920 ;
        RECT 45.180 387.570 47.210 387.900 ;
        RECT 43.410 386.770 43.760 387.530 ;
        RECT 45.120 386.710 45.820 387.330 ;
        RECT 68.570 387.570 71.560 387.920 ;
        RECT 73.770 387.570 75.800 387.900 ;
        RECT 42.380 381.480 42.800 384.650 ;
        RECT 41.410 379.660 41.930 380.180 ;
        RECT 72.000 386.770 72.350 387.530 ;
        RECT 73.710 386.710 74.410 387.330 ;
        RECT 97.160 387.570 100.150 387.920 ;
        RECT 70.970 381.480 71.390 384.650 ;
        RECT 70.000 379.660 70.520 380.180 ;
        RECT 100.590 386.770 100.940 387.530 ;
        RECT 157.790 387.570 159.820 387.900 ;
        RECT 122.520 385.980 146.320 386.240 ;
        RECT 99.560 381.480 99.980 384.650 ;
        RECT 98.590 379.660 99.110 380.180 ;
        RECT 24.160 373.210 24.490 375.240 ;
        RECT 24.730 373.150 25.350 373.850 ;
        RECT 24.530 371.440 25.290 371.790 ;
        RECT 24.140 368.010 24.490 371.000 ;
        RECT 27.410 370.410 30.580 370.830 ;
        RECT 31.880 369.440 32.400 369.960 ;
        RECT 132.290 382.070 132.680 382.460 ;
        RECT 125.780 378.660 126.040 378.920 ;
        RECT 128.640 378.710 128.900 378.970 ;
        RECT 132.370 378.620 132.760 379.010 ;
        RECT 125.770 377.630 126.030 377.890 ;
        RECT 126.440 377.650 126.700 377.910 ;
        RECT 127.180 377.640 127.440 377.900 ;
        RECT 125.770 377.180 126.030 377.440 ;
        RECT 127.180 377.200 127.440 377.460 ;
        RECT 86.320 370.730 89.550 372.980 ;
        RECT 98.510 369.450 99.030 369.820 ;
        RECT 57.730 366.240 60.960 368.490 ;
        RECT 27.310 361.970 29.560 365.200 ;
        RECT 15.780 358.570 17.640 361.800 ;
        RECT 125.770 376.760 126.030 377.020 ;
        RECT 126.440 376.810 126.700 377.070 ;
        RECT 127.200 376.780 127.460 377.040 ;
        RECT 125.770 375.410 126.030 375.670 ;
        RECT 128.330 377.330 128.590 377.590 ;
        RECT 128.140 374.910 128.400 375.170 ;
        RECT 133.750 377.450 134.010 377.710 ;
        RECT 157.730 386.710 158.430 387.330 ;
        RECT 181.180 387.570 184.170 387.920 ;
        RECT 186.380 387.570 188.410 387.900 ;
        RECT 184.610 386.770 184.960 387.530 ;
        RECT 186.320 386.710 187.020 387.330 ;
        RECT 209.770 387.570 212.760 387.920 ;
        RECT 214.970 387.570 217.000 387.900 ;
        RECT 155.200 385.980 176.060 386.240 ;
        RECT 141.830 376.910 142.090 377.170 ;
        RECT 143.190 376.990 143.450 377.250 ;
        RECT 143.880 376.980 144.140 377.240 ;
        RECT 133.670 374.750 134.090 375.170 ;
        RECT 126.420 374.010 126.680 374.270 ;
        RECT 127.850 374.030 128.110 374.290 ;
        RECT 125.630 373.430 125.890 373.690 ;
        RECT 126.560 373.430 126.820 373.690 ;
        RECT 127.260 373.430 127.520 373.690 ;
        RECT 128.000 373.430 128.260 373.690 ;
        RECT 128.710 373.420 128.970 373.680 ;
        RECT 101.850 365.070 102.260 365.480 ;
        RECT 98.370 361.130 98.890 361.650 ;
        RECT 24.160 344.620 24.490 346.650 ;
        RECT 24.730 344.560 25.350 345.260 ;
        RECT 24.530 342.850 25.290 343.200 ;
        RECT 24.140 339.420 24.490 342.410 ;
        RECT 27.410 341.820 30.580 342.240 ;
        RECT 31.880 340.850 32.400 341.370 ;
        RECT 23.830 329.980 25.910 333.210 ;
        RECT 101.900 360.280 102.310 360.690 ;
        RECT 98.470 325.110 98.990 325.630 ;
        RECT 101.900 324.170 102.310 324.610 ;
        RECT 139.620 373.350 139.910 373.930 ;
        RECT 141.110 373.250 141.370 373.510 ;
        RECT 150.970 373.270 151.230 373.530 ;
        RECT 152.910 372.290 153.170 372.550 ;
        RECT 147.330 368.610 147.590 368.870 ;
        RECT 148.420 368.620 148.680 368.880 ;
        RECT 145.790 367.700 146.050 367.960 ;
        RECT 147.340 367.620 147.600 367.880 ;
        RECT 145.770 366.780 146.030 367.040 ;
        RECT 145.750 365.790 146.010 366.050 ;
        RECT 147.340 366.630 147.600 366.890 ;
        RECT 146.830 366.040 147.090 366.300 ;
        RECT 147.250 365.900 147.510 366.160 ;
        RECT 146.800 365.120 147.060 365.380 ;
        RECT 147.340 365.200 147.600 365.460 ;
        RECT 147.250 364.910 147.510 365.170 ;
        RECT 146.810 364.200 147.070 364.460 ;
        RECT 147.340 364.210 147.600 364.470 ;
        RECT 146.160 363.180 146.420 363.440 ;
        RECT 146.120 362.220 146.380 362.480 ;
        RECT 146.160 361.260 146.420 361.520 ;
        RECT 147.250 363.920 147.510 364.180 ;
        RECT 148.430 367.630 148.690 367.890 ;
        RECT 147.340 363.220 147.600 363.480 ;
        RECT 148.430 366.640 148.690 366.900 ;
        RECT 158.700 371.860 159.010 372.170 ;
        RECT 183.580 381.480 184.000 384.650 ;
        RECT 175.280 379.500 175.700 379.920 ;
        RECT 182.610 379.660 183.130 380.180 ;
        RECT 171.430 378.740 171.850 379.160 ;
        RECT 176.950 377.130 177.390 377.570 ;
        RECT 182.670 377.130 183.110 377.570 ;
        RECT 213.200 386.770 213.550 387.530 ;
        RECT 214.910 386.710 215.610 387.330 ;
        RECT 238.360 387.570 241.350 387.920 ;
        RECT 243.560 387.570 245.590 387.900 ;
        RECT 241.790 386.770 242.140 387.530 ;
        RECT 243.500 386.710 244.200 387.330 ;
        RECT 266.950 387.570 269.940 387.920 ;
        RECT 272.150 387.570 274.180 387.900 ;
        RECT 184.490 377.100 184.930 377.540 ;
        RECT 172.530 376.110 172.970 376.550 ;
        RECT 169.770 373.090 170.030 373.350 ;
        RECT 162.700 372.400 162.960 372.660 ;
        RECT 161.530 371.410 161.800 371.670 ;
        RECT 150.200 370.630 150.550 370.980 ;
        RECT 155.450 370.940 155.710 371.200 ;
        RECT 171.380 371.070 171.640 371.330 ;
        RECT 171.380 369.320 171.640 369.580 ;
        RECT 173.480 371.910 173.740 372.170 ;
        RECT 174.420 371.430 174.680 371.690 ;
        RECT 175.460 371.470 175.720 371.730 ;
        RECT 175.520 371.190 175.780 371.450 ;
        RECT 173.480 370.160 173.740 370.420 ;
        RECT 174.420 369.680 174.680 369.940 ;
        RECT 175.460 369.720 175.720 369.980 ;
        RECT 175.520 369.440 175.780 369.700 ;
        RECT 151.220 368.390 151.480 368.780 ;
        RECT 167.620 368.400 167.950 368.660 ;
        RECT 150.580 367.570 150.840 367.970 ;
        RECT 150.600 366.460 150.860 366.720 ;
        RECT 148.550 365.800 148.810 366.060 ;
        RECT 150.600 365.540 150.860 365.800 ;
        RECT 148.550 364.810 148.810 365.070 ;
        RECT 150.570 364.620 150.830 364.880 ;
        RECT 148.550 363.820 148.810 364.080 ;
        RECT 146.120 345.980 146.380 346.450 ;
        RECT 146.760 345.980 147.020 346.450 ;
        RECT 144.760 344.950 145.020 345.210 ;
        RECT 144.240 344.550 144.500 344.810 ;
        RECT 134.960 343.300 135.620 343.960 ;
        RECT 146.840 344.930 147.100 345.190 ;
        RECT 148.600 344.940 148.870 345.210 ;
        RECT 146.180 344.570 146.440 344.830 ;
        RECT 144.260 340.640 144.520 340.900 ;
        RECT 140.170 338.780 140.540 339.150 ;
        RECT 135.000 337.440 135.660 338.100 ;
        RECT 144.120 337.400 144.380 337.660 ;
        RECT 149.100 344.550 149.360 344.810 ;
        RECT 147.430 337.840 147.690 338.100 ;
        RECT 145.220 337.410 145.480 337.670 ;
        RECT 146.310 337.410 146.570 337.670 ;
        RECT 147.440 337.370 147.700 337.630 ;
        RECT 144.670 336.730 144.930 336.990 ;
        RECT 145.770 336.730 146.030 336.990 ;
        RECT 146.870 336.730 147.130 336.990 ;
        RECT 144.670 335.360 144.930 335.620 ;
        RECT 145.770 335.360 146.030 335.620 ;
        RECT 146.870 335.360 147.130 335.620 ;
        RECT 144.120 334.630 144.380 334.890 ;
        RECT 145.220 334.630 145.480 334.890 ;
        RECT 146.310 334.630 146.570 334.890 ;
        RECT 144.110 333.290 144.370 333.550 ;
        RECT 145.220 333.280 145.480 333.540 ;
        RECT 146.310 333.260 146.570 333.520 ;
        RECT 140.160 332.540 140.530 332.910 ;
        RECT 144.670 332.590 144.930 332.850 ;
        RECT 145.770 332.580 146.030 332.840 ;
        RECT 146.860 332.580 147.120 332.840 ;
        RECT 147.700 332.120 147.960 332.480 ;
        RECT 143.150 326.880 143.440 327.170 ;
        RECT 147.470 330.280 147.730 330.540 ;
        RECT 144.160 329.840 144.420 330.100 ;
        RECT 145.260 329.850 145.520 330.110 ;
        RECT 146.350 329.850 146.610 330.110 ;
        RECT 147.480 329.810 147.740 330.070 ;
        RECT 144.710 329.170 144.970 329.430 ;
        RECT 145.810 329.170 146.070 329.430 ;
        RECT 146.910 329.170 147.170 329.430 ;
        RECT 144.710 327.800 144.970 328.060 ;
        RECT 145.810 327.800 146.070 328.060 ;
        RECT 146.910 327.800 147.170 328.060 ;
        RECT 144.160 327.070 144.420 327.330 ;
        RECT 145.260 327.070 145.520 327.330 ;
        RECT 146.350 327.070 146.610 327.330 ;
        RECT 166.990 366.680 167.320 367.010 ;
        RECT 166.420 365.200 166.750 365.530 ;
        RECT 151.210 363.530 151.470 363.790 ;
        RECT 165.780 363.600 166.110 363.930 ;
        RECT 165.140 363.030 165.470 363.360 ;
        RECT 151.220 362.570 151.480 362.830 ;
        RECT 151.210 361.610 151.470 361.870 ;
        RECT 150.570 343.950 150.830 344.210 ;
        RECT 149.950 342.800 150.210 343.060 ;
        RECT 150.520 342.190 150.780 342.450 ;
        RECT 150.020 340.890 150.280 341.150 ;
        RECT 149.530 340.190 149.790 340.450 ;
        RECT 150.020 339.340 150.280 339.600 ;
        RECT 164.530 361.460 164.860 361.790 ;
        RECT 163.900 359.930 164.230 360.260 ;
        RECT 163.340 358.360 163.670 358.690 ;
        RECT 162.720 352.890 163.050 353.220 ;
        RECT 162.090 351.300 162.420 351.630 ;
        RECT 161.470 349.750 161.800 350.080 ;
        RECT 160.870 348.270 161.200 348.600 ;
        RECT 160.230 343.100 160.560 343.430 ;
        RECT 151.740 342.630 152.000 342.890 ;
        RECT 152.390 342.630 152.650 342.890 ;
        RECT 151.220 342.190 151.480 342.450 ;
        RECT 152.760 341.610 153.020 341.870 ;
        RECT 159.560 341.530 159.890 341.860 ;
        RECT 152.420 340.390 152.680 340.650 ;
        RECT 151.210 339.620 151.470 339.880 ;
        RECT 152.430 339.850 152.690 340.110 ;
        RECT 158.940 339.890 159.270 340.220 ;
        RECT 150.550 338.310 150.810 338.570 ;
        RECT 152.740 338.990 153.000 339.250 ;
        RECT 151.240 338.300 151.500 338.560 ;
        RECT 158.260 338.450 158.590 338.780 ;
        RECT 149.970 334.500 150.230 334.920 ;
        RECT 149.930 332.120 150.190 332.480 ;
        RECT 150.550 328.490 150.810 328.820 ;
        RECT 149.520 326.870 149.810 327.160 ;
        RECT 144.150 325.730 144.410 325.990 ;
        RECT 145.260 325.720 145.520 325.980 ;
        RECT 146.350 325.700 146.610 325.960 ;
        RECT 148.360 325.860 148.960 326.460 ;
        RECT 144.710 325.030 144.970 325.290 ;
        RECT 145.810 325.020 146.070 325.280 ;
        RECT 146.900 325.020 147.160 325.280 ;
        RECT 151.720 337.530 151.980 337.790 ;
        RECT 152.430 337.470 152.690 337.730 ;
        RECT 154.220 334.090 154.800 334.800 ;
        RECT 151.140 320.930 151.400 321.270 ;
        RECT 132.230 319.990 132.620 320.380 ;
        RECT 24.160 316.030 24.490 318.060 ;
        RECT 24.730 315.970 25.350 316.670 ;
        RECT 158.230 314.620 158.660 315.050 ;
        RECT 24.530 314.260 25.290 314.610 ;
        RECT 24.140 310.830 24.490 313.820 ;
        RECT 158.880 313.830 159.310 314.260 ;
        RECT 27.410 313.230 30.580 313.650 ;
        RECT 159.550 313.150 159.950 313.550 ;
        RECT 31.880 312.260 32.400 312.780 ;
        RECT 159.380 312.210 159.890 312.720 ;
        RECT 171.380 367.570 171.640 367.830 ;
        RECT 173.480 368.410 173.740 368.670 ;
        RECT 174.420 367.930 174.680 368.190 ;
        RECT 175.460 367.970 175.720 368.230 ;
        RECT 175.520 367.690 175.780 367.950 ;
        RECT 171.380 365.820 171.640 366.080 ;
        RECT 173.480 366.660 173.740 366.920 ;
        RECT 174.420 366.180 174.680 366.440 ;
        RECT 175.460 366.220 175.720 366.480 ;
        RECT 175.520 365.940 175.780 366.200 ;
        RECT 178.240 376.110 178.680 376.550 ;
        RECT 195.050 378.740 196.400 379.160 ;
        RECT 189.630 376.100 190.580 376.510 ;
        RECT 192.640 376.110 193.080 376.550 ;
        RECT 186.890 372.330 187.150 372.590 ;
        RECT 185.010 368.800 185.270 369.060 ;
        RECT 190.480 371.420 190.740 371.680 ;
        RECT 187.350 370.400 187.610 370.660 ;
        RECT 187.770 368.310 188.030 368.570 ;
        RECT 188.830 367.830 189.090 368.090 ;
        RECT 193.650 372.340 193.910 372.600 ;
        RECT 193.210 371.430 193.470 371.690 ;
        RECT 187.320 362.520 187.580 362.780 ;
        RECT 171.380 361.050 171.640 361.310 ;
        RECT 174.420 360.690 174.680 360.950 ;
        RECT 173.480 360.210 173.740 360.470 ;
        RECT 175.520 360.930 175.780 361.190 ;
        RECT 175.460 360.650 175.720 360.910 ;
        RECT 171.380 359.300 171.640 359.560 ;
        RECT 174.420 358.940 174.680 359.200 ;
        RECT 173.480 358.460 173.740 358.720 ;
        RECT 175.520 359.180 175.780 359.440 ;
        RECT 175.460 358.900 175.720 359.160 ;
        RECT 171.380 357.550 171.640 357.810 ;
        RECT 171.380 355.800 171.640 356.060 ;
        RECT 174.420 357.190 174.680 357.450 ;
        RECT 173.480 356.710 173.740 356.970 ;
        RECT 175.520 357.430 175.780 357.690 ;
        RECT 175.460 357.150 175.720 357.410 ;
        RECT 174.420 355.440 174.680 355.700 ;
        RECT 173.480 354.960 173.740 355.220 ;
        RECT 175.520 355.680 175.780 355.940 ;
        RECT 175.460 355.400 175.720 355.660 ;
        RECT 186.230 362.000 186.490 362.260 ;
        RECT 186.230 361.630 186.490 361.890 ;
        RECT 187.320 361.110 187.580 361.370 ;
        RECT 189.730 362.520 189.990 362.780 ;
        RECT 189.730 361.110 189.990 361.370 ;
        RECT 190.470 360.730 190.740 361.000 ;
        RECT 187.320 359.320 187.580 359.580 ;
        RECT 186.230 358.800 186.490 359.060 ;
        RECT 186.230 358.430 186.490 358.690 ;
        RECT 187.320 357.910 187.580 358.170 ;
        RECT 189.730 359.320 189.990 359.580 ;
        RECT 189.730 357.910 189.990 358.170 ;
        RECT 198.440 376.070 198.880 376.510 ;
        RECT 206.770 377.100 207.050 377.540 ;
        RECT 202.990 370.440 204.210 370.700 ;
        RECT 199.750 369.790 200.010 370.050 ;
        RECT 206.080 369.250 206.340 369.510 ;
        RECT 208.420 372.340 208.680 372.600 ;
        RECT 207.530 371.470 207.790 371.730 ;
        RECT 212.170 381.480 212.590 384.650 ;
        RECT 214.940 381.440 215.310 381.810 ;
        RECT 211.200 379.660 211.720 380.180 ;
        RECT 212.630 378.230 212.890 378.490 ;
        RECT 211.090 373.050 211.350 373.320 ;
        RECT 212.630 372.660 212.890 372.920 ;
        RECT 212.880 372.200 213.140 372.460 ;
        RECT 207.530 367.260 207.790 367.520 ;
        RECT 208.550 367.270 208.810 367.530 ;
        RECT 211.300 367.150 211.730 367.580 ;
        RECT 212.880 366.630 213.140 366.890 ;
        RECT 205.050 357.510 205.310 357.770 ;
        RECT 215.760 377.980 216.130 378.350 ;
        RECT 216.860 376.430 217.120 376.690 ;
        RECT 216.200 375.550 216.460 375.810 ;
        RECT 216.850 374.740 217.110 375.000 ;
        RECT 216.530 373.270 216.900 373.640 ;
        RECT 217.350 370.970 217.610 371.230 ;
        RECT 219.860 370.660 220.360 371.160 ;
        RECT 220.810 371.150 221.310 371.650 ;
        RECT 221.890 371.620 222.390 372.120 ;
        RECT 216.460 369.810 216.720 370.070 ;
        RECT 216.460 369.210 216.720 369.470 ;
        RECT 205.050 356.960 205.310 357.220 ;
        RECT 187.110 354.090 187.390 354.370 ;
        RECT 205.050 354.850 205.310 355.110 ;
        RECT 205.050 354.270 205.310 354.560 ;
        RECT 204.460 353.520 204.720 353.780 ;
        RECT 205.050 353.720 205.310 353.980 ;
        RECT 208.770 353.000 209.030 353.080 ;
        RECT 208.770 352.820 209.260 353.000 ;
        RECT 214.950 354.070 215.320 354.440 ;
        RECT 215.720 353.480 216.090 353.850 ;
        RECT 187.300 352.050 187.560 352.310 ;
        RECT 171.380 350.920 171.640 351.180 ;
        RECT 174.420 350.560 174.680 350.820 ;
        RECT 173.480 350.080 173.740 350.340 ;
        RECT 175.520 350.800 175.780 351.060 ;
        RECT 175.460 350.520 175.720 350.780 ;
        RECT 171.380 349.170 171.640 349.430 ;
        RECT 174.420 348.810 174.680 349.070 ;
        RECT 173.480 348.330 173.740 348.590 ;
        RECT 175.520 349.050 175.780 349.310 ;
        RECT 175.460 348.770 175.720 349.030 ;
        RECT 171.380 347.420 171.640 347.680 ;
        RECT 174.420 347.060 174.680 347.320 ;
        RECT 173.480 346.580 173.740 346.840 ;
        RECT 171.380 345.670 171.640 345.930 ;
        RECT 175.520 347.300 175.780 347.560 ;
        RECT 175.460 347.020 175.720 347.280 ;
        RECT 174.420 345.310 174.680 345.570 ;
        RECT 173.480 344.830 173.740 345.090 ;
        RECT 175.520 345.550 175.780 345.810 ;
        RECT 175.460 345.270 175.720 345.530 ;
        RECT 186.210 351.530 186.470 351.790 ;
        RECT 186.210 351.160 186.470 351.420 ;
        RECT 187.300 350.640 187.560 350.900 ;
        RECT 189.710 352.050 189.970 352.310 ;
        RECT 189.710 350.640 189.970 350.900 ;
        RECT 187.300 348.850 187.560 349.110 ;
        RECT 186.210 348.330 186.470 348.590 ;
        RECT 186.210 347.960 186.470 348.220 ;
        RECT 179.740 345.900 180.000 346.310 ;
        RECT 187.300 347.440 187.560 347.700 ;
        RECT 189.710 348.850 189.970 349.110 ;
        RECT 189.710 347.440 189.970 347.700 ;
        RECT 171.340 341.860 171.600 342.120 ;
        RECT 174.380 341.500 174.640 341.760 ;
        RECT 173.440 341.020 173.700 341.280 ;
        RECT 175.480 341.740 175.740 342.000 ;
        RECT 175.420 341.460 175.680 341.720 ;
        RECT 171.340 340.110 171.600 340.370 ;
        RECT 174.380 339.750 174.640 340.010 ;
        RECT 173.440 339.270 173.700 339.530 ;
        RECT 175.480 339.990 175.740 340.250 ;
        RECT 175.420 339.710 175.680 339.970 ;
        RECT 171.340 338.360 171.600 338.620 ;
        RECT 174.380 338.000 174.640 338.260 ;
        RECT 171.340 336.610 171.600 336.870 ;
        RECT 173.440 337.520 173.700 337.780 ;
        RECT 175.480 338.240 175.740 338.500 ;
        RECT 175.420 337.960 175.680 338.220 ;
        RECT 172.580 336.170 172.890 336.480 ;
        RECT 174.380 336.250 174.640 336.510 ;
        RECT 173.440 335.770 173.700 336.030 ;
        RECT 175.480 336.490 175.740 336.750 ;
        RECT 175.420 336.210 175.680 336.470 ;
        RECT 187.330 342.780 187.590 343.040 ;
        RECT 184.140 342.180 184.400 342.440 ;
        RECT 186.240 342.260 186.500 342.520 ;
        RECT 177.560 337.050 177.820 337.310 ;
        RECT 177.020 336.680 177.310 336.970 ;
        RECT 186.240 341.890 186.500 342.150 ;
        RECT 187.330 341.370 187.590 341.630 ;
        RECT 189.740 342.780 190.000 343.040 ;
        RECT 189.740 341.370 190.000 341.630 ;
        RECT 209.000 352.740 209.260 352.820 ;
        RECT 212.930 352.700 213.190 352.960 ;
        RECT 205.050 351.620 205.310 351.880 ;
        RECT 205.050 351.070 205.310 351.330 ;
        RECT 217.410 368.470 217.780 368.570 ;
        RECT 217.350 368.210 217.780 368.470 ;
        RECT 217.410 368.200 217.780 368.210 ;
        RECT 216.460 351.150 216.830 351.520 ;
        RECT 205.650 348.670 205.910 348.930 ;
        RECT 205.650 348.120 205.910 348.380 ;
        RECT 205.650 346.030 205.910 346.290 ;
        RECT 205.650 345.430 205.910 345.740 ;
        RECT 205.650 344.880 205.910 345.140 ;
        RECT 209.720 343.820 209.980 344.080 ;
        RECT 204.020 342.160 204.280 342.420 ;
        RECT 205.650 342.780 205.910 343.040 ;
        RECT 205.650 342.230 205.910 342.490 ;
        RECT 208.730 342.150 208.990 342.410 ;
        RECT 212.020 343.700 212.280 343.960 ;
        RECT 213.740 343.800 214.010 344.060 ;
        RECT 212.000 342.650 212.260 342.910 ;
        RECT 219.680 367.960 219.940 368.220 ;
        RECT 217.390 345.900 217.760 346.310 ;
        RECT 203.500 341.230 203.760 341.490 ;
        RECT 184.770 339.400 185.030 339.660 ;
        RECT 184.170 337.090 184.430 337.350 ;
        RECT 185.200 337.080 185.460 337.340 ;
        RECT 182.770 336.680 183.030 336.940 ;
        RECT 184.740 336.760 185.000 337.020 ;
        RECT 176.390 335.460 176.810 335.880 ;
        RECT 172.540 334.500 172.960 334.920 ;
        RECT 178.450 336.140 178.710 336.400 ;
        RECT 187.330 339.580 187.590 339.840 ;
        RECT 186.240 339.060 186.500 339.320 ;
        RECT 186.240 338.690 186.500 338.950 ;
        RECT 187.330 338.170 187.590 338.430 ;
        RECT 189.740 339.580 190.000 339.840 ;
        RECT 189.740 338.170 190.000 338.430 ;
        RECT 203.030 339.390 203.290 339.650 ;
        RECT 202.530 338.460 202.790 338.720 ;
        RECT 186.980 336.700 187.240 336.960 ;
        RECT 185.780 335.450 186.110 335.780 ;
        RECT 195.820 337.010 196.170 337.360 ;
        RECT 188.970 336.280 189.230 336.540 ;
        RECT 193.010 336.250 193.280 336.520 ;
        RECT 186.930 335.380 187.270 335.720 ;
        RECT 195.860 335.240 196.120 335.560 ;
        RECT 201.850 335.460 202.110 335.800 ;
        RECT 177.070 334.410 177.390 334.730 ;
        RECT 197.280 334.530 197.660 334.910 ;
        RECT 177.360 331.430 177.620 331.690 ;
        RECT 178.450 331.430 178.710 331.690 ;
        RECT 179.550 331.420 179.810 331.680 ;
        RECT 177.910 330.750 178.170 331.010 ;
        RECT 179.000 330.730 179.260 330.990 ;
        RECT 180.110 330.720 180.370 330.980 ;
        RECT 183.390 331.420 183.650 331.680 ;
        RECT 184.490 331.430 184.750 331.690 ;
        RECT 185.580 331.430 185.840 331.690 ;
        RECT 187.170 331.460 187.430 331.720 ;
        RECT 188.260 331.460 188.520 331.720 ;
        RECT 189.360 331.450 189.620 331.710 ;
        RECT 177.910 329.380 178.170 329.640 ;
        RECT 179.000 329.380 179.260 329.640 ;
        RECT 180.100 329.380 180.360 329.640 ;
        RECT 177.170 328.630 177.630 329.090 ;
        RECT 178.450 328.650 178.710 328.910 ;
        RECT 179.550 328.650 179.810 328.910 ;
        RECT 177.350 327.280 177.610 327.540 ;
        RECT 178.450 327.280 178.710 327.540 ;
        RECT 179.550 327.280 179.810 327.540 ;
        RECT 176.780 326.640 177.040 326.900 ;
        RECT 177.910 326.600 178.170 326.860 ;
        RECT 179.000 326.600 179.260 326.860 ;
        RECT 180.100 326.610 180.360 326.870 ;
        RECT 176.790 326.170 177.050 326.430 ;
        RECT 181.090 329.660 181.370 329.940 ;
        RECT 181.830 329.680 182.110 329.960 ;
        RECT 182.830 330.720 183.090 330.980 ;
        RECT 183.940 330.730 184.200 330.990 ;
        RECT 185.030 330.750 185.290 331.010 ;
        RECT 182.840 329.380 183.100 329.640 ;
        RECT 183.940 329.380 184.200 329.640 ;
        RECT 185.030 329.380 185.290 329.640 ;
        RECT 183.390 328.650 183.650 328.910 ;
        RECT 184.490 328.650 184.750 328.910 ;
        RECT 185.590 328.650 185.850 328.910 ;
        RECT 187.720 330.780 187.980 331.040 ;
        RECT 188.810 330.760 189.070 331.020 ;
        RECT 189.920 330.750 190.180 331.010 ;
        RECT 193.200 331.450 193.460 331.710 ;
        RECT 194.300 331.460 194.560 331.720 ;
        RECT 195.390 331.460 195.650 331.720 ;
        RECT 198.940 331.430 199.200 331.690 ;
        RECT 200.040 331.440 200.300 331.700 ;
        RECT 201.130 331.440 201.390 331.700 ;
        RECT 187.720 329.410 187.980 329.670 ;
        RECT 188.810 329.410 189.070 329.670 ;
        RECT 189.910 329.410 190.170 329.670 ;
        RECT 187.160 328.680 187.420 328.940 ;
        RECT 188.260 328.680 188.520 328.940 ;
        RECT 189.360 328.680 189.620 328.940 ;
        RECT 185.550 327.680 186.010 328.140 ;
        RECT 183.390 327.280 183.650 327.540 ;
        RECT 184.490 327.280 184.750 327.540 ;
        RECT 185.590 327.280 185.850 327.540 ;
        RECT 187.160 327.310 187.420 327.570 ;
        RECT 188.260 327.310 188.520 327.570 ;
        RECT 189.360 327.310 189.620 327.570 ;
        RECT 182.840 326.610 183.100 326.870 ;
        RECT 183.940 326.600 184.200 326.860 ;
        RECT 185.030 326.600 185.290 326.860 ;
        RECT 186.160 326.640 186.420 326.900 ;
        RECT 186.590 326.670 186.850 326.930 ;
        RECT 186.980 326.790 187.440 327.250 ;
        RECT 187.720 326.630 187.980 326.890 ;
        RECT 188.810 326.630 189.070 326.890 ;
        RECT 189.910 326.640 190.170 326.900 ;
        RECT 186.150 326.170 186.410 326.430 ;
        RECT 186.600 326.200 186.860 326.460 ;
        RECT 190.900 329.660 191.180 329.940 ;
        RECT 192.640 330.750 192.900 331.010 ;
        RECT 193.750 330.760 194.010 331.020 ;
        RECT 194.840 330.780 195.100 331.040 ;
        RECT 192.650 329.410 192.910 329.670 ;
        RECT 193.750 329.410 194.010 329.670 ;
        RECT 194.840 329.410 195.100 329.670 ;
        RECT 198.380 330.730 198.640 330.990 ;
        RECT 199.490 330.740 199.750 331.000 ;
        RECT 200.580 330.760 200.840 331.020 ;
        RECT 208.710 341.140 208.970 341.400 ;
        RECT 212.000 340.770 212.260 341.030 ;
        RECT 211.870 339.590 212.130 339.850 ;
        RECT 208.710 339.150 208.970 339.410 ;
        RECT 208.760 338.190 209.020 338.450 ;
        RECT 223.080 372.220 223.580 372.720 ;
        RECT 225.670 374.010 225.930 374.270 ;
        RECT 224.610 371.380 224.870 371.640 ;
        RECT 224.640 367.690 224.900 367.950 ;
        RECT 240.760 381.480 241.180 384.650 ;
        RECT 239.790 379.660 240.310 380.180 ;
        RECT 270.380 386.770 270.730 387.530 ;
        RECT 272.090 386.710 272.790 387.330 ;
        RECT 295.540 387.570 298.530 387.920 ;
        RECT 300.740 387.570 302.770 387.900 ;
        RECT 269.350 381.480 269.770 384.650 ;
        RECT 268.380 379.660 268.900 380.180 ;
        RECT 298.970 386.770 299.320 387.530 ;
        RECT 300.680 386.710 301.380 387.330 ;
        RECT 324.130 387.570 327.120 387.920 ;
        RECT 329.330 387.570 331.360 387.900 ;
        RECT 297.940 381.480 298.360 384.650 ;
        RECT 296.970 379.660 297.490 380.180 ;
        RECT 327.560 386.770 327.910 387.530 ;
        RECT 329.270 386.710 329.970 387.330 ;
        RECT 352.720 387.570 355.710 387.920 ;
        RECT 326.530 381.480 326.950 384.650 ;
        RECT 325.560 379.660 326.080 380.180 ;
        RECT 356.150 386.770 356.500 387.530 ;
        RECT 355.120 381.480 355.540 384.650 ;
        RECT 354.150 379.660 354.670 380.180 ;
        RECT 231.890 369.280 233.170 370.560 ;
        RECT 233.890 368.330 234.150 368.590 ;
        RECT 236.210 367.120 236.470 367.550 ;
        RECT 232.380 365.840 232.640 366.260 ;
        RECT 227.920 364.890 228.180 365.150 ;
        RECT 228.380 362.640 228.780 363.040 ;
        RECT 229.360 362.000 229.720 362.360 ;
        RECT 228.170 353.000 228.430 353.090 ;
        RECT 223.990 352.700 224.250 352.960 ;
        RECT 227.920 352.830 228.430 353.000 ;
        RECT 227.920 352.740 228.180 352.830 ;
        RECT 222.990 349.940 223.490 350.440 ;
        RECT 221.910 344.750 222.410 345.220 ;
        RECT 220.840 342.740 221.100 342.990 ;
        RECT 220.690 342.730 221.100 342.740 ;
        RECT 220.690 342.480 220.950 342.730 ;
        RECT 220.690 342.060 220.950 342.310 ;
        RECT 220.690 342.050 221.100 342.060 ;
        RECT 220.840 341.800 221.100 342.050 ;
        RECT 220.840 340.060 221.100 340.220 ;
        RECT 220.780 339.970 221.280 340.060 ;
        RECT 220.690 339.710 221.280 339.970 ;
        RECT 220.780 339.560 221.280 339.710 ;
        RECT 220.690 339.290 220.950 339.540 ;
        RECT 220.690 339.280 221.100 339.290 ;
        RECT 219.730 334.260 220.230 334.760 ;
        RECT 204.000 332.750 204.260 333.250 ;
        RECT 203.460 331.850 203.720 332.350 ;
        RECT 202.990 330.950 203.250 331.450 ;
        RECT 198.390 329.390 198.650 329.650 ;
        RECT 199.490 329.390 199.750 329.650 ;
        RECT 200.580 329.390 200.840 329.650 ;
        RECT 193.200 328.680 193.460 328.940 ;
        RECT 194.300 328.680 194.560 328.940 ;
        RECT 202.510 330.050 202.770 330.550 ;
        RECT 195.400 328.680 195.660 328.940 ;
        RECT 198.940 328.660 199.200 328.920 ;
        RECT 200.040 328.660 200.300 328.920 ;
        RECT 201.140 328.660 201.400 328.920 ;
        RECT 193.200 327.310 193.460 327.570 ;
        RECT 194.300 327.310 194.560 327.570 ;
        RECT 195.400 327.310 195.660 327.570 ;
        RECT 192.650 326.640 192.910 326.900 ;
        RECT 193.750 326.630 194.010 326.890 ;
        RECT 194.840 326.630 195.100 326.890 ;
        RECT 198.940 327.290 199.200 327.550 ;
        RECT 200.040 327.290 200.300 327.550 ;
        RECT 201.140 327.290 201.400 327.550 ;
        RECT 195.970 326.670 196.230 326.930 ;
        RECT 198.390 326.620 198.650 326.880 ;
        RECT 199.490 326.610 199.750 326.870 ;
        RECT 200.580 326.610 200.840 326.870 ;
        RECT 195.370 325.880 195.830 326.340 ;
        RECT 195.960 326.200 196.220 326.460 ;
        RECT 169.300 323.650 169.560 324.770 ;
        RECT 181.410 324.710 182.530 324.730 ;
        RECT 180.670 323.610 182.530 324.710 ;
        RECT 180.670 323.590 181.790 323.610 ;
        RECT 190.480 323.560 192.340 324.750 ;
        RECT 167.620 319.360 167.950 319.690 ;
        RECT 167.000 318.740 167.330 319.070 ;
        RECT 166.370 318.110 166.700 318.440 ;
        RECT 165.770 317.480 166.100 317.810 ;
        RECT 165.130 316.800 165.460 317.130 ;
        RECT 164.530 316.180 164.860 316.510 ;
        RECT 163.930 315.540 164.260 315.870 ;
        RECT 163.350 314.970 163.680 315.300 ;
        RECT 162.770 314.280 163.100 314.610 ;
        RECT 162.120 313.640 162.450 313.970 ;
        RECT 161.480 312.990 161.810 313.330 ;
        RECT 160.900 312.350 161.270 312.720 ;
        RECT 201.710 326.650 201.970 326.910 ;
        RECT 201.700 326.180 201.960 326.440 ;
        RECT 220.840 339.030 221.100 339.280 ;
        RECT 222.290 339.500 222.560 339.770 ;
        RECT 225.970 336.780 226.470 337.280 ;
        RECT 223.100 328.670 223.600 329.170 ;
        RECT 221.910 327.720 222.410 328.180 ;
        RECT 220.780 326.850 221.280 327.310 ;
        RECT 219.850 325.940 220.350 326.400 ;
        RECT 225.390 323.650 226.330 324.770 ;
        RECT 201.180 320.020 201.510 320.350 ;
        RECT 230.280 359.630 230.670 360.020 ;
        RECT 231.110 359.070 231.490 359.330 ;
        RECT 228.440 318.830 228.840 319.230 ;
        RECT 228.050 317.990 228.310 318.250 ;
        RECT 229.350 318.030 229.740 318.420 ;
        RECT 230.280 317.210 230.670 317.600 ;
        RECT 231.870 357.510 232.130 357.770 ;
        RECT 231.870 356.960 232.130 357.220 ;
        RECT 231.870 354.850 232.130 355.110 ;
        RECT 231.870 354.270 232.130 354.560 ;
        RECT 231.870 353.720 232.130 353.980 ;
        RECT 231.870 351.620 232.130 351.880 ;
        RECT 231.870 351.070 232.130 351.330 ;
        RECT 233.620 364.830 233.880 365.090 ;
        RECT 243.160 374.610 243.870 375.320 ;
        RECT 250.210 377.000 250.470 377.260 ;
        RECT 254.680 378.230 254.940 378.490 ;
        RECT 247.940 374.010 248.200 374.270 ;
        RECT 251.100 375.840 251.360 376.100 ;
        RECT 252.040 375.560 252.300 375.820 ;
        RECT 251.100 375.240 251.360 375.500 ;
        RECT 250.210 374.240 250.470 374.500 ;
        RECT 252.750 375.070 253.010 375.330 ;
        RECT 252.700 374.420 252.960 374.680 ;
        RECT 239.630 369.500 239.890 369.760 ;
        RECT 241.860 369.490 242.120 369.750 ;
        RECT 239.320 368.630 239.580 368.890 ;
        RECT 239.690 368.330 239.950 368.590 ;
        RECT 240.990 368.630 241.250 368.890 ;
        RECT 238.920 367.750 239.180 368.010 ;
        RECT 241.880 367.950 242.140 368.210 ;
        RECT 239.630 366.300 239.890 366.560 ;
        RECT 241.860 366.290 242.120 366.550 ;
        RECT 239.320 365.430 239.580 365.690 ;
        RECT 238.920 364.440 239.180 364.810 ;
        RECT 240.990 365.430 241.250 365.690 ;
        RECT 239.320 363.560 239.580 363.820 ;
        RECT 233.620 362.310 233.880 362.570 ;
        RECT 239.630 362.690 239.890 362.950 ;
        RECT 240.990 363.560 241.250 363.820 ;
        RECT 242.160 363.580 242.420 363.840 ;
        RECT 241.860 362.700 242.120 362.960 ;
        RECT 242.310 362.750 242.570 363.010 ;
        RECT 241.480 361.920 241.740 362.180 ;
        RECT 238.920 361.240 239.180 361.500 ;
        RECT 242.600 361.490 242.860 361.750 ;
        RECT 239.320 360.360 239.580 360.620 ;
        RECT 240.990 360.360 241.250 360.620 ;
        RECT 242.210 360.640 242.470 360.900 ;
        RECT 239.630 359.490 239.890 359.750 ;
        RECT 241.860 359.500 242.120 359.760 ;
        RECT 244.170 370.970 244.430 371.230 ;
        RECT 245.060 369.810 245.320 370.070 ;
        RECT 248.640 372.200 248.900 372.460 ;
        RECT 252.700 373.150 252.960 373.410 ;
        RECT 252.750 372.500 253.010 372.760 ;
        RECT 252.750 372.070 253.010 372.330 ;
        RECT 252.700 371.420 252.960 371.680 ;
        RECT 252.700 370.150 252.960 370.410 ;
        RECT 246.000 369.530 246.260 369.790 ;
        RECT 248.200 369.610 248.460 369.870 ;
        RECT 252.750 369.500 253.010 369.760 ;
        RECT 254.410 375.030 254.670 375.290 ;
        RECT 254.460 372.920 254.720 373.070 ;
        RECT 254.460 372.810 254.940 372.920 ;
        RECT 254.680 372.660 254.940 372.810 ;
        RECT 254.450 372.090 254.710 372.350 ;
        RECT 256.110 372.040 259.340 374.100 ;
        RECT 254.370 369.840 254.630 370.100 ;
        RECT 245.060 369.210 245.320 369.470 ;
        RECT 244.170 368.210 244.430 368.470 ;
        RECT 246.710 369.040 246.970 369.300 ;
        RECT 246.660 368.390 246.920 368.650 ;
        RECT 248.370 369.040 248.630 369.260 ;
        RECT 248.350 369.000 248.630 369.040 ;
        RECT 248.350 368.780 248.610 369.000 ;
        RECT 250.080 368.480 250.340 368.740 ;
        RECT 247.520 367.950 247.780 368.210 ;
        RECT 246.660 367.120 246.920 367.380 ;
        RECT 246.710 366.470 246.970 366.730 ;
        RECT 246.710 366.040 246.970 366.300 ;
        RECT 246.660 365.390 246.920 365.650 ;
        RECT 246.660 364.120 246.920 364.380 ;
        RECT 246.710 363.470 246.970 363.730 ;
        RECT 248.640 367.520 248.900 367.780 ;
        RECT 248.420 366.930 248.680 367.040 ;
        RECT 248.250 366.890 248.680 366.930 ;
        RECT 248.250 366.780 248.900 366.890 ;
        RECT 248.250 366.670 248.510 366.780 ;
        RECT 248.640 366.630 248.900 366.780 ;
        RECT 248.410 366.060 248.670 366.320 ;
        RECT 284.700 367.150 286.760 370.450 ;
        RECT 248.330 363.810 248.590 364.070 ;
        RECT 313.290 362.900 316.520 364.960 ;
        RECT 244.060 362.440 244.330 362.700 ;
        RECT 341.880 358.490 345.110 360.540 ;
        RECT 356.220 357.850 358.210 361.080 ;
        RECT 242.970 354.820 243.680 355.530 ;
        RECT 264.480 356.870 266.700 357.190 ;
        RECT 238.770 336.770 239.280 337.280 ;
        RECT 347.670 329.260 349.760 332.490 ;
        RECT 264.320 326.480 268.600 327.570 ;
        RECT 232.880 323.280 233.140 323.540 ;
        RECT 232.880 322.610 233.140 322.870 ;
        RECT 233.150 321.320 233.410 321.580 ;
        RECT 233.150 319.710 233.410 319.970 ;
        RECT 233.140 318.100 233.400 318.360 ;
        RECT 231.100 316.420 231.480 316.800 ;
        RECT 233.150 316.480 233.410 316.740 ;
        RECT 233.140 314.870 233.400 315.130 ;
        RECT 232.380 313.390 232.640 313.650 ;
        RECT 233.140 311.670 233.400 311.930 ;
        RECT 229.900 309.960 230.160 310.220 ;
        RECT 230.840 309.960 231.100 310.220 ;
        RECT 231.790 309.940 232.050 310.200 ;
        RECT 233.100 309.960 233.360 310.220 ;
        RECT 27.730 301.390 29.810 304.620 ;
        RECT 24.160 287.440 24.490 289.470 ;
        RECT 24.730 287.380 25.350 288.080 ;
        RECT 24.530 285.670 25.290 286.020 ;
        RECT 24.140 282.240 24.490 285.230 ;
        RECT 27.410 284.640 30.580 285.060 ;
        RECT 31.880 283.670 32.400 284.190 ;
        RECT 32.360 272.800 34.440 276.030 ;
        RECT 24.160 258.850 24.490 260.880 ;
        RECT 24.730 258.790 25.350 259.490 ;
        RECT 24.530 257.080 25.290 257.430 ;
        RECT 24.140 253.650 24.490 256.640 ;
        RECT 27.410 256.050 30.580 256.470 ;
        RECT 31.880 255.080 32.400 255.600 ;
        RECT 36.770 244.210 38.850 247.440 ;
        RECT 24.160 230.260 24.490 232.290 ;
        RECT 24.730 230.200 25.350 230.900 ;
        RECT 24.530 228.490 25.290 228.840 ;
        RECT 24.140 225.060 24.490 228.050 ;
        RECT 27.410 227.460 30.580 227.880 ;
        RECT 31.880 226.490 32.400 227.010 ;
        RECT 41.110 215.620 43.190 218.850 ;
        RECT 24.160 201.670 24.490 203.700 ;
        RECT 24.730 201.610 25.350 202.310 ;
        RECT 24.530 199.900 25.290 200.250 ;
        RECT 24.140 196.470 24.490 199.460 ;
        RECT 27.410 198.870 30.580 199.290 ;
        RECT 31.880 197.900 32.400 198.420 ;
        RECT 24.160 173.080 24.490 175.110 ;
        RECT 24.730 173.020 25.350 173.720 ;
        RECT 24.530 171.310 25.290 171.660 ;
        RECT 24.140 167.880 24.490 170.870 ;
        RECT 27.410 170.280 30.580 170.700 ;
        RECT 31.880 169.310 32.400 169.830 ;
        RECT 343.420 300.670 345.510 303.900 ;
        RECT 390.330 284.950 391.090 285.300 ;
        RECT 385.040 283.920 388.210 284.340 ;
        RECT 383.220 282.950 383.740 283.470 ;
        RECT 339.440 272.080 341.530 275.310 ;
        RECT 391.130 281.520 391.480 284.510 ;
        RECT 390.270 258.070 390.890 258.770 ;
        RECT 391.130 258.130 391.460 260.160 ;
        RECT 390.330 256.360 391.090 256.710 ;
        RECT 385.040 255.330 388.210 255.750 ;
        RECT 383.220 254.360 383.740 254.880 ;
        RECT 335.190 243.490 337.280 246.720 ;
        RECT 391.130 252.930 391.480 255.920 ;
        RECT 390.270 229.480 390.890 230.180 ;
        RECT 391.130 229.540 391.460 231.570 ;
        RECT 390.330 227.770 391.090 228.120 ;
        RECT 385.040 226.740 388.210 227.160 ;
        RECT 383.220 225.770 383.740 226.290 ;
        RECT 331.250 214.900 333.340 218.130 ;
        RECT 391.130 224.340 391.480 227.330 ;
        RECT 390.270 200.890 390.890 201.590 ;
        RECT 391.130 200.950 391.460 202.980 ;
        RECT 390.330 199.180 391.090 199.530 ;
        RECT 385.040 198.150 388.210 198.570 ;
        RECT 383.220 197.180 383.740 197.700 ;
        RECT 391.130 195.750 391.480 198.740 ;
        RECT 390.270 172.300 390.890 173.000 ;
        RECT 391.130 172.360 391.460 174.390 ;
        RECT 390.330 170.590 391.090 170.940 ;
        RECT 385.040 169.560 388.210 169.980 ;
        RECT 383.220 168.590 383.740 169.110 ;
        RECT 49.650 158.440 51.730 161.670 ;
        RECT 263.500 160.540 267.920 164.960 ;
        RECT 391.130 167.160 391.480 170.150 ;
        RECT 24.160 144.490 24.490 146.520 ;
        RECT 24.730 144.430 25.350 145.130 ;
        RECT 390.270 143.710 390.890 144.410 ;
        RECT 391.130 143.770 391.460 145.800 ;
        RECT 24.530 142.720 25.290 143.070 ;
        RECT 24.140 139.290 24.490 142.280 ;
        RECT 27.410 141.690 30.580 142.110 ;
        RECT 390.330 142.000 391.090 142.350 ;
        RECT 31.880 140.720 32.400 141.240 ;
        RECT 385.040 140.970 388.210 141.390 ;
        RECT 383.220 140.000 383.740 140.520 ;
        RECT 391.130 138.570 391.480 141.560 ;
        RECT 24.160 115.900 24.490 117.930 ;
        RECT 24.730 115.840 25.350 116.540 ;
        RECT 390.270 115.120 390.890 115.820 ;
        RECT 391.130 115.180 391.460 117.210 ;
        RECT 24.530 114.130 25.290 114.480 ;
        RECT 24.140 110.700 24.490 113.690 ;
        RECT 27.410 113.100 30.580 113.520 ;
        RECT 390.330 113.410 391.090 113.760 ;
        RECT 31.880 112.130 32.400 112.650 ;
        RECT 385.040 112.380 388.210 112.800 ;
        RECT 383.220 111.410 383.740 111.930 ;
        RECT 58.270 101.260 60.350 104.490 ;
        RECT 391.130 109.980 391.480 112.970 ;
        RECT 24.160 87.310 24.490 89.340 ;
        RECT 24.730 87.250 25.350 87.950 ;
        RECT 390.270 86.530 390.890 87.230 ;
        RECT 391.130 86.590 391.460 88.620 ;
        RECT 62.240 72.670 64.320 75.900 ;
        RECT 66.680 44.080 68.760 47.310 ;
        RECT 70.980 15.490 73.060 18.720 ;
      LAYER met2 ;
        RECT 157.130 386.670 357.260 388.070 ;
        RECT 157.600 386.660 158.530 386.670 ;
        RECT 186.190 386.660 187.120 386.670 ;
        RECT 214.780 386.660 215.710 386.670 ;
        RECT 243.370 386.660 244.300 386.670 ;
        RECT 271.960 386.660 272.890 386.670 ;
        RECT 300.550 386.660 301.480 386.670 ;
        RECT 329.140 386.660 330.070 386.670 ;
        RECT 157.850 386.340 158.020 386.660 ;
        RECT 121.700 384.950 177.170 386.340 ;
        RECT 186.440 385.550 186.610 386.660 ;
        RECT 215.030 385.550 215.200 386.660 ;
        RECT 243.620 385.550 243.790 386.660 ;
        RECT 272.210 385.550 272.380 386.660 ;
        RECT 300.800 385.550 300.970 386.660 ;
        RECT 329.390 385.550 329.560 386.660 ;
        RECT 131.030 382.380 131.710 383.600 ;
        RECT 132.260 382.380 132.710 382.480 ;
        RECT 131.030 382.150 132.710 382.380 ;
        RECT 131.030 381.280 131.710 382.150 ;
        RECT 132.260 382.050 132.710 382.150 ;
        RECT 183.470 381.770 184.110 384.780 ;
        RECT 212.060 381.770 212.700 384.780 ;
        RECT 214.880 381.810 215.340 381.830 ;
        RECT 240.650 381.810 241.290 384.780 ;
        RECT 245.750 381.810 246.610 383.160 ;
        RECT 214.880 381.770 246.610 381.810 ;
        RECT 269.240 381.770 269.880 384.780 ;
        RECT 297.830 381.770 298.470 384.780 ;
        RECT 326.420 381.770 327.060 384.780 ;
        RECT 355.010 381.770 355.650 384.780 ;
        RECT 157.130 380.370 357.260 381.770 ;
        RECT 182.570 380.240 185.200 380.370 ;
        RECT 211.160 380.240 213.790 380.370 ;
        RECT 239.750 380.240 242.380 380.370 ;
        RECT 268.340 380.240 270.970 380.370 ;
        RECT 296.930 380.240 299.560 380.370 ;
        RECT 325.520 380.240 328.150 380.370 ;
        RECT 354.110 380.240 356.740 380.370 ;
        RECT 130.880 380.180 133.360 380.190 ;
        RECT 130.880 380.050 134.830 380.180 ;
        RECT 150.810 380.090 151.560 380.100 ;
        RECT 150.810 380.050 152.430 380.090 ;
        RECT 121.700 379.150 177.170 380.050 ;
        RECT 182.570 379.730 185.120 380.240 ;
        RECT 211.160 379.730 213.710 380.240 ;
        RECT 239.750 379.730 242.300 380.240 ;
        RECT 268.340 379.730 270.890 380.240 ;
        RECT 296.930 379.730 299.480 380.240 ;
        RECT 325.520 379.730 328.070 380.240 ;
        RECT 354.110 379.730 356.660 380.240 ;
        RECT 182.570 379.660 183.190 379.730 ;
        RECT 211.160 379.660 211.780 379.730 ;
        RECT 239.750 379.660 240.370 379.730 ;
        RECT 268.340 379.660 268.960 379.730 ;
        RECT 296.930 379.660 297.550 379.730 ;
        RECT 325.520 379.660 326.140 379.730 ;
        RECT 354.110 379.660 354.730 379.730 ;
        RECT 195.020 379.150 196.440 379.190 ;
        RECT 121.700 378.750 196.490 379.150 ;
        RECT 121.700 378.650 177.170 378.750 ;
        RECT 195.020 378.710 196.440 378.750 ;
        RECT 10.450 377.250 16.200 378.650 ;
        RECT 126.130 378.580 129.020 378.650 ;
        RECT 131.030 378.190 131.710 378.650 ;
        RECT 132.360 378.580 132.790 378.650 ;
        RECT 132.360 378.570 134.300 378.580 ;
        RECT 132.450 378.350 134.300 378.570 ;
        RECT 212.610 378.520 212.920 378.530 ;
        RECT 210.440 378.340 212.920 378.520 ;
        RECT 212.610 378.200 212.920 378.340 ;
        RECT 215.710 378.350 216.150 378.370 ;
        RECT 245.750 378.350 246.610 379.030 ;
        RECT 125.740 377.630 126.060 377.890 ;
        RECT 126.420 377.620 126.730 377.950 ;
        RECT 127.150 377.640 127.470 377.900 ;
        RECT 131.030 377.870 134.390 378.190 ;
        RECT 215.710 378.100 246.610 378.350 ;
        RECT 254.650 378.520 254.960 378.530 ;
        RECT 254.650 378.340 257.130 378.520 ;
        RECT 254.650 378.200 254.960 378.340 ;
        RECT 215.200 377.920 215.280 378.100 ;
        RECT 215.710 377.980 249.960 378.100 ;
        RECT 215.710 377.960 216.150 377.980 ;
        RECT 217.610 377.920 226.720 377.980 ;
        RECT 240.840 377.920 249.960 377.980 ;
        RECT 131.030 377.720 131.710 377.870 ;
        RECT 127.900 377.590 142.550 377.720 ;
        RECT 125.230 377.510 142.550 377.590 ;
        RECT 176.920 377.540 177.420 377.570 ;
        RECT 182.640 377.540 183.140 377.570 ;
        RECT 125.230 377.340 128.040 377.510 ;
        RECT 10.450 372.530 11.850 377.250 ;
        RECT 125.230 376.830 127.900 377.340 ;
        RECT 128.300 377.300 128.620 377.510 ;
        RECT 125.740 376.760 126.060 376.830 ;
        RECT 126.420 376.780 126.730 376.830 ;
        RECT 127.170 376.780 127.490 376.830 ;
        RECT 128.410 376.000 128.680 377.280 ;
        RECT 131.030 376.750 131.710 377.510 ;
        RECT 133.720 377.480 134.300 377.510 ;
        RECT 133.720 377.450 134.040 377.480 ;
        RECT 141.970 377.210 142.210 377.510 ;
        RECT 141.810 376.880 142.210 377.210 ;
        RECT 143.170 377.280 143.480 377.290 ;
        RECT 143.170 376.960 143.590 377.280 ;
        RECT 141.970 376.840 142.210 376.880 ;
        RECT 143.290 376.820 143.590 376.960 ;
        RECT 143.860 377.270 144.170 377.280 ;
        RECT 143.860 376.950 144.320 377.270 ;
        RECT 176.920 377.130 207.080 377.540 ;
        RECT 177.070 377.100 207.080 377.130 ;
        RECT 144.020 376.810 144.320 376.950 ;
        RECT 245.750 376.930 246.610 377.920 ;
        RECT 355.840 377.320 362.510 378.720 ;
        RECT 250.180 377.080 250.490 377.300 ;
        RECT 250.180 376.970 252.370 377.080 ;
        RECT 250.340 376.860 252.370 376.970 ;
        RECT 133.030 376.380 134.560 376.540 ;
        RECT 125.890 375.990 128.680 376.000 ;
        RECT 125.230 375.770 128.680 375.990 ;
        RECT 131.220 376.050 134.560 376.380 ;
        RECT 172.500 376.530 173.000 376.550 ;
        RECT 178.240 376.530 178.680 376.580 ;
        RECT 216.840 376.560 217.150 376.730 ;
        RECT 192.610 376.530 193.110 376.550 ;
        RECT 172.500 376.110 199.010 376.530 ;
        RECT 216.840 376.400 226.720 376.560 ;
        RECT 217.010 376.370 226.720 376.400 ;
        RECT 172.650 376.090 199.010 376.110 ;
        RECT 178.240 376.080 178.680 376.090 ;
        RECT 198.410 376.070 198.910 376.090 ;
        RECT 131.220 375.980 133.490 376.050 ;
        RECT 131.220 375.780 131.620 375.980 ;
        RECT 251.070 375.840 251.390 376.100 ;
        RECT 125.230 375.760 128.160 375.770 ;
        RECT 125.740 375.600 126.060 375.670 ;
        RECT 125.230 375.410 126.060 375.600 ;
        RECT 125.230 375.280 125.850 375.410 ;
        RECT 130.870 375.380 131.620 375.780 ;
        RECT 216.170 375.550 216.490 375.810 ;
        RECT 252.010 375.740 252.330 375.820 ;
        RECT 216.560 375.640 226.720 375.680 ;
        RECT 216.550 375.450 226.720 375.640 ;
        RECT 251.020 375.560 252.330 375.740 ;
        RECT 251.020 375.390 252.200 375.560 ;
        RECT 128.110 375.120 128.420 375.200 ;
        RECT 243.130 375.170 243.900 375.320 ;
        RECT 251.070 375.240 251.390 375.390 ;
        RECT 125.230 374.890 128.420 375.120 ;
        RECT 128.110 374.870 128.420 374.890 ;
        RECT 133.640 374.750 243.900 375.170 ;
        RECT 252.720 375.080 253.030 375.370 ;
        RECT 254.380 375.080 254.690 375.330 ;
        RECT 252.000 375.000 254.690 375.080 ;
        RECT 216.830 374.710 217.140 374.750 ;
        RECT 126.400 373.980 126.710 374.310 ;
        RECT 127.830 374.000 128.140 374.330 ;
        RECT 125.230 373.620 129.110 373.950 ;
        RECT 130.580 373.930 131.260 374.600 ;
        RECT 217.000 374.510 226.720 374.700 ;
        RECT 243.130 374.610 243.900 374.750 ;
        RECT 225.640 374.170 225.960 374.290 ;
        RECT 245.720 374.170 246.580 374.940 ;
        RECT 252.000 374.850 254.540 375.000 ;
        RECT 250.180 374.320 250.490 374.540 ;
        RECT 252.230 374.320 252.560 374.490 ;
        RECT 252.670 374.390 252.980 374.720 ;
        RECT 247.910 374.170 248.230 374.290 ;
        RECT 250.180 374.280 252.560 374.320 ;
        RECT 225.640 373.990 248.230 374.170 ;
        RECT 249.010 374.040 249.320 374.280 ;
        RECT 250.180 374.210 252.370 374.280 ;
        RECT 250.330 374.110 252.370 374.210 ;
        RECT 139.500 373.930 139.970 373.950 ;
        RECT 125.230 373.530 129.120 373.620 ;
        RECT 85.760 373.240 89.850 373.490 ;
        RECT 125.230 373.460 129.110 373.530 ;
        RECT 125.610 373.400 125.920 373.460 ;
        RECT 126.540 373.400 126.850 373.460 ;
        RECT 127.240 373.400 127.550 373.460 ;
        RECT 127.980 373.400 128.290 373.460 ;
        RECT 128.430 373.390 129.000 373.460 ;
        RECT 128.430 373.280 128.870 373.390 ;
        RECT 130.580 373.350 139.970 373.930 ;
        RECT 216.490 373.640 216.910 373.660 ;
        RECT 225.440 373.640 225.520 373.810 ;
        RECT 245.720 373.640 246.580 373.990 ;
        RECT 130.580 373.280 131.300 373.350 ;
        RECT 139.500 373.330 139.970 373.350 ;
        RECT 141.090 373.280 141.400 373.550 ;
        RECT 150.950 373.280 151.260 373.570 ;
        RECT 169.750 373.320 170.050 373.380 ;
        RECT 211.070 373.320 211.370 373.350 ;
        RECT 85.760 370.990 127.730 373.240 ;
        RECT 128.140 373.070 151.370 373.280 ;
        RECT 169.750 373.090 211.440 373.320 ;
        RECT 216.490 373.270 246.580 373.640 ;
        RECT 250.120 373.410 250.340 373.430 ;
        RECT 216.490 373.250 216.910 373.270 ;
        RECT 130.580 372.280 131.260 373.070 ;
        RECT 169.750 373.060 170.050 373.090 ;
        RECT 211.070 373.010 211.370 373.090 ;
        RECT 215.200 373.050 215.280 373.230 ;
        RECT 217.510 373.220 217.670 373.240 ;
        RECT 245.720 373.220 246.580 373.270 ;
        RECT 249.900 373.220 250.060 373.240 ;
        RECT 217.510 373.170 226.720 373.220 ;
        RECT 217.630 373.070 226.720 373.170 ;
        RECT 240.840 373.170 250.060 373.220 ;
        RECT 240.840 373.070 249.940 373.170 ;
        RECT 250.070 373.070 250.340 373.410 ;
        RECT 252.230 373.340 252.560 373.550 ;
        RECT 252.670 373.110 252.980 373.440 ;
        RECT 212.610 372.810 212.920 372.950 ;
        RECT 245.720 372.840 246.580 373.070 ;
        RECT 254.430 372.950 254.740 373.110 ;
        RECT 254.960 372.950 259.760 374.900 ;
        RECT 254.430 372.940 259.760 372.950 ;
        RECT 252.260 372.810 259.760 372.940 ;
        RECT 162.670 372.660 162.980 372.680 ;
        RECT 152.880 372.580 153.200 372.590 ;
        RECT 162.670 372.580 162.990 372.660 ;
        RECT 210.440 372.630 212.920 372.810 ;
        RECT 212.610 372.620 212.920 372.630 ;
        RECT 186.850 372.590 187.170 372.610 ;
        RECT 186.850 372.580 187.180 372.590 ;
        RECT 193.620 372.580 193.940 372.610 ;
        RECT 208.390 372.580 208.710 372.600 ;
        RECT 223.050 372.580 223.610 372.720 ;
        RECT 152.880 372.350 223.610 372.580 ;
        RECT 152.880 372.270 153.200 372.350 ;
        RECT 162.670 372.340 162.980 372.350 ;
        RECT 186.850 372.330 187.180 372.350 ;
        RECT 193.620 372.330 193.940 372.350 ;
        RECT 208.390 372.340 208.710 372.350 ;
        RECT 210.690 372.310 213.170 372.350 ;
        RECT 158.670 372.130 159.040 372.190 ;
        RECT 173.480 372.130 173.740 372.200 ;
        RECT 212.860 372.170 213.170 372.310 ;
        RECT 223.050 372.210 223.610 372.350 ;
        RECT 243.260 372.280 259.810 372.810 ;
        RECT 221.870 372.130 222.410 372.150 ;
        RECT 158.670 372.070 222.410 372.130 ;
        RECT 236.950 372.080 259.810 372.280 ;
        RECT 243.260 372.070 259.810 372.080 ;
        RECT 158.670 371.900 226.980 372.070 ;
        RECT 130.580 371.780 131.090 371.900 ;
        RECT 158.670 371.840 159.040 371.900 ;
        RECT 130.580 371.490 133.680 371.780 ;
        RECT 131.090 371.480 133.680 371.490 ;
        RECT 161.500 371.670 161.810 371.680 ;
        RECT 173.480 371.670 173.740 371.900 ;
        RECT 217.860 371.890 226.980 371.900 ;
        RECT 234.800 371.890 259.810 372.070 ;
        RECT 174.400 371.690 174.720 371.700 ;
        RECT 174.390 371.680 174.720 371.690 ;
        RECT 175.430 371.680 175.750 371.730 ;
        RECT 190.470 371.680 190.750 371.690 ;
        RECT 174.390 371.670 177.060 371.680 ;
        RECT 190.450 371.670 190.770 371.680 ;
        RECT 193.180 371.670 193.500 371.700 ;
        RECT 207.500 371.670 207.820 371.730 ;
        RECT 220.790 371.670 221.330 371.680 ;
        RECT 161.500 371.440 221.330 371.670 ;
        RECT 221.870 371.590 222.410 371.890 ;
        RECT 161.500 371.410 161.830 371.440 ;
        RECT 161.500 371.390 161.810 371.410 ;
        RECT 173.480 371.400 173.740 371.440 ;
        RECT 174.390 371.430 174.720 371.440 ;
        RECT 174.400 371.410 174.720 371.430 ;
        RECT 175.480 371.400 175.820 371.440 ;
        RECT 190.450 371.420 190.770 371.440 ;
        RECT 193.180 371.420 193.500 371.440 ;
        RECT 190.470 371.410 190.750 371.420 ;
        RECT 155.420 371.210 155.740 371.220 ;
        RECT 171.210 371.210 171.670 371.360 ;
        RECT 173.380 371.210 175.820 371.400 ;
        RECT 177.000 371.210 177.160 371.240 ;
        RECT 217.330 371.210 217.640 371.270 ;
        RECT 219.850 371.210 220.380 371.240 ;
        RECT 155.420 371.040 220.380 371.210 ;
        RECT 220.790 371.120 221.330 371.440 ;
        RECT 224.590 371.480 224.900 371.680 ;
        RECT 224.590 371.470 225.190 371.480 ;
        RECT 224.590 371.350 226.980 371.470 ;
        RECT 243.260 371.400 259.810 371.890 ;
        RECT 361.100 371.810 362.500 377.320 ;
        RECT 224.730 371.310 226.980 371.350 ;
        RECT 225.040 371.290 226.980 371.310 ;
        RECT 236.960 371.150 259.810 371.400 ;
        RECT 85.760 370.390 89.850 370.990 ;
        RECT 130.540 370.980 131.050 371.000 ;
        RECT 150.180 370.980 150.580 370.990 ;
        RECT 130.540 370.630 150.580 370.980 ;
        RECT 155.420 370.980 226.980 371.040 ;
        RECT 155.420 370.920 155.740 370.980 ;
        RECT 215.450 370.830 226.980 370.980 ;
        RECT 216.760 370.820 226.980 370.830 ;
        RECT 130.540 370.590 131.050 370.630 ;
        RECT 150.180 370.600 150.580 370.630 ;
        RECT 187.320 370.630 187.640 370.670 ;
        RECT 202.970 370.630 204.250 370.730 ;
        RECT 219.850 370.630 220.380 370.820 ;
        RECT 243.260 370.750 259.810 371.150 ;
        RECT 98.460 369.880 99.080 369.900 ;
        RECT 98.460 369.510 127.610 369.880 ;
        RECT 98.460 369.440 99.080 369.510 ;
        RECT 57.640 368.750 61.020 368.860 ;
        RECT 130.260 368.780 131.530 370.240 ;
        RECT 168.460 370.110 168.560 370.430 ;
        RECT 173.480 369.650 173.740 370.450 ;
        RECT 187.320 370.420 204.250 370.630 ;
        RECT 187.320 370.390 187.640 370.420 ;
        RECT 177.380 369.980 180.230 370.180 ;
        RECT 199.740 370.050 200.020 370.070 ;
        RECT 174.400 369.940 174.720 369.950 ;
        RECT 174.390 369.930 174.720 369.940 ;
        RECT 175.430 369.930 175.750 369.980 ;
        RECT 174.390 369.730 177.060 369.930 ;
        RECT 174.390 369.680 174.720 369.730 ;
        RECT 175.430 369.720 175.750 369.730 ;
        RECT 174.400 369.660 174.720 369.680 ;
        RECT 175.480 369.650 175.820 369.710 ;
        RECT 168.560 369.130 169.120 369.300 ;
        RECT 171.210 369.290 171.670 369.610 ;
        RECT 173.380 369.430 175.820 369.650 ;
        RECT 176.990 369.290 177.160 369.490 ;
        RECT 180.030 369.480 180.230 369.980 ;
        RECT 199.720 370.020 200.040 370.050 ;
        RECT 216.430 370.020 226.980 370.070 ;
        RECT 231.860 370.020 233.200 370.560 ;
        RECT 236.960 370.230 240.470 370.420 ;
        RECT 199.720 369.810 233.200 370.020 ;
        RECT 199.720 369.790 200.040 369.810 ;
        RECT 199.740 369.770 200.020 369.790 ;
        RECT 206.050 369.480 206.360 369.540 ;
        RECT 180.030 369.280 206.360 369.480 ;
        RECT 216.540 369.470 216.800 369.710 ;
        RECT 206.050 369.220 206.360 369.280 ;
        RECT 216.430 369.360 216.800 369.470 ;
        RECT 216.430 369.210 216.750 369.360 ;
        RECT 231.860 369.280 233.200 369.810 ;
        RECT 239.600 369.630 239.920 369.760 ;
        RECT 240.240 369.630 240.470 370.230 ;
        RECT 243.500 369.980 243.790 370.750 ;
        RECT 244.690 370.680 244.950 370.750 ;
        RECT 244.690 370.470 248.820 370.680 ;
        RECT 245.030 369.980 245.350 370.070 ;
        RECT 245.720 369.980 246.580 370.470 ;
        RECT 248.610 370.330 248.820 370.470 ;
        RECT 252.230 370.340 252.560 370.550 ;
        RECT 248.610 370.120 250.620 370.330 ;
        RECT 252.670 370.110 252.980 370.440 ;
        RECT 243.500 369.760 246.580 369.980 ;
        RECT 254.340 369.950 254.650 370.140 ;
        RECT 243.500 369.750 243.790 369.760 ;
        RECT 241.830 369.630 242.150 369.750 ;
        RECT 245.720 369.710 246.580 369.760 ;
        RECT 248.180 369.750 248.490 369.910 ;
        RECT 238.820 369.480 240.700 369.630 ;
        RECT 241.690 369.490 242.150 369.630 ;
        RECT 244.980 369.530 246.580 369.710 ;
        RECT 247.750 369.530 248.630 369.750 ;
        RECT 251.990 369.720 254.700 369.950 ;
        RECT 241.690 369.480 242.060 369.490 ;
        RECT 244.610 369.480 250.610 369.530 ;
        RECT 238.820 369.430 250.610 369.480 ;
        RECT 252.720 369.460 253.030 369.720 ;
        RECT 240.240 369.330 250.610 369.430 ;
        RECT 240.240 369.320 250.480 369.330 ;
        RECT 240.240 369.260 245.000 369.320 ;
        RECT 245.030 369.210 245.350 369.320 ;
        RECT 141.610 368.780 141.910 368.790 ;
        RECT 147.300 368.780 147.610 368.910 ;
        RECT 148.390 368.780 148.700 368.920 ;
        RECT 151.200 368.780 151.490 368.800 ;
        RECT 57.230 366.500 127.730 368.750 ;
        RECT 130.260 368.390 151.520 368.780 ;
        RECT 168.560 368.680 168.730 369.130 ;
        RECT 184.980 369.010 185.300 369.060 ;
        RECT 245.720 369.050 246.580 369.320 ;
        RECT 246.680 369.050 246.990 369.320 ;
        RECT 248.340 369.080 248.650 369.300 ;
        RECT 248.330 369.050 248.650 369.080 ;
        RECT 179.980 368.810 185.350 369.010 ;
        RECT 245.720 368.970 248.650 369.050 ;
        RECT 167.590 368.570 167.980 368.660 ;
        RECT 168.460 368.570 168.730 368.680 ;
        RECT 167.590 368.400 168.740 368.570 ;
        RECT 130.260 368.360 131.530 368.390 ;
        RECT 151.200 368.370 151.490 368.390 ;
        RECT 168.460 368.360 168.560 368.400 ;
        RECT 145.460 368.220 145.530 368.260 ;
        RECT 145.460 367.990 145.600 368.220 ;
        RECT 147.440 368.000 148.260 368.170 ;
        RECT 145.760 367.970 146.070 368.000 ;
        RECT 150.560 367.970 150.850 367.990 ;
        RECT 138.110 367.570 150.870 367.970 ;
        RECT 173.480 367.900 173.740 368.700 ;
        RECT 179.980 368.430 180.180 368.810 ;
        RECT 184.980 368.800 185.300 368.810 ;
        RECT 225.440 368.760 225.520 368.940 ;
        RECT 239.290 368.650 239.600 368.930 ;
        RECT 238.820 368.610 239.600 368.650 ;
        RECT 240.430 368.650 240.650 368.660 ;
        RECT 240.960 368.650 241.270 368.930 ;
        RECT 245.720 368.890 248.640 368.970 ;
        RECT 245.720 368.820 248.840 368.890 ;
        RECT 245.720 368.680 246.580 368.820 ;
        RECT 246.630 368.680 246.940 368.690 ;
        RECT 248.290 368.680 248.840 368.820 ;
        RECT 250.050 368.680 250.370 368.760 ;
        RECT 284.550 368.680 287.860 370.740 ;
        RECT 240.430 368.610 242.060 368.650 ;
        RECT 243.260 368.610 288.180 368.680 ;
        RECT 187.740 368.570 188.050 368.580 ;
        RECT 217.370 368.570 217.800 368.590 ;
        RECT 233.860 368.570 288.180 368.610 ;
        RECT 187.740 368.540 188.060 368.570 ;
        RECT 177.380 368.230 180.180 368.430 ;
        RECT 180.490 368.340 188.060 368.540 ;
        RECT 217.370 368.510 288.180 368.570 ;
        RECT 174.400 368.190 174.720 368.200 ;
        RECT 174.390 368.180 174.720 368.190 ;
        RECT 175.430 368.180 175.750 368.230 ;
        RECT 174.390 367.980 177.060 368.180 ;
        RECT 174.390 367.930 174.720 367.980 ;
        RECT 175.430 367.970 175.750 367.980 ;
        RECT 174.400 367.910 174.720 367.930 ;
        RECT 175.480 367.900 175.820 367.960 ;
        RECT 57.640 366.180 61.020 366.500 ;
        RECT 101.810 365.460 102.290 365.490 ;
        RECT 101.810 365.080 127.600 365.460 ;
        RECT 101.810 365.060 102.290 365.080 ;
        RECT 130.550 364.880 131.820 365.750 ;
        RECT 138.110 364.880 138.510 367.570 ;
        RECT 146.640 367.510 147.240 367.570 ;
        RECT 148.500 367.520 148.720 367.570 ;
        RECT 150.560 367.560 150.850 367.570 ;
        RECT 171.210 367.540 171.670 367.860 ;
        RECT 173.380 367.680 175.820 367.900 ;
        RECT 176.970 367.540 177.160 367.740 ;
        RECT 168.560 367.300 169.120 367.470 ;
        RECT 145.460 367.070 145.600 367.240 ;
        RECT 147.440 367.080 148.260 367.250 ;
        RECT 141.910 366.890 142.280 366.900 ;
        RECT 140.120 366.660 142.280 366.890 ;
        RECT 145.460 366.660 145.630 366.830 ;
        RECT 145.740 366.750 146.050 367.080 ;
        RECT 166.990 367.030 167.320 367.040 ;
        RECT 146.640 366.660 147.240 366.690 ;
        RECT 147.310 366.660 147.620 366.930 ;
        RECT 140.120 366.600 147.620 366.660 ;
        RECT 148.400 366.700 148.710 366.940 ;
        RECT 166.970 366.930 167.340 367.030 ;
        RECT 168.560 366.930 168.730 367.300 ;
        RECT 166.970 366.760 168.730 366.930 ;
        RECT 148.400 366.610 148.720 366.700 ;
        RECT 150.570 366.670 150.890 366.720 ;
        RECT 140.120 366.530 147.540 366.600 ;
        RECT 148.500 366.530 148.720 366.610 ;
        RECT 140.120 365.830 140.740 366.530 ;
        RECT 141.910 366.490 147.540 366.530 ;
        RECT 150.000 366.500 150.950 366.670 ;
        RECT 166.970 366.650 167.340 366.760 ;
        RECT 168.460 366.750 168.730 366.760 ;
        RECT 168.460 366.610 168.560 366.750 ;
        RECT 150.570 366.460 150.890 366.500 ;
        RECT 145.460 366.290 145.600 366.320 ;
        RECT 145.460 366.150 145.670 366.290 ;
        RECT 146.800 366.250 147.120 366.300 ;
        RECT 147.440 366.250 148.260 366.330 ;
        RECT 146.800 366.160 148.260 366.250 ;
        RECT 141.910 365.830 142.280 365.870 ;
        RECT 130.550 364.480 138.510 364.880 ;
        RECT 139.590 365.740 142.280 365.830 ;
        RECT 145.460 365.740 145.620 365.910 ;
        RECT 145.720 365.760 146.030 366.090 ;
        RECT 146.800 366.080 147.540 366.160 ;
        RECT 173.480 366.150 173.740 366.950 ;
        RECT 180.490 366.680 180.690 368.340 ;
        RECT 187.740 368.310 188.060 368.340 ;
        RECT 187.740 368.300 188.050 368.310 ;
        RECT 217.330 368.290 288.180 368.510 ;
        RECT 215.450 368.200 288.180 368.290 ;
        RECT 215.450 368.110 226.980 368.200 ;
        RECT 241.850 368.110 242.170 368.200 ;
        RECT 188.800 368.060 189.120 368.100 ;
        RECT 215.450 368.080 242.170 368.110 ;
        RECT 216.760 368.070 242.170 368.080 ;
        RECT 177.380 366.480 180.690 366.680 ;
        RECT 181.040 367.860 189.200 368.060 ;
        RECT 219.650 367.930 242.170 368.070 ;
        RECT 242.970 368.010 288.180 368.200 ;
        RECT 174.400 366.440 174.720 366.450 ;
        RECT 174.390 366.430 174.720 366.440 ;
        RECT 175.430 366.430 175.750 366.480 ;
        RECT 174.390 366.230 177.060 366.430 ;
        RECT 174.390 366.180 174.720 366.230 ;
        RECT 175.430 366.220 175.750 366.230 ;
        RECT 174.400 366.160 174.720 366.180 ;
        RECT 175.480 366.150 175.820 366.210 ;
        RECT 146.800 366.040 147.120 366.080 ;
        RECT 146.740 365.750 147.110 365.940 ;
        RECT 147.220 365.870 147.530 366.080 ;
        RECT 148.520 365.770 148.830 366.100 ;
        RECT 150.570 365.750 150.890 365.800 ;
        RECT 171.210 365.790 171.670 366.110 ;
        RECT 173.380 365.930 175.820 366.150 ;
        RECT 177.000 365.790 177.160 365.990 ;
        RECT 139.590 365.570 147.540 365.740 ;
        RECT 150.000 365.580 150.950 365.750 ;
        RECT 139.590 365.460 142.280 365.570 ;
        RECT 150.570 365.540 150.890 365.580 ;
        RECT 168.520 365.570 169.120 365.740 ;
        RECT 139.590 365.350 140.740 365.460 ;
        RECT 139.590 364.900 140.700 365.350 ;
        RECT 146.740 365.330 147.120 365.520 ;
        RECT 147.310 365.330 147.630 365.490 ;
        RECT 145.460 365.130 145.600 365.320 ;
        RECT 146.770 365.260 147.630 365.330 ;
        RECT 166.390 365.450 166.780 365.550 ;
        RECT 168.520 365.450 168.690 365.570 ;
        RECT 166.390 365.280 168.690 365.450 ;
        RECT 146.770 365.160 148.260 365.260 ;
        RECT 166.390 365.180 166.780 365.280 ;
        RECT 146.770 365.120 147.090 365.160 ;
        RECT 147.220 365.060 148.260 365.160 ;
        RECT 141.910 364.900 142.280 364.940 ;
        RECT 139.590 364.820 142.280 364.900 ;
        RECT 145.460 364.820 145.600 364.900 ;
        RECT 146.740 364.820 147.110 364.950 ;
        RECT 147.220 364.880 147.530 365.060 ;
        RECT 139.590 364.650 147.540 364.820 ;
        RECT 148.520 364.780 148.830 365.110 ;
        RECT 150.540 364.830 150.860 364.880 ;
        RECT 168.460 364.860 168.560 365.180 ;
        RECT 181.040 364.930 181.240 367.860 ;
        RECT 188.800 367.820 189.120 367.860 ;
        RECT 207.440 367.260 208.020 367.700 ;
        RECT 207.440 367.070 208.080 367.260 ;
        RECT 207.840 366.460 208.080 367.070 ;
        RECT 208.460 367.060 209.040 367.690 ;
        RECT 211.280 367.550 211.750 367.610 ;
        RECT 219.410 367.600 219.480 367.780 ;
        RECT 224.620 367.660 224.930 367.930 ;
        RECT 238.890 367.820 239.210 367.930 ;
        RECT 243.260 367.820 288.180 368.010 ;
        RECT 225.030 367.550 226.980 367.760 ;
        RECT 238.510 367.750 239.210 367.820 ;
        RECT 235.880 367.550 235.930 367.670 ;
        RECT 238.510 367.620 239.120 367.750 ;
        RECT 243.200 367.620 288.180 367.820 ;
        RECT 236.180 367.560 236.470 367.570 ;
        RECT 236.180 367.550 236.480 367.560 ;
        RECT 243.260 367.550 288.180 367.620 ;
        RECT 211.280 367.120 288.180 367.550 ;
        RECT 217.880 367.040 226.980 367.120 ;
        RECT 228.310 367.000 229.150 367.120 ;
        RECT 234.800 367.040 288.180 367.120 ;
        RECT 212.860 366.780 213.170 366.920 ;
        RECT 239.380 366.840 240.500 366.850 ;
        RECT 210.690 366.600 213.170 366.780 ;
        RECT 238.510 366.750 240.500 366.840 ;
        RECT 212.860 366.590 213.170 366.600 ;
        RECT 228.760 366.640 240.500 366.750 ;
        RECT 228.760 366.530 238.900 366.640 ;
        RECT 239.380 366.630 240.500 366.640 ;
        RECT 235.880 366.490 235.940 366.530 ;
        RECT 238.680 366.430 238.900 366.530 ;
        RECT 239.600 366.430 239.920 366.560 ;
        RECT 240.570 366.490 240.640 366.690 ;
        RECT 241.830 366.430 242.150 366.550 ;
        RECT 242.290 366.540 242.640 366.760 ;
        RECT 243.260 366.620 288.180 367.040 ;
        RECT 232.360 366.260 232.660 366.280 ;
        RECT 238.680 366.260 240.700 366.430 ;
        RECT 241.690 366.290 242.150 366.430 ;
        RECT 244.100 366.470 244.300 366.480 ;
        RECT 241.690 366.260 242.060 366.290 ;
        RECT 244.100 366.260 244.320 366.470 ;
        RECT 246.210 366.440 246.570 366.450 ;
        RECT 245.650 366.260 246.570 366.440 ;
        RECT 246.680 366.430 246.990 366.620 ;
        RECT 248.610 366.600 251.090 366.620 ;
        RECT 248.610 366.590 248.920 366.600 ;
        RECT 150.000 364.660 150.950 364.830 ;
        RECT 177.340 364.730 181.240 364.930 ;
        RECT 184.190 366.060 184.480 366.240 ;
        RECT 232.350 366.160 246.570 366.260 ;
        RECT 232.350 366.080 246.610 366.160 ;
        RECT 246.680 366.080 246.990 366.340 ;
        RECT 248.380 366.080 248.690 366.360 ;
        RECT 139.590 364.530 142.280 364.650 ;
        RECT 150.540 364.620 150.860 364.660 ;
        RECT 139.590 364.490 140.490 364.530 ;
        RECT 130.550 363.870 131.820 364.480 ;
        RECT 98.340 361.590 98.960 361.680 ;
        RECT 98.340 361.180 127.280 361.590 ;
        RECT 98.340 361.090 98.960 361.180 ;
        RECT 101.810 360.690 102.350 360.720 ;
        RECT 101.810 360.280 127.240 360.690 ;
        RECT 101.810 360.240 102.350 360.280 ;
        RECT 130.980 359.940 132.250 360.820 ;
        RECT 139.590 359.940 139.960 364.490 ;
        RECT 146.740 364.410 147.120 364.530 ;
        RECT 147.310 364.410 147.630 364.500 ;
        RECT 145.460 364.340 145.600 364.360 ;
        RECT 146.740 364.340 147.630 364.410 ;
        RECT 145.460 364.170 145.530 364.340 ;
        RECT 146.780 364.300 147.630 364.340 ;
        RECT 146.780 364.240 148.260 364.300 ;
        RECT 146.780 364.200 147.100 364.240 ;
        RECT 147.310 364.220 148.260 364.240 ;
        RECT 147.220 364.100 148.260 364.220 ;
        RECT 145.460 363.920 145.600 363.940 ;
        RECT 145.460 363.820 145.530 363.920 ;
        RECT 146.740 363.820 147.110 363.960 ;
        RECT 147.220 363.890 147.530 364.100 ;
        RECT 141.070 363.800 147.560 363.820 ;
        RECT 130.980 359.570 139.960 359.940 ;
        RECT 140.780 363.630 147.560 363.800 ;
        RECT 148.520 363.790 148.830 364.120 ;
        RECT 165.750 363.850 166.140 363.940 ;
        RECT 168.690 363.850 169.120 364.020 ;
        RECT 151.180 363.760 151.500 363.790 ;
        RECT 140.780 363.450 142.280 363.630 ;
        RECT 149.970 363.560 151.600 363.760 ;
        RECT 165.750 363.680 169.320 363.850 ;
        RECT 165.750 363.590 166.140 363.680 ;
        RECT 168.690 363.660 168.860 363.680 ;
        RECT 140.780 362.860 141.440 363.450 ;
        RECT 141.910 363.410 142.280 363.450 ;
        RECT 146.130 363.400 146.450 363.440 ;
        RECT 146.740 363.400 147.120 363.540 ;
        RECT 151.180 363.530 151.500 363.560 ;
        RECT 147.310 363.400 147.630 363.510 ;
        RECT 145.460 363.350 145.600 363.400 ;
        RECT 145.460 363.210 145.530 363.350 ;
        RECT 146.130 363.340 147.630 363.400 ;
        RECT 146.130 363.210 148.260 363.340 ;
        RECT 146.130 363.180 146.450 363.210 ;
        RECT 147.310 363.190 148.260 363.210 ;
        RECT 147.450 363.140 148.260 363.190 ;
        RECT 165.110 363.280 165.500 363.390 ;
        RECT 165.110 363.110 169.320 363.280 ;
        RECT 184.190 363.220 184.370 366.060 ;
        RECT 232.350 365.860 248.870 366.080 ;
        RECT 232.350 365.840 246.610 365.860 ;
        RECT 232.360 365.820 232.660 365.840 ;
        RECT 235.880 365.780 235.940 365.840 ;
        RECT 238.680 365.810 238.900 365.840 ;
        RECT 239.380 365.810 240.500 365.820 ;
        RECT 228.710 365.560 237.720 365.780 ;
        RECT 238.510 365.610 240.500 365.810 ;
        RECT 240.570 365.760 240.640 365.840 ;
        RECT 227.890 365.120 228.210 365.170 ;
        RECT 227.890 364.870 233.910 365.120 ;
        RECT 233.590 364.800 233.910 364.870 ;
        RECT 235.880 364.780 235.930 364.980 ;
        RECT 235.880 364.270 235.930 364.470 ;
        RECT 208.540 363.630 209.140 364.190 ;
        RECT 212.140 364.020 217.370 364.250 ;
        RECT 217.740 364.020 226.890 364.250 ;
        RECT 226.600 363.920 226.890 364.020 ;
        RECT 228.760 363.920 234.420 364.000 ;
        RECT 234.580 363.920 235.720 364.000 ;
        RECT 226.600 363.800 235.720 363.920 ;
        RECT 237.500 363.950 237.720 365.560 ;
        RECT 238.680 365.450 238.900 365.610 ;
        RECT 239.290 365.600 240.500 365.610 ;
        RECT 239.290 365.450 239.600 365.600 ;
        RECT 238.680 365.400 239.600 365.450 ;
        RECT 240.430 365.450 240.650 365.460 ;
        RECT 240.960 365.450 241.270 365.730 ;
        RECT 238.680 365.330 239.390 365.400 ;
        RECT 238.650 365.250 239.390 365.330 ;
        RECT 240.430 365.250 242.060 365.450 ;
        RECT 243.050 365.340 243.370 365.580 ;
        RECT 245.650 365.500 246.610 365.840 ;
        RECT 238.650 364.830 238.910 365.250 ;
        RECT 240.430 365.240 240.650 365.250 ;
        RECT 238.510 364.810 239.120 364.830 ;
        RECT 238.510 364.650 239.210 364.810 ;
        RECT 238.510 364.630 242.780 364.650 ;
        RECT 243.200 364.630 243.270 364.830 ;
        RECT 238.650 364.620 242.780 364.630 ;
        RECT 238.510 364.440 242.780 364.620 ;
        RECT 238.510 364.420 239.120 364.440 ;
        RECT 242.570 364.300 242.780 364.440 ;
        RECT 243.200 364.600 243.270 364.620 ;
        RECT 245.710 364.600 246.610 365.500 ;
        RECT 246.630 365.360 246.940 365.690 ;
        RECT 247.390 365.570 247.500 365.800 ;
        RECT 247.390 364.750 247.500 364.970 ;
        RECT 312.940 364.600 316.870 365.050 ;
        RECT 243.200 364.420 316.870 364.600 ;
        RECT 243.260 364.300 316.870 364.420 ;
        RECT 242.570 364.090 316.870 364.300 ;
        RECT 240.430 364.000 240.650 364.010 ;
        RECT 238.820 363.950 239.390 364.000 ;
        RECT 226.600 363.720 234.930 363.800 ;
        RECT 237.500 363.730 240.350 363.950 ;
        RECT 240.430 363.800 242.060 364.000 ;
        RECT 240.430 363.790 240.650 363.800 ;
        RECT 226.600 363.710 226.890 363.720 ;
        RECT 228.260 363.480 228.740 363.490 ;
        RECT 165.110 363.010 165.500 363.110 ;
        RECT 183.420 363.050 184.370 363.220 ;
        RECT 192.310 363.040 194.090 363.210 ;
        RECT 212.150 363.200 217.370 363.420 ;
        RECT 217.740 363.200 225.950 363.420 ;
        RECT 228.260 363.240 229.150 363.480 ;
        RECT 234.200 363.450 234.420 363.720 ;
        RECT 239.290 363.650 239.600 363.730 ;
        RECT 239.290 363.640 240.500 363.650 ;
        RECT 238.510 363.500 240.500 363.640 ;
        RECT 240.960 363.520 241.270 363.800 ;
        RECT 242.140 363.720 242.450 363.880 ;
        RECT 241.710 363.500 242.590 363.720 ;
        RECT 243.260 363.500 316.870 364.090 ;
        RECT 235.880 363.450 235.940 363.490 ;
        RECT 238.510 363.450 316.870 363.500 ;
        RECT 234.200 363.290 316.870 363.450 ;
        RECT 234.200 363.230 238.960 363.290 ;
        RECT 145.460 362.960 145.600 362.980 ;
        RECT 145.460 362.860 145.610 362.960 ;
        RECT 140.780 362.670 147.560 362.860 ;
        RECT 151.190 362.800 151.510 362.830 ;
        RECT 140.780 362.490 142.280 362.670 ;
        RECT 149.970 362.600 151.600 362.800 ;
        RECT 187.290 362.760 187.610 362.810 ;
        RECT 189.700 362.760 190.020 362.780 ;
        RECT 177.760 362.620 177.960 362.740 ;
        RECT 151.190 362.570 151.510 362.600 ;
        RECT 140.780 362.480 141.450 362.490 ;
        RECT 140.780 362.440 141.440 362.480 ;
        RECT 141.910 362.450 142.280 362.490 ;
        RECT 146.090 362.440 146.410 362.480 ;
        RECT 130.980 358.940 132.250 359.570 ;
        RECT 130.920 355.180 132.190 356.070 ;
        RECT 140.780 355.180 141.150 362.440 ;
        RECT 146.090 362.250 147.560 362.440 ;
        RECT 177.760 362.420 178.110 362.620 ;
        RECT 187.290 362.570 190.020 362.760 ;
        RECT 219.410 362.730 219.490 362.910 ;
        RECT 187.290 362.490 187.610 362.570 ;
        RECT 188.370 362.500 188.460 362.570 ;
        RECT 189.700 362.520 190.020 362.570 ;
        RECT 177.760 362.400 177.960 362.420 ;
        RECT 146.090 362.220 146.410 362.250 ;
        RECT 168.460 361.950 168.560 362.270 ;
        RECT 177.380 362.200 177.960 362.400 ;
        RECT 186.090 362.050 186.530 362.280 ;
        RECT 186.190 361.980 186.530 362.050 ;
        RECT 130.920 354.810 141.150 355.180 ;
        RECT 141.910 361.710 147.560 361.900 ;
        RECT 151.180 361.840 151.500 361.870 ;
        RECT 186.190 361.840 186.530 361.910 ;
        RECT 130.920 354.190 132.190 354.810 ;
        RECT 130.980 350.340 132.250 351.250 ;
        RECT 141.910 350.340 142.280 361.710 ;
        RECT 149.970 361.640 151.600 361.840 ;
        RECT 164.500 361.710 164.890 361.810 ;
        RECT 151.180 361.610 151.500 361.640 ;
        RECT 164.500 361.540 169.320 361.710 ;
        RECT 186.090 361.610 186.530 361.840 ;
        RECT 146.130 361.480 146.450 361.520 ;
        RECT 146.130 361.290 147.560 361.480 ;
        RECT 164.500 361.440 164.890 361.540 ;
        RECT 168.770 361.380 169.120 361.540 ;
        RECT 146.130 361.260 146.450 361.290 ;
        RECT 171.210 361.020 171.670 361.340 ;
        RECT 173.380 360.980 175.820 361.200 ;
        RECT 177.000 361.140 177.160 361.340 ;
        RECT 177.710 361.200 178.080 361.400 ;
        RECT 163.870 360.180 164.290 360.270 ;
        RECT 168.460 360.200 168.560 360.520 ;
        RECT 173.480 360.180 173.740 360.980 ;
        RECT 174.400 360.950 174.720 360.970 ;
        RECT 174.390 360.900 174.720 360.950 ;
        RECT 175.480 360.920 175.820 360.980 ;
        RECT 175.430 360.900 175.750 360.910 ;
        RECT 174.390 360.700 177.060 360.900 ;
        RECT 174.390 360.690 174.720 360.700 ;
        RECT 174.400 360.680 174.720 360.690 ;
        RECT 175.430 360.650 175.750 360.700 ;
        RECT 177.710 360.650 177.910 361.200 ;
        RECT 183.750 361.170 184.480 361.350 ;
        RECT 187.290 361.320 187.610 361.400 ;
        RECT 188.370 361.320 188.450 361.390 ;
        RECT 189.700 361.320 190.020 361.370 ;
        RECT 183.750 360.960 183.930 361.170 ;
        RECT 187.290 361.130 190.020 361.320 ;
        RECT 187.290 361.080 187.610 361.130 ;
        RECT 189.700 361.110 190.020 361.130 ;
        RECT 225.730 361.320 225.950 363.200 ;
        RECT 228.350 362.940 228.810 363.070 ;
        RECT 234.660 362.940 235.720 363.020 ;
        RECT 228.350 362.820 235.720 362.940 ;
        RECT 238.820 362.960 242.060 363.020 ;
        RECT 238.820 362.820 242.150 362.960 ;
        RECT 242.290 362.860 242.600 363.050 ;
        RECT 228.350 362.740 234.930 362.820 ;
        RECT 228.350 362.620 228.810 362.740 ;
        RECT 233.590 362.580 233.910 362.590 ;
        RECT 235.880 362.580 235.940 362.760 ;
        RECT 239.600 362.690 239.920 362.820 ;
        RECT 240.080 362.740 241.790 362.820 ;
        RECT 239.380 362.610 240.500 362.620 ;
        RECT 238.510 362.580 240.500 362.610 ;
        RECT 240.570 362.580 240.640 362.740 ;
        RECT 241.590 362.580 241.790 362.740 ;
        RECT 241.830 362.700 242.150 362.820 ;
        RECT 242.250 362.610 242.800 362.860 ;
        RECT 243.260 362.580 316.870 363.290 ;
        RECT 233.590 362.540 316.870 362.580 ;
        RECT 233.590 362.420 244.360 362.540 ;
        RECT 312.940 362.530 316.870 362.540 ;
        RECT 233.590 362.410 234.280 362.420 ;
        RECT 238.510 362.410 240.500 362.420 ;
        RECT 229.360 362.290 229.720 362.390 ;
        RECT 233.590 362.290 233.910 362.410 ;
        RECT 239.380 362.400 240.500 362.410 ;
        RECT 241.590 362.290 241.790 362.420 ;
        RECT 229.360 362.090 235.720 362.290 ;
        RECT 240.080 362.090 241.790 362.290 ;
        RECT 229.360 361.970 229.720 362.090 ;
        RECT 241.450 361.880 241.790 362.090 ;
        RECT 235.880 361.580 235.930 361.780 ;
        RECT 238.510 361.500 239.120 361.630 ;
        RECT 238.510 361.430 239.210 361.500 ;
        RECT 225.730 361.310 227.330 361.320 ;
        RECT 225.730 361.110 235.720 361.310 ;
        RECT 238.890 361.240 239.210 361.430 ;
        RECT 225.730 361.100 227.330 361.110 ;
        RECT 241.590 361.040 241.790 361.880 ;
        RECT 242.430 361.580 242.900 361.830 ;
        RECT 242.570 361.490 242.890 361.580 ;
        RECT 243.200 361.430 243.270 361.630 ;
        RECT 245.680 361.040 246.580 361.710 ;
        RECT 190.450 361.010 190.760 361.020 ;
        RECT 183.360 360.780 183.930 360.960 ;
        RECT 190.440 360.950 190.770 361.010 ;
        RECT 190.090 360.900 190.770 360.950 ;
        RECT 186.860 360.730 190.770 360.900 ;
        RECT 192.090 360.790 194.090 360.950 ;
        RECT 192.820 360.780 194.090 360.790 ;
        RECT 193.520 360.770 194.090 360.780 ;
        RECT 212.920 360.740 217.370 360.900 ;
        RECT 186.860 360.680 190.760 360.730 ;
        RECT 212.890 360.700 217.370 360.740 ;
        RECT 217.740 360.800 234.930 360.900 ;
        RECT 240.430 360.800 240.650 360.810 ;
        RECT 241.590 360.800 246.580 361.040 ;
        RECT 217.740 360.700 235.720 360.800 ;
        RECT 177.380 360.450 177.910 360.650 ;
        RECT 163.870 360.010 168.770 360.180 ;
        RECT 163.870 359.920 164.290 360.010 ;
        RECT 168.600 359.830 168.770 360.010 ;
        RECT 183.850 360.020 184.400 360.200 ;
        RECT 207.480 360.160 208.040 360.700 ;
        RECT 183.850 360.000 184.030 360.020 ;
        RECT 183.430 359.840 184.030 360.000 ;
        RECT 192.310 359.830 194.090 359.990 ;
        RECT 168.600 359.660 169.120 359.830 ;
        RECT 171.210 359.270 171.670 359.590 ;
        RECT 173.380 359.230 175.820 359.450 ;
        RECT 176.970 359.390 177.160 359.590 ;
        RECT 187.290 359.560 187.610 359.610 ;
        RECT 189.700 359.560 190.020 359.580 ;
        RECT 163.310 358.610 163.700 358.700 ;
        RECT 168.460 358.610 168.560 358.770 ;
        RECT 163.310 358.440 168.680 358.610 ;
        RECT 163.310 358.350 163.700 358.440 ;
        RECT 168.520 358.330 168.680 358.440 ;
        RECT 173.480 358.430 173.740 359.230 ;
        RECT 174.400 359.200 174.720 359.220 ;
        RECT 174.390 359.150 174.720 359.200 ;
        RECT 175.480 359.170 175.820 359.230 ;
        RECT 175.430 359.150 175.750 359.160 ;
        RECT 174.390 358.950 177.060 359.150 ;
        RECT 177.740 359.090 178.060 359.530 ;
        RECT 187.290 359.370 190.020 359.560 ;
        RECT 187.290 359.290 187.610 359.370 ;
        RECT 188.370 359.290 188.520 359.370 ;
        RECT 189.700 359.320 190.020 359.370 ;
        RECT 174.390 358.940 174.720 358.950 ;
        RECT 174.400 358.930 174.720 358.940 ;
        RECT 175.430 358.900 175.750 358.950 ;
        RECT 177.740 358.900 177.940 359.090 ;
        RECT 177.380 358.700 177.940 358.900 ;
        RECT 186.090 358.850 186.530 359.080 ;
        RECT 186.190 358.780 186.530 358.850 ;
        RECT 186.190 358.640 186.530 358.710 ;
        RECT 186.090 358.410 186.530 358.640 ;
        RECT 168.520 358.030 168.690 358.330 ;
        RECT 212.890 358.220 213.120 360.700 ;
        RECT 234.630 360.600 235.720 360.700 ;
        RECT 238.820 360.650 239.390 360.800 ;
        RECT 238.820 360.600 239.600 360.650 ;
        RECT 239.290 360.320 239.600 360.600 ;
        RECT 240.430 360.610 246.580 360.800 ;
        RECT 240.430 360.600 242.060 360.610 ;
        RECT 242.180 360.600 242.490 360.610 ;
        RECT 240.430 360.590 240.650 360.600 ;
        RECT 240.960 360.320 241.270 360.600 ;
        RECT 230.280 360.030 230.670 360.050 ;
        RECT 230.270 359.920 230.680 360.030 ;
        RECT 241.590 359.920 241.790 360.600 ;
        RECT 245.680 360.260 246.580 360.610 ;
        RECT 341.740 360.260 345.240 360.800 ;
        RECT 230.270 359.820 234.930 359.920 ;
        RECT 240.080 359.820 241.790 359.920 ;
        RECT 230.270 359.720 235.720 359.820 ;
        RECT 230.270 359.620 230.680 359.720 ;
        RECT 234.700 359.620 235.720 359.720 ;
        RECT 238.820 359.760 242.060 359.820 ;
        RECT 238.820 359.620 242.150 359.760 ;
        RECT 230.280 359.600 230.670 359.620 ;
        RECT 239.600 359.490 239.920 359.620 ;
        RECT 231.100 359.330 231.500 359.340 ;
        RECT 231.080 359.270 231.520 359.330 ;
        RECT 241.590 359.270 241.790 359.620 ;
        RECT 241.830 359.500 242.150 359.620 ;
        RECT 231.080 359.090 234.930 359.270 ;
        RECT 240.080 359.090 241.790 359.270 ;
        RECT 231.080 359.070 235.720 359.090 ;
        RECT 231.100 359.060 231.500 359.070 ;
        RECT 234.580 358.890 235.720 359.070 ;
        RECT 240.020 358.950 241.790 359.090 ;
        RECT 240.020 358.890 241.780 358.950 ;
        RECT 168.520 357.860 169.120 358.030 ;
        RECT 177.670 357.970 178.050 358.150 ;
        RECT 187.290 358.120 187.610 358.200 ;
        RECT 188.370 358.120 188.450 358.190 ;
        RECT 189.700 358.120 190.020 358.170 ;
        RECT 171.210 357.520 171.670 357.840 ;
        RECT 173.380 357.480 175.820 357.700 ;
        RECT 176.990 357.640 177.160 357.840 ;
        RECT 168.460 356.700 168.560 357.020 ;
        RECT 173.480 356.680 173.740 357.480 ;
        RECT 174.400 357.450 174.720 357.470 ;
        RECT 174.390 357.400 174.720 357.450 ;
        RECT 175.480 357.420 175.820 357.480 ;
        RECT 175.430 357.400 175.750 357.410 ;
        RECT 174.390 357.200 177.060 357.400 ;
        RECT 174.390 357.190 174.720 357.200 ;
        RECT 174.400 357.180 174.720 357.190 ;
        RECT 175.430 357.150 175.750 357.200 ;
        RECT 177.670 357.150 177.850 357.970 ;
        RECT 187.290 357.930 190.020 358.120 ;
        RECT 187.290 357.880 187.610 357.930 ;
        RECT 189.700 357.910 190.020 357.930 ;
        RECT 183.410 357.520 184.130 357.700 ;
        RECT 177.380 356.950 177.860 357.150 ;
        RECT 171.210 355.770 171.670 356.090 ;
        RECT 173.380 355.730 175.820 355.950 ;
        RECT 177.000 355.890 177.160 356.090 ;
        RECT 173.480 354.930 173.740 355.730 ;
        RECT 174.400 355.700 174.720 355.720 ;
        RECT 174.390 355.650 174.720 355.700 ;
        RECT 175.480 355.670 175.820 355.730 ;
        RECT 175.430 355.650 175.750 355.660 ;
        RECT 174.390 355.450 177.060 355.650 ;
        RECT 174.390 355.440 174.720 355.450 ;
        RECT 174.400 355.430 174.720 355.440 ;
        RECT 175.430 355.400 175.750 355.450 ;
        RECT 183.950 355.330 184.130 357.520 ;
        RECT 192.310 357.510 194.090 357.690 ;
        RECT 205.030 357.520 205.340 357.810 ;
        RECT 208.520 357.610 209.140 358.140 ;
        RECT 212.140 357.990 213.120 358.220 ;
        RECT 213.730 358.090 217.370 358.290 ;
        RECT 217.740 358.110 234.930 358.290 ;
        RECT 243.260 358.210 345.330 360.260 ;
        RECT 217.740 358.090 235.720 358.110 ;
        RECT 203.010 357.480 205.340 357.520 ;
        RECT 203.010 357.340 205.190 357.480 ;
        RECT 213.730 357.390 213.930 358.090 ;
        RECT 234.670 357.910 235.720 358.090 ;
        RECT 231.840 357.520 232.150 357.810 ;
        RECT 231.840 357.480 234.170 357.520 ;
        RECT 205.030 357.090 205.340 357.260 ;
        RECT 212.150 357.240 213.930 357.390 ;
        RECT 231.990 357.340 234.170 357.480 ;
        RECT 212.150 357.170 213.900 357.240 ;
        RECT 203.010 356.930 205.340 357.090 ;
        RECT 203.010 356.910 205.180 356.930 ;
        RECT 205.480 356.910 205.570 357.090 ;
        RECT 208.340 356.930 215.970 357.110 ;
        RECT 221.210 356.930 228.840 357.110 ;
        RECT 231.840 357.090 232.150 357.260 ;
        RECT 231.610 356.910 231.700 357.090 ;
        RECT 231.840 356.930 234.170 357.090 ;
        RECT 232.000 356.910 234.170 356.930 ;
        RECT 208.340 356.490 215.970 356.670 ;
        RECT 221.210 356.490 228.840 356.670 ;
        RECT 245.680 356.150 246.580 356.330 ;
        RECT 353.440 356.190 359.150 361.830 ;
        RECT 353.000 356.150 359.150 356.190 ;
        RECT 243.260 355.690 359.150 356.150 ;
        RECT 208.340 355.390 215.970 355.570 ;
        RECT 221.210 355.390 228.840 355.570 ;
        RECT 243.260 355.560 358.990 355.690 ;
        RECT 183.950 355.150 184.490 355.330 ;
        RECT 203.010 355.140 205.180 355.160 ;
        RECT 203.010 354.980 205.340 355.140 ;
        RECT 205.480 354.980 205.570 355.160 ;
        RECT 205.030 354.810 205.340 354.980 ;
        RECT 208.340 354.960 215.970 355.140 ;
        RECT 221.210 354.960 228.840 355.140 ;
        RECT 231.610 354.980 231.700 355.160 ;
        RECT 232.000 355.140 234.170 355.160 ;
        RECT 231.840 354.980 234.170 355.140 ;
        RECT 231.840 354.810 232.150 354.980 ;
        RECT 242.940 354.790 358.990 355.560 ;
        RECT 203.010 354.590 205.190 354.730 ;
        RECT 231.990 354.590 234.170 354.730 ;
        RECT 203.010 354.550 205.340 354.590 ;
        RECT 187.090 354.390 187.410 354.400 ;
        RECT 205.030 354.390 205.340 354.550 ;
        RECT 231.840 354.550 234.170 354.590 ;
        RECT 214.900 354.390 215.360 354.460 ;
        RECT 187.090 354.110 215.360 354.390 ;
        RECT 231.840 354.280 232.150 354.550 ;
        RECT 231.840 354.240 234.170 354.280 ;
        RECT 187.090 354.060 187.410 354.110 ;
        RECT 203.010 354.100 205.190 354.110 ;
        RECT 214.900 354.050 215.360 354.110 ;
        RECT 231.990 354.100 234.170 354.240 ;
        RECT 205.030 353.850 205.340 354.020 ;
        RECT 203.010 353.790 205.340 353.850 ;
        RECT 205.480 353.790 205.570 353.850 ;
        RECT 208.350 353.790 216.120 353.870 ;
        RECT 203.010 353.670 216.120 353.790 ;
        RECT 221.210 353.690 228.830 353.870 ;
        RECT 231.840 353.850 232.150 354.020 ;
        RECT 231.610 353.670 231.700 353.850 ;
        RECT 231.840 353.690 234.170 353.850 ;
        RECT 243.260 353.790 358.990 354.790 ;
        RECT 232.000 353.670 234.170 353.690 ;
        RECT 204.430 353.530 216.120 353.670 ;
        RECT 204.430 353.520 204.750 353.530 ;
        RECT 215.690 353.460 216.120 353.530 ;
        RECT 208.340 353.260 215.970 353.440 ;
        RECT 221.210 353.260 228.840 353.440 ;
        RECT 162.700 353.140 163.070 353.260 ;
        RECT 162.700 352.970 169.020 353.140 ;
        RECT 162.700 352.860 163.070 352.970 ;
        RECT 208.730 352.940 228.470 353.120 ;
        RECT 208.730 352.800 213.220 352.940 ;
        RECT 208.970 352.770 213.220 352.800 ;
        RECT 183.870 352.730 184.050 352.740 ;
        RECT 183.530 352.620 184.050 352.730 ;
        RECT 183.530 352.550 185.880 352.620 ;
        RECT 192.290 352.570 194.070 352.740 ;
        RECT 208.970 352.720 209.290 352.770 ;
        RECT 212.900 352.700 213.220 352.770 ;
        RECT 223.960 352.810 228.470 352.940 ;
        RECT 223.960 352.770 228.210 352.810 ;
        RECT 223.960 352.700 224.280 352.770 ;
        RECT 227.890 352.720 228.210 352.770 ;
        RECT 183.870 352.440 185.880 352.550 ;
        RECT 208.530 352.480 208.590 352.660 ;
        RECT 228.560 352.480 228.650 352.660 ;
        RECT 187.270 352.290 187.590 352.340 ;
        RECT 189.680 352.290 190.000 352.310 ;
        RECT 168.460 351.820 168.560 352.140 ;
        RECT 177.450 352.070 178.050 352.270 ;
        RECT 187.270 352.100 190.000 352.290 ;
        RECT 208.350 352.160 215.970 352.340 ;
        RECT 221.210 352.160 228.830 352.340 ;
        RECT 187.270 352.020 187.590 352.100 ;
        RECT 188.350 352.030 188.440 352.100 ;
        RECT 189.680 352.050 190.000 352.100 ;
        RECT 208.530 352.050 208.600 352.160 ;
        RECT 228.560 352.050 228.650 352.160 ;
        RECT 203.010 351.910 205.180 351.930 ;
        RECT 162.060 351.550 162.450 351.640 ;
        RECT 186.070 351.580 186.510 351.810 ;
        RECT 203.010 351.750 205.340 351.910 ;
        RECT 205.480 351.750 205.570 351.930 ;
        RECT 205.030 351.580 205.340 351.750 ;
        RECT 208.370 351.740 215.970 351.910 ;
        RECT 221.210 351.740 228.810 351.910 ;
        RECT 231.610 351.750 231.700 351.930 ;
        RECT 232.000 351.910 234.170 351.930 ;
        RECT 231.840 351.750 234.170 351.910 ;
        RECT 231.840 351.580 232.150 351.750 ;
        RECT 162.060 351.430 169.020 351.550 ;
        RECT 186.170 351.510 186.510 351.580 ;
        RECT 162.060 351.380 169.120 351.430 ;
        RECT 162.060 351.290 162.450 351.380 ;
        RECT 168.730 351.260 169.120 351.380 ;
        RECT 186.170 351.370 186.510 351.440 ;
        RECT 171.210 350.890 171.670 351.210 ;
        RECT 173.380 350.850 175.820 351.070 ;
        RECT 177.000 351.010 177.160 351.210 ;
        RECT 186.070 351.140 186.510 351.370 ;
        RECT 203.010 351.360 205.190 351.500 ;
        RECT 216.430 351.420 216.870 351.540 ;
        RECT 203.010 351.320 205.340 351.360 ;
        RECT 205.030 351.030 205.340 351.320 ;
        RECT 216.300 351.240 216.870 351.420 ;
        RECT 231.990 351.360 234.170 351.500 ;
        RECT 245.680 351.410 246.580 351.450 ;
        RECT 347.660 351.410 349.750 351.590 ;
        RECT 216.420 351.140 216.870 351.240 ;
        RECT 231.840 351.320 234.170 351.360 ;
        RECT 208.530 351.080 208.590 351.120 ;
        RECT 216.420 351.080 216.820 351.140 ;
        RECT 177.650 350.870 178.030 350.880 ;
        RECT 130.980 349.970 142.280 350.340 ;
        RECT 161.440 350.000 161.830 350.080 ;
        RECT 168.460 350.070 168.560 350.390 ;
        RECT 173.480 350.050 173.740 350.850 ;
        RECT 174.400 350.820 174.720 350.840 ;
        RECT 174.390 350.770 174.720 350.820 ;
        RECT 175.480 350.790 175.820 350.850 ;
        RECT 175.430 350.770 175.750 350.780 ;
        RECT 174.390 350.570 177.060 350.770 ;
        RECT 177.630 350.700 178.030 350.870 ;
        RECT 187.270 350.850 187.590 350.930 ;
        RECT 188.350 350.850 188.430 350.920 ;
        RECT 205.590 350.900 216.820 351.080 ;
        RECT 228.590 350.940 228.650 351.120 ;
        RECT 231.840 351.030 232.150 351.320 ;
        RECT 189.680 350.850 190.000 350.900 ;
        RECT 174.390 350.560 174.720 350.570 ;
        RECT 174.400 350.550 174.720 350.560 ;
        RECT 175.430 350.520 175.750 350.570 ;
        RECT 177.630 350.520 177.830 350.700 ;
        RECT 187.270 350.660 190.000 350.850 ;
        RECT 177.380 350.320 177.830 350.520 ;
        RECT 183.610 350.490 185.940 350.650 ;
        RECT 187.270 350.610 187.590 350.660 ;
        RECT 189.680 350.640 190.000 350.660 ;
        RECT 208.530 350.510 208.660 350.690 ;
        RECT 228.590 350.510 228.650 350.690 ;
        RECT 183.390 350.470 185.940 350.490 ;
        RECT 183.390 350.310 183.790 350.470 ;
        RECT 192.070 350.320 194.070 350.480 ;
        RECT 192.800 350.310 194.070 350.320 ;
        RECT 193.500 350.300 194.070 350.310 ;
        RECT 222.960 350.420 223.560 350.480 ;
        RECT 243.260 350.420 349.750 351.410 ;
        RECT 130.980 349.370 132.250 349.970 ;
        RECT 161.440 349.830 168.620 350.000 ;
        RECT 222.960 349.950 349.750 350.420 ;
        RECT 222.960 349.900 223.560 349.950 ;
        RECT 161.440 349.750 161.830 349.830 ;
        RECT 168.470 349.760 168.620 349.830 ;
        RECT 168.470 349.650 168.640 349.760 ;
        RECT 168.470 349.480 169.120 349.650 ;
        RECT 183.410 349.520 183.810 349.530 ;
        RECT 171.210 349.140 171.670 349.460 ;
        RECT 173.380 349.100 175.820 349.320 ;
        RECT 176.970 349.260 177.160 349.460 ;
        RECT 183.410 349.380 183.820 349.520 ;
        RECT 183.410 349.370 185.920 349.380 ;
        RECT 183.640 349.200 185.920 349.370 ;
        RECT 192.290 349.360 194.070 349.520 ;
        RECT 208.530 349.240 208.600 349.420 ;
        RECT 228.560 349.240 228.650 349.420 ;
        RECT 243.260 349.320 349.750 349.950 ;
        RECT 160.830 348.520 161.250 348.610 ;
        RECT 168.460 348.520 168.560 348.640 ;
        RECT 160.830 348.350 168.640 348.520 ;
        RECT 160.830 348.250 161.250 348.350 ;
        RECT 168.460 348.320 168.640 348.350 ;
        RECT 168.470 347.860 168.640 348.320 ;
        RECT 173.480 348.300 173.740 349.100 ;
        RECT 174.400 349.070 174.720 349.090 ;
        RECT 174.390 349.020 174.720 349.070 ;
        RECT 175.480 349.040 175.820 349.100 ;
        RECT 187.270 349.090 187.590 349.140 ;
        RECT 189.680 349.090 190.000 349.110 ;
        RECT 175.430 349.020 175.750 349.030 ;
        RECT 174.390 348.820 177.060 349.020 ;
        RECT 177.580 348.920 178.030 349.050 ;
        RECT 174.390 348.810 174.720 348.820 ;
        RECT 174.400 348.800 174.720 348.810 ;
        RECT 175.430 348.770 175.750 348.820 ;
        RECT 177.580 348.770 178.070 348.920 ;
        RECT 187.270 348.900 190.000 349.090 ;
        RECT 187.270 348.820 187.590 348.900 ;
        RECT 188.350 348.820 188.500 348.900 ;
        RECT 189.680 348.850 190.000 348.900 ;
        RECT 177.380 348.720 178.070 348.770 ;
        RECT 177.380 348.570 177.930 348.720 ;
        RECT 205.630 348.680 205.940 348.970 ;
        RECT 208.530 348.810 208.600 348.990 ;
        RECT 228.560 348.810 228.650 348.990 ;
        RECT 203.610 348.640 205.940 348.680 ;
        RECT 186.070 348.380 186.510 348.610 ;
        RECT 203.610 348.500 205.790 348.640 ;
        RECT 186.170 348.310 186.510 348.380 ;
        RECT 205.630 348.250 205.940 348.420 ;
        RECT 215.230 348.320 221.990 348.500 ;
        RECT 186.170 348.170 186.510 348.240 ;
        RECT 186.070 347.940 186.510 348.170 ;
        RECT 203.610 348.090 205.940 348.250 ;
        RECT 203.610 348.070 205.780 348.090 ;
        RECT 206.080 348.070 206.170 348.250 ;
        RECT 206.500 348.090 206.590 348.270 ;
        RECT 168.470 347.690 169.120 347.860 ;
        RECT 171.210 347.390 171.670 347.710 ;
        RECT 173.380 347.350 175.820 347.570 ;
        RECT 176.990 347.510 177.160 347.710 ;
        RECT 130.920 346.190 132.190 347.030 ;
        RECT 168.460 346.570 168.560 346.890 ;
        RECT 173.480 346.550 173.740 347.350 ;
        RECT 174.400 347.320 174.720 347.340 ;
        RECT 174.390 347.270 174.720 347.320 ;
        RECT 175.480 347.290 175.820 347.350 ;
        RECT 177.620 347.500 178.050 347.730 ;
        RECT 187.270 347.650 187.590 347.730 ;
        RECT 188.350 347.650 188.430 347.720 ;
        RECT 189.680 347.650 190.000 347.700 ;
        RECT 206.500 347.660 206.590 347.840 ;
        RECT 208.530 347.710 208.600 347.890 ;
        RECT 208.960 347.650 216.570 347.840 ;
        RECT 228.560 347.710 228.650 347.890 ;
        RECT 175.430 347.270 175.750 347.280 ;
        RECT 174.390 347.070 177.060 347.270 ;
        RECT 174.390 347.060 174.720 347.070 ;
        RECT 174.400 347.050 174.720 347.060 ;
        RECT 175.430 347.020 175.750 347.070 ;
        RECT 177.620 347.020 177.820 347.500 ;
        RECT 187.270 347.460 190.000 347.650 ;
        RECT 183.600 347.240 185.900 347.420 ;
        RECT 187.270 347.410 187.590 347.460 ;
        RECT 189.680 347.440 190.000 347.460 ;
        RECT 208.530 347.280 208.600 347.460 ;
        RECT 228.560 347.280 228.650 347.460 ;
        RECT 183.600 347.230 183.800 347.240 ;
        RECT 183.390 347.050 183.800 347.230 ;
        RECT 192.290 347.040 194.070 347.220 ;
        RECT 177.380 346.820 177.820 347.020 ;
        RECT 206.500 346.570 206.590 346.750 ;
        RECT 208.940 346.570 216.570 346.750 ;
        RECT 146.090 346.450 146.400 346.470 ;
        RECT 146.750 346.450 147.060 346.470 ;
        RECT 130.920 345.820 140.620 346.190 ;
        RECT 146.090 345.980 153.410 346.450 ;
        RECT 146.090 345.960 146.400 345.980 ;
        RECT 146.750 345.960 147.060 345.980 ;
        RECT 130.920 345.150 132.190 345.820 ;
        RECT 140.250 344.470 140.620 345.820 ;
        RECT 152.940 345.300 153.410 345.980 ;
        RECT 179.710 346.310 180.020 346.330 ;
        RECT 203.610 346.320 205.780 346.340 ;
        RECT 203.610 346.310 205.940 346.320 ;
        RECT 206.080 346.310 206.170 346.340 ;
        RECT 206.500 346.310 206.590 346.320 ;
        RECT 217.350 346.310 217.800 346.340 ;
        RECT 171.210 345.640 171.670 345.960 ;
        RECT 173.380 345.600 175.820 345.820 ;
        RECT 177.000 345.760 177.160 345.960 ;
        RECT 179.710 345.900 217.800 346.310 ;
        RECT 245.710 346.010 246.610 346.270 ;
        RECT 179.710 345.880 180.020 345.900 ;
        RECT 203.610 345.770 205.790 345.900 ;
        RECT 217.350 345.880 217.800 345.900 ;
        RECT 203.610 345.730 205.940 345.770 ;
        RECT 173.480 345.300 173.740 345.600 ;
        RECT 174.400 345.570 174.720 345.590 ;
        RECT 174.390 345.520 174.720 345.570 ;
        RECT 175.480 345.540 175.820 345.600 ;
        RECT 175.430 345.520 175.750 345.530 ;
        RECT 174.390 345.320 177.060 345.520 ;
        RECT 205.630 345.440 205.940 345.730 ;
        RECT 203.610 345.400 205.940 345.440 ;
        RECT 174.390 345.310 174.720 345.320 ;
        RECT 174.400 345.300 174.720 345.310 ;
        RECT 175.430 345.300 175.750 345.320 ;
        RECT 203.610 345.300 205.790 345.400 ;
        RECT 243.260 345.300 345.610 346.010 ;
        RECT 144.760 345.170 145.020 345.240 ;
        RECT 146.810 345.170 147.130 345.190 ;
        RECT 148.570 345.170 148.900 345.210 ;
        RECT 144.760 344.980 148.900 345.170 ;
        RECT 144.760 344.920 145.020 344.980 ;
        RECT 146.810 344.930 147.130 344.980 ;
        RECT 148.570 344.940 148.900 344.980 ;
        RECT 152.940 344.830 345.610 345.300 ;
        RECT 144.210 344.770 144.530 344.810 ;
        RECT 146.150 344.770 146.470 344.830 ;
        RECT 149.070 344.770 149.390 344.810 ;
        RECT 173.480 344.800 173.740 344.830 ;
        RECT 144.210 344.580 149.390 344.770 ;
        RECT 221.870 344.710 222.440 344.830 ;
        RECT 144.210 344.550 144.530 344.580 ;
        RECT 146.150 344.570 146.470 344.580 ;
        RECT 149.070 344.550 149.390 344.580 ;
        RECT 140.250 344.460 142.280 344.470 ;
        RECT 140.250 344.280 142.500 344.460 ;
        RECT 206.500 344.420 206.610 344.600 ;
        RECT 208.940 344.430 215.800 344.600 ;
        RECT 216.100 344.460 216.570 344.620 ;
        RECT 216.100 344.450 216.560 344.460 ;
        RECT 140.250 344.220 143.900 344.280 ;
        RECT 140.250 344.100 145.230 344.220 ;
        RECT 150.550 344.210 150.850 344.230 ;
        RECT 150.540 344.190 150.860 344.210 ;
        RECT 141.910 344.060 145.230 344.100 ;
        RECT 142.280 344.000 145.230 344.060 ;
        RECT 134.910 343.810 135.680 344.000 ;
        RECT 148.320 343.970 150.860 344.190 ;
        RECT 141.910 343.810 142.300 343.830 ;
        RECT 134.910 343.770 142.300 343.810 ;
        RECT 134.910 343.560 145.220 343.770 ;
        RECT 134.910 343.440 142.290 343.560 ;
        RECT 148.320 343.530 148.540 343.970 ;
        RECT 150.540 343.950 150.860 343.970 ;
        RECT 150.550 343.930 150.850 343.950 ;
        RECT 168.660 343.890 169.080 344.060 ;
        RECT 209.690 344.030 210.010 344.090 ;
        RECT 213.710 344.030 214.040 344.060 ;
        RECT 168.660 343.790 169.040 343.890 ;
        RECT 209.690 343.860 214.040 344.030 ;
        RECT 243.260 343.920 345.610 344.830 ;
        RECT 168.660 343.570 168.940 343.790 ;
        RECT 208.590 343.680 209.320 343.860 ;
        RECT 209.690 343.810 210.010 343.860 ;
        RECT 211.990 343.840 212.310 343.860 ;
        RECT 213.710 343.840 214.040 343.860 ;
        RECT 211.990 343.700 219.820 343.840 ;
        RECT 212.170 343.650 219.820 343.700 ;
        RECT 212.170 343.640 219.990 343.650 ;
        RECT 208.940 343.630 219.990 343.640 ;
        RECT 134.910 343.260 135.680 343.440 ;
        RECT 141.910 343.420 142.280 343.440 ;
        RECT 160.190 343.350 160.600 343.450 ;
        RECT 168.660 343.350 168.930 343.570 ;
        RECT 160.190 343.180 168.930 343.350 ;
        RECT 183.420 343.290 183.730 343.470 ;
        RECT 192.320 343.300 194.100 343.470 ;
        RECT 206.500 343.320 206.610 343.500 ;
        RECT 208.940 343.470 216.570 343.630 ;
        RECT 219.610 343.440 219.990 343.630 ;
        RECT 219.100 343.430 219.240 343.440 ;
        RECT 160.190 343.090 160.600 343.180 ;
        RECT 168.660 343.170 168.830 343.180 ;
        RECT 149.930 343.060 150.220 343.080 ;
        RECT 149.920 343.030 150.240 343.060 ;
        RECT 149.680 343.020 151.670 343.030 ;
        RECT 130.980 342.160 132.250 342.930 ;
        RECT 148.350 342.830 151.670 343.020 ;
        RECT 152.520 342.920 153.210 343.000 ;
        RECT 149.680 342.810 151.670 342.830 ;
        RECT 149.920 342.800 150.240 342.810 ;
        RECT 149.930 342.780 150.220 342.800 ;
        RECT 151.710 342.590 152.020 342.920 ;
        RECT 152.360 342.790 153.210 342.920 ;
        RECT 152.360 342.590 152.670 342.790 ;
        RECT 168.420 342.760 168.520 343.080 ;
        RECT 177.340 343.010 177.950 343.210 ;
        RECT 183.550 343.110 185.900 343.290 ;
        RECT 203.610 343.070 205.780 343.090 ;
        RECT 177.750 342.970 177.950 343.010 ;
        RECT 187.300 343.020 187.620 343.070 ;
        RECT 189.710 343.020 190.030 343.040 ;
        RECT 177.750 342.770 178.170 342.970 ;
        RECT 187.300 342.830 190.030 343.020 ;
        RECT 203.610 342.910 205.940 343.070 ;
        RECT 206.080 342.910 206.170 343.090 ;
        RECT 187.300 342.750 187.620 342.830 ;
        RECT 188.380 342.760 188.470 342.830 ;
        RECT 189.710 342.780 190.030 342.830 ;
        RECT 205.630 342.740 205.940 342.910 ;
        RECT 206.500 342.890 206.610 343.070 ;
        RECT 208.630 342.800 208.780 343.220 ;
        RECT 219.100 343.100 219.250 343.430 ;
        RECT 208.630 342.710 211.900 342.800 ;
        RECT 211.970 342.710 212.290 342.910 ;
        RECT 219.100 342.900 220.310 343.100 ;
        RECT 149.680 342.370 150.390 342.580 ;
        RECT 151.340 342.480 153.210 342.560 ;
        RECT 184.190 342.480 185.360 342.630 ;
        RECT 130.980 341.790 136.970 342.160 ;
        RECT 150.490 342.150 150.800 342.480 ;
        RECT 151.190 342.340 153.210 342.480 ;
        RECT 151.190 342.150 151.500 342.340 ;
        RECT 168.600 342.130 169.080 342.300 ;
        RECT 184.130 342.150 184.410 342.480 ;
        RECT 186.100 342.310 186.540 342.540 ;
        RECT 203.610 342.520 205.790 342.660 ;
        RECT 208.630 342.650 212.290 342.710 ;
        RECT 220.420 342.670 220.540 342.880 ;
        RECT 220.810 342.770 221.120 343.030 ;
        RECT 221.450 342.790 222.710 342.950 ;
        RECT 211.760 342.550 212.060 342.650 ;
        RECT 220.660 342.610 223.250 342.770 ;
        RECT 203.610 342.480 205.940 342.520 ;
        RECT 186.200 342.240 186.540 342.310 ;
        RECT 205.630 342.190 205.940 342.480 ;
        RECT 220.660 342.440 220.970 342.610 ;
        RECT 208.700 342.320 209.020 342.410 ;
        RECT 36.770 339.000 127.730 341.080 ;
        RECT 130.980 341.050 132.250 341.790 ;
        RECT 136.600 340.130 136.970 341.790 ;
        RECT 152.730 341.840 153.050 341.900 ;
        RECT 152.730 341.630 153.210 341.840 ;
        RECT 159.530 341.780 159.920 341.890 ;
        RECT 168.600 341.840 168.770 342.130 ;
        RECT 168.600 341.780 168.760 341.840 ;
        RECT 171.170 341.830 171.630 342.150 ;
        RECT 173.340 341.790 175.780 342.010 ;
        RECT 176.960 341.950 177.120 342.150 ;
        RECT 186.200 342.100 186.540 342.170 ;
        RECT 186.100 341.870 186.540 342.100 ;
        RECT 208.610 342.150 209.020 342.320 ;
        RECT 219.210 342.240 220.410 342.340 ;
        RECT 219.200 342.160 220.410 342.240 ;
        RECT 208.610 342.050 208.930 342.150 ;
        RECT 220.130 342.040 220.410 342.160 ;
        RECT 220.660 342.180 220.970 342.350 ;
        RECT 220.130 342.020 220.160 342.040 ;
        RECT 220.420 341.910 220.540 342.120 ;
        RECT 220.660 342.020 223.250 342.180 ;
        RECT 152.730 341.580 153.050 341.630 ;
        RECT 159.530 341.620 168.760 341.780 ;
        RECT 159.530 341.610 168.410 341.620 ;
        RECT 159.530 341.510 159.920 341.610 ;
        RECT 149.680 341.010 149.930 341.230 ;
        RECT 144.240 340.900 144.530 340.910 ;
        RECT 144.230 340.880 144.550 340.900 ;
        RECT 149.990 340.890 150.310 341.150 ;
        RECT 168.420 341.010 168.520 341.330 ;
        RECT 173.440 340.990 173.700 341.790 ;
        RECT 174.360 341.760 174.680 341.780 ;
        RECT 174.350 341.710 174.680 341.760 ;
        RECT 175.440 341.730 175.780 341.790 ;
        RECT 208.560 341.730 209.140 341.910 ;
        RECT 220.810 341.760 221.120 342.020 ;
        RECT 221.450 341.860 222.710 342.020 ;
        RECT 175.390 341.710 175.710 341.720 ;
        RECT 174.350 341.510 177.020 341.710 ;
        RECT 174.350 341.500 174.680 341.510 ;
        RECT 174.360 341.490 174.680 341.500 ;
        RECT 175.390 341.460 175.710 341.510 ;
        RECT 177.740 341.460 178.060 341.620 ;
        RECT 177.340 341.260 178.060 341.460 ;
        RECT 187.300 341.580 187.620 341.660 ;
        RECT 188.380 341.580 188.460 341.650 ;
        RECT 189.710 341.580 190.030 341.630 ;
        RECT 187.300 341.390 190.030 341.580 ;
        RECT 211.840 341.570 212.070 341.580 ;
        RECT 211.840 341.540 219.410 341.570 ;
        RECT 187.300 341.340 187.620 341.390 ;
        RECT 189.710 341.370 190.030 341.390 ;
        RECT 183.530 341.210 185.320 341.340 ;
        RECT 208.680 341.270 209.000 341.400 ;
        RECT 211.840 341.370 219.470 341.540 ;
        RECT 211.840 341.270 212.080 341.370 ;
        RECT 183.390 341.160 185.320 341.210 ;
        RECT 183.390 341.010 183.710 341.160 ;
        RECT 192.100 341.050 194.100 341.210 ;
        RECT 208.630 341.090 212.080 341.270 ;
        RECT 219.280 341.170 219.990 341.370 ;
        RECT 245.680 341.130 246.580 341.190 ;
        RECT 208.630 341.070 212.000 341.090 ;
        RECT 192.830 341.040 194.100 341.050 ;
        RECT 193.530 341.030 194.100 341.040 ;
        RECT 183.390 340.930 183.570 341.010 ;
        RECT 211.970 340.890 212.290 341.030 ;
        RECT 144.230 340.660 145.230 340.880 ;
        RECT 211.970 340.870 219.430 340.890 ;
        RECT 211.970 340.770 219.990 340.870 ;
        RECT 144.230 340.640 144.550 340.660 ;
        RECT 152.390 340.650 152.710 340.680 ;
        RECT 211.980 340.670 219.990 340.770 ;
        RECT 211.980 340.660 212.300 340.670 ;
        RECT 144.240 340.620 144.530 340.640 ;
        RECT 149.680 340.470 152.710 340.650 ;
        RECT 149.500 340.440 152.710 340.470 ;
        RECT 149.500 340.420 149.820 340.440 ;
        RECT 148.330 340.250 149.820 340.420 ;
        RECT 152.390 340.360 152.710 340.440 ;
        RECT 168.520 340.320 169.080 340.490 ;
        RECT 208.590 340.440 209.140 340.620 ;
        RECT 168.520 340.280 168.690 340.320 ;
        RECT 148.330 340.210 152.660 340.250 ;
        RECT 149.500 340.170 152.660 340.210 ;
        RECT 149.680 340.140 152.660 340.170 ;
        RECT 158.920 340.240 159.290 340.250 ;
        RECT 168.520 340.240 168.680 340.280 ;
        RECT 136.600 339.950 142.550 340.130 ;
        RECT 149.680 340.040 152.720 340.140 ;
        RECT 136.600 339.880 142.620 339.950 ;
        RECT 144.010 339.880 145.230 339.890 ;
        RECT 151.190 339.880 151.480 339.900 ;
        RECT 136.600 339.760 145.230 339.880 ;
        RECT 151.180 339.850 151.500 339.880 ;
        RECT 141.910 339.720 145.230 339.760 ;
        RECT 142.270 339.670 145.230 339.720 ;
        RECT 148.330 339.640 151.500 339.850 ;
        RECT 152.400 339.820 152.720 340.040 ;
        RECT 158.920 340.070 168.680 340.240 ;
        RECT 171.170 340.080 171.630 340.400 ;
        RECT 158.920 339.860 159.290 340.070 ;
        RECT 173.340 340.040 175.780 340.260 ;
        RECT 176.930 340.200 177.120 340.400 ;
        RECT 183.440 340.100 183.640 340.260 ;
        RECT 140.140 339.150 140.550 339.170 ;
        RECT 141.910 339.150 143.900 339.170 ;
        RECT 140.140 339.110 143.900 339.150 ;
        RECT 36.770 247.590 38.850 339.000 ;
        RECT 140.140 338.890 145.230 339.110 ;
        RECT 130.980 338.020 132.250 338.840 ;
        RECT 140.140 338.780 142.290 338.890 ;
        RECT 148.330 338.820 148.540 339.640 ;
        RECT 149.680 339.470 149.930 339.640 ;
        RECT 151.180 339.620 151.500 339.640 ;
        RECT 151.190 339.600 151.480 339.620 ;
        RECT 149.990 339.340 150.310 339.600 ;
        RECT 152.710 339.230 153.030 339.280 ;
        RECT 168.420 339.260 168.520 339.580 ;
        RECT 173.440 339.240 173.700 340.040 ;
        RECT 174.360 340.010 174.680 340.030 ;
        RECT 174.350 339.960 174.680 340.010 ;
        RECT 175.440 339.980 175.780 340.040 ;
        RECT 183.460 340.050 183.640 340.100 ;
        RECT 192.320 340.090 194.100 340.250 ;
        RECT 175.390 339.960 175.710 339.970 ;
        RECT 174.350 339.760 177.020 339.960 ;
        RECT 183.460 339.870 185.350 340.050 ;
        RECT 187.300 339.820 187.620 339.870 ;
        RECT 189.710 339.820 190.030 339.840 ;
        RECT 174.350 339.750 174.680 339.760 ;
        RECT 174.360 339.740 174.680 339.750 ;
        RECT 175.390 339.710 175.710 339.760 ;
        RECT 177.340 339.690 178.030 339.710 ;
        RECT 177.340 339.510 178.110 339.690 ;
        RECT 177.820 339.420 178.110 339.510 ;
        RECT 184.740 339.640 185.060 339.680 ;
        RECT 184.740 339.430 185.350 339.640 ;
        RECT 187.300 339.630 190.030 339.820 ;
        RECT 187.300 339.550 187.620 339.630 ;
        RECT 188.380 339.550 188.530 339.630 ;
        RECT 189.710 339.580 190.030 339.630 ;
        RECT 208.570 339.710 208.770 340.210 ;
        RECT 219.190 340.050 220.190 340.210 ;
        RECT 220.420 339.900 220.540 340.110 ;
        RECT 220.810 340.070 221.120 340.260 ;
        RECT 220.750 340.060 221.300 340.070 ;
        RECT 220.750 340.040 221.310 340.060 ;
        RECT 221.450 340.040 222.710 340.180 ;
        RECT 243.260 340.040 341.530 341.130 ;
        RECT 220.750 340.000 341.530 340.040 ;
        RECT 211.840 339.710 212.160 339.850 ;
        RECT 208.570 339.590 212.160 339.710 ;
        RECT 220.660 339.690 341.530 340.000 ;
        RECT 208.570 339.510 212.120 339.590 ;
        RECT 215.910 339.570 341.530 339.690 ;
        RECT 215.910 339.520 222.590 339.570 ;
        RECT 184.740 339.360 185.200 339.430 ;
        RECT 152.710 339.020 153.210 339.230 ;
        RECT 186.100 339.110 186.540 339.340 ;
        RECT 208.680 339.270 208.990 339.450 ;
        RECT 220.660 339.410 220.970 339.520 ;
        RECT 222.260 339.490 222.590 339.520 ;
        RECT 186.200 339.040 186.540 339.110 ;
        RECT 208.560 339.120 208.990 339.270 ;
        RECT 152.710 338.960 153.030 339.020 ;
        RECT 208.560 339.000 208.840 339.120 ;
        RECT 219.200 339.070 220.200 339.240 ;
        RECT 220.420 339.140 220.540 339.350 ;
        RECT 220.660 339.250 223.250 339.410 ;
        RECT 219.200 339.060 220.140 339.070 ;
        RECT 220.810 338.990 221.120 339.250 ;
        RECT 221.470 339.090 222.710 339.250 ;
        RECT 243.260 339.040 341.530 339.570 ;
        RECT 186.200 338.900 186.540 338.970 ;
        RECT 140.140 338.760 140.550 338.780 ;
        RECT 141.910 338.760 142.280 338.780 ;
        RECT 158.230 338.700 158.620 338.800 ;
        RECT 168.430 338.700 169.080 338.770 ;
        RECT 149.680 338.690 149.950 338.700 ;
        RECT 149.680 338.480 150.430 338.690 ;
        RECT 134.910 338.020 135.710 338.160 ;
        RECT 147.560 338.130 148.160 338.280 ;
        RECT 150.520 338.270 150.830 338.600 ;
        RECT 151.380 338.590 153.210 338.670 ;
        RECT 151.210 338.460 153.210 338.590 ;
        RECT 158.230 338.600 169.080 338.700 ;
        RECT 186.100 338.670 186.540 338.900 ;
        RECT 158.230 338.530 168.720 338.600 ;
        RECT 151.210 338.260 151.520 338.460 ;
        RECT 158.230 338.430 158.620 338.530 ;
        RECT 168.550 338.510 168.720 338.530 ;
        RECT 171.170 338.330 171.630 338.650 ;
        RECT 173.340 338.290 175.780 338.510 ;
        RECT 176.950 338.450 177.120 338.650 ;
        RECT 177.800 338.540 178.100 338.580 ;
        RECT 130.980 337.520 135.710 338.020 ;
        RECT 144.020 337.830 146.730 337.840 ;
        RECT 130.980 336.960 132.250 337.520 ;
        RECT 134.910 337.390 135.710 337.520 ;
        RECT 143.790 337.510 146.730 337.830 ;
        RECT 147.410 337.800 148.160 338.130 ;
        RECT 147.560 337.660 148.160 337.800 ;
        RECT 149.680 337.700 151.640 337.920 ;
        RECT 143.790 337.360 144.410 337.510 ;
        RECT 145.200 337.370 145.510 337.510 ;
        RECT 146.290 337.370 146.600 337.510 ;
        RECT 147.420 337.460 148.160 337.660 ;
        RECT 151.690 337.490 152.000 337.820 ;
        RECT 152.530 337.760 153.210 337.840 ;
        RECT 152.400 337.630 153.210 337.760 ;
        RECT 41.120 334.740 127.730 336.820 ;
        RECT 143.790 335.890 144.140 337.360 ;
        RECT 147.420 337.330 147.730 337.460 ;
        RECT 152.400 337.430 152.710 337.630 ;
        RECT 168.420 337.510 168.520 337.830 ;
        RECT 173.440 337.490 173.700 338.290 ;
        RECT 174.360 338.260 174.680 338.280 ;
        RECT 174.350 338.210 174.680 338.260 ;
        RECT 175.440 338.230 175.780 338.290 ;
        RECT 177.790 338.300 178.100 338.540 ;
        RECT 208.570 338.480 209.140 338.660 ;
        RECT 219.430 338.610 219.980 338.620 ;
        RECT 187.300 338.380 187.620 338.460 ;
        RECT 188.380 338.380 188.460 338.450 ;
        RECT 189.710 338.380 190.030 338.430 ;
        RECT 175.390 338.210 175.710 338.220 ;
        RECT 174.350 338.010 177.020 338.210 ;
        RECT 174.350 338.000 174.680 338.010 ;
        RECT 174.360 337.990 174.680 338.000 ;
        RECT 175.390 337.960 175.710 338.010 ;
        RECT 177.790 337.960 177.990 338.300 ;
        RECT 187.300 338.190 190.030 338.380 ;
        RECT 208.730 338.330 209.040 338.480 ;
        RECT 187.300 338.140 187.620 338.190 ;
        RECT 189.710 338.170 190.030 338.190 ;
        RECT 208.610 338.200 209.040 338.330 ;
        RECT 211.850 338.390 219.980 338.610 ;
        RECT 211.850 338.380 219.440 338.390 ;
        RECT 211.850 338.370 212.620 338.380 ;
        RECT 211.850 338.200 212.090 338.370 ;
        RECT 208.610 338.120 212.090 338.200 ;
        RECT 183.700 337.960 185.330 338.090 ;
        RECT 208.720 337.960 212.090 338.120 ;
        RECT 177.340 337.760 177.990 337.960 ;
        RECT 183.390 337.910 185.330 337.960 ;
        RECT 183.390 337.780 183.880 337.910 ;
        RECT 192.320 337.770 194.100 337.950 ;
        RECT 177.530 337.260 177.850 337.310 ;
        RECT 184.140 337.260 184.460 337.360 ;
        RECT 144.760 337.020 147.920 337.160 ;
        RECT 177.530 337.100 184.460 337.260 ;
        RECT 177.530 337.050 177.850 337.100 ;
        RECT 184.140 337.080 184.460 337.100 ;
        RECT 185.170 337.240 185.490 337.550 ;
        RECT 195.790 337.260 196.200 337.370 ;
        RECT 188.820 337.240 196.200 337.260 ;
        RECT 185.170 337.100 196.200 337.240 ;
        RECT 185.170 337.070 185.490 337.100 ;
        RECT 188.740 337.030 196.200 337.100 ;
        RECT 184.730 337.020 185.010 337.030 ;
        RECT 144.650 336.840 147.920 337.020 ;
        RECT 177.000 336.970 177.330 336.990 ;
        RECT 176.990 336.900 177.340 336.970 ;
        RECT 144.650 336.690 144.960 336.840 ;
        RECT 145.750 336.690 146.060 336.840 ;
        RECT 146.850 336.690 147.160 336.840 ;
        RECT 147.600 335.890 147.920 336.840 ;
        RECT 171.170 336.580 171.630 336.900 ;
        RECT 176.960 336.890 177.340 336.900 ;
        RECT 182.740 336.890 183.060 336.950 ;
        RECT 184.710 336.930 185.030 337.020 ;
        RECT 195.790 337.000 196.200 337.030 ;
        RECT 225.940 337.230 226.500 337.300 ;
        RECT 238.660 337.230 239.340 337.290 ;
        RECT 246.190 337.230 246.850 337.870 ;
        RECT 186.950 336.930 187.270 336.960 ;
        RECT 173.340 336.540 175.780 336.760 ;
        RECT 176.960 336.730 183.060 336.890 ;
        RECT 184.680 336.770 187.270 336.930 ;
        RECT 225.940 336.820 246.850 337.230 ;
        RECT 225.940 336.770 226.500 336.820 ;
        RECT 184.710 336.760 185.030 336.770 ;
        RECT 184.730 336.750 185.010 336.760 ;
        RECT 176.960 336.700 177.340 336.730 ;
        RECT 176.990 336.660 177.340 336.700 ;
        RECT 182.740 336.680 183.060 336.730 ;
        RECT 186.950 336.700 187.270 336.770 ;
        RECT 238.660 336.760 239.340 336.820 ;
        RECT 246.190 336.720 246.850 336.820 ;
        RECT 186.970 336.690 187.250 336.700 ;
        RECT 172.570 336.270 172.900 336.510 ;
        RECT 173.440 336.270 173.700 336.540 ;
        RECT 174.360 336.510 174.680 336.530 ;
        RECT 174.350 336.460 174.680 336.510 ;
        RECT 175.440 336.480 175.780 336.540 ;
        RECT 175.390 336.460 175.710 336.470 ;
        RECT 174.350 336.270 177.020 336.460 ;
        RECT 178.430 336.400 178.730 336.410 ;
        RECT 178.420 336.270 178.740 336.400 ;
        RECT 188.960 336.270 189.240 336.570 ;
        RECT 192.990 336.270 193.290 336.550 ;
        RECT 172.570 336.250 193.290 336.270 ;
        RECT 172.570 336.220 193.280 336.250 ;
        RECT 172.570 336.110 193.220 336.220 ;
        RECT 173.440 335.890 173.700 336.110 ;
        RECT 176.380 335.890 176.820 335.900 ;
        RECT 131.060 335.880 176.820 335.890 ;
        RECT 131.060 335.470 176.840 335.880 ;
        RECT 143.790 335.070 144.140 335.470 ;
        RECT 144.650 335.320 144.960 335.470 ;
        RECT 145.750 335.320 146.060 335.470 ;
        RECT 146.850 335.320 147.160 335.470 ;
        RECT 143.790 334.920 146.740 335.070 ;
        RECT 147.600 334.920 147.920 335.470 ;
        RECT 169.530 335.460 170.010 335.470 ;
        RECT 176.360 335.460 176.840 335.470 ;
        RECT 176.380 335.450 176.820 335.460 ;
        RECT 185.750 335.420 186.130 335.810 ;
        RECT 201.830 335.800 202.130 335.820 ;
        RECT 186.900 335.380 187.300 335.720 ;
        RECT 195.490 335.220 196.150 335.580 ;
        RECT 201.120 335.460 202.140 335.800 ;
        RECT 201.830 335.440 202.140 335.460 ;
        RECT 36.610 244.020 39.000 247.590 ;
        RECT 36.770 243.490 38.850 244.020 ;
        RECT 41.120 218.980 43.200 334.740 ;
        RECT 131.040 334.500 173.020 334.920 ;
        RECT 143.790 333.870 144.140 334.500 ;
        RECT 143.790 333.740 144.170 333.870 ;
        RECT 143.790 333.700 144.540 333.740 ;
        RECT 130.920 332.910 132.190 333.690 ;
        RECT 143.790 333.400 146.730 333.700 ;
        RECT 144.090 333.250 144.400 333.400 ;
        RECT 145.200 333.240 145.510 333.400 ;
        RECT 146.290 333.220 146.600 333.400 ;
        RECT 147.600 333.020 147.920 334.500 ;
        RECT 154.090 334.000 154.920 334.500 ;
        RECT 177.050 334.380 177.430 334.760 ;
        RECT 197.240 334.500 197.690 334.930 ;
        RECT 219.700 334.740 220.300 334.790 ;
        RECT 243.260 334.740 337.440 335.930 ;
        RECT 219.700 334.270 337.440 334.740 ;
        RECT 219.700 334.230 220.300 334.270 ;
        RECT 243.260 333.840 337.440 334.270 ;
        RECT 246.110 333.600 248.210 333.840 ;
        RECT 246.130 333.590 246.900 333.600 ;
        RECT 140.150 332.910 140.560 332.930 ;
        RECT 45.460 330.670 127.730 332.750 ;
        RECT 130.920 332.540 140.560 332.910 ;
        RECT 144.770 332.880 147.920 333.020 ;
        RECT 144.650 332.690 147.920 332.880 ;
        RECT 144.650 332.680 147.830 332.690 ;
        RECT 144.650 332.550 144.960 332.680 ;
        RECT 145.750 332.540 146.060 332.680 ;
        RECT 146.840 332.540 147.150 332.680 ;
        RECT 130.920 331.810 132.190 332.540 ;
        RECT 140.150 332.520 140.560 332.540 ;
        RECT 147.680 332.480 147.970 332.500 ;
        RECT 149.910 332.480 150.220 332.500 ;
        RECT 147.670 332.120 150.220 332.480 ;
        RECT 147.680 332.100 147.970 332.120 ;
        RECT 149.910 332.100 150.220 332.120 ;
        RECT 177.330 331.590 177.640 331.730 ;
        RECT 178.420 331.590 178.730 331.730 ;
        RECT 179.520 331.590 179.830 331.720 ;
        RECT 176.650 331.580 179.830 331.590 ;
        RECT 176.560 331.390 179.830 331.580 ;
        RECT 183.370 331.590 183.680 331.720 ;
        RECT 184.470 331.590 184.780 331.730 ;
        RECT 185.560 331.590 185.870 331.730 ;
        RECT 187.140 331.620 187.450 331.760 ;
        RECT 188.230 331.620 188.540 331.760 ;
        RECT 189.330 331.620 189.640 331.750 ;
        RECT 186.460 331.610 189.640 331.620 ;
        RECT 186.370 331.590 189.640 331.610 ;
        RECT 183.370 331.420 189.640 331.590 ;
        RECT 193.180 331.620 193.490 331.750 ;
        RECT 194.280 331.620 194.590 331.760 ;
        RECT 195.370 331.620 195.680 331.760 ;
        RECT 193.180 331.610 196.360 331.620 ;
        RECT 193.180 331.420 196.450 331.610 ;
        RECT 183.370 331.390 189.520 331.420 ;
        RECT 176.560 331.250 179.710 331.390 ;
        RECT 183.490 331.280 189.520 331.390 ;
        RECT 193.300 331.280 196.450 331.420 ;
        RECT 198.920 331.600 199.230 331.730 ;
        RECT 200.020 331.600 200.330 331.740 ;
        RECT 201.110 331.600 201.420 331.740 ;
        RECT 198.920 331.590 202.100 331.600 ;
        RECT 198.920 331.400 202.190 331.590 ;
        RECT 183.490 331.250 186.690 331.280 ;
        RECT 40.940 215.460 43.390 218.980 ;
        RECT 41.120 215.340 43.200 215.460 ;
        RECT 45.460 190.470 47.540 330.670 ;
        RECT 147.600 330.570 148.200 330.720 ;
        RECT 144.060 330.270 146.770 330.280 ;
        RECT 143.830 329.950 146.770 330.270 ;
        RECT 147.450 330.240 148.200 330.570 ;
        RECT 147.600 330.100 148.200 330.240 ;
        RECT 143.830 329.800 144.450 329.950 ;
        RECT 145.240 329.810 145.550 329.950 ;
        RECT 146.330 329.810 146.640 329.950 ;
        RECT 147.460 329.900 148.200 330.100 ;
        RECT 141.870 329.520 142.240 329.530 ;
        RECT 130.980 328.700 132.250 329.400 ;
        RECT 140.550 329.140 143.160 329.520 ;
        RECT 140.550 328.700 140.930 329.140 ;
        RECT 141.870 329.120 142.240 329.140 ;
        RECT 49.620 326.520 127.730 328.600 ;
        RECT 130.980 328.320 140.930 328.700 ;
        RECT 130.980 327.520 132.250 328.320 ;
        RECT 143.830 327.510 144.180 329.800 ;
        RECT 147.460 329.770 147.770 329.900 ;
        RECT 144.800 329.460 147.960 329.600 ;
        RECT 144.690 329.280 147.960 329.460 ;
        RECT 144.690 329.130 145.000 329.280 ;
        RECT 145.790 329.130 146.100 329.280 ;
        RECT 146.890 329.130 147.200 329.280 ;
        RECT 147.640 328.820 147.960 329.280 ;
        RECT 150.540 328.820 150.820 328.830 ;
        RECT 146.950 328.490 150.840 328.820 ;
        RECT 176.560 328.800 176.880 331.250 ;
        RECT 177.880 330.870 178.190 331.050 ;
        RECT 178.970 330.870 179.280 331.030 ;
        RECT 180.080 330.870 180.390 331.020 ;
        RECT 182.810 330.870 183.120 331.020 ;
        RECT 183.920 330.870 184.230 331.030 ;
        RECT 185.010 330.870 185.320 331.050 ;
        RECT 177.750 330.570 180.690 330.870 ;
        RECT 179.940 330.530 180.690 330.570 ;
        RECT 180.310 330.400 180.690 330.530 ;
        RECT 180.340 329.680 180.690 330.400 ;
        RECT 182.510 330.570 185.450 330.870 ;
        RECT 182.510 330.530 183.260 330.570 ;
        RECT 182.510 330.400 182.890 330.530 ;
        RECT 182.510 329.970 182.860 330.400 ;
        RECT 186.320 329.970 186.690 331.250 ;
        RECT 187.690 330.900 188.000 331.080 ;
        RECT 188.780 330.900 189.090 331.060 ;
        RECT 189.890 330.900 190.200 331.050 ;
        RECT 192.620 330.900 192.930 331.050 ;
        RECT 193.730 330.900 194.040 331.060 ;
        RECT 194.820 330.900 195.130 331.080 ;
        RECT 187.560 330.600 190.500 330.900 ;
        RECT 189.750 330.560 190.500 330.600 ;
        RECT 190.120 330.430 190.500 330.560 ;
        RECT 190.150 329.970 190.500 330.430 ;
        RECT 192.320 330.600 195.260 330.900 ;
        RECT 192.320 330.560 193.070 330.600 ;
        RECT 192.320 330.430 192.700 330.560 ;
        RECT 181.070 329.940 191.970 329.970 ;
        RECT 177.880 329.530 178.190 329.680 ;
        RECT 178.970 329.530 179.280 329.680 ;
        RECT 180.070 329.530 180.690 329.680 ;
        RECT 181.060 329.690 191.970 329.940 ;
        RECT 192.320 329.710 192.670 330.430 ;
        RECT 181.060 329.660 181.400 329.690 ;
        RECT 181.800 329.680 182.140 329.690 ;
        RECT 182.510 329.680 182.860 329.690 ;
        RECT 177.740 329.200 180.690 329.530 ;
        RECT 177.140 329.150 177.640 329.160 ;
        RECT 180.340 329.150 180.690 329.200 ;
        RECT 182.510 329.530 183.130 329.680 ;
        RECT 183.920 329.530 184.230 329.680 ;
        RECT 185.010 329.530 185.320 329.680 ;
        RECT 182.510 329.200 185.460 329.530 ;
        RECT 182.510 329.150 182.860 329.200 ;
        RECT 186.320 329.150 186.690 329.690 ;
        RECT 187.690 329.560 188.000 329.690 ;
        RECT 188.780 329.560 189.090 329.690 ;
        RECT 189.880 329.560 190.500 329.690 ;
        RECT 190.870 329.660 191.210 329.690 ;
        RECT 187.550 329.230 190.500 329.560 ;
        RECT 190.150 329.150 190.500 329.230 ;
        RECT 192.320 329.560 192.940 329.710 ;
        RECT 193.730 329.560 194.040 329.710 ;
        RECT 194.820 329.560 195.130 329.710 ;
        RECT 192.320 329.230 195.270 329.560 ;
        RECT 192.320 329.150 192.670 329.230 ;
        RECT 196.130 329.150 196.450 331.280 ;
        RECT 199.040 331.260 202.190 331.400 ;
        RECT 198.360 330.880 198.670 331.030 ;
        RECT 199.470 330.880 199.780 331.040 ;
        RECT 200.560 330.880 200.870 331.060 ;
        RECT 198.060 330.580 201.000 330.880 ;
        RECT 198.060 330.540 198.810 330.580 ;
        RECT 198.060 330.410 198.440 330.540 ;
        RECT 198.060 329.690 198.410 330.410 ;
        RECT 198.060 329.540 198.680 329.690 ;
        RECT 199.470 329.540 199.780 329.690 ;
        RECT 200.560 329.540 200.870 329.690 ;
        RECT 198.060 329.210 201.010 329.540 ;
        RECT 198.060 329.150 198.410 329.210 ;
        RECT 201.870 329.150 202.190 331.260 ;
        RECT 223.070 329.150 223.630 329.170 ;
        RECT 177.140 328.800 223.630 329.150 ;
        RECT 176.560 328.690 223.630 328.800 ;
        RECT 176.560 328.620 179.830 328.690 ;
        RECT 147.640 328.240 147.960 328.490 ;
        RECT 150.540 328.470 150.820 328.490 ;
        RECT 176.560 328.470 179.720 328.620 ;
        RECT 144.800 328.090 147.960 328.240 ;
        RECT 144.690 327.910 147.960 328.090 ;
        RECT 144.690 327.760 145.000 327.910 ;
        RECT 145.790 327.760 146.100 327.910 ;
        RECT 146.890 327.760 147.200 327.910 ;
        RECT 143.830 327.180 146.780 327.510 ;
        RECT 143.120 327.140 143.470 327.170 ;
        RECT 143.830 327.140 144.450 327.180 ;
        RECT 145.240 327.140 145.550 327.180 ;
        RECT 146.330 327.140 146.640 327.180 ;
        RECT 147.640 327.140 147.960 327.910 ;
        RECT 176.560 327.430 176.880 328.470 ;
        RECT 177.320 327.430 177.630 327.580 ;
        RECT 178.420 327.430 178.730 327.580 ;
        RECT 179.520 327.430 179.830 327.580 ;
        RECT 176.560 327.250 179.830 327.430 ;
        RECT 149.500 327.160 149.830 327.200 ;
        RECT 149.490 327.140 149.840 327.160 ;
        RECT 143.120 326.880 153.150 327.140 ;
        RECT 176.560 327.110 179.720 327.250 ;
        RECT 143.160 326.850 153.150 326.880 ;
        RECT 45.210 186.740 47.810 190.470 ;
        RECT 45.460 186.410 47.540 186.740 ;
        RECT 49.620 161.840 51.700 326.520 ;
        RECT 143.830 326.310 144.180 326.850 ;
        RECT 147.640 326.510 147.960 326.850 ;
        RECT 149.500 326.830 149.830 326.850 ;
        RECT 143.830 326.180 144.210 326.310 ;
        RECT 143.830 326.140 144.580 326.180 ;
        RECT 146.960 326.170 149.300 326.510 ;
        RECT 143.830 325.840 146.770 326.140 ;
        RECT 146.960 325.930 149.340 326.170 ;
        RECT 146.960 325.910 149.300 325.930 ;
        RECT 144.130 325.690 144.440 325.840 ;
        RECT 145.240 325.680 145.550 325.840 ;
        RECT 146.330 325.660 146.640 325.840 ;
        RECT 98.440 325.590 99.040 325.640 ;
        RECT 98.440 325.150 127.780 325.590 ;
        RECT 147.640 325.460 147.960 325.910 ;
        RECT 148.330 325.840 148.990 325.910 ;
        RECT 148.360 325.830 148.960 325.840 ;
        RECT 144.810 325.320 147.960 325.460 ;
        RECT 98.440 325.080 99.040 325.150 ;
        RECT 144.690 325.130 147.960 325.320 ;
        RECT 144.690 325.120 147.870 325.130 ;
        RECT 144.690 324.990 145.000 325.120 ;
        RECT 145.790 324.980 146.100 325.120 ;
        RECT 146.880 324.980 147.190 325.120 ;
        RECT 152.850 324.770 153.140 326.850 ;
        RECT 176.750 326.810 177.060 326.940 ;
        RECT 180.340 326.910 180.690 328.690 ;
        RECT 176.320 326.610 177.060 326.810 ;
        RECT 177.880 326.760 178.190 326.900 ;
        RECT 178.970 326.760 179.280 326.900 ;
        RECT 180.070 326.760 180.690 326.910 ;
        RECT 176.320 326.470 176.920 326.610 ;
        RECT 176.320 326.140 177.070 326.470 ;
        RECT 177.750 326.440 180.690 326.760 ;
        RECT 182.510 326.910 182.860 328.690 ;
        RECT 183.370 328.650 189.640 328.690 ;
        RECT 183.370 328.620 189.530 328.650 ;
        RECT 183.480 328.500 189.530 328.620 ;
        RECT 183.480 328.470 186.690 328.500 ;
        RECT 186.320 328.240 186.690 328.470 ;
        RECT 190.150 328.240 190.500 328.690 ;
        RECT 192.320 328.240 192.670 328.690 ;
        RECT 193.180 328.650 196.450 328.690 ;
        RECT 193.290 328.500 196.450 328.650 ;
        RECT 196.130 328.240 196.450 328.500 ;
        RECT 198.060 328.240 198.410 328.690 ;
        RECT 198.920 328.630 202.190 328.690 ;
        RECT 223.070 328.670 223.630 328.690 ;
        RECT 199.030 328.480 202.190 328.630 ;
        RECT 201.870 328.240 202.190 328.480 ;
        RECT 185.450 327.780 222.530 328.240 ;
        RECT 185.520 327.680 186.040 327.780 ;
        RECT 183.370 327.430 183.680 327.580 ;
        RECT 184.470 327.430 184.780 327.580 ;
        RECT 185.570 327.430 185.880 327.580 ;
        RECT 186.320 327.460 186.690 327.780 ;
        RECT 187.130 327.460 187.440 327.610 ;
        RECT 188.230 327.460 188.540 327.610 ;
        RECT 189.330 327.460 189.640 327.610 ;
        RECT 186.320 327.430 189.640 327.460 ;
        RECT 183.370 327.330 189.640 327.430 ;
        RECT 190.150 327.330 190.500 327.780 ;
        RECT 192.320 327.330 192.670 327.780 ;
        RECT 193.180 327.460 193.490 327.610 ;
        RECT 194.280 327.460 194.590 327.610 ;
        RECT 195.380 327.460 195.690 327.610 ;
        RECT 196.130 327.460 196.450 327.780 ;
        RECT 193.180 327.330 196.450 327.460 ;
        RECT 198.060 327.330 198.410 327.780 ;
        RECT 198.920 327.440 199.230 327.590 ;
        RECT 200.020 327.440 200.330 327.590 ;
        RECT 201.120 327.440 201.430 327.590 ;
        RECT 201.870 327.440 202.190 327.780 ;
        RECT 221.880 327.720 222.440 327.780 ;
        RECT 198.920 327.330 202.190 327.440 ;
        RECT 183.370 327.250 221.440 327.330 ;
        RECT 183.480 327.140 221.440 327.250 ;
        RECT 183.480 327.110 186.640 327.140 ;
        RECT 182.510 326.760 183.130 326.910 ;
        RECT 183.920 326.760 184.230 326.900 ;
        RECT 185.010 326.760 185.320 326.900 ;
        RECT 186.140 326.840 186.450 326.940 ;
        RECT 186.560 326.840 186.870 326.970 ;
        RECT 186.130 326.810 186.870 326.840 ;
        RECT 186.880 326.870 221.440 327.140 ;
        RECT 186.880 326.810 187.530 326.870 ;
        RECT 182.510 326.440 185.450 326.760 ;
        RECT 177.750 326.430 180.460 326.440 ;
        RECT 182.740 326.430 185.450 326.440 ;
        RECT 186.130 326.740 187.530 326.810 ;
        RECT 187.690 326.790 188.000 326.870 ;
        RECT 188.780 326.790 189.090 326.870 ;
        RECT 189.880 326.790 190.500 326.870 ;
        RECT 176.320 325.990 176.920 326.140 ;
        RECT 186.130 326.020 186.880 326.740 ;
        RECT 187.560 326.470 190.500 326.790 ;
        RECT 192.320 326.790 192.940 326.870 ;
        RECT 193.730 326.790 194.040 326.870 ;
        RECT 194.820 326.790 195.130 326.870 ;
        RECT 195.950 326.840 196.260 326.870 ;
        RECT 192.320 326.470 195.260 326.790 ;
        RECT 195.950 326.640 196.690 326.840 ;
        RECT 196.090 326.500 196.690 326.640 ;
        RECT 187.560 326.460 190.270 326.470 ;
        RECT 192.550 326.460 195.260 326.470 ;
        RECT 186.280 325.990 186.880 326.020 ;
        RECT 195.330 326.390 195.850 326.410 ;
        RECT 195.940 326.390 196.690 326.500 ;
        RECT 198.060 326.770 198.680 326.870 ;
        RECT 199.470 326.770 199.780 326.870 ;
        RECT 200.560 326.770 200.870 326.870 ;
        RECT 201.690 326.820 202.000 326.870 ;
        RECT 220.750 326.850 221.310 326.870 ;
        RECT 198.060 326.450 201.000 326.770 ;
        RECT 201.690 326.620 202.430 326.820 ;
        RECT 201.830 326.480 202.430 326.620 ;
        RECT 198.290 326.440 201.000 326.450 ;
        RECT 201.680 326.390 202.430 326.480 ;
        RECT 219.820 326.390 220.380 326.400 ;
        RECT 195.330 325.930 220.470 326.390 ;
        RECT 195.330 325.880 195.860 325.930 ;
        RECT 195.330 325.830 195.850 325.880 ;
        RECT 169.270 324.770 169.590 324.790 ;
        RECT 225.270 324.770 226.430 324.800 ;
        RECT 101.870 324.610 102.330 324.620 ;
        RECT 101.870 324.170 127.740 324.610 ;
        RECT 101.870 324.150 102.330 324.170 ;
        RECT 130.980 323.470 132.250 324.380 ;
        RECT 152.660 323.650 226.430 324.770 ;
        RECT 169.270 323.630 169.590 323.650 ;
        RECT 180.640 323.570 182.560 323.650 ;
        RECT 190.450 323.540 192.380 323.650 ;
        RECT 225.270 323.620 226.430 323.650 ;
        RECT 53.870 321.370 127.730 323.450 ;
        RECT 130.980 323.090 140.950 323.470 ;
        RECT 232.850 323.250 233.180 323.560 ;
        RECT 130.980 322.500 132.250 323.090 ;
        RECT 140.570 322.240 140.950 323.090 ;
        RECT 232.870 323.070 233.160 323.250 ;
        RECT 232.880 322.890 233.160 323.070 ;
        RECT 232.850 322.580 233.180 322.890 ;
        RECT 232.880 322.320 233.160 322.580 ;
        RECT 141.870 322.240 142.240 322.250 ;
        RECT 140.570 321.860 143.290 322.240 ;
        RECT 141.870 321.840 142.240 321.860 ;
        RECT 229.100 321.470 229.300 321.480 ;
        RECT 49.200 158.170 51.910 161.840 ;
        RECT 49.620 157.450 51.700 158.170 ;
        RECT 53.870 133.220 55.950 321.370 ;
        RECT 229.100 321.320 233.040 321.470 ;
        RECT 151.120 321.270 151.430 321.290 ;
        RECT 146.890 320.930 151.430 321.270 ;
        RECT 151.120 320.910 151.430 320.930 ;
        RECT 132.190 320.320 132.690 320.430 ;
        RECT 201.160 320.350 201.550 320.360 ;
        RECT 201.150 320.320 201.550 320.350 ;
        RECT 132.190 320.040 201.550 320.320 ;
        RECT 132.190 319.960 132.690 320.040 ;
        RECT 201.150 320.020 201.550 320.040 ;
        RECT 201.160 320.010 201.550 320.020 ;
        RECT 167.570 319.690 167.990 319.700 ;
        RECT 167.570 319.440 207.840 319.690 ;
        RECT 167.570 319.360 207.850 319.440 ;
        RECT 167.570 319.350 167.990 319.360 ;
        RECT 201.810 319.340 207.850 319.360 ;
        RECT 58.130 317.110 127.730 319.190 ;
        RECT 166.970 319.070 167.350 319.080 ;
        RECT 53.540 129.740 56.280 133.220 ;
        RECT 53.870 128.930 55.950 129.740 ;
        RECT 58.130 104.930 60.210 317.110 ;
        RECT 130.850 316.960 132.120 318.840 ;
        RECT 166.970 318.740 203.770 319.070 ;
        RECT 166.970 318.730 167.350 318.740 ;
        RECT 197.700 318.730 203.770 318.740 ;
        RECT 166.330 318.440 166.750 318.450 ;
        RECT 166.330 318.110 199.690 318.440 ;
        RECT 166.330 318.100 166.750 318.110 ;
        RECT 165.740 317.800 166.140 317.820 ;
        RECT 165.740 317.470 195.680 317.800 ;
        RECT 165.740 317.460 166.140 317.470 ;
        RECT 165.080 317.130 165.490 317.140 ;
        RECT 165.070 316.800 191.590 317.130 ;
        RECT 165.080 316.780 165.490 316.800 ;
        RECT 164.500 316.510 164.910 316.520 ;
        RECT 164.500 316.490 187.570 316.510 ;
        RECT 164.500 316.180 187.580 316.490 ;
        RECT 164.500 316.170 164.910 316.180 ;
        RECT 163.900 315.860 164.290 315.870 ;
        RECT 163.900 315.540 183.590 315.860 ;
        RECT 164.000 315.530 183.590 315.540 ;
        RECT 163.320 315.250 163.710 315.300 ;
        RECT 158.180 315.040 158.720 315.080 ;
        RECT 145.350 315.000 158.720 315.040 ;
        RECT 145.300 314.610 158.720 315.000 ;
        RECT 163.320 314.970 179.680 315.250 ;
        RECT 163.580 314.920 179.680 314.970 ;
        RECT 62.280 312.070 127.730 314.150 ;
        RECT 130.920 312.210 132.190 314.090 ;
        RECT 145.300 312.730 147.310 314.610 ;
        RECT 158.180 314.580 158.720 314.610 ;
        RECT 162.740 314.280 175.480 314.610 ;
        RECT 158.830 314.200 159.370 314.270 ;
        RECT 149.400 313.770 159.370 314.200 ;
        RECT 169.350 313.980 171.370 314.000 ;
        RECT 162.190 313.970 171.400 313.980 ;
        RECT 149.400 312.760 151.380 313.770 ;
        RECT 162.090 313.650 171.400 313.970 ;
        RECT 162.090 313.640 162.480 313.650 ;
        RECT 159.510 313.390 160.000 313.590 ;
        RECT 153.900 313.370 160.000 313.390 ;
        RECT 153.330 313.090 160.000 313.370 ;
        RECT 153.330 312.990 159.910 313.090 ;
        RECT 161.450 312.990 167.430 313.330 ;
        RECT 153.330 312.760 155.310 312.990 ;
        RECT 159.340 312.760 159.990 312.770 ;
        RECT 145.280 312.070 147.310 312.730 ;
        RECT 149.350 312.100 151.380 312.760 ;
        RECT 153.310 312.100 155.340 312.760 ;
        RECT 157.310 312.130 159.990 312.760 ;
        RECT 160.840 312.740 161.390 312.760 ;
        RECT 160.840 312.310 163.390 312.740 ;
        RECT 165.400 312.730 167.440 312.990 ;
        RECT 157.310 312.100 159.340 312.130 ;
        RECT 161.360 312.080 163.390 312.310 ;
        RECT 165.390 312.070 167.440 312.730 ;
        RECT 169.320 312.100 171.400 313.650 ;
        RECT 173.430 312.980 175.460 314.280 ;
        RECT 173.430 312.690 175.470 312.980 ;
        RECT 173.440 312.080 175.470 312.690 ;
        RECT 177.610 312.100 179.640 314.920 ;
        RECT 181.600 312.820 183.590 315.530 ;
        RECT 181.590 312.070 183.620 312.820 ;
        RECT 185.580 312.800 187.580 316.180 ;
        RECT 185.550 312.100 187.580 312.800 ;
        RECT 189.680 312.730 191.590 316.800 ;
        RECT 193.720 312.750 195.670 317.470 ;
        RECT 197.700 312.750 199.690 318.110 ;
        RECT 201.810 318.410 203.770 318.730 ;
        RECT 205.910 318.840 207.850 319.340 ;
        RECT 228.430 319.230 228.860 319.250 ;
        RECT 209.930 319.200 211.890 319.230 ;
        RECT 228.410 319.200 228.870 319.230 ;
        RECT 209.930 318.850 228.870 319.200 ;
        RECT 201.810 312.750 203.760 318.410 ;
        RECT 205.910 312.770 207.840 318.840 ;
        RECT 189.600 312.080 191.630 312.730 ;
        RECT 193.670 312.100 195.700 312.750 ;
        RECT 197.700 312.100 199.730 312.750 ;
        RECT 201.750 312.100 203.780 312.750 ;
        RECT 57.910 100.880 60.700 104.930 ;
        RECT 58.130 100.600 60.210 100.880 ;
        RECT 62.280 76.150 64.360 312.070 ;
        RECT 205.820 311.990 207.850 312.770 ;
        RECT 209.930 312.750 211.890 318.850 ;
        RECT 228.410 318.830 228.870 318.850 ;
        RECT 228.430 318.820 228.860 318.830 ;
        RECT 229.100 318.410 229.300 321.320 ;
        RECT 233.120 321.290 233.440 321.610 ;
        RECT 230.070 319.720 232.880 319.920 ;
        RECT 229.330 318.420 229.760 318.440 ;
        RECT 229.320 318.410 229.770 318.420 ;
        RECT 213.860 318.030 229.770 318.410 ;
        RECT 209.900 312.100 211.930 312.750 ;
        RECT 213.860 312.730 215.820 318.030 ;
        RECT 227.980 317.960 228.310 318.030 ;
        RECT 227.980 317.590 228.180 317.960 ;
        RECT 229.100 317.590 229.300 318.030 ;
        RECT 229.330 318.010 229.760 318.030 ;
        RECT 230.070 317.600 230.280 319.720 ;
        RECT 233.120 319.680 233.440 320.000 ;
        RECT 231.850 318.260 232.160 318.290 ;
        RECT 231.850 318.010 232.920 318.260 ;
        RECT 233.110 318.070 233.430 318.390 ;
        RECT 230.070 317.590 230.700 317.600 ;
        RECT 218.010 317.210 230.700 317.590 ;
        RECT 218.010 312.750 219.990 317.210 ;
        RECT 227.980 316.800 228.180 317.210 ;
        RECT 229.100 316.800 229.300 317.210 ;
        RECT 230.070 316.800 230.280 317.210 ;
        RECT 231.090 316.800 231.510 316.830 ;
        RECT 222.120 316.420 231.510 316.800 ;
        RECT 213.850 312.080 215.880 312.730 ;
        RECT 217.970 312.100 220.000 312.750 ;
        RECT 222.120 312.720 224.100 316.420 ;
        RECT 227.980 313.630 228.180 316.420 ;
        RECT 229.100 313.630 229.300 316.420 ;
        RECT 230.070 313.630 230.280 316.420 ;
        RECT 231.090 316.390 231.510 316.420 ;
        RECT 231.850 313.630 232.150 318.010 ;
        RECT 233.120 316.660 233.440 316.770 ;
        RECT 232.970 316.450 233.440 316.660 ;
        RECT 232.970 315.160 233.160 316.450 ;
        RECT 232.970 314.840 233.430 315.160 ;
        RECT 232.350 313.630 232.670 313.680 ;
        RECT 232.970 313.630 233.160 314.840 ;
        RECT 227.190 313.430 233.430 313.630 ;
        RECT 227.190 312.750 227.390 313.430 ;
        RECT 227.980 312.750 228.180 313.430 ;
        RECT 222.110 312.070 224.140 312.720 ;
        RECT 226.100 312.100 228.180 312.750 ;
        RECT 227.980 309.610 228.180 312.100 ;
        RECT 229.100 309.750 229.300 313.430 ;
        RECT 230.070 312.750 230.280 313.430 ;
        RECT 231.850 313.310 232.150 313.430 ;
        RECT 232.350 313.360 232.670 313.430 ;
        RECT 231.850 313.220 232.610 313.310 ;
        RECT 232.970 313.220 233.160 313.430 ;
        RECT 234.350 313.220 234.550 313.630 ;
        RECT 231.850 313.020 234.550 313.220 ;
        RECT 231.850 312.750 232.320 313.020 ;
        RECT 230.070 312.450 232.320 312.750 ;
        RECT 230.070 312.100 232.150 312.450 ;
        RECT 230.070 310.250 230.280 312.100 ;
        RECT 231.850 311.670 232.150 312.100 ;
        RECT 232.970 311.960 233.160 313.020 ;
        RECT 235.320 312.750 235.530 313.640 ;
        RECT 234.200 312.100 236.230 312.750 ;
        RECT 237.250 312.660 237.460 313.640 ;
        RECT 238.220 313.450 238.410 313.620 ;
        RECT 238.220 313.260 243.220 313.450 ;
        RECT 243.030 312.800 243.220 313.260 ;
        RECT 238.380 312.660 240.410 312.750 ;
        RECT 243.030 312.730 244.060 312.800 ;
        RECT 237.250 312.450 240.410 312.660 ;
        RECT 238.380 312.100 240.410 312.450 ;
        RECT 242.360 312.080 244.390 312.730 ;
        RECT 231.850 311.510 232.210 311.670 ;
        RECT 229.870 309.930 230.280 310.250 ;
        RECT 230.810 309.930 231.130 310.250 ;
        RECT 232.000 310.230 232.210 311.510 ;
        RECT 229.090 309.610 229.300 309.750 ;
        RECT 230.070 309.610 230.280 309.930 ;
        RECT 231.760 309.870 232.210 310.230 ;
        RECT 232.970 311.640 233.430 311.960 ;
        RECT 232.970 310.250 233.160 311.640 ;
        RECT 232.970 309.930 233.390 310.250 ;
        RECT 232.970 309.900 233.160 309.930 ;
        RECT 232.000 309.610 232.210 309.870 ;
        RECT 232.950 309.610 233.160 309.900 ;
        RECT 66.630 306.460 127.730 308.540 ;
        RECT 61.790 72.370 64.620 76.150 ;
        RECT 62.280 71.810 64.360 72.370 ;
        RECT 66.630 47.570 68.710 306.460 ;
        RECT 70.790 301.760 127.730 303.840 ;
        RECT 66.280 43.850 68.930 47.570 ;
        RECT 66.630 43.840 68.710 43.850 ;
        RECT 70.790 18.870 72.870 301.760 ;
        RECT 70.600 15.340 73.270 18.870 ;
        RECT 132.330 9.510 135.670 301.900 ;
        RECT 335.350 246.810 337.440 333.840 ;
        RECT 339.440 275.580 341.530 339.040 ;
        RECT 343.520 304.080 345.610 343.920 ;
        RECT 347.660 332.640 349.750 349.320 ;
        RECT 347.460 329.100 349.890 332.640 ;
        RECT 347.660 328.430 349.750 329.100 ;
        RECT 343.280 300.510 345.790 304.080 ;
        RECT 383.930 285.540 385.330 286.060 ;
        RECT 383.800 285.460 385.330 285.540 ;
        RECT 383.290 284.450 385.330 285.460 ;
        RECT 383.290 283.810 388.340 284.450 ;
        RECT 383.290 283.530 385.330 283.810 ;
        RECT 383.220 282.910 385.330 283.530 ;
        RECT 339.240 271.870 341.760 275.580 ;
        RECT 339.440 271.840 341.530 271.870 ;
        RECT 383.930 256.950 385.330 282.910 ;
        RECT 390.230 258.870 391.630 286.060 ;
        RECT 390.220 258.360 391.630 258.870 ;
        RECT 389.110 258.190 391.630 258.360 ;
        RECT 390.220 257.940 391.630 258.190 ;
        RECT 383.800 256.870 385.330 256.950 ;
        RECT 383.290 255.860 385.330 256.870 ;
        RECT 383.290 255.220 388.340 255.860 ;
        RECT 383.290 254.940 385.330 255.220 ;
        RECT 383.220 254.320 385.330 254.940 ;
        RECT 335.080 243.390 337.440 246.810 ;
        RECT 335.350 242.680 337.440 243.390 ;
        RECT 383.930 228.360 385.330 254.320 ;
        RECT 390.230 230.280 391.630 257.940 ;
        RECT 390.220 229.770 391.630 230.280 ;
        RECT 389.110 229.600 391.630 229.770 ;
        RECT 390.220 229.350 391.630 229.600 ;
        RECT 383.800 228.280 385.330 228.360 ;
        RECT 383.290 227.270 385.330 228.280 ;
        RECT 383.290 226.630 388.340 227.270 ;
        RECT 383.290 226.350 385.330 226.630 ;
        RECT 383.220 225.730 385.330 226.350 ;
        RECT 383.930 199.770 385.330 225.730 ;
        RECT 390.230 201.690 391.630 229.350 ;
        RECT 390.220 201.180 391.630 201.690 ;
        RECT 389.110 201.010 391.630 201.180 ;
        RECT 390.220 200.760 391.630 201.010 ;
        RECT 383.800 199.690 385.330 199.770 ;
        RECT 383.290 198.680 385.330 199.690 ;
        RECT 383.290 198.040 388.340 198.680 ;
        RECT 383.290 197.760 385.330 198.040 ;
        RECT 383.220 197.140 385.330 197.760 ;
        RECT 383.930 171.180 385.330 197.140 ;
        RECT 390.230 173.100 391.630 200.760 ;
        RECT 390.220 172.590 391.630 173.100 ;
        RECT 389.110 172.420 391.630 172.590 ;
        RECT 390.220 172.170 391.630 172.420 ;
        RECT 383.800 171.100 385.330 171.180 ;
        RECT 383.290 170.090 385.330 171.100 ;
        RECT 383.290 169.450 388.340 170.090 ;
        RECT 383.290 169.170 385.330 169.450 ;
        RECT 383.220 168.550 385.330 169.170 ;
        RECT 383.930 142.590 385.330 168.550 ;
        RECT 390.230 144.510 391.630 172.170 ;
        RECT 390.220 144.000 391.630 144.510 ;
        RECT 389.110 143.830 391.630 144.000 ;
        RECT 390.220 143.580 391.630 143.830 ;
        RECT 383.800 142.510 385.330 142.590 ;
        RECT 383.290 141.500 385.330 142.510 ;
        RECT 383.290 140.860 388.340 141.500 ;
        RECT 383.290 140.580 385.330 140.860 ;
        RECT 383.220 139.960 385.330 140.580 ;
        RECT 383.930 114.000 385.330 139.960 ;
        RECT 390.230 115.920 391.630 143.580 ;
        RECT 390.220 115.410 391.630 115.920 ;
        RECT 389.110 115.240 391.630 115.410 ;
        RECT 390.220 114.990 391.630 115.240 ;
        RECT 383.800 113.920 385.330 114.000 ;
        RECT 383.290 112.910 385.330 113.920 ;
        RECT 383.290 112.270 388.340 112.910 ;
        RECT 383.290 111.990 385.330 112.270 ;
        RECT 383.220 111.370 385.330 111.990 ;
        RECT 383.930 85.930 385.330 111.370 ;
        RECT 390.230 87.330 391.630 114.990 ;
        RECT 390.220 86.820 391.630 87.330 ;
        RECT 389.110 86.650 391.630 86.820 ;
        RECT 390.220 86.400 391.630 86.650 ;
        RECT 390.230 85.930 391.630 86.400 ;
      LAYER via2 ;
        RECT 207.560 367.230 207.880 367.550 ;
        RECT 208.590 367.220 208.910 367.540 ;
        RECT 208.670 363.740 209.010 364.080 ;
        RECT 207.600 360.260 207.930 360.610 ;
        RECT 208.690 357.690 209.030 358.050 ;
      LAYER met3 ;
        RECT 207.490 366.860 207.940 367.610 ;
        RECT 207.490 360.700 207.860 366.860 ;
        RECT 208.530 366.850 208.980 367.600 ;
        RECT 208.610 364.210 208.980 366.850 ;
        RECT 208.610 363.610 209.050 364.210 ;
        RECT 207.490 360.370 207.980 360.700 ;
        RECT 207.540 360.210 207.980 360.370 ;
        RECT 208.610 358.500 208.980 363.610 ;
        RECT 208.600 357.630 209.070 358.500 ;
  END
END sky130_hilas_TopProtectStructure

MACRO sky130_hilas_nFETLarge
  CLASS CORE ;
  FOREIGN sky130_hilas_nFETLarge ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.570 BY 6.030 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    USE ANALOG ;
    ANTENNAGATEAREA 2.642500 ;
    PORT
      LAYER met2 ;
        RECT 0.430 0.820 0.740 0.950 ;
        RECT 0.000 0.620 0.740 0.820 ;
        RECT 0.000 0.480 0.600 0.620 ;
        RECT 0.000 0.150 0.750 0.480 ;
        RECT 0.000 0.000 0.600 0.150 ;
    END
  END GATE
  PIN SOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 1.343400 ;
    PORT
      LAYER met2 ;
        RECT 1.010 5.600 1.320 5.740 ;
        RECT 2.100 5.600 2.410 5.740 ;
        RECT 3.200 5.600 3.510 5.730 ;
        RECT 0.330 5.590 3.510 5.600 ;
        RECT 0.240 5.400 3.510 5.590 ;
        RECT 0.240 5.260 3.390 5.400 ;
        RECT 0.240 2.810 0.560 5.260 ;
        RECT 1.000 2.810 1.310 2.960 ;
        RECT 2.100 2.810 2.410 2.960 ;
        RECT 3.200 2.810 3.510 2.960 ;
        RECT 0.240 2.630 3.510 2.810 ;
        RECT 0.240 2.480 3.400 2.630 ;
        RECT 0.240 1.440 0.560 2.480 ;
        RECT 1.000 1.440 1.310 1.590 ;
        RECT 2.100 1.440 2.410 1.590 ;
        RECT 3.200 1.440 3.510 1.590 ;
        RECT 0.240 1.260 3.510 1.440 ;
        RECT 0.240 1.120 3.400 1.260 ;
    END
  END SOURCE
  PIN DRAIN
    USE ANALOG ;
    ANTENNADIFFAREA 2.723900 ;
    PORT
      LAYER met2 ;
        RECT 1.560 4.880 1.870 5.060 ;
        RECT 2.650 4.880 2.960 5.040 ;
        RECT 3.760 4.880 4.070 5.030 ;
        RECT 1.430 4.580 4.370 4.880 ;
        RECT 3.620 4.540 4.370 4.580 ;
        RECT 3.990 4.410 4.370 4.540 ;
        RECT 4.020 3.690 4.370 4.410 ;
        RECT 1.560 3.540 1.870 3.690 ;
        RECT 2.650 3.540 2.960 3.690 ;
        RECT 3.750 3.540 4.370 3.690 ;
        RECT 1.420 3.210 4.370 3.540 ;
        RECT 4.020 0.920 4.370 3.210 ;
        RECT 1.560 0.770 1.870 0.910 ;
        RECT 2.650 0.770 2.960 0.910 ;
        RECT 3.750 0.770 4.370 0.920 ;
        RECT 1.430 0.450 4.370 0.770 ;
        RECT 1.430 0.440 4.140 0.450 ;
    END
  END DRAIN
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.180 2.450 0.450 2.480 ;
        RECT 0.180 1.920 0.460 2.450 ;
        RECT 0.000 1.620 0.460 1.920 ;
        RECT 0.000 1.600 0.470 1.620 ;
        RECT 0.180 1.170 0.470 1.600 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.020 5.660 1.340 5.700 ;
        RECT 2.110 5.660 2.430 5.700 ;
        RECT 1.020 5.470 1.350 5.660 ;
        RECT 2.110 5.470 2.440 5.660 ;
        RECT 1.020 5.440 1.340 5.470 ;
        RECT 2.110 5.440 2.430 5.470 ;
        RECT 1.570 4.980 1.890 5.020 ;
        RECT 2.600 5.000 2.770 5.890 ;
        RECT 3.150 5.690 3.320 5.890 ;
        RECT 3.150 5.650 3.530 5.690 ;
        RECT 3.150 5.460 3.540 5.650 ;
        RECT 3.150 5.430 3.530 5.460 ;
        RECT 1.570 4.790 1.900 4.980 ;
        RECT 2.600 4.960 2.980 5.000 ;
        RECT 1.570 4.760 1.890 4.790 ;
        RECT 2.600 4.770 2.990 4.960 ;
        RECT 2.600 4.740 2.980 4.770 ;
        RECT 2.600 3.650 2.770 4.740 ;
        RECT 1.570 3.610 1.890 3.650 ;
        RECT 2.600 3.610 2.980 3.650 ;
        RECT 1.570 3.420 1.900 3.610 ;
        RECT 2.600 3.490 2.990 3.610 ;
        RECT 3.150 3.490 3.320 5.430 ;
        RECT 3.700 4.990 3.870 5.890 ;
        RECT 3.700 4.950 4.090 4.990 ;
        RECT 3.700 4.760 4.100 4.950 ;
        RECT 3.700 4.730 4.090 4.760 ;
        RECT 3.700 3.650 3.870 4.730 ;
        RECT 3.700 3.610 4.080 3.650 ;
        RECT 3.700 3.490 4.090 3.610 ;
        RECT 4.250 3.490 4.420 5.890 ;
        RECT 4.800 3.490 4.970 5.890 ;
        RECT 5.350 3.490 5.520 5.890 ;
        RECT 2.660 3.420 2.990 3.490 ;
        RECT 3.760 3.420 4.090 3.490 ;
        RECT 1.570 3.390 1.890 3.420 ;
        RECT 2.660 3.390 2.980 3.420 ;
        RECT 3.760 3.390 4.080 3.420 ;
        RECT 0.950 2.920 1.120 3.180 ;
        RECT 0.950 2.880 1.330 2.920 ;
        RECT 0.950 2.800 1.340 2.880 ;
        RECT 1.500 2.800 1.670 3.180 ;
        RECT 2.050 2.920 2.220 3.180 ;
        RECT 2.050 2.880 2.430 2.920 ;
        RECT 2.050 2.800 2.440 2.880 ;
        RECT 1.010 2.690 1.340 2.800 ;
        RECT 2.110 2.690 2.440 2.800 ;
        RECT 1.010 2.660 1.330 2.690 ;
        RECT 2.110 2.660 2.430 2.690 ;
        RECT 0.240 1.200 0.410 2.420 ;
        RECT 1.010 1.510 1.330 1.550 ;
        RECT 2.110 1.510 2.430 1.550 ;
        RECT 1.010 1.320 1.340 1.510 ;
        RECT 2.110 1.320 2.440 1.510 ;
        RECT 1.010 1.290 1.330 1.320 ;
        RECT 2.110 1.290 2.430 1.320 ;
        RECT 0.190 0.910 0.700 1.010 ;
        RECT 0.190 0.870 0.760 0.910 ;
        RECT 2.600 0.870 2.770 3.180 ;
        RECT 3.150 2.920 3.320 3.180 ;
        RECT 3.150 2.880 3.530 2.920 ;
        RECT 3.150 2.690 3.540 2.880 ;
        RECT 3.150 2.660 3.530 2.690 ;
        RECT 3.150 1.550 3.320 2.660 ;
        RECT 3.150 1.510 3.530 1.550 ;
        RECT 3.150 1.320 3.540 1.510 ;
        RECT 3.150 1.290 3.530 1.320 ;
        RECT 0.190 0.680 0.770 0.870 ;
        RECT 1.570 0.830 1.890 0.870 ;
        RECT 2.600 0.830 2.980 0.870 ;
        RECT 0.200 0.650 0.760 0.680 ;
        RECT 0.200 0.440 0.710 0.650 ;
        RECT 1.570 0.640 1.900 0.830 ;
        RECT 2.600 0.710 2.990 0.830 ;
        RECT 3.150 0.710 3.320 1.290 ;
        RECT 3.700 0.880 3.870 3.180 ;
        RECT 3.700 0.840 4.080 0.880 ;
        RECT 3.700 0.710 4.090 0.840 ;
        RECT 4.250 0.710 4.420 3.110 ;
        RECT 4.800 0.710 4.970 3.110 ;
        RECT 5.350 0.710 5.520 3.110 ;
        RECT 2.660 0.640 2.990 0.710 ;
        RECT 3.760 0.650 4.090 0.710 ;
        RECT 1.570 0.610 1.890 0.640 ;
        RECT 2.660 0.610 2.980 0.640 ;
        RECT 3.760 0.620 4.080 0.650 ;
        RECT 0.200 0.400 0.770 0.440 ;
        RECT 0.200 0.210 0.780 0.400 ;
        RECT 0.200 0.180 0.770 0.210 ;
        RECT 0.200 0.000 0.710 0.180 ;
      LAYER mcon ;
        RECT 1.080 5.480 1.250 5.650 ;
        RECT 2.170 5.480 2.340 5.650 ;
        RECT 3.270 5.470 3.440 5.640 ;
        RECT 1.630 4.800 1.800 4.970 ;
        RECT 2.720 4.780 2.890 4.950 ;
        RECT 1.630 3.430 1.800 3.600 ;
        RECT 2.720 3.430 2.890 3.600 ;
        RECT 3.830 4.770 4.000 4.940 ;
        RECT 3.820 3.430 3.990 3.600 ;
        RECT 1.070 2.700 1.240 2.870 ;
        RECT 2.170 2.700 2.340 2.870 ;
        RECT 0.240 2.250 0.410 2.420 ;
        RECT 0.240 1.890 0.410 2.060 ;
        RECT 1.070 1.330 1.240 1.500 ;
        RECT 2.170 1.330 2.340 1.500 ;
        RECT 3.270 2.700 3.440 2.870 ;
        RECT 3.270 1.330 3.440 1.500 ;
        RECT 0.500 0.690 0.670 0.860 ;
        RECT 1.630 0.650 1.800 0.820 ;
        RECT 2.720 0.650 2.890 0.820 ;
        RECT 3.820 0.660 3.990 0.830 ;
        RECT 0.510 0.220 0.680 0.390 ;
      LAYER met1 ;
        RECT 1.010 5.410 1.330 5.730 ;
        RECT 2.100 5.410 2.420 5.730 ;
        RECT 3.200 5.400 3.520 5.720 ;
        RECT 1.560 4.730 1.880 5.050 ;
        RECT 2.650 4.710 2.970 5.030 ;
        RECT 3.760 4.700 4.080 5.020 ;
        RECT 1.560 3.360 1.880 3.680 ;
        RECT 2.650 3.360 2.970 3.680 ;
        RECT 3.750 3.360 4.070 3.680 ;
        RECT 1.000 2.630 1.320 2.950 ;
        RECT 2.100 2.630 2.420 2.950 ;
        RECT 3.200 2.630 3.520 2.950 ;
        RECT 1.000 1.260 1.320 1.580 ;
        RECT 2.100 1.260 2.420 1.580 ;
        RECT 3.200 1.260 3.520 1.580 ;
        RECT 0.430 0.620 0.750 0.940 ;
        RECT 1.560 0.580 1.880 0.900 ;
        RECT 2.650 0.580 2.970 0.900 ;
        RECT 3.750 0.590 4.070 0.910 ;
        RECT 0.440 0.150 0.760 0.470 ;
      LAYER via ;
        RECT 1.040 5.440 1.300 5.700 ;
        RECT 2.130 5.440 2.390 5.700 ;
        RECT 3.230 5.430 3.490 5.690 ;
        RECT 1.590 4.760 1.850 5.020 ;
        RECT 2.680 4.740 2.940 5.000 ;
        RECT 3.790 4.730 4.050 4.990 ;
        RECT 1.590 3.390 1.850 3.650 ;
        RECT 2.680 3.390 2.940 3.650 ;
        RECT 3.780 3.390 4.040 3.650 ;
        RECT 1.030 2.660 1.290 2.920 ;
        RECT 2.130 2.660 2.390 2.920 ;
        RECT 3.230 2.660 3.490 2.920 ;
        RECT 1.030 1.290 1.290 1.550 ;
        RECT 2.130 1.290 2.390 1.550 ;
        RECT 3.230 1.290 3.490 1.550 ;
        RECT 0.460 0.650 0.720 0.910 ;
        RECT 1.590 0.610 1.850 0.870 ;
        RECT 2.680 0.610 2.940 0.870 ;
        RECT 3.780 0.620 4.040 0.880 ;
        RECT 0.470 0.180 0.730 0.440 ;
  END
END sky130_hilas_nFETLarge

END LIBRARY