magic
tech sky130A
timestamp 1634057778
<< checkpaint >>
rect 33 1301 1710 1351
rect -279 999 1710 1301
rect -280 -578 1710 999
rect 33 -630 1710 -578
<< error_s >>
rect 1 640 400 646
rect 1 598 400 604
rect 1 572 400 578
rect 1 530 400 536
rect 1 489 400 495
rect 1 447 400 453
rect 1 421 400 427
rect 1 379 400 385
rect 0 338 399 344
rect 0 296 399 302
rect 0 270 399 276
rect 0 228 399 234
rect 0 187 399 193
rect 0 145 399 151
rect 0 119 399 125
rect 0 77 399 83
<< nwell >>
rect 490 333 907 388
<< locali >>
rect 518 572 547 617
<< metal1 >>
rect 428 76 462 648
rect 824 589 867 653
rect 824 72 866 589
<< metal2 >>
rect 333 605 549 628
rect 359 391 924 414
rect 333 309 923 331
rect 332 92 560 115
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1634057699
transform 1 0 527 0 1 110
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1634057699
transform 1 0 525 0 1 409
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1634057699
transform 1 0 523 0 1 313
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1634057699
transform 1 0 524 0 1 605
box 0 0 34 33
use sky130_hilas_nMirror03_LongL  sky130_hilas_nMirror03_LongL_2
timestamp 1634057736
transform 1 0 350 0 1 227
box 0 0 562 142
use sky130_hilas_nMirror03_LongL  sky130_hilas_nMirror03_LongL_3
timestamp 1634057736
transform 1 0 350 0 -1 194
box 0 0 562 142
use sky130_hilas_nMirror03_LongL  sky130_hilas_nMirror03_LongL_1
timestamp 1634057736
transform 1 0 351 0 -1 496
box 0 0 562 142
use sky130_hilas_nMirror03_LongL  sky130_hilas_nMirror03_LongL_0
timestamp 1634057736
transform 1 0 351 0 1 529
box 0 0 562 142
use sky130_hilas_pFETmirror02_LongL  sky130_hilas_pFETmirror02_LongL_1
timestamp 1634057735
transform 1 0 663 0 1 0
box 0 0 417 235
use sky130_hilas_pFETmirror02_LongL  sky130_hilas_pFETmirror02_LongL_0
timestamp 1634057735
transform 1 0 663 0 -1 721
box 0 0 417 235
<< labels >>
rlabel metal2 613 391 624 414 0 output1
rlabel space 613 309 624 332 0 output2
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
