magic
tech sky130A
timestamp 1634057825
<< checkpaint >>
rect 359 2064 2168 2133
rect -234 -248 2680 2064
rect 1007 -589 2625 -248
<< error_s >>
rect 964 577 1014 583
rect 1036 577 1086 583
rect 964 535 1014 541
rect 1036 535 1086 541
rect 286 322 303 324
rect 286 303 303 305
rect 286 288 303 289
rect 1550 281 1577 287
rect 286 269 303 270
rect 1550 239 1577 245
rect 1550 214 1577 220
rect 1550 172 1577 178
rect 1550 131 1577 137
rect 1550 89 1577 95
rect 964 64 1014 70
rect 1036 64 1086 70
rect 1550 64 1577 70
rect 964 22 1014 28
rect 1036 22 1086 28
rect 1550 22 1577 28
<< nwell >>
rect 1145 431 1311 453
rect 1664 0 1792 19
<< locali >>
rect 283 339 329 348
rect 283 322 286 339
rect 303 322 329 339
rect 1324 330 1342 353
rect 283 270 329 322
rect 1236 295 1342 330
rect 1256 278 1262 295
rect 283 253 286 270
rect 303 253 329 270
rect 283 247 329 253
<< viali >>
rect 286 322 303 339
rect 286 253 303 270
<< metal1 >>
rect 35 598 77 605
rect 405 597 428 605
rect 1057 597 1076 605
rect 1101 597 1129 605
rect 1596 591 1630 605
rect 1663 590 1690 605
rect 1600 439 1626 465
rect 1595 392 1638 395
rect 1595 358 1600 392
rect 1634 358 1638 392
rect 1595 356 1638 358
rect 1600 355 1634 356
rect 279 344 317 348
rect 279 251 283 344
rect 312 251 317 344
rect 279 247 317 251
rect 1596 0 1630 19
rect 1663 0 1690 21
<< via1 >>
rect 1600 358 1634 392
rect 283 339 312 344
rect 283 322 286 339
rect 286 322 303 339
rect 303 322 312 339
rect 283 270 312 322
rect 283 253 286 270
rect 286 253 303 270
rect 303 253 312 270
rect 283 251 312 253
<< metal2 >>
rect 0 537 7 555
rect 1145 431 1792 453
rect 1597 392 1637 393
rect 1597 384 1600 392
rect 282 365 1600 384
rect 282 347 301 365
rect 1431 351 1470 365
rect 1597 358 1600 365
rect 1634 358 1637 392
rect 1597 357 1637 358
rect 280 344 315 347
rect 280 251 283 344
rect 312 251 315 344
rect 1411 252 1508 294
rect 280 248 315 251
rect 1296 187 1473 207
rect 1139 138 1155 178
rect 1267 106 1473 127
rect 0 52 8 67
rect 1187 2 1213 27
use sky130_hilas_pTransistorSingle  sky130_hilas_pTransistorSingle_0
timestamp 1634057769
transform 1 0 1150 0 1 440
box 0 0 549 779
use sky130_hilas_SingleTACore01  sky130_hilas_SingleTACore01_0
timestamp 1634057770
transform 1 0 1637 0 1 41
box 0 0 358 661
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_0
timestamp 1634057767
transform 1 0 989 0 1 440
box 0 0 549 1063
use sky130_hilas_FGBias2x1cell  sky130_hilas_FGBias2x1cell_0
timestamp 1634057765
transform 1 0 396 0 1 382
box 0 0 1654 1052
<< labels >>
rlabel metal1 1596 0 1630 6 0 VGND
port 7 nsew ground default
rlabel metal1 1663 0 1690 6 0 VPWR
port 8 nsew power default
rlabel metal1 1596 600 1630 605 0 VGND
port 7 nsew ground default
rlabel metal1 1663 600 1690 605 0 VPWR
port 8 nsew power default
rlabel metal2 1187 2 1210 27 0 VIN
port 2 nsew analog default
rlabel metal1 1057 597 1076 605 0 COLSEL1
port 1 nsew
rlabel metal2 0 537 7 555 0 DRAIN1
port 9 nsew
rlabel metal2 0 52 8 67 0 DRAIN2
port 10 nsew
rlabel metal1 35 598 77 605 0 VTUN
port 11 nsew
rlabel metal1 405 597 428 605 0 GATE1
port 12 nsew
rlabel metal1 1101 597 1129 605 0 VINJ
port 13 nsew
rlabel metal2 1776 431 1792 453 0 OUTPUT
port 14 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
