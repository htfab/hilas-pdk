magic
tech sky130A
timestamp 1629137251
<< checkpaint >>
rect -629 -630 2655 1720
<< error_s >>
rect 432 605 438 611
rect 537 605 543 611
rect 58 595 64 601
rect 111 595 117 601
rect 52 545 58 551
rect 117 545 123 551
rect 426 541 432 547
rect 543 541 549 547
rect 58 486 64 492
rect 111 486 117 492
rect 432 488 438 494
rect 537 488 543 494
rect 52 436 58 442
rect 117 436 123 442
rect 426 424 432 430
rect 543 424 549 430
rect 3635 348 3637 376
rect 432 303 438 309
rect 537 303 543 309
rect 58 297 64 303
rect 111 297 117 303
rect 52 247 58 253
rect 117 247 123 253
rect 426 239 432 245
rect 543 239 549 245
rect 432 187 438 193
rect 537 187 543 193
rect 58 180 64 186
rect 111 180 117 186
rect 52 130 58 136
rect 117 130 123 136
rect 426 123 432 129
rect 543 123 549 129
<< nwell >>
rect 1007 667 3542 668
rect 1008 660 3542 667
rect 1 600 12 618
rect 0 414 12 432
rect 2 115 12 132
rect 1006 69 3542 660
rect 1007 64 3542 69
rect 1200 63 3542 64
<< metal1 >>
rect 36 654 76 668
rect 280 662 304 668
rect 442 660 479 668
rect 673 661 697 668
rect 912 663 931 668
rect 956 663 972 668
rect 441 655 479 660
rect 440 76 441 78
rect 36 63 75 75
rect 280 63 304 70
rect 440 64 479 76
rect 440 63 441 64
rect 673 63 697 70
rect 875 64 891 70
rect 912 64 931 70
rect 956 64 972 70
<< metal2 >>
rect 1074 665 1125 668
rect 1074 663 1167 665
rect 1074 656 1130 663
rect 888 637 1130 656
rect 1117 635 1130 637
rect 1158 635 1167 663
rect 1 600 12 618
rect 898 600 3670 618
rect 892 557 3670 575
rect 898 457 3670 475
rect 3569 432 3670 433
rect 0 414 12 432
rect 894 414 3670 432
rect 3601 376 3670 383
rect 3601 348 3608 376
rect 3637 348 3670 376
rect 3601 342 3670 348
rect 2 299 12 316
rect 877 299 3670 316
rect 887 257 3670 274
rect 885 159 3670 176
rect 2 115 12 132
rect 881 115 3670 132
<< via2 >>
rect 1130 635 1158 663
rect 3608 348 3637 376
<< metal3 >>
rect 1125 663 1163 666
rect 1125 637 1130 663
rect 1117 635 1130 637
rect 1158 637 1163 663
rect 1158 635 1171 637
rect 1117 512 1171 635
rect 3523 376 3638 447
rect 3523 348 3608 376
rect 3637 348 3638 376
rect 1037 263 1055 293
rect 3523 283 3638 348
rect 3568 282 3638 283
rect 1146 142 1164 172
<< metal4 >>
rect 1279 601 1689 631
rect 1110 540 1380 551
rect 1110 510 1401 540
rect 1350 476 1401 510
rect 1651 481 1689 601
rect 1935 484 2263 514
rect 1041 438 1177 468
rect 1147 382 1177 438
rect 1935 382 1965 484
rect 2233 382 2263 484
rect 1147 352 2263 382
rect 2503 482 3392 512
rect 1371 293 1690 296
rect 1935 293 1965 296
rect 1037 263 2257 293
rect 1371 226 1401 263
rect 1660 229 1690 263
rect 1935 229 1965 263
rect 1660 226 1965 229
rect 2227 226 2257 263
rect 1371 196 2257 226
rect 2503 230 2533 482
rect 2786 479 3097 482
rect 2786 230 2816 479
rect 3067 230 3097 479
rect 3362 230 3392 482
rect 2503 200 3398 230
rect 3067 199 3398 200
rect 1134 142 1185 172
rect 1155 118 1185 142
rect 3368 118 3398 199
rect 1155 88 3398 118
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_1
timestamp 1629137207
transform 1 0 264 0 1 445
box -263 -445 1761 645
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_0
timestamp 1629137207
transform 1 0 264 0 1 445
box -263 -445 1761 645
use sky130_hilas_m22m4  sky130_hilas_m22m4_1
timestamp 1629137164
transform 1 0 1002 0 1 468
box 0 0 79 75
use sky130_hilas_m22m4  sky130_hilas_m22m4_2
timestamp 1629137164
transform 1 0 998 0 1 259
box 0 0 79 75
use sky130_hilas_m22m4  sky130_hilas_m22m4_3
timestamp 1629137164
transform 1 0 1107 0 1 172
box 0 0 79 75
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1629137154
transform 1 0 876 0 1 644
box 0 0 32 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1629137154
transform 1 0 876 0 1 644
box 0 0 32 32
<< labels >>
rlabel metal2 3658 342 3670 383 0 CAPTERM2
port 1 nsew analog default
rlabel metal2 1074 655 1125 668 0 CAPTERM1
port 2 nsew analog default
rlabel metal1 912 663 931 668 0 GATESELECT
port 4 nsew
rlabel metal1 956 663 972 668 0 VINJ
port 3 nsew power default
rlabel metal1 442 655 479 668 0 GATE
port 6 nsew analog default
rlabel metal1 36 654 76 668 0 VTUN
port 5 nsew
rlabel metal1 36 63 75 75 0 VTUN
port 5 nsew
rlabel metal1 440 64 479 76 0 GATE
port 6 nsew
rlabel metal1 956 64 972 70 0 VINJ
rlabel metal1 875 64 891 70 0 CAPTERM1
rlabel metal1 912 64 931 70 0 GATESELECT
rlabel metal2 1 600 12 618 0 DRAIN1
port 8 nsew
rlabel metal2 0 414 12 432 0 DRAIN2
port 7 nsew
rlabel metal2 3660 115 3670 132 0 DRAIN4
port 10 nsew
rlabel metal2 3660 600 3670 618 0 DRAIN1
port 8 nsew
rlabel metal2 3659 414 3670 433 0 DRAIN2
port 7 nsew
rlabel metal2 3659 299 3670 316 0 DRAIN3
port 11 nsew
rlabel metal2 2 299 12 316 0 DRAIN3
port 11 nsew
rlabel metal2 2 115 12 132 0 DRAIN4
port 10 nsew
rlabel metal1 280 662 304 668 0 VGND
port 12 nsew
rlabel metal1 673 661 697 668 0 VGND
port 12 nsew
rlabel metal1 280 63 304 70 0 VGND
port 12 nsew
rlabel metal1 673 63 697 70 0 VGND
port 12 nsew
<< end >>
