magic
tech sky130A
timestamp 1625359887
<< psubdiff >>
rect 671 88 672 171
<< locali >>
rect 646 547 665 636
rect 646 82 672 171
<< metal1 >>
rect 341 598 376 661
rect 341 582 603 598
rect 637 607 744 661
rect 637 598 656 607
rect 629 582 656 598
rect 341 581 656 582
rect 682 581 744 607
rect 341 567 744 581
rect 341 566 656 567
rect 341 540 601 566
rect 627 541 656 566
rect 682 541 744 567
rect 627 540 744 541
rect 341 530 744 540
rect 341 476 744 499
rect 341 449 392 476
rect 419 449 447 476
rect 474 449 744 476
rect 341 419 744 449
rect 341 418 447 419
rect 341 391 391 418
rect 418 392 447 418
rect 474 392 744 419
rect 418 391 744 392
rect 341 335 744 391
rect 341 334 447 335
rect 341 307 392 334
rect 419 308 447 334
rect 474 308 744 335
rect 419 307 744 308
rect 341 284 744 307
rect 341 257 392 284
rect 419 282 744 284
rect 419 257 445 282
rect 341 255 445 257
rect 472 255 744 282
rect 341 220 744 255
rect 341 157 744 184
rect 341 131 617 157
rect 643 131 665 157
rect 691 131 744 157
rect 341 116 744 131
rect 341 90 615 116
rect 641 90 664 116
rect 690 90 744 116
rect 341 60 744 90
rect 341 57 377 60
rect 646 58 744 60
rect 645 57 744 58
<< via1 >>
rect 603 582 629 608
rect 656 581 682 607
rect 601 540 627 566
rect 656 541 682 567
rect 392 449 419 476
rect 447 449 474 476
rect 391 391 418 418
rect 447 392 474 419
rect 392 307 419 334
rect 447 308 474 335
rect 392 257 419 284
rect 445 255 472 282
rect 617 131 643 157
rect 665 131 691 157
rect 615 90 641 116
rect 664 90 690 116
<< metal2 >>
rect 377 476 507 661
rect 377 449 392 476
rect 419 449 447 476
rect 474 449 507 476
rect 377 419 507 449
rect 377 418 447 419
rect 377 391 391 418
rect 418 392 447 418
rect 474 392 507 419
rect 418 391 507 392
rect 377 335 507 391
rect 377 334 447 335
rect 377 307 392 334
rect 419 308 447 334
rect 474 308 507 335
rect 419 307 507 308
rect 377 284 507 307
rect 377 257 392 284
rect 419 282 507 284
rect 419 257 445 282
rect 377 255 445 257
rect 472 255 507 282
rect 377 57 507 255
rect 585 608 715 661
rect 585 582 603 608
rect 629 607 715 608
rect 629 582 656 607
rect 585 581 656 582
rect 682 581 715 607
rect 585 567 715 581
rect 585 566 656 567
rect 585 540 601 566
rect 627 541 656 566
rect 682 541 715 567
rect 627 540 715 541
rect 585 519 715 540
rect 585 189 714 519
rect 585 157 715 189
rect 585 131 617 157
rect 643 131 665 157
rect 691 131 715 157
rect 585 116 715 131
rect 585 90 615 116
rect 641 90 664 116
rect 690 90 715 116
rect 585 57 715 90
use sky130_hilas_DecoupVinj00  CapDeco_1
timestamp 1625358249
transform 1 0 273 0 1 170
box 68 -113 473 189
use sky130_hilas_DecoupVinj00  CapDeco_0
timestamp 1625358249
transform 1 0 273 0 -1 548
box 68 -113 473 189
<< labels >>
rlabel metal1 355 57 364 120 0 VGND 
port 1 nsew
rlabel metal1 729 57 744 120 0 VGND 
port 1 nsew
rlabel metal2 377 651 507 661 0 VINJ
port 1 nsew
rlabel metal2 585 653 715 661 0 VGND
port 2 nsew
rlabel metal2 377 57 507 69 0 VINJ
port 1 nsew
rlabel metal2 585 57 715 69 0 VGND
port 2 nsew
rlabel metal1 727 313 744 407 0 VINJ
port 1 nsew
rlabel metal1 341 311 358 407 0 VINJ
port 1 nsew
rlabel metal1 355 598 363 661 0 VGND
port 3 nsew
rlabel metal1 734 598 744 661 0 VGND
port 2 nsew
<< end >>
