magic
tech sky130A
timestamp 1634057710
<< error_p >>
rect 31 49 430 55
rect 31 7 430 13
<< nmos >>
rect 31 13 430 49
<< ndiff >>
rect 0 39 31 49
rect 0 22 5 39
rect 25 22 31 39
rect 0 13 31 22
rect 430 39 463 49
rect 430 22 436 39
rect 456 22 463 39
rect 430 13 463 22
<< ndiffc >>
rect 5 22 25 39
rect 436 22 456 39
<< poly >>
rect 31 49 430 62
rect 31 0 430 13
<< locali >>
rect 5 39 25 47
rect 5 14 25 22
rect 436 39 456 47
rect 436 14 456 22
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
