magic
tech sky130A
timestamp 1629137189
<< checkpaint >>
rect -895 1265 765 1289
rect 1032 1265 2692 1289
rect -895 -575 2692 1265
rect -895 -576 886 -575
rect -630 -635 886 -576
rect 911 -576 2692 -575
rect 911 -635 2427 -576
<< error_s >>
rect 323 572 352 588
rect 402 572 431 588
rect 481 572 510 588
rect 560 572 589 588
rect 806 574 835 592
rect 962 574 991 592
rect 1208 572 1237 588
rect 1287 572 1316 588
rect 1366 572 1395 588
rect 1445 572 1474 588
rect 806 542 807 543
rect 834 542 835 543
rect 962 542 963 543
rect 990 542 991 543
rect 323 538 324 539
rect 351 538 352 539
rect 402 538 403 539
rect 430 538 431 539
rect 481 538 482 539
rect 509 538 510 539
rect 560 538 561 539
rect 588 538 589 539
rect 273 509 290 538
rect 322 537 353 538
rect 401 537 432 538
rect 480 537 511 538
rect 559 537 590 538
rect 323 530 352 537
rect 402 530 431 537
rect 481 530 510 537
rect 560 530 589 537
rect 323 516 332 530
rect 579 516 589 530
rect 323 510 352 516
rect 402 510 431 516
rect 481 510 510 516
rect 560 510 589 516
rect 322 509 353 510
rect 401 509 432 510
rect 480 509 511 510
rect 559 509 590 510
rect 621 509 639 538
rect 756 513 774 542
rect 805 541 836 542
rect 806 532 835 541
rect 806 523 816 532
rect 825 523 835 532
rect 806 514 835 523
rect 805 513 836 514
rect 867 513 885 542
rect 912 513 930 542
rect 961 541 992 542
rect 962 532 991 541
rect 962 523 972 532
rect 981 523 991 532
rect 962 514 991 523
rect 961 513 992 514
rect 1023 513 1041 542
rect 1208 538 1209 539
rect 1236 538 1237 539
rect 1287 538 1288 539
rect 1315 538 1316 539
rect 1366 538 1367 539
rect 1394 538 1395 539
rect 1445 538 1446 539
rect 1473 538 1474 539
rect 806 512 807 513
rect 834 512 835 513
rect 962 512 963 513
rect 990 512 991 513
rect 1158 509 1176 538
rect 1207 537 1238 538
rect 1286 537 1317 538
rect 1365 537 1396 538
rect 1444 537 1475 538
rect 1208 530 1237 537
rect 1287 530 1316 537
rect 1366 530 1395 537
rect 1445 530 1474 537
rect 1208 516 1218 530
rect 1465 516 1474 530
rect 1208 510 1237 516
rect 1287 510 1316 516
rect 1366 510 1395 516
rect 1445 510 1474 516
rect 1207 509 1238 510
rect 1286 509 1317 510
rect 1365 509 1396 510
rect 1444 509 1475 510
rect 1507 509 1524 538
rect 1541 516 1543 517
rect 323 508 324 509
rect 351 508 352 509
rect 402 508 403 509
rect 430 508 431 509
rect 481 508 482 509
rect 509 508 510 509
rect 560 508 561 509
rect 588 508 589 509
rect 1208 508 1209 509
rect 1236 508 1237 509
rect 1287 508 1288 509
rect 1315 508 1316 509
rect 1366 508 1367 509
rect 1394 508 1395 509
rect 1445 508 1446 509
rect 1473 508 1474 509
rect 323 459 352 474
rect 402 459 431 474
rect 481 459 510 474
rect 560 459 589 474
rect 806 463 835 481
rect 962 463 991 481
rect 1208 459 1237 474
rect 1287 459 1316 474
rect 1366 459 1395 474
rect 1445 459 1474 474
rect 323 425 352 441
rect 402 425 431 441
rect 481 425 510 441
rect 560 425 589 441
rect 806 422 835 440
rect 962 422 991 440
rect 1208 425 1237 441
rect 1287 425 1316 441
rect 1366 425 1395 441
rect 1445 425 1474 441
rect 323 391 324 392
rect 351 391 352 392
rect 402 391 403 392
rect 430 391 431 392
rect 481 391 482 392
rect 509 391 510 392
rect 560 391 561 392
rect 588 391 589 392
rect 1208 391 1209 392
rect 1236 391 1237 392
rect 1287 391 1288 392
rect 1315 391 1316 392
rect 1366 391 1367 392
rect 1394 391 1395 392
rect 1445 391 1446 392
rect 1473 391 1474 392
rect 273 362 290 391
rect 322 390 353 391
rect 401 390 432 391
rect 480 390 511 391
rect 559 390 590 391
rect 323 383 352 390
rect 402 383 431 390
rect 481 383 510 390
rect 560 383 589 390
rect 323 369 332 383
rect 579 369 589 383
rect 323 363 352 369
rect 402 363 431 369
rect 481 363 510 369
rect 560 363 589 369
rect 322 362 353 363
rect 401 362 432 363
rect 480 362 511 363
rect 559 362 590 363
rect 621 362 639 391
rect 806 390 807 391
rect 834 390 835 391
rect 962 390 963 391
rect 990 390 991 391
rect 323 361 324 362
rect 351 361 352 362
rect 402 361 403 362
rect 430 361 431 362
rect 481 361 482 362
rect 509 361 510 362
rect 560 361 561 362
rect 588 361 589 362
rect 756 361 774 390
rect 805 389 836 390
rect 806 380 835 389
rect 806 371 816 380
rect 825 371 835 380
rect 806 362 835 371
rect 805 361 836 362
rect 867 361 885 390
rect 912 361 930 390
rect 961 389 992 390
rect 962 380 991 389
rect 962 371 972 380
rect 981 371 991 380
rect 962 362 991 371
rect 961 361 992 362
rect 1023 361 1041 390
rect 1158 362 1176 391
rect 1207 390 1238 391
rect 1286 390 1317 391
rect 1365 390 1396 391
rect 1444 390 1475 391
rect 1208 383 1237 390
rect 1287 383 1316 390
rect 1366 383 1395 390
rect 1445 383 1474 390
rect 1208 369 1218 383
rect 1465 369 1474 383
rect 1208 363 1237 369
rect 1287 363 1316 369
rect 1366 363 1395 369
rect 1445 363 1474 369
rect 1207 362 1238 363
rect 1286 362 1317 363
rect 1365 362 1396 363
rect 1444 362 1475 363
rect 1507 362 1524 391
rect 1208 361 1209 362
rect 1236 361 1237 362
rect 1287 361 1288 362
rect 1315 361 1316 362
rect 1366 361 1367 362
rect 1394 361 1395 362
rect 1445 361 1446 362
rect 1473 361 1474 362
rect 806 360 807 361
rect 834 360 835 361
rect 962 360 963 361
rect 990 360 991 361
rect 323 312 352 327
rect 402 312 431 327
rect 481 312 510 327
rect 560 312 589 327
rect 806 311 835 329
rect 962 311 991 329
rect 1208 312 1237 327
rect 1287 312 1316 327
rect 1366 312 1395 327
rect 1445 312 1474 327
rect 323 278 352 294
rect 402 278 431 294
rect 481 278 510 294
rect 560 278 589 294
rect 806 277 835 295
rect 962 277 991 295
rect 1208 278 1237 294
rect 1287 278 1316 294
rect 1366 278 1395 294
rect 1445 278 1474 294
rect 806 245 807 246
rect 834 245 835 246
rect 962 245 963 246
rect 990 245 991 246
rect 323 244 324 245
rect 351 244 352 245
rect 402 244 403 245
rect 430 244 431 245
rect 481 244 482 245
rect 509 244 510 245
rect 560 244 561 245
rect 588 244 589 245
rect 273 215 290 244
rect 322 243 353 244
rect 401 243 432 244
rect 480 243 511 244
rect 559 243 590 244
rect 323 236 352 243
rect 402 236 431 243
rect 481 236 510 243
rect 560 236 589 243
rect 323 222 332 236
rect 579 222 589 236
rect 323 216 352 222
rect 402 216 431 222
rect 481 216 510 222
rect 560 216 589 222
rect 322 215 353 216
rect 401 215 432 216
rect 480 215 511 216
rect 559 215 590 216
rect 621 215 639 244
rect 756 216 774 245
rect 805 244 836 245
rect 806 235 835 244
rect 806 226 816 235
rect 825 226 835 235
rect 806 217 835 226
rect 805 216 836 217
rect 867 216 885 245
rect 912 216 930 245
rect 961 244 992 245
rect 962 235 991 244
rect 962 226 972 235
rect 981 226 991 235
rect 962 217 991 226
rect 961 216 992 217
rect 1023 216 1041 245
rect 1208 244 1209 245
rect 1236 244 1237 245
rect 1287 244 1288 245
rect 1315 244 1316 245
rect 1366 244 1367 245
rect 1394 244 1395 245
rect 1445 244 1446 245
rect 1473 244 1474 245
rect 806 215 807 216
rect 834 215 835 216
rect 962 215 963 216
rect 990 215 991 216
rect 1158 215 1176 244
rect 1207 243 1238 244
rect 1286 243 1317 244
rect 1365 243 1396 244
rect 1444 243 1475 244
rect 1208 236 1237 243
rect 1287 236 1316 243
rect 1366 236 1395 243
rect 1445 236 1474 243
rect 1208 222 1218 236
rect 1465 222 1474 236
rect 1208 216 1237 222
rect 1287 216 1316 222
rect 1366 216 1395 222
rect 1445 216 1474 222
rect 1207 215 1238 216
rect 1286 215 1317 216
rect 1365 215 1396 216
rect 1444 215 1475 216
rect 1507 215 1524 244
rect 323 214 324 215
rect 351 214 352 215
rect 402 214 403 215
rect 430 214 431 215
rect 481 214 482 215
rect 509 214 510 215
rect 560 214 561 215
rect 588 214 589 215
rect 1208 214 1209 215
rect 1236 214 1237 215
rect 1287 214 1288 215
rect 1315 214 1316 215
rect 1366 214 1367 215
rect 1394 214 1395 215
rect 1445 214 1446 215
rect 1473 214 1474 215
rect 323 165 352 180
rect 402 165 431 180
rect 481 165 510 180
rect 560 165 589 180
rect 806 166 835 184
rect 962 166 991 184
rect 1208 165 1237 180
rect 1287 165 1316 180
rect 1366 165 1395 180
rect 1445 165 1474 180
rect 323 131 352 147
rect 402 131 431 147
rect 481 131 510 147
rect 560 131 589 147
rect 806 123 835 141
rect 962 123 991 141
rect 1208 131 1237 147
rect 1287 131 1316 147
rect 1366 131 1395 147
rect 1445 131 1474 147
rect 323 97 324 98
rect 351 97 352 98
rect 402 97 403 98
rect 430 97 431 98
rect 481 97 482 98
rect 509 97 510 98
rect 560 97 561 98
rect 588 97 589 98
rect 1208 97 1209 98
rect 1236 97 1237 98
rect 1287 97 1288 98
rect 1315 97 1316 98
rect 1366 97 1367 98
rect 1394 97 1395 98
rect 1445 97 1446 98
rect 1473 97 1474 98
rect 273 68 290 97
rect 322 96 353 97
rect 401 96 432 97
rect 480 96 511 97
rect 559 96 590 97
rect 323 89 352 96
rect 402 89 431 96
rect 481 89 510 96
rect 560 89 589 96
rect 323 75 332 89
rect 579 75 589 89
rect 323 69 352 75
rect 402 69 431 75
rect 481 69 510 75
rect 560 69 589 75
rect 322 68 353 69
rect 401 68 432 69
rect 480 68 511 69
rect 559 68 590 69
rect 621 68 639 97
rect 806 91 807 92
rect 834 91 835 92
rect 962 91 963 92
rect 990 91 991 92
rect 323 67 324 68
rect 351 67 352 68
rect 402 67 403 68
rect 430 67 431 68
rect 481 67 482 68
rect 509 67 510 68
rect 560 67 561 68
rect 588 67 589 68
rect 756 62 774 91
rect 805 90 836 91
rect 806 81 835 90
rect 806 72 816 81
rect 825 72 835 81
rect 806 63 835 72
rect 805 62 836 63
rect 867 62 885 91
rect 912 62 930 91
rect 961 90 992 91
rect 962 81 991 90
rect 962 72 972 81
rect 981 72 991 81
rect 962 63 991 72
rect 961 62 992 63
rect 1023 62 1041 91
rect 1158 68 1176 97
rect 1207 96 1238 97
rect 1286 96 1317 97
rect 1365 96 1396 97
rect 1444 96 1475 97
rect 1208 89 1237 96
rect 1287 89 1316 96
rect 1366 89 1395 96
rect 1445 89 1474 96
rect 1208 75 1218 89
rect 1465 75 1474 89
rect 1208 69 1237 75
rect 1287 69 1316 75
rect 1366 69 1395 75
rect 1445 69 1474 75
rect 1207 68 1238 69
rect 1286 68 1317 69
rect 1365 68 1396 69
rect 1444 68 1475 69
rect 1507 68 1524 97
rect 1208 67 1209 68
rect 1236 67 1237 68
rect 1287 67 1288 68
rect 1315 67 1316 68
rect 1366 67 1367 68
rect 1394 67 1395 68
rect 1445 67 1446 68
rect 1473 67 1474 68
rect 806 61 807 62
rect 834 61 835 62
rect 962 61 963 62
rect 990 61 991 62
rect 323 18 352 33
rect 402 18 431 33
rect 481 18 510 33
rect 560 18 589 33
rect 806 12 835 30
rect 962 12 991 30
rect 1208 18 1237 33
rect 1287 18 1316 33
rect 1366 18 1395 33
rect 1445 18 1474 33
<< metal1 >>
rect 36 599 52 605
rect 77 599 96 605
rect 117 599 133 605
rect 36 1 52 8
rect 77 1 96 8
rect 117 1 133 8
rect 444 0 469 605
rect 805 0 835 605
rect 963 0 993 605
rect 1329 0 1353 605
rect 1664 598 1680 605
rect 1701 598 1720 605
rect 1745 598 1761 605
rect 1664 1 1680 8
rect 1701 1 1720 8
rect 1745 1 1761 8
<< metal2 >>
rect 0 537 8 555
rect 1786 537 1797 555
rect 0 494 8 512
rect 1787 494 1798 512
rect 0 394 8 412
rect 1787 394 1798 412
rect 0 351 8 369
rect 240 361 252 369
rect 1549 355 1561 369
rect 1787 351 1798 369
rect 0 236 7 254
rect 1786 236 1797 254
rect 0 193 7 211
rect 1786 193 1797 211
rect 0 94 7 112
rect 1786 94 1797 112
rect 0 51 7 69
rect 1786 51 1797 69
use sky130_hilas_swc4x1cellOverlap2  sky130_hilas_swc4x1cellOverlap2_0
timestamp 1607392100
transform 1 0 1053 0 1 382
box -191 -387 1009 277
use sky130_hilas_swc4x1cellOverlap2  sky130_hilas_swc4x1cellOverlap2_1
timestamp 1607392100
transform -1 0 744 0 1 382
box -191 -387 1009 277
<< labels >>
rlabel metal1 117 599 133 605 0 VERT1
port 1 nsew analog default
rlabel metal1 36 599 52 605 0 VINJ
port 10 nsew
rlabel metal1 77 599 96 605 0 GATESELECT1
port 11 nsew analog default
rlabel metal2 0 537 8 555 0 DRAIN1
port 3 nsew analog default
rlabel metal2 0 494 8 512 0 HORIZ1
port 2 nsew analog default
rlabel metal2 0 394 8 412 0 HORIZ2
port 4 nsew analog default
rlabel metal2 0 351 8 369 0 DRAIN2
port 5 nsew analog default
rlabel metal2 0 236 7 254 0 DRAIN3
port 6 nsew analog default
rlabel metal2 0 193 7 211 0 HORIZ3
port 7 nsew analog default
rlabel metal2 0 94 7 112 0 HORIZ4
port 8 nsew analog default
rlabel metal2 0 51 7 69 0 DRAIN4
port 9 nsew analog default
rlabel metal1 36 1 52 8 0 VINJ
port 10 nsew power default
rlabel metal1 117 1 133 8 0 VERT1
port 1 nsew analog default
rlabel metal1 77 1 96 8 0 GATESELECT1
port 11 nsew analog default
rlabel metal1 1745 1 1761 8 0 VINJ
port 10 nsew power default
rlabel metal1 1664 598 1680 605 0 VERT2
port 12 nsew analog default
rlabel metal1 1701 598 1720 605 0 GATESELECT2
port 13 nsew analog default
rlabel metal1 1745 598 1761 605 0 VINJ
port 10 nsew power default
rlabel metal1 1664 1 1680 8 0 VERT2
port 12 nsew analog default
rlabel metal1 1701 1 1720 8 0 GATESELECT2
port 13 nsew analog default
rlabel metal2 1786 537 1797 555 0 DRAIN1
port 3 nsew analog default
rlabel metal2 1787 494 1798 512 0 HORIZ1
port 2 nsew analog default
rlabel metal2 1787 394 1798 412 0 HORIZ2
port 4 nsew analog default
rlabel metal2 1787 351 1798 369 0 DRAIN2
port 5 nsew analog default
rlabel metal2 1786 236 1797 254 0 DRAIN3
port 6 nsew analog default
rlabel metal2 1786 193 1797 211 0 HORIZ3
port 7 nsew analog default
rlabel metal2 1786 94 1797 112 0 HORIZ4
port 8 nsew analog default
rlabel metal2 1786 51 1797 69 0 DRAIN
port 14 nsew analog default
rlabel metal1 1329 600 1353 605 0 GATE2
port 15 nsew analog default
rlabel metal1 1329 0 1353 6 0 GATE2
port 15 nsew analog default
rlabel metal1 444 599 469 605 0 GATE1
port 16 nsew analog default
rlabel metal1 444 0 469 6 0 GATE1
port 16 nsew analog default
rlabel metal1 805 597 835 605 0 VTUN
port 17 nsew analog default
rlabel metal1 963 597 993 605 0 VTUN
rlabel metal1 805 0 835 8 0 VTUN
port 17 nsew analog default
rlabel metal1 963 0 993 8 0 VTUN
port 17 nsew analog default
<< end >>
