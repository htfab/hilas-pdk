magic
tech sky130A
timestamp 1628707358
<< error_s >>
rect 84 660 134 666
rect 407 661 457 667
rect 564 660 592 667
rect 706 661 734 667
rect 84 618 134 624
rect 407 619 457 625
rect 564 618 592 625
rect 706 619 734 625
rect 155 594 205 600
rect 335 589 386 595
rect 515 589 543 595
rect 755 589 783 595
rect 155 552 205 558
rect 335 547 386 553
rect 515 547 543 553
rect 755 547 783 553
rect 84 485 134 491
rect 407 486 457 492
rect 564 485 592 492
rect 706 486 734 492
rect 84 443 134 449
rect 407 444 457 450
rect 564 443 592 450
rect 706 444 734 450
rect 155 419 205 425
rect 335 414 386 420
rect 515 414 543 420
rect 755 414 783 420
rect 155 377 205 383
rect 335 372 386 378
rect 515 372 543 378
rect 755 372 783 378
rect 84 310 134 316
rect 407 311 457 317
rect 564 310 592 317
rect 706 311 734 317
rect 84 268 134 274
rect 407 269 457 275
rect 564 268 592 275
rect 706 269 734 275
rect 155 244 205 250
rect 335 239 386 245
rect 515 239 543 245
rect 755 239 783 245
rect 155 202 205 208
rect 335 197 386 203
rect 515 197 543 203
rect 755 197 783 203
rect 84 135 134 141
rect 407 136 457 142
rect 564 135 592 142
rect 706 136 734 142
rect 84 93 134 99
rect 407 94 457 100
rect 564 93 592 100
rect 706 94 734 100
rect 155 69 205 75
rect 335 64 386 70
rect 515 64 543 70
rect 755 64 783 70
rect 155 27 205 33
rect 335 22 386 28
rect 515 22 543 28
rect 755 22 783 28
<< nwell >>
rect 19 576 30 596
<< metal1 >>
rect 53 691 82 700
rect 484 694 515 700
rect 785 695 809 700
rect 53 0 82 12
rect 484 0 515 6
rect 785 0 809 5
<< metal2 >>
rect 19 636 35 656
rect 879 543 889 575
rect 19 461 36 481
rect 879 368 889 400
rect 19 286 38 306
rect 879 193 889 225
rect 19 111 35 131
rect 879 18 889 50
use sky130_hilas_StepUpDigital  StepUpDigital_2
timestamp 1628707339
transform 1 0 0 0 1 569
box 0 0 836 218
use sky130_hilas_StepUpDigital  StepUpDigital_1
timestamp 1628707339
transform 1 0 0 0 1 394
box 0 0 836 218
use sky130_hilas_StepUpDigital  StepUpDigital_3
timestamp 1628707339
transform 1 0 0 0 1 44
box 0 0 836 218
use sky130_hilas_StepUpDigital  StepUpDigital_0
timestamp 1628707339
transform 1 0 0 0 1 219
box 0 0 836 218
<< labels >>
rlabel metal1 53 4 82 9 0 VINJ
port 6 nsew
rlabel metal2 19 111 30 131 0 OUTPUT4
port 10 nsew
rlabel metal2 879 543 889 575 0 INPUT1
port 12 nsew
rlabel metal2 879 368 889 400 0 INPUT2
port 13 nsew
rlabel metal2 879 193 889 225 0 INPUT3
port 14 nsew
rlabel metal2 879 18 889 50 0 INPUT4
port 15 nsew
rlabel metal2 19 286 27 306 0 OUTPUT3
port 9 nsew
rlabel metal2 19 461 26 481 0 OUTPUT2
port 8 nsew
rlabel metal2 19 636 26 656 0 OUTPUT1
port 7 nsew
rlabel metal1 484 0 515 6 0 VGND
port 11 nsew
rlabel metal1 484 694 515 700 0 VGND
port 11 nsew
rlabel metal1 53 691 82 700 0 VINJ
port 6 nsew
rlabel metal1 785 695 809 700 0 VPWR
port 5 nsew
rlabel metal1 785 0 809 5 0 VPWR
port 5 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
