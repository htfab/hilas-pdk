magic
tech sky130A
magscale 1 2
timestamp 1627400561
<< error_s >>
rect 106 1318 164 1346
rect 988 1314 1050 1342
rect 1590 1318 1638 1346
rect 38 1224 66 1264
rect 130 1182 230 1204
rect 230 1171 298 1182
rect 796 1176 896 1194
rect 896 1165 958 1176
rect 1110 1164 1166 1196
rect 1394 1164 1450 1196
rect 130 1098 230 1120
rect 428 1096 462 1105
rect 796 1092 896 1110
rect 82 1080 116 1082
rect 1110 1080 1166 1112
rect 1394 1080 1450 1112
rect 272 1058 372 1080
rect 82 1042 116 1044
rect 652 1040 754 1060
rect 588 1031 625 1040
rect 1012 1038 1068 1072
rect 1492 1038 1548 1072
rect 372 996 436 1005
rect 272 974 372 996
rect 588 976 597 1031
rect 1780 1028 1808 1092
rect 1752 1006 1760 1012
rect 754 976 816 987
rect 652 956 754 976
rect 1012 954 1068 988
rect 1492 954 1548 988
rect 38 914 66 954
rect 130 872 230 894
rect 230 861 298 872
rect 796 866 896 884
rect 896 855 958 866
rect 1110 854 1166 886
rect 1394 854 1450 886
rect 130 788 230 810
rect 428 786 462 795
rect 796 782 896 800
rect 82 770 116 772
rect 1110 770 1166 802
rect 1394 770 1450 802
rect 272 748 372 770
rect 82 732 116 734
rect 652 730 754 750
rect 588 721 625 730
rect 1012 728 1068 762
rect 1492 728 1548 762
rect 372 686 436 695
rect 272 664 372 686
rect 588 666 597 721
rect 1780 718 1808 782
rect 1752 696 1760 702
rect 754 666 816 677
rect 652 646 754 666
rect 1012 644 1068 678
rect 1492 644 1548 678
rect 38 604 66 644
rect 130 562 230 584
rect 230 551 298 562
rect 796 556 896 574
rect 896 545 958 556
rect 1110 544 1166 576
rect 1394 544 1450 576
rect 130 478 230 500
rect 428 476 462 485
rect 796 472 896 490
rect 82 460 116 462
rect 1110 460 1166 492
rect 1394 460 1450 492
rect 272 438 372 460
rect 82 422 116 424
rect 652 420 754 440
rect 588 411 625 420
rect 1012 418 1068 452
rect 1492 418 1548 452
rect 372 376 436 385
rect 272 354 372 376
rect 588 356 597 411
rect 1780 408 1808 472
rect 1752 386 1760 392
rect 754 356 816 367
rect 652 336 754 356
rect 1012 334 1068 368
rect 1492 334 1548 368
rect 38 294 66 334
rect 130 252 230 274
rect 230 241 298 252
rect 796 246 896 264
rect 896 235 958 246
rect 1110 234 1166 266
rect 1394 234 1450 266
rect 130 168 230 190
rect 428 166 462 175
rect 796 162 896 180
rect 82 150 116 152
rect 1110 150 1166 182
rect 1394 150 1450 182
rect 272 128 372 150
rect 82 112 116 114
rect 652 110 754 130
rect 126 90 164 108
rect 588 101 625 110
rect 1012 108 1068 142
rect 1492 108 1548 142
rect 372 66 436 75
rect 272 44 372 66
rect 588 46 597 101
rect 1012 92 1050 108
rect 1600 90 1638 108
rect 1780 98 1808 162
rect 1752 76 1760 82
rect 754 46 816 57
rect 652 26 754 46
rect 1012 24 1068 58
rect 1492 24 1548 58
<< metal1 >>
rect 106 1318 164 1328
rect 988 1314 1050 1328
rect 1590 1318 1638 1328
rect 106 80 164 90
rect 988 80 1050 92
rect 1590 80 1638 90
<< metal2 >>
rect 38 1224 60 1264
rect 1780 1028 1798 1092
rect 38 914 60 954
rect 1780 718 1798 782
rect 38 604 60 644
rect 1780 408 1798 472
rect 38 294 60 334
rect 1780 98 1798 162
use sky130_hilas_StepUpDigital  StepUpDigital_3
timestamp 1627063084
transform 1 0 0 0 1 160
box 0 -160 1760 158
use sky130_hilas_StepUpDigital  StepUpDigital_0
timestamp 1627063084
transform 1 0 0 0 1 470
box 0 -160 1760 158
use sky130_hilas_StepUpDigital  StepUpDigital_1
timestamp 1627063084
transform 1 0 0 0 1 780
box 0 -160 1760 158
use sky130_hilas_StepUpDigital  StepUpDigital_2
timestamp 1627063084
transform 1 0 0 0 1 1090
box 0 -160 1760 158
<< labels >>
rlabel metal2 1780 1028 1798 1092 0 INPUT1
port 1 nsew
rlabel metal2 1780 718 1798 782 0 INPUT2
port 2 nsew
rlabel metal2 1780 408 1798 472 0 INPUT3
port 3 nsew
rlabel metal2 1780 98 1798 162 0 INPUT4
port 4 nsew
rlabel metal1 1590 1318 1638 1328 0 VPWR
port 5 nsew
rlabel metal1 1590 80 1638 90 0 VPWR
port 5 nsew
rlabel metal1 106 1318 164 1328 0 VINJ
port 6 nsew
rlabel metal1 106 80 164 90 0 VINJ
port 6 nsew
rlabel metal2 38 1224 60 1264 0 OUTPUT1
port 7 nsew
rlabel metal2 38 914 60 954 0 OUTPUT2
port 8 nsew
rlabel metal2 38 604 60 644 0 OUTPUT3
port 9 nsew
rlabel metal2 38 294 60 334 0 OUTPUT4
port 10 nsew
rlabel metal1 988 1314 1050 1328 0 VGND
port 11 nsew
rlabel metal1 988 80 1050 92 0 VGND
port 11 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
