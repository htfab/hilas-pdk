magic
tech sky130A
timestamp 1628707347
<< checkpaint >>
rect -544 657 749 666
rect -544 -621 763 657
rect -530 -630 763 -621
<< nwell >>
rect 0 8 128 292
<< pmos >>
rect 21 214 89 244
rect 21 83 89 113
<< pdiff >>
rect 21 268 89 273
rect 21 250 28 268
rect 46 250 64 268
rect 82 250 89 268
rect 21 244 89 250
rect 21 208 89 214
rect 21 190 29 208
rect 46 190 65 208
rect 83 190 89 208
rect 21 184 89 190
rect 21 137 89 143
rect 21 120 29 137
rect 47 120 65 137
rect 83 120 89 137
rect 21 113 89 120
rect 21 76 89 83
rect 21 59 29 76
rect 47 59 65 76
rect 83 59 89 76
rect 21 55 89 59
<< pdiffc >>
rect 28 250 46 268
rect 64 250 82 268
rect 29 190 46 208
rect 65 190 83 208
rect 29 120 47 137
rect 65 120 83 137
rect 29 59 47 76
rect 65 59 83 76
<< nsubdiff >>
rect 21 172 89 184
rect 21 155 29 172
rect 47 155 65 172
rect 83 155 89 172
rect 21 143 89 155
<< nsubdiffcont >>
rect 29 155 47 172
rect 65 155 83 172
<< poly >>
rect 8 214 21 244
rect 89 214 114 244
rect 97 113 114 214
rect 8 83 21 113
rect 89 83 114 113
rect 97 31 114 83
<< locali >>
rect 20 250 28 268
rect 46 250 64 268
rect 82 250 90 268
rect 21 190 29 208
rect 46 190 65 208
rect 83 190 91 208
rect 21 172 91 190
rect 21 155 29 172
rect 47 155 65 172
rect 83 155 91 172
rect 21 137 91 155
rect 21 120 29 137
rect 47 120 65 137
rect 83 120 91 137
rect 21 59 29 76
rect 47 59 65 76
rect 83 59 92 76
rect 56 31 92 59
rect 56 14 89 31
use sky130_hilas_poly2li  sky130_hilas_poly2li_0
timestamp 1628707323
transform 0 1 100 -1 0 27
box 0 0 27 33
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
