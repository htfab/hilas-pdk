magic
tech sky130A
timestamp 1634057780
<< nwell >>
rect 0 139 969 599
rect 0 0 1029 139
<< mvvaractor >>
rect 56 74 912 540
<< mvnsubdiff >>
rect 56 540 912 566
rect 960 89 996 106
rect 56 50 912 74
rect 960 72 966 89
rect 983 72 996 89
rect 960 55 996 72
rect 960 50 966 55
rect 56 38 966 50
rect 983 38 996 55
rect 56 33 996 38
<< mvnsubdiffcont >>
rect 966 72 983 89
rect 966 38 983 55
<< poly >>
rect 16 74 56 540
rect 912 74 951 540
<< locali >>
rect 966 89 983 97
rect 966 30 983 38
<< viali >>
rect 966 55 983 72
<< metal1 >>
rect 963 72 987 82
rect 963 55 966 72
rect 983 55 987 72
rect 963 46 987 55
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
