magic
tech sky130A
timestamp 1627737364
<< error_s >>
rect 489 970 506 972
rect 489 951 506 953
rect 154 503 158 537
rect 154 455 159 503
<< nwell >>
rect 145 728 213 729
rect 145 725 221 728
rect 428 725 429 729
rect 466 437 528 1007
<< nsubdiff >>
rect 484 970 510 989
rect 484 953 489 970
rect 506 953 510 970
rect 484 936 510 953
rect 484 919 489 936
rect 506 919 510 936
rect 484 907 510 919
<< nsubdiffcont >>
rect 489 953 506 970
rect 489 919 506 936
<< poly >>
rect 126 1001 429 1018
rect 126 729 145 1001
rect 126 714 429 729
rect 126 523 146 714
rect 78 513 146 523
rect 78 496 83 513
rect 100 496 117 513
rect 134 496 146 513
rect 78 479 146 496
rect 78 462 84 479
rect 101 462 118 479
rect 135 462 146 479
rect 78 447 146 462
rect 78 445 428 447
rect 78 428 84 445
rect 101 428 118 445
rect 135 430 428 445
rect 135 428 161 430
rect 78 423 161 428
rect 78 420 147 423
<< polycont >>
rect 83 496 100 513
rect 117 496 134 513
rect 84 462 101 479
rect 118 462 135 479
rect 84 428 101 445
rect 118 428 135 445
<< locali >>
rect 489 911 506 919
rect 160 735 176 738
rect 160 701 177 735
rect 215 734 231 738
rect 215 701 232 734
rect 270 701 287 741
rect 325 734 341 738
rect 380 734 396 738
rect 435 736 451 738
rect 325 701 342 734
rect 380 701 397 734
rect 435 701 452 736
rect 160 700 176 701
rect 215 700 231 701
rect 270 700 286 701
rect 325 700 341 701
rect 380 700 396 701
rect 435 700 451 701
rect 83 513 134 521
rect 100 496 117 513
rect 83 495 134 496
rect 83 488 135 495
rect 84 479 135 488
rect 101 462 118 479
rect 84 445 135 462
rect 101 428 118 445
rect 84 420 135 428
<< viali >>
rect 489 970 506 987
rect 489 936 506 953
<< metal1 >>
rect 478 998 504 1018
rect 478 987 509 998
rect 478 970 489 987
rect 506 970 509 987
rect 478 953 509 970
rect 478 936 489 953
rect 506 936 509 953
rect 478 917 509 936
rect 478 419 504 917
<< metal2 >>
rect 97 979 403 980
rect 88 946 403 979
rect 88 701 120 946
rect 207 878 501 908
rect 426 874 501 878
rect 463 861 501 874
rect 466 774 501 861
rect 206 741 501 774
rect 88 668 404 701
rect 88 564 120 668
rect 88 532 404 564
rect 64 420 124 502
rect 466 497 501 741
rect 207 465 501 497
rect 207 464 478 465
use sky130_hilas_li2m2  sky130_hilas_li2m2_10
timestamp 1627737364
transform 1 0 274 0 1 546
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_6
timestamp 1627737364
transform 1 0 384 0 1 546
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_15
timestamp 1627737364
transform 1 0 220 0 1 478
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_17
timestamp 1627737364
transform 1 0 329 0 1 478
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_19
timestamp 1627737364
transform 1 0 439 0 1 479
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_9
timestamp 1627737364
transform 1 0 164 0 1 546
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_7
timestamp 1627737364
transform 1 0 108 0 1 435
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_8
timestamp 1627737364
transform 1 0 107 0 1 482
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1627737364
transform 1 0 274 0 1 683
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1627737364
transform 1 0 384 0 1 683
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1627737364
transform 1 0 164 0 1 683
box -14 -15 20 18
use sky130_hilas_pFETLargePart1  sky130_hilas_pFETLargePart1_1
timestamp 1627737364
transform 1 0 142 0 1 446
box -6 -9 333 278
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1627737364
transform 1 0 329 0 1 756
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_4
timestamp 1627737364
transform 1 0 220 0 1 756
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_5
timestamp 1627737364
transform 1 0 439 0 1 756
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_14
timestamp 1627737364
transform 1 0 274 0 1 961
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_18
timestamp 1627737364
transform 1 0 384 0 1 960
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_11
timestamp 1627737364
transform 1 0 165 0 1 961
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_16
timestamp 1627737364
transform 1 0 220 0 1 893
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_12
timestamp 1627737364
transform 1 0 329 0 1 891
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_13
timestamp 1627737364
transform 1 0 440 0 1 890
box -14 -15 20 18
use sky130_hilas_pFETLargePart1  sky130_hilas_pFETLargePart1_0
timestamp 1627737364
transform 1 0 142 0 1 729
box -6 -9 333 278
<< labels >>
rlabel metal2 486 834 500 908 0 DRAIN
port 3 nsew analog default
rlabel metal2 88 905 102 979 0 SOURCE
port 2 nsew analog default
rlabel metal2 64 420 74 502 0 GATE
port 1 nsew
rlabel metal1 478 1010 504 1018 0 WELL
port 4 nsew analog default
rlabel metal1 478 419 504 427 0 WELL
port 4 nsew analog default
<< end >>
