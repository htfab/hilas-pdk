magic
tech sky130A
timestamp 1607257541
<< error_p >>
rect -237 109 -208 137
rect -158 109 -129 137
rect -79 109 -50 137
rect -259 102 -29 109
rect -259 87 -252 102
rect -237 96 -208 102
rect -158 96 -129 102
rect -79 96 -50 102
rect -237 87 -236 88
rect -209 87 -208 88
rect -158 87 -157 88
rect -130 87 -129 88
rect -79 87 -78 88
rect -51 87 -50 88
rect -36 87 -29 102
rect -287 58 -246 87
rect -238 86 -207 87
rect -159 86 -128 87
rect -80 86 -49 87
rect -237 59 -208 86
rect -158 59 -129 86
rect -79 59 -50 86
rect -238 58 -207 59
rect -159 58 -128 59
rect -80 58 -49 59
rect -42 58 0 87
rect -259 8 -252 58
rect -237 57 -236 58
rect -209 57 -208 58
rect -158 57 -157 58
rect -130 57 -129 58
rect -79 57 -78 58
rect -51 57 -50 58
rect -237 8 -236 9
rect -209 8 -208 9
rect -158 8 -157 9
rect -130 8 -129 9
rect -79 8 -78 9
rect -51 8 -50 9
rect -36 8 -29 58
rect -287 -21 -246 8
rect -238 7 -207 8
rect -159 7 -128 8
rect -80 7 -49 8
rect -237 -20 -208 7
rect -158 -20 -129 7
rect -79 -20 -50 7
rect -238 -21 -207 -20
rect -159 -21 -128 -20
rect -80 -21 -49 -20
rect -42 -21 0 8
rect -259 -36 -252 -21
rect -237 -22 -236 -21
rect -209 -22 -208 -21
rect -158 -22 -157 -21
rect -130 -22 -129 -21
rect -79 -22 -78 -21
rect -51 -22 -50 -21
rect -237 -36 -208 -30
rect -158 -36 -129 -30
rect -79 -36 -50 -30
rect -36 -36 -29 -21
rect -259 -43 -29 -36
rect -237 -71 -208 -43
rect -158 -71 -129 -43
rect -79 -71 -50 -43
<< nwell >>
rect -281 -65 -9 131
<< mvpmos >>
rect -246 87 -42 96
rect -246 58 -237 87
rect -208 58 -158 87
rect -129 58 -79 87
rect -50 58 -42 87
rect -246 8 -42 58
rect -246 -21 -237 8
rect -208 -21 -158 8
rect -129 -21 -79 8
rect -50 -21 -42 8
rect -246 -30 -42 -21
<< mvpdiff >>
rect -237 81 -208 87
rect -237 64 -231 81
rect -214 64 -208 81
rect -237 58 -208 64
rect -158 81 -129 87
rect -158 64 -152 81
rect -135 64 -129 81
rect -158 58 -129 64
rect -79 81 -50 87
rect -79 64 -73 81
rect -56 64 -50 81
rect -79 58 -50 64
rect -237 1 -208 8
rect -237 -15 -231 1
rect -214 -15 -208 1
rect -237 -21 -208 -15
rect -158 1 -129 8
rect -158 -15 -152 1
rect -135 -15 -129 1
rect -158 -21 -129 -15
rect -79 2 -50 8
rect -79 -15 -73 2
rect -56 -15 -50 2
rect -79 -21 -50 -15
<< mvpdiffc >>
rect -231 64 -214 81
rect -152 64 -135 81
rect -73 64 -56 81
rect -231 -15 -214 1
rect -152 -15 -135 1
rect -73 -15 -56 2
<< poly >>
rect -252 96 -36 102
rect -252 -30 -246 96
rect -42 -30 -36 96
rect -252 -36 -36 -30
<< locali >>
rect -241 81 -46 91
rect -241 64 -231 81
rect -214 74 -152 81
rect -214 64 -193 74
rect -241 57 -193 64
rect -176 64 -152 74
rect -135 64 -73 81
rect -56 64 -46 81
rect -176 57 -46 64
rect -241 40 -46 57
rect -241 23 -193 40
rect -176 23 -46 40
rect -241 6 -46 23
rect -241 1 -193 6
rect -241 -15 -231 1
rect -214 -11 -193 1
rect -176 2 -46 6
rect -176 1 -73 2
rect -176 -11 -152 1
rect -214 -15 -152 -11
rect -135 -15 -73 1
rect -56 -15 -46 2
rect -241 -26 -46 -15
<< viali >>
rect -193 57 -176 74
rect -193 23 -176 40
rect -193 -11 -176 6
<< metal1 >>
rect -197 74 -171 80
rect -197 57 -193 74
rect -176 57 -171 74
rect -197 40 -171 57
rect -197 32 -193 40
rect -198 23 -193 32
rect -176 23 -171 40
rect -198 6 -171 23
rect -198 -11 -193 6
rect -176 -11 -171 6
rect -198 -20 -171 -11
rect -198 -65 -172 -20
<< end >>
