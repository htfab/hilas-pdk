magic
tech sky130A
timestamp 1607993916
<< error_s >>
rect -401 342 -395 348
rect -296 342 -290 348
rect -407 278 -401 284
rect -290 278 -284 284
rect -457 219 -234 220
rect -31 195 44 213
rect -31 131 -13 195
rect 26 131 44 195
rect -31 113 44 131
rect -36 64 59 82
rect -374 20 -368 26
rect -321 20 -315 26
rect -8 -18 -7 64
rect 25 47 59 64
rect -3 39 25 47
rect -3 28 38 39
rect -3 -18 19 28
rect 25 10 59 28
rect 68 21 74 27
rect 173 21 179 27
rect 20 -18 59 10
rect -8 -19 59 -18
rect -380 -30 -374 -24
rect -315 -30 -309 -24
rect 62 -29 68 -23
rect 179 -29 185 -23
<< nmos >>
rect -8 10 25 39
<< ndiff >>
rect -8 39 25 64
rect -8 4 25 10
rect -8 -13 0 4
rect 17 -13 25 4
rect -8 -19 25 -13
<< pdiff >>
rect -13 131 26 195
<< ndiffc >>
rect 0 -13 17 4
<< poly >>
rect -21 10 -8 39
rect 25 10 38 39
<< locali >>
rect -8 -13 0 4
rect 17 -13 25 4
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_0
timestamp 1607993916
transform 1 0 1020 0 1 303
box -1451 -400 -784 -210
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_0
timestamp 1607386385
transform 1 0 530 0 1 165
box -289 47 -33 232
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_0
timestamp 1606741561
transform 1 0 500 0 1 614
box -957 -395 -734 -209
<< end >>
