magic
tech sky130A
timestamp 1607480432
use sky130_hilas_pFETdevice01a  sky130_hilas_pFETdevice01a_0
timestamp 1607477942
transform 1 0 108 0 1 -132
box -80 -42 81 43
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_0
timestamp 1607471549
transform 1 0 107 0 1 -36
box -79 -78 82 43
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_4
timestamp 1607471549
transform 1 0 107 0 1 60
box -79 -78 82 43
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_3
timestamp 1607471549
transform 1 0 107 0 1 156
box -79 -78 82 43
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_6
timestamp 1607471549
transform 1 0 107 0 1 252
box -79 -78 82 43
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_0
timestamp 1607478455
transform 1 0 108 0 1 348
box -80 -78 92 43
<< end >>
