magic
tech sky130A
timestamp 1625321931
<< nwell >>
rect 663 213 744 505
<< psubdiff >>
rect 670 619 714 643
rect 670 602 683 619
rect 700 602 714 619
rect 670 585 714 602
rect 670 568 683 585
rect 700 568 714 585
rect 670 551 714 568
rect 670 534 683 551
rect 700 534 714 551
rect 670 525 714 534
rect 671 161 714 187
rect 671 144 684 161
rect 701 144 714 161
rect 671 127 714 144
rect 671 110 684 127
rect 701 110 714 127
rect 671 93 714 110
rect 671 76 684 93
rect 701 76 714 93
rect 671 71 714 76
<< nsubdiff >>
rect 671 462 713 474
rect 671 444 682 462
rect 700 444 713 462
rect 671 425 713 444
rect 671 407 682 425
rect 700 407 713 425
rect 671 389 713 407
rect 671 371 682 389
rect 700 371 713 389
rect 671 353 713 371
rect 671 335 682 353
rect 700 335 713 353
rect 671 318 713 335
rect 671 300 683 318
rect 701 300 713 318
rect 671 282 713 300
rect 671 264 683 282
rect 701 264 713 282
rect 671 255 713 264
<< psubdiffcont >>
rect 683 602 700 619
rect 683 568 700 585
rect 683 534 700 551
rect 684 144 701 161
rect 684 110 701 127
rect 684 76 701 93
<< nsubdiffcont >>
rect 682 444 700 462
rect 682 407 700 425
rect 682 371 700 389
rect 682 335 700 353
rect 683 300 701 318
rect 683 264 701 282
<< locali >>
rect 646 619 708 636
rect 646 602 683 619
rect 700 602 708 619
rect 646 585 708 602
rect 646 568 683 585
rect 700 568 708 585
rect 646 551 708 568
rect 646 547 683 551
rect 672 534 683 547
rect 700 534 708 551
rect 672 532 708 534
rect 644 462 702 470
rect 644 444 682 462
rect 700 444 702 462
rect 644 431 702 444
rect 644 425 707 431
rect 644 407 682 425
rect 700 407 707 425
rect 644 389 707 407
rect 644 385 682 389
rect 644 368 647 385
rect 664 368 681 385
rect 700 371 707 389
rect 698 368 707 371
rect 644 353 707 368
rect 644 350 682 353
rect 644 333 647 350
rect 664 333 681 350
rect 700 335 707 353
rect 698 333 707 335
rect 644 318 707 333
rect 644 300 683 318
rect 701 300 707 318
rect 644 293 707 300
rect 644 282 702 293
rect 644 264 683 282
rect 701 264 702 282
rect 644 256 702 264
rect 646 161 701 171
rect 646 144 684 161
rect 646 127 701 144
rect 646 110 684 127
rect 646 93 701 110
rect 646 82 684 93
rect 684 68 701 76
<< viali >>
rect 647 368 664 385
rect 681 371 682 385
rect 682 371 698 385
rect 681 368 698 371
rect 647 333 664 350
rect 681 335 682 350
rect 682 335 698 350
rect 681 333 698 335
<< metal1 >>
rect 355 598 376 661
rect 637 598 744 661
rect 355 530 744 598
rect 355 385 744 499
rect 355 379 647 385
rect 355 314 372 379
rect 607 368 647 379
rect 664 368 681 385
rect 698 368 744 385
rect 607 350 744 368
rect 607 333 647 350
rect 664 333 681 350
rect 698 333 744 350
rect 607 314 744 333
rect 355 220 744 314
rect 355 60 744 184
rect 355 57 372 60
rect 646 58 744 60
rect 645 57 744 58
use sky130_hilas_decoup_cap_00  CapDeco_0
timestamp 1623107852
transform 1 0 273 0 -1 548
box 82 -113 390 189
use sky130_hilas_decoup_cap_00  CapDeco_1
timestamp 1623107852
transform 1 0 273 0 1 170
box 82 -113 390 189
<< labels >>
rlabel metal1 355 311 372 407 0 VPWR
rlabel metal1 727 313 744 407 0 VPWR
rlabel metal1 734 598 744 661 0 VPWR
rlabel metal1 355 598 363 661 0 VPWR
rlabel metal1 355 57 364 120 0 VPWR
rlabel metal1 729 57 744 120 0 VPWR
<< end >>
