* Copyright 2020 The Hilas PDK Authors
* 
* This file is part of HILAS.
* 
* HILAS is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published by
* the Free Software Foundation, version 3 of the License.
* 
* HILAS is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
* 
* You should have received a copy of the GNU Lesser General Public License
* along with HILAS.  If not, see <https://www.gnu.org/licenses/>.
* 
* Licensed under the Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
* https://www.gnu.org/licenses/lgpl-3.0.en.html
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
* SPDX-License-Identifier: LGPL-3.0
* 
* 

* NGSPICE file created from sky130_hilas_WTAblockSample01.ext - technology: sky130A

.subckt sky130_hilas_TunCap01 $SUB a_n2872_n666# w_n2902_n800#
X0 a_n2872_n666# w_n2902_n800# w_n2902_n800# sky130_fd_pr__cap_var w=590000u l=500000u
.ends

.subckt sky130_hilas_horizPcell01 a_n502_286# a_n508_162# w_n578_94# $SUB a_n578_238#
+ m1_n258_94# a_n300_94# a_n344_286#
X0 w_n578_94# a_n300_94# a_n344_162# w_n578_94# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
X1 a_n344_286# a_n578_238# a_n502_286# w_n578_94# sky130_fd_pr__pfet_g5v0d10v5 w=300000u l=500000u
X2 a_n344_162# a_n578_238# a_n508_162# w_n578_94# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
.ends

.subckt sky130_hilas_FGVaractorCapacitor m1_n1784_n790# $SUB a_n1882_n672# w_n1914_n790#
X0 a_n1882_n672# w_n1914_n790# w_n1914_n790# sky130_fd_pr__cap_var w=1.11e+06u l=640000u
.ends

.subckt sky130_hilas_cellAttempt01 m1_n456_n764# a_1264_n176# m2_n524_n660# m2_n524_n572#
+ m2_n528_n62# sky130_hilas_wellContact_0/w_n2898_n880# sky130_hilas_horizPcell01_3/a_n344_286#
+ m2_n524_n376# $SUB m2_n524_n292# w_1264_n176# m2_n528_24# m2_n528_310# m2_n528_224#
Xsky130_hilas_TunCap01_0 $SUB a_640_n334# m1_n456_n764# sky130_hilas_TunCap01
Xsky130_hilas_TunCap01_1 $SUB a_640_n618# m1_n456_n764# sky130_hilas_TunCap01
Xsky130_hilas_TunCap01_2 $SUB a_n214_10# m1_n456_n764# sky130_hilas_TunCap01
Xsky130_hilas_TunCap01_3 $SUB a_638_270# m1_n456_n764# sky130_hilas_TunCap01
Xsky130_hilas_horizPcell01_0 m2_n528_24# m2_n528_n62# w_1264_n176# $SUB a_n214_10#
+ a_1264_n176# a_1264_n176# sky130_hilas_horizPcell01_3/a_n344_286# sky130_hilas_horizPcell01
Xsky130_hilas_horizPcell01_1 m2_n524_n572# m2_n524_n660# w_1264_n176# $SUB a_640_n618#
+ a_1264_n176# a_1264_n176# sky130_hilas_horizPcell01_3/a_n344_286# sky130_hilas_horizPcell01
Xsky130_hilas_horizPcell01_2 m2_n524_n376# m2_n524_n292# w_1264_n176# $SUB a_640_n334#
+ a_1264_n176# a_1264_n176# sky130_hilas_horizPcell01_3/a_n344_286# sky130_hilas_horizPcell01
Xsky130_hilas_horizPcell01_3 m2_n528_224# m2_n528_310# w_1264_n176# $SUB a_638_270#
+ a_1264_n176# a_1264_n176# sky130_hilas_horizPcell01_3/a_n344_286# sky130_hilas_horizPcell01
Xsky130_hilas_FGVaractorCapacitor_0 sky130_hilas_wellContact_0/w_n2898_n880# $SUB
+ a_640_n618# sky130_hilas_wellContact_0/w_n2898_n880# sky130_hilas_FGVaractorCapacitor
Xsky130_hilas_FGVaractorCapacitor_2 sky130_hilas_wellContact_0/w_n2898_n880# $SUB
+ a_n214_10# sky130_hilas_wellContact_0/w_n2898_n880# sky130_hilas_FGVaractorCapacitor
Xsky130_hilas_FGVaractorCapacitor_1 sky130_hilas_wellContact_0/w_n2898_n880# $SUB
+ a_640_n334# sky130_hilas_wellContact_0/w_n2898_n880# sky130_hilas_FGVaractorCapacitor
Xsky130_hilas_FGVaractorCapacitor_3 sky130_hilas_wellContact_0/w_n2898_n880# $SUB
+ a_638_270# sky130_hilas_wellContact_0/w_n2898_n880# sky130_hilas_FGVaractorCapacitor
.ends

.subckt sky130_hilas_swc4x2cell GATE2 VTUN GATE1 VPWR GATESELECT1 SelectGate2 VERT1
+ VERT2 HORIZ1 HORIZ2 DRAIN1 DRAIN4 DRAIN3 HORIZ3 HORIZ4 $SUB
Xsky130_hilas_cellAttempt01_0 VTUN SelectGate2 DRAIN4 HORIZ4 DRAIN4 GATE2 VERT2 HORIZ3
+ $SUB DRAIN3 VPWR HORIZ2 DRAIN1 HORIZ1 sky130_hilas_cellAttempt01
Xsky130_hilas_cellAttempt01_1 VTUN GATESELECT1 DRAIN4 HORIZ4 DRAIN4 GATE1 VERT1 HORIZ3
+ $SUB DRAIN3 VPWR HORIZ2 DRAIN1 HORIZ1 sky130_hilas_cellAttempt01
.ends

.subckt sky130_hilas_WTAsinglestage01 a_4_n68# a_216_n68# $SUB
X0 a_4_n68# a_n126_n150# a_n94_n68# $SUB sky130_fd_pr__nfet_01v8 w=590000u l=200000u
X1 $SUB a_4_n68# a_n126_n150# $SUB sky130_fd_pr__nfet_01v8 w=590000u l=200000u
.ends

.subckt sky130_hilas_WTA4stage01 $SUB
Xsky130_hilas_WTAsinglestage01_0 a_284_2# m1_380_516# $SUB sky130_hilas_WTAsinglestage01
Xsky130_hilas_WTAsinglestage01_1 a_284_2# m1_380_516# $SUB sky130_hilas_WTAsinglestage01
Xsky130_hilas_WTAsinglestage01_2 a_284_2# m1_380_516# $SUB sky130_hilas_WTAsinglestage01
Xsky130_hilas_WTAsinglestage01_3 a_284_2# m1_380_516# $SUB sky130_hilas_WTAsinglestage01
.ends


* Top level circuit sky130_hilas_WTAblockSample01

Xsky130_hilas_swc4x2cell_0 sky130_hilas_swc4x2cell_1/GATE2 sky130_hilas_swc4x2cell_1/VTUN
+ sky130_hilas_swc4x2cell_1/GATE1 sky130_hilas_swc4x2cell_1/VPWR sky130_hilas_swc4x2cell_1/GATESELECT1
+ sky130_hilas_swc4x2cell_1/SelectGate2 sky130_hilas_swc4x2cell_1/VERT1 sky130_hilas_swc4x2cell_1/VERT2
+ sky130_hilas_swc4x2cell_0/HORIZ1 sky130_hilas_swc4x2cell_0/HORIZ2 sky130_hilas_swc4x2cell_0/DRAIN1
+ sky130_hilas_swc4x2cell_0/DRAIN4 sky130_hilas_swc4x2cell_0/DRAIN3 sky130_hilas_swc4x2cell_0/HORIZ3
+ sky130_hilas_swc4x2cell_0/HORIZ4 $SUB sky130_hilas_swc4x2cell
Xsky130_hilas_swc4x2cell_1 sky130_hilas_swc4x2cell_1/GATE2 sky130_hilas_swc4x2cell_1/VTUN
+ sky130_hilas_swc4x2cell_1/GATE1 sky130_hilas_swc4x2cell_1/VPWR sky130_hilas_swc4x2cell_1/GATESELECT1
+ sky130_hilas_swc4x2cell_1/SelectGate2 sky130_hilas_swc4x2cell_1/VERT1 sky130_hilas_swc4x2cell_1/VERT2
+ sky130_hilas_swc4x2cell_1/HORIZ1 sky130_hilas_swc4x2cell_1/HORIZ2 sky130_hilas_swc4x2cell_1/DRAIN1
+ sky130_hilas_swc4x2cell_1/DRAIN4 sky130_hilas_swc4x2cell_1/DRAIN3 sky130_hilas_swc4x2cell_1/HORIZ3
+ sky130_hilas_swc4x2cell_1/HORIZ4 $SUB sky130_hilas_swc4x2cell
Xsky130_hilas_WTA4stage01_0 $SUB sky130_hilas_WTA4stage01
Xsky130_hilas_WTA4stage01_1 $SUB sky130_hilas_WTA4stage01
.end

