magic
tech sky130A
timestamp 1629137229
<< checkpaint >>
rect -612 -512 820 1253
rect -612 -608 809 -512
<< error_s >>
rect 0 522 39 525
rect 0 480 39 483
rect 0 426 39 429
rect 0 384 39 387
rect 0 330 39 333
rect 0 288 39 291
rect 0 234 39 237
rect 0 192 39 195
rect 0 138 39 141
rect 0 96 39 99
rect 0 42 39 45
rect 0 0 39 3
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_3
timestamp 1629137127
transform 1 0 18 0 1 502
box 0 0 172 121
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_2
timestamp 1629137127
transform 1 0 18 0 1 406
box 0 0 172 121
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_4
timestamp 1629137127
transform 1 0 18 0 1 310
box 0 0 172 121
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_1
timestamp 1629137127
transform 1 0 18 0 1 214
box 0 0 172 121
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_0
timestamp 1629137127
transform 1 0 18 0 1 118
box 0 0 172 121
use sky130_hilas_pFETdevice01a  sky130_hilas_pFETdevice01a_0
timestamp 1629137174
transform 1 0 18 0 1 22
box 0 0 161 85
<< end >>
