magic
tech sky130A
timestamp 1623423324
<< metal1 >>
rect 1108 604 1133 610
rect 1407 605 1430 610
rect 1542 605 1561 610
<< metal2 >>
rect 1107 559 1180 560
rect 1107 543 1249 559
rect 1107 542 1180 543
rect 1107 372 1174 374
rect 1107 356 1246 372
rect 1107 257 1177 258
rect 1107 241 1250 257
rect 1107 57 1253 74
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_2
timestamp 1607907894
transform 1 0 1282 0 1 45
box -210 -40 332 119
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_1
timestamp 1607907894
transform 1 0 1282 0 -1 570
box -210 -40 332 119
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_3
timestamp 1607907894
transform 1 0 1282 0 -1 277
box -210 -40 332 119
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_0
timestamp 1607907894
transform 1 0 1282 0 1 338
box -210 -40 332 119
<< labels >>
rlabel metal2 1107 542 1112 560 0 drain1
rlabel metal2 1107 356 1112 374 0 drain2
rlabel metal2 1107 241 1112 258 0 drain3
rlabel metal2 1107 57 1112 74 0 drain4
rlabel metal1 1108 604 1133 610 0 Vinj
port 1 nsew
rlabel metal1 1407 605 1430 610 0 SelectDrain
port 2 nsew
rlabel metal1 1542 605 1561 610 0 GND
port 3 nsew
<< end >>
