magic
tech sky130A
timestamp 1634057762
<< checkpaint >>
rect -607 -548 687 745
<< nwell >>
rect 0 0 256 191
<< mvpmos >>
rect 67 85 117 139
<< mvpdiff >>
rect 38 133 67 139
rect 38 91 42 133
rect 60 91 67 133
rect 38 85 67 91
rect 117 128 146 139
rect 117 111 123 128
rect 142 111 146 128
rect 117 85 146 111
<< mvpdiffc >>
rect 42 91 60 133
rect 123 111 142 128
<< mvnsubdiff >>
rect 189 128 223 142
rect 189 110 196 128
rect 216 110 223 128
rect 189 98 223 110
<< mvnsubdiffcont >>
rect 196 110 216 128
<< poly >>
rect 67 139 117 152
rect 67 76 117 85
rect 0 59 117 76
<< locali >>
rect 34 133 68 135
rect 34 91 42 133
rect 60 91 68 133
rect 123 128 143 136
rect 142 111 143 128
rect 123 97 143 111
rect 123 80 124 97
rect 141 80 143 97
rect 123 76 143 80
rect 195 128 217 136
rect 195 110 196 128
rect 216 110 217 128
rect 195 94 217 110
rect 195 77 197 94
rect 214 77 217 94
rect 196 74 217 77
rect 196 70 216 74
<< viali >>
rect 124 80 141 97
rect 197 77 214 94
<< metal1 >>
rect 123 105 139 191
rect 204 140 220 191
rect 204 131 221 140
rect 193 126 221 131
rect 123 100 144 105
rect 121 97 144 100
rect 121 80 124 97
rect 141 80 144 97
rect 121 76 144 80
rect 193 94 220 126
rect 193 77 197 94
rect 214 77 220 94
rect 123 74 143 76
rect 123 1 139 74
rect 193 71 220 77
rect 204 1 220 71
<< metal2 >>
rect 0 99 9 117
rect 39 99 256 117
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1634057699
transform 1 0 23 0 -1 115
box 0 0 34 33
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
