VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_swc4x2cellOverlap
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc4x2cellOverlap ;
  ORIGIN 10.010 -7.280 ;
  SIZE 17.980 BY 6.050 ;
  PIN Vert1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT -8.840 12.590 -8.680 13.330 ;
    END
    PORT
      LAYER met1 ;
        RECT -8.840 7.290 -8.680 8.030 ;
    END
  END Vert1
  PIN Horiz1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -10.010 12.220 -7.830 12.400 ;
    END
    PORT
      LAYER met2 ;
        RECT 5.780 12.220 7.970 12.400 ;
    END
  END Horiz1
  PIN drain1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -10.010 12.650 -7.830 12.830 ;
    END
    PORT
      LAYER met2 ;
        RECT 5.780 12.650 7.960 12.830 ;
    END
  END drain1
  PIN Horiz2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -10.010 11.220 -7.830 11.400 ;
    END
    PORT
      LAYER met2 ;
        RECT 5.780 11.220 7.970 11.400 ;
    END
  END Horiz2
  PIN drain2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -10.010 10.790 -7.830 10.970 ;
    END
    PORT
      LAYER met2 ;
        RECT 5.780 10.790 7.970 10.970 ;
    END
  END drain2
  PIN drain3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -10.010 9.640 -7.830 9.820 ;
    END
    PORT
      LAYER met2 ;
        RECT 5.780 9.640 7.960 9.820 ;
    END
  END drain3
  PIN Horiz3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -10.010 9.210 -7.830 9.390 ;
    END
    PORT
      LAYER met2 ;
        RECT 5.780 9.210 7.960 9.390 ;
    END
  END Horiz3
  PIN Horiz4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -10.010 8.220 -7.830 8.400 ;
    END
    PORT
      LAYER met2 ;
        RECT 5.780 8.220 7.960 8.400 ;
    END
  END Horiz4
  PIN drain4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -10.010 7.790 -7.830 7.970 ;
    END
  END drain4
  PIN Vinj
    PORT
      LAYER met1 ;
        RECT -9.650 12.620 -9.490 13.330 ;
    END
    PORT
      LAYER met1 ;
        RECT -9.650 7.290 -9.490 8.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 7.440 7.290 7.600 8.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 7.440 12.620 7.600 13.330 ;
    END
  END Vinj
  PIN GateSelect1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT -9.240 12.340 -9.050 13.330 ;
    END
    PORT
      LAYER met1 ;
        RECT -9.240 7.290 -9.050 8.280 ;
    END
  END GateSelect1
  PIN Vert2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 6.630 12.590 6.790 13.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.630 7.290 6.790 8.030 ;
    END
  END Vert2
  PIN GateSelect2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 7.000 12.340 7.190 13.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 7.000 7.290 7.190 8.280 ;
    END
  END GateSelect2
  PIN drain
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.780 7.790 7.960 7.970 ;
    END
  END drain
  PIN Gate2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 3.280 12.940 3.520 13.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.280 7.280 3.520 7.670 ;
    END
  END Gate2
  PIN Gate1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT -5.570 12.940 -5.320 13.330 ;
    END
    PORT
      LAYER met1 ;
        RECT -5.570 7.280 -5.320 7.670 ;
    END
  END Gate1
  PIN Vtun
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT -1.960 12.980 -1.660 13.330 ;
    END
    PORT
      LAYER met1 ;
        RECT -1.960 7.280 -1.660 7.610 ;
    END
    PORT
      LAYER met1 ;
        RECT -0.380 7.280 -0.080 7.610 ;
    END
  END Vtun
  OBS
      LAYER li1 ;
        RECT -9.620 7.610 7.570 13.010 ;
      LAYER met1 ;
        RECT -8.400 12.660 -5.850 13.330 ;
        RECT -5.040 12.700 -2.240 13.330 ;
        RECT -1.380 12.700 3.000 13.330 ;
        RECT -5.040 12.660 3.000 12.700 ;
        RECT 3.800 12.660 6.350 13.330 ;
        RECT -9.660 12.060 -9.520 12.340 ;
        RECT -8.400 12.310 6.350 12.660 ;
        RECT -8.770 12.060 6.720 12.310 ;
        RECT 7.470 12.060 7.610 12.340 ;
        RECT -9.660 8.560 7.610 12.060 ;
        RECT -9.660 8.280 -9.520 8.560 ;
        RECT -8.770 8.310 6.720 8.560 ;
        RECT -8.400 7.950 6.350 8.310 ;
        RECT 7.470 8.280 7.610 8.560 ;
        RECT -8.400 7.470 -5.850 7.950 ;
        RECT -5.040 7.890 3.000 7.950 ;
        RECT -5.040 7.470 -2.240 7.890 ;
        RECT -1.380 7.470 -0.660 7.890 ;
        RECT 0.200 7.470 3.000 7.890 ;
        RECT 3.800 7.470 6.350 7.950 ;
      LAYER met2 ;
        RECT -7.550 11.940 5.500 12.970 ;
        RECT -7.850 11.680 5.800 11.940 ;
        RECT -7.550 10.510 5.500 11.680 ;
        RECT -7.850 10.100 5.800 10.510 ;
        RECT -7.550 8.930 5.500 10.100 ;
        RECT -7.850 8.680 5.800 8.930 ;
        RECT -7.550 7.650 5.500 8.680 ;
  END
END sky130_hilas_swc4x2cellOverlap
END LIBRARY

