magic
tech sky130A
timestamp 1608229393
<< metal1 >>
rect 1108 603 1133 610
rect 1407 603 1430 610
rect 1542 605 1561 610
rect 1607 498 1614 522
rect 1607 386 1614 410
rect 1608 205 1614 229
rect 1608 93 1614 117
rect 1407 5 1430 13
rect 1542 5 1561 12
<< metal2 >>
rect 1107 559 1180 560
rect 1107 543 1249 559
rect 1107 542 1180 543
rect 1107 372 1174 374
rect 1107 356 1246 372
rect 1107 257 1177 258
rect 1107 241 1250 257
rect 1107 57 1253 74
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_2
timestamp 1607907894
transform 1 0 1282 0 1 45
box -210 -40 332 119
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_1
timestamp 1607907894
transform 1 0 1282 0 -1 570
box -210 -40 332 119
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_3
timestamp 1607907894
transform 1 0 1282 0 -1 277
box -210 -40 332 119
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_0
timestamp 1607907894
transform 1 0 1282 0 1 338
box -210 -40 332 119
<< labels >>
rlabel metal2 1107 542 1112 560 0 DRAIN1
port 4 nsew analog default
rlabel metal2 1107 356 1112 374 0 DRAIN2
port 3 nsew analog default
rlabel metal2 1107 241 1112 258 0 DRAIN3
port 2 nsew
rlabel metal2 1107 57 1112 74 0 DRAIN4
port 1 nsew
rlabel metal1 1607 498 1614 522 0 DRAINSELECT1
port 5 nsew analog default
rlabel metal1 1607 386 1614 410 0 DRAINSELECT2
port 6 nsew analog default
rlabel metal1 1608 205 1614 229 0 DRAINSELECT3
port 7 nsew analog default
rlabel metal1 1608 93 1614 117 0 DRAINSELECT4
port 8 nsew analog default
rlabel metal1 1108 603 1133 610 0 VINJ
port 9 nsew power default
rlabel metal1 1407 603 1430 610 0 DRAIN_MUX
port 10 nsew analog default
rlabel metal1 1407 5 1430 13 0 DRAIN_MUX
port 10 nsew analog default
rlabel metal1 1542 5 1561 12 0 VGND
port 11 nsew ground default
rlabel metal1 1542 605 1561 610 0 VGND
port 11 nsew ground default
<< end >>
