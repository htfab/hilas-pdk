magic
tech sky130A
timestamp 1632489745
<< error_s >>
rect -87 540 -60 546
rect -87 498 -60 504
rect -87 473 -60 479
rect -87 431 -60 437
rect -87 390 -60 396
rect -87 348 -60 354
rect -87 323 -60 329
rect -87 281 -60 287
rect -87 240 -60 246
rect -87 198 -60 204
rect -87 173 -60 179
rect -87 131 -60 137
rect -87 90 -60 96
rect -87 48 -60 54
rect -87 23 -60 29
rect -87 -19 -60 -13
<< metal1 >>
rect -41 -22 -7 550
rect 26 -21 53 549
<< metal2 >>
rect -136 507 118 530
rect -110 293 155 316
rect -136 211 155 233
rect -137 -6 134 17
use sky130_hilas_pFETmirror02  sky130_hilas_pFETmirror02_0
timestamp 1632489745
transform 1 0 88 0 1 -111
box -61 89 67 373
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_1
timestamp 1632489745
transform 1 0 -113 0 1 130
box -59 -6 125 123
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_0
timestamp 1632489745
transform 1 0 -113 0 -1 97
box -59 -6 125 123
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1632488964
transform 1 0 41 0 1 126
box -10 -8 13 21
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1632488964
transform 1 0 106 0 1 228
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1632488964
transform 1 0 98 0 1 3
box -14 -15 20 18
use sky130_hilas_pFETmirror02  sky130_hilas_pFETmirror02_1
timestamp 1632489745
transform 1 0 88 0 -1 635
box -61 89 67 373
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_3
timestamp 1632489745
transform 1 0 -113 0 -1 397
box -59 -6 125 123
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_2
timestamp 1632489745
transform 1 0 -113 0 1 430
box -59 -6 125 123
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1632488964
transform 1 0 41 0 1 385
box -10 -8 13 21
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1632488964
transform 1 0 107 0 1 300
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1632488964
transform 1 0 102 0 1 522
box -14 -15 20 18
<< labels >>
rlabel metal2 144 293 155 316 0 output1
rlabel space 144 211 155 234 0 output2
<< end >>
