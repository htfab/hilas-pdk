VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_Trans4small
  CLASS BLOCK ;
  FOREIGN sky130_hilas_Trans4small ;
  ORIGIN -1.910 1.500 ;
  SIZE 2.800 BY 5.880 ;
  PIN nFET_Source1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 3.980 2.540 4.150 ;
    END
  END nFET_Source1
  PIN nFET_Gate1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 3.570 2.070 3.740 ;
    END
  END nFET_Gate1
  PIN nFET_Source2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 3.060 2.540 3.230 ;
    END
  END nFET_Source2
  PIN nFET_Gate2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 2.650 2.070 2.820 ;
    END
  END nFET_Gate2
  PIN nFET_Source3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 2.140 2.540 2.310 ;
    END
  END nFET_Source3
  PIN nFET_Gate3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 1.730 2.070 1.900 ;
    END
  END nFET_Gate3
  PIN pFET_Source1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 1.120 2.350 1.310 ;
    END
  END pFET_Source1
  PIN pFET_Gate1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 0.700 2.350 0.890 ;
    END
  END pFET_Gate1
  PIN pFET_Source2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 0.160 2.350 0.350 ;
    END
  END pFET_Source2
  PIN pFET_Gate2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 -0.260 2.350 -0.070 ;
    END
  END pFET_Gate2
  PIN pFET_Source3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 -0.800 2.350 -0.610 ;
    END
  END pFET_Source3
  PIN pFET_Gate3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 -1.220 2.350 -1.030 ;
    END
  END pFET_Gate3
  PIN Well
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 4.090 -1.500 4.310 -1.300 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.090 -1.130 4.310 4.380 ;
    END
  END Well
  PIN GND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 4.490 -1.500 4.710 3.520 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.490 3.690 4.710 4.380 ;
    END
  END GND
  PIN pFET_Drain3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 3.910 -0.870 4.710 -0.670 ;
    END
  END pFET_Drain3
  PIN pFET_Drain2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 3.910 0.090 4.710 0.290 ;
    END
  END pFET_Drain2
  PIN pFET_Drain1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 3.910 1.050 4.710 1.250 ;
    END
  END pFET_Drain1
  PIN nFET_Drain3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 3.890 2.150 4.710 2.320 ;
    END
  END nFET_Drain3
  PIN nFET_Drain2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 3.890 3.070 4.710 3.240 ;
    END
  END nFET_Drain2
  PIN nFET_Drain1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 3.890 3.990 4.710 4.160 ;
    END
  END nFET_Drain1
  OBS
      LAYER li1 ;
        RECT 2.080 -1.310 4.690 4.240 ;
      LAYER met1 ;
        RECT 2.040 -1.330 3.810 4.240 ;
      LAYER met2 ;
        RECT 2.820 3.710 3.610 4.250 ;
        RECT 2.820 3.700 3.930 3.710 ;
        RECT 2.350 3.520 3.930 3.700 ;
        RECT 2.350 3.510 3.610 3.520 ;
        RECT 2.820 2.790 3.610 3.510 ;
        RECT 2.820 2.780 3.930 2.790 ;
        RECT 2.350 2.600 3.930 2.780 ;
        RECT 2.350 2.590 3.610 2.600 ;
        RECT 2.820 1.870 3.610 2.590 ;
        RECT 2.820 1.860 3.930 1.870 ;
        RECT 2.350 1.590 3.930 1.860 ;
        RECT 2.630 1.530 3.930 1.590 ;
        RECT 2.630 0.770 3.630 1.530 ;
        RECT 2.630 0.570 3.930 0.770 ;
        RECT 2.630 -0.190 3.630 0.570 ;
        RECT 2.630 -0.390 3.930 -0.190 ;
        RECT 2.630 -1.150 3.630 -0.390 ;
        RECT 2.630 -1.290 3.930 -1.150 ;
  END
END sky130_hilas_Trans4small
END LIBRARY

