magic
tech sky130A
timestamp 1627063197
<< error_s >>
rect 434 542 440 548
rect 539 542 545 548
rect 60 532 66 538
rect 113 532 119 538
rect 54 482 60 488
rect 119 482 125 488
rect 428 478 434 484
rect 545 478 551 484
rect 60 423 66 429
rect 113 423 119 429
rect 434 425 440 431
rect 539 425 545 431
rect 54 373 60 379
rect 119 373 125 379
rect 428 361 434 367
rect 545 361 551 367
rect 434 240 440 246
rect 539 240 545 246
rect 60 234 66 240
rect 113 234 119 240
rect 265 235 282 239
rect 54 184 60 190
rect 119 184 125 190
rect 428 176 434 182
rect 545 176 551 182
rect 434 124 440 130
rect 539 124 545 130
rect 60 117 66 123
rect 113 117 119 123
rect 54 67 60 73
rect 119 67 125 73
rect 428 60 434 66
rect 545 60 551 66
<< nwell >>
rect 378 602 601 605
rect 2 419 3 542
rect 754 361 763 369
rect 898 310 933 311
rect 898 294 915 310
rect 932 294 933 310
rect 378 0 601 2
<< psubdiff >>
rect 260 464 285 487
rect 260 447 264 464
rect 281 447 285 464
rect 260 419 285 447
rect 662 461 687 489
rect 662 444 666 461
rect 683 444 687 461
rect 662 418 687 444
rect 260 337 286 379
rect 260 320 265 337
rect 282 320 286 337
rect 260 303 286 320
rect 260 286 265 303
rect 282 286 286 303
rect 260 269 286 286
rect 260 252 265 269
rect 282 252 286 269
rect 260 239 286 252
rect 662 343 689 364
rect 662 326 667 343
rect 684 326 689 343
rect 662 309 689 326
rect 662 292 667 309
rect 684 292 689 309
rect 662 275 689 292
rect 662 258 667 275
rect 684 258 689 275
rect 662 240 689 258
rect 265 235 282 239
<< psubdiffcont >>
rect 264 447 281 464
rect 666 444 683 461
rect 265 320 282 337
rect 265 286 282 303
rect 265 252 282 269
rect 667 326 684 343
rect 667 292 684 309
rect 667 258 684 275
<< poly >>
rect 585 529 755 533
rect 159 496 396 520
rect 585 517 754 529
rect 159 387 394 411
rect 585 373 754 390
rect 915 310 933 311
rect 931 294 933 310
rect 159 207 396 231
rect 586 215 754 232
rect 161 87 398 111
rect 586 73 754 90
<< polycont >>
rect 898 294 915 311
<< locali >>
rect 889 294 898 311
<< viali >>
rect 264 464 281 481
rect 264 430 281 447
rect 666 461 683 478
rect 666 427 683 444
rect 265 337 282 354
rect 265 303 282 320
rect 265 269 282 286
rect 265 235 282 252
rect 667 343 684 360
rect 667 309 684 326
rect 915 294 933 311
rect 667 275 684 292
rect 667 241 684 258
<< metal1 >>
rect 38 0 78 605
rect 259 481 286 605
rect 443 595 481 605
rect 259 464 264 481
rect 281 464 286 481
rect 259 447 286 464
rect 259 430 264 447
rect 281 430 286 447
rect 259 354 286 430
rect 259 337 265 354
rect 282 337 286 354
rect 259 320 286 337
rect 259 303 265 320
rect 282 303 286 320
rect 259 286 286 303
rect 259 269 265 286
rect 282 269 286 286
rect 259 252 286 269
rect 259 235 265 252
rect 282 235 286 252
rect 259 158 286 235
rect 662 478 687 605
rect 877 598 893 605
rect 914 598 933 605
rect 958 598 974 605
rect 662 461 666 478
rect 683 461 687 478
rect 662 444 687 461
rect 662 427 666 444
rect 683 427 687 444
rect 662 360 687 427
rect 662 343 667 360
rect 684 343 687 360
rect 662 326 687 343
rect 662 309 667 326
rect 684 309 687 326
rect 920 314 933 316
rect 662 292 687 309
rect 662 275 667 292
rect 684 275 687 292
rect 912 311 936 314
rect 912 294 915 311
rect 933 294 936 311
rect 912 291 936 294
rect 922 287 933 291
rect 662 258 687 275
rect 662 241 667 258
rect 684 241 687 258
rect 662 161 687 241
rect 661 158 689 161
rect 257 155 288 158
rect 257 129 259 155
rect 286 129 288 155
rect 660 157 690 158
rect 660 131 662 157
rect 688 131 690 157
rect 660 130 690 131
rect 257 127 288 129
rect 661 128 689 130
rect 259 0 286 127
rect 443 0 481 10
rect 662 0 687 128
rect 877 1 893 8
rect 914 1 933 8
rect 958 1 974 8
<< via1 >>
rect 259 129 286 155
rect 662 131 688 157
<< metal2 >>
rect 753 548 763 555
rect 753 537 766 548
rect 1001 537 1010 555
rect 2 494 806 512
rect 1001 494 1010 512
rect 2 493 17 494
rect 0 412 14 414
rect 0 406 763 412
rect 0 394 766 406
rect 1002 394 1011 412
rect 754 362 763 365
rect 754 351 766 362
rect 1001 351 1010 369
rect 751 236 766 253
rect 1000 236 1011 254
rect 3 195 766 211
rect 4 194 766 195
rect 999 193 1010 211
rect 659 157 691 158
rect 256 129 259 155
rect 286 152 289 155
rect 659 152 662 157
rect 286 135 662 152
rect 286 129 289 135
rect 659 131 662 135
rect 688 131 691 157
rect 659 130 691 131
rect 3 96 766 113
rect 82 87 236 96
rect 999 94 1010 112
rect 753 52 766 69
rect 999 51 1010 69
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_1
timestamp 1608066871
transform 1 0 1454 0 1 400
box -1451 -400 -1278 -210
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_0
timestamp 1608066871
transform 1 0 1454 0 1 517
box -1451 -400 -1278 -210
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_0
timestamp 1606741561
transform 1 0 1335 0 1 396
box -957 -395 -734 -209
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_1
timestamp 1606741561
transform 1 0 1335 0 1 512
box -957 -395 -734 -209
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_1
timestamp 1607386385
transform 1 0 1043 0 1 -46
box -289 47 -33 232
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_2
timestamp 1607386385
transform 1 0 1043 0 -1 351
box -289 47 -33 232
use sky130_hilas_wellContact  sky130_hilas_wellContact_1
timestamp 1606753443
transform 1 0 1451 0 1 675
box -1449 -441 -1275 -255
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_2
timestamp 1608066871
transform 1 0 1454 0 1 706
box -1451 -400 -1278 -210
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_2
timestamp 1606741561
transform 1 0 1335 0 1 697
box -957 -395 -734 -209
use sky130_hilas_wellContact  sky130_hilas_wellContact_0
timestamp 1606753443
transform 1 0 1854 0 1 668
box -1449 -441 -1275 -255
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_0
timestamp 1607386385
transform 1 0 1043 0 1 254
box -289 47 -33 232
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_3
timestamp 1608066871
transform 1 0 1454 0 1 815
box -1451 -400 -1278 -210
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_3
timestamp 1606741561
transform 1 0 1335 0 1 814
box -957 -395 -734 -209
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_3
timestamp 1607386385
transform 1 0 1043 0 -1 652
box -289 47 -33 232
<< labels >>
rlabel metal2 2 493 14 512 0 ROW1
port 1 nsew analog default
rlabel metal2 0 395 12 414 0 ROW2
port 2 nsew analog default
rlabel metal2 3 195 15 211 0 ROW3
port 3 nsew analog default
rlabel metal2 3 97 17 112 0 ROW4
port 4 nsew analog default
rlabel metal1 38 591 78 605 0 VTUN
port 5 nsew analog default
rlabel metal1 38 0 78 10 0 VTUN
port 5 nsew analog default
rlabel metal1 443 0 481 10 0 GATE1
port 6 nsew analog default
rlabel metal1 443 595 481 605 0 GATE1
port 6 nsew analog default
rlabel metal1 958 598 974 605 0 VINJ
port 7 nsew power default
rlabel metal1 877 598 893 605 0 VPWR
port 8 nsew power default
rlabel metal1 914 598 933 605 0 COLSEL1
rlabel metal1 958 1 974 8 0 VINJ
port 7 nsew power default
rlabel metal1 877 1 893 8 0 VPWR
port 8 nsew power default
rlabel metal1 914 1 933 8 0 COLSEL1
port 9 nsew analog default
rlabel metal2 1001 537 1010 555 0 DRAIN1
port 10 nsew analog default
rlabel metal2 1001 494 1010 512 0 ROW1
port 11 nsew analog default
rlabel metal2 1001 351 1010 369 0 DRAIN2
port 13 nsew
rlabel metal2 1002 394 1011 412 0 ROW2
port 12 nsew analog default
rlabel metal2 1000 236 1011 254 0 DRAIN3
port 14 nsew analog default
rlabel metal2 999 193 1010 211 0 ROW3
port 15 nsew analog default
rlabel metal2 999 94 1010 112 0 ROW4
port 16 nsew analog default
rlabel metal2 999 51 1010 69 0 DRAIN4
port 17 nsew analog default
rlabel metal1 259 597 286 605 0 VGND
port 18 nsew
rlabel metal1 662 600 687 605 0 VGND
port 18 nsew
rlabel metal1 259 0 286 7 0 VGND
port 18 nsew
rlabel metal1 662 0 687 7 0 VGND
port 18 nsew
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
