* Copyright 2020 The Hilas PDK Authors
* 
* This file is part of HILAS.
* 
* HILAS is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published by
* the Free Software Foundation, version 3 of the License.
* 
* HILAS is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
* 
* You should have received a copy of the GNU Lesser General Public License
* along with HILAS.  If not, see <https://www.gnu.org/licenses/>.
* 
* Licensed under the Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
* https://www.gnu.org/licenses/lgpl-3.0.en.html
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
* SPDX-License-Identifier: LGPL-3.0
* 
* 

* NGSPICE file created from sky130_hilas_capacitorSize04.ext - technology: sky130A

.subckt sky130_hilas_CapModule01a VSUBS m3_n832_n432# c1_n802_n404#
X0 c1_n802_n404# m3_n832_n432# sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
.ends

.subckt sky130_hilas_capacitorSize04 CAP1TERM02 CAP2TERM02 CAP2TERM01 CAP1TERM01
Xsky130_hilas_CapModule01a_0 VSUBS CAP2TERM02 CAP2TERM01 sky130_hilas_CapModule01a
Xsky130_hilas_CapModule01a_1 VSUBS CAP1TERM02 CAP1TERM01 sky130_hilas_CapModule01a
.ends

