* NGSPICE file created from /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_DAC6TransistorStack01b.ext - technology: sky130A

.subckt sky130_hilas_pFETdevice01d VSUBS w_n158_n156#
X0 a_42_n38# a_n36_n84# a_n90_n38# w_n158_n156# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends

.subckt sky130_hilas_pFETdevice01 VSUBS w_n158_n156#
X0 a_42_n38# a_n158_36# a_n90_n38# w_n158_n156# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends

.subckt sky130_hilas_pFETdevice01aa VSUBS w_n160_n156#
X0 a_42_n38# a_n160_36# a_n92_n38# w_n160_n156# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends

.subckt sky130_hilas_pFETdevice01a VSUBS w_n160_n84#
X0 a_42_n38# a_n160_36# a_n92_n38# w_n160_n84# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends


* Top level circuit /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_DAC6TransistorStack01b

Xsky130_hilas_pFETdevice01d_0 VSUBS sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01d
Xsky130_hilas_pFETdevice01_0 VSUBS sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01_4 VSUBS sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01_6 VSUBS sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01aa_0 VSUBS sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01aa
Xsky130_hilas_pFETdevice01a_0 VSUBS sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01a
.end

