magic
tech sky130A
timestamp 1627742263
<< error_s >>
rect -222 173 -172 185
rect -251 143 -222 144
rect -145 143 -141 173
rect -222 131 -172 143
rect -222 112 -172 123
rect -150 112 -100 123
rect -254 111 -222 112
rect -222 70 -172 81
rect -150 70 -100 81
<< nwell >>
rect -289 48 -33 232
rect -289 47 -34 48
<< mvpmos >>
rect -222 143 -172 173
rect -222 81 -172 112
rect -150 81 -100 112
<< mvpdiff >>
rect -251 167 -222 173
rect -251 150 -247 167
rect -229 150 -222 167
rect -251 143 -222 150
rect -172 166 -141 173
rect -172 149 -165 166
rect -146 149 -141 166
rect -172 143 -141 149
rect -254 105 -222 112
rect -254 88 -247 105
rect -229 88 -222 105
rect -254 81 -222 88
rect -172 81 -150 112
rect -100 105 -66 112
rect -100 88 -93 105
rect -73 88 -66 105
rect -100 81 -66 88
<< mvpdiffc >>
rect -247 150 -229 167
rect -165 149 -146 166
rect -247 88 -229 105
rect -93 88 -73 105
<< mvnsubdiff >>
rect -100 169 -66 183
rect -100 151 -93 169
rect -73 151 -66 169
rect -100 139 -66 151
<< mvnsubdiffcont >>
rect -93 151 -73 169
<< poly >>
rect -222 173 -172 188
rect -137 158 -117 199
rect -222 136 -172 143
rect -289 119 -172 136
rect -137 127 -116 158
rect -222 112 -172 119
rect -150 112 -100 127
rect -222 66 -172 81
rect -150 47 -100 81
<< locali >>
rect -255 150 -247 167
rect -229 150 -221 167
rect -166 166 -146 174
rect -166 149 -165 166
rect -166 138 -146 149
rect -166 121 -165 138
rect -148 121 -146 138
rect -166 117 -146 121
rect -94 169 -72 177
rect -94 151 -93 169
rect -73 151 -72 169
rect -94 135 -72 151
rect -94 118 -92 135
rect -75 118 -72 135
rect -93 115 -72 118
rect -93 105 -73 115
rect -255 88 -247 105
rect -229 88 -221 105
rect -93 80 -73 88
<< viali >>
rect -165 121 -148 138
rect -92 118 -75 135
<< metal1 >>
rect -166 163 -150 232
rect -166 141 -146 163
rect -126 158 -110 232
rect -85 181 -69 232
rect -85 172 -68 181
rect -127 146 -110 158
rect -168 138 -145 141
rect -168 121 -165 138
rect -148 121 -145 138
rect -168 117 -145 121
rect -166 115 -146 117
rect -166 47 -150 115
rect -129 47 -110 146
rect -96 167 -68 172
rect -96 135 -69 167
rect -96 118 -92 135
rect -75 118 -69 135
rect -96 112 -69 118
rect -85 47 -69 112
<< metal2 >>
rect -289 140 -280 158
rect -250 140 -33 158
rect -251 97 -33 115
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1627742263
transform 1 0 -266 0 -1 101
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1627742263
transform 1 0 -266 0 -1 156
box -14 -15 20 18
<< end >>
