magic
tech sky130A
timestamp 1628704327
<< error_s >>
rect 62 542 101 545
rect 62 500 101 503
rect 62 446 101 449
rect 62 404 101 407
rect 62 350 101 353
rect 62 308 101 311
rect 62 254 101 257
rect 62 212 101 215
rect 62 158 101 161
rect 62 116 101 119
rect 62 62 101 65
rect 62 20 101 23
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_0
timestamp 1628704221
transform 1 0 80 0 1 138
box 0 0 172 121
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_1
timestamp 1628704221
transform 1 0 80 0 1 234
box 0 0 172 121
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_4
timestamp 1628704221
transform 1 0 80 0 1 330
box 0 0 172 121
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_2
timestamp 1628704221
transform 1 0 80 0 1 426
box 0 0 172 121
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_3
timestamp 1628704221
transform 1 0 80 0 1 522
box 0 0 172 121
use sky130_hilas_pFETdevice01a  sky130_hilas_pFETdevice01a_0
timestamp 1628285143
transform 1 0 80 0 1 42
box -80 -42 81 43
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
