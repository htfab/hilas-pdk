magic
tech sky130A
timestamp 1629137215
<< checkpaint >>
rect -630 -630 969 917
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_2
timestamp 1629137178
transform 1 0 165 0 1 0
box 0 0 119 287
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_1
timestamp 1629137178
transform 1 0 110 0 1 0
box 0 0 119 287
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_0
timestamp 1629137178
transform 1 0 55 0 1 0
box 0 0 119 287
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_4
timestamp 1629137178
transform 1 0 0 0 1 0
box 0 0 119 287
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_3
timestamp 1629137178
transform 1 0 220 0 1 0
box 0 0 119 287
<< end >>
