* Copyright 2020 The Hilas PDK Authors
* 
* This file is part of HILAS.
* 
* HILAS is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published by
* the Free Software Foundation, version 3 of the License.
* 
* HILAS is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
* 
* You should have received a copy of the GNU Lesser General Public License
* along with HILAS.  If not, see <https://www.gnu.org/licenses/>.
* 
* Licensed under the Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
* https://www.gnu.org/licenses/lgpl-3.0.en.html
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
* SPDX-License-Identifier: LGPL-3.0
* 
* 

* NGSPICE file created from sky130_hilas_Tgate4Single01.ext - technology: sky130A

.subckt sky130_hilas_TgateSingle01Part1 sky130_hilas_m12m2_3/SUB a_582_n188# output
+ a_582_n314# a_514_n112#
X0 sky130_hilas_m12m2_3/SUB a_514_n112# a_582_n188# sky130_hilas_m12m2_3/SUB sky130_fd_pr__nfet_01v8 w=300000u l=400000u
X1 output a_514_n112# a_582_n314# sky130_hilas_m12m2_3/SUB sky130_fd_pr__nfet_01v8 w=310000u l=400000u
.ends

.subckt sky130_hilas_TgateSingle01Part2 a_18_n340# a_n40_n314# SUB w_n134_n362# li_n36_n176#
+ a_98_n314# a_n36_n112#
X0 a_98_n314# a_18_n340# a_n40_n314# w_n134_n362# sky130_fd_pr__pfet_01v8 w=310000u l=400000u
.ends

.subckt sky130_hilas_TgateSingle01 m2_n526_n340# a_n468_n112# SUB w_n502_n362# sky130_hilas_TgateSingle01Part1_0/output
Xsky130_hilas_TgateSingle01Part1_0 SUB a_n196_n192# sky130_hilas_TgateSingle01Part1_0/output
+ m2_n526_n340# a_n468_n112# sky130_hilas_TgateSingle01Part1
Xsky130_hilas_TgateSingle01Part2_0 a_n196_n192# m2_n526_n340# SUB w_n502_n362# a_n196_n192#
+ sky130_hilas_TgateSingle01Part1_0/output a_n468_n112# sky130_hilas_TgateSingle01Part2
X0 a_n196_n192# a_n468_n112# w_n502_n362# w_n502_n362# sky130_fd_pr__pfet_01v8 w=320000u l=400000u
.ends

.subckt sky130_hilas_Tgate4Single01 INPUT1_4 VPWR SELECT4 SELECT3 INPUT1_3 INPUT1_2
+ SELECT2 SELECT1 INPUT1_1 VGND OUTPUT1 OUTPUT2 OUTPUT3 OUTPUT4
Xsky130_hilas_TgateSingle01_0 INPUT1_1 SELECT1 VGND VPWR OUTPUT1 sky130_hilas_TgateSingle01
Xsky130_hilas_TgateSingle01_1 INPUT1_4 SELECT4 VGND VPWR OUTPUT4 sky130_hilas_TgateSingle01
Xsky130_hilas_TgateSingle01_2 INPUT1_3 SELECT3 VGND VPWR OUTPUT3 sky130_hilas_TgateSingle01
Xsky130_hilas_TgateSingle01_3 INPUT1_2 SELECT2 VGND VPWR OUTPUT2 sky130_hilas_TgateSingle01
.ends

