magic
tech sky130A
timestamp 1606871823
<< error_s >>
rect -338 150 -332 156
rect -285 150 -279 156
rect -344 100 -338 106
rect -279 100 -273 106
rect 85 91 91 97
rect 190 91 196 97
rect 79 41 85 47
rect 196 41 202 47
rect 85 -210 91 -204
rect 190 -210 196 -204
rect -338 -265 -332 -259
rect -285 -265 -279 -259
rect 79 -260 85 -254
rect 196 -260 202 -254
rect -344 -315 -338 -309
rect -279 -315 -273 -309
rect 514 -314 524 -313
<< nwell >>
rect -337 -242 -281 0
<< mvnsubdiff >>
rect -337 -242 -281 0
<< poly >>
rect -237 134 331 151
rect -237 126 -185 134
rect 45 91 64 134
rect 220 90 237 134
rect 46 -293 63 -260
rect 220 -293 237 -260
rect -280 -310 331 -293
<< metal1 >>
rect -361 -382 -319 223
<< metal2 >>
rect 484 173 516 175
rect -396 155 516 173
rect 510 -315 514 -313
rect -394 -330 514 -315
use FGVaractorCapacitor02  FGVaractorCapacitor02_2
timestamp 1606868103
transform 1 0 986 0 -1 -231
box -1005 -380 -733 -211
use FGVaractorCapacitor02  FGVaractorCapacitor02_0
timestamp 1606868103
transform 1 0 986 0 1 62
box -1005 -380 -733 -211
use horizTransCell01  horizTransCell01_1
timestamp 1606869277
transform 1 0 790 0 -1 270
box -476 47 -33 359
use horizTransCell01  horizTransCell01_0
timestamp 1606869277
transform 1 0 790 0 1 -429
box -476 47 -33 359
use TunCap01  TunCap01_1
timestamp 1606740587
transform 1 0 1056 0 1 18
box -1451 -400 -1278 -210
use wellContact  wellContact_0
timestamp 1606753443
transform 1 0 1054 0 1 231
box -1449 -441 -1275 -255
use wellContact  wellContact_1
timestamp 1606753443
transform 1 0 1054 0 1 404
box -1449 -441 -1275 -255
use TunCap01  TunCap01_3
timestamp 1606740587
transform 1 0 1056 0 1 433
box -1451 -400 -1278 -210
<< end >>
