magic
tech sky130A
timestamp 1627060558
<< metal2 >>
rect 0 528 1042 546
rect 0 485 1042 503
rect 3 385 1042 403
rect 851 360 1042 361
rect 3 342 1042 360
rect 2 280 29 308
rect 1006 281 1042 309
rect 3 227 1042 244
rect 3 185 1042 202
rect 3 87 1042 104
rect 3 43 1042 60
<< metal3 >>
rect 823 255 1019 330
<< metal4 >>
rect 116 320 217 321
rect 45 270 380 320
rect 45 269 152 270
rect 316 158 379 270
rect 316 128 531 158
rect 349 127 531 128
use sky130_hilas_m22m4  sky130_hilas_m22m4_1
timestamp 1607701799
transform 1 0 987 0 1 291
box -36 -36 43 39
use sky130_hilas_m22m4  sky130_hilas_m22m4_0
timestamp 1607701799
transform 1 0 38 0 1 290
box -36 -36 43 39
use sky130_hilas_CapModule02  sky130_hilas_CapModule02_0
timestamp 1607802006
transform 1 0 589 0 1 247
box -443 -247 277 336
<< labels >>
rlabel metal2 2 280 9 308 0 CAPTERM01
port 2 nsew analog default
rlabel metal2 1030 281 1042 309 0 CAPTERM02
port 1 nsew analog default
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
