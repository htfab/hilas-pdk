magic
tech sky130A
timestamp 1637801776
<< error_p >>
rect -178 275 -126 283
rect -126 270 -98 275
rect 176 271 226 281
rect 145 270 176 271
rect -178 233 -126 241
rect 176 229 226 239
rect -252 210 -199 219
rect -105 210 -53 220
rect -279 204 -252 210
rect -53 205 -26 210
rect 105 209 155 220
rect 247 209 297 220
rect 76 205 105 209
rect -279 185 -276 204
rect -252 168 -199 177
rect -105 168 -53 178
rect 105 167 155 178
rect 247 167 297 178
<< nwell >>
rect -336 144 8 308
<< mvnmos >>
rect 176 239 226 271
rect 105 178 155 209
rect 247 178 297 209
<< mvpmos >>
rect -178 241 -126 275
rect -252 177 -199 210
rect -105 178 -53 210
<< mvndiff >>
rect 145 263 176 271
rect 145 246 152 263
rect 169 246 176 263
rect 145 239 176 246
rect 226 263 253 271
rect 226 246 232 263
rect 249 246 253 263
rect 226 239 253 246
rect 76 202 105 209
rect 76 185 81 202
rect 98 185 105 202
rect 76 178 105 185
rect 155 202 183 209
rect 155 185 161 202
rect 178 185 183 202
rect 155 178 183 185
rect 219 202 247 209
rect 219 185 224 202
rect 241 185 247 202
rect 219 178 247 185
rect 297 202 326 209
rect 297 185 303 202
rect 320 185 326 202
rect 297 178 326 185
<< mvpdiff >>
rect -206 267 -178 275
rect -206 250 -201 267
rect -184 250 -178 267
rect -206 241 -178 250
rect -126 267 -98 275
rect -126 250 -120 267
rect -103 250 -98 267
rect -126 241 -98 250
rect -279 202 -252 210
rect -279 185 -275 202
rect -258 185 -252 202
rect -279 177 -252 185
rect -199 202 -171 210
rect -199 185 -193 202
rect -176 185 -171 202
rect -199 177 -171 185
rect -132 202 -105 210
rect -132 185 -128 202
rect -111 185 -105 202
rect -132 178 -105 185
rect -53 202 -26 210
rect -53 185 -47 202
rect -30 185 -26 202
rect -53 178 -26 185
<< mvndiffc >>
rect 152 246 169 263
rect 232 246 249 263
rect 81 185 98 202
rect 161 185 178 202
rect 224 185 241 202
rect 303 185 320 202
<< mvpdiffc >>
rect -201 250 -184 267
rect -120 250 -103 267
rect -275 185 -258 202
rect -193 185 -176 202
rect -128 185 -111 202
rect -47 185 -30 202
<< psubdiff >>
rect 292 264 333 271
rect 292 247 304 264
rect 321 247 333 264
rect 292 239 333 247
<< mvnsubdiff >>
rect -286 267 -245 275
rect -286 250 -274 267
rect -257 250 -245 267
rect -286 241 -245 250
<< psubdiffcont >>
rect 304 247 321 264
<< mvnsubdiffcont >>
rect -274 250 -257 267
<< poly >>
rect -143 289 194 295
rect -178 284 194 289
rect -178 278 226 284
rect -178 275 -126 278
rect 25 275 60 278
rect 25 258 34 275
rect 51 258 60 275
rect 176 271 226 278
rect -74 251 -39 257
rect 25 251 60 258
rect -322 226 -236 227
rect -322 212 -199 226
rect -178 225 -126 241
rect -74 234 -64 251
rect -47 234 -39 251
rect -74 230 -39 234
rect -74 225 123 230
rect 176 225 226 239
rect -322 202 -295 212
rect -252 210 -199 212
rect -105 223 123 225
rect -105 213 155 223
rect -105 210 -53 213
rect -322 185 -317 202
rect -300 185 -295 202
rect -322 177 -295 185
rect 105 209 155 213
rect 247 209 297 223
rect -252 164 -199 177
rect -105 165 -53 178
rect 105 165 155 178
rect 247 165 297 178
<< polycont >>
rect 34 258 51 275
rect -64 234 -47 251
rect -317 185 -300 202
<< locali >>
rect -274 267 -257 279
rect 34 275 51 283
rect -201 267 -184 275
rect -120 267 -103 275
rect -274 248 -272 250
rect -184 250 -180 267
rect -274 238 -257 248
rect -201 210 -180 250
rect -124 250 -120 267
rect -124 242 -103 250
rect -64 251 -47 259
rect 223 264 249 271
rect 303 264 321 277
rect 223 263 304 264
rect 47 254 51 258
rect 34 250 51 254
rect -124 210 -107 242
rect -50 232 -47 234
rect -64 222 -47 232
rect 90 246 152 263
rect 169 246 177 263
rect 223 246 232 263
rect 249 247 304 263
rect 249 246 321 247
rect -317 202 -300 210
rect -302 183 -300 185
rect -317 177 -300 183
rect -275 204 -258 210
rect -275 202 -250 204
rect -258 197 -250 202
rect -275 180 -271 185
rect -254 180 -250 197
rect -201 202 -176 210
rect -201 185 -193 202
rect -275 177 -250 180
rect -274 175 -250 177
rect -193 176 -176 185
rect -128 202 -107 210
rect 90 202 107 246
rect 223 232 249 246
rect 303 235 321 246
rect 223 214 226 232
rect 244 214 249 232
rect 223 202 249 214
rect -111 185 -107 202
rect -56 185 -47 202
rect -30 198 81 202
rect -30 185 21 198
rect -128 177 -111 185
rect 38 185 81 198
rect 98 185 107 202
rect 152 185 161 202
rect 178 185 224 202
rect 241 185 249 202
rect 294 185 303 202
rect 320 185 328 202
<< viali >>
rect -272 250 -257 265
rect -257 250 -255 265
rect -272 248 -255 250
rect 30 258 34 271
rect 34 258 47 271
rect 30 254 47 258
rect -67 234 -64 249
rect -64 234 -50 249
rect -67 232 -50 234
rect -319 185 -317 200
rect -317 185 -302 200
rect -319 183 -302 185
rect -271 185 -258 197
rect -258 185 -254 197
rect -271 180 -254 185
rect 226 214 244 232
rect 21 181 38 198
<< metal1 >>
rect -275 270 -253 304
rect -275 265 -252 270
rect -275 248 -272 265
rect -255 248 -252 265
rect -275 244 -252 248
rect -328 205 -297 211
rect -328 179 -325 205
rect -299 179 -297 205
rect -328 176 -297 179
rect -275 204 -253 244
rect -73 228 -69 254
rect -43 228 -40 254
rect 24 253 30 279
rect 56 253 67 279
rect 24 250 67 253
rect 222 232 249 305
rect 222 214 226 232
rect 244 214 249 232
rect -275 197 -250 204
rect -275 180 -271 197
rect -254 180 -250 197
rect -275 173 -250 180
rect 11 201 50 202
rect 11 175 17 201
rect 43 175 50 201
rect -275 153 -253 173
rect 222 153 249 214
rect 304 205 335 208
rect 304 179 307 205
rect 333 179 335 205
rect 304 176 335 179
<< via1 >>
rect -325 200 -299 205
rect -325 183 -319 200
rect -319 183 -302 200
rect -302 183 -299 200
rect -325 179 -299 183
rect -69 249 -43 254
rect -69 232 -67 249
rect -67 232 -50 249
rect -50 232 -43 249
rect -69 228 -43 232
rect 30 271 56 279
rect 30 254 47 271
rect 47 254 56 271
rect 30 253 56 254
rect 17 198 43 201
rect 17 181 21 198
rect 21 181 38 198
rect 38 181 43 198
rect 17 175 43 181
rect 307 179 333 205
<< metal2 >>
rect -337 279 67 289
rect -337 273 30 279
rect -73 246 -69 254
rect -100 244 -69 246
rect -336 228 -69 244
rect -43 228 -40 254
rect 25 253 30 273
rect 56 253 67 279
rect 25 250 67 253
rect 304 205 335 208
rect -328 195 -325 205
rect -336 179 -325 195
rect -299 179 -296 205
rect 13 175 17 201
rect 43 193 50 201
rect 43 192 116 193
rect 304 192 307 205
rect 43 179 307 192
rect 333 192 335 205
rect 333 179 351 192
rect 43 175 351 179
<< labels >>
rlabel metal2 345 175 351 192 0 Output
rlabel metal2 -337 273 -331 289 0 Input1
rlabel space -337 228 -331 244 0 Input2
rlabel space -337 179 -331 195 0 Input3
rlabel metal1 222 299 249 305 0 GND
rlabel metal1 222 153 249 158 0 GND
rlabel metal1 -275 153 -253 159 0 Vinj
rlabel metal1 -275 297 -253 304 0 Vinj
<< end >>
