magic
tech sky130A
timestamp 1628704414
<< checkpaint >>
rect -630 -622 719 910
<< error_s >>
rect 394 173 411 174
rect 418 162 419 203
rect 382 150 386 162
rect 418 150 423 162
rect 418 134 419 150
rect 418 102 419 133
rect 418 44 419 73
<< nwell >>
rect 248 304 467 477
<< nmos >>
rect 301 203 334 232
rect 386 203 419 232
rect 301 73 334 102
rect 386 73 419 102
<< pmos >>
rect 269 356 337 386
rect 373 356 441 386
<< ndiff >>
rect 301 256 334 260
rect 301 239 309 256
rect 326 239 334 256
rect 301 232 334 239
rect 386 256 419 260
rect 386 239 394 256
rect 411 239 419 256
rect 386 232 419 239
rect 301 196 334 203
rect 301 179 309 196
rect 326 179 334 196
rect 301 173 334 179
rect 301 125 334 132
rect 301 108 309 125
rect 326 108 334 125
rect 301 102 334 108
rect 386 196 419 203
rect 386 179 394 196
rect 411 179 419 196
rect 386 173 419 179
rect 386 126 419 133
rect 386 109 394 126
rect 411 109 419 126
rect 386 102 419 109
rect 301 66 334 73
rect 301 49 308 66
rect 326 49 334 66
rect 301 45 334 49
rect 386 67 419 73
rect 386 50 393 67
rect 412 50 419 67
rect 386 44 419 50
<< pdiff >>
rect 269 410 337 416
rect 269 393 277 410
rect 295 393 313 410
rect 331 393 337 410
rect 269 386 337 393
rect 373 410 441 416
rect 373 393 381 410
rect 399 393 418 410
rect 437 393 441 410
rect 373 386 441 393
rect 269 349 337 356
rect 269 332 277 349
rect 295 332 313 349
rect 331 332 337 349
rect 269 323 337 332
rect 373 349 441 356
rect 373 332 379 349
rect 397 332 415 349
rect 433 332 441 349
rect 373 328 441 332
rect 380 323 441 328
<< ndiffc >>
rect 309 239 326 256
rect 394 239 411 256
rect 309 179 326 196
rect 309 108 326 125
rect 394 179 411 196
rect 394 109 411 126
rect 308 49 326 66
rect 393 50 412 67
<< pdiffc >>
rect 277 393 295 410
rect 313 393 331 410
rect 381 393 399 410
rect 418 393 437 410
rect 277 332 295 349
rect 313 332 331 349
rect 379 332 397 349
rect 415 332 433 349
<< psubdiff >>
rect 301 161 334 173
rect 301 144 309 161
rect 326 144 334 161
rect 301 132 334 144
rect 386 162 419 173
rect 386 145 394 162
rect 411 145 419 162
rect 386 134 419 145
rect 386 133 418 134
<< nsubdiff >>
rect 269 445 337 457
rect 269 428 277 445
rect 295 428 313 445
rect 331 428 337 445
rect 269 416 337 428
rect 373 445 441 457
rect 373 428 381 445
rect 399 428 418 445
rect 437 428 441 445
rect 373 416 441 428
<< psubdiffcont >>
rect 309 144 326 161
rect 394 145 411 162
<< nsubdiffcont >>
rect 277 428 295 445
rect 313 428 331 445
rect 381 428 399 445
rect 418 428 437 445
<< poly >>
rect 256 356 269 386
rect 337 356 373 386
rect 441 356 454 386
rect 345 312 362 356
rect 339 304 366 312
rect 339 287 344 304
rect 361 287 366 304
rect 339 279 366 287
rect 31 215 58 219
rect 276 203 301 232
rect 334 203 347 232
rect 372 203 386 232
rect 419 203 442 232
rect 276 102 292 203
rect 426 102 442 203
rect 276 73 301 102
rect 334 73 347 102
rect 371 73 386 102
rect 419 73 442 102
rect 31 69 58 72
rect 276 34 292 73
rect 276 26 335 34
rect 426 33 442 73
rect 276 9 308 26
rect 326 9 335 26
rect 276 3 335 9
rect 386 25 442 33
rect 386 8 395 25
rect 412 8 442 25
rect 386 3 442 8
<< polycont >>
rect 344 287 361 304
rect 308 9 326 26
rect 395 8 412 25
<< locali >>
rect 269 428 277 445
rect 295 428 313 445
rect 331 428 381 445
rect 399 428 418 445
rect 437 428 445 445
rect 269 410 445 428
rect 269 393 277 410
rect 295 393 313 410
rect 331 393 381 410
rect 399 393 418 410
rect 437 393 445 410
rect 269 332 277 349
rect 295 332 313 349
rect 331 332 340 349
rect 371 332 379 349
rect 397 332 415 349
rect 433 332 441 349
rect 304 315 340 332
rect 304 304 369 315
rect 304 287 344 304
rect 361 287 369 304
rect 304 279 369 287
rect 304 256 331 279
rect 394 257 419 332
rect 386 256 419 257
rect 301 239 309 256
rect 326 239 334 256
rect 386 239 394 256
rect 411 239 419 256
rect 297 179 309 196
rect 326 179 338 196
rect 297 172 338 179
rect 382 179 394 196
rect 411 179 423 196
rect 382 172 423 179
rect 297 162 423 172
rect 297 161 394 162
rect 297 144 309 161
rect 326 145 394 161
rect 411 145 423 162
rect 326 144 423 145
rect 297 134 423 144
rect 297 125 338 134
rect 297 108 309 125
rect 326 108 338 125
rect 382 126 423 134
rect 382 109 394 126
rect 411 109 423 126
rect 300 49 308 66
rect 326 49 334 66
rect 385 50 393 67
rect 412 50 421 67
rect 385 49 421 50
rect 308 26 326 49
rect 308 0 326 9
rect 393 25 412 49
rect 393 8 395 25
rect 393 0 412 8
use sky130_hilas_nFET03  sky130_hilas_nFET03_3
timestamp 1628285143
transform 1 0 31 0 1 238
box -31 -19 58 42
use sky130_hilas_nFET03  sky130_hilas_nFET03_2
timestamp 1628285143
transform 1 0 31 0 1 173
box -31 -19 58 42
use sky130_hilas_nFET03  sky130_hilas_nFET03_1
timestamp 1628285143
transform 1 0 31 0 1 91
box -31 -19 58 42
use sky130_hilas_nFET03  sky130_hilas_nFET03_0
timestamp 1628285143
transform 1 0 31 0 1 27
box -31 -19 58 42
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
