magic
tech sky130A
magscale 1 2
timestamp 1632256330
<< error_s >>
rect 4264 1878 4274 1886
rect 4264 1858 4392 1878
rect 4264 1847 4275 1858
rect 4294 1344 4306 1414
rect 4322 1344 4334 1386
rect 4136 1332 4236 1344
rect 4280 1332 4380 1344
rect 3370 1292 3408 1320
rect 3458 1294 3490 1322
rect 4294 1320 4306 1332
rect 4322 1292 4334 1332
rect 4136 1248 4236 1260
rect 4280 1248 4380 1260
rect 3014 1234 3052 1240
rect 2980 1184 2996 1218
rect 3014 1200 3030 1234
rect 3014 1194 3052 1200
rect 3546 1168 3574 1204
rect 4274 1198 4379 1202
rect 2958 1106 2970 1116
rect 3650 1044 3654 1144
rect 3734 1044 3738 1144
rect 3920 1044 3926 1144
rect 4004 1044 4010 1144
rect 4274 1130 4290 1198
rect 4311 1191 4379 1198
rect 4322 1130 4368 1191
rect 4437 1130 4448 1141
rect 4234 1116 4290 1130
rect 4392 1116 4448 1130
rect 4192 1030 4290 1116
rect 1308 308 1552 924
rect 3650 886 3654 986
rect 3734 886 3738 986
rect 3920 888 3926 986
rect 4004 888 4010 986
rect 4274 962 4290 1030
rect 4300 1020 4392 1030
rect 4314 986 4392 1020
rect 4314 970 4384 986
rect 2874 710 2882 812
rect 2902 682 2910 840
rect 3014 836 3052 842
rect 3014 824 3016 836
rect 3014 802 3026 824
rect 3014 796 3052 802
rect 2976 756 3010 790
rect 3852 764 4514 888
rect 3304 740 3318 746
rect 3276 712 3290 720
rect 3276 674 3292 712
rect 3304 694 3320 740
rect 2726 662 2758 672
rect 2724 642 2758 662
rect 2920 658 2958 664
rect 2920 654 2936 658
rect 2942 654 2958 658
rect 2920 638 2958 654
rect 2760 636 2794 638
rect 2892 636 2958 638
rect 2760 630 2792 636
rect 2742 608 2792 630
rect 2886 630 2902 636
rect 2886 596 2910 630
rect 2920 618 2958 636
rect 2976 608 3010 642
rect 3012 622 3050 628
rect 3012 588 3020 622
rect 3012 582 3050 588
rect 3174 526 3230 552
rect 3146 498 3202 524
rect 3650 412 3654 512
rect 3734 412 3738 512
rect 3920 412 3926 512
rect 4004 412 4010 512
rect 2774 326 2810 328
rect 2960 326 2972 336
rect 2774 324 2776 326
rect 1326 110 1410 264
rect 3650 254 3654 354
rect 3734 254 3738 354
rect 3920 254 3926 354
rect 4004 254 4010 354
rect 2988 224 3008 234
rect 3048 232 3100 246
rect 3048 228 3068 232
rect 3092 196 3094 222
rect 3092 194 3120 196
rect 3546 194 3574 230
rect 4136 138 4236 150
rect 4280 138 4380 150
rect 1410 96 1494 110
rect 3370 94 3408 122
rect 3458 94 3490 122
rect 4136 54 4236 66
rect 4280 54 4380 66
<< nwell >>
rect 1374 374 1486 858
rect 1326 96 1410 110
<< psubdiff >>
rect 1858 774 1908 1100
rect 1858 740 1864 774
rect 1902 740 1908 774
rect 1858 714 1908 740
rect 1858 708 2584 714
rect 1858 706 2340 708
rect 1858 672 1906 706
rect 1944 672 1992 706
rect 2030 672 2080 706
rect 2118 672 2160 706
rect 2198 672 2248 706
rect 2286 674 2340 706
rect 2378 706 2584 708
rect 2378 674 2428 706
rect 2286 672 2428 674
rect 2466 672 2520 706
rect 2558 672 2584 706
rect 1858 664 2584 672
rect 1858 638 1908 664
rect 1858 604 1864 638
rect 1902 604 1908 638
rect 1858 296 1908 604
<< mvnsubdiff >>
rect 1374 374 1486 858
<< psubdiffcont >>
rect 1864 740 1902 774
rect 1906 672 1944 706
rect 1992 672 2030 706
rect 2080 672 2118 706
rect 2160 672 2198 706
rect 2248 672 2286 706
rect 2340 674 2378 708
rect 2428 672 2466 706
rect 2520 672 2558 706
rect 1864 604 1902 638
<< poly >>
rect 1574 1130 2710 1160
rect 1574 1126 2686 1130
rect 1574 1110 1678 1126
rect 2044 1040 2088 1126
rect 2380 1040 2424 1126
rect 2600 960 2676 1060
rect 2600 438 2630 960
rect 2816 802 2844 804
rect 2816 596 2860 802
rect 2600 392 2680 438
rect 2592 382 2680 392
rect 2592 348 2608 382
rect 2642 348 2680 382
rect 2592 338 2680 348
rect 2042 272 2082 338
rect 2386 272 2426 338
rect 2592 332 2648 338
rect 1488 268 2682 272
rect 1488 238 2710 268
<< polycont >>
rect 2608 348 2642 382
<< locali >>
rect 2820 1184 2996 1218
rect 2820 1106 2854 1184
rect 2776 1072 2854 1106
rect 2936 1072 2980 1106
rect 2490 914 2706 948
rect 2772 914 2988 948
rect 1864 774 1902 790
rect 2976 756 2992 790
rect 1864 708 1902 740
rect 1864 706 2340 708
rect 1864 672 1906 706
rect 1944 672 1992 706
rect 2030 672 2080 706
rect 2118 672 2160 706
rect 2198 672 2248 706
rect 2286 674 2340 706
rect 2378 706 2574 708
rect 2378 674 2428 706
rect 2286 672 2428 674
rect 2466 672 2520 706
rect 2558 672 2574 706
rect 1864 638 1902 672
rect 2724 642 2758 756
rect 2760 636 2776 638
rect 2892 636 2902 638
rect 2760 628 2902 636
rect 2756 620 2902 628
rect 1864 588 1902 604
rect 2742 596 2910 620
rect 2976 608 2986 642
rect 2460 450 2708 484
rect 2772 450 2988 484
rect 2608 386 2642 398
rect 2608 330 2642 344
rect 2776 324 2868 326
rect 2774 294 2868 324
rect 2776 292 2868 294
rect 2938 292 2980 326
rect 2830 224 2868 292
rect 2830 188 3022 224
<< viali >>
rect 2604 382 2646 386
rect 2604 348 2608 382
rect 2608 348 2642 382
rect 2642 348 2646 382
rect 2604 344 2646 348
<< metal1 >>
rect 1326 94 1410 1304
rect 1822 94 1868 1304
rect 2606 398 2642 1304
rect 2596 386 2654 398
rect 2596 344 2604 386
rect 2646 344 2654 386
rect 2596 330 2654 344
rect 2606 94 2642 330
rect 2816 94 2858 1304
rect 2902 94 2940 1304
rect 2992 746 3034 1304
rect 3370 1292 3408 1304
rect 3458 1294 3490 1304
rect 3290 656 3338 740
rect 2992 194 3030 644
rect 3092 194 3094 196
rect 2986 94 3032 194
rect 3370 94 3408 104
rect 3458 94 3490 104
<< metal2 >>
rect 3016 1204 3080 1208
rect 1258 1168 3080 1204
rect 3546 1168 3562 1204
rect 1258 858 3200 896
rect 1258 712 3290 720
rect 1258 674 3292 712
rect 1258 486 3202 524
rect 3068 228 3100 232
rect 1258 218 3100 228
rect 1258 198 3076 218
rect 3546 194 3562 230
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_2
timestamp 1632251432
transform -1 0 544 0 -1 396
box 0 0 544 338
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1632251332
transform 1 0 1842 0 1 674
box 0 0 46 58
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1632251356
transform 1 0 3174 0 1 526
box 0 0 68 66
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1632251332
transform 1 0 2916 0 1 612
box 0 0 46 58
use sky130_hilas_li2m1  sky130_hilas_li2m1_3
timestamp 1632251332
transform 1 0 3008 0 1 576
box 0 0 46 58
use sky130_hilas_li2m1  sky130_hilas_li2m1_2
timestamp 1632251332
transform 1 0 2918 0 1 296
box 0 0 46 58
use sky130_hilas_li2m1  sky130_hilas_li2m1_5
timestamp 1632251332
transform 1 0 3004 0 1 194
box 0 0 46 58
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1632251372
transform 1 0 3304 0 1 688
box 0 0 64 64
use sky130_hilas_horizTransCell01a  sky130_hilas_horizTransCell01a_0
timestamp 1632251381
transform 1 0 3628 0 1 0
box 0 0 886 634
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_0
timestamp 1632251432
transform -1 0 544 0 1 982
box 0 0 544 338
use sky130_hilas_poly2m1  sky130_hilas_poly2m1_0
timestamp 1632251319
transform 1 0 2826 0 1 710
box 0 0 66 102
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1632251356
transform 1 0 3172 0 1 864
box 0 0 68 66
use sky130_hilas_li2m1  sky130_hilas_li2m1_6
timestamp 1632251332
transform 1 0 3010 0 1 1188
box 0 0 46 58
use sky130_hilas_li2m1  sky130_hilas_li2m1_4
timestamp 1632251332
transform 1 0 2916 0 1 1076
box 0 0 46 58
use sky130_hilas_li2m1  sky130_hilas_li2m1_7
timestamp 1632251332
transform 1 0 3010 0 1 790
box 0 0 46 58
use sky130_hilas_horizTransCell01a  sky130_hilas_horizTransCell01a_1
timestamp 1632251381
transform 1 0 3628 0 -1 1398
box 0 0 886 634
use sky130_hilas_wellContact  sky130_hilas_wellContact_0
timestamp 1632251355
transform 1 0 4156 0 1 1320
box 0 0 346 372
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_1
timestamp 1632251302
transform 1 0 4160 0 1 896
box 0 0 346 380
use sky130_hilas_wellContact  sky130_hilas_wellContact_1
timestamp 1632251355
transform 1 0 4156 0 1 1666
box 0 0 346 372
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_3
timestamp 1632251302
transform 1 0 4160 0 1 1724
box 0 0 346 380
<< labels >>
rlabel metal1 1326 1290 1410 1304 0 VTUN
port 11 nsew analog default
rlabel metal1 1822 1290 1868 1304 0 VGND
port 10 nsew ground default
rlabel space 3458 1292 3490 1302 0 VINJ
port 2 nsew analog default
rlabel metal2 1258 198 1266 228 3 DRAIN2
port 12 e analog default
rlabel metal2 1258 1168 1270 1204 0 DRAIN1
port 15 nsew analog default
rlabel metal1 2902 1292 2940 1304 0 GATE1
port 9 nsew analog default
rlabel metal1 2986 96 3032 144 0 VIN2
port 7 nsew analog default
rlabel metal1 2606 94 2642 108 0 RUN
port 6 nsew analog default
rlabel metal1 2816 94 2858 108 0 PROG
port 5 nsew analog default
rlabel metal1 2606 1290 2642 1304 0 RUN
port 6 nsew analog default
rlabel metal1 2816 1292 2858 1304 0 PROG
port 5 nsew analog default
rlabel metal1 2992 1240 3034 1302 0 VIN1
port 8 nsew analog default
rlabel metal1 3370 1292 3408 1304 0 COLSEL1
port 1 nsew analog default
rlabel metal1 3370 94 3408 104 0 COLSEL1
port 1 nsew analog default
rlabel metal1 3458 94 3490 104 0 VINJ
port 2 nsew analog default
rlabel metal2 3546 1168 3562 1204 0 DRAIN1
port 3 nsew analog default
rlabel metal2 3546 194 3562 230 0 DRAIN2
port 4 nsew analog default
rlabel metal1 2902 96 2940 106 0 GATE1
port 9 nsew analog default
rlabel metal1 1822 94 1868 108 0 VGND
port 10 nsew ground default
rlabel metal1 1326 96 1410 110 0 VTUN
port 11 nsew analog default
rlabel metal2 1258 674 1270 720 0 COL1
port 16 nsew
rlabel metal2 1258 858 1270 896 0 ROW1
port 17 nsew
rlabel metal2 1258 486 1270 524 0 ROW2
port 18 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
