magic
tech sky130A
timestamp 1637801776
<< error_p >>
rect -10 15 13 21
rect -10 -2 -7 15
rect -10 -8 13 -2
<< locali >>
rect -8 15 11 18
rect -8 -2 -7 15
rect 10 -2 11 15
rect -8 -5 11 -2
<< viali >>
rect -7 -2 10 15
<< metal1 >>
rect -10 15 13 21
rect -10 -2 -7 15
rect 10 -2 13 15
rect -10 -8 13 -2
<< end >>
