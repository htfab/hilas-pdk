* Copyright 2020 The Hilas PDK Authors
* 
* This file is part of HILAS.
* 
* HILAS is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published by
* the Free Software Foundation, version 3 of the License.
* 
* HILAS is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
* 
* You should have received a copy of the GNU Lesser General Public License
* along with HILAS.  If not, see <https://www.gnu.org/licenses/>.
* 
* Licensed under the Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
* https://www.gnu.org/licenses/lgpl-3.0.en.html
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
* SPDX-License-Identifier: LGPL-3.0
* 
* 

* NGSPICE file created from sky130_hilas_pFETLarge.ext - technology: sky130A

.subckt sky130_hilas_pFETmed VSUBS a_440_n8# w_294_n44# a_388_n34# a_330_n8#
X0 a_440_n8# a_388_n34# a_330_n8# w_294_n44# sky130_fd_pr__pfet_01v8 w=2.51e+06u l=260000u
.ends

.subckt sky130_hilas_pFETLargePart1 VSUBS sky130_hilas_pFETmed_2/a_388_n34# sky130_hilas_pFETmed_4/a_330_n8#
+ sky130_hilas_pFETmed_1/a_388_n34# sky130_hilas_pFETmed_0/a_388_n34# sky130_hilas_pFETmed_3/a_330_n8#
+ sky130_hilas_pFETmed_2/a_330_n8# sky130_hilas_pFETmed_1/a_330_n8# sky130_hilas_pFETmed_4/a_440_n8#
+ sky130_hilas_pFETmed_4/a_388_n34# sky130_hilas_pFETmed_4/w_294_n44# sky130_hilas_pFETmed_3/a_388_n34#
+ sky130_hilas_pFETmed_3/a_440_n8#
Xsky130_hilas_pFETmed_0 VSUBS sky130_hilas_pFETmed_1/a_330_n8# sky130_hilas_pFETmed_4/w_294_n44#
+ sky130_hilas_pFETmed_0/a_388_n34# sky130_hilas_pFETmed_4/a_440_n8# sky130_hilas_pFETmed
Xsky130_hilas_pFETmed_2 VSUBS sky130_hilas_pFETmed_3/a_330_n8# sky130_hilas_pFETmed_4/w_294_n44#
+ sky130_hilas_pFETmed_2/a_388_n34# sky130_hilas_pFETmed_2/a_330_n8# sky130_hilas_pFETmed
Xsky130_hilas_pFETmed_1 VSUBS sky130_hilas_pFETmed_2/a_330_n8# sky130_hilas_pFETmed_4/w_294_n44#
+ sky130_hilas_pFETmed_1/a_388_n34# sky130_hilas_pFETmed_1/a_330_n8# sky130_hilas_pFETmed
Xsky130_hilas_pFETmed_3 VSUBS sky130_hilas_pFETmed_3/a_440_n8# sky130_hilas_pFETmed_4/w_294_n44#
+ sky130_hilas_pFETmed_3/a_388_n34# sky130_hilas_pFETmed_3/a_330_n8# sky130_hilas_pFETmed
Xsky130_hilas_pFETmed_4 VSUBS sky130_hilas_pFETmed_4/a_440_n8# sky130_hilas_pFETmed_4/w_294_n44#
+ sky130_hilas_pFETmed_4/a_388_n34# sky130_hilas_pFETmed_4/a_330_n8# sky130_hilas_pFETmed
.ends

.subckt sky130_hilas_pFETLarge GATE SOURCE DRAIN WELL
Xsky130_hilas_pFETLargePart1_0 VSUBS GATE SOURCE GATE GATE SOURCE DRAIN SOURCE DRAIN
+ GATE WELL GATE DRAIN sky130_hilas_pFETLargePart1
Xsky130_hilas_pFETLargePart1_1 VSUBS GATE SOURCE GATE GATE SOURCE DRAIN SOURCE DRAIN
+ GATE WELL GATE DRAIN sky130_hilas_pFETLargePart1
.ends

