magic
tech sky130A
timestamp 1628707355
<< checkpaint >>
rect -621 1197 2278 1429
rect -621 -454 2288 1197
rect -593 -628 2288 -454
rect -329 -631 2081 -628
<< error_s >>
rect 99 544 138 547
rect 260 544 299 547
rect 421 544 460 547
rect 582 544 621 547
rect 743 544 782 547
rect 904 544 943 547
rect 1065 544 1104 547
rect 1226 544 1265 547
rect 1387 544 1426 547
rect 1548 544 1587 547
rect 99 502 138 505
rect 260 502 299 505
rect 421 502 460 505
rect 582 502 621 505
rect 743 502 782 505
rect 904 502 943 505
rect 1065 502 1104 505
rect 1226 502 1265 505
rect 1387 502 1426 505
rect 1548 502 1587 505
rect 99 448 138 451
rect 259 448 298 451
rect 420 448 459 451
rect 581 448 620 451
rect 742 448 781 451
rect 903 448 942 451
rect 1064 448 1103 451
rect 1225 448 1264 451
rect 1386 448 1425 451
rect 1548 448 1587 451
rect 99 406 138 409
rect 259 406 298 409
rect 420 406 459 409
rect 581 406 620 409
rect 742 406 781 409
rect 903 406 942 409
rect 1064 406 1103 409
rect 1225 406 1264 409
rect 1386 406 1425 409
rect 1548 406 1587 409
rect 99 352 138 355
rect 259 352 298 355
rect 420 352 459 355
rect 581 352 620 355
rect 742 352 781 355
rect 903 352 942 355
rect 1064 352 1103 355
rect 1225 352 1264 355
rect 1386 352 1425 355
rect 1548 352 1587 355
rect 99 310 138 313
rect 259 310 298 313
rect 420 310 459 313
rect 581 310 620 313
rect 742 310 781 313
rect 903 310 942 313
rect 1064 310 1103 313
rect 1225 310 1264 313
rect 1386 310 1425 313
rect 1548 310 1587 313
rect 853 290 854 294
rect 99 256 138 259
rect 259 256 298 259
rect 420 256 459 259
rect 581 256 620 259
rect 742 256 781 259
rect 903 256 942 259
rect 1064 256 1103 259
rect 1225 256 1264 259
rect 1386 256 1425 259
rect 1548 256 1587 259
rect 99 214 138 217
rect 259 214 298 217
rect 420 214 459 217
rect 581 214 620 217
rect 742 214 781 217
rect 903 214 942 217
rect 1064 214 1103 217
rect 1225 214 1264 217
rect 1386 214 1425 217
rect 1548 214 1587 217
rect 99 160 138 163
rect 259 160 298 163
rect 420 160 459 163
rect 581 160 620 163
rect 742 160 781 163
rect 903 160 942 163
rect 1064 160 1103 163
rect 1225 160 1264 163
rect 1386 160 1425 163
rect 1548 160 1587 163
rect 99 118 138 121
rect 259 118 298 121
rect 420 118 459 121
rect 581 118 620 121
rect 742 118 781 121
rect 903 118 942 121
rect 1064 118 1103 121
rect 1225 118 1264 121
rect 1386 118 1425 121
rect 1548 118 1587 121
rect 99 64 138 67
rect 260 64 299 67
rect 421 64 460 67
rect 582 64 621 67
rect 743 64 782 67
rect 904 64 943 67
rect 1065 64 1104 67
rect 1226 64 1265 67
rect 1387 64 1426 67
rect 1548 64 1587 67
rect 99 22 138 25
rect 260 22 299 25
rect 421 22 460 25
rect 582 22 621 25
rect 743 22 782 25
rect 904 22 943 25
rect 1065 22 1104 25
rect 1226 22 1265 25
rect 1387 22 1426 25
rect 1548 22 1587 25
<< nwell >>
rect 237 495 1380 502
<< poly >>
rect 198 557 224 560
rect 520 557 546 560
rect 681 557 707 561
rect 842 557 868 560
rect 1003 557 1029 562
rect 1164 557 1190 561
<< locali >>
rect 398 502 415 503
rect 1295 502 1316 580
rect 1362 502 1379 570
rect 237 479 1380 502
rect 237 123 254 479
rect 303 0 320 446
rect 398 123 415 479
rect 466 0 483 442
rect 557 123 574 479
rect 626 0 643 450
rect 719 123 736 479
rect 788 0 805 445
rect 881 125 898 479
rect 948 0 965 450
rect 1041 126 1058 479
rect 1110 0 1127 450
rect 1202 125 1219 479
rect 1270 0 1287 448
rect 1363 122 1380 479
rect 1431 0 1448 466
<< metal1 >>
rect 674 355 1019 372
rect 829 102 847 256
rect 999 171 1019 355
rect 304 0 1658 23
<< metal2 >>
rect 0 577 705 596
rect 0 575 29 577
rect 0 495 206 501
rect 348 495 370 541
rect 840 496 865 572
rect 840 495 868 496
rect 0 480 868 495
rect 26 456 46 480
rect 190 465 868 480
rect 1011 308 1031 568
rect 0 287 1031 308
rect 1171 210 1186 584
rect 1271 568 1387 596
rect 1346 567 1387 568
rect 0 190 1187 210
rect 0 189 14 190
rect 0 78 854 98
use sky130_hilas_DAC6TransistorStack01a  sky130_hilas_DAC6TransistorStack01a_0
timestamp 1628707318
transform 1 0 9 0 1 176
box 0 0 190 623
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_8
timestamp 1628707353
transform 1 0 202 0 1 568
box 0 0 33 55
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_10
timestamp 1628707353
transform 1 0 29 0 1 433
box 0 0 33 55
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_12
timestamp 1628707353
transform 1 0 31 0 1 244
box 0 0 33 55
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_11
timestamp 1628707353
transform 1 0 31 0 1 338
box 0 0 33 55
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_9
timestamp 1628707353
transform 1 0 31 0 1 564
box 0 0 33 55
use sky130_hilas_li2m1  sky130_hilas_li2m1_6
timestamp 1628707287
transform 1 0 473 0 1 7
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1628707287
transform 1 0 311 0 1 7
box 0 0 23 29
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_6
timestamp 1628707353
transform 1 0 522 0 1 568
box 0 0 33 55
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_7
timestamp 1628707353
transform 0 1 352 -1 0 548
box 0 0 33 55
use sky130_hilas_DAC6TransistorStack01  sky130_hilas_DAC6TransistorStack01_0
array 0 2 161 0 0 566
timestamp 1628707266
transform 1 0 170 0 1 176
box 0 0 191 623
use sky130_hilas_li2m1  sky130_hilas_li2m1_7
timestamp 1628707287
transform 1 0 633 0 1 7
box 0 0 23 29
use sky130_hilas_DAC6TransistorStack01b  sky130_hilas_DAC6TransistorStack01b_0
timestamp 1628707317
transform 1 0 653 0 1 176
box 0 0 209 623
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_5
timestamp 1628707353
transform 1 0 683 0 1 569
box 0 0 33 55
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1628707287
transform 1 0 795 0 1 7
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_5
timestamp 1628707287
transform 1 0 955 0 1 7
box 0 0 23 29
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1628707321
transform 1 0 835 0 1 82
box 0 0 32 32
use sky130_hilas_DAC6TransistorStack01c  sky130_hilas_DAC6TransistorStack01c_0
timestamp 1628707348
transform 1 0 814 0 1 176
box 0 0 206 623
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_4
timestamp 1628707353
transform 1 0 845 0 1 568
box 0 0 33 55
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_3
timestamp 1628707353
transform 1 0 1006 0 1 569
box 0 0 33 55
use sky130_hilas_DAC6TransistorStack01  sky130_hilas_DAC6TransistorStack01_2
array 0 2 161 0 0 566
timestamp 1628707266
transform 1 0 975 0 1 176
box 0 0 191 623
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_2
timestamp 1628707353
transform 1 0 1167 0 1 569
box 0 0 33 55
use sky130_hilas_DAC6TransistorStack01a  sky130_hilas_DAC6TransistorStack01a_1
timestamp 1628707318
transform 1 0 1458 0 1 176
box 0 0 190 623
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628707307
transform 1 0 1297 0 1 565
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628707307
transform 1 0 1364 0 1 565
box 0 0 34 33
use sky130_hilas_li2m1  sky130_hilas_li2m1_3
timestamp 1628707287
transform 1 0 1277 0 1 7
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_4
timestamp 1628707287
transform 1 0 1438 0 1 7
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_2
timestamp 1628707287
transform 1 0 1117 0 1 7
box 0 0 23 29
<< labels >>
rlabel metal2 1 575 11 596 0 A4
port 5 nsew analog default
rlabel metal2 0 480 10 501 0 A3
port 4 nsew analog default
rlabel metal2 1 287 11 308 0 A2
port 3 nsew analog default
rlabel metal2 1 189 11 210 0 A1
port 2 nsew analog default
rlabel metal2 0 78 8 98 0 A0
port 1 nsew analog default
rlabel metal2 1271 582 1346 596 0 VPWR
port 6 nsew analog default
rlabel metal1 1646 0 1658 23 0 OUT
port 7 nsew analog default
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
