magic
tech sky130A
timestamp 1634057839
<< checkpaint >>
rect -630 1190 867 1223
rect -630 951 1023 1190
rect -630 -324 1044 951
rect -531 -342 1044 -324
rect -531 -396 1043 -342
rect -531 -397 1019 -396
rect -512 -445 1019 -397
rect -462 -575 1019 -445
rect -453 -610 1019 -575
rect -340 -619 1019 -610
<< nwell >>
rect 384 304 440 501
<< psubdiff >>
rect 393 153 422 182
rect 393 136 399 153
rect 416 136 422 153
rect 393 119 422 136
rect 393 102 399 119
rect 416 102 422 119
rect 393 89 422 102
<< nsubdiff >>
rect 394 417 422 429
rect 394 400 398 417
rect 415 400 422 417
rect 394 383 422 400
rect 394 366 398 383
rect 415 366 422 383
rect 394 337 422 366
<< psubdiffcont >>
rect 399 136 416 153
rect 399 102 416 119
<< nsubdiffcont >>
rect 398 400 415 417
rect 398 366 415 383
<< poly >>
rect 141 279 220 294
rect 312 279 391 294
rect 140 243 219 258
rect 312 243 391 258
<< locali >>
rect 398 417 415 425
rect 398 358 415 366
rect 399 119 416 136
<< viali >>
rect 398 383 415 400
rect 399 153 416 170
rect 399 85 416 102
<< metal1 >>
rect 392 407 419 424
rect 390 404 422 407
rect 390 378 393 404
rect 419 378 422 404
rect 390 375 422 378
rect 392 357 419 375
rect 439 230 440 253
rect 393 170 422 173
rect 393 153 399 170
rect 416 153 422 170
rect 393 142 422 153
rect 393 116 395 142
rect 421 116 422 142
rect 393 102 422 116
rect 393 85 399 102
rect 416 85 422 102
rect 393 82 422 85
<< via1 >>
rect 393 400 419 404
rect 393 383 398 400
rect 398 383 415 400
rect 415 383 419 400
rect 393 378 419 383
rect 395 116 421 142
<< metal2 >>
rect 87 511 283 533
rect 372 519 440 540
rect 87 434 162 455
rect 257 436 440 457
rect 87 433 114 434
rect 390 404 422 407
rect 390 378 393 404
rect 419 401 422 404
rect 419 380 440 401
rect 419 378 422 380
rect 390 375 422 378
rect 87 334 112 356
rect 87 278 385 299
rect 87 238 385 259
rect 87 180 112 202
rect 392 142 424 145
rect 392 116 395 142
rect 421 140 424 142
rect 421 119 440 140
rect 421 116 424 119
rect 392 113 424 116
rect 87 45 158 66
rect 253 47 440 69
rect 87 0 286 22
rect 371 3 440 24
use sky130_hilas_poly2m1  sky130_hilas_poly2m1_0
timestamp 1634057706
transform 1 0 118 0 -1 304
box 0 0 33 51
use sky130_hilas_poly2m1  sky130_hilas_poly2m1_1
timestamp 1634057706
transform -1 0 132 0 1 233
box 0 0 33 51
use sky130_hilas_nFETmed  sky130_hilas_nFETmed_1
timestamp 1634057737
transform 1 0 177 0 1 20
box 0 0 82 272
use sky130_hilas_nFETmed  sky130_hilas_nFETmed_0
timestamp 1634057737
transform 1 0 296 0 1 20
box 0 0 82 272
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_0
timestamp 1634057713
transform 0 -1 413 1 0 234
box 0 0 33 55
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_1
timestamp 1634057713
transform 0 -1 414 1 0 288
box 0 0 33 55
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_1
timestamp 1634057714
transform 1 0 118 0 1 306
box 0 0 119 287
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_0
timestamp 1634057714
transform 1 0 0 0 1 306
box 0 0 119 287
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1634057711
transform 1 0 118 0 1 185
box 0 0 32 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1634057711
transform 1 0 118 0 1 340
box 0 0 32 32
use sky130_hilas_li2m2  sky130_hilas_li2m2_4
timestamp 1634057699
transform 1 0 168 0 1 55
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_5
timestamp 1634057699
transform 1 0 238 0 1 55
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_7
timestamp 1634057699
transform 1 0 290 0 1 11
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_6
timestamp 1634057699
transform 1 0 355 0 1 11
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1634057699
transform 1 0 171 0 1 443
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1634057699
transform 1 0 288 0 1 521
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1634057699
transform 1 0 240 0 1 444
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1634057699
transform 1 0 359 0 1 527
box 0 0 34 33
<< labels >>
rlabel metal2 87 334 96 356 0 GATE1P
port 3 nsew analog default
rlabel metal2 87 278 95 299 0 GATE2P
port 2 nsew analog default
rlabel metal2 87 238 95 259 0 GATE2N
port 4 nsew analog default
rlabel metal2 87 181 95 202 0 GATE1N
port 1 nsew analog default
rlabel metal2 430 519 440 540 0 DRAIN2P
port 12 nsew analog default
rlabel metal2 430 436 440 457 0 DRAIN1P
port 11 nsew analog default
rlabel metal2 87 433 95 455 0 SOURCE1P
port 5 nsew analog default
rlabel metal2 87 511 95 533 0 SOURCE2P
port 6 nsew analog default
rlabel metal2 87 45 94 66 0 SOURCE1N
port 8 nsew analog default
rlabel metal2 87 0 94 22 0 SOURCE2N
port 7 nsew analog default
rlabel metal2 433 47 440 69 0 DRAIN1N
port 9 nsew analog default
rlabel metal2 433 3 440 24 0 DRAIN2N
port 10 nsew analog default
rlabel metal2 429 119 440 140 0 VGND
port 14 nsew
rlabel metal2 431 380 440 401 0 WELL
port 15 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
