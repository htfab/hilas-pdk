magic
tech sky130A
timestamp 1628707319
<< nmos >>
rect 8 15 14 18
<< pmos >>
rect 39 15 45 18
<< ndiff >>
rect 8 24 14 25
rect 8 20 9 24
rect 13 20 14 24
rect 8 18 14 20
rect 8 13 14 15
rect 8 9 9 13
rect 13 9 14 13
rect 8 8 14 9
<< pdiff >>
rect 39 25 45 26
rect 39 21 40 25
rect 44 21 45 25
rect 39 18 45 21
rect 39 12 45 15
rect 39 8 40 12
rect 44 8 45 12
rect 39 7 45 8
<< ndiffc >>
rect 9 20 13 24
rect 9 9 13 13
<< pdiffc >>
rect 40 21 44 25
rect 40 8 44 12
<< poly >>
rect 5 15 8 18
rect 14 15 39 18
rect 45 15 47 18
rect 24 12 27 15
rect 22 11 28 12
rect 22 7 23 11
rect 27 7 28 11
rect 22 6 28 7
<< metal1 >>
rect 23 24 27 31
rect 13 21 40 24
rect 13 20 44 21
rect 5 9 9 13
rect 44 8 47 12
rect 23 0 27 7
<< via1 >>
rect 1 9 5 13
rect 47 8 51 12
<< metal2 >>
rect 0 13 6 30
rect 0 9 1 13
rect 5 9 6 13
rect 0 3 6 9
rect 46 12 52 30
rect 46 8 47 12
rect 51 8 52 12
rect 46 3 52 8
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
