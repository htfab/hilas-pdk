magic
tech sky130A
timestamp 1632151084
<< mvnmos >>
rect 1679 316 1729 556
rect 1679 40 1729 280
<< mvndiff >>
rect 1650 551 1679 556
rect 1650 336 1656 551
rect 1673 336 1679 551
rect 1650 316 1679 336
rect 1729 550 1766 556
rect 1729 336 1735 550
rect 1752 345 1766 550
rect 1752 336 1778 345
rect 1729 318 1778 336
rect 1729 316 1755 318
rect 1749 280 1755 316
rect 1650 260 1679 280
rect 1650 50 1656 260
rect 1673 50 1679 260
rect 1650 40 1679 50
rect 1729 277 1755 280
rect 1772 277 1778 318
rect 1729 260 1778 277
rect 1729 50 1735 260
rect 1752 251 1778 260
rect 1752 50 1766 251
rect 1729 40 1766 50
<< mvndiffc >>
rect 1656 336 1673 551
rect 1735 336 1752 550
rect 1656 50 1673 260
rect 1755 277 1772 318
rect 1735 50 1752 260
<< psubdiff >>
rect 1766 537 1809 556
rect 1766 361 1779 537
rect 1797 361 1809 537
rect 1766 345 1809 361
rect 1766 244 1809 251
rect 1766 52 1779 244
rect 1797 52 1809 244
rect 1766 40 1809 52
<< psubdiffcont >>
rect 1779 361 1797 537
rect 1779 52 1797 244
<< poly >>
rect 1183 575 1270 597
rect 1183 29 1216 31
rect 1183 12 1191 29
rect 1208 12 1216 29
rect 1183 7 1216 12
rect 1292 575 1380 597
rect 1237 7 1325 31
rect 1402 575 1490 597
rect 1347 7 1435 31
rect 1512 575 1600 597
rect 1457 7 1545 31
rect 1679 592 1729 597
rect 1679 575 1695 592
rect 1712 575 1729 592
rect 1679 556 1729 575
rect 1679 280 1729 316
rect 1567 29 1600 31
rect 1567 12 1575 29
rect 1592 12 1600 29
rect 1567 7 1600 12
rect 1679 7 1729 40
<< polycont >>
rect 1191 12 1208 29
rect 1695 575 1712 592
rect 1575 12 1592 29
<< npolyres >>
rect 1183 31 1216 575
rect 1237 31 1270 575
rect 1292 31 1325 575
rect 1347 31 1380 575
rect 1402 31 1435 575
rect 1457 31 1490 575
rect 1512 31 1545 575
rect 1567 31 1600 575
<< locali >>
rect 1627 575 1695 592
rect 1712 575 1720 592
rect 1627 551 1675 575
rect 1627 546 1656 551
rect 1627 336 1631 546
rect 1649 336 1656 546
rect 1673 336 1675 551
rect 1627 328 1675 336
rect 1733 550 1797 558
rect 1733 336 1735 550
rect 1752 537 1797 550
rect 1752 361 1779 537
rect 1752 336 1797 361
rect 1733 318 1797 336
rect 1733 277 1755 318
rect 1772 277 1797 318
rect 1624 260 1675 268
rect 1537 76 1573 86
rect 1537 59 1548 76
rect 1565 59 1573 76
rect 1537 48 1573 59
rect 1162 29 1216 30
rect 1162 28 1191 29
rect 1162 11 1165 28
rect 1182 12 1191 28
rect 1208 12 1216 29
rect 1547 29 1573 48
rect 1624 50 1631 260
rect 1649 50 1656 260
rect 1673 50 1675 260
rect 1624 43 1675 50
rect 1654 42 1675 43
rect 1733 260 1797 277
rect 1733 50 1735 260
rect 1752 244 1797 260
rect 1752 107 1779 244
rect 1752 90 1760 107
rect 1777 90 1779 107
rect 1752 70 1779 90
rect 1752 53 1760 70
rect 1777 53 1779 70
rect 1752 52 1779 53
rect 1752 50 1797 52
rect 1733 43 1797 50
rect 1733 42 1784 43
rect 1752 33 1784 42
rect 1547 12 1575 29
rect 1592 12 1600 29
rect 1752 16 1760 33
rect 1777 16 1784 33
rect 1752 13 1784 16
rect 1182 11 1216 12
rect 1162 8 1216 11
<< viali >>
rect 1631 336 1649 546
rect 1548 59 1565 76
rect 1165 11 1182 28
rect 1631 50 1649 260
rect 1760 90 1777 107
rect 1760 53 1777 70
rect 1760 16 1777 33
<< metal1 >>
rect 1625 546 1665 553
rect 1625 539 1631 546
rect 1649 539 1665 546
rect 1625 345 1630 539
rect 1659 345 1665 539
rect 1625 336 1631 345
rect 1649 336 1665 345
rect 1625 332 1665 336
rect 1155 323 1181 326
rect 1155 294 1181 297
rect 1159 45 1180 294
rect 1626 261 1657 266
rect 1626 260 1669 261
rect 1537 82 1573 86
rect 1537 56 1543 82
rect 1569 56 1573 82
rect 1537 48 1573 56
rect 1626 50 1631 260
rect 1649 254 1669 260
rect 1663 144 1669 254
rect 1649 50 1669 144
rect 1626 49 1669 50
rect 1750 107 1786 110
rect 1750 90 1760 107
rect 1777 90 1786 107
rect 1750 70 1786 90
rect 1750 53 1760 70
rect 1777 53 1786 70
rect 1159 39 1181 45
rect 1626 44 1657 49
rect 1159 31 1184 39
rect 1750 33 1786 53
rect 1159 28 1188 31
rect 1159 11 1165 28
rect 1182 11 1188 28
rect 1159 8 1188 11
rect 1750 21 1760 33
rect 1777 21 1786 33
rect 1750 -5 1755 21
rect 1781 -5 1786 21
rect 1750 -10 1786 -5
<< via1 >>
rect 1630 345 1631 539
rect 1631 345 1649 539
rect 1649 345 1659 539
rect 1155 297 1181 323
rect 1543 76 1569 82
rect 1543 59 1548 76
rect 1548 59 1565 76
rect 1565 59 1569 76
rect 1543 56 1569 59
rect 1637 144 1649 254
rect 1649 144 1663 254
rect 1755 16 1760 21
rect 1760 16 1777 21
rect 1777 16 1781 21
rect 1755 -5 1781 16
<< metal2 >>
rect 1627 539 1661 544
rect 1627 415 1630 539
rect 1128 396 1630 415
rect 1627 345 1630 396
rect 1659 395 1661 539
rect 1659 369 1833 395
rect 1659 345 1661 369
rect 1627 335 1661 345
rect 1154 323 1182 327
rect 1152 321 1155 323
rect 1124 298 1155 321
rect 1152 297 1155 298
rect 1181 297 1184 323
rect 1154 293 1182 297
rect 1626 254 1670 268
rect 1626 229 1637 254
rect 1128 210 1637 229
rect 1626 144 1637 210
rect 1663 237 1670 254
rect 1663 211 1833 237
rect 1663 210 1712 211
rect 1663 144 1670 210
rect 1626 141 1670 144
rect 1539 82 1573 86
rect 1539 56 1543 82
rect 1569 81 1573 82
rect 1569 56 1833 81
rect 1539 55 1833 56
rect 1539 52 1573 55
rect 1642 21 1833 29
rect 1642 -5 1755 21
rect 1781 -5 1833 21
rect 1642 -11 1833 -5
use sky130_hilas_FGtrans2x1cell2  sky130_hilas_FGtrans2x1cell2_0
timestamp 1631886322
transform -1 0 752 0 -1 229
box -395 -387 757 228
<< labels >>
rlabel metal2 1820 369 1833 395 0 NBIAS
port 1 nsew
rlabel metal2 1821 211 1833 237 0 PBIAS
port 2 nsew
rlabel metal2 1823 -11 1833 29 0 VGND
port 3 nsew
rlabel metal2 1823 55 1833 81 0 RESIST
port 4 nsew
<< end >>
