magic
tech sky130A
timestamp 1629137192
<< checkpaint >>
rect -652 -635 1176 1240
<< metal2 >>
rect 35 554 108 555
rect 35 538 177 554
rect 35 537 108 538
rect 35 367 102 369
rect 35 351 174 367
rect 35 252 105 253
rect 35 236 178 252
rect 35 52 181 69
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_0
timestamp 1628285143
transform 1 0 210 0 1 333
box -232 -45 336 125
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_3
timestamp 1628285143
transform 1 0 210 0 -1 272
box -232 -45 336 125
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_1
timestamp 1628285143
transform 1 0 210 0 -1 565
box -232 -45 336 125
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_2
timestamp 1628285143
transform 1 0 210 0 1 40
box -232 -45 336 125
<< labels >>
rlabel metal2 35 537 40 555 0 drain1
rlabel metal2 35 351 40 369 0 drain2
rlabel metal2 35 236 40 253 0 drain3
rlabel metal2 35 52 40 69 0 drain4
<< end >>
