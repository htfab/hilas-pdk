magic
tech sky130A
timestamp 1628704292
<< error_s >>
rect 307 540 308 543
rect 307 389 308 392
rect 307 238 308 241
rect 839 171 891 172
rect 1049 171 1099 172
<< nwell >>
rect 669 605 691 611
rect 669 10 691 15
<< metal1 >>
rect 61 604 83 612
rect 318 603 341 612
rect 367 577 394 606
rect 669 605 691 611
rect 1166 607 1193 612
rect 363 550 366 577
rect 393 550 396 577
rect 459 558 486 563
rect 367 472 394 550
rect 366 469 394 472
rect 393 442 394 469
rect 366 439 394 442
rect 367 436 394 439
rect 413 509 440 516
rect 413 304 440 482
rect 459 417 486 531
rect 554 513 583 518
rect 552 510 583 513
rect 581 481 583 510
rect 552 478 583 481
rect 454 390 457 417
rect 484 390 487 417
rect 412 301 440 304
rect 439 274 440 301
rect 412 271 440 274
rect 413 154 440 271
rect 459 259 486 390
rect 457 256 486 259
rect 484 229 486 256
rect 457 226 486 229
rect 459 224 486 226
rect 506 363 533 369
rect 506 360 534 363
rect 506 333 507 360
rect 506 330 534 333
rect 554 356 583 478
rect 554 330 556 356
rect 582 330 583 356
rect 413 151 443 154
rect 413 124 416 151
rect 413 121 443 124
rect 413 116 440 121
rect 506 109 533 330
rect 504 106 533 109
rect 531 79 533 106
rect 504 76 533 79
rect 506 73 533 76
rect 554 213 583 330
rect 554 210 584 213
rect 554 181 555 210
rect 554 178 584 181
rect 554 56 583 178
rect 554 24 583 27
rect 669 10 691 15
rect 1166 10 1193 15
<< via1 >>
rect 366 550 393 577
rect 459 531 486 558
rect 366 442 393 469
rect 413 482 440 509
rect 552 481 581 510
rect 457 390 484 417
rect 412 274 439 301
rect 457 229 484 256
rect 507 333 534 360
rect 556 330 582 356
rect 416 124 443 151
rect 504 79 531 106
rect 555 181 584 210
rect 554 27 583 56
<< metal2 >>
rect 371 596 608 597
rect 369 581 608 596
rect 369 580 396 581
rect 366 577 396 580
rect 0 555 11 573
rect 343 555 366 573
rect 393 555 396 577
rect 366 547 393 550
rect 456 531 459 558
rect 486 552 489 558
rect 486 536 608 552
rect 486 531 489 536
rect 410 506 413 509
rect 343 488 413 506
rect 410 482 413 488
rect 440 506 443 509
rect 440 487 445 506
rect 440 482 443 487
rect 549 481 552 510
rect 581 503 584 510
rect 581 487 608 503
rect 581 481 584 487
rect 1282 483 1295 500
rect 363 442 366 469
rect 393 463 396 469
rect 393 447 527 463
rect 393 442 396 447
rect 511 446 527 447
rect 511 430 607 446
rect 0 404 11 422
rect 343 420 479 422
rect 343 417 484 420
rect 343 404 457 417
rect 484 390 485 401
rect 457 387 485 390
rect 462 385 485 387
rect 512 385 608 401
rect 512 360 528 385
rect 504 355 507 360
rect 343 337 507 355
rect 504 333 507 337
rect 534 333 537 360
rect 553 330 556 356
rect 582 352 585 356
rect 582 336 608 352
rect 582 330 585 336
rect 1282 332 1295 349
rect 409 274 412 301
rect 439 295 442 301
rect 439 279 608 295
rect 439 274 442 279
rect 0 253 11 271
rect 454 229 457 256
rect 484 250 487 256
rect 484 234 608 250
rect 484 229 487 234
rect 552 204 555 210
rect 343 186 555 204
rect 552 181 555 186
rect 584 204 587 210
rect 584 201 601 204
rect 584 185 608 201
rect 584 181 587 185
rect 1282 181 1295 198
rect 413 124 416 151
rect 443 145 446 151
rect 443 129 608 145
rect 443 124 446 129
rect 501 79 504 106
rect 531 100 534 106
rect 531 84 608 100
rect 531 79 534 84
rect 551 27 554 56
rect 583 51 586 56
rect 583 35 608 51
rect 583 27 586 35
rect 1282 31 1295 48
use sky130_hilas_VinjNOR3  VinjNOR3_2
timestamp 1624138502
transform 1 0 944 0 1 157
box -337 144 351 308
use sky130_hilas_VinjNOR3  VinjNOR3_1
timestamp 1624138502
transform 1 0 944 0 1 6
box -337 144 351 308
use sky130_hilas_VinjNOR3  VinjNOR3_3
timestamp 1624138502
transform 1 0 944 0 1 308
box -337 144 351 308
use sky130_hilas_VinjNOR3  VinjNOR3_0
timestamp 1624138502
transform 1 0 944 0 1 -144
box -337 144 351 308
use sky130_hilas_VinjInv2  VinjInv2_0
timestamp 1624141468
transform 1 0 336 0 1 308
box -336 144 25 308
use sky130_hilas_VinjInv2  VinjInv2_1
timestamp 1624141468
transform 1 0 336 0 1 157
box -336 144 25 308
use sky130_hilas_VinjInv2  VinjInv2_2
timestamp 1624141468
transform 1 0 336 0 1 6
box -336 144 25 308
<< labels >>
rlabel metal2 1282 483 1295 500 0 OUTPUT00
port 1 nsew
rlabel metal2 1282 332 1295 349 0 OUTPUT01
port 2 nsew
rlabel metal2 1282 181 1295 198 0 OUTPUT10
port 3 nsew
rlabel metal2 1282 31 1295 48 0 OUTPUT11
port 4 nsew
rlabel metal1 1166 607 1193 612 0 VGND
port 5 nsew
rlabel metal1 1166 10 1193 15 0 VGND
port 5 nsew
rlabel metal1 669 10 691 15 0 VINJ
port 6 nsew
rlabel metal1 669 605 691 611 0 VINJ
port 6 nsew
rlabel metal2 0 555 11 573 0 IN1
port 8 nsew
rlabel metal2 0 404 11 422 0 IN2
port 7 nsew
rlabel metal2 0 253 11 271 0 ENABLE
port 9 nsew
rlabel metal1 61 604 83 612 0 VINJ
port 6 nsew
rlabel metal1 318 603 341 612 0 VGND
port 5 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
