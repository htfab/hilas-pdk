magic
tech sky130A
timestamp 1606955279
<< error_s >>
rect -338 150 -332 156
rect -285 150 -279 156
rect -344 100 -338 106
rect -279 100 -273 106
rect 85 91 91 97
rect 190 91 196 97
rect 79 41 85 47
rect 196 41 202 47
rect 364 -188 379 -187
rect 453 -188 466 -187
rect 85 -210 91 -204
rect 190 -210 196 -204
rect -338 -265 -332 -259
rect -285 -265 -279 -259
rect 79 -260 85 -254
rect 196 -260 202 -254
rect -344 -315 -338 -309
rect -279 -315 -273 -309
rect 514 -314 524 -313
<< nwell >>
rect 9 24 10 27
rect -337 -242 -281 0
rect 7 -11 39 24
<< psubdiff >>
rect -95 -42 -70 121
rect -95 -59 -92 -42
rect -73 -59 -70 -42
rect -95 -72 -70 -59
rect -95 -75 268 -72
rect -95 -76 146 -75
rect -95 -93 -71 -76
rect -52 -93 -28 -76
rect -9 -93 16 -76
rect 35 -93 56 -76
rect 75 -93 100 -76
rect 119 -92 146 -76
rect 165 -76 268 -75
rect 165 -92 190 -76
rect 119 -93 190 -92
rect 209 -93 236 -76
rect 255 -93 268 -76
rect -95 -97 268 -93
rect -95 -110 -70 -97
rect -95 -127 -92 -110
rect -73 -127 -70 -110
rect -95 -281 -70 -127
<< mvnsubdiff >>
rect -337 -242 -281 0
<< psubdiffcont >>
rect -92 -59 -73 -42
rect -71 -93 -52 -76
rect -28 -93 -9 -76
rect 16 -93 35 -76
rect 56 -93 75 -76
rect 100 -93 119 -76
rect 146 -92 165 -75
rect 190 -93 209 -76
rect 236 -93 255 -76
rect -92 -127 -73 -110
<< poly >>
rect -237 134 331 151
rect -237 126 -185 134
rect 45 91 64 134
rect 220 90 237 134
rect 276 52 319 102
rect 276 -210 291 52
rect 381 -131 398 -27
rect 276 -233 316 -210
rect 272 -238 316 -233
rect 272 -255 280 -238
rect 297 -255 316 -238
rect 272 -260 316 -255
rect 46 -293 63 -260
rect 220 -293 237 -260
rect 272 -263 300 -260
rect -280 -310 331 -293
<< polycont >>
rect 280 -255 297 -238
<< locali >>
rect 362 28 470 45
rect -92 -42 -73 -34
rect 464 -51 472 -34
rect -92 -75 -73 -59
rect -92 -76 146 -75
rect -92 -93 -71 -76
rect -52 -93 -28 -76
rect -9 -93 16 -76
rect 35 -93 56 -76
rect 75 -93 100 -76
rect 119 -92 146 -76
rect 165 -76 263 -75
rect 165 -92 190 -76
rect 119 -93 190 -92
rect 209 -93 236 -76
rect 255 -93 263 -76
rect -92 -110 -73 -93
rect 338 -108 355 -51
rect 474 -108 491 -51
rect 361 -125 363 -124
rect 464 -125 469 -108
rect -92 -135 -73 -127
rect 362 -205 470 -188
rect 280 -236 297 -230
rect 280 -264 297 -257
<< viali >>
rect 278 -238 299 -236
rect 278 -255 280 -238
rect 280 -255 297 -238
rect 297 -255 299 -238
rect 278 -257 299 -255
<< metal1 >>
rect -361 -382 -319 223
rect 9 25 10 27
rect 9 24 34 25
rect 9 18 39 24
rect 9 -8 12 18
rect 38 -8 39 18
rect 9 -11 39 -8
rect 279 -230 297 223
rect 274 -236 303 -230
rect 274 -257 278 -236
rect 299 -257 303 -236
rect 274 -264 303 -257
rect 279 -383 297 -264
<< via1 >>
rect 12 -8 38 18
<< metal2 >>
rect 484 173 516 175
rect -396 155 516 173
rect 7 19 38 24
rect -255 18 269 19
rect -255 0 12 18
rect 7 -8 12 0
rect 38 0 269 18
rect 7 -11 38 -8
rect 510 -315 514 -313
rect -394 -330 514 -315
use TunCap01  TunCap01_3
timestamp 1606740587
transform 1 0 1056 0 1 433
box -1451 -400 -1278 -210
use wellContact  wellContact_1
timestamp 1606753443
transform 1 0 1054 0 1 404
box -1449 -441 -1275 -255
use wellContact  wellContact_0
timestamp 1606753443
transform 1 0 1054 0 1 231
box -1449 -441 -1275 -255
use TunCap01  TunCap01_1
timestamp 1606740587
transform 1 0 1056 0 1 18
box -1451 -400 -1278 -210
use horizTransCell01  horizTransCell01_0
timestamp 1606869277
transform 1 0 790 0 1 -429
box -476 47 -33 359
use horizTransCell01  horizTransCell01_1
timestamp 1606869277
transform 1 0 790 0 -1 270
box -476 47 -33 359
use FGVaractorCapacitor02  FGVaractorCapacitor02_0
timestamp 1606868103
transform 1 0 986 0 1 62
box -1005 -380 -733 -211
use FGVaractorCapacitor02  FGVaractorCapacitor02_2
timestamp 1606868103
transform 1 0 986 0 -1 -231
box -1005 -380 -733 -211
<< end >>
