magic
tech sky130A
timestamp 1628616696
<< checkpaint >>
rect -630 2577 1354 3031
rect -630 2331 1487 2577
rect -630 708 1811 2331
rect -497 309 1811 708
rect -497 268 1643 309
rect -389 254 1643 268
rect -299 -176 1643 254
rect -299 -630 1510 -176
<< error_s >>
rect 873 1286 874 1287
<< nwell >>
rect 90 1502 281 1503
rect 90 942 650 1502
rect 850 1485 978 1503
rect 90 924 133 942
rect 90 901 161 924
rect 90 899 133 901
rect 850 898 978 917
<< nsubdiff >>
rect 109 1419 140 1456
rect 109 1402 115 1419
rect 132 1402 140 1419
rect 109 1385 140 1402
rect 109 1368 115 1385
rect 132 1368 140 1385
rect 109 1351 140 1368
rect 109 1334 115 1351
rect 132 1334 140 1351
rect 109 1317 140 1334
rect 109 1300 115 1317
rect 132 1300 140 1317
rect 109 1283 140 1300
rect 109 1266 115 1283
rect 132 1266 140 1283
rect 109 1251 140 1266
rect 108 1116 140 1149
rect 108 1099 116 1116
rect 133 1099 140 1116
rect 108 1082 140 1099
rect 108 1065 116 1082
rect 133 1065 140 1082
rect 108 1048 140 1065
rect 108 1031 116 1048
rect 133 1031 140 1048
rect 108 1014 140 1031
rect 108 997 116 1014
rect 133 997 140 1014
rect 108 980 140 997
rect 108 963 116 980
rect 133 963 140 980
rect 108 948 140 963
<< nsubdiffcont >>
rect 115 1402 132 1419
rect 115 1368 132 1385
rect 115 1334 132 1351
rect 115 1300 132 1317
rect 115 1266 132 1283
rect 116 1099 133 1116
rect 116 1065 133 1082
rect 116 1031 133 1048
rect 116 997 133 1014
rect 116 963 133 980
<< locali >>
rect 157 1455 191 1456
rect 132 1431 191 1455
rect 132 1382 174 1431
rect 855 1356 857 1373
rect 874 1356 880 1373
rect 855 1319 880 1356
rect 855 1303 876 1319
rect 855 1286 857 1303
rect 874 1286 876 1303
rect 855 1284 876 1286
rect 115 1249 132 1266
rect 116 955 133 963
<< viali >>
rect 115 1419 132 1436
rect 115 1385 132 1402
rect 174 1414 191 1431
rect 174 1380 191 1397
rect 115 1351 132 1368
rect 115 1317 132 1334
rect 115 1283 132 1300
rect 857 1356 874 1373
rect 857 1286 874 1303
rect 116 1116 133 1133
rect 116 1082 133 1099
rect 116 1048 133 1065
rect 116 1014 133 1031
rect 116 980 133 997
<< metal1 >>
rect 782 1489 816 1503
rect 849 1488 876 1503
rect 112 1456 165 1457
rect 112 1455 191 1456
rect 112 1449 194 1455
rect 112 1436 124 1449
rect 112 1419 115 1436
rect 183 1431 194 1449
rect 112 1402 124 1419
rect 191 1425 194 1431
rect 191 1414 197 1425
rect 112 1385 115 1402
rect 183 1397 197 1414
rect 112 1377 124 1385
rect 191 1396 197 1397
rect 191 1380 194 1396
rect 183 1377 194 1380
rect 112 1371 194 1377
rect 852 1373 884 1377
rect 112 1368 176 1371
rect 112 1351 115 1368
rect 132 1351 176 1368
rect 112 1334 176 1351
rect 112 1317 115 1334
rect 132 1317 176 1334
rect 112 1300 176 1317
rect 112 1283 115 1300
rect 132 1283 176 1300
rect 852 1287 853 1373
rect 879 1287 884 1373
rect 852 1286 857 1287
rect 874 1286 884 1287
rect 852 1285 884 1286
rect 855 1284 884 1285
rect 112 1133 176 1283
rect 112 1116 116 1133
rect 133 1116 176 1133
rect 112 1099 176 1116
rect 112 1082 116 1099
rect 133 1082 176 1099
rect 112 1065 176 1082
rect 112 1048 116 1065
rect 133 1048 176 1065
rect 112 1031 176 1048
rect 112 1014 116 1031
rect 133 1014 176 1031
rect 112 997 176 1014
rect 112 980 116 997
rect 133 980 176 997
rect 112 953 176 980
rect 134 952 176 953
rect 782 898 816 917
rect 849 898 876 919
<< via1 >>
rect 124 1436 183 1449
rect 124 1419 132 1436
rect 132 1431 183 1436
rect 132 1419 174 1431
rect 124 1414 174 1419
rect 174 1414 183 1431
rect 124 1402 183 1414
rect 124 1385 132 1402
rect 132 1397 183 1402
rect 132 1385 174 1397
rect 124 1380 174 1385
rect 174 1380 183 1397
rect 124 1377 183 1380
rect 853 1356 857 1373
rect 857 1356 874 1373
rect 874 1356 879 1373
rect 853 1303 879 1356
rect 853 1287 857 1303
rect 857 1287 874 1303
rect 874 1287 879 1303
<< metal2 >>
rect 169 1456 193 1503
rect 529 1476 554 1502
rect 117 1449 193 1456
rect 117 1377 124 1449
rect 183 1421 193 1449
rect 183 1398 571 1421
rect 183 1377 193 1398
rect 117 1374 193 1377
rect 117 1373 162 1374
rect 548 1362 571 1398
rect 635 1378 660 1415
rect 850 1373 883 1377
rect 850 1362 853 1373
rect 278 1329 497 1351
rect 548 1342 853 1362
rect 574 1341 853 1342
rect 638 1293 659 1322
rect 850 1287 853 1341
rect 879 1287 883 1373
rect 850 1284 883 1287
rect 963 1232 978 1254
rect 533 1209 558 1232
rect 91 1168 237 1192
rect 377 1168 405 1192
rect 91 1167 155 1168
rect 963 1150 978 1172
rect 482 1085 659 1105
rect 325 1050 341 1068
rect 323 1049 341 1050
rect 301 1036 341 1049
rect 301 987 337 1036
rect 453 1004 659 1025
rect 95 901 260 924
rect 373 900 399 925
<< rmetal2 >>
rect 162 1373 193 1374
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1628616688
transform 1 0 823 0 1 939
box 0 0 358 746
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_2
timestamp 1628616688
transform 1 0 0 0 1 1338
box 0 0 549 1063
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1628616688
transform 1 0 331 0 -1 1063
box 0 0 549 1063
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_0
timestamp 1628616688
transform 1 0 175 0 1 1338
box 0 0 549 1063
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628616688
transform 1 0 179 0 1 1467
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628616688
transform 1 0 263 0 1 1339
box 0 0 34 33
<< labels >>
rlabel metal1 782 898 816 904 0 VGND
port 3 nsew ground default
rlabel metal1 849 898 876 904 0 VPWR
port 4 nsew power default
rlabel metal1 782 1498 816 1503 0 VGND
port 3 nsew ground default
rlabel metal1 849 1498 876 1503 0 VPWR
port 4 nsew power default
rlabel metal2 377 1168 400 1192 0 VIN11
port 7 nsew analog default
rlabel metal2 533 1209 558 1232 0 VIN21
port 6 nsew analog default
rlabel metal2 373 900 396 925 0 VIN12
port 8 nsew analog default
rlabel metal2 529 1476 554 1502 0 VIN22
port 5 nsew analog default
rlabel metal2 963 1150 978 1172 0 VOUT_AMP1
port 2 nsew analog default
rlabel metal2 963 1232 978 1254 0 VOUT_AMP2
port 1 nsew analog default
rlabel metal2 169 1495 193 1503 0 VPWR
port 4 nsew power default
rlabel metal2 133 1168 140 1192 0 VBIAS1
port 10 nsew analog default
rlabel metal2 133 901 140 924 0 VBIAS2
port 9 nsew analog default
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
