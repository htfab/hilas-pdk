magic
tech sky130A
timestamp 1627400275
<< error_s >>
rect 2146 7164 2175 7180
rect 2225 7164 2254 7180
rect 2304 7164 2333 7180
rect 2383 7164 2412 7180
rect 1008 7140 1015 7146
rect 1859 7140 1865 7146
rect 2691 7140 2697 7146
rect 2796 7140 2802 7146
rect 3211 7135 3217 7141
rect 3266 7135 3272 7141
rect 2146 7130 2147 7131
rect 2174 7130 2175 7131
rect 2225 7130 2226 7131
rect 2253 7130 2254 7131
rect 2304 7130 2305 7131
rect 2332 7130 2333 7131
rect 2383 7130 2384 7131
rect 2411 7130 2412 7131
rect 2096 7101 2113 7130
rect 2145 7129 2176 7130
rect 2224 7129 2255 7130
rect 2303 7129 2334 7130
rect 2382 7129 2413 7130
rect 2146 7122 2175 7129
rect 2225 7122 2254 7129
rect 2304 7122 2333 7129
rect 2383 7122 2412 7129
rect 2146 7108 2155 7122
rect 2402 7108 2412 7122
rect 2146 7102 2175 7108
rect 2225 7102 2254 7108
rect 2304 7102 2333 7108
rect 2383 7102 2412 7108
rect 2145 7101 2176 7102
rect 2224 7101 2255 7102
rect 2303 7101 2334 7102
rect 2382 7101 2413 7102
rect 2444 7101 2462 7130
rect 2146 7100 2147 7101
rect 2174 7100 2175 7101
rect 2225 7100 2226 7101
rect 2253 7100 2254 7101
rect 2304 7100 2305 7101
rect 2332 7100 2333 7101
rect 2383 7100 2384 7101
rect 2411 7100 2412 7101
rect 2685 7090 2691 7096
rect 2802 7090 2808 7096
rect 3205 7085 3211 7091
rect 3272 7085 3278 7091
rect 2146 7051 2175 7066
rect 2225 7051 2254 7066
rect 2304 7051 2333 7066
rect 2383 7051 2412 7066
rect 2146 6884 2175 6900
rect 2225 6884 2254 6900
rect 2304 6884 2333 6900
rect 2383 6884 2412 6900
rect 700 6881 705 6882
rect 2146 6850 2147 6851
rect 2174 6850 2175 6851
rect 2225 6850 2226 6851
rect 2253 6850 2254 6851
rect 2304 6850 2305 6851
rect 2332 6850 2333 6851
rect 2383 6850 2384 6851
rect 2411 6850 2412 6851
rect 2096 6821 2113 6850
rect 2145 6849 2176 6850
rect 2224 6849 2255 6850
rect 2303 6849 2334 6850
rect 2382 6849 2413 6850
rect 2146 6842 2175 6849
rect 2225 6842 2254 6849
rect 2304 6842 2333 6849
rect 2383 6842 2412 6849
rect 2146 6828 2155 6842
rect 2402 6828 2412 6842
rect 2146 6822 2175 6828
rect 2225 6822 2254 6828
rect 2304 6822 2333 6828
rect 2383 6822 2412 6828
rect 2145 6821 2176 6822
rect 2224 6821 2255 6822
rect 2303 6821 2334 6822
rect 2382 6821 2413 6822
rect 2444 6821 2462 6850
rect 2691 6841 2697 6847
rect 2796 6841 2802 6847
rect 2146 6820 2147 6821
rect 2174 6820 2175 6821
rect 2225 6820 2226 6821
rect 2253 6820 2254 6821
rect 2304 6820 2305 6821
rect 2332 6820 2333 6821
rect 2383 6820 2384 6821
rect 2411 6820 2412 6821
rect 3242 6802 3271 6820
rect 2685 6791 2691 6797
rect 2802 6791 2808 6797
rect 2146 6771 2175 6786
rect 2225 6771 2254 6786
rect 2304 6771 2333 6786
rect 2383 6771 2412 6786
rect 3242 6770 3243 6771
rect 3270 6770 3271 6771
rect 412 6714 413 6769
rect 2146 6729 2175 6745
rect 2225 6729 2254 6745
rect 2304 6729 2333 6745
rect 2383 6729 2412 6745
rect 2691 6740 2697 6746
rect 2796 6740 2802 6746
rect 3192 6741 3210 6770
rect 3241 6769 3272 6770
rect 3242 6760 3271 6769
rect 3242 6751 3252 6760
rect 3261 6751 3271 6760
rect 3242 6742 3271 6751
rect 3241 6741 3272 6742
rect 3303 6741 3321 6770
rect 3242 6740 3243 6741
rect 3270 6740 3271 6741
rect 2146 6695 2147 6696
rect 2174 6695 2175 6696
rect 2225 6695 2226 6696
rect 2253 6695 2254 6696
rect 2304 6695 2305 6696
rect 2332 6695 2333 6696
rect 2383 6695 2384 6696
rect 2411 6695 2412 6696
rect 1003 6674 1009 6680
rect 1865 6674 1871 6680
rect 2096 6666 2113 6695
rect 2145 6694 2176 6695
rect 2224 6694 2255 6695
rect 2303 6694 2334 6695
rect 2382 6694 2413 6695
rect 2146 6687 2175 6694
rect 2225 6687 2254 6694
rect 2304 6687 2333 6694
rect 2383 6687 2412 6694
rect 2146 6673 2155 6687
rect 2402 6673 2412 6687
rect 2146 6667 2175 6673
rect 2225 6667 2254 6673
rect 2304 6667 2333 6673
rect 2383 6667 2412 6673
rect 2145 6666 2176 6667
rect 2224 6666 2255 6667
rect 2303 6666 2334 6667
rect 2382 6666 2413 6667
rect 2444 6666 2462 6695
rect 2685 6690 2691 6696
rect 2802 6690 2808 6696
rect 3242 6691 3271 6709
rect 2146 6665 2147 6666
rect 2174 6665 2175 6666
rect 2225 6665 2226 6666
rect 2253 6665 2254 6666
rect 2304 6665 2305 6666
rect 2332 6665 2333 6666
rect 2383 6665 2384 6666
rect 2411 6665 2412 6666
rect 2146 6616 2175 6631
rect 2225 6616 2254 6631
rect 2304 6616 2333 6631
rect 2383 6616 2412 6631
rect 6818 5860 6831 5861
rect 6437 5639 6443 5645
rect 6490 5639 6496 5645
rect 6603 5639 6609 5645
rect 6656 5639 6662 5645
rect 6431 5589 6437 5595
rect 6496 5589 6502 5595
rect 6597 5589 6603 5595
rect 6662 5589 6668 5595
rect 6009 5580 6015 5586
rect 6114 5580 6120 5586
rect 7026 5580 7032 5586
rect 7131 5580 7137 5586
rect 6003 5530 6009 5536
rect 6120 5530 6126 5536
rect 7020 5530 7026 5536
rect 7137 5530 7143 5536
rect 3870 5400 4233 5401
rect 4290 5400 4413 5401
rect 4488 5394 4518 5513
rect 6009 5279 6015 5285
rect 6114 5279 6120 5285
rect 7026 5279 7032 5285
rect 7131 5279 7137 5285
rect 6003 5229 6009 5235
rect 6120 5229 6126 5235
rect 6437 5225 6443 5231
rect 6490 5225 6496 5231
rect 6603 5225 6609 5231
rect 6656 5225 6662 5231
rect 7020 5229 7026 5235
rect 7137 5229 7143 5235
rect 6431 5175 6437 5181
rect 6496 5175 6502 5181
rect 6597 5175 6603 5181
rect 6662 5175 6668 5181
rect 6271 5112 6275 5123
rect 6271 5098 6272 5109
rect 6380 5108 6381 5161
rect 6438 5036 6444 5042
rect 6491 5036 6497 5042
rect 6603 5036 6609 5042
rect 6656 5036 6662 5042
rect 6432 4986 6438 4992
rect 6497 4986 6503 4992
rect 6597 4986 6603 4992
rect 6662 4986 6668 4992
rect 5963 4977 5969 4983
rect 6068 4977 6074 4983
rect 7026 4977 7032 4983
rect 7131 4977 7137 4983
rect 5957 4927 5963 4933
rect 6074 4927 6080 4933
rect 7020 4927 7026 4933
rect 7137 4927 7143 4933
rect 6831 4792 6848 4793
rect 6831 4775 6848 4776
rect 6269 4758 6270 4771
rect 5963 4676 5969 4682
rect 6068 4676 6074 4682
rect 7026 4676 7032 4682
rect 7131 4676 7137 4682
rect 5957 4626 5963 4632
rect 6074 4626 6080 4632
rect 6438 4622 6444 4628
rect 6491 4622 6497 4628
rect 6603 4622 6609 4628
rect 6656 4622 6662 4628
rect 7020 4626 7026 4632
rect 7137 4626 7143 4632
rect 6432 4572 6438 4578
rect 6497 4572 6503 4578
rect 6597 4572 6603 4578
rect 6662 4572 6668 4578
rect 6011 4311 6017 4317
rect 6116 4311 6122 4317
rect 6982 4311 6988 4317
rect 7087 4311 7093 4317
rect 6437 4301 6443 4307
rect 6490 4301 6496 4307
rect 6608 4301 6614 4307
rect 6661 4301 6667 4307
rect 6005 4247 6011 4253
rect 6122 4247 6128 4253
rect 6431 4251 6437 4257
rect 6496 4251 6502 4257
rect 6602 4251 6608 4257
rect 6667 4251 6673 4257
rect 6976 4247 6982 4253
rect 7093 4247 7099 4253
rect 6011 4194 6017 4200
rect 6116 4194 6122 4200
rect 6437 4192 6443 4198
rect 6490 4192 6496 4198
rect 6608 4192 6614 4198
rect 6661 4192 6667 4198
rect 6982 4194 6988 4200
rect 7087 4194 7093 4200
rect 6431 4142 6437 4148
rect 6496 4142 6502 4148
rect 6602 4142 6608 4148
rect 6667 4142 6673 4148
rect 6005 4130 6011 4136
rect 6122 4130 6128 4136
rect 6976 4130 6982 4136
rect 7093 4130 7099 4136
rect 6011 4009 6017 4015
rect 6116 4009 6122 4015
rect 6982 4009 6988 4015
rect 7087 4009 7093 4015
rect 6437 4003 6443 4009
rect 6490 4003 6496 4009
rect 6608 4003 6614 4009
rect 6661 4003 6667 4009
rect 6431 3953 6437 3959
rect 6496 3953 6502 3959
rect 6602 3953 6608 3959
rect 6667 3953 6673 3959
rect 6005 3945 6011 3951
rect 6122 3945 6128 3951
rect 6976 3945 6982 3951
rect 7093 3945 7099 3951
rect 6011 3893 6017 3899
rect 6116 3893 6122 3899
rect 6982 3893 6988 3899
rect 7087 3893 7093 3899
rect 6437 3886 6443 3892
rect 6490 3886 6496 3892
rect 6608 3886 6614 3892
rect 6661 3886 6667 3892
rect 6431 3836 6437 3842
rect 6496 3836 6502 3842
rect 6602 3836 6608 3842
rect 6667 3836 6673 3842
rect 6005 3829 6011 3835
rect 6122 3829 6128 3835
rect 6976 3829 6982 3835
rect 7093 3829 7099 3835
rect 6011 3333 6017 3339
rect 6116 3333 6122 3339
rect 6437 3323 6443 3329
rect 6490 3323 6496 3329
rect 6005 3269 6011 3275
rect 6122 3269 6128 3275
rect 6431 3273 6437 3279
rect 6496 3273 6502 3279
rect 6011 3216 6017 3222
rect 6116 3216 6122 3222
rect 6437 3214 6443 3220
rect 6490 3214 6496 3220
rect 6431 3164 6437 3170
rect 6496 3164 6502 3170
rect 6005 3152 6011 3158
rect 6122 3152 6128 3158
rect 6011 3031 6017 3037
rect 6116 3031 6122 3037
rect 6274 3026 6291 3030
rect 6437 3025 6443 3031
rect 6490 3025 6496 3031
rect 6431 2975 6437 2981
rect 6496 2975 6502 2981
rect 6005 2967 6011 2973
rect 6122 2967 6128 2973
rect 6011 2915 6017 2921
rect 6116 2915 6122 2921
rect 6437 2908 6443 2914
rect 6490 2908 6496 2914
rect 6431 2858 6437 2864
rect 6496 2858 6502 2864
rect 6005 2851 6011 2857
rect 6122 2851 6128 2857
rect 11573 2112 11574 2125
rect 11573 2111 11587 2112
rect 1275 1953 1282 1991
rect 1289 1959 1296 2005
rect 1841 1569 1853 1572
rect 1829 1548 1834 1560
rect 6164 1520 6165 1538
rect 6178 1520 6179 1524
rect 1822 1208 1834 1216
rect 2053 1208 2055 1216
rect 10583 1063 10584 1065
rect 3516 313 3683 326
rect 4109 316 4111 329
rect 3513 299 3683 312
rect 4109 302 4112 315
rect 4519 314 4520 327
rect 4519 300 4521 313
<< nwell >>
rect 3969 5395 3993 5400
rect 3945 5394 4092 5395
rect 3915 5386 4092 5394
rect 4518 5386 4739 5395
rect 5333 5370 5401 5371
rect 5332 4765 5402 5370
rect 7722 5055 7778 5109
rect 5332 2790 5507 3390
rect 5522 2077 5724 2646
rect 10786 465 10921 2012
rect 10785 418 10921 465
<< psubdiff >>
rect 668 6247 2470 6260
rect 668 6176 2040 6247
rect 2129 6176 2470 6247
rect 668 6169 2470 6176
rect 2379 2439 2470 6169
rect 6774 5942 8385 5947
rect 6774 5860 6787 5942
rect 6813 5941 8385 5942
rect 6813 5863 8120 5941
rect 8209 5863 8385 5941
rect 6813 5860 8385 5863
rect 6774 5856 8385 5860
rect 8294 4037 8385 5856
rect 2379 2405 2390 2439
rect 2407 2422 2424 2439
rect 2441 2422 2470 2439
rect 2458 2405 2470 2422
rect 2379 2387 2470 2405
rect 2379 2326 2393 2387
rect 2446 2326 2470 2387
rect 1834 1560 2052 1569
rect 1834 1208 1841 1560
rect 1858 1208 1877 1560
rect 1894 1208 1912 1560
rect 1929 1208 1947 1560
rect 1964 1208 1983 1560
rect 2000 1208 2018 1560
rect 2035 1208 2053 1560
rect 2379 1276 2470 2326
rect 8045 3946 8385 4037
rect 8045 1276 8136 3946
rect 1822 1201 2055 1208
rect 1834 1195 2052 1201
rect 2379 1185 9537 1276
rect 2379 788 2470 1185
<< nsubdiff >>
rect 10827 1981 10884 1989
rect 10827 486 10840 1981
rect 10857 486 10884 1981
rect 10827 480 10884 486
<< psubdiffcont >>
rect 2040 6176 2129 6247
rect 6787 5860 6813 5942
rect 8120 5863 8209 5941
rect 2390 2422 2407 2439
rect 2424 2422 2441 2439
rect 2390 2405 2458 2422
rect 2393 2326 2446 2387
rect 1841 1208 1858 1560
rect 1877 1208 1894 1560
rect 1912 1208 1929 1560
rect 1947 1208 1964 1560
rect 1983 1208 2000 1560
rect 2018 1208 2035 1560
<< nsubdiffcont >>
rect 10840 486 10857 1981
<< locali >>
rect 1982 6252 2134 6253
rect 1982 6250 2137 6252
rect 1982 6176 1989 6250
rect 2032 6247 2137 6250
rect 2032 6176 2040 6247
rect 2129 6176 2137 6247
rect 1982 6173 2137 6176
rect 6779 5942 6846 5944
rect 6779 5860 6787 5942
rect 6813 5860 6818 5942
rect 6844 5860 6846 5942
rect 6779 5857 6846 5860
rect 8007 5942 8217 5944
rect 8007 5863 8013 5942
rect 8045 5941 8217 5942
rect 8045 5863 8120 5941
rect 8209 5863 8217 5941
rect 8007 5859 8217 5863
rect 2382 2405 2390 2439
rect 2382 2397 2458 2405
rect 2384 2387 2458 2397
rect 2384 2326 2393 2387
rect 2446 2326 2458 2387
rect 2384 2318 2458 2326
rect 10840 1982 10877 1989
rect 10840 1981 10860 1982
rect 1817 1560 2056 1565
rect 1817 1528 1823 1560
rect 1822 1208 1823 1528
rect 1840 1208 1841 1560
rect 1858 1208 1860 1560
rect 1894 1208 1895 1560
rect 1946 1208 1947 1560
rect 1981 1208 1983 1560
rect 2017 1208 2018 1560
rect 2035 1208 2036 1560
rect 2053 1208 2056 1560
rect 1822 1202 2056 1208
rect 1822 1201 2055 1202
rect 10857 487 10860 1981
rect 10877 487 10878 502
rect 10857 486 10878 487
rect 10840 477 10878 486
<< viali >>
rect 1989 6176 2032 6250
rect 6818 5860 6844 5942
rect 8013 5863 8045 5942
rect 2407 2422 2424 2439
rect 2407 2405 2424 2422
rect 2441 2422 2458 2439
rect 2441 2405 2458 2422
rect 1823 1208 1840 1560
rect 1860 1208 1877 1560
rect 1895 1208 1912 1560
rect 1929 1208 1946 1560
rect 1964 1208 1981 1560
rect 2000 1208 2017 1560
rect 2036 1208 2053 1560
rect 10860 487 10877 1982
<< metal1 >>
rect 8015 7642 8049 7656
rect 8803 7642 8875 7816
rect 8015 7570 8875 7642
rect 2808 7325 2942 7370
rect 198 7285 248 7289
rect 198 7246 203 7285
rect 242 7246 248 7285
rect 2808 7283 4160 7325
rect 4339 7316 4658 7428
rect 2808 7269 2942 7283
rect 198 7241 248 7246
rect 208 6945 247 7241
rect 2267 7209 2544 7233
rect 2267 7168 2291 7209
rect 208 6940 255 6945
rect 208 6901 211 6940
rect 250 6901 255 6940
rect 208 6896 255 6901
rect 208 6895 253 6896
rect 208 1084 247 6895
rect 349 6810 375 6813
rect 349 6781 375 6784
rect 350 6559 374 6781
rect 341 6556 383 6559
rect 341 6511 383 6514
rect 930 6435 959 6627
rect 928 6432 969 6435
rect 928 6374 936 6432
rect 965 6374 969 6432
rect 928 6368 969 6374
rect 2266 6299 2290 6622
rect 2261 6294 2295 6299
rect 2261 6268 2265 6294
rect 2291 6268 2295 6294
rect 2261 6265 2295 6268
rect 1986 6255 2035 6256
rect 1985 6250 2036 6255
rect 1985 6176 1989 6250
rect 2032 6176 2036 6250
rect 1593 5386 1616 5734
rect 1660 5672 1682 5734
rect 1929 5706 1951 6161
rect 1985 6140 2036 6176
rect 2520 6162 2544 7209
rect 2851 7176 3154 7203
rect 3322 7177 3348 7283
rect 2848 6259 2879 6629
rect 2840 6256 2879 6259
rect 2840 6225 2844 6256
rect 2875 6225 2879 6256
rect 2840 6222 2879 6225
rect 3127 6208 3154 7176
rect 4118 6958 4160 7283
rect 4499 7034 4541 7316
rect 4499 7031 4546 7034
rect 4499 6989 4502 7031
rect 4544 6989 4546 7031
rect 4499 6986 4546 6989
rect 4114 6955 4162 6958
rect 4114 6913 4117 6955
rect 4159 6913 4162 6955
rect 4114 6910 4162 6913
rect 4669 6796 4713 6799
rect 4669 6749 4713 6752
rect 5241 6796 5285 6799
rect 5241 6749 5285 6752
rect 5420 6793 5493 7432
rect 5935 7417 6033 7432
rect 5420 6749 5423 6793
rect 5467 6749 5493 6793
rect 4227 6694 4271 6697
rect 4227 6647 4271 6650
rect 3244 6308 3269 6623
rect 3948 6374 3980 6378
rect 3948 6373 3951 6374
rect 3939 6348 3951 6373
rect 3977 6348 3980 6374
rect 3939 6344 3980 6348
rect 3240 6305 3273 6308
rect 3240 6279 3244 6305
rect 3270 6279 3273 6305
rect 3240 6272 3273 6279
rect 3123 6206 3157 6208
rect 3123 6180 3127 6206
rect 3154 6180 3157 6206
rect 3123 6177 3157 6180
rect 1980 6137 2036 6140
rect 1980 6130 1994 6137
rect 1969 6102 1994 6130
rect 2029 6102 2036 6137
rect 2515 6159 2549 6162
rect 2515 6133 2519 6159
rect 2545 6133 2549 6159
rect 2515 6130 2549 6133
rect 1969 6090 2036 6102
rect 1969 6087 2035 6090
rect 1969 5706 1991 6087
rect 3939 5994 3963 6344
rect 4233 5987 4264 6647
rect 4676 5989 4705 6749
rect 4795 6650 4798 6694
rect 4842 6650 4845 6694
rect 2091 5917 2126 5921
rect 2091 5878 2096 5917
rect 2122 5878 2126 5917
rect 2091 5875 2126 5878
rect 3734 5905 3771 5908
rect 3734 5879 3736 5905
rect 3769 5879 3771 5905
rect 3734 5877 3771 5879
rect 2031 5839 2056 5851
rect 2028 5836 2060 5839
rect 2028 5796 2032 5836
rect 2058 5796 2060 5836
rect 2028 5793 2060 5796
rect 2031 5714 2056 5793
rect 2031 5711 2060 5714
rect 2031 5685 2034 5711
rect 2031 5682 2060 5685
rect 1657 5669 1683 5672
rect 1657 5640 1683 5643
rect 1660 5580 1682 5640
rect 1654 5577 1682 5580
rect 1680 5551 1682 5577
rect 1654 5548 1682 5551
rect 1660 5488 1682 5548
rect 1655 5485 1682 5488
rect 1681 5459 1682 5485
rect 1655 5456 1682 5459
rect 1590 5383 1616 5386
rect 1590 5354 1616 5357
rect 1593 5290 1616 5354
rect 1586 5287 1616 5290
rect 1612 5261 1616 5287
rect 1586 5258 1616 5261
rect 1593 5194 1616 5258
rect 1590 5191 1616 5194
rect 1590 5162 1616 5165
rect 1593 3687 1616 5162
rect 1660 3687 1682 5456
rect 2031 5622 2056 5682
rect 2031 5619 2060 5622
rect 2031 5593 2034 5619
rect 2031 5590 2060 5593
rect 2031 5530 2056 5590
rect 2031 5527 2057 5530
rect 2031 5498 2057 5501
rect 1582 3684 1616 3687
rect 1582 3637 1586 3684
rect 1612 3637 1616 3684
rect 1582 3634 1616 3637
rect 1648 3684 1682 3687
rect 1648 3637 1650 3684
rect 1676 3637 1682 3684
rect 1648 3634 1682 3637
rect 1451 3560 1474 3567
rect 1447 3534 1450 3560
rect 1476 3534 1479 3560
rect 1402 3523 1425 3527
rect 1398 3520 1425 3523
rect 1424 3494 1425 3520
rect 1398 3491 1425 3494
rect 467 3435 539 3437
rect 467 3369 470 3435
rect 536 3369 539 3435
rect 467 3367 539 3369
rect 468 2852 534 3367
rect 1402 3139 1425 3491
rect 1451 3287 1474 3534
rect 1593 3525 1616 3634
rect 1660 3561 1682 3634
rect 1836 3563 1863 3567
rect 1658 3558 1684 3561
rect 1658 3529 1684 3532
rect 1834 3560 1863 3563
rect 1861 3533 1863 3560
rect 1834 3530 1863 3533
rect 1592 3522 1618 3525
rect 1592 3493 1618 3496
rect 1781 3376 1810 3379
rect 1451 3250 1524 3287
rect 1402 3132 1428 3139
rect 1400 3131 1428 3132
rect 1397 3129 1429 3131
rect 1397 3103 1400 3129
rect 1426 3103 1429 3129
rect 1397 3100 1429 3103
rect 987 2954 1030 2957
rect 987 2917 991 2954
rect 1028 2917 1030 2954
rect 987 2914 1030 2917
rect 468 2849 542 2852
rect 468 2783 474 2849
rect 540 2783 542 2849
rect 468 2780 542 2783
rect 992 2333 1029 2914
rect 1451 2500 1474 3250
rect 1836 3233 1863 3530
rect 1824 3208 1863 3233
rect 1884 3523 1908 3527
rect 1884 3520 1910 3523
rect 1884 3491 1910 3494
rect 1884 3177 1908 3491
rect 1824 3154 1908 3177
rect 1451 2477 1696 2500
rect 1664 2444 1696 2477
rect 988 2330 1031 2333
rect 988 2293 990 2330
rect 1027 2293 1031 2330
rect 988 2290 1031 2293
rect 1740 2287 1773 2290
rect 1726 2279 1744 2287
rect 1702 2255 1744 2279
rect 1740 2251 1744 2255
rect 1770 2251 1773 2287
rect 1740 2248 1773 2251
rect 1289 1756 1318 1759
rect 1289 1724 1318 1727
rect 1290 1667 1316 1724
rect 1884 1688 1908 3154
rect 1929 3087 1951 5162
rect 1969 3348 1991 5162
rect 2031 3463 2056 5498
rect 2093 5421 2119 5875
rect 3670 5740 3709 5742
rect 3670 5707 3673 5740
rect 3706 5707 3709 5740
rect 3670 5705 3709 5707
rect 3612 5592 3651 5595
rect 3612 5559 3616 5592
rect 3649 5559 3651 5592
rect 3612 5556 3651 5559
rect 3548 5432 3587 5435
rect 2093 5418 2121 5421
rect 2093 5392 2095 5418
rect 3548 5399 3552 5432
rect 3585 5399 3587 5432
rect 3548 5397 3587 5399
rect 2093 5389 2121 5392
rect 3551 5396 3585 5397
rect 2093 5325 2119 5389
rect 3487 5377 3521 5378
rect 3486 5375 3522 5377
rect 3486 5342 3488 5375
rect 3521 5342 3522 5375
rect 3486 5338 3522 5342
rect 2093 5322 2122 5325
rect 2093 5296 2096 5322
rect 2093 5293 2122 5296
rect 2093 5229 2119 5293
rect 2093 5226 2121 5229
rect 2093 5200 2095 5226
rect 2093 5197 2121 5200
rect 3425 5218 3461 5221
rect 2031 3461 2057 3463
rect 2030 3460 2058 3461
rect 2030 3434 2031 3460
rect 2057 3434 2058 3460
rect 2030 3433 2058 3434
rect 2031 3431 2057 3433
rect 1965 3345 1997 3348
rect 1965 3319 1969 3345
rect 1995 3319 1997 3345
rect 1965 3316 1997 3319
rect 1925 3084 1953 3087
rect 1925 3058 1927 3084
rect 1925 3055 1953 3058
rect 1929 1758 1951 3055
rect 1969 2534 1991 3316
rect 1969 2531 1998 2534
rect 1969 2489 1971 2531
rect 1997 2489 1998 2531
rect 1969 2486 1998 2489
rect 1969 2290 1991 2486
rect 1967 2287 1993 2290
rect 1967 2248 1993 2251
rect 1969 1786 1991 2248
rect 2031 1924 2056 3431
rect 2093 3030 2119 5197
rect 3425 5185 3427 5218
rect 3460 5185 3461 5218
rect 3425 5182 3461 5185
rect 3360 5065 3401 5068
rect 3360 5032 3364 5065
rect 3397 5032 3401 5065
rect 3360 5028 3401 5032
rect 3307 4908 3343 4911
rect 3307 4875 3308 4908
rect 3341 4875 3343 4908
rect 3307 4872 3343 4875
rect 3249 4366 3282 4368
rect 3243 4361 3282 4366
rect 3243 4328 3246 4361
rect 3279 4328 3282 4361
rect 3243 4324 3282 4328
rect 3186 4205 3219 4207
rect 3181 4202 3220 4205
rect 3181 4169 3183 4202
rect 3216 4169 3220 4202
rect 3181 4166 3220 4169
rect 3124 4050 3157 4051
rect 3121 4047 3157 4050
rect 3154 4014 3157 4047
rect 3121 4011 3157 4014
rect 3059 3899 3098 3903
rect 3059 3866 3061 3899
rect 3094 3866 3098 3899
rect 3059 3863 3098 3866
rect 2992 3382 3035 3386
rect 2992 3349 2997 3382
rect 3030 3349 3035 3382
rect 2992 3346 3035 3349
rect 2926 3225 2967 3229
rect 2926 3192 2930 3225
rect 2963 3192 2967 3225
rect 2926 3189 2967 3192
rect 2865 3061 2904 3065
rect 2092 3027 2123 3030
rect 2092 3001 2095 3027
rect 2121 3001 2123 3027
rect 2865 3028 2868 3061
rect 2901 3028 2904 3061
rect 2865 3025 2904 3028
rect 2092 2998 2123 3001
rect 2027 1921 2057 1924
rect 2027 1888 2029 1921
rect 2055 1888 2057 1921
rect 2027 1884 2057 1888
rect 1969 1772 1993 1786
rect 1925 1755 1956 1758
rect 1925 1726 1926 1755
rect 1955 1726 1956 1755
rect 1925 1723 1956 1726
rect 1970 1709 1993 1772
rect 1805 1685 1908 1688
rect 1805 1625 1810 1685
rect 1870 1632 1908 1685
rect 1969 1706 1993 1709
rect 1870 1625 1884 1632
rect 1805 1621 1884 1625
rect 1969 1567 1991 1706
rect 1816 1560 2058 1567
rect 1816 1208 1823 1560
rect 1840 1208 1860 1560
rect 1877 1208 1895 1560
rect 1912 1208 1929 1560
rect 1946 1208 1964 1560
rect 1981 1208 2000 1560
rect 2017 1208 2036 1560
rect 2053 1208 2058 1560
rect 1816 1199 2058 1208
rect 2093 1170 2119 2998
rect 2796 2917 2837 2920
rect 2796 2884 2800 2917
rect 2833 2884 2837 2917
rect 2796 2881 2837 2884
rect 2375 2519 2468 2531
rect 2375 2448 2396 2519
rect 2454 2448 2468 2519
rect 2375 2439 2468 2448
rect 2375 2405 2407 2439
rect 2424 2405 2441 2439
rect 2458 2405 2468 2439
rect 2375 2366 2468 2405
rect 2384 2318 2458 2366
rect 2084 1166 2119 1170
rect 2084 1132 2088 1166
rect 2114 1132 2119 1166
rect 2084 1129 2119 1132
rect 191 1077 247 1084
rect 191 1038 197 1077
rect 236 1038 247 1077
rect 191 1032 247 1038
rect 2802 547 2835 2881
rect 2797 546 2840 547
rect 2794 544 2843 546
rect 2794 501 2797 544
rect 2840 501 2843 544
rect 2794 500 2843 501
rect 2797 498 2840 500
rect 2867 468 2900 3025
rect 2858 465 2907 468
rect 2858 422 2862 465
rect 2905 422 2907 465
rect 2858 419 2907 422
rect 2932 397 2965 3189
rect 2929 394 2969 397
rect 2929 351 2969 354
rect 2908 311 2966 313
rect 2908 260 2912 311
rect 2963 302 2966 311
rect 2999 302 3032 3346
rect 3063 760 3096 3863
rect 3063 314 3095 760
rect 3124 375 3157 4011
rect 3186 436 3219 4166
rect 3249 503 3282 4324
rect 3309 569 3342 4872
rect 3367 626 3400 5028
rect 3428 693 3461 5182
rect 3487 754 3520 5338
rect 3551 821 3584 5396
rect 3613 886 3646 5556
rect 3673 949 3706 5705
rect 3736 1010 3769 5877
rect 4263 5394 4264 5395
rect 3939 5386 3963 5394
rect 4233 5386 4264 5394
rect 4676 5386 4705 5394
rect 4822 5350 4841 6650
rect 5250 5346 5275 6749
rect 5420 6745 5493 6749
rect 5436 5706 5453 6745
rect 5936 6692 6033 7417
rect 7198 7315 7517 7427
rect 6475 6955 6622 6961
rect 6475 6913 6479 6955
rect 6614 6913 6622 6955
rect 6475 6908 6622 6913
rect 6238 6694 6282 6697
rect 5934 6690 6035 6692
rect 5934 6649 5937 6690
rect 6032 6649 6035 6690
rect 5934 6645 6035 6649
rect 6238 6647 6282 6650
rect 5658 6298 5692 6301
rect 5658 6272 5663 6298
rect 5689 6272 5692 6298
rect 5663 6269 5689 6272
rect 5475 5945 5501 5948
rect 5475 5916 5501 5919
rect 5478 5693 5497 5916
rect 5665 5691 5686 6269
rect 6022 6209 6048 6210
rect 6020 6207 6050 6209
rect 6020 6181 6022 6207
rect 6048 6181 6050 6207
rect 6020 6179 6050 6181
rect 6022 6178 6048 6179
rect 5705 6105 5739 6108
rect 5705 6079 5709 6105
rect 5735 6079 5739 6105
rect 5705 6076 5739 6079
rect 5712 5693 5731 6076
rect 5749 5896 5778 5899
rect 5749 5870 5751 5896
rect 5777 5870 5778 5896
rect 5749 5867 5778 5870
rect 5753 5691 5774 5867
rect 5853 5848 5887 5851
rect 5853 5822 5857 5848
rect 5883 5822 5887 5848
rect 5853 5819 5887 5822
rect 5861 5694 5879 5819
rect 6025 5155 6045 6178
rect 6248 5689 6271 6647
rect 6338 6299 6366 6302
rect 6338 6273 6339 6299
rect 6365 6273 6366 6299
rect 6338 6270 6366 6273
rect 6294 6208 6322 6211
rect 6294 6182 6295 6208
rect 6321 6182 6322 6208
rect 6294 6179 6322 6182
rect 6023 5142 6045 5155
rect 6018 5139 6051 5142
rect 6018 5112 6021 5139
rect 6048 5112 6051 5139
rect 6018 5109 6051 5112
rect 6297 5025 6319 6179
rect 6296 5018 6319 5025
rect 6295 4958 6315 5018
rect 6340 4973 6363 6270
rect 6477 5670 6519 6908
rect 6580 5670 6622 6908
rect 6818 6690 6862 6693
rect 6818 6643 6862 6646
rect 6828 5945 6851 6643
rect 7270 6118 7398 7315
rect 7646 6796 7674 6808
rect 7646 6793 7679 6796
rect 7646 6749 7651 6793
rect 7646 6746 7679 6749
rect 7270 6110 7400 6118
rect 7269 6109 7400 6110
rect 7269 6083 7273 6109
rect 7395 6083 7400 6109
rect 7269 6080 7400 6083
rect 6947 6044 6977 6047
rect 6947 6018 6949 6044
rect 6975 6018 6977 6044
rect 6947 6015 6977 6018
rect 6815 5944 6851 5945
rect 6812 5942 6851 5944
rect 6812 5860 6818 5942
rect 6844 5860 6851 5942
rect 6812 5859 6851 5860
rect 6815 5858 6851 5859
rect 6828 5689 6851 5858
rect 6950 5689 6973 6015
rect 7578 5990 7621 5994
rect 7578 5964 7582 5990
rect 7608 5964 7621 5990
rect 7578 5960 7621 5964
rect 7602 5693 7621 5960
rect 7646 5684 7674 6746
rect 7816 6299 7842 6302
rect 7816 6270 7842 6273
rect 7727 6212 7753 6215
rect 7727 6183 7753 6186
rect 7730 5811 7749 6183
rect 7818 5811 7840 6270
rect 8015 5948 8049 7570
rect 10055 7318 10374 7430
rect 8465 7224 8502 7225
rect 8460 7220 8510 7224
rect 8460 7183 8468 7220
rect 8505 7183 8510 7220
rect 8460 7179 8510 7183
rect 8080 6371 8112 6375
rect 8080 6344 8083 6371
rect 8109 6344 8112 6371
rect 8080 6338 8112 6344
rect 8010 5942 8049 5948
rect 8010 5940 8013 5942
rect 8009 5863 8013 5940
rect 8045 5863 8049 5942
rect 8010 5856 8049 5863
rect 7713 5791 7781 5811
rect 7713 5765 7727 5791
rect 7753 5765 7781 5791
rect 7713 5742 7781 5765
rect 7817 5792 7885 5811
rect 7817 5766 7829 5792
rect 7855 5766 7885 5792
rect 7817 5742 7885 5766
rect 8015 5678 8049 5856
rect 8082 5800 8109 6338
rect 8082 5797 8150 5800
rect 8082 5754 8104 5797
rect 8147 5754 8150 5797
rect 8082 5750 8150 5754
rect 8082 5685 8109 5750
rect 6296 4955 6319 4958
rect 3939 4349 3963 4786
rect 4233 4342 4264 4793
rect 4676 4344 4705 4791
rect 4822 4345 4841 4785
rect 4953 4364 4976 4789
rect 5250 4364 5275 4791
rect 6297 4635 6319 4955
rect 6297 4626 6332 4635
rect 6297 4604 6348 4626
rect 5426 4421 5454 4532
rect 5479 4463 5498 4523
rect 5679 4479 5718 4481
rect 5678 4476 5718 4479
rect 5678 4470 5685 4476
rect 5479 4444 5642 4463
rect 5426 4393 5598 4421
rect 5570 4370 5598 4393
rect 5623 4366 5642 4444
rect 5663 4448 5685 4470
rect 5713 4448 5718 4476
rect 5663 4445 5718 4448
rect 5663 4443 5717 4445
rect 5663 4358 5679 4443
rect 6075 4436 6113 4438
rect 6127 4436 6150 4527
rect 6075 4413 6150 4436
rect 6249 4427 6272 4527
rect 6580 4428 6622 4546
rect 6828 4429 6851 4527
rect 6950 4438 6973 4527
rect 6075 4336 6113 4413
rect 6249 4397 6274 4427
rect 6250 4350 6274 4397
rect 6580 4389 6626 4428
rect 6828 4394 6854 4429
rect 6948 4400 7029 4438
rect 7602 4425 7621 4523
rect 6586 4334 6626 4389
rect 6830 4350 6854 4394
rect 6991 4336 7029 4400
rect 7419 4417 7447 4420
rect 7419 4391 7420 4417
rect 7446 4391 7447 4417
rect 7419 4388 7447 4391
rect 7462 4406 7621 4425
rect 7425 4358 7441 4388
rect 7462 4371 7481 4406
rect 7646 4387 7674 4532
rect 8465 4488 8502 7179
rect 8544 6874 8590 6877
rect 8544 6837 8550 6874
rect 8587 6837 8590 6874
rect 8544 6834 8590 6837
rect 8462 4483 8507 4488
rect 8462 4446 8469 4483
rect 8506 4446 8507 4483
rect 8462 4442 8507 4446
rect 8465 4438 8502 4442
rect 8546 4429 8583 6834
rect 8621 6403 8666 6406
rect 8621 6366 8627 6403
rect 8664 6366 8666 6403
rect 8621 6363 8666 6366
rect 7507 4359 7674 4387
rect 8543 4424 8587 4429
rect 8543 4387 8546 4424
rect 8583 4387 8587 4424
rect 8543 4383 8587 4387
rect 8546 4378 8583 4383
rect 8623 4194 8660 6363
rect 9278 6311 9336 6314
rect 9278 6261 9282 6311
rect 9332 6261 9336 6311
rect 9278 6258 9336 6261
rect 9160 6251 9216 6255
rect 9052 6204 9108 6208
rect 8957 6155 9013 6166
rect 8957 6105 8960 6155
rect 9010 6105 9013 6155
rect 8957 6101 9013 6105
rect 9052 6154 9055 6204
rect 9105 6154 9108 6204
rect 9160 6201 9163 6251
rect 9213 6201 9216 6251
rect 9160 6196 9216 6201
rect 9052 6150 9108 6154
rect 8710 5896 8753 5899
rect 8710 5859 8715 5896
rect 8752 5859 8753 5896
rect 8710 5855 8753 5859
rect 8620 4193 8660 4194
rect 8619 4191 8661 4193
rect 8619 4154 8620 4191
rect 8657 4154 8661 4191
rect 8619 4151 8661 4154
rect 8623 4150 8660 4151
rect 3939 3396 3963 3773
rect 4233 3396 4264 3780
rect 4676 3396 4705 3778
rect 4822 3369 4841 3778
rect 4953 3674 4976 3782
rect 4944 3670 4977 3674
rect 4944 3629 4948 3670
rect 4974 3629 4977 3670
rect 4944 3626 4977 3629
rect 4953 3365 4976 3626
rect 5250 3386 5275 3784
rect 5582 3380 5598 3785
rect 5857 3421 5881 3793
rect 5855 3396 5894 3421
rect 5869 3371 5894 3396
rect 6075 3358 6113 3807
rect 6250 3419 6274 3793
rect 6250 3392 6297 3419
rect 6270 3369 6297 3392
rect 6478 3356 6518 3809
rect 6830 3542 6854 3793
rect 8711 3676 8748 5855
rect 8707 3670 8756 3676
rect 8707 3629 8713 3670
rect 8750 3629 8756 3670
rect 8707 3625 8756 3629
rect 8711 3622 8748 3625
rect 6830 3518 6888 3542
rect 6864 3384 6888 3518
rect 5385 3283 5417 3287
rect 5385 3257 5388 3283
rect 5414 3257 5417 3283
rect 7376 3281 7402 3284
rect 5385 3253 5417 3257
rect 7375 3255 7376 3278
rect 3939 1533 3963 2796
rect 4233 2688 4264 2803
rect 4676 2739 4705 2801
rect 4726 2770 4760 2773
rect 4726 2744 4730 2770
rect 4756 2744 4760 2770
rect 4726 2741 4760 2744
rect 4673 2736 4708 2739
rect 4673 2707 4676 2736
rect 4705 2707 4708 2736
rect 4673 2704 4708 2707
rect 4229 2687 4266 2688
rect 4229 2656 4232 2687
rect 4263 2656 4266 2687
rect 4676 2658 4705 2704
rect 4726 2680 4751 2741
rect 4822 2682 4841 2802
rect 5250 2735 5275 2808
rect 5393 2777 5414 3253
rect 7375 3252 7402 3255
rect 7324 3188 7350 3191
rect 7324 3159 7350 3162
rect 5519 3084 5558 3109
rect 5447 3005 5481 3008
rect 5447 2979 5451 3005
rect 5477 2979 5481 3005
rect 5447 2974 5481 2979
rect 5451 2972 5473 2974
rect 5390 2774 5418 2777
rect 5390 2748 5391 2774
rect 5417 2748 5418 2774
rect 5390 2745 5418 2748
rect 5451 2744 5471 2972
rect 5497 2776 5516 2826
rect 5493 2773 5521 2776
rect 5493 2747 5494 2773
rect 5520 2747 5521 2773
rect 5447 2741 5475 2744
rect 5493 2743 5521 2747
rect 5247 2733 5281 2735
rect 5247 2707 5251 2733
rect 5277 2707 5281 2733
rect 5447 2715 5448 2741
rect 5474 2715 5475 2741
rect 5447 2712 5475 2715
rect 5247 2706 5281 2707
rect 4229 2655 4266 2656
rect 4233 2534 4264 2655
rect 4619 2630 4705 2658
rect 4611 2629 4705 2630
rect 4721 2669 4751 2680
rect 4816 2679 4848 2682
rect 4611 2627 4657 2629
rect 4611 2585 4613 2627
rect 4655 2585 4657 2627
rect 4611 2582 4657 2585
rect 4228 2531 4270 2534
rect 4721 2518 4740 2669
rect 4816 2653 4819 2679
rect 4845 2653 4848 2679
rect 4816 2650 4848 2653
rect 5084 2629 5159 2648
rect 5109 2545 5159 2629
rect 5540 2621 5558 3084
rect 7277 3004 7303 3007
rect 7277 2975 7303 2978
rect 7227 2911 7253 2914
rect 7227 2882 7253 2885
rect 5672 2737 5698 2740
rect 5670 2735 5700 2737
rect 5670 2709 5672 2735
rect 5698 2709 5700 2735
rect 5670 2707 5700 2709
rect 5672 2706 5698 2707
rect 5540 2617 5588 2621
rect 5540 2591 5552 2617
rect 5548 2584 5552 2591
rect 5585 2584 5588 2617
rect 5673 2614 5695 2706
rect 5869 2693 5894 2816
rect 6270 2695 6297 2818
rect 6552 2775 6595 2778
rect 6552 2740 6556 2775
rect 6591 2740 6595 2775
rect 6552 2738 6595 2740
rect 5868 2667 5871 2693
rect 5897 2667 5900 2693
rect 6270 2691 6305 2695
rect 6270 2664 6275 2691
rect 6302 2664 6305 2691
rect 5548 2580 5588 2584
rect 5667 2611 5701 2614
rect 5667 2574 5701 2577
rect 5673 2566 5695 2574
rect 6068 2547 6162 2640
rect 6556 2595 6591 2738
rect 6738 2682 6760 2814
rect 6864 2742 6887 2814
rect 6864 2719 7185 2742
rect 6864 2718 6887 2719
rect 6556 2563 6560 2595
rect 6586 2563 6591 2595
rect 6556 2559 6591 2563
rect 6709 2658 6760 2682
rect 4228 2486 4270 2489
rect 4677 2512 4740 2518
rect 5060 2513 5084 2545
rect 5184 2513 5208 2545
rect 6041 2515 6065 2547
rect 6165 2515 6189 2547
rect 6709 2533 6732 2658
rect 7162 2622 7185 2719
rect 7157 2619 7188 2622
rect 7157 2585 7159 2619
rect 7185 2585 7188 2619
rect 7157 2582 7188 2585
rect 6698 2530 6744 2533
rect 4677 2480 4681 2512
rect 4713 2486 4740 2512
rect 6698 2492 6702 2530
rect 6740 2492 6744 2530
rect 6698 2489 6744 2492
rect 4713 2480 4721 2486
rect 4677 2476 4721 2480
rect 5060 2379 5084 2411
rect 5184 2378 5208 2410
rect 6041 2381 6065 2413
rect 6165 2380 6189 2412
rect 7162 2265 7185 2582
rect 7149 2243 7185 2265
rect 7129 2220 7185 2243
rect 7129 2219 7183 2220
rect 4698 1958 4730 2133
rect 5060 2102 5084 2134
rect 5184 2101 5208 2133
rect 5084 2036 5110 2082
rect 5158 2038 5184 2082
rect 5083 2033 5111 2036
rect 5083 2002 5111 2005
rect 5157 2035 5185 2038
rect 5157 2004 5185 2007
rect 4686 1948 4740 1958
rect 4686 1902 4691 1948
rect 4737 1902 4740 1948
rect 4686 1898 4740 1902
rect 5084 1861 5110 2002
rect 5158 1861 5184 2004
rect 3899 1516 3964 1533
rect 5084 1518 5184 1861
rect 5535 1856 5569 2135
rect 5529 1853 5575 1856
rect 5529 1804 5575 1807
rect 5678 1767 5712 2134
rect 6041 2104 6065 2136
rect 6165 2104 6189 2136
rect 6065 2036 6091 2085
rect 6064 2033 6092 2036
rect 6064 2002 6092 2005
rect 6065 1884 6091 2002
rect 6139 1884 6165 2085
rect 5669 1764 5721 1767
rect 5669 1718 5672 1764
rect 5718 1718 5721 1764
rect 5669 1715 5721 1718
rect 6065 1520 6165 1884
rect 6520 1679 6547 2138
rect 7227 2098 7252 2882
rect 7277 2188 7302 2975
rect 7325 2279 7350 3159
rect 7375 2368 7400 3252
rect 8959 2518 9009 6101
rect 9052 3046 9102 6150
rect 9165 3569 9215 6196
rect 9278 4086 9328 6258
rect 10164 6098 10292 7318
rect 10163 6095 10292 6098
rect 10291 5967 10292 6095
rect 10163 5964 10292 5967
rect 10164 5915 10292 5964
rect 10600 5797 10620 5800
rect 10591 5794 10622 5797
rect 10591 5751 10595 5794
rect 10621 5751 10622 5794
rect 10591 5747 10622 5751
rect 10209 5665 10244 5668
rect 10209 5623 10212 5665
rect 10238 5623 10244 5665
rect 10209 5620 10244 5623
rect 9810 5343 9857 5349
rect 9810 5303 9812 5343
rect 9852 5303 9857 5343
rect 9810 5300 9857 5303
rect 9273 4083 9328 4086
rect 9323 4033 9328 4083
rect 9273 4030 9328 4033
rect 9164 3561 9216 3569
rect 9164 3514 9165 3561
rect 9215 3514 9216 3561
rect 9164 3513 9216 3514
rect 9051 3045 9103 3046
rect 9051 2995 9052 3045
rect 9102 2995 9103 3045
rect 9051 2994 9103 2995
rect 8943 2515 9009 2518
rect 8943 2465 8947 2515
rect 8997 2465 9009 2515
rect 8943 2461 9009 2465
rect 7370 2364 7407 2368
rect 7370 2314 7374 2364
rect 7400 2314 7407 2364
rect 7370 2310 7407 2314
rect 7317 2274 7354 2279
rect 7317 2224 7320 2274
rect 7346 2224 7354 2274
rect 7317 2221 7354 2224
rect 7268 2184 7305 2188
rect 7268 2134 7273 2184
rect 7299 2134 7305 2184
rect 7268 2130 7305 2134
rect 7221 2094 7256 2098
rect 6509 1673 6558 1679
rect 6509 1627 6511 1673
rect 6557 1627 6558 1673
rect 6509 1623 6558 1627
rect 6178 1520 6267 1524
rect 3899 1404 3904 1516
rect 3930 1404 3964 1516
rect 5036 1514 5229 1518
rect 3899 1401 3964 1404
rect 4982 1512 5229 1514
rect 4982 1510 5115 1512
rect 4982 1398 5041 1510
rect 5227 1400 5229 1512
rect 5153 1398 5229 1400
rect 4982 1395 5229 1398
rect 6017 1514 6267 1520
rect 6017 1395 6022 1514
rect 6208 1395 6267 1514
rect 3734 1008 3771 1010
rect 3734 975 3736 1008
rect 3769 975 3771 1008
rect 3734 972 3771 975
rect 3669 946 3708 949
rect 3669 913 3674 946
rect 3707 913 3708 946
rect 3669 910 3708 913
rect 3609 883 3647 886
rect 3609 850 3611 883
rect 3644 850 3647 883
rect 3609 847 3647 850
rect 3550 820 3585 821
rect 3550 787 3551 820
rect 3584 787 3585 820
rect 3550 784 3585 787
rect 3486 752 3522 754
rect 3486 719 3487 752
rect 3520 719 3522 752
rect 3486 716 3522 719
rect 3427 692 3461 693
rect 3425 690 3463 692
rect 3425 657 3427 690
rect 3460 657 3463 690
rect 3425 655 3463 657
rect 3427 654 3460 655
rect 3367 590 3400 593
rect 3309 533 3342 536
rect 3249 500 3284 503
rect 3249 470 3251 500
rect 3251 464 3284 467
rect 3186 400 3219 403
rect 3122 372 3157 375
rect 3155 342 3157 372
rect 3122 335 3155 338
rect 2963 269 3032 302
rect 3061 311 3105 314
rect 3061 274 3064 311
rect 3101 274 3105 311
rect 3061 272 3105 274
rect 2963 260 2966 269
rect 2908 258 2966 260
rect 4982 246 5076 1395
rect 6017 1392 6267 1395
rect 6178 392 6267 1392
rect 7094 1077 7127 2076
rect 7221 2044 7225 2094
rect 7251 2044 7256 2094
rect 7221 2041 7256 2044
rect 8959 1679 9009 2461
rect 9052 1770 9102 2994
rect 9165 1857 9215 3513
rect 9278 1959 9328 4030
rect 9567 2767 9625 2771
rect 9567 2717 9571 2767
rect 9621 2717 9625 2767
rect 9567 2715 9625 2717
rect 9570 2714 9621 2715
rect 9278 1956 9334 1959
rect 9278 1906 9284 1956
rect 9278 1903 9334 1906
rect 9278 1890 9328 1903
rect 9165 1808 9215 1811
rect 9052 1721 9102 1724
rect 8959 1630 9009 1633
rect 9570 1527 9620 2714
rect 9507 1516 9620 1527
rect 9507 1404 9513 1516
rect 9607 1404 9620 1516
rect 9507 1399 9620 1404
rect 7088 1074 7131 1077
rect 7088 1041 7092 1074
rect 7125 1041 7131 1074
rect 7088 1038 7131 1041
rect 9815 965 9855 5300
rect 9907 5239 9910 5275
rect 9946 5239 9949 5275
rect 9814 962 9861 965
rect 9814 922 9818 962
rect 9858 922 9861 962
rect 9814 919 9861 922
rect 9908 885 9947 5239
rect 9999 5041 10044 5043
rect 9999 5002 10002 5041
rect 10041 5002 10044 5041
rect 9999 5000 10044 5002
rect 9905 881 9951 885
rect 9905 842 9909 881
rect 9948 842 9951 881
rect 9905 838 9951 842
rect 10001 803 10040 5000
rect 10085 4974 10123 4975
rect 10083 4972 10125 4974
rect 10083 4946 10085 4972
rect 10123 4946 10125 4972
rect 10083 4944 10125 4946
rect 9999 799 10046 803
rect 9999 760 10002 799
rect 10041 760 10046 799
rect 9999 757 10046 760
rect 10085 723 10123 4944
rect 10219 2621 10242 5620
rect 10600 5422 10620 5747
rect 10951 5423 10970 7450
rect 11285 6571 11367 6574
rect 11285 6565 11290 6571
rect 11279 6500 11290 6565
rect 11361 6500 11367 6571
rect 11279 6496 11367 6500
rect 11279 4596 11350 6496
rect 11266 4592 11350 4596
rect 11266 4521 11271 4592
rect 11342 4521 11350 4592
rect 11266 4517 11350 4521
rect 10838 2767 10910 2770
rect 10838 2716 10851 2767
rect 10902 2716 10910 2767
rect 10838 2713 10910 2716
rect 10219 2598 10243 2621
rect 10219 2017 10242 2598
rect 10844 2012 10895 2713
rect 10830 2007 10895 2012
rect 10829 1989 10895 2007
rect 10826 1988 10895 1989
rect 10826 1982 10886 1988
rect 10826 1764 10860 1982
rect 10791 1665 10860 1764
rect 10826 1587 10860 1665
rect 10827 1526 10860 1587
rect 10826 1426 10860 1526
rect 10827 1366 10860 1426
rect 10082 719 10126 723
rect 10082 681 10084 719
rect 10122 681 10126 719
rect 10082 677 10126 681
rect 10826 622 10860 1366
rect 10827 562 10860 622
rect 10826 487 10860 562
rect 10877 1951 10886 1982
rect 10877 487 10884 1951
rect 10826 480 10884 487
rect 10826 479 10880 480
rect 6178 319 6270 392
rect 6175 246 6267 319
<< via1 >>
rect 203 7246 242 7285
rect 211 6901 250 6940
rect 349 6784 375 6810
rect 341 6514 383 6556
rect 936 6374 965 6432
rect 2265 6268 2291 6294
rect 2844 6225 2875 6256
rect 4502 6989 4544 7031
rect 4117 6913 4159 6955
rect 4669 6752 4713 6796
rect 5241 6752 5285 6796
rect 5423 6749 5467 6793
rect 4227 6650 4271 6694
rect 3951 6348 3977 6374
rect 3244 6279 3270 6305
rect 3127 6180 3154 6206
rect 1994 6102 2029 6137
rect 2519 6133 2545 6159
rect 4798 6650 4842 6694
rect 2096 5878 2122 5917
rect 3736 5879 3769 5905
rect 2032 5796 2058 5836
rect 2034 5685 2060 5711
rect 1657 5643 1683 5669
rect 1654 5551 1680 5577
rect 1655 5459 1681 5485
rect 1590 5357 1616 5383
rect 1586 5261 1612 5287
rect 1590 5165 1616 5191
rect 2034 5593 2060 5619
rect 2031 5501 2057 5527
rect 1586 3637 1612 3684
rect 1650 3637 1676 3684
rect 1450 3534 1476 3560
rect 1398 3494 1424 3520
rect 470 3369 536 3435
rect 1658 3532 1684 3558
rect 1834 3533 1861 3560
rect 1592 3496 1618 3522
rect 1400 3103 1426 3129
rect 991 2917 1028 2954
rect 474 2783 540 2849
rect 1884 3494 1910 3520
rect 990 2293 1027 2330
rect 1744 2251 1770 2287
rect 1289 1727 1318 1756
rect 3673 5707 3706 5740
rect 3616 5559 3649 5592
rect 2095 5392 2121 5418
rect 3552 5399 3585 5432
rect 3488 5342 3521 5375
rect 2096 5296 2122 5322
rect 2095 5200 2121 5226
rect 2031 3434 2057 3460
rect 1969 3319 1995 3345
rect 1927 3058 1953 3084
rect 1971 2489 1997 2531
rect 1967 2251 1993 2287
rect 3427 5185 3460 5218
rect 3364 5032 3397 5065
rect 3308 4875 3341 4908
rect 3246 4328 3279 4361
rect 3183 4169 3216 4202
rect 3121 4014 3154 4047
rect 3061 3866 3094 3899
rect 2997 3349 3030 3382
rect 2930 3192 2963 3225
rect 2095 3001 2121 3027
rect 2868 3028 2901 3061
rect 2029 1888 2055 1921
rect 1926 1726 1955 1755
rect 1810 1625 1870 1685
rect 2800 2884 2833 2917
rect 2396 2448 2454 2519
rect 2088 1132 2114 1166
rect 197 1038 236 1077
rect 2797 501 2840 544
rect 2862 422 2905 465
rect 2929 354 2969 394
rect 2912 260 2963 311
rect 6479 6913 6614 6955
rect 5937 6649 6032 6690
rect 6238 6650 6282 6694
rect 5663 6272 5689 6298
rect 5475 5919 5501 5945
rect 6022 6181 6048 6207
rect 5709 6079 5735 6105
rect 5751 5870 5777 5896
rect 5857 5822 5883 5848
rect 6339 6273 6365 6299
rect 6295 6182 6321 6208
rect 6021 5112 6048 5139
rect 6818 6646 6862 6690
rect 7651 6749 7679 6793
rect 7273 6083 7395 6109
rect 6949 6018 6975 6044
rect 7582 5964 7608 5990
rect 7816 6273 7842 6299
rect 7727 6186 7753 6212
rect 8468 7183 8505 7220
rect 8083 6344 8109 6371
rect 7727 5765 7753 5791
rect 7829 5766 7855 5792
rect 8104 5754 8147 5797
rect 5685 4448 5713 4476
rect 7420 4391 7446 4417
rect 8550 6837 8587 6874
rect 8469 4446 8506 4483
rect 8627 6366 8664 6403
rect 8546 4387 8583 4424
rect 9282 6261 9332 6311
rect 8960 6105 9010 6155
rect 9055 6154 9105 6204
rect 9163 6201 9213 6251
rect 8715 5859 8752 5896
rect 8620 4154 8657 4191
rect 4948 3629 4974 3670
rect 8713 3629 8750 3670
rect 5388 3257 5414 3283
rect 7376 3255 7402 3281
rect 4730 2744 4756 2770
rect 4676 2707 4705 2736
rect 4232 2656 4263 2687
rect 7324 3162 7350 3188
rect 5451 2979 5477 3005
rect 5391 2748 5417 2774
rect 5494 2747 5520 2773
rect 5251 2707 5277 2733
rect 5448 2715 5474 2741
rect 4613 2585 4655 2627
rect 4228 2489 4270 2531
rect 4819 2653 4845 2679
rect 7277 2978 7303 3004
rect 7227 2885 7253 2911
rect 5672 2709 5698 2735
rect 5552 2584 5585 2617
rect 6556 2740 6591 2775
rect 5871 2667 5897 2693
rect 6275 2664 6302 2691
rect 5667 2577 5701 2611
rect 6560 2563 6586 2595
rect 7159 2585 7185 2619
rect 4681 2480 4713 2512
rect 6702 2492 6740 2530
rect 5083 2005 5111 2033
rect 5157 2007 5185 2035
rect 4691 1902 4737 1948
rect 5529 1807 5575 1853
rect 6064 2005 6092 2033
rect 5672 1718 5718 1764
rect 10163 5967 10291 6095
rect 10595 5751 10621 5794
rect 10212 5623 10238 5665
rect 9812 5303 9852 5343
rect 9273 4033 9323 4083
rect 9165 3514 9215 3561
rect 9052 2995 9102 3045
rect 8947 2465 8997 2515
rect 7374 2314 7400 2364
rect 7320 2224 7346 2274
rect 7273 2134 7299 2184
rect 6511 1627 6557 1673
rect 3904 1404 3930 1516
rect 5115 1510 5227 1512
rect 5041 1400 5227 1510
rect 5041 1398 5153 1400
rect 6022 1395 6208 1514
rect 3736 975 3769 1008
rect 3674 913 3707 946
rect 3611 850 3644 883
rect 3551 787 3584 820
rect 3487 719 3520 752
rect 3427 657 3460 690
rect 3367 593 3400 626
rect 3309 536 3342 569
rect 3251 467 3284 500
rect 3186 403 3219 436
rect 3122 338 3155 372
rect 3064 274 3101 311
rect 7225 2044 7251 2094
rect 9571 2717 9621 2767
rect 9284 1906 9334 1956
rect 9165 1811 9215 1857
rect 9052 1724 9102 1770
rect 8959 1633 9009 1679
rect 9513 1404 9607 1516
rect 7092 1041 7125 1074
rect 9910 5239 9946 5275
rect 9818 922 9858 962
rect 10002 5002 10041 5041
rect 9909 842 9948 881
rect 10085 4946 10123 4972
rect 10002 760 10041 799
rect 11290 6500 11361 6571
rect 11271 4521 11342 4592
rect 10851 2716 10902 2767
rect 10084 681 10122 719
<< metal2 >>
rect 77 7277 145 7399
rect 200 7285 245 7287
rect 200 7277 203 7285
rect 77 7254 203 7277
rect 77 7167 145 7254
rect 200 7246 203 7254
rect 242 7246 245 7285
rect 200 7244 245 7246
rect 8462 7220 8508 7222
rect 11549 7220 11635 7355
rect 8462 7183 8468 7220
rect 8505 7183 11635 7220
rect 8462 7181 8508 7183
rect 11549 7145 11635 7183
rect 62 7057 310 7058
rect 62 7018 457 7057
rect 289 6981 457 7018
rect 2055 7048 2130 7049
rect 2055 7018 2217 7048
rect 4500 7031 4545 7033
rect 4499 7025 4502 7031
rect 2055 7001 2079 7018
rect 2187 6996 2217 7018
rect 2260 6995 4502 7025
rect 4499 6989 4502 6995
rect 4544 6989 4547 7031
rect 4500 6987 4545 6989
rect 4115 6955 4160 6957
rect 6476 6955 6618 6958
rect 77 6858 145 6946
rect 210 6940 253 6944
rect 210 6901 211 6940
rect 250 6901 253 6940
rect 4114 6913 4117 6955
rect 4159 6954 4162 6955
rect 6476 6954 6479 6955
rect 4159 6914 6479 6954
rect 4159 6913 4162 6914
rect 6476 6913 6479 6914
rect 6614 6954 6618 6955
rect 6614 6914 6623 6954
rect 6614 6913 6618 6914
rect 4115 6911 4160 6913
rect 6476 6910 6618 6913
rect 210 6897 253 6901
rect 210 6896 404 6897
rect 219 6874 404 6896
rect 8545 6874 8589 6876
rect 11549 6874 11635 6942
rect 77 6826 413 6858
rect 8545 6837 8550 6874
rect 8587 6837 11635 6874
rect 8545 6835 8589 6837
rect 77 6714 145 6826
rect 346 6784 349 6810
rect 375 6787 404 6810
rect 375 6784 378 6787
rect 4666 6752 4669 6796
rect 4713 6793 4716 6796
rect 5238 6793 5241 6796
rect 4713 6752 5241 6793
rect 5285 6793 5288 6796
rect 5285 6752 5423 6793
rect 4681 6749 5423 6752
rect 5467 6749 7651 6793
rect 7679 6749 7682 6793
rect 11549 6732 11635 6837
rect 4798 6694 4842 6697
rect 277 6677 430 6693
rect 96 6644 430 6677
rect 4224 6650 4227 6694
rect 4271 6692 4274 6694
rect 4271 6650 4798 6692
rect 6235 6692 6238 6694
rect 4842 6690 6238 6692
rect 4842 6650 5937 6690
rect 4239 6649 5937 6650
rect 6032 6650 6238 6690
rect 6282 6692 6285 6694
rect 6282 6690 6875 6692
rect 6282 6650 6818 6690
rect 6032 6649 6818 6650
rect 4239 6648 6818 6649
rect 4798 6647 4842 6648
rect 6815 6646 6818 6648
rect 6862 6648 6875 6690
rect 6862 6646 6865 6648
rect 96 6637 323 6644
rect 96 6617 136 6637
rect 61 6577 136 6617
rect 11287 6556 11290 6571
rect 338 6514 341 6556
rect 383 6514 11290 6556
rect 11287 6500 11290 6514
rect 11361 6500 11364 6571
rect 32 6432 100 6499
rect 924 6432 971 6434
rect 32 6374 936 6432
rect 965 6374 971 6432
rect 8623 6403 8665 6405
rect 11546 6403 11632 6533
rect 32 6350 104 6374
rect 924 6372 971 6374
rect 3949 6374 3979 6377
rect 32 6267 100 6350
rect 3949 6348 3951 6374
rect 3977 6371 3979 6374
rect 8081 6371 8111 6374
rect 3977 6348 8083 6371
rect 3949 6345 3979 6348
rect 8081 6344 8083 6348
rect 8109 6348 8118 6371
rect 8623 6366 8627 6403
rect 8664 6366 11632 6403
rect 8623 6364 8665 6366
rect 8109 6344 8111 6348
rect 8081 6340 8111 6344
rect 11546 6323 11632 6366
rect 3241 6305 3272 6307
rect 2262 6297 2294 6298
rect 3241 6297 3244 6305
rect 2262 6294 3244 6297
rect 2262 6268 2265 6294
rect 2291 6279 3244 6294
rect 3270 6297 3273 6305
rect 5659 6298 5691 6300
rect 6336 6299 6368 6300
rect 5659 6297 5663 6298
rect 3270 6279 5663 6297
rect 2291 6274 5663 6279
rect 2291 6268 2294 6274
rect 3241 6273 3272 6274
rect 5659 6272 5663 6274
rect 5689 6297 5692 6298
rect 6336 6297 6339 6299
rect 5689 6274 6339 6297
rect 5689 6272 5692 6274
rect 6336 6273 6339 6274
rect 6365 6297 6368 6299
rect 7813 6297 7816 6299
rect 6365 6274 7816 6297
rect 6365 6273 6368 6274
rect 7813 6273 7816 6274
rect 7842 6297 7845 6299
rect 9279 6297 9282 6311
rect 7842 6274 9282 6297
rect 7842 6273 7845 6274
rect 6336 6272 6368 6273
rect 2262 6266 2294 6268
rect 9279 6261 9282 6274
rect 9332 6261 9335 6311
rect 9279 6260 9335 6261
rect 2841 6256 2878 6258
rect 32 6217 83 6229
rect 2841 6225 2844 6256
rect 2875 6252 2878 6256
rect 9161 6252 9215 6254
rect 2875 6251 9215 6252
rect 2875 6229 9163 6251
rect 2875 6225 2878 6229
rect 2841 6223 2878 6225
rect 32 6188 342 6217
rect 6292 6208 6324 6209
rect 6021 6207 6049 6208
rect 83 6187 342 6188
rect 3124 6206 3155 6207
rect 6019 6206 6022 6207
rect 3124 6180 3127 6206
rect 3154 6183 6022 6206
rect 3154 6180 3157 6183
rect 6019 6181 6022 6183
rect 6048 6206 6051 6207
rect 6292 6206 6295 6208
rect 6048 6183 6295 6206
rect 6048 6181 6051 6183
rect 6292 6182 6295 6183
rect 6321 6206 6324 6208
rect 7724 6206 7727 6212
rect 6321 6186 7727 6206
rect 7753 6206 7756 6212
rect 9053 6206 9107 6207
rect 7753 6204 9107 6206
rect 7753 6186 9055 6204
rect 6321 6183 9055 6186
rect 6321 6182 6324 6183
rect 6292 6181 6324 6182
rect 6021 6180 6049 6181
rect 3124 6178 3155 6180
rect 2516 6160 2548 6161
rect 8959 6160 9012 6163
rect 2516 6159 9012 6160
rect 28 6137 79 6139
rect 1992 6137 2032 6138
rect 28 6102 1994 6137
rect 2029 6102 2032 6137
rect 2516 6133 2519 6159
rect 2545 6155 9012 6159
rect 2545 6137 8960 6155
rect 2545 6133 2548 6137
rect 2516 6131 2548 6133
rect 7271 6109 7399 6112
rect 28 6098 79 6102
rect 1992 6099 2032 6102
rect 5706 6105 5738 6106
rect 5706 6079 5709 6105
rect 5735 6102 5738 6105
rect 7271 6102 7273 6109
rect 5735 6083 7273 6102
rect 7395 6083 7399 6109
rect 8959 6105 8960 6137
rect 9010 6105 9012 6155
rect 9053 6154 9055 6183
rect 9105 6154 9107 6204
rect 9161 6201 9163 6229
rect 9213 6201 9215 6251
rect 9161 6198 9215 6201
rect 9053 6151 9107 6154
rect 8959 6102 9012 6105
rect 5735 6081 7399 6083
rect 5735 6079 5738 6081
rect 5706 6078 5738 6079
rect 0 5917 127 6063
rect 6948 6044 6976 6046
rect 6946 6018 6949 6044
rect 6975 6041 6978 6044
rect 10160 6041 10163 6095
rect 6975 6020 10163 6041
rect 6975 6018 6978 6020
rect 6948 6016 6976 6018
rect 7579 5990 7610 5993
rect 7579 5987 7582 5990
rect 4749 5986 7582 5987
rect 4716 5967 7582 5986
rect 4716 5966 4774 5967
rect 7579 5964 7582 5967
rect 7608 5964 7610 5990
rect 10160 5967 10163 6020
rect 10291 5967 10294 6095
rect 7579 5961 7610 5964
rect 5472 5940 5475 5945
rect 4972 5920 5475 5940
rect 1135 5917 1165 5918
rect 2094 5917 2123 5919
rect 0 5878 2096 5917
rect 2122 5878 2126 5917
rect 3733 5879 3736 5905
rect 3769 5896 3772 5905
rect 3769 5879 3906 5896
rect 0 5875 127 5878
rect 2094 5876 2123 5878
rect 2030 5836 2059 5838
rect 785 5796 2032 5836
rect 2058 5796 2061 5836
rect 4972 5832 4992 5920
rect 5472 5919 5475 5920
rect 5501 5940 5504 5945
rect 5501 5920 5509 5940
rect 5501 5919 5504 5920
rect 5748 5896 5779 5897
rect 8711 5896 8754 5898
rect 11546 5896 11632 6094
rect 5748 5893 5751 5896
rect 4748 5831 4992 5832
rect 4719 5812 4992 5831
rect 5023 5873 5751 5893
rect 4719 5811 4768 5812
rect 29 5527 156 5614
rect 785 5527 825 5796
rect 2030 5795 2059 5796
rect 3673 5742 3706 5743
rect 3671 5740 3708 5742
rect 1165 5728 1202 5729
rect 986 5705 1202 5728
rect 2031 5706 2034 5711
rect 986 5692 1728 5705
rect 986 5622 1048 5692
rect 1165 5688 1728 5692
rect 1974 5689 2034 5706
rect 2031 5685 2034 5689
rect 2060 5706 2063 5711
rect 3671 5707 3673 5740
rect 3706 5732 3708 5740
rect 3706 5715 3906 5732
rect 3706 5707 3708 5715
rect 2060 5689 2069 5706
rect 3671 5704 3708 5707
rect 2060 5685 2063 5689
rect 5023 5677 5043 5873
rect 5748 5870 5751 5873
rect 5777 5870 5780 5896
rect 5748 5869 5779 5870
rect 8711 5859 8715 5896
rect 8752 5884 11632 5896
rect 8752 5859 11621 5884
rect 8711 5856 8752 5859
rect 5854 5848 5886 5849
rect 5854 5845 5857 5848
rect 4748 5676 5043 5677
rect 1654 5643 1657 5669
rect 1683 5664 1686 5669
rect 1683 5647 1728 5664
rect 4719 5657 5043 5676
rect 5078 5825 5857 5845
rect 4719 5656 4769 5657
rect 1683 5643 1686 5647
rect 1165 5622 1202 5626
rect 29 5487 825 5527
rect 933 5613 1202 5622
rect 2031 5614 2034 5619
rect 933 5596 1728 5613
rect 1974 5597 2034 5614
rect 933 5585 1202 5596
rect 2031 5593 2034 5597
rect 2060 5614 2063 5619
rect 2060 5597 2069 5614
rect 2060 5593 2063 5597
rect 3613 5592 3652 5594
rect 933 5574 1048 5585
rect 933 5529 1044 5574
rect 1651 5551 1654 5577
rect 1680 5572 1683 5577
rect 1680 5555 1728 5572
rect 3613 5559 3616 5592
rect 3649 5584 3652 5592
rect 3649 5567 3906 5584
rect 3649 5559 3652 5567
rect 3613 5557 3652 5559
rect 1680 5551 1683 5555
rect 1165 5529 1202 5533
rect 933 5521 1202 5529
rect 2028 5522 2031 5527
rect 933 5504 1728 5521
rect 1974 5505 2031 5522
rect 933 5492 1202 5504
rect 2028 5501 2031 5505
rect 2057 5522 2060 5527
rect 5078 5522 5098 5825
rect 5854 5822 5857 5825
rect 5883 5845 5886 5848
rect 5883 5825 5894 5845
rect 5883 5822 5886 5825
rect 5854 5821 5886 5822
rect 7718 5794 7776 5809
rect 7718 5791 7730 5794
rect 7718 5765 7727 5791
rect 7762 5765 7776 5794
rect 7820 5793 7878 5808
rect 7820 5792 7833 5793
rect 7820 5766 7829 5792
rect 7718 5762 7730 5765
rect 7762 5762 7782 5765
rect 7718 5746 7782 5762
rect 7758 5685 7782 5746
rect 7820 5761 7833 5766
rect 7865 5761 7878 5793
rect 7820 5745 7878 5761
rect 8102 5797 8149 5800
rect 8102 5754 8104 5797
rect 8147 5794 8149 5797
rect 10592 5795 10621 5796
rect 10592 5794 10622 5795
rect 11645 5794 11690 5796
rect 8147 5754 10595 5794
rect 8102 5751 10595 5754
rect 10621 5751 11691 5794
rect 10592 5750 10622 5751
rect 10592 5748 10621 5750
rect 11595 5683 11631 5684
rect 10210 5665 10240 5667
rect 11539 5665 11631 5683
rect 2057 5505 2069 5522
rect 4749 5521 5098 5522
rect 2057 5501 2060 5505
rect 4719 5502 5098 5521
rect 5393 5645 5422 5663
rect 4719 5501 4765 5502
rect 933 5488 1023 5492
rect 29 5426 156 5487
rect 72 5033 199 5121
rect 933 5033 970 5488
rect 1652 5459 1655 5485
rect 1681 5480 1684 5485
rect 1681 5463 1728 5480
rect 1681 5459 1684 5463
rect 3549 5432 3588 5433
rect 1081 5419 1730 5421
rect 72 4996 970 5033
rect 1052 5402 1730 5419
rect 2092 5415 2095 5418
rect 1052 5384 1202 5402
rect 1971 5395 2095 5415
rect 2092 5392 2095 5395
rect 2121 5415 2124 5418
rect 2121 5395 2134 5415
rect 3549 5399 3552 5432
rect 3585 5424 3588 5432
rect 3585 5407 3906 5424
rect 3585 5399 3588 5407
rect 3549 5398 3588 5399
rect 2121 5392 2124 5395
rect 1052 5325 1118 5384
rect 1165 5380 1202 5384
rect 1587 5357 1590 5383
rect 1616 5379 1619 5383
rect 1616 5360 1730 5379
rect 3485 5375 3524 5378
rect 1616 5357 1619 5360
rect 3485 5342 3488 5375
rect 3521 5367 3524 5375
rect 3521 5350 3906 5367
rect 3521 5342 3524 5350
rect 3485 5340 3524 5342
rect 1052 5306 1730 5325
rect 2093 5319 2096 5322
rect 1052 5288 1202 5306
rect 1971 5299 2096 5319
rect 2093 5296 2096 5299
rect 2122 5319 2125 5322
rect 5393 5319 5411 5645
rect 10209 5623 10212 5665
rect 10238 5655 11631 5665
rect 10238 5623 11635 5655
rect 10210 5621 10240 5623
rect 11539 5589 11635 5623
rect 7828 5447 7888 5458
rect 7828 5413 7841 5447
rect 7875 5413 7888 5447
rect 8188 5441 8711 5464
rect 8748 5441 9663 5464
rect 11545 5446 11635 5589
rect 7828 5402 7888 5413
rect 9634 5431 9663 5441
rect 9634 5411 10546 5431
rect 9634 5410 9663 5411
rect 8189 5359 8711 5381
rect 8748 5359 9569 5381
rect 2122 5299 2134 5319
rect 5310 5301 5411 5319
rect 2122 5296 2125 5299
rect 1052 5287 1119 5288
rect 1052 5283 1118 5287
rect 1165 5284 1202 5288
rect 72 4933 199 4996
rect 66 4557 193 4646
rect 1052 4557 1089 5283
rect 1583 5261 1586 5287
rect 1612 5283 1615 5287
rect 1612 5264 1730 5283
rect 4749 5280 4779 5283
rect 4749 5279 4788 5280
rect 1612 5261 1615 5264
rect 4719 5259 4788 5279
rect 66 4520 1089 4557
rect 1165 5210 1730 5229
rect 2092 5223 2095 5226
rect 66 4458 193 4520
rect 72 4073 199 4164
rect 1165 4073 1202 5210
rect 1971 5203 2095 5223
rect 2092 5200 2095 5203
rect 2121 5223 2124 5226
rect 2121 5203 2134 5223
rect 3424 5218 3463 5220
rect 2121 5200 2124 5203
rect 1587 5165 1590 5191
rect 1616 5187 1619 5191
rect 1616 5168 1730 5187
rect 3424 5185 3427 5218
rect 3460 5210 3463 5218
rect 3460 5193 3906 5210
rect 3460 5185 3463 5193
rect 3424 5183 3463 5185
rect 1616 5165 1619 5168
rect 4746 5148 4779 5168
rect 5349 5156 5422 5174
rect 9547 5171 9569 5359
rect 9809 5343 9855 5346
rect 9809 5303 9812 5343
rect 9852 5333 9855 5343
rect 9852 5313 10546 5333
rect 10982 5313 11153 5333
rect 9852 5303 9855 5313
rect 9809 5301 9855 5303
rect 9910 5275 9946 5278
rect 11133 5268 11153 5313
rect 9946 5248 10546 5268
rect 10982 5248 11153 5268
rect 9910 5236 9946 5239
rect 9547 5170 9707 5171
rect 4746 5126 4764 5148
rect 5349 5135 5367 5156
rect 9547 5150 10546 5170
rect 9547 5149 9707 5150
rect 11133 5143 11153 5248
rect 11542 5143 11632 5210
rect 6019 5140 6050 5141
rect 4744 5124 4764 5126
rect 4719 5104 4764 5124
rect 5310 5117 5367 5135
rect 6018 5139 6051 5140
rect 6018 5134 6021 5139
rect 5983 5129 6021 5134
rect 5660 5112 6021 5129
rect 6048 5112 6051 5139
rect 8266 5113 8711 5129
rect 5660 5107 6050 5112
rect 8263 5109 8711 5113
rect 8748 5109 10546 5129
rect 7722 5100 7778 5109
rect 3361 5065 3403 5066
rect 3361 5032 3364 5065
rect 3397 5057 3403 5065
rect 7722 5065 7734 5100
rect 7767 5065 7778 5100
rect 3397 5040 3906 5057
rect 5359 5041 5414 5059
rect 7722 5055 7778 5065
rect 3397 5032 3403 5040
rect 3361 5031 3403 5032
rect 5359 5020 5377 5041
rect 5310 5002 5377 5020
rect 4744 4985 4779 4992
rect 4744 4969 4783 4985
rect 4725 4962 4783 4969
rect 4725 4949 4764 4962
rect 3305 4908 3344 4909
rect 3305 4875 3308 4908
rect 3341 4900 3344 4908
rect 3341 4883 3906 4900
rect 3341 4875 3344 4883
rect 3305 4874 3344 4875
rect 4753 4854 4779 4875
rect 8263 4861 8286 5109
rect 11133 5100 11632 5143
rect 10002 5042 10041 5044
rect 10001 5041 10042 5042
rect 10001 5002 10002 5041
rect 10041 5031 10042 5041
rect 11133 5031 11153 5100
rect 10041 5011 10546 5031
rect 10982 5011 11153 5031
rect 10041 5002 10042 5011
rect 10001 5001 10042 5002
rect 10002 4999 10041 5001
rect 10084 4972 10124 4973
rect 10082 4946 10085 4972
rect 10123 4966 10126 4972
rect 11133 4966 11153 5011
rect 11542 5001 11632 5100
rect 10123 4946 10546 4966
rect 10982 4954 11153 4966
rect 10982 4946 11150 4954
rect 10084 4945 10124 4946
rect 4753 4814 4773 4854
rect 7826 4844 7888 4853
rect 5310 4816 5387 4834
rect 4739 4794 4773 4814
rect 4753 4793 4773 4794
rect 5369 4572 5387 4816
rect 7826 4808 7843 4844
rect 7877 4808 7888 4844
rect 8188 4838 8286 4861
rect 8347 4848 8711 4868
rect 8748 4848 10546 4868
rect 7826 4800 7888 4808
rect 8347 4778 8367 4848
rect 8189 4763 8367 4778
rect 8189 4756 8364 4763
rect 11268 4592 11346 4595
rect 5369 4554 5423 4572
rect 11268 4521 11271 4592
rect 11342 4580 11346 4592
rect 11542 4580 11632 4672
rect 11342 4533 11632 4580
rect 11342 4521 11346 4533
rect 11268 4518 11346 4521
rect 8464 4483 8510 4485
rect 5683 4478 5715 4479
rect 8464 4478 8469 4483
rect 5683 4476 8469 4478
rect 5683 4448 5685 4476
rect 5713 4450 8469 4476
rect 5713 4448 5715 4450
rect 5683 4445 5715 4448
rect 8464 4446 8469 4450
rect 8506 4446 8510 4483
rect 11542 4463 11632 4533
rect 8464 4444 8510 4446
rect 8543 4424 8586 4426
rect 8543 4418 8546 4424
rect 7417 4417 8546 4418
rect 7417 4391 7420 4417
rect 7446 4392 8546 4417
rect 7446 4391 7449 4392
rect 8543 4387 8546 4392
rect 8583 4387 8586 4424
rect 8543 4385 8586 4387
rect 3244 4361 3281 4365
rect 3244 4328 3246 4361
rect 3279 4353 3281 4361
rect 3279 4336 3876 4353
rect 3279 4328 3281 4336
rect 3244 4325 3281 4328
rect 5386 4312 5564 4324
rect 5327 4306 5564 4312
rect 5327 4294 5411 4306
rect 4753 4276 4778 4278
rect 4753 4266 4779 4276
rect 4719 4246 4779 4266
rect 7540 4263 7596 4281
rect 3180 4202 3219 4203
rect 3180 4169 3183 4202
rect 3216 4194 3219 4202
rect 3216 4177 3876 4194
rect 8617 4191 8661 4193
rect 8617 4181 8620 4191
rect 3216 4169 3219 4177
rect 3180 4168 3219 4169
rect 7541 4163 8620 4181
rect 4738 4141 4776 4161
rect 8617 4154 8620 4163
rect 8657 4154 8661 4191
rect 8617 4153 8661 4154
rect 4738 4138 4775 4141
rect 4738 4111 4758 4138
rect 5388 4128 5564 4138
rect 4719 4091 4758 4111
rect 5328 4120 5564 4128
rect 5328 4110 5416 4120
rect 72 4036 1202 4073
rect 9270 4083 9330 4087
rect 72 3976 199 4036
rect 3118 4014 3121 4047
rect 3154 4039 3157 4047
rect 3154 4022 3876 4039
rect 9270 4033 9273 4083
rect 9323 4081 9330 4083
rect 11542 4081 11632 4184
rect 9323 4034 11632 4081
rect 9323 4033 9330 4034
rect 9270 4029 9330 4033
rect 3154 4014 3157 4022
rect 5389 4013 5564 4023
rect 5328 4005 5564 4013
rect 5328 3995 5416 4005
rect 4759 3956 4779 3984
rect 11542 3975 11632 4034
rect 4719 3936 4779 3956
rect 3057 3899 3099 3900
rect 3057 3866 3061 3899
rect 3094 3891 3099 3899
rect 3094 3874 3876 3891
rect 3094 3866 3099 3874
rect 3057 3864 3099 3866
rect 4759 3801 4779 3868
rect 5386 3827 5564 3838
rect 5328 3820 5564 3827
rect 5328 3809 5416 3820
rect 4719 3781 4779 3801
rect 66 3658 193 3742
rect 1583 3684 1614 3686
rect 1649 3684 1680 3686
rect 66 3621 1036 3658
rect 1583 3637 1586 3684
rect 1612 3637 1650 3684
rect 1676 3637 2315 3684
rect 1583 3635 1614 3637
rect 1649 3635 1680 3637
rect 66 3554 193 3621
rect 999 3486 1036 3621
rect 2268 3569 2315 3637
rect 4945 3670 4976 3672
rect 8709 3670 8754 3673
rect 4945 3629 4948 3670
rect 4974 3629 8713 3670
rect 8750 3629 8754 3670
rect 4945 3627 4976 3629
rect 8709 3627 8754 3629
rect 11545 3569 11635 3666
rect 1450 3560 1476 3563
rect 2268 3561 11635 3569
rect 1655 3556 1658 3558
rect 1476 3537 1658 3556
rect 1450 3531 1476 3534
rect 1655 3532 1658 3537
rect 1684 3556 1687 3558
rect 1831 3556 1834 3560
rect 1684 3537 1834 3556
rect 1684 3532 1687 3537
rect 1831 3533 1834 3537
rect 1861 3533 1864 3560
rect 2268 3522 9165 3561
rect 1395 3494 1398 3520
rect 1424 3516 1427 3520
rect 1589 3516 1592 3522
rect 1424 3497 1592 3516
rect 1424 3494 1427 3497
rect 1589 3496 1592 3497
rect 1618 3516 1621 3522
rect 1881 3516 1884 3520
rect 1618 3497 1884 3516
rect 1618 3496 1621 3497
rect 1881 3494 1884 3497
rect 1910 3494 1913 3520
rect 9161 3514 9165 3522
rect 9215 3522 11635 3561
rect 9215 3514 9218 3522
rect 9161 3510 9218 3514
rect 999 3485 1202 3486
rect 999 3467 1224 3485
rect 999 3461 1364 3467
rect 999 3449 1497 3461
rect 2029 3460 2059 3462
rect 2028 3458 2031 3460
rect 1165 3445 1497 3449
rect 1202 3439 1497 3445
rect 465 3435 542 3439
rect 465 3369 470 3435
rect 536 3420 542 3435
rect 1806 3436 2031 3458
rect 1165 3420 1204 3422
rect 536 3416 1204 3420
rect 536 3395 1496 3416
rect 536 3383 1203 3395
rect 1806 3392 1828 3436
rect 2028 3434 2031 3436
rect 2057 3434 2060 3460
rect 11545 3457 11635 3522
rect 2029 3432 2059 3434
rect 536 3369 542 3383
rect 1165 3381 1202 3383
rect 2993 3382 3034 3384
rect 465 3365 542 3369
rect 2993 3349 2997 3382
rect 3030 3374 3034 3382
rect 3030 3357 3876 3374
rect 3030 3349 3034 3357
rect 2993 3348 3034 3349
rect 1967 3345 1996 3347
rect 1966 3341 1969 3345
rect 72 3255 199 3332
rect 1809 3322 1969 3341
rect 1966 3319 1969 3322
rect 1995 3319 1998 3345
rect 5313 3328 5509 3346
rect 1967 3317 1996 3319
rect 4717 3269 4782 3289
rect 5393 3287 5510 3302
rect 5387 3283 5415 3287
rect 5387 3257 5388 3283
rect 5414 3257 5415 3283
rect 7373 3276 7376 3281
rect 6766 3260 7376 3276
rect 72 3218 671 3255
rect 5387 3254 5415 3257
rect 7373 3255 7376 3260
rect 7402 3255 7405 3281
rect 72 3144 199 3218
rect 634 3052 671 3218
rect 2927 3225 2966 3228
rect 2927 3192 2930 3225
rect 2963 3217 2966 3225
rect 2963 3200 3876 3217
rect 2963 3192 2966 3200
rect 2927 3190 2966 3192
rect 4755 3164 4780 3187
rect 7321 3183 7324 3188
rect 6767 3167 7324 3183
rect 4755 3134 4775 3164
rect 7321 3162 7324 3167
rect 7350 3162 7353 3188
rect 1398 3129 1427 3130
rect 1397 3103 1400 3129
rect 1426 3127 1429 3129
rect 1426 3105 1497 3127
rect 4719 3114 4775 3134
rect 5313 3142 5547 3160
rect 5313 3132 5331 3142
rect 1426 3103 1429 3105
rect 1398 3101 1427 3103
rect 1924 3084 1956 3086
rect 1924 3081 1927 3084
rect 1807 3060 1927 3081
rect 1924 3058 1927 3060
rect 1953 3058 1956 3084
rect 1924 3056 1956 3058
rect 2866 3063 2903 3064
rect 2866 3061 3876 3063
rect 634 3034 1229 3052
rect 634 3027 1236 3034
rect 1375 3027 1497 3028
rect 2093 3027 2122 3029
rect 2866 3028 2868 3061
rect 2901 3046 3876 3061
rect 2901 3028 2903 3046
rect 9049 3045 9104 3046
rect 634 3015 1497 3027
rect 2092 3024 2095 3027
rect 1165 3011 1497 3015
rect 1201 3006 1497 3011
rect 1807 3003 2095 3024
rect 988 2954 1029 2956
rect 1165 2954 1364 2956
rect 72 2841 199 2923
rect 988 2917 991 2954
rect 1028 2950 1364 2954
rect 1028 2928 1497 2950
rect 1028 2917 1203 2928
rect 1807 2921 1828 3003
rect 2092 3001 2095 3003
rect 2121 3001 2124 3027
rect 2866 3025 2903 3028
rect 5314 3027 5510 3045
rect 4756 3008 4776 3009
rect 2093 2999 2122 3001
rect 4756 2981 4785 3008
rect 5448 3005 5480 3007
rect 4756 2979 4776 2981
rect 4715 2959 4776 2979
rect 5448 2979 5451 3005
rect 5477 3002 5480 3005
rect 5477 2982 5509 3002
rect 7274 2999 7277 3004
rect 6766 2983 7277 2999
rect 5477 2979 5494 2982
rect 5448 2975 5494 2979
rect 7274 2978 7277 2983
rect 7303 2978 7306 3004
rect 9049 2995 9052 3045
rect 9102 3043 9105 3045
rect 11542 3043 11632 3158
rect 9102 2996 11632 3043
rect 9102 2995 9105 2996
rect 9049 2993 9104 2995
rect 11542 2949 11632 2996
rect 2797 2917 2836 2919
rect 988 2915 1029 2917
rect 1165 2915 1202 2917
rect 2797 2884 2800 2917
rect 2833 2909 2836 2917
rect 2833 2892 3876 2909
rect 7224 2906 7227 2911
rect 4754 2893 4784 2897
rect 2833 2884 2836 2892
rect 2797 2882 2836 2884
rect 4753 2869 4784 2893
rect 6772 2890 7227 2906
rect 7224 2885 7227 2890
rect 7253 2885 7256 2911
rect 465 2849 545 2855
rect 465 2841 474 2849
rect 72 2791 474 2841
rect 72 2735 199 2791
rect 465 2783 474 2791
rect 540 2783 545 2849
rect 4753 2824 4773 2869
rect 5314 2842 5543 2860
rect 4718 2804 4773 2824
rect 465 2778 545 2783
rect 6553 2775 6594 2776
rect 5388 2774 5420 2775
rect 4727 2744 4730 2770
rect 4756 2765 4759 2770
rect 5388 2765 5391 2774
rect 4756 2749 5391 2765
rect 4756 2744 4759 2749
rect 5388 2748 5391 2749
rect 5417 2748 5420 2774
rect 5388 2747 5420 2748
rect 5491 2773 5523 2774
rect 5491 2747 5494 2773
rect 5520 2765 5523 2773
rect 6553 2765 6556 2775
rect 5520 2749 6556 2765
rect 5520 2747 5523 2749
rect 5491 2746 5523 2747
rect 5447 2741 5475 2742
rect 4674 2736 4707 2738
rect 4673 2707 4676 2736
rect 4705 2728 4708 2736
rect 5248 2733 5280 2734
rect 5248 2728 5251 2733
rect 4705 2712 5251 2728
rect 4705 2707 4708 2712
rect 5248 2707 5251 2712
rect 5277 2707 5280 2733
rect 5445 2732 5448 2741
rect 5442 2716 5448 2732
rect 5445 2715 5448 2716
rect 5474 2732 5477 2741
rect 6553 2740 6556 2749
rect 6591 2740 6594 2775
rect 6553 2739 6594 2740
rect 9568 2767 9624 2769
rect 5669 2732 5672 2735
rect 5474 2716 5672 2732
rect 5474 2715 5477 2716
rect 5447 2714 5475 2715
rect 5669 2709 5672 2716
rect 5698 2709 5701 2735
rect 9568 2717 9571 2767
rect 9621 2762 9624 2767
rect 10840 2767 10908 2768
rect 10840 2762 10851 2767
rect 9621 2721 10851 2762
rect 9621 2717 9624 2721
rect 9568 2716 9624 2717
rect 10840 2716 10851 2721
rect 10902 2762 10908 2767
rect 11593 2762 11659 2826
rect 10902 2721 11659 2762
rect 10902 2716 10908 2721
rect 10840 2715 10908 2716
rect 11593 2711 11659 2721
rect 5671 2708 5699 2709
rect 4673 2705 4708 2707
rect 5870 2693 5898 2696
rect 4231 2687 4264 2690
rect 4231 2656 4232 2687
rect 4263 2666 4264 2687
rect 4817 2679 4847 2680
rect 4816 2666 4819 2679
rect 4263 2656 4819 2666
rect 4231 2653 4819 2656
rect 4845 2666 4848 2679
rect 5870 2667 5871 2693
rect 5897 2667 5898 2693
rect 5870 2666 5898 2667
rect 6273 2691 6303 2694
rect 6273 2666 6275 2691
rect 4845 2664 6275 2666
rect 6302 2664 6303 2691
rect 4845 2661 6302 2664
rect 4845 2653 6296 2661
rect 4231 2650 6296 2653
rect 4612 2628 4656 2629
rect 80 2627 4656 2628
rect 80 2586 4613 2627
rect 3927 2585 3975 2586
rect 4610 2585 4613 2586
rect 4655 2585 4658 2627
rect 5549 2617 5587 2620
rect 7157 2619 7187 2621
rect 4612 2584 4656 2585
rect 5549 2584 5552 2617
rect 5585 2584 5587 2617
rect 5549 2581 5587 2584
rect 5664 2577 5667 2611
rect 5701 2577 5704 2611
rect 6523 2595 6589 2597
rect 6523 2563 6560 2595
rect 6586 2563 6589 2595
rect 7086 2585 7159 2619
rect 7185 2585 7188 2619
rect 7157 2583 7188 2585
rect 6523 2561 6589 2563
rect 78 2489 1971 2531
rect 1997 2519 4228 2531
rect 1997 2489 2396 2519
rect 2383 2448 2396 2489
rect 2454 2489 4228 2519
rect 4270 2489 4276 2531
rect 6698 2530 6743 2532
rect 4679 2512 4717 2515
rect 2454 2448 2466 2489
rect 4679 2480 4681 2512
rect 4713 2480 4717 2512
rect 6698 2492 6702 2530
rect 6740 2492 6743 2530
rect 6698 2489 6743 2492
rect 8944 2515 9004 2518
rect 4679 2477 4717 2480
rect 8944 2465 8947 2515
rect 8997 2513 9004 2515
rect 11585 2513 11795 2607
rect 8997 2466 11795 2513
rect 8997 2465 9004 2466
rect 8944 2462 9004 2465
rect 2383 2439 2466 2448
rect 66 2330 193 2408
rect 11585 2399 11795 2466
rect 11587 2398 11664 2399
rect 989 2330 1030 2332
rect 66 2293 990 2330
rect 1027 2293 1030 2330
rect 7371 2314 7374 2364
rect 7400 2360 12954 2364
rect 7400 2314 13025 2360
rect 66 2220 193 2293
rect 989 2291 1030 2293
rect 1742 2287 1771 2289
rect 1965 2287 1996 2289
rect 1741 2251 1744 2287
rect 1770 2251 1967 2287
rect 1993 2251 1996 2287
rect 12415 2274 12616 2276
rect 1742 2249 1771 2251
rect 1965 2249 1996 2251
rect 7317 2224 7320 2274
rect 7346 2224 12616 2274
rect 7270 2134 7273 2184
rect 7299 2182 12197 2184
rect 7299 2134 12208 2182
rect 11573 2111 11574 2112
rect 7222 2044 7225 2094
rect 7251 2093 11801 2094
rect 7251 2044 11822 2093
rect 5081 2035 6171 2036
rect 5081 2033 5157 2035
rect 5080 2005 5083 2033
rect 5111 2008 5157 2033
rect 5111 2005 5114 2008
rect 5154 2007 5157 2008
rect 5185 2033 6171 2035
rect 5185 2008 6064 2033
rect 5185 2007 5188 2008
rect 6061 2005 6064 2008
rect 6092 2008 6171 2033
rect 6092 2005 6095 2008
rect 1161 1991 1198 1992
rect 72 1909 199 1979
rect 1029 1953 1282 1991
rect 4688 1954 4738 1955
rect 9281 1954 9284 1956
rect 1029 1909 1067 1953
rect 1161 1951 1198 1953
rect 4688 1948 9284 1954
rect 2028 1921 2056 1922
rect 72 1871 1067 1909
rect 1669 1888 2029 1921
rect 2055 1888 2058 1921
rect 4688 1902 4691 1948
rect 4737 1908 9284 1948
rect 4737 1902 4740 1908
rect 9281 1906 9284 1908
rect 9334 1906 9337 1956
rect 4688 1900 4738 1902
rect 2028 1886 2056 1888
rect 72 1791 199 1871
rect 5519 1857 9227 1863
rect 5519 1853 9165 1857
rect 5519 1817 5529 1853
rect 5526 1807 5529 1817
rect 5575 1817 9165 1853
rect 5575 1807 5578 1817
rect 9162 1811 9165 1817
rect 9215 1817 9227 1857
rect 9215 1811 9218 1817
rect 5663 1770 9118 1772
rect 5663 1765 9052 1770
rect 5662 1764 9052 1765
rect 1286 1727 1289 1756
rect 1318 1753 1321 1756
rect 1924 1755 1957 1759
rect 1923 1753 1926 1755
rect 1318 1727 1926 1753
rect 1290 1726 1926 1727
rect 1955 1753 1958 1755
rect 1955 1726 2289 1753
rect 1290 1724 2289 1726
rect 1924 1722 1957 1724
rect 1670 1685 1904 1690
rect 1670 1630 1810 1685
rect 1807 1625 1810 1630
rect 1870 1656 1904 1685
rect 1870 1632 1908 1656
rect 1870 1630 1904 1632
rect 1870 1625 1873 1630
rect 1807 1623 1873 1625
rect 1810 1622 1870 1623
rect 2259 1516 2288 1724
rect 5662 1718 5672 1764
rect 5718 1726 9052 1764
rect 5718 1718 5727 1726
rect 9049 1724 9052 1726
rect 9102 1726 9118 1770
rect 9102 1724 9105 1726
rect 5662 1713 5727 1718
rect 6507 1678 6559 1680
rect 8956 1678 8959 1679
rect 6507 1673 8959 1678
rect 6507 1627 6511 1673
rect 6557 1633 8959 1673
rect 9009 1678 9012 1679
rect 9009 1633 9021 1678
rect 6557 1632 9021 1633
rect 6557 1627 6560 1632
rect 6507 1622 6559 1627
rect 3901 1516 3933 1518
rect 9501 1516 9617 1519
rect 72 1386 199 1477
rect 2240 1404 3904 1516
rect 3930 1514 9513 1516
rect 3930 1512 6022 1514
rect 3930 1510 5115 1512
rect 3930 1404 5041 1510
rect 3901 1402 3933 1404
rect 5038 1398 5041 1404
rect 5227 1404 6022 1512
rect 5227 1400 5230 1404
rect 5153 1398 5230 1400
rect 5038 1396 5230 1398
rect 6019 1395 6022 1404
rect 6208 1404 9513 1514
rect 9607 1404 9617 1516
rect 6208 1395 6212 1404
rect 9501 1401 9617 1404
rect 6019 1393 6212 1395
rect 72 1348 1069 1386
rect 72 1289 199 1348
rect 1031 1263 1069 1348
rect 1161 1263 1198 1264
rect 1031 1225 1303 1263
rect 1161 1223 1198 1225
rect 2086 1166 2117 1168
rect 1663 1132 2088 1166
rect 2114 1132 2117 1166
rect 2086 1130 2117 1132
rect 193 1077 243 1082
rect 193 1038 197 1077
rect 236 1071 243 1077
rect 7090 1074 7129 1075
rect 7089 1071 7092 1074
rect 236 1043 7092 1071
rect 236 1038 243 1043
rect 7089 1041 7092 1043
rect 7125 1041 7129 1074
rect 7090 1040 7129 1041
rect 193 1035 243 1038
rect 3731 1008 3773 1009
rect 3731 975 3736 1008
rect 3769 983 7758 1008
rect 3769 975 7759 983
rect 3731 974 3773 975
rect 7155 973 7759 975
rect 3671 946 3709 947
rect 59 735 186 923
rect 3671 913 3674 946
rect 3707 913 7351 946
rect 3671 912 3709 913
rect 6744 912 7351 913
rect 3607 883 3649 884
rect 3607 850 3611 883
rect 3644 850 6943 883
rect 3607 849 3649 850
rect 3548 820 3588 821
rect 3548 787 3551 820
rect 3584 819 3588 820
rect 3584 787 6542 819
rect 3548 786 6542 787
rect 3548 785 3588 786
rect 3482 752 3523 753
rect 3481 719 3487 752
rect 3520 719 6133 752
rect 3482 717 3523 719
rect 3424 690 3465 691
rect 3424 657 3427 690
rect 3460 688 5731 690
rect 3460 657 5732 688
rect 3424 656 3465 657
rect 3364 593 3367 626
rect 3400 625 3403 626
rect 3400 593 5333 625
rect 3374 592 5333 593
rect 2792 544 2846 547
rect 2792 543 2797 544
rect 1509 539 2797 543
rect 1504 501 2797 539
rect 2840 501 2846 544
rect 3306 536 3309 569
rect 3342 564 3345 569
rect 3342 536 4942 564
rect 3332 531 4942 536
rect 1504 500 2846 501
rect 66 260 193 448
rect 1504 312 1705 500
rect 2792 497 2846 500
rect 3248 467 3251 500
rect 3284 467 4522 500
rect 2857 465 2911 466
rect 2857 459 2862 465
rect 1914 422 2862 459
rect 2905 422 2911 465
rect 3909 437 4111 439
rect 3193 436 4111 437
rect 1914 416 2911 422
rect 1914 315 2112 416
rect 3183 403 3186 436
rect 3219 404 4111 436
rect 3219 403 3222 404
rect 2925 394 2974 398
rect 2925 378 2929 394
rect 2364 376 2929 378
rect 2307 354 2929 376
rect 2969 354 2974 394
rect 2307 348 2974 354
rect 2307 338 2965 348
rect 3119 338 3122 372
rect 3155 338 3717 372
rect 2307 315 2505 338
rect 2908 315 2973 316
rect 1502 246 1705 312
rect 1909 249 2112 315
rect 2305 249 2508 315
rect 2705 311 2973 315
rect 2705 260 2912 311
rect 2963 260 2973 311
rect 3058 313 3113 315
rect 3516 313 3717 338
rect 3058 311 3313 313
rect 3683 312 3717 313
rect 3058 274 3064 311
rect 3101 274 3313 311
rect 3058 270 3313 274
rect 2705 252 2973 260
rect 2705 249 2908 252
rect 3110 247 3313 270
rect 3513 294 3717 312
rect 3907 316 4111 404
rect 3907 315 4109 316
rect 3907 308 4112 315
rect 4317 314 4520 467
rect 4317 313 4519 314
rect 4317 308 4521 313
rect 3513 246 3716 294
rect 3909 249 4112 308
rect 4318 247 4521 308
rect 4735 249 4938 531
rect 5134 321 5333 592
rect 5133 246 5336 321
rect 5532 319 5732 657
rect 5529 249 5732 319
rect 5942 312 6133 719
rect 6346 314 6541 786
rect 6744 314 6943 850
rect 7155 880 7351 912
rect 7565 923 7759 973
rect 9817 962 9860 964
rect 7967 959 8163 962
rect 9815 959 9818 962
rect 7967 924 9818 959
rect 7155 314 7350 880
rect 7565 316 7758 923
rect 5934 247 6137 312
rect 6341 249 6544 314
rect 6744 249 6947 314
rect 7149 249 7352 314
rect 7556 238 7759 316
rect 7967 314 8163 924
rect 9815 922 9818 924
rect 9858 922 9861 962
rect 9817 921 9860 922
rect 9907 881 9950 883
rect 9906 880 9909 881
rect 8360 842 9909 880
rect 9948 842 9951 881
rect 7964 249 8167 314
rect 8360 312 8556 842
rect 9907 840 9950 842
rect 9999 798 10002 799
rect 8775 760 10002 798
rect 10041 760 10044 799
rect 8775 314 8973 760
rect 10083 719 10125 722
rect 9186 681 10084 719
rect 10122 681 10125 719
rect 8359 247 8562 312
rect 8771 249 8974 314
rect 9186 311 9384 681
rect 10083 678 10125 681
rect 9693 382 10317 402
rect 9693 314 9713 382
rect 10409 361 10429 402
rect 10186 341 10429 361
rect 10186 314 10206 341
rect 10506 314 10527 403
rect 9185 246 9388 311
rect 9584 249 9787 314
rect 9986 284 10206 314
rect 9986 249 10189 284
rect 10394 249 10597 314
rect 10699 305 10720 403
rect 10796 384 10815 401
rect 10796 365 11296 384
rect 10812 305 11015 314
rect 11277 312 11296 365
rect 11361 312 11380 319
rect 11621 314 11822 2044
rect 10699 284 11015 305
rect 10812 249 11015 284
rect 11210 247 11413 312
rect 11615 262 11822 314
rect 12007 314 12208 2134
rect 11615 249 11818 262
rect 12007 249 12214 314
rect 12415 312 12616 2224
rect 12824 314 13025 2314
rect 12007 245 12208 249
rect 12415 247 12619 312
rect 12821 256 13025 314
rect 12821 249 13024 256
rect 12415 239 12616 247
<< via2 >>
rect 7730 5791 7762 5794
rect 7730 5765 7753 5791
rect 7753 5765 7762 5791
rect 7833 5792 7865 5793
rect 7833 5766 7855 5792
rect 7855 5766 7865 5792
rect 7730 5762 7762 5765
rect 7833 5761 7865 5766
rect 7841 5413 7875 5447
rect 7734 5065 7767 5100
rect 7843 4808 7877 4844
<< metal3 >>
rect 7723 5794 7768 5800
rect 7723 5762 7730 5794
rect 7762 5762 7768 5794
rect 7723 5725 7768 5762
rect 7827 5793 7872 5799
rect 7827 5761 7833 5793
rect 7865 5761 7872 5793
rect 7723 5109 7760 5725
rect 7827 5724 7872 5761
rect 7835 5460 7872 5724
rect 7835 5447 7879 5460
rect 7835 5413 7841 5447
rect 7875 5413 7879 5447
rect 7835 5400 7879 5413
rect 7723 5100 7772 5109
rect 7723 5076 7734 5100
rect 7728 5065 7734 5076
rect 7767 5065 7772 5100
rect 7728 5060 7772 5065
rect 7835 4889 7872 5400
rect 7834 4844 7881 4889
rect 7834 4808 7843 4844
rect 7877 4808 7881 4844
rect 7834 4802 7881 4808
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_0
timestamp 1608245216
transform -1 0 1794 0 -1 2112
box 64 419 528 1018
use sky130_hilas_nFETLarge  sky130_hilas_nFETLarge_0
timestamp 1625426387
transform -1 0 1790 0 -1 2867
box 64 420 501 1003
use sky130_hilas_DAC5bit01  sky130_hilas_DAC5bit01_0
timestamp 1625056879
transform 0 1 9694 1 0 0
box 382 524 2040 1121
use sky130_hilas_Trans2med  sky130_hilas_Trans2med_0
timestamp 1626027626
transform 1 0 1855 0 -1 3342
box -380 -143 -27 452
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_3
timestamp 1624113741
transform -1 0 4709 0 -1 3294
box -30 -102 850 522
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_3
timestamp 1625970648
transform -1 0 6383 0 -1 3393
box 1050 5 1622 610
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_1
timestamp 1608245216
transform 1 0 4606 0 1 1637
box 64 419 528 1018
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_2
timestamp 1608245216
transform -1 0 5662 0 1 1637
box 64 419 528 1018
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_3
timestamp 1608245216
transform 1 0 5587 0 1 1640
box 64 419 528 1018
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_4
timestamp 1608245216
transform -1 0 6643 0 1 1640
box 64 419 528 1018
use sky130_hilas_WTA4Stage01  sky130_hilas_WTA4Stage01_0
timestamp 1625404155
transform 1 0 6607 0 1 2834
box -1121 -43 296 562
use sky130_hilas_nFETLarge  sky130_hilas_nFETLarge_1
timestamp 1625426387
transform -1 0 7217 0 1 1639
box 64 420 501 1003
use sky130_hilas_Trans4small  sky130_hilas_Trans4small_0
timestamp 1608234847
transform 1 0 1520 0 1 5290
box 191 -150 471 438
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_2
timestamp 1624113741
transform -1 0 4709 0 -1 4271
box -30 -102 850 522
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_1
timestamp 1624113741
transform -1 0 4709 0 -1 5284
box -30 -102 850 522
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_2
timestamp 1625970648
transform -1 0 6383 0 -1 4369
box 1050 5 1622 610
use sky130_hilas_swc4x2cell  sky130_hilas_swc4x2cell_0
timestamp 1625491916
transform 1 0 6550 0 1 3773
box -1004 -4 1009 601
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_1
timestamp 1625970648
transform -1 0 6383 0 -1 5376
box 1050 5 1622 610
use sky130_hilas_TA2Cell_1FG  sky130_hilas_TA2Cell_1FG_0
timestamp 1625491133
transform 1 0 8018 0 1 4364
box -2616 140 193 745
use sky130_hilas_TA2Cell_1FG_Strong  sky130_hilas_TA2Cell_1FG_Strong_0
timestamp 1626460134
transform 1 0 8018 0 1 4967
box -2617 140 193 745
use sky130_hilas_Tgate4Single01  sky130_hilas_Tgate4Single01_0
timestamp 1608226321
transform 1 0 10562 0 1 4978
box -36 -141 440 464
use sky130_hilas_FGcharacterization01  sky130_hilas_FGcharacterization01_0
timestamp 1625074044
transform -1 0 2464 0 1 6339
box -912 259 2083 864
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_0
timestamp 1624113741
transform -1 0 4709 0 1 5496
box -30 -102 850 522
<< labels >>
rlabel metal2 12821 249 13024 314 1 DIG24 
port 1 n
rlabel metal2 12416 247 12619 312 0 DIG23
port 2 nsew
rlabel metal2 12011 249 12214 314 0 DIG22
port 3 nsew
rlabel metal2 11615 249 11818 314 0 DIG21
port 4 nsew
rlabel metal2 11210 247 11413 312 0 DIG29
port 5 nsew
rlabel metal2 10812 249 11015 314 0 DIG28
port 6 nsew
rlabel metal2 10394 249 10597 314 0 DIG27
port 7 nsew
rlabel metal2 9986 249 10189 314 0 DIG26
port 8 nsew
rlabel metal2 9584 249 9787 314 0 DIG25
port 9 nsew
rlabel metal2 9185 246 9388 311 0 DIG20
port 10 nsew
rlabel metal2 8771 249 8974 314 0 DIG19
port 11 nsew
rlabel metal2 8359 247 8562 312 0 DIG18
port 12 nsew
rlabel metal2 7964 249 8167 314 0 DIG17
port 13 nsew
rlabel metal2 7556 251 7759 316 0 DIG16
port 14 nsew
rlabel metal2 7149 249 7352 314 0 DIG15
port 15 nsew
rlabel metal2 6744 249 6947 314 0 DIG14
port 16 nsew
rlabel metal2 6341 249 6544 314 0 DIG13
port 17 nsew
rlabel metal2 5934 247 6137 312 0 DIG12
port 18 nsew
rlabel metal2 5529 253 5732 319 0 DIG11
port 19 nsew
rlabel metal2 5133 255 5336 321 0 DIG10
port 20 nsew
rlabel metal2 4735 249 4938 315 0 DIG09
port 21 nsew
rlabel metal2 4318 247 4521 313 0 DIG08
port 22 nsew
rlabel metal2 3909 249 4112 315 0 DIG07
port 23 nsew
rlabel metal2 3513 246 3716 312 0 DIG06
port 24 nsew
rlabel metal2 3110 247 3313 313 0 DIG05
port 25 nsew
rlabel metal2 2705 249 2908 315 0 DIG04
port 26 nsew
rlabel metal2 2305 249 2508 315 0 DIG03
port 27 nsew
rlabel metal2 1909 249 2112 315 0 DIG02
port 28 nsew
rlabel metal2 1502 246 1705 312 0 DIG01
port 29 nsew
rlabel metal2 11587 2398 11664 2607 0 CAP2    
port 30 nsew
rlabel metal2 11542 2949 11632 3158 0 GENERALGATE01   
port 31 nsew
rlabel metal2 11545 3457 11635 3666 0 GATEANDCAP1    
port 32 nsew
rlabel metal2 11542 3975 11632 4184 0 GENERALGATE02
port 33 nsew
rlabel metal2 11542 4463 11632 4672 0 OUTPUTTA1    
port 34 nsew
rlabel metal2 11542 5001 11632 5210 0 GATENFET1   
port 35 nsew
rlabel metal2 11545 5446 11635 5655 0 DACOUTPUT  
port 36 nsew
rlabel metal2 11546 5884 11632 6094 0 DRAINOUT
port 37 nsew
rlabel metal2 11546 6323 11632 6533 0 ROWTERM2
port 38 nsew
rlabel metal2 11549 6732 11635 6942 0 COLUMN2
port 39 nsew
rlabel metal2 11549 7145 11635 7355 0 COLUMN1
port 40 nsew
rlabel metal1 10055 7318 10374 7430 0 GATE2
port 41 nsew
rlabel metal1 7198 7315 7517 7427 0 GATE1
port 61 nsew
rlabel metal1 4339 7316 4658 7428 0 DRAININJECT
port 42 nsew
rlabel metal1 2808 7269 2942 7370 0 VTUN
port 43 nsew
rlabel metal2 77 7167 145 7399 0 VREFCHAR
port 44 nsew
rlabel metal2 77 6714 145 6946 0 CHAROUTPUT
port 45 nsew
rlabel metal2 32 6267 100 6499 0 LARGECAPACITOR
port 46 nsew
rlabel metal2 1161 1951 1198 1992 0 DRAIN6N
port 47 nsew
rlabel metal2 1161 1223 1198 1264 0 DRAIN6P
port 48 nsew
rlabel metal2 1165 2915 1202 2956 0 DRAIN5P
port 49 nsew
rlabel metal2 1165 3011 1202 3052 0 DARIN4P
port 50 nsew
rlabel metal2 1165 3381 1202 3422 0 DRAIN5N
port 51 nsew
rlabel metal2 1165 3445 1202 3486 0 DRAIN4N
port 52 nsew
rlabel metal2 1165 5188 1202 5229 0 DRAIN3P
port 53 nsew
rlabel metal2 1165 5284 1202 5325 0 DRAIN2P
port 54 nsew
rlabel metal2 1165 5380 1202 5421 0 DRAIN1P
port 55 nsew
rlabel metal2 1165 5492 1202 5533 0 DRAIN3N
port 56 nsew
rlabel metal2 1165 5585 1202 5626 0 DRAIN2N
port 57 nsew
rlabel metal2 1165 5688 1202 5729 0 DRAIN1N
port 58 nsew
rlabel metal2 1135 5796 1165 5836 0 SOURCEN
port 59 nsew
rlabel metal2 1135 5878 1165 5918 0 SOURCEP
port 60 nsew
rlabel metal2 61 6577 106 6617 0 VGND
port 63 nsew
rlabel metal2 65 7018 110 7058 0 VINJ
port 62 nsew
rlabel metal2 32 6188 83 6229 0 VINJ
port 62 nsew
rlabel metal2 28 6098 79 6139 0 VGND
port 63 nsew
rlabel metal2 80 2586 143 2628 0 VINJ
port 62 nsew
rlabel metal2 78 2489 141 2531 0 VGND
port 63 nsew
rlabel metal2 11645 5751 11690 5796 0 VPWR
port 64 nsew
rlabel metal1 5420 7402 5493 7432 0 VINJ
port 62 nsew
rlabel metal1 5936 7411 6033 7432 0 VGND
port 63 nsew
rlabel metal2 11593 2711 11659 2826 0 VPWR
port 64 nsew
rlabel metal1 4982 246 5074 319 0 VPWR
port 64 nsew
rlabel metal1 6175 246 6267 319 0 VPWR
port 64 nsew
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
