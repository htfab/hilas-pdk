magic
tech sky130A
timestamp 1608072649
<< metal2 >>
rect 1417 480 1992 498
rect 1417 437 1992 455
rect 1417 385 1444 413
rect 1957 385 1992 413
rect 1417 337 1992 355
rect 1417 294 1992 312
rect 1417 179 1992 196
rect 1417 137 1992 154
rect 1417 85 1445 113
rect 1957 85 1993 113
rect 1417 39 1992 56
rect 1417 -5 1992 12
<< metal3 >>
rect 1801 359 1904 434
rect 1800 60 1906 133
<< metal4 >>
rect 1441 365 1720 406
rect 1472 64 1684 105
use sky130_hilas_m22m4  sky130_hilas_m22m4_4
timestamp 1607701799
transform 1 0 1938 0 1 95
box -36 -36 43 39
use sky130_hilas_m22m4  sky130_hilas_m22m4_3
timestamp 1607701799
transform 1 0 1938 0 1 395
box -36 -36 43 39
use sky130_hilas_m22m4  sky130_hilas_m22m4_5
timestamp 1607701799
transform 1 0 1454 0 1 95
box -36 -36 43 39
use sky130_hilas_m22m4  sky130_hilas_m22m4_2
timestamp 1607701799
transform 1 0 1451 0 1 395
box -36 -36 43 39
use sky130_hilas_CapModule01a  sky130_hilas_CapModule01a_0
timestamp 1607818356
transform 1 0 2002 0 1 198
box -416 -216 -186 12
use sky130_hilas_CapModule01a  sky130_hilas_CapModule01a_1
timestamp 1607818356
transform 1 0 2002 0 1 499
box -416 -216 -186 12
<< labels >>
rlabel metal2 1982 385 1992 413 0 Cap1Term02
port 1 nsew analog default
rlabel metal2 1417 385 1424 413 0 Cap1Term01
port 4 nsew analog default
rlabel metal2 1417 85 1423 113 0 Cap2Term01
port 3 nsew analog default
rlabel metal2 1986 85 1993 113 0 Cap2Term02
port 2 nsew analog default
<< end >>
