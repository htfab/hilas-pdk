magic
tech sky130A
timestamp 1607258550
<< error_s >>
rect 267 230 296 258
rect 346 230 375 258
rect 425 230 454 258
rect 245 223 475 230
rect 245 208 252 223
rect 267 217 296 223
rect 346 217 375 223
rect 425 217 454 223
rect 267 208 268 209
rect 295 208 296 209
rect 346 208 347 209
rect 374 208 375 209
rect 425 208 426 209
rect 453 208 454 209
rect 468 208 475 223
rect 217 179 258 208
rect 266 207 297 208
rect 345 207 376 208
rect 424 207 455 208
rect 267 180 296 207
rect 346 180 375 207
rect 425 180 454 207
rect 266 179 297 180
rect 345 179 376 180
rect 424 179 455 180
rect 462 179 504 208
rect -206 150 -200 156
rect -153 150 -147 156
rect 245 129 252 179
rect 267 178 268 179
rect 295 178 296 179
rect 346 178 347 179
rect 374 178 375 179
rect 425 178 426 179
rect 453 178 454 179
rect 468 151 475 179
rect 267 129 268 130
rect 295 129 296 130
rect 346 129 347 130
rect 374 129 375 130
rect 425 129 426 130
rect 453 129 454 130
rect 468 129 475 135
rect 488 134 489 135
rect -212 100 -206 106
rect -147 100 -141 106
rect 217 100 258 129
rect 266 128 297 129
rect 345 128 376 129
rect 424 128 455 129
rect 267 101 296 128
rect 346 101 375 128
rect 425 101 454 128
rect 266 100 297 101
rect 345 100 376 101
rect 424 100 455 101
rect 462 100 504 129
rect 245 91 252 100
rect 267 99 268 100
rect 295 99 296 100
rect 346 99 347 100
rect 374 99 375 100
rect 425 99 426 100
rect 453 99 454 100
rect 258 91 462 94
rect 468 91 475 100
rect 245 78 475 91
rect 267 77 296 78
rect 346 77 375 78
rect 425 77 454 78
rect 245 70 475 77
rect 245 55 252 70
rect 267 64 296 70
rect 346 64 375 70
rect 425 64 454 70
rect 306 56 332 62
rect 267 55 268 56
rect 295 55 296 56
rect 346 55 347 56
rect 374 55 375 56
rect 425 55 426 56
rect 453 55 454 56
rect 468 55 475 70
rect -206 41 -200 47
rect -153 41 -147 47
rect 217 26 258 55
rect 266 54 297 55
rect 345 54 376 55
rect 424 54 455 55
rect 267 27 296 54
rect 307 42 333 48
rect 346 27 375 54
rect 425 27 454 54
rect 266 26 297 27
rect 345 26 376 27
rect 424 26 455 27
rect 462 26 504 55
rect -212 -9 -206 -3
rect -147 -9 -141 -3
rect 245 -24 252 26
rect 267 25 268 26
rect 295 25 296 26
rect 346 25 347 26
rect 374 25 375 26
rect 425 25 426 26
rect 453 25 454 26
rect 468 8 475 26
rect 267 -24 268 -23
rect 295 -24 296 -23
rect 346 -24 347 -23
rect 374 -24 375 -23
rect 425 -24 426 -23
rect 453 -24 454 -23
rect 468 -24 475 -9
rect 217 -53 258 -24
rect 266 -25 297 -24
rect 345 -25 376 -24
rect 424 -25 455 -24
rect 267 -52 296 -25
rect 346 -52 375 -25
rect 425 -52 454 -25
rect 266 -53 297 -52
rect 345 -53 376 -52
rect 424 -53 455 -52
rect 462 -53 504 -24
rect 245 -65 252 -53
rect 267 -54 268 -53
rect 295 -54 296 -53
rect 346 -54 347 -53
rect 374 -54 375 -53
rect 425 -54 426 -53
rect 453 -54 454 -53
rect 266 -65 296 -62
rect 345 -65 375 -62
rect 424 -65 454 -62
rect 468 -65 475 -53
rect 245 -75 475 -65
rect 266 -79 296 -75
rect 345 -79 375 -75
rect 424 -79 454 -75
rect 244 -86 474 -79
rect 244 -101 251 -86
rect 266 -92 296 -86
rect 345 -92 375 -86
rect 424 -92 454 -86
rect 306 -97 332 -94
rect 266 -101 267 -100
rect 294 -101 295 -100
rect 345 -101 346 -100
rect 373 -101 374 -100
rect 424 -101 425 -100
rect 452 -101 453 -100
rect 467 -101 474 -86
rect 216 -130 257 -101
rect 265 -102 296 -101
rect 344 -102 375 -101
rect 423 -102 454 -101
rect 266 -129 295 -102
rect 306 -111 332 -108
rect 345 -129 374 -102
rect 424 -129 453 -102
rect 265 -130 296 -129
rect 344 -130 375 -129
rect 423 -130 454 -129
rect 461 -130 503 -101
rect -206 -148 -200 -142
rect -153 -148 -147 -142
rect 244 -180 251 -130
rect 266 -131 267 -130
rect 294 -131 295 -130
rect 345 -131 346 -130
rect 373 -131 374 -130
rect 424 -131 425 -130
rect 452 -131 453 -130
rect 467 -150 474 -130
rect 266 -180 267 -179
rect 294 -180 295 -179
rect 345 -180 346 -179
rect 373 -180 374 -179
rect 424 -180 425 -179
rect 452 -180 453 -179
rect 467 -180 474 -167
rect -212 -198 -206 -192
rect -147 -198 -141 -192
rect 216 -209 257 -180
rect 265 -181 296 -180
rect 344 -181 375 -180
rect 423 -181 454 -180
rect 266 -208 295 -181
rect 345 -208 374 -181
rect 424 -208 453 -181
rect 265 -209 296 -208
rect 344 -209 375 -208
rect 423 -209 454 -208
rect 461 -209 503 -180
rect 244 -219 251 -209
rect 266 -210 267 -209
rect 294 -210 295 -209
rect 345 -210 346 -209
rect 373 -210 374 -209
rect 424 -210 425 -209
rect 452 -210 453 -209
rect 257 -218 461 -216
rect 266 -219 295 -218
rect 345 -219 374 -218
rect 424 -219 453 -218
rect 467 -219 474 -209
rect 244 -231 474 -219
rect 266 -233 295 -231
rect 345 -233 374 -231
rect 424 -233 453 -231
rect 244 -240 474 -233
rect 244 -255 251 -240
rect 266 -246 295 -240
rect 345 -246 374 -240
rect 424 -246 453 -240
rect 305 -253 331 -248
rect 266 -255 267 -254
rect 294 -255 295 -254
rect 345 -255 346 -254
rect 373 -255 374 -254
rect 424 -255 425 -254
rect 452 -255 453 -254
rect 467 -255 474 -240
rect -206 -265 -200 -259
rect -153 -265 -147 -259
rect 216 -284 257 -255
rect 265 -256 296 -255
rect 344 -256 375 -255
rect 423 -256 454 -255
rect 266 -283 295 -256
rect 306 -267 332 -262
rect 345 -283 374 -256
rect 424 -283 453 -256
rect 265 -284 296 -283
rect 344 -284 375 -283
rect 423 -284 454 -283
rect 461 -284 503 -255
rect -212 -315 -206 -309
rect -147 -315 -141 -309
rect 244 -334 251 -284
rect 266 -285 267 -284
rect 294 -285 295 -284
rect 345 -285 346 -284
rect 373 -285 374 -284
rect 424 -285 425 -284
rect 452 -285 453 -284
rect 467 -292 474 -284
rect 266 -334 267 -333
rect 294 -334 295 -333
rect 345 -334 346 -333
rect 373 -334 374 -333
rect 424 -334 425 -333
rect 452 -334 453 -333
rect 467 -334 474 -309
rect 216 -363 257 -334
rect 265 -335 296 -334
rect 344 -335 375 -334
rect 423 -335 454 -334
rect 266 -362 295 -335
rect 345 -362 374 -335
rect 424 -362 453 -335
rect 265 -363 296 -362
rect 344 -363 375 -362
rect 423 -363 454 -362
rect 461 -363 503 -334
rect 244 -378 251 -363
rect 266 -364 267 -363
rect 294 -364 295 -363
rect 345 -364 346 -363
rect 373 -364 374 -363
rect 424 -364 425 -363
rect 452 -364 453 -363
rect 266 -378 295 -372
rect 345 -378 374 -372
rect 424 -378 453 -372
rect 467 -378 474 -363
rect 244 -385 474 -378
rect 266 -413 295 -385
rect 345 -413 374 -385
rect 424 -413 453 -385
<< nwell >>
rect 632 -72 667 -71
rect 632 -88 649 -72
rect 666 -88 667 -72
<< poly >>
rect 453 147 489 151
rect -107 114 130 138
rect 453 135 488 147
rect -107 5 128 29
rect 453 -9 488 8
rect 649 -72 667 -71
rect 665 -88 667 -72
rect -107 -175 130 -151
rect 320 -167 488 -150
rect -105 -295 132 -271
rect 320 -309 488 -292
<< polycont >>
rect 632 -88 649 -71
<< locali >>
rect 623 -88 632 -71
<< viali >>
rect 649 -88 667 -71
<< metal1 >>
rect -228 -382 -188 217
rect 654 -68 667 -66
rect 646 -71 670 -68
rect 646 -88 649 -71
rect 667 -88 670 -71
rect 646 -91 670 -88
rect 656 -95 667 -91
<< metal2 >>
rect -264 166 497 173
rect -264 155 500 166
rect -264 112 710 130
rect -264 24 497 30
rect -264 12 500 24
rect -264 -20 496 -13
rect -264 -31 500 -20
rect -262 -146 500 -129
rect -262 -188 500 -171
rect -262 -286 500 -269
rect -184 -295 -30 -286
rect -262 -330 500 -313
use TunCap01  TunCap01_0
timestamp 1606740587
transform 1 0 1188 0 1 135
box -1451 -400 -1278 -210
use TunCap01  TunCap01_1
timestamp 1606740587
transform 1 0 1188 0 1 18
box -1451 -400 -1278 -210
use overlapCap01  overlapCap01_2
timestamp 1607257541
transform 1 0 503 0 1 -188
box -287 -71 0 137
use overlapCap01  overlapCap01_3
timestamp 1607257541
transform 1 0 503 0 1 -342
box -287 -71 0 137
use horizPcell01  horizPcell01_1
timestamp 1606750506
transform 1 0 777 0 1 -428
box -289 47 -33 232
use horizPcell01  horizPcell01_2
timestamp 1606750506
transform 1 0 777 0 -1 -31
box -289 47 -33 232
use TunCap01  TunCap01_2
timestamp 1606740587
transform 1 0 1188 0 1 324
box -1451 -400 -1278 -210
use wellContact  wellContact_1
timestamp 1606753443
transform 1 0 1185 0 1 293
box -1449 -441 -1275 -255
use TunCap01  TunCap01_3
timestamp 1606740587
transform 1 0 1188 0 1 433
box -1451 -400 -1278 -210
use overlapCap01  overlapCap01_1
timestamp 1607257541
transform 1 0 504 0 1 -32
box -287 -71 0 137
use horizPcell01  horizPcell01_0
timestamp 1606750506
transform 1 0 777 0 1 -128
box -289 47 -33 232
use overlapCap01  overlapCap01_0
timestamp 1607257541
transform 1 0 504 0 1 121
box -287 -71 0 137
use horizPcell01  horizPcell01_3
timestamp 1606750506
transform 1 0 777 0 -1 270
box -289 47 -33 232
<< end >>
