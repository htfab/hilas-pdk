magic
tech sky130A
timestamp 1629420194
<< error_p >>
rect -12 68 17 86
rect -12 36 -11 37
rect 16 36 17 37
rect -62 7 -44 36
rect -13 35 18 36
rect -12 26 17 35
rect -12 17 -2 26
rect 7 17 17 26
rect -12 8 17 17
rect -13 7 18 8
rect 49 7 67 36
rect -12 6 -11 7
rect 16 6 17 7
rect -12 -43 17 -25
<< mvnmos >>
rect -44 36 49 68
rect -44 7 -12 36
rect 17 7 49 36
rect -44 -25 49 7
<< mvndiff >>
rect -12 30 17 36
rect -12 13 -6 30
rect 11 13 17 30
rect -12 7 17 13
<< mvndiffc >>
rect -6 13 11 30
<< poly >>
rect -57 68 62 81
rect -57 -25 -44 68
rect 49 -25 62 68
rect -57 -38 62 -25
<< locali >>
rect -6 64 11 67
rect -6 30 11 47
rect -6 -5 11 13
<< viali >>
rect -6 47 11 64
rect -6 -22 11 -5
<< metal1 >>
rect -9 64 14 86
rect -9 47 -6 64
rect 11 47 14 64
rect -9 -5 14 47
rect -9 -22 -6 -5
rect 11 -22 14 -5
rect -9 -43 14 -22
<< end >>
