magic
tech sky130A
timestamp 1626460134
<< error_s >>
rect -626 12757 -597 12773
rect -547 12757 -518 12773
rect -468 12757 -439 12773
rect -389 12757 -360 12773
rect -1764 12733 -1757 12739
rect -913 12733 -907 12739
rect -81 12733 -75 12739
rect 24 12733 30 12739
rect 439 12728 445 12734
rect 494 12728 500 12734
rect -626 12723 -625 12724
rect -598 12723 -597 12724
rect -547 12723 -546 12724
rect -519 12723 -518 12724
rect -468 12723 -467 12724
rect -440 12723 -439 12724
rect -389 12723 -388 12724
rect -361 12723 -360 12724
rect -676 12694 -659 12723
rect -627 12722 -596 12723
rect -548 12722 -517 12723
rect -469 12722 -438 12723
rect -390 12722 -359 12723
rect -626 12715 -597 12722
rect -547 12715 -518 12722
rect -468 12715 -439 12722
rect -389 12715 -360 12722
rect -626 12701 -617 12715
rect -370 12701 -360 12715
rect -626 12695 -597 12701
rect -547 12695 -518 12701
rect -468 12695 -439 12701
rect -389 12695 -360 12701
rect -627 12694 -596 12695
rect -548 12694 -517 12695
rect -469 12694 -438 12695
rect -390 12694 -359 12695
rect -328 12694 -310 12723
rect -626 12693 -625 12694
rect -598 12693 -597 12694
rect -547 12693 -546 12694
rect -519 12693 -518 12694
rect -468 12693 -467 12694
rect -440 12693 -439 12694
rect -389 12693 -388 12694
rect -361 12693 -360 12694
rect -87 12683 -81 12689
rect 30 12683 36 12689
rect 433 12678 439 12684
rect 500 12678 506 12684
rect -626 12644 -597 12659
rect -547 12644 -518 12659
rect -468 12644 -439 12659
rect -389 12644 -360 12659
rect -626 12477 -597 12493
rect -547 12477 -518 12493
rect -468 12477 -439 12493
rect -389 12477 -360 12493
rect -2072 12474 -2067 12475
rect -626 12443 -625 12444
rect -598 12443 -597 12444
rect -547 12443 -546 12444
rect -519 12443 -518 12444
rect -468 12443 -467 12444
rect -440 12443 -439 12444
rect -389 12443 -388 12444
rect -361 12443 -360 12444
rect -676 12414 -659 12443
rect -627 12442 -596 12443
rect -548 12442 -517 12443
rect -469 12442 -438 12443
rect -390 12442 -359 12443
rect -626 12435 -597 12442
rect -547 12435 -518 12442
rect -468 12435 -439 12442
rect -389 12435 -360 12442
rect -626 12421 -617 12435
rect -370 12421 -360 12435
rect -626 12415 -597 12421
rect -547 12415 -518 12421
rect -468 12415 -439 12421
rect -389 12415 -360 12421
rect -627 12414 -596 12415
rect -548 12414 -517 12415
rect -469 12414 -438 12415
rect -390 12414 -359 12415
rect -328 12414 -310 12443
rect -81 12434 -75 12440
rect 24 12434 30 12440
rect -626 12413 -625 12414
rect -598 12413 -597 12414
rect -547 12413 -546 12414
rect -519 12413 -518 12414
rect -468 12413 -467 12414
rect -440 12413 -439 12414
rect -389 12413 -388 12414
rect -361 12413 -360 12414
rect 470 12395 499 12413
rect -87 12384 -81 12390
rect 30 12384 36 12390
rect -626 12364 -597 12379
rect -547 12364 -518 12379
rect -468 12364 -439 12379
rect -389 12364 -360 12379
rect 470 12363 471 12364
rect 498 12363 499 12364
rect -2360 12307 -2359 12362
rect -626 12322 -597 12338
rect -547 12322 -518 12338
rect -468 12322 -439 12338
rect -389 12322 -360 12338
rect -81 12333 -75 12339
rect 24 12333 30 12339
rect 420 12334 438 12363
rect 469 12362 500 12363
rect 470 12353 499 12362
rect 470 12344 480 12353
rect 489 12344 499 12353
rect 470 12335 499 12344
rect 469 12334 500 12335
rect 531 12334 549 12363
rect 470 12333 471 12334
rect 498 12333 499 12334
rect -626 12288 -625 12289
rect -598 12288 -597 12289
rect -547 12288 -546 12289
rect -519 12288 -518 12289
rect -468 12288 -467 12289
rect -440 12288 -439 12289
rect -389 12288 -388 12289
rect -361 12288 -360 12289
rect -1769 12267 -1763 12273
rect -907 12267 -901 12273
rect -676 12259 -659 12288
rect -627 12287 -596 12288
rect -548 12287 -517 12288
rect -469 12287 -438 12288
rect -390 12287 -359 12288
rect -626 12280 -597 12287
rect -547 12280 -518 12287
rect -468 12280 -439 12287
rect -389 12280 -360 12287
rect -626 12266 -617 12280
rect -370 12266 -360 12280
rect -626 12260 -597 12266
rect -547 12260 -518 12266
rect -468 12260 -439 12266
rect -389 12260 -360 12266
rect -627 12259 -596 12260
rect -548 12259 -517 12260
rect -469 12259 -438 12260
rect -390 12259 -359 12260
rect -328 12259 -310 12288
rect -87 12283 -81 12289
rect 30 12283 36 12289
rect 470 12284 499 12302
rect -626 12258 -625 12259
rect -598 12258 -597 12259
rect -547 12258 -546 12259
rect -519 12258 -518 12259
rect -468 12258 -467 12259
rect -440 12258 -439 12259
rect -389 12258 -388 12259
rect -361 12258 -360 12259
rect -626 12209 -597 12224
rect -547 12209 -518 12224
rect -468 12209 -439 12224
rect -389 12209 -360 12224
rect 3665 11232 3671 11238
rect 3718 11232 3724 11238
rect 3831 11232 3837 11238
rect 3884 11232 3890 11238
rect 3659 11182 3665 11188
rect 3724 11182 3730 11188
rect 3825 11182 3831 11188
rect 3890 11182 3896 11188
rect 3237 11173 3243 11179
rect 3342 11173 3348 11179
rect 4254 11173 4260 11179
rect 4359 11173 4365 11179
rect 3231 11123 3237 11129
rect 3348 11123 3354 11129
rect 4248 11123 4254 11129
rect 4365 11123 4371 11129
rect 1098 10993 1461 10994
rect 1518 10993 1641 10994
rect 1716 10987 1746 11106
rect 3237 10872 3243 10878
rect 3342 10872 3348 10878
rect 4254 10872 4260 10878
rect 4359 10872 4365 10878
rect 3231 10822 3237 10828
rect 3348 10822 3354 10828
rect 3665 10818 3671 10824
rect 3718 10818 3724 10824
rect 3831 10818 3837 10824
rect 3884 10818 3890 10824
rect 4248 10822 4254 10828
rect 4365 10822 4371 10828
rect 3659 10768 3665 10774
rect 3724 10768 3730 10774
rect 3825 10768 3831 10774
rect 3890 10768 3896 10774
rect 3499 10705 3503 10716
rect 3499 10691 3500 10702
rect 3608 10701 3609 10754
rect 3666 10629 3672 10635
rect 3719 10629 3725 10635
rect 3831 10629 3837 10635
rect 3884 10629 3890 10635
rect 3660 10579 3666 10585
rect 3725 10579 3731 10585
rect 3825 10579 3831 10585
rect 3890 10579 3896 10585
rect 3191 10570 3197 10576
rect 3296 10570 3302 10576
rect 4254 10570 4260 10576
rect 4359 10570 4365 10576
rect 3185 10520 3191 10526
rect 3302 10520 3308 10526
rect 4248 10520 4254 10526
rect 4365 10520 4371 10526
rect 4059 10385 4076 10386
rect 4059 10368 4076 10369
rect 3497 10351 3498 10364
rect 3191 10269 3197 10275
rect 3296 10269 3302 10275
rect 4254 10269 4260 10275
rect 4359 10269 4365 10275
rect 3185 10219 3191 10225
rect 3302 10219 3308 10225
rect 3666 10215 3672 10221
rect 3719 10215 3725 10221
rect 3831 10215 3837 10221
rect 3884 10215 3890 10221
rect 4248 10219 4254 10225
rect 4365 10219 4371 10225
rect 3660 10165 3666 10171
rect 3725 10165 3731 10171
rect 3825 10165 3831 10171
rect 3890 10165 3896 10171
rect 3239 9904 3245 9910
rect 3344 9904 3350 9910
rect 4210 9904 4216 9910
rect 4315 9904 4321 9910
rect 3665 9894 3671 9900
rect 3718 9894 3724 9900
rect 3836 9894 3842 9900
rect 3889 9894 3895 9900
rect 3233 9840 3239 9846
rect 3350 9840 3356 9846
rect 3659 9844 3665 9850
rect 3724 9844 3730 9850
rect 3830 9844 3836 9850
rect 3895 9844 3901 9850
rect 4204 9840 4210 9846
rect 4321 9840 4327 9846
rect 3239 9787 3245 9793
rect 3344 9787 3350 9793
rect 3665 9785 3671 9791
rect 3718 9785 3724 9791
rect 3836 9785 3842 9791
rect 3889 9785 3895 9791
rect 4210 9787 4216 9793
rect 4315 9787 4321 9793
rect 3659 9735 3665 9741
rect 3724 9735 3730 9741
rect 3830 9735 3836 9741
rect 3895 9735 3901 9741
rect 3233 9723 3239 9729
rect 3350 9723 3356 9729
rect 4204 9723 4210 9729
rect 4321 9723 4327 9729
rect 3239 9602 3245 9608
rect 3344 9602 3350 9608
rect 4210 9602 4216 9608
rect 4315 9602 4321 9608
rect 3665 9596 3671 9602
rect 3718 9596 3724 9602
rect 3836 9596 3842 9602
rect 3889 9596 3895 9602
rect 3659 9546 3665 9552
rect 3724 9546 3730 9552
rect 3830 9546 3836 9552
rect 3895 9546 3901 9552
rect 3233 9538 3239 9544
rect 3350 9538 3356 9544
rect 4204 9538 4210 9544
rect 4321 9538 4327 9544
rect 3239 9486 3245 9492
rect 3344 9486 3350 9492
rect 4210 9486 4216 9492
rect 4315 9486 4321 9492
rect 3665 9479 3671 9485
rect 3718 9479 3724 9485
rect 3836 9479 3842 9485
rect 3889 9479 3895 9485
rect 3659 9429 3665 9435
rect 3724 9429 3730 9435
rect 3830 9429 3836 9435
rect 3895 9429 3901 9435
rect 3233 9422 3239 9428
rect 3350 9422 3356 9428
rect 4204 9422 4210 9428
rect 4321 9422 4327 9428
rect 3239 8926 3245 8932
rect 3344 8926 3350 8932
rect 3665 8916 3671 8922
rect 3718 8916 3724 8922
rect 3233 8862 3239 8868
rect 3350 8862 3356 8868
rect 3659 8866 3665 8872
rect 3724 8866 3730 8872
rect 3239 8809 3245 8815
rect 3344 8809 3350 8815
rect 3665 8807 3671 8813
rect 3718 8807 3724 8813
rect 3659 8757 3665 8763
rect 3724 8757 3730 8763
rect 3233 8745 3239 8751
rect 3350 8745 3356 8751
rect 3239 8624 3245 8630
rect 3344 8624 3350 8630
rect 3502 8619 3519 8623
rect 3665 8618 3671 8624
rect 3718 8618 3724 8624
rect 3659 8568 3665 8574
rect 3724 8568 3730 8574
rect 3233 8560 3239 8566
rect 3350 8560 3356 8566
rect 3239 8508 3245 8514
rect 3344 8508 3350 8514
rect 3665 8501 3671 8507
rect 3718 8501 3724 8507
rect 3659 8451 3665 8457
rect 3724 8451 3730 8457
rect 3233 8444 3239 8450
rect 3350 8444 3356 8450
rect 8801 7705 8802 7718
rect 8801 7704 8815 7705
rect -1497 7546 -1490 7584
rect -1483 7552 -1476 7598
rect -817 7316 -816 7351
rect -803 7302 -802 7365
rect -931 7162 -919 7165
rect -943 7141 -938 7153
rect -950 6801 -938 6809
rect -719 6801 -717 6809
rect 7811 6656 7812 6658
rect 744 5906 911 5919
rect 1337 5909 1339 5922
rect 741 5892 911 5905
rect 1337 5895 1340 5908
rect 1747 5907 1748 5920
rect 1747 5893 1749 5906
<< metal1 >>
rect -13106 14454 -12717 14571
rect -10247 14453 -9858 14570
rect -7388 14453 -6999 14570
rect -3198 14456 -2809 14573
rect 1014 14454 1403 14571
rect 3873 14454 4262 14571
rect 6733 14454 7122 14571
rect 9592 14454 9981 14571
rect 12451 14454 12840 14571
rect 15310 14453 15699 14570
rect 18169 14453 18558 14570
rect -12554 12222 -12231 13533
rect -9695 12563 -9372 13533
rect -6836 12992 -6513 13533
rect -5582 13312 -5565 13324
rect -6879 12961 -6496 12992
rect -6879 12736 -6836 12961
rect -6513 12736 -6496 12961
rect -6879 12718 -6496 12736
rect -5617 12656 -5565 13312
rect -5623 12645 -5558 12656
rect -5623 12608 -5617 12645
rect -5565 12608 -5558 12645
rect -5623 12605 -5558 12608
rect -9711 12512 -9361 12563
rect -9711 12287 -9695 12512
rect -9372 12287 -9361 12512
rect -9711 12274 -9361 12287
rect -12771 12183 -12231 12222
rect -12771 11860 -12737 12183
rect -12512 11860 -12231 12183
rect -14015 11852 -13676 11859
rect -14112 11843 -13676 11852
rect -14435 11520 -13890 11843
rect -13704 11520 -13676 11843
rect -12771 11842 -12477 11860
rect -5617 11837 -5565 12605
rect -5277 12214 -5236 13335
rect -2566 13135 -2450 13326
rect -2566 13022 170 13135
rect -2566 13002 189 13022
rect 37 12862 170 13002
rect 1566 12911 1889 13534
rect 2730 13326 2791 13340
rect 2728 13130 2846 13326
rect 2648 13039 2846 13130
rect 2648 13021 2829 13039
rect 3172 13023 3244 13409
rect 2648 12952 2721 13021
rect 4425 12911 4748 13533
rect 7284 12911 7607 13533
rect 8177 13272 8196 13273
rect 8890 13272 8962 13409
rect 8177 13237 8962 13272
rect 8177 13024 8196 13237
rect 10143 13218 10466 13533
rect 10067 13190 10466 13218
rect 10065 13170 10466 13190
rect 10047 13073 10482 13170
rect 10047 12867 10143 13073
rect 10466 12867 10482 13073
rect 10047 12800 10482 12867
rect 13002 12752 13325 13533
rect 12972 12708 13327 12752
rect 12972 12378 13002 12708
rect 13208 12378 13327 12708
rect 12972 12347 13327 12378
rect -5289 12211 -5236 12214
rect -5289 12170 -5283 12211
rect -5242 12170 -5236 12211
rect 15861 12189 16184 13533
rect -5289 12167 -5236 12170
rect -5637 11828 -5565 11837
rect -5637 11776 -5631 11828
rect -5579 11776 -5565 11828
rect -5637 11764 -5565 11776
rect -14112 11452 -13676 11520
rect -15468 10968 -15343 11357
rect -13098 8984 -12872 8988
rect -14435 8661 -13085 8984
rect -12877 8661 -12872 8984
rect -13098 8657 -12872 8661
rect -15467 8110 -15342 8499
rect -5617 8229 -5565 11764
rect -5277 11742 -5236 12167
rect 15841 12159 16200 12189
rect 15841 11953 15861 12159
rect 16184 11953 16200 12159
rect 15841 11936 16200 11953
rect 18720 11840 19043 13533
rect -5291 11732 -5229 11742
rect -5291 11691 -5278 11732
rect -5237 11691 -5229 11732
rect -5291 11683 -5229 11691
rect 18689 11717 19065 11840
rect -5625 8226 -5562 8229
rect -5625 8174 -5621 8226
rect -5569 8174 -5562 8226
rect -5625 8169 -5562 8174
rect -5277 8127 -5236 11683
rect 18689 11512 18720 11717
rect 19043 11512 19065 11717
rect 18689 11478 19065 11512
rect 20124 11771 20465 11803
rect 20124 11448 20154 11771
rect 20353 11448 20788 11771
rect 10956 11382 11398 11443
rect 20124 11399 20465 11448
rect 10956 11350 10980 11382
rect 11202 11350 11398 11382
rect 10956 8432 11398 11350
rect 21692 10898 21817 11287
rect 19283 8912 19515 8920
rect 19283 8589 19299 8912
rect 19508 8589 20787 8912
rect 19283 8583 19515 8589
rect 10953 8420 11400 8432
rect 10953 8311 10964 8420
rect 11392 8311 11400 8420
rect 10953 8300 11400 8311
rect -5282 8124 -5234 8127
rect -5282 8080 -5278 8124
rect -5237 8080 -5234 8124
rect -5282 8077 -5234 8080
rect -12707 6125 -12484 6133
rect -14434 5802 -12695 6125
rect -12487 5802 -12484 6125
rect -12707 5787 -12484 5802
rect -15468 5250 -15343 5639
rect -12256 3266 -12015 3276
rect -14435 2943 -12232 3266
rect -12024 2943 -12015 3266
rect -12256 2933 -12015 2943
rect -15466 2391 -15341 2780
rect -11800 407 -11573 414
rect -14434 84 -11791 407
rect -11583 84 -11573 407
rect -11800 74 -11573 84
rect -15467 -467 -15342 -78
rect -11364 -2452 -11139 -2446
rect -14435 -2775 -11357 -2452
rect -11149 -2775 -11139 -2452
rect -11364 -2783 -11139 -2775
rect -15468 -3327 -15343 -2938
rect -10932 -5311 -10707 -5300
rect -14435 -5634 -10692 -5311
rect -10932 -5645 -10707 -5634
rect -15467 -6185 -15342 -5796
rect 10956 -7830 11398 8300
rect 21691 8038 21816 8427
rect 18866 6053 19102 6066
rect 18866 5730 18874 6053
rect 19083 5730 20789 6053
rect 18866 5720 19102 5730
rect 21691 5178 21816 5567
rect 18465 3194 18693 3210
rect 18465 2871 18476 3194
rect 18685 2871 20787 3194
rect 18465 2860 18693 2871
rect 21692 2322 21817 2711
rect 18035 335 18277 347
rect 18035 12 18051 335
rect 18260 12 20787 335
rect 18035 -4 18277 12
rect 21690 -539 21815 -150
rect 17646 -2524 17873 -2513
rect 17646 -2847 17657 -2524
rect 17866 -2847 20788 -2524
rect 17646 -2860 17873 -2847
rect 21692 -3397 21817 -3008
rect 17206 -5383 17436 -5375
rect 17206 -5706 20788 -5383
rect 17206 -5716 17436 -5706
rect 21692 -6258 21817 -5869
rect 10864 -7841 11398 -7830
rect -10526 -8170 -10285 -8160
rect -14435 -8493 -10503 -8170
rect -10295 -8493 -10285 -8170
rect 10864 -8283 10882 -7841
rect 11324 -8204 11398 -7841
rect 11324 -8283 11340 -8204
rect 10864 -8300 11340 -8283
rect -10526 -8511 -10285 -8493
rect -15464 -9043 -15339 -8654
rect -10098 -11029 -9852 -11022
rect -14435 -11352 -9852 -11029
rect -10098 -11357 -9852 -11352
rect -15466 -11904 -15341 -11515
rect -9661 -13888 -9421 -13874
rect -14436 -14211 -9641 -13888
rect -9433 -14211 -9421 -13888
rect -9661 -14221 -9421 -14211
rect -15467 -14763 -15342 -14374
rect -9267 -16747 -9018 -16739
rect -14436 -17070 -9244 -16747
rect -9036 -17070 -9018 -16747
rect -9267 -17089 -9018 -17070
rect -15467 -17622 -15342 -17233
rect -8820 -19606 -8585 -19596
rect -14434 -19929 -8800 -19606
rect -8592 -19929 -8585 -19606
rect -8820 -19942 -8585 -19929
rect -15466 -20481 -15341 -20092
rect -8420 -22465 -8149 -22459
rect -14434 -22788 -8370 -22465
rect -8162 -22788 -8149 -22465
rect -8420 -22800 -8149 -22788
rect -15466 -23339 -15341 -22950
<< via1 >>
rect -6836 12736 -6513 12961
rect -5617 12608 -5565 12645
rect -9695 12287 -9372 12512
rect -12737 11860 -12512 12183
rect -13890 11520 -13704 11843
rect 10143 12867 10466 13073
rect 13002 12378 13208 12708
rect -5283 12170 -5242 12211
rect -5631 11776 -5579 11828
rect -13085 8661 -12877 8984
rect 15861 11953 16184 12159
rect -5278 11691 -5237 11732
rect -5621 8174 -5569 8226
rect 18720 11512 19043 11717
rect 20154 11448 20353 11771
rect 10980 11350 11202 11382
rect 19299 8589 19508 8912
rect 10964 8311 11392 8420
rect -5278 8080 -5237 8124
rect -12695 5802 -12487 6125
rect -12232 2943 -12024 3266
rect -11791 84 -11583 407
rect -11357 -2775 -11149 -2452
rect 18874 5730 19083 6053
rect 18476 2871 18685 3194
rect 18051 12 18260 335
rect 17657 -2847 17866 -2524
rect -10503 -8493 -10295 -8170
rect 10882 -8283 11324 -7841
rect -9641 -14211 -9433 -13888
rect -9244 -17070 -9036 -16747
rect -8800 -19929 -8592 -19606
rect -8370 -22788 -8162 -22465
<< metal2 >>
rect 21381 14165 21500 14166
rect -15126 14164 -13833 14165
rect -15139 14025 -13833 14164
rect 20201 14113 21500 14165
rect 20180 14037 21500 14113
rect -15139 13873 -14910 14025
rect -15094 13869 -14910 13873
rect -15050 13017 -14910 13869
rect 21284 13905 21500 14037
rect -14423 13388 -13848 13528
rect 20116 13395 20783 13535
rect -14423 12916 -14283 13388
rect 10028 13073 10508 13153
rect -6892 12987 -6483 13012
rect -6892 12961 -2695 12987
rect -6892 12736 -6836 12961
rect -6513 12762 -2695 12961
rect 10028 12944 10143 13073
rect 8858 12867 10143 12944
rect 10466 12944 10508 13073
rect 10466 12867 10513 12944
rect -6513 12736 -6483 12762
rect 8858 12738 10513 12867
rect 20642 12844 20782 13395
rect 21284 12982 21412 13905
rect 21336 12908 21412 12982
rect -6892 12702 -6483 12736
rect 12987 12708 13318 12737
rect -5622 12651 -5560 12653
rect -5622 12645 -2707 12651
rect -5622 12608 -5617 12645
rect -5565 12614 -2707 12645
rect -5565 12608 -5560 12614
rect -5622 12607 -5560 12608
rect -9704 12538 -9366 12549
rect -9745 12512 -2695 12538
rect 12987 12531 13002 12708
rect -9745 12313 -9695 12512
rect -9704 12287 -9695 12313
rect -9372 12313 -2695 12512
rect 8858 12378 13002 12531
rect 13208 12531 13318 12708
rect 13208 12378 13350 12531
rect 8858 12325 13350 12378
rect -9372 12287 -9366 12313
rect -9704 12281 -9366 12287
rect -5287 12211 -5239 12212
rect -12758 12183 -12494 12207
rect -12758 12089 -12737 12183
rect -12766 11864 -12737 12089
rect -12758 11860 -12737 11864
rect -12512 12089 -12494 12183
rect -5287 12170 -5283 12211
rect -5242 12209 -5239 12211
rect -5242 12171 -2708 12209
rect -5242 12170 -5239 12171
rect -5287 12169 -5239 12170
rect 15826 12159 16219 12168
rect 15826 12123 15861 12159
rect -12512 11864 -2735 12089
rect 8858 11953 15861 12123
rect 16184 11953 16219 12159
rect 8858 11917 16219 11953
rect 15826 11916 16219 11917
rect -12512 11860 -12494 11864
rect -13981 11843 -13692 11851
rect -12758 11847 -12494 11860
rect -13981 11655 -13890 11843
rect -13984 11520 -13890 11655
rect -13704 11655 -13692 11843
rect -5634 11828 -5572 11831
rect -5634 11776 -5631 11828
rect -5579 11822 -5572 11828
rect -5579 11781 -2740 11822
rect -5579 11776 -5572 11781
rect -5634 11772 -5572 11776
rect 19876 11771 20447 11846
rect -5287 11732 -5233 11735
rect -5287 11691 -5278 11732
rect -5237 11691 -2744 11732
rect 18706 11717 19056 11743
rect -5287 11687 -5233 11691
rect 18706 11689 18720 11717
rect -13704 11520 -2772 11655
rect -13984 11469 -2772 11520
rect 8858 11512 18720 11689
rect 19043 11689 19056 11717
rect 19043 11512 19065 11689
rect 8858 11484 19065 11512
rect 19876 11448 20154 11771
rect 20353 11448 20447 11771
rect 8876 11382 11209 11387
rect 8876 11350 10980 11382
rect 11202 11350 11209 11382
rect 8876 11344 11209 11350
rect 19876 11282 20447 11448
rect 19832 11278 20447 11282
rect 8858 11232 20447 11278
rect -13095 11003 -2743 11211
rect 8858 11042 20431 11232
rect -13095 8992 -12887 11003
rect 19298 10804 19507 10822
rect -12679 10515 -2695 10723
rect 8858 10595 19507 10804
rect -13102 8984 -12868 8992
rect -13102 8661 -13085 8984
rect -12877 8661 -12868 8984
rect -13102 8655 -12868 8661
rect -13095 8568 -12887 8655
rect -12679 6132 -12471 10515
rect -12701 6125 -12471 6132
rect -12701 5802 -12695 6125
rect -12487 5802 -12471 6125
rect -12701 5791 -12471 5802
rect -12679 5758 -12471 5791
rect -12245 10033 -2695 10241
rect 8858 10055 19093 10264
rect -12245 3284 -12037 10033
rect -11791 9563 -2695 9771
rect 8858 9567 18685 9776
rect -12266 3266 -12009 3284
rect -12266 2943 -12232 3266
rect -12024 2943 -12009 3266
rect -12266 2924 -12009 2943
rect -12245 2920 -12037 2924
rect -11791 422 -11583 9563
rect -11356 9137 -2695 9345
rect -11807 407 -11568 422
rect -11807 84 -11791 407
rect -11583 84 -11568 407
rect -11807 65 -11568 84
rect -11791 12 -11583 65
rect -11356 -2439 -11148 9137
rect 8858 9047 18276 9256
rect -10922 8730 -2695 8938
rect -11374 -2452 -11129 -2439
rect -11374 -2775 -11357 -2452
rect -11149 -2775 -11129 -2452
rect -11374 -2791 -11129 -2775
rect -11356 -2803 -11148 -2791
rect -10922 -5290 -10714 8730
rect 8858 8543 17863 8752
rect -10506 8315 -2695 8523
rect 10955 8421 11408 8429
rect 8886 8420 11415 8421
rect -10947 -5663 -10687 -5290
rect -10922 -5696 -10714 -5663
rect -10506 -8153 -10298 8315
rect 8886 8311 10964 8420
rect 11392 8311 11415 8420
rect 8886 8306 11415 8311
rect 10955 8304 11408 8306
rect -5624 8226 -5564 8227
rect -5624 8174 -5621 8226
rect -5569 8222 -5564 8226
rect -5569 8178 -2690 8222
rect -5569 8174 -5564 8178
rect -5624 8171 -5564 8174
rect -5281 8124 -5235 8125
rect -5281 8080 -5278 8124
rect -5237 8080 -2694 8124
rect -5281 8078 -5235 8080
rect -10081 7800 -2695 8008
rect 8890 7992 17439 8201
rect -10548 -8170 -10277 -8153
rect -10548 -8493 -10503 -8170
rect -10295 -8493 -10277 -8170
rect -10548 -8520 -10277 -8493
rect -10506 -8592 -10298 -8520
rect -10081 -11015 -9873 7800
rect -9655 7374 -2695 7582
rect -10114 -11363 -9840 -11015
rect -10081 -11444 -9873 -11363
rect -9655 -13844 -9447 7374
rect -9240 6870 -2695 7078
rect -9677 -13888 -9398 -13844
rect -9677 -14211 -9641 -13888
rect -9433 -14211 -9398 -13888
rect -9677 -14249 -9398 -14211
rect -9655 -14277 -9447 -14249
rect -9240 -16722 -9032 6870
rect -8805 6309 -2695 6517
rect -9289 -16747 -9006 -16722
rect -9289 -17070 -9244 -16747
rect -9036 -17070 -9006 -16747
rect -9289 -17100 -9006 -17070
rect -9240 -17156 -9032 -17100
rect -8805 -19580 -8597 6309
rect -8389 5839 -2695 6047
rect -8840 -19606 -8575 -19580
rect -8840 -19929 -8800 -19606
rect -8592 -19929 -8575 -19606
rect -8840 -19952 -8575 -19929
rect -8805 -19953 -8597 -19952
rect -8389 -22450 -8181 5839
rect -8408 -22465 -8141 -22450
rect -8408 -22788 -8370 -22465
rect -8162 -22788 -8141 -22465
rect -8408 -22803 -8141 -22788
rect -2235 -23386 -1901 5853
rect -1269 -23816 -1067 5843
rect -863 -23659 -661 5843
rect -863 -23815 -660 -23659
rect -466 -23660 -264 5843
rect -66 -23660 136 5843
rect -863 -23816 -661 -23815
rect -467 -23816 -264 -23660
rect -67 -23816 136 -23660
rect 339 -23816 541 5843
rect 740 -23659 942 5843
rect 739 -23815 942 -23659
rect 740 -23816 942 -23815
rect 1140 -23816 1342 5843
rect 1549 -23816 1751 5843
rect 1962 -23660 2164 5843
rect 2362 -23660 2564 5843
rect 2758 -23660 2960 5843
rect 1961 -23816 2164 -23660
rect 2361 -23816 2564 -23660
rect 2757 -23816 2960 -23660
rect 3163 -23659 3365 5843
rect 3163 -23815 3366 -23659
rect 3163 -23816 3365 -23815
rect 3572 -23816 3774 5843
rect 3973 -23661 4175 5843
rect 4377 -23660 4579 5843
rect 3973 -23816 4176 -23661
rect 4377 -23816 4580 -23660
rect 4786 -23662 4988 5843
rect 4786 -23816 4989 -23662
rect 5191 -23816 5393 5843
rect 5588 -23816 5790 5843
rect 6000 -23816 6202 5843
rect 3974 -23817 4176 -23816
rect 4787 -23818 4989 -23816
rect 6413 -23817 6615 5843
rect 6814 -23816 7016 5843
rect 7215 -23648 7417 5843
rect 7215 -23814 7419 -23648
rect 7624 -23650 7826 5843
rect 7624 -23816 7827 -23650
rect 8041 -23816 8243 5843
rect 8441 -23650 8643 5843
rect 8842 -23650 9044 5843
rect 9238 -23650 9440 5843
rect 8441 -23816 8644 -23650
rect 8839 -23816 9044 -23650
rect 9237 -23816 9440 -23650
rect 9643 -23650 9845 5843
rect 10049 -23650 10251 5843
rect 17230 -5151 17439 7992
rect 17654 -2504 17863 8543
rect 18067 344 18276 9047
rect 18476 3221 18685 9567
rect 18884 6071 19093 10055
rect 19298 8927 19507 10595
rect 19278 8912 19521 8927
rect 19278 8589 19299 8912
rect 19508 8589 19521 8912
rect 19278 8573 19521 8589
rect 19298 8506 19507 8573
rect 18860 6053 19111 6071
rect 18860 5730 18874 6053
rect 19083 5730 19111 6053
rect 18860 5714 19111 5730
rect 18456 3194 18708 3221
rect 18456 2871 18476 3194
rect 18685 2871 18708 3194
rect 18456 2850 18708 2871
rect 18476 2847 18685 2850
rect 18040 335 18276 344
rect 18040 12 18051 335
rect 18260 12 18276 335
rect 18040 2 18276 12
rect 18067 -69 18276 2
rect 17637 -2524 17880 -2504
rect 17637 -2847 17657 -2524
rect 17866 -2847 17880 -2524
rect 17637 -2875 17880 -2847
rect 17231 -5341 17439 -5151
rect 17231 -5353 17440 -5341
rect 17220 -5359 17440 -5353
rect 17194 -5727 17447 -5359
rect 17220 -5729 17429 -5727
rect 21338 -6998 21412 -6964
rect 20640 -7101 20780 -7023
rect 21272 -7038 21413 -6998
rect 20639 -7113 20780 -7101
rect 21274 -7107 21412 -7038
rect 20638 -7128 20780 -7113
rect 20638 -7218 20779 -7128
rect 21273 -7224 21413 -7107
rect 10871 -7841 11331 -7836
rect 10871 -8283 10882 -7841
rect 11324 -7914 11331 -7841
rect 11324 -8082 20786 -7914
rect 11324 -8211 20799 -8082
rect 11324 -8283 11331 -8211
rect 10871 -8293 11331 -8283
rect 9643 -23816 9847 -23650
rect 10049 -23816 10253 -23650
rect -15053 -24304 -14913 -24107
rect -14423 -24337 -14283 -23971
use sky130_hilas_TopLevelTextStructure  sky130_hilas_TopLevelTextStructure_0
timestamp 1626460134
transform 1 0 -2990 0 1 6624
box 218 -793 13243 6785
use sky130_hilas_RightProtection  sky130_hilas_RightProtection_0
timestamp 1626060794
transform 1 0 22518 0 1 -15744
box -2054 8715 -826 28728
use sky130_hilas_LeftProtection  sky130_hilas_LeftProtection_0
timestamp 1626060794
transform 1 0 -13278 0 1 -15672
box -2065 -8439 -833 28728
use sky130_hilas_TopProtection  sky130_hilas_TopProtection_0
timestamp 1626100607
transform 1 0 -13875 0 1 13286
box -2 -76 34131 1170
<< labels >>
rlabel metal1 21692 -6258 21817 -5869 0 IO07
port 1 nsew
rlabel metal1 21692 -3397 21817 -3008 0 IO08
port 2 nsew
rlabel metal1 21690 -539 21815 -150 0 IO09
port 3 nsew
rlabel metal1 21692 2322 21817 2711 0 IO10
port 4 nsew
rlabel metal1 21691 5178 21816 5567 0 IO11
port 5 nsew
rlabel metal1 21691 8038 21816 8427 0 IO12
port 6 nsew
rlabel metal1 21692 10898 21817 11287 0 IO13
port 7 nsew
rlabel metal1 -15468 10968 -15343 11357 0 IO25
port 8 nsew
rlabel metal1 -15467 8110 -15342 8499 0 IO26
port 9 nsew
rlabel metal1 -15468 5250 -15343 5639 0 IO27
port 10 nsew
rlabel metal1 -15466 2391 -15341 2780 0 IO28
port 11 nsew
rlabel metal1 -15467 -467 -15342 -78 0 IO29
port 12 nsew
rlabel metal1 -15468 -3327 -15343 -2938 0 IO30
port 13 nsew
rlabel metal1 -15467 -6185 -15342 -5796 0 IO31
port 14 nsew
rlabel metal1 -15464 -9043 -15339 -8654 0 IO32
port 15 nsew
rlabel metal1 -15466 -11904 -15341 -11515 0 IO33
port 16 nsew
rlabel metal1 -15467 -14763 -15342 -14374 0 IO34
port 17 nsew
rlabel metal1 -15467 -17622 -15342 -17233 0 IO35
port 18 nsew
rlabel metal1 -15466 -20481 -15341 -20092 0 IO36
port 19 nsew
rlabel metal1 -15466 -23339 -15341 -22950 0 IO37
port 20 nsew
rlabel metal2 -15139 13873 -14971 14164 0 Vssa1
port 21 nsew
rlabel metal1 -13106 14454 -12717 14571 0 ANALOG10
port 22 nsew
rlabel metal1 -10247 14453 -9858 14570 0 ANALOG09
port 23 nsew
rlabel metal1 -7388 14453 -6999 14570 0 ANALOG08
port 24 nsew
rlabel metal1 -3198 14456 -2809 14573 0 ANALOG07
port 25 nsew
rlabel metal1 1014 14454 1403 14571 0 ANALOG06
port 26 nsew
rlabel metal1 3873 14454 4262 14571 0 ANALOG05
port 27 nsew
rlabel metal1 6733 14454 7122 14571 0 ANALOG04
port 28 nsew
rlabel metal1 9592 14454 9981 14571 0 ANALOG03
port 29 nsew
rlabel metal1 12451 14454 12840 14571 0 ANALOG02
port 30 nsew
rlabel metal1 15310 14453 15699 14570 0 ANALOG01
port 31 nsew
rlabel metal1 18169 14453 18558 14570 0 ANALOG00
port 32 nsew
rlabel metal2 21381 13908 21500 14166 0 VSSA1
port 33 nsew
rlabel metal2 -14423 -24337 -14283 -24197 0 VDDA1
port 34 nsew
rlabel metal2 -15053 -24304 -14913 -24164 0 VSSA1
port 33 nsew
rlabel metal2 20639 -7218 20779 -7101 0 VDDA1
port 34 nsew
rlabel metal2 21273 -7224 21413 -7107 0 VSSA1
port 33 nsew
rlabel metal2 -1269 -23816 -1067 -23660 0 LADATAOUT00
port 36 nsew
rlabel metal2 -862 -23815 -660 -23659 0 LADATAOUT01
port 35 nsew
rlabel metal2 -467 -23816 -265 -23660 0 LADATAOUT02
port 37 nsew
rlabel metal2 -67 -23816 135 -23660 0 LADATAOUT03
port 38 nsew
rlabel metal2 339 -23816 541 -23660 0 LADATAOUT04
port 39 nsew
rlabel metal2 739 -23815 941 -23659 0 LADATAOUT05
port 40 nsew
rlabel metal2 1140 -23816 1342 -23660 0 LADATAOUT06
port 41 nsew
rlabel metal2 1549 -23816 1751 -23660 0 LADATAOUT07
port 42 nsew
rlabel metal2 1961 -23816 2163 -23660 0 LADATAOUT08
port 43 nsew
rlabel metal2 2361 -23816 2563 -23660 0 LADATAOUT09
port 44 nsew
rlabel metal2 2757 -23816 2959 -23660 0 LADATAOUT10
port 45 nsew
rlabel metal2 3164 -23815 3366 -23659 0 LADATAOUT11
port 46 nsew
rlabel metal2 3572 -23816 3774 -23660 0 LADATAOUT12
port 47 nsew
rlabel metal2 3974 -23817 4176 -23661 0 LADATAOUT13
port 48 nsew
rlabel metal2 4378 -23816 4580 -23660 0 LADATAOUT14
port 49 nsew
rlabel metal2 4787 -23818 4989 -23662 0 LADATAOUT15
port 50 nsew
rlabel metal2 5191 -23816 5393 -23660 0 LADATA16
port 51 nsew
rlabel metal2 5588 -23816 5790 -23660 0 LADATAOUT17
port 52 nsew
rlabel metal2 6000 -23815 6202 -23659 0 LADATAOUT18
port 53 nsew
rlabel metal2 6413 -23817 6615 -23661 0 LADATAOUT19
port 54 nsew
rlabel metal2 6814 -23816 7016 -23660 0 LADATAOUT20
port 55 nsew
rlabel metal2 7215 -23814 7419 -23648 0 LADATAOUT21
port 56 nsew
rlabel metal2 7624 -23816 7827 -23650 0 LADATAOUT22
port 57 nsew
rlabel space 8039 -23816 8242 -23650 0 LADATAOUT23
port 58 nsew
rlabel metal2 8441 -23816 8644 -23650 0 LADATAOUT24
port 59 nsew
rlabel metal2 8839 -23816 9042 -23650 0 LADATAIN00
port 60 nsew
rlabel metal2 9237 -23816 9440 -23650 0 LADATAIN01
port 61 nsew
rlabel metal2 9644 -23816 9847 -23650 0 LADATAIN02
port 62 nsew
rlabel metal2 10050 -23816 10253 -23650 0 LADATAIN03
port 63 nsew
rlabel metal2 20683 -8211 20799 -8085 0 VCCA
port 64 nsew
<< end >>
