VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_TA2Cell_1FG_Strong
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TA2Cell_1FG_Strong ;
  ORIGIN 26.170 -1.400 ;
  SIZE 28.100 BY 6.050 ;
  PIN Vin+_Amp2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -2.520 4.510 -2.170 4.750 ;
    END
  END Vin+_Amp2
  PIN Vin-_Amp2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -2.600 7.180 -1.940 7.420 ;
    END
  END Vin-_Amp2
  PIN Vdd
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.630 7.300 0.910 7.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.640 1.400 0.910 3.050 ;
    END
  END Vdd
  PIN GateColSelect
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT -4.160 5.920 -3.970 7.450 ;
    END
    PORT
      LAYER met1 ;
        RECT -4.160 1.400 -3.970 2.930 ;
    END
  END GateColSelect
  PIN Vin+_Amp1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT -23.530 7.020 -23.320 7.450 ;
    END
  END Vin+_Amp1
  PIN GND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT -0.030 6.750 0.310 7.450 ;
    END
    PORT
      LAYER met1 ;
        RECT -0.030 1.400 0.310 2.140 ;
    END
  END GND
  PIN output2
    PORT
      LAYER met2 ;
        RECT 1.750 3.920 1.930 4.150 ;
    END
  END output2
  PIN output1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.600 4.740 1.930 4.970 ;
    END
  END output1
  PIN Vinj
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT -3.720 6.740 -3.440 7.450 ;
    END
    PORT
      LAYER met1 ;
        RECT -3.720 1.400 -3.440 2.110 ;
    END
  END Vinj
  OBS
      LAYER nwell ;
        RECT -26.170 1.410 -22.860 7.440 ;
      LAYER li1 ;
        RECT -25.780 1.650 1.790 7.450 ;
      LAYER met1 ;
        RECT -25.820 6.740 -23.810 7.450 ;
        RECT -23.040 6.740 -4.440 7.450 ;
        RECT -25.820 5.640 -4.440 6.740 ;
        RECT -3.160 6.470 -0.310 7.450 ;
        RECT 1.190 7.020 1.630 7.450 ;
        RECT 0.590 6.470 1.630 7.020 ;
        RECT -3.160 6.460 1.630 6.470 ;
        RECT -3.690 5.640 1.630 6.460 ;
        RECT -25.820 3.330 1.630 5.640 ;
        RECT -25.820 3.210 0.360 3.330 ;
        RECT -25.820 1.400 -4.440 3.210 ;
        RECT -3.690 2.420 0.360 3.210 ;
        RECT -3.690 2.390 -0.310 2.420 ;
        RECT -3.160 1.400 -0.310 2.390 ;
        RECT 1.190 1.400 1.630 3.330 ;
      LAYER met2 ;
        RECT -26.170 6.900 -2.880 7.440 ;
        RECT -1.660 6.900 1.750 7.440 ;
        RECT -26.170 5.250 1.750 6.900 ;
        RECT -26.170 5.030 1.320 5.250 ;
        RECT -26.170 4.230 -2.800 5.030 ;
        RECT -1.890 4.460 1.320 5.030 ;
        RECT -1.890 4.430 1.750 4.460 ;
        RECT -1.890 4.230 1.470 4.430 ;
        RECT -26.170 3.640 1.470 4.230 ;
        RECT -26.170 1.690 1.750 3.640 ;
  END
END sky130_hilas_TA2Cell_1FG_Strong
END LIBRARY

