magic
tech sky130A
timestamp 1637951121
<< error_p >>
rect -239 308 -65 310
rect -178 277 -126 283
rect -206 275 -98 277
rect 176 276 226 281
rect -178 235 -126 241
rect 176 234 226 239
rect -252 210 -199 215
rect -105 210 -53 215
rect 105 209 155 215
rect 247 209 297 215
rect -279 173 -171 177
rect -132 173 -26 177
rect -252 168 -199 173
rect -105 168 -53 173
rect 105 167 155 173
rect 247 167 297 173
rect -312 140 7 144
<< nwell >>
rect -336 144 8 308
<< mvnmos >>
rect 176 239 226 276
rect 105 173 155 209
rect 247 173 297 209
<< mvpmos >>
rect -178 241 -126 277
rect -252 173 -199 210
rect -105 173 -53 210
<< mvndiff >>
rect 145 263 176 276
rect 145 246 152 263
rect 169 246 176 263
rect 145 239 176 246
rect 226 263 253 276
rect 226 246 232 263
rect 249 246 253 263
rect 226 239 253 246
rect 76 202 105 209
rect 76 185 81 202
rect 98 185 105 202
rect 76 173 105 185
rect 155 202 183 209
rect 155 185 161 202
rect 178 185 183 202
rect 155 173 183 185
rect 219 202 247 209
rect 219 185 224 202
rect 241 185 247 202
rect 219 173 247 185
rect 297 202 326 209
rect 297 185 303 202
rect 320 185 326 202
rect 297 173 326 185
<< mvpdiff >>
rect -206 267 -178 277
rect -206 250 -201 267
rect -184 250 -178 267
rect -206 241 -178 250
rect -126 267 -98 277
rect -126 250 -120 267
rect -103 250 -98 267
rect -126 241 -98 250
rect -279 202 -252 210
rect -279 185 -275 202
rect -258 185 -252 202
rect -279 173 -252 185
rect -199 202 -171 210
rect -199 185 -193 202
rect -176 185 -171 202
rect -199 173 -171 185
rect -132 202 -105 210
rect -132 185 -128 202
rect -111 185 -105 202
rect -132 173 -105 185
rect -53 202 -26 210
rect -53 185 -47 202
rect -30 185 -26 202
rect -53 173 -26 185
<< mvndiffc >>
rect 152 246 169 263
rect 232 246 249 263
rect 81 185 98 202
rect 161 185 178 202
rect 224 185 241 202
rect 303 185 320 202
<< mvpdiffc >>
rect -201 250 -184 267
rect -120 250 -103 267
rect -275 185 -258 202
rect -193 185 -176 202
rect -128 185 -111 202
rect -47 185 -30 202
<< psubdiff >>
rect 292 264 333 271
rect 292 247 304 264
rect 321 247 333 264
rect 292 239 333 247
<< mvnsubdiff >>
rect -286 267 -245 275
rect -286 250 -274 267
rect -257 250 -245 267
rect -286 241 -245 250
<< psubdiffcont >>
rect 304 247 321 264
<< mvnsubdiffcont >>
rect -274 250 -257 267
<< poly >>
rect -141 295 195 299
rect -143 294 195 295
rect -143 290 -13 294
rect -178 284 -13 290
rect -178 277 -126 284
rect -19 283 -13 284
rect -18 277 -13 283
rect 4 289 195 294
rect 4 284 226 289
rect 4 277 9 284
rect -18 269 9 277
rect 176 276 226 284
rect -74 251 -39 257
rect -327 226 -236 233
rect -327 218 -199 226
rect -178 225 -126 241
rect -74 234 -64 251
rect -47 234 -39 251
rect -74 233 -39 234
rect -74 230 120 233
rect -74 225 123 230
rect 176 225 226 239
rect -327 197 -300 218
rect -252 210 -199 218
rect -105 223 123 225
rect -105 218 155 223
rect -105 210 -53 218
rect -327 180 -322 197
rect -305 180 -300 197
rect -327 172 -300 180
rect 105 209 155 218
rect 247 209 297 223
rect 334 178 367 200
rect -252 160 -199 173
rect -105 160 -53 173
rect 105 160 155 173
rect 247 165 297 173
rect 334 165 345 178
rect 247 161 345 165
rect 362 161 367 178
rect 247 155 367 161
rect 266 150 367 155
<< polycont >>
rect -13 277 4 294
rect -64 234 -47 251
rect -322 180 -305 197
rect 345 161 362 178
<< locali >>
rect -17 294 4 303
rect -17 292 -13 294
rect -274 267 -257 279
rect -17 275 -15 292
rect 2 275 4 277
rect -201 267 -184 275
rect -120 267 -103 275
rect -17 269 4 275
rect -274 248 -272 250
rect -184 250 -180 267
rect -274 238 -257 248
rect -201 210 -180 250
rect -124 250 -120 267
rect 81 268 108 269
rect -124 242 -103 250
rect -64 251 -47 259
rect -124 210 -107 242
rect 81 251 84 268
rect 101 263 108 268
rect 223 264 249 271
rect 303 264 321 265
rect 223 263 304 264
rect 101 251 152 263
rect 81 246 152 251
rect 169 246 177 263
rect 223 246 232 263
rect 249 247 304 263
rect 321 247 329 264
rect 249 246 321 247
rect 81 245 108 246
rect -50 232 -47 234
rect -64 222 -47 232
rect -326 197 -301 205
rect -326 195 -322 197
rect -326 178 -324 195
rect -305 180 -301 197
rect -307 178 -301 180
rect -326 172 -301 178
rect -275 204 -258 210
rect -275 202 -250 204
rect -258 197 -250 202
rect -275 180 -271 185
rect -254 180 -250 197
rect -201 202 -176 210
rect -201 185 -193 202
rect -275 177 -250 180
rect -274 175 -250 177
rect -193 176 -176 185
rect -128 202 -107 210
rect 90 202 107 245
rect 223 232 249 246
rect 223 214 226 232
rect 244 214 249 232
rect 343 223 368 225
rect 343 220 349 223
rect 223 202 249 214
rect -111 185 -107 202
rect -56 185 -47 202
rect -30 185 81 202
rect 98 185 107 202
rect 152 185 161 202
rect 178 185 224 202
rect 241 185 249 202
rect 303 206 349 220
rect 366 206 368 223
rect 303 203 368 206
rect 303 202 320 203
rect -128 177 -111 185
rect 303 177 320 185
rect 340 178 362 186
rect 340 176 345 178
rect 340 159 343 176
rect 360 159 362 161
rect 340 153 362 159
<< viali >>
rect -15 277 -13 292
rect -13 277 2 292
rect -15 275 2 277
rect -272 250 -257 265
rect -257 250 -255 265
rect -272 248 -255 250
rect -67 234 -64 249
rect -64 234 -50 249
rect 84 251 101 268
rect -67 232 -50 234
rect -324 180 -322 195
rect -322 180 -307 195
rect -324 178 -307 180
rect -271 185 -258 197
rect -258 185 -254 197
rect -271 180 -254 185
rect 226 214 244 232
rect 349 206 366 223
rect 343 161 345 176
rect 345 161 360 176
rect 343 159 360 161
<< metal1 >>
rect -275 270 -253 308
rect -22 298 10 299
rect -22 272 -19 298
rect 7 272 10 298
rect -275 265 -252 270
rect -22 269 10 272
rect 76 273 110 274
rect -275 248 -272 265
rect -255 248 -252 265
rect -275 244 -252 248
rect -275 204 -253 244
rect -73 228 -69 254
rect -43 228 -40 254
rect 76 247 80 273
rect 106 269 110 273
rect 106 247 117 269
rect 76 244 117 247
rect 76 243 110 244
rect 222 232 249 310
rect 222 214 226 232
rect 244 214 249 232
rect -331 201 -297 204
rect -331 175 -327 201
rect -301 175 -297 201
rect -331 172 -297 175
rect -275 197 -250 204
rect -275 180 -271 197
rect -254 180 -250 197
rect -275 173 -250 180
rect -275 148 -253 173
rect 222 148 249 214
rect 343 231 377 234
rect 343 205 348 231
rect 374 205 377 231
rect 343 202 377 205
rect 332 182 362 186
rect 332 156 333 182
rect 359 179 362 182
rect 359 176 363 179
rect 360 159 363 176
rect 359 156 363 159
rect 332 153 362 156
<< via1 >>
rect -19 292 7 298
rect -19 275 -15 292
rect -15 275 2 292
rect 2 275 7 292
rect -19 272 7 275
rect -69 249 -43 254
rect -69 232 -67 249
rect -67 232 -50 249
rect -50 232 -43 249
rect -69 228 -43 232
rect 80 268 106 273
rect 80 251 84 268
rect 84 251 101 268
rect 101 251 106 268
rect 80 247 106 251
rect -327 195 -301 201
rect -327 178 -324 195
rect -324 178 -307 195
rect -307 178 -301 195
rect -327 175 -301 178
rect 348 223 374 231
rect 348 206 349 223
rect 349 206 366 223
rect 366 206 374 223
rect 348 205 374 206
rect 333 176 359 182
rect 333 159 343 176
rect 343 159 359 176
rect 333 156 359 159
<< metal2 >>
rect -22 289 -19 298
rect -337 273 -19 289
rect -22 272 -19 273
rect 7 272 10 298
rect -22 269 10 272
rect -73 246 -69 254
rect -100 244 -69 246
rect -337 228 -69 244
rect -43 228 -40 254
rect 77 247 80 273
rect 106 266 109 273
rect 106 249 387 266
rect 106 247 109 249
rect 77 244 109 247
rect 373 232 387 249
rect 345 231 387 232
rect 345 205 348 231
rect 374 205 387 231
rect 345 203 387 205
rect -330 201 -298 203
rect -330 195 -327 201
rect -337 179 -327 195
rect -330 175 -327 179
rect -301 181 -298 201
rect 333 182 359 185
rect -301 175 333 181
rect -330 173 333 175
rect -329 165 333 173
rect 373 175 387 203
rect 333 153 359 156
<< labels >>
rlabel metal2 -337 273 -331 289 0 Input1
rlabel metal2 -337 228 -331 244 0 Input2
rlabel metal2 -337 179 -331 195 0 Input3
rlabel metal1 222 299 249 305 0 GND
rlabel metal1 222 153 249 158 0 GND
rlabel metal1 -275 153 -253 159 0 Vinj
rlabel metal1 -275 297 -253 304 0 Vinj
rlabel metal2 381 175 387 192 0 OUTPUT
port 1 nsew
<< end >>
