magic
tech sky130A
timestamp 1628704276
<< checkpaint >>
rect 822 1272 2255 1666
rect 122 1081 2255 1272
rect -629 -199 2255 1081
rect -629 -365 1638 -199
rect 122 -604 1638 -365
<< error_s >>
rect 531 643 560 671
rect 610 643 639 671
rect 689 643 718 671
rect 509 636 739 643
rect 509 621 516 636
rect 531 630 560 636
rect 610 630 639 636
rect 689 630 718 636
rect 531 621 532 622
rect 559 621 560 622
rect 610 621 611 622
rect 638 621 639 622
rect 689 621 690 622
rect 717 621 718 622
rect 732 621 739 636
rect 481 592 522 621
rect 530 620 561 621
rect 609 620 640 621
rect 688 620 719 621
rect 531 593 560 620
rect 610 593 639 620
rect 689 593 718 620
rect 530 592 561 593
rect 609 592 640 593
rect 688 592 719 593
rect 726 592 768 621
rect 58 563 64 569
rect 111 563 117 569
rect 509 542 516 592
rect 531 591 532 592
rect 559 591 560 592
rect 610 591 611 592
rect 638 591 639 592
rect 689 591 690 592
rect 717 591 718 592
rect 732 564 739 592
rect 531 542 532 543
rect 559 542 560 543
rect 610 542 611 543
rect 638 542 639 543
rect 689 542 690 543
rect 717 542 718 543
rect 732 542 739 548
rect 752 547 753 548
rect 52 513 58 519
rect 117 513 123 519
rect 481 513 522 542
rect 530 541 561 542
rect 609 541 640 542
rect 688 541 719 542
rect 531 514 560 541
rect 610 514 639 541
rect 689 514 718 541
rect 530 513 561 514
rect 609 513 640 514
rect 688 513 719 514
rect 726 513 768 542
rect 509 504 516 513
rect 531 512 532 513
rect 559 512 560 513
rect 610 512 611 513
rect 638 512 639 513
rect 689 512 690 513
rect 717 512 718 513
rect 522 504 726 507
rect 732 504 739 513
rect 509 491 739 504
rect 531 490 560 491
rect 610 490 639 491
rect 689 490 718 491
rect 509 483 739 490
rect 509 468 516 483
rect 531 477 560 483
rect 610 477 639 483
rect 689 477 718 483
rect 570 469 596 475
rect 531 468 532 469
rect 559 468 560 469
rect 610 468 611 469
rect 638 468 639 469
rect 689 468 690 469
rect 717 468 718 469
rect 732 468 739 483
rect 58 454 64 460
rect 111 454 117 460
rect 481 439 522 468
rect 530 467 561 468
rect 609 467 640 468
rect 688 467 719 468
rect 531 440 560 467
rect 571 455 597 461
rect 610 440 639 467
rect 689 440 718 467
rect 530 439 561 440
rect 609 439 640 440
rect 688 439 719 440
rect 726 439 768 468
rect 52 404 58 410
rect 117 404 123 410
rect 509 389 516 439
rect 531 438 532 439
rect 559 438 560 439
rect 610 438 611 439
rect 638 438 639 439
rect 689 438 690 439
rect 717 438 718 439
rect 732 421 739 439
rect 531 389 532 390
rect 559 389 560 390
rect 610 389 611 390
rect 638 389 639 390
rect 689 389 690 390
rect 717 389 718 390
rect 732 389 739 404
rect 481 360 522 389
rect 530 388 561 389
rect 609 388 640 389
rect 688 388 719 389
rect 531 361 560 388
rect 610 361 639 388
rect 689 361 718 388
rect 530 360 561 361
rect 609 360 640 361
rect 688 360 719 361
rect 726 360 768 389
rect 509 348 516 360
rect 531 359 532 360
rect 559 359 560 360
rect 610 359 611 360
rect 638 359 639 360
rect 689 359 690 360
rect 717 359 718 360
rect 530 348 560 351
rect 609 348 639 351
rect 688 348 718 351
rect 732 348 739 360
rect 509 338 739 348
rect 530 334 560 338
rect 609 334 639 338
rect 688 334 718 338
rect 508 327 738 334
rect 508 312 515 327
rect 530 321 560 327
rect 609 321 639 327
rect 688 321 718 327
rect 570 316 596 319
rect 530 312 531 313
rect 558 312 559 313
rect 609 312 610 313
rect 637 312 638 313
rect 688 312 689 313
rect 716 312 717 313
rect 731 312 738 327
rect 480 283 521 312
rect 529 311 560 312
rect 608 311 639 312
rect 687 311 718 312
rect 530 284 559 311
rect 570 302 596 305
rect 609 284 638 311
rect 688 284 717 311
rect 529 283 560 284
rect 608 283 639 284
rect 687 283 718 284
rect 725 283 767 312
rect 58 265 64 271
rect 111 265 117 271
rect 508 233 515 283
rect 530 282 531 283
rect 558 282 559 283
rect 609 282 610 283
rect 637 282 638 283
rect 688 282 689 283
rect 716 282 717 283
rect 731 263 738 283
rect 530 233 531 234
rect 558 233 559 234
rect 609 233 610 234
rect 637 233 638 234
rect 688 233 689 234
rect 716 233 717 234
rect 731 233 738 246
rect 52 215 58 221
rect 117 215 123 221
rect 480 204 521 233
rect 529 232 560 233
rect 608 232 639 233
rect 687 232 718 233
rect 530 205 559 232
rect 609 205 638 232
rect 688 205 717 232
rect 529 204 560 205
rect 608 204 639 205
rect 687 204 718 205
rect 725 204 767 233
rect 508 194 515 204
rect 530 203 531 204
rect 558 203 559 204
rect 609 203 610 204
rect 637 203 638 204
rect 688 203 689 204
rect 716 203 717 204
rect 521 195 725 197
rect 530 194 559 195
rect 609 194 638 195
rect 688 194 717 195
rect 731 194 738 204
rect 508 182 738 194
rect 530 180 559 182
rect 609 180 638 182
rect 688 180 717 182
rect 508 173 738 180
rect 508 158 515 173
rect 530 167 559 173
rect 609 167 638 173
rect 688 167 717 173
rect 569 160 595 165
rect 530 158 531 159
rect 558 158 559 159
rect 609 158 610 159
rect 637 158 638 159
rect 688 158 689 159
rect 716 158 717 159
rect 731 158 738 173
rect 58 148 64 154
rect 111 148 117 154
rect 480 129 521 158
rect 529 157 560 158
rect 608 157 639 158
rect 687 157 718 158
rect 530 130 559 157
rect 570 146 596 151
rect 609 130 638 157
rect 688 130 717 157
rect 529 129 560 130
rect 608 129 639 130
rect 687 129 718 130
rect 725 129 767 158
rect 52 98 58 104
rect 117 98 123 104
rect 508 79 515 129
rect 530 128 531 129
rect 558 128 559 129
rect 609 128 610 129
rect 637 128 638 129
rect 688 128 689 129
rect 716 128 717 129
rect 731 121 738 129
rect 530 79 531 80
rect 558 79 559 80
rect 609 79 610 80
rect 637 79 638 80
rect 688 79 689 80
rect 716 79 717 80
rect 731 79 738 104
rect 480 50 521 79
rect 529 78 560 79
rect 608 78 639 79
rect 687 78 718 79
rect 530 51 559 78
rect 609 51 638 78
rect 688 51 717 78
rect 529 50 560 51
rect 608 50 639 51
rect 687 50 718 51
rect 725 50 767 79
rect 508 35 515 50
rect 530 49 531 50
rect 558 49 559 50
rect 609 49 610 50
rect 637 49 638 50
rect 688 49 689 50
rect 716 49 717 50
rect 530 35 559 41
rect 609 35 638 41
rect 688 35 717 41
rect 731 35 738 50
rect 508 28 738 35
rect 530 0 559 28
rect 609 0 638 28
rect 688 0 717 28
<< nwell >>
rect 896 341 931 342
rect 896 325 913 341
rect 930 325 931 341
<< poly >>
rect 717 560 753 564
rect 157 527 394 551
rect 717 548 752 560
rect 157 418 392 442
rect 717 404 752 421
rect 913 341 931 342
rect 929 325 931 341
rect 157 238 394 262
rect 584 246 752 263
rect 159 118 396 142
rect 584 104 752 121
<< polycont >>
rect 896 325 913 342
<< locali >>
rect 887 325 896 342
<< viali >>
rect 913 325 931 342
<< metal1 >>
rect 36 31 76 630
rect 918 345 931 347
rect 910 342 934 345
rect 910 325 913 342
rect 931 325 934 342
rect 910 322 934 325
rect 920 318 931 322
<< metal2 >>
rect 0 579 761 586
rect 0 568 764 579
rect 0 525 974 543
rect 0 437 761 443
rect 0 425 764 437
rect 0 393 760 400
rect 0 382 764 393
rect 2 267 764 284
rect 2 225 764 242
rect 2 127 764 144
rect 80 118 234 127
rect 2 83 764 100
use sky130_hilas_wellContact  sky130_hilas_wellContact_1
timestamp 1628285143
transform 1 0 1449 0 1 706
box -1448 -441 -1275 -255
use sky130_hilas_overlapCap01  sky130_hilas_overlapCap01_2
timestamp 1607257541
transform 1 0 767 0 1 225
box -287 -71 0 137
use sky130_hilas_overlapCap01  sky130_hilas_overlapCap01_3
timestamp 1607257541
transform 1 0 767 0 1 71
box -287 -71 0 137
use sky130_hilas_overlapCap01  sky130_hilas_overlapCap01_1
timestamp 1607257541
transform 1 0 768 0 1 381
box -287 -71 0 137
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_0
timestamp 1628285143
transform 1 0 1041 0 1 285
box -289 41 -33 232
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_2
timestamp 1628285143
transform 1 0 1041 0 -1 382
box -289 41 -33 232
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_1
timestamp 1628285143
transform 1 0 1041 0 1 -15
box -289 41 -33 232
use sky130_hilas_overlapCap01  sky130_hilas_overlapCap01_0
timestamp 1607257541
transform 1 0 768 0 1 534
box -287 -71 0 137
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_3
timestamp 1628285143
transform 1 0 1041 0 -1 683
box -289 41 -33 232
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_1
timestamp 1628704213
transform 1 0 1452 0 1 431
box 0 0 173 190
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_0
timestamp 1628704213
transform 1 0 1452 0 1 548
box 0 0 173 190
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_3
timestamp 1628704213
transform 1 0 1452 0 1 846
box 0 0 173 190
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_2
timestamp 1628704213
transform 1 0 1452 0 1 737
box 0 0 173 190
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
