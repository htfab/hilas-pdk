VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_poly2li
  CLASS BLOCK ;
  FOREIGN /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_poly2li ;
  ORIGIN 0.090 0.140 ;
  SIZE 0.270 BY 0.330 ;
  OBS
      LAYER li1 ;
        RECT -0.040 -0.140 0.130 0.190 ;
  END
END /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_poly2li
END LIBRARY

