magic
tech sky130A
timestamp 1629137195
<< checkpaint >>
rect -1247 1675 186 1679
rect 1826 1675 3259 1679
rect -1247 1506 305 1675
rect -1647 60 305 1506
rect -1247 -230 305 60
rect -1178 -235 305 -230
rect 1707 1506 3259 1675
rect 1707 60 3659 1506
rect 1707 -230 3259 60
rect 1707 -235 3190 -230
<< error_s >>
rect 67 616 117 622
rect 139 616 189 622
rect 1823 616 1873 622
rect 1895 616 1945 622
rect 67 574 117 580
rect 139 574 189 580
rect 1823 574 1873 580
rect 1895 574 1945 580
rect 139 547 189 553
rect 1823 547 1873 553
rect 139 505 189 511
rect 1823 505 1873 511
rect 139 462 189 468
rect 1823 462 1873 468
rect 139 420 189 426
rect 1823 420 1873 426
rect 67 393 117 399
rect 139 393 189 399
rect 1823 393 1873 399
rect 1895 393 1945 399
rect 67 351 117 357
rect 139 351 189 357
rect 1823 351 1873 357
rect 1895 351 1945 357
rect 67 292 117 298
rect 139 292 189 298
rect 1823 292 1873 298
rect 1895 292 1945 298
rect 67 250 117 256
rect 139 250 189 256
rect 1823 250 1873 256
rect 1895 250 1945 256
rect 139 223 189 229
rect 1823 223 1873 229
rect 139 181 189 187
rect 1823 181 1873 187
rect 139 139 189 145
rect 1823 139 1873 145
rect 139 97 189 103
rect 1823 97 1873 103
rect 67 70 117 76
rect 139 70 189 76
rect 1823 70 1873 76
rect 1895 70 1945 76
rect 67 28 117 34
rect 139 28 189 34
rect 1823 28 1873 34
rect 1895 28 1945 34
<< nwell >>
rect 1984 609 1993 639
rect 0 391 13 397
rect 0 379 7 391
<< metal1 >>
rect 1961 637 1993 638
rect 21 636 52 637
rect 21 623 24 636
rect 20 610 24 623
rect 50 610 52 636
rect 1961 627 1964 637
rect 77 622 96 627
rect 117 622 133 627
rect 311 618 335 627
rect 529 617 567 627
rect 704 621 728 627
rect 932 614 972 627
rect 1040 617 1080 627
rect 1284 622 1308 627
rect 1445 617 1483 627
rect 1677 620 1701 627
rect 1879 622 1895 627
rect 1916 622 1935 627
rect 20 608 52 610
rect 36 593 52 608
rect 972 591 1040 613
rect 1960 611 1964 627
rect 1990 611 1993 637
rect 1960 610 1993 611
rect 1960 593 1976 610
rect 36 22 52 28
rect 77 23 96 29
rect 117 23 133 29
rect 311 22 335 30
rect 529 22 567 31
rect 704 22 728 29
rect 932 22 972 34
rect 1040 22 1080 34
rect 1284 22 1308 29
rect 1445 22 1483 37
rect 1677 22 1701 28
rect 1879 23 1895 29
rect 1916 23 1935 29
rect 1960 23 1976 29
<< via1 >>
rect 24 610 50 636
rect 1964 611 1990 637
<< metal2 >>
rect 20 637 1994 640
rect 20 636 1964 637
rect 20 610 24 636
rect 50 622 1964 636
rect 50 610 62 622
rect 20 608 62 610
rect 1960 611 1964 622
rect 1990 611 1994 637
rect 1960 609 1994 611
rect 0 576 6 594
rect 2003 576 2012 594
rect 0 533 7 551
rect 2003 533 2012 551
rect 0 422 6 440
rect 2006 422 2012 440
rect 0 379 13 397
rect 2006 379 2012 397
rect 0 252 7 270
rect 2003 252 2012 270
rect 0 209 7 227
rect 2003 209 2012 227
rect 670 160 1346 178
rect 0 99 7 117
rect 2003 99 2012 117
rect 0 56 7 74
rect 2003 56 2012 74
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_0
timestamp 1628285143
transform 1 0 1268 0 1 404
box -263 -404 744 246
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_1
timestamp 1628285143
transform -1 0 744 0 1 404
box -263 -404 744 246
<< labels >>
rlabel metal1 1445 617 1483 627 0 GATE2
port 1 nsew analog default
rlabel metal1 932 22 972 34 0 VTUN
port 2 nsew power default
rlabel metal1 1040 22 1080 34 0 VTUN
port 2 nsew power default
rlabel metal1 1040 617 1080 627 0 VTUN
port 2 nsew power default
rlabel metal1 932 614 972 627 0 VTUN
port 2 nsew power default
rlabel metal1 529 617 567 627 0 GATE1
port 3 nsew analog default
rlabel metal1 529 22 567 31 0 GATE1
port 3 nsew analog default
rlabel metal1 1960 23 1976 29 0 VINJ
port 4 nsew power default
rlabel metal1 1445 22 1483 37 0 GATE2
port 1 nsew analog default
rlabel metal1 1916 622 1935 627 0 SelectGate2
rlabel metal1 1960 622 1976 627 0 VINJ
port 6 nsew power default
rlabel metal1 36 622 52 627 0 VINJ
port 6 nsew power default
rlabel metal1 77 622 96 627 0 GATESELECT1
port 10 nsew analog default
rlabel metal1 36 22 52 28 0 VINJ
port 6 nsew power default
rlabel metal1 77 23 96 29 0 GATESELECT1
port 10 nsew analog default
rlabel metal1 117 622 133 627 0 COL1
port 12 nsew analog default
rlabel metal1 117 23 133 29 0 COL1
port 12 nsew analog default
rlabel metal1 1916 23 1935 29 0 GATESELECT2
port 11 nsew analog default
rlabel metal1 1879 23 1895 29 0 COL2
port 13 nsew analog default
rlabel metal1 1879 622 1895 627 0 COL2
port 13 nsew analog default
rlabel metal1 311 621 335 627 0 VGND
port 22 nsew
rlabel metal1 311 22 335 30 0 VGND
port 22 nsew
rlabel metal1 704 22 728 29 0 VGND
port 22 nsew
rlabel metal1 704 621 728 627 0 VGND
port 22 nsew
rlabel metal1 1284 22 1308 29 0 VGND
port 22 nsew
rlabel metal1 1677 22 1701 28 0 VGND
port 22 nsew
rlabel metal1 1284 622 1308 627 0 VGND
port 22 nsew
rlabel metal1 1677 620 1701 627 0 VGND
port 22 nsew
rlabel metal2 0 56 7 74 0 DRAIN4
port 21 nsew
rlabel metal2 0 99 7 117 0 ROW4
port 20 nsew
rlabel metal2 0 209 7 227 0 ROW3
port 19 nsew
rlabel metal2 0 252 7 270 0 DRAIN3
port 18 nsew
rlabel metal2 0 379 7 397 0 DRAIN2
port 17 nsew
rlabel metal2 0 422 6 440 0 ROW2
port 15 nsew
rlabel metal2 0 533 7 551 0 ROW1
port 14 nsew
rlabel metal2 0 576 6 594 0 DRAIN1
port 16 nsew
rlabel metal2 2003 533 2012 551 0 ROW1
port 14 nsew
rlabel metal2 2006 422 2012 440 0 ROW2
port 15 nsew
rlabel metal2 2006 379 2012 397 0 DRAIN2
port 17 nsew
rlabel metal2 2003 252 2012 270 0 DRAIN3
port 18 nsew
rlabel metal2 2003 209 2012 227 0 ROW3
port 19 nsew
rlabel metal2 2003 99 2012 117 0 ROW4
port 20 nsew
rlabel metal2 2003 56 2012 74 0 DRAIN4
port 21 nsew
rlabel metal2 2003 576 2012 594 0 DRAIN1
port 16 nsew
<< end >>
