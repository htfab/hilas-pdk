magic
tech sky130A
timestamp 1628704266
<< checkpaint >>
rect -630 1240 886 1246
rect 911 1240 2427 1246
rect -630 -625 2427 1240
rect -630 -630 886 -625
rect 911 -630 2427 -625
<< error_s >>
rect 323 577 352 593
rect 402 577 431 593
rect 481 577 510 593
rect 560 577 589 593
rect 806 579 835 597
rect 962 579 991 597
rect 1208 577 1237 593
rect 1287 577 1316 593
rect 1366 577 1395 593
rect 1445 577 1474 593
rect 806 547 807 548
rect 834 547 835 548
rect 962 547 963 548
rect 990 547 991 548
rect 323 543 324 544
rect 351 543 352 544
rect 402 543 403 544
rect 430 543 431 544
rect 481 543 482 544
rect 509 543 510 544
rect 560 543 561 544
rect 588 543 589 544
rect 273 514 290 543
rect 322 542 353 543
rect 401 542 432 543
rect 480 542 511 543
rect 559 542 590 543
rect 323 535 352 542
rect 402 535 431 542
rect 481 535 510 542
rect 560 535 589 542
rect 323 521 332 535
rect 579 521 589 535
rect 323 515 352 521
rect 402 515 431 521
rect 481 515 510 521
rect 560 515 589 521
rect 322 514 353 515
rect 401 514 432 515
rect 480 514 511 515
rect 559 514 590 515
rect 621 514 639 543
rect 756 518 774 547
rect 805 546 836 547
rect 806 537 835 546
rect 806 528 816 537
rect 825 528 835 537
rect 806 519 835 528
rect 805 518 836 519
rect 867 518 885 547
rect 912 518 930 547
rect 961 546 992 547
rect 962 537 991 546
rect 962 528 972 537
rect 981 528 991 537
rect 962 519 991 528
rect 961 518 992 519
rect 1023 518 1041 547
rect 1208 543 1209 544
rect 1236 543 1237 544
rect 1287 543 1288 544
rect 1315 543 1316 544
rect 1366 543 1367 544
rect 1394 543 1395 544
rect 1445 543 1446 544
rect 1473 543 1474 544
rect 806 517 807 518
rect 834 517 835 518
rect 962 517 963 518
rect 990 517 991 518
rect 1158 514 1176 543
rect 1207 542 1238 543
rect 1286 542 1317 543
rect 1365 542 1396 543
rect 1444 542 1475 543
rect 1208 535 1237 542
rect 1287 535 1316 542
rect 1366 535 1395 542
rect 1445 535 1474 542
rect 1208 521 1218 535
rect 1465 521 1474 535
rect 1208 515 1237 521
rect 1287 515 1316 521
rect 1366 515 1395 521
rect 1445 515 1474 521
rect 1207 514 1238 515
rect 1286 514 1317 515
rect 1365 514 1396 515
rect 1444 514 1475 515
rect 1507 514 1524 543
rect 1541 521 1543 522
rect 323 513 324 514
rect 351 513 352 514
rect 402 513 403 514
rect 430 513 431 514
rect 481 513 482 514
rect 509 513 510 514
rect 560 513 561 514
rect 588 513 589 514
rect 1208 513 1209 514
rect 1236 513 1237 514
rect 1287 513 1288 514
rect 1315 513 1316 514
rect 1366 513 1367 514
rect 1394 513 1395 514
rect 1445 513 1446 514
rect 1473 513 1474 514
rect 323 464 352 479
rect 402 464 431 479
rect 481 464 510 479
rect 560 464 589 479
rect 806 468 835 486
rect 962 468 991 486
rect 1208 464 1237 479
rect 1287 464 1316 479
rect 1366 464 1395 479
rect 1445 464 1474 479
rect 323 430 352 446
rect 402 430 431 446
rect 481 430 510 446
rect 560 430 589 446
rect 806 427 835 445
rect 962 427 991 445
rect 1208 430 1237 446
rect 1287 430 1316 446
rect 1366 430 1395 446
rect 1445 430 1474 446
rect 323 396 324 397
rect 351 396 352 397
rect 402 396 403 397
rect 430 396 431 397
rect 481 396 482 397
rect 509 396 510 397
rect 560 396 561 397
rect 588 396 589 397
rect 1208 396 1209 397
rect 1236 396 1237 397
rect 1287 396 1288 397
rect 1315 396 1316 397
rect 1366 396 1367 397
rect 1394 396 1395 397
rect 1445 396 1446 397
rect 1473 396 1474 397
rect 273 367 290 396
rect 322 395 353 396
rect 401 395 432 396
rect 480 395 511 396
rect 559 395 590 396
rect 323 388 352 395
rect 402 388 431 395
rect 481 388 510 395
rect 560 388 589 395
rect 323 374 332 388
rect 579 374 589 388
rect 323 368 352 374
rect 402 368 431 374
rect 481 368 510 374
rect 560 368 589 374
rect 322 367 353 368
rect 401 367 432 368
rect 480 367 511 368
rect 559 367 590 368
rect 621 367 639 396
rect 806 395 807 396
rect 834 395 835 396
rect 962 395 963 396
rect 990 395 991 396
rect 323 366 324 367
rect 351 366 352 367
rect 402 366 403 367
rect 430 366 431 367
rect 481 366 482 367
rect 509 366 510 367
rect 560 366 561 367
rect 588 366 589 367
rect 756 366 774 395
rect 805 394 836 395
rect 806 385 835 394
rect 806 376 816 385
rect 825 376 835 385
rect 806 367 835 376
rect 805 366 836 367
rect 867 366 885 395
rect 912 366 930 395
rect 961 394 992 395
rect 962 385 991 394
rect 962 376 972 385
rect 981 376 991 385
rect 962 367 991 376
rect 961 366 992 367
rect 1023 366 1041 395
rect 1158 367 1176 396
rect 1207 395 1238 396
rect 1286 395 1317 396
rect 1365 395 1396 396
rect 1444 395 1475 396
rect 1208 388 1237 395
rect 1287 388 1316 395
rect 1366 388 1395 395
rect 1445 388 1474 395
rect 1208 374 1218 388
rect 1465 374 1474 388
rect 1208 368 1237 374
rect 1287 368 1316 374
rect 1366 368 1395 374
rect 1445 368 1474 374
rect 1207 367 1238 368
rect 1286 367 1317 368
rect 1365 367 1396 368
rect 1444 367 1475 368
rect 1507 367 1524 396
rect 1208 366 1209 367
rect 1236 366 1237 367
rect 1287 366 1288 367
rect 1315 366 1316 367
rect 1366 366 1367 367
rect 1394 366 1395 367
rect 1445 366 1446 367
rect 1473 366 1474 367
rect 806 365 807 366
rect 834 365 835 366
rect 962 365 963 366
rect 990 365 991 366
rect 323 317 352 332
rect 402 317 431 332
rect 481 317 510 332
rect 560 317 589 332
rect 806 316 835 334
rect 962 316 991 334
rect 1208 317 1237 332
rect 1287 317 1316 332
rect 1366 317 1395 332
rect 1445 317 1474 332
rect 323 283 352 299
rect 402 283 431 299
rect 481 283 510 299
rect 560 283 589 299
rect 806 282 835 300
rect 962 282 991 300
rect 1208 283 1237 299
rect 1287 283 1316 299
rect 1366 283 1395 299
rect 1445 283 1474 299
rect 806 250 807 251
rect 834 250 835 251
rect 962 250 963 251
rect 990 250 991 251
rect 323 249 324 250
rect 351 249 352 250
rect 402 249 403 250
rect 430 249 431 250
rect 481 249 482 250
rect 509 249 510 250
rect 560 249 561 250
rect 588 249 589 250
rect 273 220 290 249
rect 322 248 353 249
rect 401 248 432 249
rect 480 248 511 249
rect 559 248 590 249
rect 323 241 352 248
rect 402 241 431 248
rect 481 241 510 248
rect 560 241 589 248
rect 323 227 332 241
rect 579 227 589 241
rect 323 221 352 227
rect 402 221 431 227
rect 481 221 510 227
rect 560 221 589 227
rect 322 220 353 221
rect 401 220 432 221
rect 480 220 511 221
rect 559 220 590 221
rect 621 220 639 249
rect 756 221 774 250
rect 805 249 836 250
rect 806 240 835 249
rect 806 231 816 240
rect 825 231 835 240
rect 806 222 835 231
rect 805 221 836 222
rect 867 221 885 250
rect 912 221 930 250
rect 961 249 992 250
rect 962 240 991 249
rect 962 231 972 240
rect 981 231 991 240
rect 962 222 991 231
rect 961 221 992 222
rect 1023 221 1041 250
rect 1208 249 1209 250
rect 1236 249 1237 250
rect 1287 249 1288 250
rect 1315 249 1316 250
rect 1366 249 1367 250
rect 1394 249 1395 250
rect 1445 249 1446 250
rect 1473 249 1474 250
rect 806 220 807 221
rect 834 220 835 221
rect 962 220 963 221
rect 990 220 991 221
rect 1158 220 1176 249
rect 1207 248 1238 249
rect 1286 248 1317 249
rect 1365 248 1396 249
rect 1444 248 1475 249
rect 1208 241 1237 248
rect 1287 241 1316 248
rect 1366 241 1395 248
rect 1445 241 1474 248
rect 1208 227 1218 241
rect 1465 227 1474 241
rect 1208 221 1237 227
rect 1287 221 1316 227
rect 1366 221 1395 227
rect 1445 221 1474 227
rect 1207 220 1238 221
rect 1286 220 1317 221
rect 1365 220 1396 221
rect 1444 220 1475 221
rect 1507 220 1524 249
rect 323 219 324 220
rect 351 219 352 220
rect 402 219 403 220
rect 430 219 431 220
rect 481 219 482 220
rect 509 219 510 220
rect 560 219 561 220
rect 588 219 589 220
rect 1208 219 1209 220
rect 1236 219 1237 220
rect 1287 219 1288 220
rect 1315 219 1316 220
rect 1366 219 1367 220
rect 1394 219 1395 220
rect 1445 219 1446 220
rect 1473 219 1474 220
rect 323 170 352 185
rect 402 170 431 185
rect 481 170 510 185
rect 560 170 589 185
rect 806 171 835 189
rect 962 171 991 189
rect 1208 170 1237 185
rect 1287 170 1316 185
rect 1366 170 1395 185
rect 1445 170 1474 185
rect 323 136 352 152
rect 402 136 431 152
rect 481 136 510 152
rect 560 136 589 152
rect 806 128 835 146
rect 962 128 991 146
rect 1208 136 1237 152
rect 1287 136 1316 152
rect 1366 136 1395 152
rect 1445 136 1474 152
rect 323 102 324 103
rect 351 102 352 103
rect 402 102 403 103
rect 430 102 431 103
rect 481 102 482 103
rect 509 102 510 103
rect 560 102 561 103
rect 588 102 589 103
rect 1208 102 1209 103
rect 1236 102 1237 103
rect 1287 102 1288 103
rect 1315 102 1316 103
rect 1366 102 1367 103
rect 1394 102 1395 103
rect 1445 102 1446 103
rect 1473 102 1474 103
rect 273 73 290 102
rect 322 101 353 102
rect 401 101 432 102
rect 480 101 511 102
rect 559 101 590 102
rect 323 94 352 101
rect 402 94 431 101
rect 481 94 510 101
rect 560 94 589 101
rect 323 80 332 94
rect 579 80 589 94
rect 323 74 352 80
rect 402 74 431 80
rect 481 74 510 80
rect 560 74 589 80
rect 322 73 353 74
rect 401 73 432 74
rect 480 73 511 74
rect 559 73 590 74
rect 621 73 639 102
rect 806 96 807 97
rect 834 96 835 97
rect 962 96 963 97
rect 990 96 991 97
rect 323 72 324 73
rect 351 72 352 73
rect 402 72 403 73
rect 430 72 431 73
rect 481 72 482 73
rect 509 72 510 73
rect 560 72 561 73
rect 588 72 589 73
rect 756 67 774 96
rect 805 95 836 96
rect 806 86 835 95
rect 806 77 816 86
rect 825 77 835 86
rect 806 68 835 77
rect 805 67 836 68
rect 867 67 885 96
rect 912 67 930 96
rect 961 95 992 96
rect 962 86 991 95
rect 962 77 972 86
rect 981 77 991 86
rect 962 68 991 77
rect 961 67 992 68
rect 1023 67 1041 96
rect 1158 73 1176 102
rect 1207 101 1238 102
rect 1286 101 1317 102
rect 1365 101 1396 102
rect 1444 101 1475 102
rect 1208 94 1237 101
rect 1287 94 1316 101
rect 1366 94 1395 101
rect 1445 94 1474 101
rect 1208 80 1218 94
rect 1465 80 1474 94
rect 1208 74 1237 80
rect 1287 74 1316 80
rect 1366 74 1395 80
rect 1445 74 1474 80
rect 1207 73 1238 74
rect 1286 73 1317 74
rect 1365 73 1396 74
rect 1444 73 1475 74
rect 1507 73 1524 102
rect 1208 72 1209 73
rect 1236 72 1237 73
rect 1287 72 1288 73
rect 1315 72 1316 73
rect 1366 72 1367 73
rect 1394 72 1395 73
rect 1445 72 1446 73
rect 1473 72 1474 73
rect 806 66 807 67
rect 834 66 835 67
rect 962 66 963 67
rect 990 66 991 67
rect 323 23 352 38
rect 402 23 431 38
rect 481 23 510 38
rect 560 23 589 38
rect 806 17 835 35
rect 962 17 991 35
rect 1208 23 1237 38
rect 1287 23 1316 38
rect 1366 23 1395 38
rect 1445 23 1474 38
<< metal1 >>
rect 36 604 52 610
rect 77 604 96 610
rect 117 604 133 610
rect 36 6 52 13
rect 77 6 96 13
rect 117 6 133 13
rect 444 5 469 610
rect 805 5 835 610
rect 963 5 993 610
rect 1329 5 1353 610
rect 1664 603 1680 610
rect 1701 603 1720 610
rect 1745 603 1761 610
rect 1664 6 1680 13
rect 1701 6 1720 13
rect 1745 6 1761 13
<< metal2 >>
rect 0 542 8 560
rect 1786 542 1797 560
rect 0 499 8 517
rect 1787 499 1798 517
rect 0 399 8 417
rect 1787 399 1798 417
rect 0 356 8 374
rect 240 366 252 374
rect 1549 360 1561 374
rect 1787 356 1798 374
rect 0 241 7 259
rect 1786 241 1797 259
rect 0 198 7 216
rect 1786 198 1797 216
rect 0 99 7 117
rect 1786 99 1797 117
rect 0 56 7 74
rect 1786 56 1797 74
use sky130_hilas_swc4x1cellOverlap2  sky130_hilas_swc4x1cellOverlap2_0
timestamp 1607392100
transform 1 0 1053 0 1 387
box -191 -387 744 229
use sky130_hilas_swc4x1cellOverlap2  sky130_hilas_swc4x1cellOverlap2_1
timestamp 1607392100
transform -1 0 744 0 1 387
box -191 -387 744 229
<< labels >>
rlabel metal1 117 604 133 610 0 VERT1
port 1 nsew analog default
rlabel metal1 36 604 52 610 0 VINJ
port 10 nsew
rlabel metal1 77 604 96 610 0 GATESELECT1
port 11 nsew analog default
rlabel metal2 0 542 8 560 0 DRAIN1
port 3 nsew analog default
rlabel metal2 0 499 8 517 0 HORIZ1
port 2 nsew analog default
rlabel metal2 0 399 8 417 0 HORIZ2
port 4 nsew analog default
rlabel metal2 0 356 8 374 0 DRAIN2
port 5 nsew analog default
rlabel metal2 0 241 7 259 0 DRAIN3
port 6 nsew analog default
rlabel metal2 0 198 7 216 0 HORIZ3
port 7 nsew analog default
rlabel metal2 0 99 7 117 0 HORIZ4
port 8 nsew analog default
rlabel metal2 0 56 7 74 0 DRAIN4
port 9 nsew analog default
rlabel metal1 36 6 52 13 0 VINJ
port 10 nsew power default
rlabel metal1 117 6 133 13 0 VERT1
port 1 nsew analog default
rlabel metal1 77 6 96 13 0 GATESELECT1
port 11 nsew analog default
rlabel metal1 1745 6 1761 13 0 VINJ
port 10 nsew power default
rlabel metal1 1664 603 1680 610 0 VERT2
port 12 nsew analog default
rlabel metal1 1701 603 1720 610 0 GATESELECT2
port 13 nsew analog default
rlabel metal1 1745 603 1761 610 0 VINJ
port 10 nsew power default
rlabel metal1 1664 6 1680 13 0 VERT2
port 12 nsew analog default
rlabel metal1 1701 6 1720 13 0 GATESELECT2
port 13 nsew analog default
rlabel metal2 1786 542 1797 560 0 DRAIN1
port 3 nsew analog default
rlabel metal2 1787 499 1798 517 0 HORIZ1
port 2 nsew analog default
rlabel metal2 1787 399 1798 417 0 HORIZ2
port 4 nsew analog default
rlabel metal2 1787 356 1798 374 0 DRAIN2
port 5 nsew analog default
rlabel metal2 1786 241 1797 259 0 DRAIN3
port 6 nsew analog default
rlabel metal2 1786 198 1797 216 0 HORIZ3
port 7 nsew analog default
rlabel metal2 1786 99 1797 117 0 HORIZ4
port 8 nsew analog default
rlabel metal2 1786 56 1797 74 0 DRAIN
port 14 nsew analog default
rlabel metal1 1329 605 1353 610 0 GATE2
port 15 nsew analog default
rlabel metal1 1329 5 1353 11 0 GATE2
port 15 nsew analog default
rlabel metal1 444 604 469 610 0 GATE1
port 16 nsew analog default
rlabel metal1 444 5 469 11 0 GATE1
port 16 nsew analog default
rlabel metal1 805 602 835 610 0 VTUN
port 17 nsew analog default
rlabel metal1 963 602 993 610 0 VTUN
rlabel metal1 805 5 835 13 0 VTUN
port 17 nsew analog default
rlabel metal1 963 5 993 13 0 VTUN
port 17 nsew analog default
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
