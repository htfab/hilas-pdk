magic
tech sky130A
timestamp 1627737364
<< error_s >>
rect 555 189 605 200
rect 627 189 677 200
rect 523 158 555 159
rect 555 147 605 158
rect 627 147 677 158
rect 555 127 605 139
rect 526 126 555 127
rect 632 97 636 127
rect 555 85 605 97
rect -2 82 15 84
rect 400 79 417 81
rect -2 63 15 65
rect 400 60 417 62
rect 555 45 605 57
rect 526 15 555 16
rect 632 15 636 45
rect 555 3 605 15
rect 555 -16 605 -5
rect 627 -16 677 -5
rect 523 -17 555 -16
rect 401 -39 418 -37
rect -1 -45 16 -43
rect 401 -58 418 -56
rect 555 -58 605 -47
rect 627 -58 677 -47
rect -1 -64 16 -62
rect 401 -73 418 -71
rect -1 -79 16 -77
rect 401 -92 418 -90
rect -1 -98 16 -96
rect 401 -107 418 -105
rect -1 -113 16 -111
rect 555 -112 605 -101
rect 627 -112 677 -101
rect 401 -126 418 -124
rect -1 -132 16 -130
rect 523 -143 555 -142
rect -1 -147 16 -145
rect 555 -154 605 -143
rect 627 -154 677 -143
rect 555 -174 605 -162
rect 526 -175 555 -174
rect 632 -204 636 -174
rect 555 -216 605 -204
rect 555 -255 605 -243
rect 526 -285 555 -284
rect 632 -285 636 -255
rect 555 -297 605 -285
rect 555 -316 605 -305
rect 627 -316 677 -305
rect 523 -317 555 -316
rect 555 -358 605 -347
rect 627 -358 677 -347
<< nwell >>
rect 112 220 335 223
rect -264 37 -263 160
rect 488 -21 497 -13
rect 632 -72 667 -71
rect 632 -88 649 -72
rect 666 -88 667 -72
rect 112 -382 335 -380
<< psubdiff >>
rect -6 82 19 105
rect -6 65 -2 82
rect 15 65 19 82
rect -6 37 19 65
rect 396 79 421 107
rect 396 62 400 79
rect 417 62 421 79
rect 396 36 421 62
rect -6 -45 20 -3
rect -6 -62 -1 -45
rect 16 -62 20 -45
rect -6 -79 20 -62
rect -6 -96 -1 -79
rect 16 -96 20 -79
rect -6 -113 20 -96
rect -6 -130 -1 -113
rect 16 -130 20 -113
rect -6 -143 20 -130
rect 396 -39 423 -18
rect 396 -56 401 -39
rect 418 -56 423 -39
rect 396 -73 423 -56
rect 396 -90 401 -73
rect 418 -90 423 -73
rect 396 -107 423 -90
rect 396 -124 401 -107
rect 418 -124 423 -107
rect 396 -142 423 -124
rect -1 -147 16 -143
<< psubdiffcont >>
rect -2 65 15 82
rect 400 62 417 79
rect -1 -62 16 -45
rect -1 -96 16 -79
rect -1 -130 16 -113
rect 401 -56 418 -39
rect 401 -90 418 -73
rect 401 -124 418 -107
<< poly >>
rect 319 147 489 151
rect -107 114 130 138
rect 319 135 488 147
rect -107 5 128 29
rect 319 -9 488 8
rect 649 -72 667 -71
rect 665 -88 667 -72
rect -107 -175 130 -151
rect 320 -167 488 -150
rect -105 -295 132 -271
rect 320 -309 488 -292
<< polycont >>
rect 632 -88 649 -71
<< locali >>
rect 623 -88 632 -71
<< viali >>
rect -2 82 15 99
rect -2 48 15 65
rect 400 79 417 96
rect 400 45 417 62
rect -1 -45 16 -28
rect -1 -79 16 -62
rect -1 -113 16 -96
rect -1 -147 16 -130
rect 401 -39 418 -22
rect 401 -73 418 -56
rect 649 -88 667 -71
rect 401 -107 418 -90
rect 401 -141 418 -124
<< metal1 >>
rect -228 -382 -188 223
rect -7 99 20 223
rect 177 213 215 223
rect -7 82 -2 99
rect 15 82 20 99
rect -7 65 20 82
rect -7 48 -2 65
rect 15 48 20 65
rect -7 -28 20 48
rect -7 -45 -1 -28
rect 16 -45 20 -28
rect -7 -62 20 -45
rect -7 -79 -1 -62
rect 16 -79 20 -62
rect -7 -96 20 -79
rect -7 -113 -1 -96
rect 16 -113 20 -96
rect -7 -130 20 -113
rect -7 -147 -1 -130
rect 16 -147 20 -130
rect -7 -224 20 -147
rect 396 96 421 223
rect 611 216 627 223
rect 648 216 667 223
rect 692 216 708 223
rect 396 79 400 96
rect 417 79 421 96
rect 396 62 421 79
rect 396 45 400 62
rect 417 45 421 62
rect 396 -22 421 45
rect 396 -39 401 -22
rect 418 -39 421 -22
rect 396 -56 421 -39
rect 396 -73 401 -56
rect 418 -73 421 -56
rect 654 -68 667 -66
rect 396 -90 421 -73
rect 396 -107 401 -90
rect 418 -107 421 -90
rect 646 -71 670 -68
rect 646 -88 649 -71
rect 667 -88 670 -71
rect 646 -91 670 -88
rect 656 -95 667 -91
rect 396 -124 421 -107
rect 396 -141 401 -124
rect 418 -141 421 -124
rect 396 -221 421 -141
rect 395 -224 423 -221
rect -9 -227 22 -224
rect -9 -253 -7 -227
rect 20 -253 22 -227
rect 394 -225 424 -224
rect 394 -251 396 -225
rect 422 -251 424 -225
rect 394 -252 424 -251
rect -9 -255 22 -253
rect 395 -254 423 -252
rect -7 -382 20 -255
rect 177 -382 215 -372
rect 396 -382 421 -254
rect 611 -381 627 -374
rect 648 -381 667 -374
rect 692 -381 708 -374
<< via1 >>
rect -7 -253 20 -227
rect 396 -251 422 -225
<< metal2 >>
rect 487 166 497 173
rect 487 155 500 166
rect 735 155 744 173
rect -264 112 540 130
rect 735 112 744 130
rect -264 111 -249 112
rect -266 30 -252 32
rect -266 24 497 30
rect -266 12 500 24
rect 736 12 745 30
rect 488 -20 497 -17
rect 488 -31 500 -20
rect 735 -31 744 -13
rect 485 -146 500 -129
rect 734 -146 745 -128
rect -263 -187 500 -171
rect -262 -188 500 -187
rect 733 -189 744 -171
rect 393 -225 425 -224
rect -10 -253 -7 -227
rect 20 -230 23 -227
rect 393 -230 396 -225
rect 20 -247 396 -230
rect 20 -253 23 -247
rect 393 -251 396 -247
rect 422 -251 425 -225
rect 393 -252 425 -251
rect -263 -286 500 -269
rect -184 -295 -30 -286
rect 733 -288 744 -270
rect 487 -330 500 -313
rect 733 -331 744 -313
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_1
timestamp 1627737364
transform 1 0 1188 0 1 18
box -1451 -400 -1278 -210
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_0
timestamp 1627737364
transform 1 0 1188 0 1 135
box -1451 -400 -1278 -210
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_0
timestamp 1627737364
transform 1 0 1069 0 1 14
box -957 -395 -734 -209
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_1
timestamp 1627737364
transform 1 0 1069 0 1 130
box -957 -395 -734 -209
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_1
timestamp 1627737364
transform 1 0 777 0 1 -428
box -289 47 -33 232
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_2
timestamp 1627737364
transform 1 0 777 0 -1 -31
box -289 47 -33 232
use sky130_hilas_wellContact  sky130_hilas_wellContact_1
timestamp 1627737364
transform 1 0 1185 0 1 293
box -1449 -441 -1275 -255
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_2
timestamp 1627737364
transform 1 0 1188 0 1 324
box -1451 -400 -1278 -210
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_2
timestamp 1627737364
transform 1 0 1069 0 1 315
box -957 -395 -734 -209
use sky130_hilas_wellContact  sky130_hilas_wellContact_0
timestamp 1627737364
transform 1 0 1588 0 1 286
box -1449 -441 -1275 -255
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_0
timestamp 1627737364
transform 1 0 777 0 1 -128
box -289 47 -33 232
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_3
timestamp 1627737364
transform 1 0 1188 0 1 433
box -1451 -400 -1278 -210
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_3
timestamp 1627737364
transform 1 0 1069 0 1 432
box -957 -395 -734 -209
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_3
timestamp 1627737364
transform 1 0 777 0 -1 270
box -289 47 -33 232
<< labels >>
rlabel metal2 -264 111 -252 130 0 ROW1
port 1 nsew analog default
rlabel metal2 -266 13 -254 32 0 ROW2
port 2 nsew analog default
rlabel metal2 -263 -187 -251 -171 0 ROW3
port 3 nsew analog default
rlabel metal2 -263 -285 -249 -270 0 ROW4
port 4 nsew analog default
rlabel metal1 -228 209 -188 223 0 VTUN
port 5 nsew analog default
rlabel metal1 -228 -382 -188 -372 0 VTUN
port 5 nsew analog default
rlabel metal1 177 -382 215 -372 0 GATE1
port 6 nsew analog default
rlabel metal1 177 213 215 223 0 GATE1
port 6 nsew analog default
rlabel metal1 692 216 708 223 0 VINJ
port 7 nsew power default
rlabel metal1 611 216 627 223 0 VPWR
port 8 nsew power default
rlabel metal1 648 216 667 223 0 COLSEL1
rlabel metal1 692 -381 708 -374 0 VINJ
port 7 nsew power default
rlabel metal1 611 -381 627 -374 0 VPWR
port 8 nsew power default
rlabel metal1 648 -381 667 -374 0 COLSEL1
port 9 nsew analog default
rlabel metal2 735 155 744 173 0 DRAIN1
port 10 nsew analog default
rlabel metal2 735 112 744 130 0 ROW1
port 11 nsew analog default
rlabel metal2 735 -31 744 -13 0 DRAIN2
port 13 nsew
rlabel metal2 736 12 745 30 0 ROW2
port 12 nsew analog default
rlabel metal2 734 -146 745 -128 0 DRAIN3
port 14 nsew analog default
rlabel metal2 733 -189 744 -171 0 ROW3
port 15 nsew analog default
rlabel metal2 733 -288 744 -270 0 ROW4
port 16 nsew analog default
rlabel metal2 733 -331 744 -313 0 DRAIN4
port 17 nsew analog default
rlabel metal1 -7 215 20 223 0 VGND
port 18 nsew
rlabel metal1 396 218 421 223 0 VGND
port 18 nsew
rlabel metal1 -7 -382 20 -375 0 VGND
port 18 nsew
rlabel metal1 396 -382 421 -375 0 VGND
port 18 nsew
<< end >>
