magic
tech sky130A
timestamp 1627062261
<< error_s >>
rect 59 532 65 538
rect 112 532 118 538
rect 53 482 59 488
rect 118 482 124 488
rect 482 473 488 479
rect 587 473 593 479
rect 476 423 482 429
rect 593 423 599 429
rect 482 172 488 178
rect 587 172 593 178
rect 59 118 65 124
rect 112 118 118 124
rect 476 122 482 128
rect 593 122 599 128
rect 53 68 59 74
rect 118 68 124 74
<< nwell >>
rect 60 140 116 382
<< psubdiff >>
rect 302 340 327 483
rect 302 323 305 340
rect 324 323 327 340
rect 302 310 327 323
rect 302 307 664 310
rect 302 306 543 307
rect 302 289 326 306
rect 345 289 369 306
rect 388 289 413 306
rect 432 289 453 306
rect 472 289 497 306
rect 516 290 543 306
rect 562 306 664 307
rect 562 290 587 306
rect 516 289 587 290
rect 606 289 633 306
rect 652 289 664 306
rect 302 285 664 289
rect 302 272 327 285
rect 302 255 305 272
rect 324 255 327 272
rect 302 101 327 255
<< mvnsubdiff >>
rect 60 140 116 382
<< psubdiffcont >>
rect 305 323 324 340
rect 326 289 345 306
rect 369 289 388 306
rect 413 289 432 306
rect 453 289 472 306
rect 497 289 516 306
rect 543 290 562 307
rect 587 289 606 306
rect 633 289 652 306
rect 305 255 324 272
<< poly >>
rect 191 533 690 583
rect 160 516 729 533
rect 160 508 718 516
rect 442 473 461 508
rect 617 472 634 508
rect 443 89 460 122
rect 617 89 634 122
rect 117 72 728 89
rect 195 15 695 72
<< locali >>
rect 188 504 694 587
rect 195 496 243 504
rect 228 471 243 496
rect 864 410 867 427
rect 305 340 324 348
rect 864 331 869 348
rect 305 307 324 323
rect 305 306 543 307
rect 305 289 326 306
rect 345 289 369 306
rect 388 289 413 306
rect 432 289 453 306
rect 472 289 497 306
rect 516 290 543 306
rect 562 306 660 307
rect 562 290 587 306
rect 516 289 587 290
rect 606 289 633 306
rect 652 289 660 306
rect 305 272 324 289
rect 871 274 888 331
rect 864 257 866 274
rect 305 247 324 255
rect 408 185 431 189
rect 864 178 867 195
rect 225 103 227 128
rect 192 95 227 103
rect 192 10 697 95
<< metal1 >>
rect 36 1 78 605
rect 284 508 307 605
rect 284 483 308 508
rect 284 0 307 483
rect 406 0 429 605
rect 1058 599 1077 605
rect 1058 0 1077 6
rect 1102 0 1130 605
<< metal2 >>
rect 1 537 913 555
rect 180 495 226 496
rect 1 479 226 495
rect 1 477 195 479
rect 951 452 1154 453
rect 1 431 1154 452
rect 1 430 1023 431
rect 1 333 1047 355
rect 1019 284 1045 319
rect 1 156 1154 177
rect 1 155 1023 156
rect 1 103 196 124
rect 907 67 923 69
rect 1 62 923 67
rect 1 52 911 62
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_1
timestamp 1608066871
transform 1 0 1453 0 1 401
box -1451 -400 -1278 -210
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_3
timestamp 1608066871
transform 1 0 1453 0 1 815
box -1451 -400 -1278 -210
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1607089160
transform 1 0 206 0 1 114
box -14 -15 20 18
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_0
timestamp 1606868103
transform 1 0 1383 0 1 444
box -1005 -380 -733 -211
use sky130_hilas_wellContact  sky130_hilas_wellContact_0
timestamp 1606753443
transform 1 0 1451 0 1 613
box -1449 -441 -1275 -255
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_2
timestamp 1606868103
transform 1 0 1383 0 -1 151
box -1005 -380 -733 -211
use sky130_hilas_wellContact  sky130_hilas_wellContact_1
timestamp 1606753443
transform 1 0 1451 0 1 786
box -1449 -441 -1275 -255
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1607179295
transform 1 0 294 0 1 290
box -10 -8 13 21
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1607089160
transform 1 0 209 0 1 483
box -14 -15 20 18
use sky130_hilas_horizTransCell01  sky130_hilas_horizTransCell01_1
timestamp 1625488390
transform 1 0 1187 0 -1 652
box -476 48 -33 359
use sky130_hilas_horizTransCell01  sky130_hilas_horizTransCell01_0
timestamp 1625488390
transform 1 0 1187 0 1 -47
box -476 48 -33 359
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1607949437
transform 1 0 1024 0 1 326
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1607949437
transform 1 0 1024 0 1 266
box -9 -10 23 22
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1607089160
transform 1 0 935 0 1 166
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1607089160
transform 1 0 935 0 1 442
box -14 -15 20 18
<< labels >>
rlabel metal1 36 598 78 605 0 VTUN
port 9 nsew analog default
rlabel metal1 284 598 307 605 0 VGND
port 7 nsew ground default
rlabel metal1 406 597 429 605 0 GATE1
port 8 nsew analog default
rlabel metal1 1102 598 1130 605 0 VINJ
port 5 nsew power default
rlabel metal2 1146 431 1154 453 0 ROW1
port 3 nsew analog default
rlabel metal2 1147 156 1154 177 0 ROW2
port 4 nsew analog default
rlabel metal2 1 537 8 555 0 DRAIN1
port 1 nsew analog default
rlabel metal2 1 477 6 495 0 VIN11
port 2 nsew
rlabel metal1 1058 599 1077 604 0 COLSEL1
port 6 nsew analog default
rlabel metal1 1058 0 1077 6 0 COLSEL1
port 6 nsew analog default
rlabel metal1 1102 0 1130 7 0 VINJ
port 5 nsew power default
rlabel metal1 284 0 307 10 0 VGND
port 7 nsew ground default
rlabel metal1 406 0 429 8 0 GATE1
port 10 nsew analog default
rlabel metal2 1 52 6 67 0 DRAIN2
port 11 nsew analog default
rlabel metal2 1 103 7 124 0 VIN12
port 12 nsew analog default
rlabel metal2 1 333 7 355 0 COMMONSOURCE
port 13 nsew analog default
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
