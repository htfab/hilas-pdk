magic
tech sky130A
timestamp 1628616981
<< checkpaint >>
rect -687 1155 1141 1200
rect -687 -630 1373 1155
rect -687 -675 1141 -630
<< metal2 >>
rect 0 514 73 515
rect 0 498 142 514
rect 0 497 73 498
rect 0 327 67 329
rect 0 311 139 327
rect 0 212 70 213
rect 0 196 143 212
rect 0 12 146 29
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_0
timestamp 1628616972
transform 1 0 175 0 1 293
box 0 0 568 170
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_3
timestamp 1628616972
transform 1 0 175 0 -1 232
box 0 0 568 170
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_1
timestamp 1628616972
transform 1 0 175 0 -1 525
box 0 0 568 170
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_2
timestamp 1628616972
transform 1 0 175 0 1 0
box 0 0 568 170
<< labels >>
rlabel metal2 0 497 5 515 0 drain1
rlabel metal2 0 311 5 329 0 drain2
rlabel metal2 0 196 5 213 0 drain3
rlabel metal2 0 12 5 29 0 drain4
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
