VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_WTA4Stage01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_WTA4Stage01 ;
  ORIGIN 11.210 0.430 ;
  SIZE 14.170 BY 6.050 ;
  PIN GND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2.570 4.530 2.800 5.620 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.570 -0.430 2.800 0.450 ;
    END
  END GND
  PIN CommonNode
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 1.310 3.960 1.540 5.620 ;
    END
  END CommonNode
  PIN CommonMode
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 1.310 -0.430 1.540 1.020 ;
    END
  END CommonMode
  PIN output1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.670 4.260 2.960 4.420 ;
    END
  END output1
  PIN output2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.670 3.330 2.960 3.490 ;
    END
  END output2
  PIN output3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.670 1.490 2.960 1.650 ;
    END
  END output3
  PIN output4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.670 0.560 2.960 0.720 ;
    END
  END output4
  PIN input1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -11.120 4.020 -10.970 4.690 ;
    END
  END input1
  PIN input2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -11.120 3.520 -10.860 3.780 ;
    END
  END input2
  PIN input3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -11.180 0.980 -10.980 1.680 ;
    END
  END input3
  PIN input4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -11.190 0.470 -10.910 0.740 ;
    END
  END input4
  OBS
      LAYER li1 ;
        RECT -11.200 -0.380 2.940 5.290 ;
      LAYER met1 ;
        RECT -11.210 3.680 1.030 5.620 ;
        RECT 1.820 4.250 2.290 5.620 ;
        RECT 1.820 3.680 2.800 4.250 ;
        RECT -11.210 1.300 2.800 3.680 ;
        RECT -11.210 -0.430 1.030 1.300 ;
        RECT 1.820 0.730 2.800 1.300 ;
        RECT 1.820 -0.430 2.290 0.730 ;
      LAYER met2 ;
        RECT -11.210 4.970 0.690 5.340 ;
        RECT -10.690 4.700 0.690 4.970 ;
        RECT -10.690 4.060 0.390 4.700 ;
        RECT -10.580 3.980 0.390 4.060 ;
        RECT -10.580 3.770 0.690 3.980 ;
        RECT -10.580 3.240 0.390 3.770 ;
        RECT -11.210 3.050 0.390 3.240 ;
        RECT -11.210 1.960 0.690 3.050 ;
        RECT -10.700 1.930 0.690 1.960 ;
        RECT -10.700 1.210 0.390 1.930 ;
        RECT -10.700 1.020 0.690 1.210 ;
        RECT -10.630 1.000 0.690 1.020 ;
        RECT -10.630 0.280 0.390 1.000 ;
        RECT -10.630 0.190 0.690 0.280 ;
        RECT -11.210 -0.410 0.690 0.190 ;
  END
END sky130_hilas_WTA4Stage01
END LIBRARY

