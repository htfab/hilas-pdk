magic
tech sky130A
timestamp 1628616757
<< checkpaint >>
rect -337 1270 957 1271
rect -446 1235 957 1270
rect -624 1172 957 1235
rect -624 1001 958 1172
rect -624 -115 970 1001
rect -623 -562 970 -115
rect -623 -617 840 -562
<< nwell >>
rect 210 132 264 309
rect 204 105 264 132
rect 210 63 264 105
rect 192 18 264 63
rect 7 0 264 18
<< psubdiff >>
rect 206 518 250 525
rect 206 501 221 518
rect 238 501 250 518
rect 206 494 250 501
<< nsubdiff >>
rect 204 127 246 132
rect 204 110 216 127
rect 233 110 246 127
rect 204 105 246 110
<< psubdiffcont >>
rect 221 501 238 518
<< nsubdiffcont >>
rect 216 110 233 127
<< locali >>
rect 33 512 54 537
rect 220 526 237 531
rect 219 523 237 526
rect 219 518 262 523
rect 219 501 221 518
rect 238 501 262 518
rect 219 498 262 501
rect 219 495 238 498
rect 220 492 238 495
rect 208 110 216 127
rect 233 110 241 127
<< metal1 >>
rect 218 127 240 588
rect 216 110 240 127
rect 218 0 240 110
rect 258 0 280 588
<< metal2 >>
rect 0 571 7 575
rect 0 548 14 571
rect 198 549 280 566
rect 0 507 16 524
rect 0 456 14 473
rect 198 457 280 474
rect 0 415 17 432
rect 0 378 14 381
rect 0 364 21 378
rect 198 365 280 382
rect 0 323 16 340
rect 0 262 14 281
rect 200 255 280 275
rect 0 220 14 239
rect 0 183 14 185
rect 0 166 7 183
rect 200 159 280 179
rect 0 141 14 143
rect 0 124 7 141
rect 0 84 14 89
rect 0 70 7 84
rect 199 63 280 83
rect 0 45 14 47
rect 0 28 15 45
use sky130_hilas_pFETdevice01e  sky130_hilas_pFETdevice01e_2
timestamp 1628616734
transform 1 0 128 0 1 68
box 0 0 212 105
use sky130_hilas_pFETdevice01e  sky130_hilas_pFETdevice01e_1
timestamp 1628616734
transform 1 0 128 0 1 167
box 0 0 212 105
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1628616665
transform 0 1 221 -1 0 120
box 0 0 23 29
use sky130_hilas_pFETdevice01e  sky130_hilas_pFETdevice01e_0
timestamp 1628616734
transform 1 0 128 0 1 266
box 0 0 212 105
use sky130_hilas_nFET03a  sky130_hilas_nFET03a_0
timestamp 1628616711
transform 1 0 118 0 1 358
box 0 0 210 90
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1628616688
transform 1 0 26 0 1 325
box 0 0 34 33
use sky130_hilas_nFET03a  sky130_hilas_nFET03a_1
timestamp 1628616711
transform 1 0 118 0 1 457
box 0 0 210 90
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628616688
transform 1 0 28 0 1 424
box 0 0 34 33
use sky130_hilas_nFET03a  sky130_hilas_nFET03a_3
timestamp 1628616711
transform 1 0 117 0 1 556
box 0 0 210 90
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628616688
transform 1 0 30 0 1 516
box 0 0 34 33
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1628616665
transform 1 0 267 0 1 504
box 0 0 23 29
<< labels >>
rlabel metal1 218 0 240 9 0 WELL
port 13 nsew power default
rlabel metal1 258 0 280 9 0 VGND
port 14 nsew ground default
rlabel metal1 218 579 240 588 0 WELL
port 13 nsew ground default
rlabel metal1 258 579 280 588 0 VGND
port 14 nsew power default
rlabel metal2 0 548 7 565 0 NFET_SOURCE1
port 1 nsew analog default
rlabel metal2 0 507 7 524 0 NFET_GATE1
port 2 nsew analog default
rlabel metal2 0 456 7 473 0 NFET_SOURCE2
port 3 nsew analog default
rlabel metal2 0 415 7 432 0 NFET_GATE2
port 4 nsew analog default
rlabel metal2 0 364 7 381 0 NFET_SOURCE3
port 5 nsew analog default
rlabel metal2 0 323 7 340 0 NFET_GATE3
port 6 nsew analog default
rlabel metal2 0 220 7 239 0 PFET_GATE1
port 8 nsew analog default
rlabel metal2 0 262 7 281 0 PFET_SOURCE1
port 7 nsew analog default
rlabel metal2 0 166 7 185 0 PFET_SOURCE2
port 9 nsew analog default
rlabel metal2 0 124 7 143 0 PFET_GATE2
port 10 nsew analog default
rlabel metal2 0 70 7 89 0 PFET_SOURCE3
port 11 nsew analog default
rlabel metal2 0 28 7 47 0 PFET_GATE3
port 12 nsew analog default
rlabel metal2 274 255 280 275 0 PFET_DRAIN1
port 17 nsew analog default
rlabel metal2 274 159 280 179 0 PFET_DRAIN2
port 16 nsew analog default
rlabel metal2 274 63 280 83 0 PFET_DRAIN3
port 15 nsew analog default
rlabel metal2 275 549 280 566 0 NFET_DRAIN1
port 20 nsew analog default
rlabel metal2 275 457 280 474 0 NFET_DRAIN2
port 19 nsew analog default
rlabel metal2 275 365 280 382 0 NFET_DRAIN3
port 18 nsew analog default
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
