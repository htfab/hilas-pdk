magic
tech sky130A
magscale 1 2
timestamp 1627063414
<< error_s >>
rect 134 1906 234 1928
rect 278 1906 378 1928
rect 4702 1906 4802 1928
rect 4846 1906 4946 1928
rect 378 1844 442 1845
rect 4638 1844 4702 1845
rect 134 1822 234 1844
rect 278 1822 378 1844
rect 4702 1822 4802 1844
rect 4846 1822 4946 1844
rect 278 1782 378 1806
rect 4702 1782 4802 1806
rect 216 1722 223 1782
rect 378 1781 436 1782
rect 4644 1781 4702 1782
rect 4857 1722 4864 1782
rect 278 1698 378 1722
rect 4702 1698 4802 1722
rect 628 1690 662 1694
rect 1416 1692 1450 1696
rect 3630 1692 3664 1696
rect 4418 1690 4452 1694
rect 628 1652 662 1656
rect 1416 1654 1450 1658
rect 3630 1654 3664 1658
rect 4418 1652 4452 1656
rect 278 1618 378 1642
rect 4702 1618 4802 1642
rect 216 1558 223 1618
rect 378 1558 436 1559
rect 4644 1558 4702 1559
rect 4857 1558 4864 1618
rect 278 1534 378 1558
rect 4702 1534 4802 1558
rect 134 1496 234 1518
rect 278 1496 378 1518
rect 4702 1496 4802 1518
rect 4846 1496 4946 1518
rect 378 1495 442 1496
rect 4638 1495 4702 1496
rect 134 1412 234 1434
rect 278 1412 378 1434
rect 4702 1412 4802 1434
rect 4846 1412 4946 1434
rect 1414 1400 1448 1404
rect 3632 1400 3666 1404
rect 628 1372 662 1376
rect 4418 1372 4452 1376
rect 1414 1362 1448 1366
rect 3632 1362 3666 1366
rect 628 1334 662 1338
rect 4418 1334 4452 1338
rect 134 1304 234 1326
rect 278 1304 378 1326
rect 4702 1304 4802 1326
rect 4846 1304 4946 1326
rect 378 1242 442 1243
rect 4638 1242 4702 1243
rect 134 1220 234 1242
rect 278 1220 378 1242
rect 278 1180 378 1204
rect 216 1120 223 1180
rect 378 1179 436 1180
rect 654 1172 670 1238
rect 682 1200 720 1228
rect 762 1200 794 1228
rect 1122 1218 1136 1238
rect 1122 1164 1134 1218
rect 1150 1192 1198 1220
rect 1586 1190 1662 1218
rect 1944 1210 1984 1226
rect 2392 1184 2472 1212
rect 2608 1190 2688 1218
rect 3096 1210 3136 1228
rect 3418 1190 3494 1218
rect 3882 1196 3930 1224
rect 3944 1218 3958 1238
rect 2472 1156 2500 1182
rect 2580 1162 2608 1182
rect 3946 1168 3958 1218
rect 4286 1200 4318 1228
rect 4360 1200 4398 1228
rect 4410 1172 4426 1238
rect 4702 1220 4802 1242
rect 4846 1220 4946 1242
rect 4702 1180 4802 1204
rect 4644 1179 4702 1180
rect 4857 1120 4864 1180
rect 278 1096 378 1120
rect 528 1074 556 1112
rect 4534 1074 4562 1110
rect 4702 1096 4802 1120
rect 278 1018 378 1042
rect 216 958 223 1018
rect 4552 990 4562 1024
rect 4702 1018 4802 1042
rect 378 958 436 959
rect 4644 958 4702 959
rect 4857 958 4864 1018
rect 278 934 378 958
rect 4702 934 4802 958
rect 134 896 234 918
rect 278 896 378 918
rect 4702 896 4802 918
rect 4846 896 4946 918
rect 378 895 442 896
rect 4638 895 4702 896
rect 134 812 234 834
rect 278 812 378 834
rect 528 788 558 826
rect 4528 788 4556 824
rect 4702 812 4802 834
rect 4846 812 4946 834
rect 528 702 556 738
rect 4526 702 4554 738
rect 528 472 556 508
rect 4536 472 4564 508
rect 528 386 556 422
rect 4536 386 4564 422
rect 528 188 556 224
rect 4536 188 4564 224
rect 528 102 556 138
rect 4536 102 4564 138
rect 600 0 632 28
rect 682 2 720 30
rect 762 2 794 30
rect 1150 0 1198 28
rect 1586 0 1662 28
rect 1936 0 1984 28
rect 2392 0 2472 28
rect 2608 0 2688 28
rect 3096 0 3144 28
rect 3418 0 3494 30
rect 3882 0 3930 28
rect 4286 2 4318 30
rect 4360 2 4398 30
rect 4448 2 4480 30
<< metal1 >>
rect 600 1202 632 1210
rect 568 1198 632 1202
rect 682 1200 720 1210
rect 762 1200 794 1210
rect 568 1146 574 1198
rect 626 1146 632 1198
rect 1150 1192 1198 1210
rect 1586 1190 1662 1210
rect 1936 1198 1984 1210
rect 2392 1184 2472 1210
rect 2608 1190 2688 1210
rect 3096 1200 3144 1210
rect 3418 1190 3494 1210
rect 3882 1196 3930 1210
rect 4286 1200 4318 1210
rect 4360 1200 4398 1210
rect 4448 1202 4480 1210
rect 4448 1198 4512 1202
rect 568 1142 632 1146
rect 2472 1138 2608 1182
rect 4448 1146 4454 1198
rect 4506 1146 4512 1198
rect 4448 1142 4512 1146
rect 600 0 632 12
rect 682 2 720 14
rect 762 2 794 14
rect 1150 0 1198 16
rect 1586 0 1662 18
rect 1936 0 1984 14
rect 2392 0 2472 24
rect 2608 0 2688 24
rect 3096 0 3144 14
rect 3418 0 3494 30
rect 3882 0 3930 12
rect 4286 2 4318 14
rect 4360 2 4398 14
rect 4448 2 4480 14
<< via1 >>
rect 574 1146 626 1198
rect 4454 1146 4506 1198
<< metal2 >>
rect 568 1198 1138 1202
rect 568 1146 574 1198
rect 626 1182 1138 1198
rect 3946 1198 4512 1202
rect 3946 1182 4454 1198
rect 626 1166 4454 1182
rect 626 1146 652 1166
rect 1050 1146 3986 1166
rect 4448 1146 4454 1166
rect 4506 1146 4512 1198
rect 568 1142 652 1146
rect 4448 1142 4512 1146
rect 528 1074 556 1112
rect 4534 1074 4552 1110
rect 528 988 556 1026
rect 4534 988 4552 1024
rect 528 788 558 826
rect 4528 788 4554 824
rect 528 702 554 738
rect 4526 702 4554 738
rect 528 472 542 508
rect 4536 472 4554 508
rect 528 386 542 422
rect 4536 386 4554 422
rect 1868 276 3220 312
rect 528 188 542 224
rect 4536 188 4554 224
rect 528 102 542 138
rect 4536 102 4554 138
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_1
timestamp 1627063299
transform -1 0 2016 0 1 764
box 0 0 2016 1210
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_0
timestamp 1627063299
transform 1 0 3064 0 1 764
box 0 0 2016 1210
<< labels >>
rlabel metal1 3418 1190 3494 1210 0 GATE2
port 1 nsew analog default
rlabel metal1 2392 0 2472 24 0 VTUN
port 2 nsew power default
rlabel metal1 2608 0 2688 24 0 VTUN
port 2 nsew power default
rlabel metal1 2608 1190 2688 1210 0 VTUN
port 2 nsew power default
rlabel metal1 2392 1184 2472 1210 0 VTUN
port 2 nsew power default
rlabel metal1 1586 1190 1662 1210 0 GATE1
port 3 nsew analog default
rlabel metal1 1586 0 1662 18 0 GATE1
port 3 nsew analog default
rlabel metal1 4448 2 4480 14 0 VINJ
port 4 nsew power default
rlabel metal1 3418 0 3494 30 0 GATE2
port 1 nsew analog default
rlabel metal1 4360 1200 4398 1210 0 SelectGate2
rlabel metal1 4448 1200 4480 1210 0 VINJ
port 6 nsew power default
rlabel metal1 600 1200 632 1210 0 VINJ
port 6 nsew power default
rlabel metal1 682 1200 720 1210 0 GATESELECT1
port 10 nsew analog default
rlabel metal1 600 0 632 12 0 VINJ
port 6 nsew power default
rlabel metal1 682 2 720 14 0 GATESELECT1
port 10 nsew analog default
rlabel metal1 762 1200 794 1210 0 COL1
port 12 nsew analog default
rlabel metal1 762 2 794 14 0 COL1
port 12 nsew analog default
rlabel metal1 4360 2 4398 14 0 GATESELECT2
port 11 nsew analog default
rlabel metal1 4286 2 4318 14 0 COL2
port 13 nsew analog default
rlabel metal1 4286 1200 4318 1210 0 COL2
port 13 nsew analog default
rlabel metal2 528 988 542 1026 0 ROW1
port 14 nsew analog default
rlabel metal2 528 788 542 826 0 ROW2
port 15 nsew analog default
rlabel metal2 528 1074 542 1112 0 DRAIN1
port 16 nsew analog default
rlabel metal2 528 702 542 738 0 DRAIN2
port 17 nsew analog default
rlabel metal2 528 472 542 508 0 DRAIN3
port 18 nsew analog default
rlabel metal2 528 386 542 422 0 ROW3
port 19 nsew analog default
rlabel metal2 528 188 542 224 0 ROW4
port 20 nsew analog default
rlabel metal2 528 102 542 138 0 DRAIN4
port 21 nsew analog default
rlabel metal2 4534 1074 4552 1110 0 DRAIN1
port 16 nsew analog default
rlabel metal2 4534 988 4552 1024 0 ROW1
port 14 nsew analog default
rlabel metal2 4536 788 4554 824 0 ROW2
port 15 nsew
rlabel metal2 4536 702 4554 738 0 DRAIN2
port 17 nsew analog default
rlabel metal2 4536 472 4554 508 0 DRAIN3
port 18 nsew analog default
rlabel metal2 4536 386 4554 422 0 ROW3
port 19 nsew analog default
rlabel metal2 4536 188 4554 224 0 ROW4
port 20 nsew analog default
rlabel metal2 4536 102 4554 138 0 DRAIN4
port 21 nsew
rlabel metal1 1150 1198 1198 1210 0 VGND
port 22 nsew
rlabel metal1 1150 0 1198 16 0 VGND
port 22 nsew
rlabel metal1 1936 0 1984 14 0 VGND
port 22 nsew
rlabel metal1 1936 1198 1984 1210 0 VGND
port 22 nsew
rlabel metal1 3096 0 3144 14 0 VGND
port 22 nsew
rlabel metal1 3882 0 3930 12 0 VGND
port 22 nsew
rlabel metal1 3096 1200 3144 1210 0 VGND
port 22 nsew
rlabel metal1 3882 1196 3930 1210 0 VGND
port 22 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
