VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_pfetmirror02
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pfetmirror02 ;
  ORIGIN 0.610 -0.890 ;
  SIZE 1.280 BY 2.840 ;
  OBS
      LAYER nwell ;
        RECT -0.610 0.890 0.670 3.730 ;
      LAYER li1 ;
        RECT -0.410 3.310 0.290 3.490 ;
        RECT -0.400 2.010 0.300 2.890 ;
        RECT -0.400 1.400 0.310 1.570 ;
        RECT -0.050 1.120 0.310 1.400 ;
        RECT -0.050 0.950 0.280 1.120 ;
  END
END sky130_hilas_pfetmirror02
END LIBRARY

