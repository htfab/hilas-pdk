VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_hilas_invert01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_invert01 ;
  ORIGIN 0.130 0.150 ;
  SIZE 0.520 BY 0.310 ;
  OBS
      LAYER li1 ;
        RECT -0.040 0.050 0.000 0.090 ;
        RECT 0.270 0.060 0.310 0.100 ;
        RECT -0.040 -0.060 0.000 -0.020 ;
        RECT 0.270 -0.070 0.310 -0.030 ;
      LAYER met1 ;
        RECT 0.100 0.090 0.140 0.160 ;
        RECT 0.000 0.060 0.270 0.090 ;
        RECT 0.000 0.050 0.310 0.060 ;
        RECT -0.120 -0.060 -0.040 -0.020 ;
        RECT 0.310 -0.070 0.380 -0.030 ;
        RECT 0.100 -0.150 0.140 -0.080 ;
      LAYER via ;
        RECT 0.340 -0.070 0.380 -0.030 ;
      LAYER met2 ;
        RECT -0.130 -0.120 -0.070 0.150 ;
        RECT 0.330 -0.120 0.390 0.150 ;
  END
END sky130_hilas_invert01

MACRO sky130_hilas_CapModule02
  CLASS BLOCK ;
  FOREIGN sky130_hilas_CapModule02 ;
  ORIGIN 4.430 2.470 ;
  SIZE 7.200 BY 5.830 ;
  OBS
      LAYER met3 ;
        RECT -4.430 3.330 -1.610 3.360 ;
        RECT -4.430 -2.450 2.770 3.330 ;
        RECT -1.640 -2.470 2.770 -2.450 ;
      LAYER met4 ;
        RECT -3.540 -1.370 -0.500 -0.900 ;
  END
END sky130_hilas_CapModule02

MACRO sky130_hilas_poly2m1
  CLASS BLOCK ;
  FOREIGN sky130_hilas_poly2m1 ;
  ORIGIN 0.090 0.260 ;
  SIZE 0.330 BY 0.510 ;
  OBS
      LAYER li1 ;
        RECT -0.030 -0.180 0.180 0.250 ;
        RECT -0.010 -0.200 0.160 -0.180 ;
      LAYER met1 ;
        RECT -0.030 0.030 0.190 0.250 ;
        RECT -0.040 -0.260 0.190 0.030 ;
  END
END sky130_hilas_poly2m1

MACRO sky130_hilas_FGVaractorCapacitor02
  CLASS BLOCK ;
  FOREIGN sky130_hilas_FGVaractorCapacitor02 ;
  ORIGIN 10.050 3.800 ;
  SIZE 2.720 BY 1.690 ;
  OBS
      LAYER nwell ;
        RECT -10.050 -2.150 -7.340 -2.110 ;
        RECT -10.050 -3.800 -7.330 -2.150 ;
      LAYER li1 ;
        RECT -9.750 -3.280 -9.520 -2.590 ;
      LAYER mcon ;
        RECT -9.720 -2.800 -9.550 -2.630 ;
        RECT -9.720 -3.250 -9.550 -3.080 ;
      LAYER met1 ;
        RECT -9.770 -3.330 -9.510 -2.540 ;
  END
END sky130_hilas_FGVaractorCapacitor02

MACRO sky130_hilas_poly2m2
  CLASS BLOCK ;
  FOREIGN sky130_hilas_poly2m2 ;
  ORIGIN 0.090 0.260 ;
  SIZE 0.330 BY 0.550 ;
  OBS
      LAYER li1 ;
        RECT -0.030 -0.180 0.180 0.250 ;
        RECT -0.010 -0.200 0.160 -0.180 ;
      LAYER met1 ;
        RECT -0.080 -0.030 0.240 0.290 ;
        RECT -0.040 -0.260 0.190 -0.030 ;
      LAYER via ;
        RECT -0.050 0.000 0.210 0.260 ;
      LAYER met2 ;
        RECT -0.080 -0.030 0.240 0.290 ;
  END
END sky130_hilas_poly2m2

MACRO sky130_hilas_Trans4small
  CLASS BLOCK ;
  FOREIGN sky130_hilas_Trans4small ;
  ORIGIN -1.910 1.500 ;
  SIZE 2.800 BY 5.880 ;
  PIN NFET_SOURCE1
    USE ANALOG ;
    ANTENNADIFFAREA 0.108500 ;
    PORT
      LAYER li1 ;
        RECT 2.830 4.200 3.030 4.240 ;
        RECT 2.520 3.940 3.030 4.200 ;
        RECT 2.830 3.910 3.030 3.940 ;
      LAYER mcon ;
        RECT 2.580 3.980 2.750 4.150 ;
      LAYER met1 ;
        RECT 2.510 3.910 2.830 4.230 ;
      LAYER via ;
        RECT 2.540 3.940 2.800 4.200 ;
      LAYER met2 ;
        RECT 2.510 4.150 2.820 4.240 ;
        RECT 1.910 3.980 2.820 4.150 ;
        RECT 2.510 3.910 2.820 3.980 ;
    END
  END NFET_SOURCE1
  PIN NFET_GATE1
    USE ANALOG ;
    ANTENNAGATEAREA 0.094500 ;
    PORT
      LAYER li1 ;
        RECT 2.080 3.740 2.510 3.760 ;
        RECT 2.080 3.570 2.530 3.740 ;
        RECT 2.080 3.550 2.510 3.570 ;
      LAYER mcon ;
        RECT 2.360 3.570 2.530 3.740 ;
      LAYER met1 ;
        RECT 2.040 3.770 2.360 3.820 ;
        RECT 2.040 3.540 2.590 3.770 ;
        RECT 2.040 3.500 2.360 3.540 ;
      LAYER via ;
        RECT 2.070 3.530 2.330 3.790 ;
      LAYER met2 ;
        RECT 2.040 3.740 2.360 3.820 ;
        RECT 1.910 3.570 2.360 3.740 ;
        RECT 2.040 3.500 2.360 3.570 ;
    END
  END NFET_GATE1
  PIN NFET_SOURCE2
    USE ANALOG ;
    ANTENNADIFFAREA 0.108500 ;
    PORT
      LAYER li1 ;
        RECT 2.830 3.280 3.030 3.320 ;
        RECT 2.520 3.020 3.030 3.280 ;
        RECT 2.830 2.990 3.030 3.020 ;
      LAYER mcon ;
        RECT 2.580 3.060 2.750 3.230 ;
      LAYER met1 ;
        RECT 2.510 2.990 2.830 3.310 ;
      LAYER via ;
        RECT 2.540 3.020 2.800 3.280 ;
      LAYER met2 ;
        RECT 2.510 3.230 2.820 3.320 ;
        RECT 1.910 3.060 2.820 3.230 ;
        RECT 2.510 2.990 2.820 3.060 ;
    END
  END NFET_SOURCE2
  PIN NFET_GATE2
    USE ANALOG ;
    ANTENNAGATEAREA 0.094500 ;
    PORT
      LAYER li1 ;
        RECT 2.080 2.820 2.510 2.840 ;
        RECT 2.080 2.650 2.530 2.820 ;
        RECT 2.080 2.630 2.510 2.650 ;
      LAYER mcon ;
        RECT 2.360 2.650 2.530 2.820 ;
      LAYER met1 ;
        RECT 2.040 2.850 2.360 2.900 ;
        RECT 2.040 2.620 2.590 2.850 ;
        RECT 2.040 2.580 2.360 2.620 ;
      LAYER via ;
        RECT 2.070 2.610 2.330 2.870 ;
      LAYER met2 ;
        RECT 2.040 2.820 2.360 2.900 ;
        RECT 1.910 2.650 2.360 2.820 ;
        RECT 2.040 2.580 2.360 2.650 ;
    END
  END NFET_GATE2
  PIN NFET_SOURCE3
    USE ANALOG ;
    ANTENNADIFFAREA 0.108500 ;
    PORT
      LAYER li1 ;
        RECT 2.830 2.360 3.030 2.400 ;
        RECT 2.520 2.100 3.030 2.360 ;
        RECT 2.830 2.070 3.030 2.100 ;
      LAYER mcon ;
        RECT 2.580 2.140 2.750 2.310 ;
      LAYER met1 ;
        RECT 2.510 2.070 2.830 2.390 ;
      LAYER via ;
        RECT 2.540 2.100 2.800 2.360 ;
      LAYER met2 ;
        RECT 2.510 2.310 2.820 2.400 ;
        RECT 1.910 2.140 2.820 2.310 ;
        RECT 2.510 2.070 2.820 2.140 ;
    END
  END NFET_SOURCE3
  PIN NFET_GATE3
    USE ANALOG ;
    ANTENNAGATEAREA 0.094500 ;
    PORT
      LAYER li1 ;
        RECT 2.080 1.900 2.510 1.920 ;
        RECT 2.080 1.730 2.530 1.900 ;
        RECT 2.080 1.710 2.510 1.730 ;
      LAYER mcon ;
        RECT 2.360 1.730 2.530 1.900 ;
      LAYER met1 ;
        RECT 2.040 1.930 2.360 1.980 ;
        RECT 2.040 1.700 2.590 1.930 ;
        RECT 2.040 1.660 2.360 1.700 ;
      LAYER via ;
        RECT 2.070 1.690 2.330 1.950 ;
      LAYER met2 ;
        RECT 2.040 1.900 2.360 1.980 ;
        RECT 1.910 1.730 2.360 1.900 ;
        RECT 2.040 1.660 2.360 1.730 ;
    END
  END NFET_GATE3
  PIN PFET_SOURCE1
    USE ANALOG ;
    ANTENNADIFFAREA 0.109200 ;
    PORT
      LAYER li1 ;
        RECT 2.330 1.340 2.650 1.380 ;
        RECT 2.330 1.320 2.660 1.340 ;
        RECT 2.330 1.120 2.950 1.320 ;
        RECT 2.780 0.990 2.950 1.120 ;
      LAYER mcon ;
        RECT 2.390 1.160 2.560 1.330 ;
      LAYER met1 ;
        RECT 2.320 1.090 2.640 1.410 ;
      LAYER via ;
        RECT 2.350 1.120 2.610 1.380 ;
      LAYER met2 ;
        RECT 2.320 1.310 2.630 1.420 ;
        RECT 1.910 1.120 2.630 1.310 ;
        RECT 2.320 1.090 2.630 1.120 ;
    END
  END PFET_SOURCE1
  PIN PFET_GATE1
    USE ANALOG ;
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER li1 ;
        RECT 2.170 0.880 2.600 0.900 ;
        RECT 2.150 0.710 2.600 0.880 ;
        RECT 2.170 0.690 2.600 0.710 ;
      LAYER met1 ;
        RECT 2.320 0.910 2.640 0.950 ;
        RECT 2.090 0.680 2.640 0.910 ;
        RECT 2.320 0.630 2.640 0.680 ;
      LAYER via ;
        RECT 2.350 0.660 2.610 0.920 ;
      LAYER met2 ;
        RECT 2.320 0.890 2.640 0.950 ;
        RECT 1.910 0.700 2.640 0.890 ;
        RECT 2.320 0.630 2.640 0.700 ;
    END
  END PFET_GATE1
  PIN PFET_SOURCE2
    USE ANALOG ;
    ANTENNADIFFAREA 0.109200 ;
    PORT
      LAYER li1 ;
        RECT 2.330 0.380 2.650 0.420 ;
        RECT 2.330 0.360 2.660 0.380 ;
        RECT 2.330 0.160 2.950 0.360 ;
        RECT 2.780 0.030 2.950 0.160 ;
      LAYER mcon ;
        RECT 2.390 0.200 2.560 0.370 ;
      LAYER met1 ;
        RECT 2.320 0.130 2.640 0.450 ;
      LAYER via ;
        RECT 2.350 0.160 2.610 0.420 ;
      LAYER met2 ;
        RECT 2.320 0.350 2.630 0.460 ;
        RECT 1.910 0.160 2.630 0.350 ;
        RECT 2.320 0.130 2.630 0.160 ;
    END
  END PFET_SOURCE2
  PIN PFET_GATE2
    USE ANALOG ;
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER li1 ;
        RECT 2.170 -0.080 2.600 -0.060 ;
        RECT 2.150 -0.250 2.600 -0.080 ;
        RECT 2.170 -0.270 2.600 -0.250 ;
      LAYER met1 ;
        RECT 2.320 -0.050 2.640 -0.010 ;
        RECT 2.090 -0.280 2.640 -0.050 ;
        RECT 2.320 -0.330 2.640 -0.280 ;
      LAYER via ;
        RECT 2.350 -0.300 2.610 -0.040 ;
      LAYER met2 ;
        RECT 2.320 -0.070 2.640 -0.010 ;
        RECT 1.910 -0.260 2.640 -0.070 ;
        RECT 2.320 -0.330 2.640 -0.260 ;
    END
  END PFET_GATE2
  PIN PFET_SOURCE3
    USE ANALOG ;
    ANTENNADIFFAREA 0.109200 ;
    PORT
      LAYER li1 ;
        RECT 2.330 -0.580 2.650 -0.540 ;
        RECT 2.330 -0.600 2.660 -0.580 ;
        RECT 2.330 -0.800 2.950 -0.600 ;
        RECT 2.780 -0.930 2.950 -0.800 ;
      LAYER mcon ;
        RECT 2.390 -0.760 2.560 -0.590 ;
      LAYER met1 ;
        RECT 2.320 -0.830 2.640 -0.510 ;
      LAYER via ;
        RECT 2.350 -0.800 2.610 -0.540 ;
      LAYER met2 ;
        RECT 2.320 -0.610 2.630 -0.500 ;
        RECT 1.910 -0.800 2.630 -0.610 ;
        RECT 2.320 -0.830 2.630 -0.800 ;
    END
  END PFET_SOURCE3
  PIN PFET_GATE3
    USE ANALOG ;
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER li1 ;
        RECT 2.170 -1.040 2.600 -1.020 ;
        RECT 2.150 -1.210 2.600 -1.040 ;
        RECT 2.170 -1.230 2.600 -1.210 ;
      LAYER met1 ;
        RECT 2.320 -1.010 2.640 -0.970 ;
        RECT 2.090 -1.240 2.640 -1.010 ;
        RECT 2.320 -1.290 2.640 -1.240 ;
      LAYER via ;
        RECT 2.350 -1.260 2.610 -1.000 ;
      LAYER met2 ;
        RECT 2.320 -1.030 2.640 -0.970 ;
        RECT 1.910 -1.220 2.640 -1.030 ;
        RECT 2.320 -1.290 2.640 -1.220 ;
    END
  END PFET_GATE3
  PIN WELL
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 1.980 -1.500 4.550 1.590 ;
      LAYER li1 ;
        RECT 3.960 -1.270 4.380 -1.100 ;
        RECT 4.060 -1.310 4.290 -1.270 ;
      LAYER mcon ;
        RECT 4.090 -1.300 4.260 -1.130 ;
      LAYER met1 ;
        RECT 4.090 -1.100 4.310 4.380 ;
        RECT 4.030 -1.330 4.320 -1.100 ;
        RECT 4.090 -1.500 4.310 -1.330 ;
    END
  END WELL
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 4.110 3.760 4.280 3.810 ;
        RECT 4.100 3.730 4.280 3.760 ;
        RECT 4.100 3.720 4.530 3.730 ;
        RECT 4.100 3.490 4.690 3.720 ;
        RECT 4.100 3.480 4.530 3.490 ;
        RECT 4.100 3.420 4.270 3.480 ;
      LAYER mcon ;
        RECT 4.510 3.520 4.680 3.690 ;
      LAYER met1 ;
        RECT 4.490 3.750 4.710 4.380 ;
        RECT 4.480 3.460 4.710 3.750 ;
        RECT 4.490 -1.500 4.710 3.460 ;
    END
  END VGND
  PIN PFET_DRAIN3
    USE ANALOG ;
    ANTENNADIFFAREA 0.105300 ;
    PORT
      LAYER li1 ;
        RECT 3.460 -0.640 3.630 -0.600 ;
        RECT 3.460 -0.680 3.950 -0.640 ;
        RECT 3.460 -0.870 3.960 -0.680 ;
        RECT 3.460 -0.900 3.950 -0.870 ;
        RECT 3.460 -0.930 3.630 -0.900 ;
      LAYER mcon ;
        RECT 3.690 -0.860 3.860 -0.690 ;
      LAYER met1 ;
        RECT 3.620 -0.930 3.940 -0.610 ;
      LAYER via ;
        RECT 3.650 -0.900 3.910 -0.640 ;
      LAYER met2 ;
        RECT 3.620 -0.670 3.930 -0.600 ;
        RECT 3.620 -0.870 4.710 -0.670 ;
        RECT 3.620 -0.930 3.930 -0.870 ;
    END
  END PFET_DRAIN3
  PIN PFET_DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.105300 ;
    PORT
      LAYER li1 ;
        RECT 3.460 0.320 3.630 0.360 ;
        RECT 3.460 0.280 3.950 0.320 ;
        RECT 3.460 0.090 3.960 0.280 ;
        RECT 3.460 0.060 3.950 0.090 ;
        RECT 3.460 0.030 3.630 0.060 ;
      LAYER mcon ;
        RECT 3.690 0.100 3.860 0.270 ;
      LAYER met1 ;
        RECT 3.620 0.030 3.940 0.350 ;
      LAYER via ;
        RECT 3.650 0.060 3.910 0.320 ;
      LAYER met2 ;
        RECT 3.620 0.290 3.930 0.360 ;
        RECT 3.620 0.090 4.710 0.290 ;
        RECT 3.620 0.030 3.930 0.090 ;
    END
  END PFET_DRAIN2
  PIN PFET_DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.105300 ;
    PORT
      LAYER li1 ;
        RECT 3.460 1.280 3.630 1.320 ;
        RECT 3.460 1.240 3.950 1.280 ;
        RECT 3.460 1.050 3.960 1.240 ;
        RECT 3.460 1.020 3.950 1.050 ;
        RECT 3.460 0.990 3.630 1.020 ;
      LAYER mcon ;
        RECT 3.690 1.060 3.860 1.230 ;
      LAYER met1 ;
        RECT 3.620 0.990 3.940 1.310 ;
      LAYER via ;
        RECT 3.650 1.020 3.910 1.280 ;
      LAYER met2 ;
        RECT 3.620 1.250 3.930 1.320 ;
        RECT 3.620 1.050 4.710 1.250 ;
        RECT 3.620 0.990 3.930 1.050 ;
    END
  END PFET_DRAIN1
  PIN NFET_DRAIN3
    USE ANALOG ;
    ANTENNADIFFAREA 0.108500 ;
    PORT
      LAYER li1 ;
        RECT 3.420 2.370 3.620 2.400 ;
        RECT 3.420 2.330 3.930 2.370 ;
        RECT 3.420 2.140 3.940 2.330 ;
        RECT 3.420 2.110 3.930 2.140 ;
        RECT 3.420 2.070 3.620 2.110 ;
      LAYER mcon ;
        RECT 3.670 2.150 3.840 2.320 ;
      LAYER met1 ;
        RECT 3.600 2.080 3.920 2.400 ;
      LAYER via ;
        RECT 3.630 2.110 3.890 2.370 ;
      LAYER met2 ;
        RECT 3.600 2.320 3.910 2.410 ;
        RECT 3.600 2.150 4.710 2.320 ;
        RECT 3.600 2.080 3.910 2.150 ;
    END
  END NFET_DRAIN3
  PIN NFET_DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.108500 ;
    PORT
      LAYER li1 ;
        RECT 3.420 3.290 3.620 3.320 ;
        RECT 3.420 3.250 3.930 3.290 ;
        RECT 3.420 3.060 3.940 3.250 ;
        RECT 3.420 3.030 3.930 3.060 ;
        RECT 3.420 2.990 3.620 3.030 ;
      LAYER mcon ;
        RECT 3.670 3.070 3.840 3.240 ;
      LAYER met1 ;
        RECT 3.600 3.000 3.920 3.320 ;
      LAYER via ;
        RECT 3.630 3.030 3.890 3.290 ;
      LAYER met2 ;
        RECT 3.600 3.240 3.910 3.330 ;
        RECT 3.600 3.070 4.710 3.240 ;
        RECT 3.600 3.000 3.910 3.070 ;
    END
  END NFET_DRAIN2
  PIN NFET_DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.108500 ;
    PORT
      LAYER li1 ;
        RECT 3.420 4.210 3.620 4.240 ;
        RECT 3.420 4.170 3.930 4.210 ;
        RECT 3.420 3.980 3.940 4.170 ;
        RECT 3.420 3.950 3.930 3.980 ;
        RECT 3.420 3.910 3.620 3.950 ;
      LAYER mcon ;
        RECT 3.670 3.990 3.840 4.160 ;
      LAYER met1 ;
        RECT 3.600 3.920 3.920 4.240 ;
      LAYER via ;
        RECT 3.630 3.950 3.890 4.210 ;
      LAYER met2 ;
        RECT 3.600 4.160 3.910 4.250 ;
        RECT 3.600 3.990 4.710 4.160 ;
        RECT 3.600 3.920 3.910 3.990 ;
    END
  END NFET_DRAIN1
END sky130_hilas_Trans4small

MACRO sky130_hilas_horizPcell01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_horizPcell01 ;
  ORIGIN 2.890 -0.470 ;
  SIZE 2.560 BY 1.850 ;
  OBS
      LAYER nwell ;
        RECT -2.890 0.480 -0.330 2.320 ;
        RECT -2.890 0.470 -0.340 0.480 ;
      LAYER li1 ;
        RECT -2.790 1.670 -2.470 1.680 ;
        RECT -2.790 1.500 -2.210 1.670 ;
        RECT -2.790 1.460 -2.460 1.500 ;
        RECT -2.790 1.420 -2.470 1.460 ;
        RECT -1.660 1.170 -1.460 1.740 ;
        RECT -0.940 1.180 -0.720 1.770 ;
        RECT -0.930 1.150 -0.720 1.180 ;
        RECT -2.790 1.100 -2.470 1.130 ;
        RECT -2.790 1.050 -2.460 1.100 ;
        RECT -2.790 0.880 -2.210 1.050 ;
        RECT -2.790 0.870 -2.470 0.880 ;
        RECT -0.930 0.800 -0.730 1.150 ;
      LAYER mcon ;
        RECT -2.730 1.470 -2.560 1.640 ;
        RECT -1.650 1.210 -1.480 1.380 ;
        RECT -0.920 1.180 -0.750 1.350 ;
        RECT -2.730 0.920 -2.560 1.090 ;
      LAYER met1 ;
        RECT -2.800 1.390 -2.480 1.710 ;
        RECT -1.660 1.630 -1.500 2.320 ;
        RECT -1.660 1.410 -1.460 1.630 ;
        RECT -1.260 1.580 -1.100 2.320 ;
        RECT -0.850 1.810 -0.690 2.320 ;
        RECT -0.850 1.720 -0.680 1.810 ;
        RECT -1.270 1.460 -1.100 1.580 ;
        RECT -1.680 1.170 -1.450 1.410 ;
        RECT -2.800 0.840 -2.480 1.160 ;
        RECT -1.660 1.150 -1.460 1.170 ;
        RECT -1.660 0.470 -1.500 1.150 ;
        RECT -1.290 0.470 -1.100 1.460 ;
        RECT -0.960 1.670 -0.680 1.720 ;
        RECT -0.960 1.120 -0.690 1.670 ;
        RECT -0.850 0.470 -0.690 1.120 ;
      LAYER via ;
        RECT -2.770 1.420 -2.510 1.680 ;
        RECT -2.770 0.870 -2.510 1.130 ;
      LAYER met2 ;
        RECT -2.800 1.580 -2.490 1.710 ;
        RECT -2.890 1.400 -0.330 1.580 ;
        RECT -2.800 1.380 -2.490 1.400 ;
        RECT -2.800 1.150 -2.490 1.160 ;
        RECT -2.800 0.970 -0.330 1.150 ;
        RECT -2.800 0.830 -2.490 0.970 ;
  END
END sky130_hilas_horizPcell01

MACRO sky130_hilas_Trans2med
  CLASS BLOCK ;
  FOREIGN sky130_hilas_Trans2med ;
  ORIGIN 3.800 1.430 ;
  SIZE 3.530 BY 5.950 ;
  PIN NFET_GATE01
    USE ANALOG ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER li1 ;
        RECT -3.530 0.960 -3.320 1.390 ;
        RECT -3.510 0.940 -3.340 0.960 ;
      LAYER met1 ;
        RECT -3.540 1.170 -3.320 1.390 ;
        RECT -3.540 0.880 -3.310 1.170 ;
        RECT -3.550 0.560 -3.290 0.880 ;
      LAYER via ;
        RECT -3.550 0.590 -3.290 0.850 ;
      LAYER met2 ;
        RECT -3.580 0.830 -3.260 0.850 ;
        RECT -3.800 0.610 -3.260 0.830 ;
        RECT -3.580 0.590 -3.260 0.610 ;
    END
  END NFET_GATE01
  PIN PET_GATE02
    USE ANALOG ;
    ANTENNAGATEAREA 0.652600 ;
    PORT
      LAYER li1 ;
        RECT -0.780 1.850 -0.350 1.870 ;
        RECT -0.780 1.680 -0.330 1.850 ;
        RECT -0.780 1.660 -0.350 1.680 ;
      LAYER mcon ;
        RECT -0.500 1.680 -0.330 1.850 ;
      LAYER met1 ;
        RECT -0.820 1.880 -0.500 1.930 ;
        RECT -0.820 1.650 -0.270 1.880 ;
        RECT -0.820 1.610 -0.500 1.650 ;
      LAYER via ;
        RECT -0.790 1.640 -0.530 1.900 ;
      LAYER met2 ;
        RECT -0.820 1.800 -0.500 1.930 ;
        RECT -3.800 1.610 -0.500 1.800 ;
        RECT -3.800 1.590 -0.820 1.610 ;
    END
  END PET_GATE02
  PIN PFET_GATE01
    USE ANALOG ;
    ANTENNAGATEAREA 0.652600 ;
    PORT
      LAYER li1 ;
        RECT -3.500 2.030 -3.330 2.050 ;
        RECT -3.520 1.600 -3.310 2.030 ;
      LAYER mcon ;
        RECT -3.500 1.880 -3.330 2.050 ;
      LAYER met1 ;
        RECT -3.550 2.110 -3.290 2.430 ;
        RECT -3.530 1.820 -3.300 2.110 ;
        RECT -3.520 1.600 -3.300 1.820 ;
      LAYER via ;
        RECT -3.550 2.140 -3.290 2.400 ;
      LAYER met2 ;
        RECT -3.580 2.370 -3.260 2.400 ;
        RECT -3.800 2.150 -3.260 2.370 ;
        RECT -3.580 2.140 -3.260 2.150 ;
    END
  END PFET_GATE01
  PIN NFET_GATE02
    USE ANALOG ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER li1 ;
        RECT -0.790 1.310 -0.360 1.330 ;
        RECT -0.790 1.140 -0.340 1.310 ;
        RECT -0.790 1.120 -0.360 1.140 ;
      LAYER mcon ;
        RECT -0.510 1.140 -0.340 1.310 ;
      LAYER met1 ;
        RECT -0.830 1.340 -0.510 1.390 ;
        RECT -0.830 1.110 -0.280 1.340 ;
        RECT -0.830 1.070 -0.510 1.110 ;
      LAYER via ;
        RECT -0.800 1.100 -0.540 1.360 ;
      LAYER met2 ;
        RECT -3.800 1.390 -0.820 1.400 ;
        RECT -3.800 1.190 -0.510 1.390 ;
        RECT -0.830 1.070 -0.510 1.190 ;
    END
  END NFET_GATE02
  PIN PFET_SOURCE1
    USE ANALOG ;
    ANTENNADIFFAREA 0.727900 ;
    PORT
      LAYER li1 ;
        RECT -2.960 3.380 -2.790 4.290 ;
        RECT -3.090 3.340 -2.770 3.380 ;
        RECT -3.090 3.150 -2.760 3.340 ;
        RECT -3.090 3.120 -2.770 3.150 ;
        RECT -2.960 1.800 -2.790 3.120 ;
      LAYER mcon ;
        RECT -3.030 3.160 -2.860 3.330 ;
      LAYER met1 ;
        RECT -3.100 3.090 -2.780 3.410 ;
      LAYER via ;
        RECT -3.070 3.120 -2.810 3.380 ;
      LAYER met2 ;
        RECT -3.100 3.360 -2.790 3.420 ;
        RECT -3.800 3.150 -2.790 3.360 ;
        RECT -3.800 3.140 -3.530 3.150 ;
        RECT -3.100 3.090 -2.790 3.150 ;
    END
  END PFET_SOURCE1
  PIN PFET_SOURCE2
    USE ANALOG ;
    ANTENNADIFFAREA 0.727900 ;
    PORT
      LAYER li1 ;
        RECT -1.780 4.160 -1.610 4.290 ;
        RECT -1.920 4.120 -1.600 4.160 ;
        RECT -1.920 3.930 -1.590 4.120 ;
        RECT -1.920 3.900 -1.600 3.930 ;
        RECT -1.780 1.800 -1.610 3.900 ;
      LAYER mcon ;
        RECT -1.860 3.940 -1.690 4.110 ;
      LAYER met1 ;
        RECT -1.930 3.870 -1.610 4.190 ;
      LAYER via ;
        RECT -1.900 3.900 -1.640 4.160 ;
      LAYER met2 ;
        RECT -1.930 4.140 -1.620 4.200 ;
        RECT -3.800 3.920 -1.620 4.140 ;
        RECT -1.930 3.870 -1.620 3.920 ;
    END
  END PFET_SOURCE2
  PIN NFET_SOURCE2
    USE ANALOG ;
    ANTENNADIFFAREA 0.688800 ;
    PORT
      LAYER li1 ;
        RECT -1.780 -0.940 -1.610 1.150 ;
        RECT -1.900 -0.980 -1.580 -0.940 ;
        RECT -1.900 -1.170 -1.570 -0.980 ;
        RECT -1.900 -1.200 -1.580 -1.170 ;
        RECT -1.780 -1.250 -1.610 -1.200 ;
      LAYER mcon ;
        RECT -1.840 -1.160 -1.670 -0.990 ;
      LAYER met1 ;
        RECT -1.910 -1.230 -1.590 -0.910 ;
      LAYER via ;
        RECT -1.880 -1.200 -1.620 -0.940 ;
      LAYER met2 ;
        RECT -1.910 -0.970 -1.600 -0.900 ;
        RECT -3.800 -1.190 -1.600 -0.970 ;
        RECT -1.910 -1.230 -1.600 -1.190 ;
    END
  END NFET_SOURCE2
  PIN NFET_SOURCE1
    USE ANALOG ;
    ANTENNADIFFAREA 0.688800 ;
    PORT
      LAYER li1 ;
        RECT -2.970 -0.500 -2.800 1.150 ;
        RECT -3.120 -0.540 -2.800 -0.500 ;
        RECT -3.120 -0.730 -2.790 -0.540 ;
        RECT -3.120 -0.760 -2.800 -0.730 ;
        RECT -2.970 -1.250 -2.800 -0.760 ;
      LAYER mcon ;
        RECT -3.060 -0.720 -2.890 -0.550 ;
      LAYER met1 ;
        RECT -3.130 -0.790 -2.810 -0.470 ;
      LAYER via ;
        RECT -3.100 -0.760 -2.840 -0.500 ;
      LAYER met2 ;
        RECT -3.130 -0.530 -2.820 -0.460 ;
        RECT -3.800 -0.740 -2.820 -0.530 ;
        RECT -3.130 -0.790 -2.820 -0.740 ;
    END
  END NFET_SOURCE1
  PIN NFET_DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.688800 ;
    PORT
      LAYER li1 ;
        RECT -2.420 -0.500 -2.250 1.150 ;
        RECT -2.420 -0.540 -2.100 -0.500 ;
        RECT -2.420 -0.730 -2.090 -0.540 ;
        RECT -2.420 -0.760 -2.100 -0.730 ;
        RECT -2.420 -1.250 -2.250 -0.760 ;
      LAYER mcon ;
        RECT -2.360 -0.720 -2.190 -0.550 ;
      LAYER met1 ;
        RECT -2.430 -0.790 -2.110 -0.470 ;
      LAYER via ;
        RECT -2.400 -0.760 -2.140 -0.500 ;
      LAYER met2 ;
        RECT -2.430 -0.500 -2.120 -0.460 ;
        RECT -2.430 -0.720 -0.270 -0.500 ;
        RECT -2.430 -0.790 -2.120 -0.720 ;
    END
  END NFET_DRAIN1
  PIN NFET_DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.688800 ;
    PORT
      LAYER li1 ;
        RECT -1.230 -0.940 -1.060 1.150 ;
        RECT -1.250 -0.980 -0.930 -0.940 ;
        RECT -1.250 -1.170 -0.920 -0.980 ;
        RECT -1.250 -1.200 -0.930 -1.170 ;
        RECT -1.230 -1.250 -1.060 -1.200 ;
      LAYER mcon ;
        RECT -1.190 -1.160 -1.020 -0.990 ;
      LAYER met1 ;
        RECT -1.260 -1.230 -0.940 -0.910 ;
      LAYER via ;
        RECT -1.230 -1.200 -0.970 -0.940 ;
      LAYER met2 ;
        RECT -1.260 -0.950 -0.950 -0.900 ;
        RECT -1.260 -1.160 -0.270 -0.950 ;
        RECT -1.260 -1.230 -0.950 -1.160 ;
    END
  END NFET_DRAIN2
  PIN PFET_DRAIN01
    USE ANALOG ;
    ANTENNADIFFAREA 0.702800 ;
    PORT
      LAYER li1 ;
        RECT -2.410 3.390 -2.240 4.290 ;
        RECT -2.410 3.350 -2.080 3.390 ;
        RECT -2.410 3.160 -2.070 3.350 ;
        RECT -2.410 3.130 -2.080 3.160 ;
        RECT -2.410 1.790 -2.240 3.130 ;
      LAYER mcon ;
        RECT -2.340 3.170 -2.170 3.340 ;
      LAYER met1 ;
        RECT -2.410 3.100 -2.090 3.420 ;
      LAYER via ;
        RECT -2.380 3.130 -2.120 3.390 ;
      LAYER met2 ;
        RECT -2.410 3.380 -2.100 3.430 ;
        RECT -2.410 3.170 -0.270 3.380 ;
        RECT -2.410 3.100 -2.100 3.170 ;
    END
  END PFET_DRAIN01
  PIN PFET_DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.702800 ;
    PORT
      LAYER li1 ;
        RECT -1.230 4.220 -1.060 4.290 ;
        RECT -1.230 4.180 -0.890 4.220 ;
        RECT -1.230 3.990 -0.880 4.180 ;
        RECT -1.230 3.960 -0.890 3.990 ;
        RECT -1.230 1.790 -1.060 3.960 ;
      LAYER mcon ;
        RECT -1.150 4.000 -0.980 4.170 ;
      LAYER met1 ;
        RECT -1.220 3.930 -0.900 4.250 ;
      LAYER via ;
        RECT -1.190 3.960 -0.930 4.220 ;
      LAYER met2 ;
        RECT -1.220 4.210 -0.910 4.260 ;
        RECT -1.220 4.000 -0.270 4.210 ;
        RECT -1.220 3.930 -0.910 4.000 ;
    END
  END PFET_DRAIN2
  OBS
      LAYER nwell ;
        RECT -3.200 1.650 -0.830 4.520 ;
  END
END sky130_hilas_Trans2med

MACRO sky130_hilas_FGBiasWeakGate2x1cell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_FGBiasWeakGate2x1cell ;
  ORIGIN 3.960 3.820 ;
  SIZE 11.530 BY 6.050 ;
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.105400 ;
    PORT
      LAYER li1 ;
        RECT 5.160 1.650 5.690 1.820 ;
      LAYER met1 ;
        RECT 5.090 1.550 5.390 1.930 ;
      LAYER via ;
        RECT 5.110 1.610 5.370 1.880 ;
      LAYER met2 ;
        RECT 5.090 1.750 5.390 1.930 ;
        RECT 4.840 1.730 5.390 1.750 ;
        RECT -3.960 1.550 7.570 1.730 ;
    END
  END DRAIN1
  PIN INPUT1
    PORT
      LAYER li1 ;
        RECT -2.090 1.220 2.970 2.050 ;
        RECT -2.020 1.140 -1.540 1.220 ;
        RECT -2.010 0.890 -1.540 1.140 ;
      LAYER mcon ;
        RECT -1.950 0.930 -1.780 1.100 ;
      LAYER met1 ;
        RECT -2.020 0.860 -1.700 1.180 ;
      LAYER via ;
        RECT -1.990 0.890 -1.730 1.150 ;
      LAYER met2 ;
        RECT -2.020 1.140 -1.710 1.190 ;
        RECT -2.170 1.130 -1.710 1.140 ;
        RECT -3.960 0.950 -1.710 1.130 ;
        RECT -2.020 0.860 -1.710 0.950 ;
    END
  END INPUT1
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER li1 ;
        RECT 5.410 0.740 5.580 1.260 ;
        RECT 5.250 0.480 5.580 0.740 ;
        RECT 5.410 -0.430 5.580 0.480 ;
      LAYER mcon ;
        RECT 5.310 0.520 5.480 0.690 ;
      LAYER met1 ;
        RECT 5.240 0.450 5.560 0.770 ;
      LAYER via ;
        RECT 5.270 0.480 5.530 0.740 ;
      LAYER met2 ;
        RECT 5.240 0.710 5.550 0.780 ;
        RECT 5.240 0.700 7.570 0.710 ;
        RECT -3.960 0.490 7.570 0.700 ;
        RECT -3.960 0.480 6.260 0.490 ;
        RECT 5.240 0.450 5.550 0.480 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER li1 ;
        RECT 5.410 -2.020 5.580 -1.160 ;
        RECT 5.250 -2.280 5.580 -2.020 ;
        RECT 5.410 -2.850 5.580 -2.280 ;
      LAYER mcon ;
        RECT 5.310 -2.240 5.480 -2.070 ;
      LAYER met1 ;
        RECT 5.240 -2.310 5.560 -1.990 ;
      LAYER via ;
        RECT 5.270 -2.280 5.530 -2.020 ;
      LAYER met2 ;
        RECT 5.240 -2.050 5.550 -1.980 ;
        RECT -3.960 -2.260 7.570 -2.050 ;
        RECT -3.960 -2.270 6.260 -2.260 ;
        RECT 5.240 -2.310 5.550 -2.270 ;
    END
  END OUTPUT2
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 4.260 -3.810 7.570 2.220 ;
      LAYER li1 ;
        RECT 6.970 1.550 7.170 1.900 ;
        RECT 6.970 1.520 7.180 1.550 ;
        RECT 6.960 0.940 7.180 1.520 ;
        RECT 6.970 0.930 7.180 0.940 ;
        RECT 6.970 -2.530 7.180 -2.520 ;
        RECT 6.960 -3.110 7.180 -2.530 ;
        RECT 6.970 -3.140 7.180 -3.110 ;
        RECT 6.970 -3.490 7.170 -3.140 ;
      LAYER mcon ;
        RECT 6.980 1.350 7.150 1.520 ;
        RECT 6.980 -3.110 7.150 -2.940 ;
      LAYER met1 ;
        RECT 7.050 1.580 7.330 2.230 ;
        RECT 6.940 0.980 7.330 1.580 ;
        RECT 7.050 -2.570 7.330 0.980 ;
        RECT 6.940 -3.170 7.330 -2.570 ;
        RECT 7.050 -3.820 7.330 -3.170 ;
    END
  END VINJ
  PIN GATESELECT
    USE ANALOG ;
    ANTENNAGATEAREA 0.310000 ;
    PORT
      LAYER li1 ;
        RECT 6.610 0.760 6.800 0.770 ;
        RECT 6.610 0.470 6.810 0.760 ;
        RECT 6.600 0.140 6.840 0.470 ;
        RECT 6.600 -2.060 6.840 -1.730 ;
        RECT 6.610 -2.350 6.810 -2.060 ;
        RECT 6.610 -2.360 6.800 -2.350 ;
      LAYER mcon ;
        RECT 6.620 0.510 6.800 0.700 ;
        RECT 6.620 -2.290 6.800 -2.100 ;
      LAYER met1 ;
        RECT 6.610 0.770 6.800 2.230 ;
        RECT 6.610 0.740 6.830 0.770 ;
        RECT 6.590 0.470 6.840 0.740 ;
        RECT 6.600 0.460 6.840 0.470 ;
        RECT 6.600 0.220 6.830 0.460 ;
        RECT 6.640 -1.810 6.800 0.220 ;
        RECT 6.600 -2.050 6.830 -1.810 ;
        RECT 6.600 -2.060 6.840 -2.050 ;
        RECT 6.590 -2.330 6.840 -2.060 ;
        RECT 6.610 -2.360 6.830 -2.330 ;
        RECT 6.610 -3.820 6.800 -2.360 ;
    END
  END GATESELECT
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT -0.920 -0.740 -0.730 -0.340 ;
        RECT -1.110 -0.750 -0.730 -0.740 ;
        RECT -1.110 -0.930 2.630 -0.750 ;
        RECT -1.110 -0.970 -0.730 -0.930 ;
        RECT -0.920 -1.350 -0.730 -0.970 ;
      LAYER mcon ;
        RECT -1.100 -0.940 -0.930 -0.770 ;
      LAYER met1 ;
        RECT -1.130 1.260 -0.900 2.230 ;
        RECT -1.130 1.010 -0.890 1.260 ;
        RECT -1.130 -3.820 -0.900 1.010 ;
    END
  END VGND
  PIN GATE_CONTROL
    USE ANALOG ;
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT -0.190 -0.160 2.530 1.490 ;
        RECT -0.190 -0.200 2.520 -0.160 ;
        RECT -0.190 -1.530 2.520 -1.490 ;
        RECT -0.190 -3.180 2.530 -1.530 ;
      LAYER li1 ;
        RECT 0.110 0.280 0.340 0.970 ;
        RECT 0.110 -2.660 0.340 -1.930 ;
      LAYER mcon ;
        RECT 0.140 0.770 0.310 0.940 ;
        RECT 0.140 0.320 0.310 0.490 ;
        RECT 0.140 -2.180 0.310 -2.010 ;
        RECT 0.140 -2.630 0.310 -2.460 ;
      LAYER met1 ;
        RECT 0.090 1.020 0.320 2.230 ;
        RECT 0.090 0.230 0.350 1.020 ;
        RECT 0.090 -1.920 0.320 0.230 ;
        RECT 0.090 -2.710 0.350 -1.920 ;
        RECT 0.090 -3.820 0.320 -2.710 ;
    END
  END GATE_CONTROL
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 2.516100 ;
    PORT
      LAYER nwell ;
        RECT -3.950 1.480 -2.220 2.230 ;
        RECT -3.950 -2.090 -2.210 1.480 ;
        RECT -3.950 -3.810 -2.220 -2.090 ;
      LAYER li1 ;
        RECT -3.520 0.090 -2.970 0.520 ;
        RECT -3.520 -1.640 -2.970 -1.210 ;
      LAYER mcon ;
        RECT -3.520 0.170 -3.250 0.440 ;
        RECT -3.520 -1.560 -3.250 -1.290 ;
      LAYER met1 ;
        RECT -3.610 -3.810 -3.190 2.230 ;
    END
  END VTUN
  PIN DRAIN4
    USE ANALOG ;
    ANTENNADIFFAREA 0.105400 ;
    PORT
      LAYER li1 ;
        RECT 5.160 -3.410 5.690 -3.240 ;
      LAYER met1 ;
        RECT 5.090 -3.520 5.390 -3.140 ;
      LAYER via ;
        RECT 5.110 -3.470 5.370 -3.200 ;
      LAYER met2 ;
        RECT 5.100 -3.140 5.260 -3.130 ;
        RECT 5.010 -3.150 7.570 -3.140 ;
        RECT -3.960 -3.300 7.570 -3.150 ;
        RECT 5.010 -3.320 7.570 -3.300 ;
        RECT 5.090 -3.520 5.390 -3.320 ;
    END
  END DRAIN4
  PIN INPUT2
    USE ANALOG ;
    PORT
      LAYER li1 ;
        RECT -2.040 -2.790 -1.700 -2.540 ;
        RECT -2.050 -2.870 -1.700 -2.790 ;
        RECT -2.050 -3.720 3.000 -2.870 ;
      LAYER mcon ;
        RECT -1.980 -2.760 -1.810 -2.590 ;
      LAYER met1 ;
        RECT -2.050 -2.830 -1.730 -2.510 ;
      LAYER via ;
        RECT -2.020 -2.800 -1.760 -2.540 ;
      LAYER met2 ;
        RECT -2.050 -2.580 -1.740 -2.500 ;
        RECT -3.960 -2.790 -1.740 -2.580 ;
        RECT -2.050 -2.830 -1.740 -2.790 ;
    END
  END INPUT2
  PIN COMMONSOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 1.030400 ;
    PORT
      LAYER li1 ;
        RECT 6.240 -0.340 6.410 1.270 ;
        RECT 6.240 -0.530 6.420 -0.340 ;
        RECT 6.240 -1.250 6.420 -1.060 ;
        RECT 6.240 -2.860 6.410 -1.250 ;
      LAYER met1 ;
        RECT 6.210 -0.340 6.450 -0.210 ;
        RECT 6.210 -0.660 6.470 -0.340 ;
        RECT 6.210 -1.260 6.470 -0.940 ;
        RECT 6.210 -1.380 6.450 -1.260 ;
      LAYER via ;
        RECT 6.210 -0.630 6.470 -0.370 ;
        RECT 6.210 -1.230 6.470 -0.970 ;
      LAYER met2 ;
        RECT -3.960 -0.490 6.500 -0.270 ;
        RECT 6.180 -0.630 6.500 -0.490 ;
        RECT 6.220 -0.970 6.480 -0.630 ;
        RECT 6.180 -1.230 6.500 -0.970 ;
    END
  END COMMONSOURCE
  OBS
      LAYER li1 ;
        RECT 3.290 1.070 3.640 1.240 ;
        RECT 4.660 1.070 4.990 1.240 ;
        RECT 3.290 0.280 3.640 0.450 ;
        RECT 4.660 0.280 4.990 0.450 ;
        RECT 3.300 -0.510 3.640 -0.340 ;
        RECT 4.660 -0.510 4.990 -0.340 ;
        RECT 4.740 -1.080 4.910 -0.510 ;
        RECT 3.300 -1.250 3.640 -1.080 ;
        RECT 4.660 -1.250 4.990 -1.080 ;
        RECT 3.290 -2.040 3.640 -1.870 ;
        RECT 4.660 -2.040 4.990 -1.870 ;
        RECT 3.290 -2.830 3.640 -2.660 ;
        RECT 4.660 -2.830 4.990 -2.660 ;
  END
END sky130_hilas_FGBiasWeakGate2x1cell

MACRO sky130_hilas_pFETdevice01a
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pFETdevice01a ;
  ORIGIN 0.800 0.420 ;
  SIZE 1.610 BY 0.850 ;
  OBS
      LAYER nwell ;
        RECT -0.800 -0.420 0.810 0.430 ;
  END
END sky130_hilas_pFETdevice01a

MACRO sky130_hilas_CapModule01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_CapModule01 ;
  ORIGIN 4.430 2.450 ;
  SIZE 2.840 BY 2.860 ;
  OBS
      LAYER met3 ;
        RECT -4.430 -2.450 -1.590 0.410 ;
      LAYER met4 ;
        RECT -3.310 -0.930 -2.860 -0.920 ;
        RECT -3.330 -1.420 -2.810 -0.930 ;
  END
END sky130_hilas_CapModule01

MACRO sky130_hilas_overlapCap02
  CLASS BLOCK ;
  FOREIGN sky130_hilas_overlapCap02 ;
  ORIGIN 5.370 0.690 ;
  SIZE 4.320 BY 1.950 ;
  OBS
      LAYER nwell ;
        RECT -5.370 -0.690 -1.050 1.260 ;
      LAYER li1 ;
        RECT -5.120 -0.430 -1.320 0.980 ;
      LAYER mcon ;
        RECT -3.290 0.540 -3.120 0.710 ;
        RECT -3.290 0.190 -3.120 0.360 ;
        RECT -3.290 -0.150 -3.120 0.020 ;
      LAYER met1 ;
        RECT -3.330 0.130 -3.090 0.770 ;
        RECT -3.320 -0.520 -3.090 0.130 ;
  END
END sky130_hilas_overlapCap02

MACRO sky130_hilas_pTransistorVert01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pTransistorVert01 ;
  ORIGIN 3.630 4.440 ;
  SIZE 1.860 BY 2.990 ;
  OBS
      LAYER nwell ;
        RECT -3.630 -4.440 -1.770 -1.450 ;
      LAYER li1 ;
        RECT -3.220 -3.970 -3.040 -1.920 ;
        RECT -2.410 -3.710 -2.240 -1.930 ;
        RECT -2.490 -3.880 -2.160 -3.710 ;
  END
END sky130_hilas_pTransistorVert01

MACRO sky130_hilas_Tgate4Double01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_Tgate4Double01 ;
  ORIGIN 0.360 1.410 ;
  SIZE 7.080 BY 6.050 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER nwell ;
        RECT -0.240 -1.410 3.230 4.640 ;
      LAYER li1 ;
        RECT 0.070 4.130 0.240 4.410 ;
        RECT 0.070 4.090 0.280 4.130 ;
        RECT 0.070 4.070 0.300 4.090 ;
        RECT 0.070 4.050 0.330 4.070 ;
        RECT 0.070 4.000 0.410 4.050 ;
        RECT 0.070 3.940 0.560 4.000 ;
        RECT 0.070 3.910 0.580 3.940 ;
        RECT 0.110 3.880 0.580 3.910 ;
        RECT 0.240 3.830 0.580 3.880 ;
        RECT 0.360 3.820 0.580 3.830 ;
        RECT 0.370 3.790 0.580 3.820 ;
        RECT 0.390 3.710 0.580 3.790 ;
        RECT 0.390 3.540 0.910 3.710 ;
        RECT 0.390 3.510 0.580 3.540 ;
        RECT 0.390 2.710 0.580 2.740 ;
        RECT 0.390 2.540 0.910 2.710 ;
        RECT 0.390 2.460 0.580 2.540 ;
        RECT 0.370 2.430 0.580 2.460 ;
        RECT 0.360 2.420 0.580 2.430 ;
        RECT 0.240 2.370 0.580 2.420 ;
        RECT 0.110 2.340 0.580 2.370 ;
        RECT 0.070 2.310 0.580 2.340 ;
        RECT 0.070 2.250 0.560 2.310 ;
        RECT 0.070 2.200 0.410 2.250 ;
        RECT 0.070 2.180 0.330 2.200 ;
        RECT 0.070 2.160 0.300 2.180 ;
        RECT 0.070 2.120 0.280 2.160 ;
        RECT 0.070 1.840 0.240 2.120 ;
        RECT 0.070 1.110 0.240 1.390 ;
        RECT 0.070 1.070 0.280 1.110 ;
        RECT 0.070 1.050 0.300 1.070 ;
        RECT 0.070 1.030 0.330 1.050 ;
        RECT 0.070 0.980 0.410 1.030 ;
        RECT 0.070 0.920 0.560 0.980 ;
        RECT 0.070 0.890 0.580 0.920 ;
        RECT 0.110 0.860 0.580 0.890 ;
        RECT 0.240 0.810 0.580 0.860 ;
        RECT 0.360 0.800 0.580 0.810 ;
        RECT 0.370 0.770 0.580 0.800 ;
        RECT 0.390 0.690 0.580 0.770 ;
        RECT 0.390 0.520 0.910 0.690 ;
        RECT 0.390 0.490 0.580 0.520 ;
        RECT 0.390 -0.310 0.580 -0.280 ;
        RECT 0.390 -0.480 0.910 -0.310 ;
        RECT 0.390 -0.560 0.580 -0.480 ;
        RECT 0.370 -0.590 0.580 -0.560 ;
        RECT 0.360 -0.600 0.580 -0.590 ;
        RECT 0.240 -0.650 0.580 -0.600 ;
        RECT 0.110 -0.680 0.580 -0.650 ;
        RECT 0.070 -0.710 0.580 -0.680 ;
        RECT 0.070 -0.770 0.560 -0.710 ;
        RECT 0.070 -0.820 0.410 -0.770 ;
        RECT 0.070 -0.840 0.330 -0.820 ;
        RECT 0.070 -0.860 0.300 -0.840 ;
        RECT 0.070 -0.900 0.280 -0.860 ;
        RECT 0.070 -1.180 0.240 -0.900 ;
      LAYER mcon ;
        RECT 0.400 3.540 0.570 3.710 ;
        RECT 0.400 2.540 0.570 2.710 ;
        RECT 0.400 0.520 0.570 0.690 ;
        RECT 0.400 -0.480 0.570 -0.310 ;
      LAYER met1 ;
        RECT 0.380 3.770 0.580 4.640 ;
        RECT 0.370 3.480 0.600 3.770 ;
        RECT 0.380 2.770 0.580 3.480 ;
        RECT 0.370 2.480 0.600 2.770 ;
        RECT 0.380 0.750 0.580 2.480 ;
        RECT 0.370 0.460 0.600 0.750 ;
        RECT 0.380 -0.250 0.580 0.460 ;
        RECT 0.370 -0.540 0.600 -0.250 ;
        RECT 0.380 -1.410 0.580 -0.540 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.470 3.740 6.640 4.420 ;
        RECT 6.210 3.700 6.640 3.740 ;
        RECT 5.860 3.540 6.640 3.700 ;
        RECT 5.860 3.530 6.400 3.540 ;
        RECT 6.210 3.510 6.400 3.530 ;
        RECT 6.210 2.720 6.400 2.740 ;
        RECT 5.860 2.710 6.400 2.720 ;
        RECT 5.860 2.550 6.640 2.710 ;
        RECT 6.210 2.510 6.640 2.550 ;
        RECT 6.470 1.830 6.640 2.510 ;
        RECT 6.470 0.720 6.640 1.400 ;
        RECT 6.210 0.680 6.640 0.720 ;
        RECT 5.860 0.520 6.640 0.680 ;
        RECT 5.860 0.510 6.400 0.520 ;
        RECT 6.210 0.490 6.400 0.510 ;
        RECT 6.210 -0.300 6.400 -0.280 ;
        RECT 5.860 -0.310 6.400 -0.300 ;
        RECT 5.860 -0.470 6.640 -0.310 ;
        RECT 6.210 -0.510 6.640 -0.470 ;
        RECT 6.470 -1.190 6.640 -0.510 ;
      LAYER mcon ;
        RECT 6.220 3.540 6.390 3.710 ;
        RECT 6.220 2.540 6.390 2.710 ;
        RECT 6.220 0.520 6.390 0.690 ;
        RECT 6.220 -0.480 6.390 -0.310 ;
      LAYER met1 ;
        RECT 6.210 3.770 6.400 4.640 ;
        RECT 6.190 3.480 6.420 3.770 ;
        RECT 6.210 2.770 6.400 3.480 ;
        RECT 6.190 2.480 6.420 2.770 ;
        RECT 6.210 0.750 6.400 2.480 ;
        RECT 6.190 0.460 6.420 0.750 ;
        RECT 6.210 -0.250 6.400 0.460 ;
        RECT 6.190 -0.540 6.420 -0.250 ;
        RECT 6.210 -1.410 6.400 -0.540 ;
    END
  END VGND
  PIN INPUT1_1
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER li1 ;
        RECT 2.100 4.480 2.420 4.510 ;
        RECT 2.100 4.290 2.430 4.480 ;
        RECT 5.180 4.470 5.500 4.500 ;
        RECT 2.100 4.250 2.420 4.290 ;
        RECT 5.180 4.280 5.510 4.470 ;
        RECT 2.130 4.080 2.300 4.250 ;
        RECT 5.180 4.240 5.500 4.280 ;
        RECT 5.240 4.080 5.410 4.240 ;
      LAYER mcon ;
        RECT 2.160 4.300 2.330 4.470 ;
        RECT 5.240 4.290 5.410 4.460 ;
      LAYER met1 ;
        RECT 2.090 4.220 2.410 4.540 ;
        RECT 5.170 4.210 5.490 4.530 ;
      LAYER via ;
        RECT 2.120 4.250 2.380 4.510 ;
        RECT 5.200 4.240 5.460 4.500 ;
      LAYER met2 ;
        RECT 2.090 4.530 2.400 4.540 ;
        RECT -0.360 4.330 5.480 4.530 ;
        RECT 2.090 4.210 2.400 4.330 ;
        RECT 5.170 4.200 5.480 4.330 ;
    END
  END INPUT1_1
  PIN INPUT2_1
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER li1 ;
        RECT 0.580 4.170 0.930 4.340 ;
        RECT 0.750 4.140 0.930 4.170 ;
        RECT 3.780 4.140 3.950 4.420 ;
        RECT 0.750 4.110 1.070 4.140 ;
        RECT 3.670 4.110 3.990 4.140 ;
        RECT 0.750 3.920 1.080 4.110 ;
        RECT 3.670 3.920 4.000 4.110 ;
        RECT 0.750 3.880 1.070 3.920 ;
        RECT 3.670 3.880 3.990 3.920 ;
      LAYER mcon ;
        RECT 0.810 3.930 0.980 4.100 ;
        RECT 3.730 3.930 3.900 4.100 ;
      LAYER met1 ;
        RECT 0.740 3.850 1.060 4.170 ;
        RECT 3.660 3.850 3.980 4.170 ;
      LAYER via ;
        RECT 0.770 3.880 1.030 4.140 ;
        RECT 3.690 3.880 3.950 4.140 ;
      LAYER met2 ;
        RECT 0.740 4.050 1.050 4.170 ;
        RECT 3.660 4.050 3.970 4.170 ;
        RECT -0.360 3.850 4.010 4.050 ;
        RECT 0.740 3.840 1.050 3.850 ;
        RECT 3.660 3.840 3.970 3.850 ;
    END
  END INPUT2_1
  PIN SELECT1
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER li1 ;
        RECT -0.100 3.660 0.070 3.680 ;
        RECT -0.120 3.230 0.090 3.660 ;
      LAYER mcon ;
        RECT -0.100 3.510 0.070 3.680 ;
      LAYER met1 ;
        RECT -0.130 3.550 0.100 3.740 ;
        RECT -0.130 3.450 0.220 3.550 ;
        RECT -0.120 3.230 0.220 3.450 ;
      LAYER via ;
        RECT -0.040 3.260 0.220 3.520 ;
      LAYER met2 ;
        RECT -0.360 3.350 0.250 3.550 ;
        RECT -0.070 3.260 0.250 3.350 ;
    END
  END SELECT1
  PIN SELECT2
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER li1 ;
        RECT -0.120 2.590 0.090 3.020 ;
        RECT -0.100 2.570 0.070 2.590 ;
      LAYER met1 ;
        RECT -0.120 2.800 0.220 3.020 ;
        RECT -0.130 2.700 0.220 2.800 ;
        RECT -0.130 2.510 0.100 2.700 ;
      LAYER via ;
        RECT -0.040 2.730 0.220 2.990 ;
      LAYER met2 ;
        RECT -0.070 2.900 0.250 2.990 ;
        RECT -0.360 2.700 0.250 2.900 ;
    END
  END SELECT2
  PIN INPUT2_2
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER li1 ;
        RECT 0.750 2.330 1.070 2.370 ;
        RECT 3.670 2.330 3.990 2.370 ;
        RECT 0.750 2.140 1.080 2.330 ;
        RECT 3.670 2.140 4.000 2.330 ;
        RECT 0.750 2.110 1.070 2.140 ;
        RECT 3.670 2.110 3.990 2.140 ;
        RECT 0.750 2.080 0.930 2.110 ;
        RECT 0.580 1.910 0.930 2.080 ;
        RECT 3.780 1.830 3.950 2.110 ;
      LAYER mcon ;
        RECT 0.810 2.150 0.980 2.320 ;
        RECT 3.730 2.150 3.900 2.320 ;
      LAYER met1 ;
        RECT 0.740 2.080 1.060 2.400 ;
        RECT 3.660 2.080 3.980 2.400 ;
      LAYER via ;
        RECT 0.770 2.110 1.030 2.370 ;
        RECT 3.690 2.110 3.950 2.370 ;
      LAYER met2 ;
        RECT 0.740 2.400 1.050 2.410 ;
        RECT 3.660 2.400 3.970 2.410 ;
        RECT -0.360 2.200 4.010 2.400 ;
        RECT 0.740 2.080 1.050 2.200 ;
        RECT 3.660 2.080 3.970 2.200 ;
    END
  END INPUT2_2
  PIN INPUT1_2
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER li1 ;
        RECT 2.130 2.000 2.300 2.170 ;
        RECT 5.240 2.010 5.410 2.170 ;
        RECT 2.100 1.960 2.420 2.000 ;
        RECT 5.180 1.970 5.500 2.010 ;
        RECT 2.100 1.770 2.430 1.960 ;
        RECT 5.180 1.780 5.510 1.970 ;
        RECT 2.100 1.740 2.420 1.770 ;
        RECT 5.180 1.750 5.500 1.780 ;
      LAYER mcon ;
        RECT 2.160 1.780 2.330 1.950 ;
        RECT 5.240 1.790 5.410 1.960 ;
      LAYER met1 ;
        RECT 2.090 1.710 2.410 2.030 ;
        RECT 5.170 1.720 5.490 2.040 ;
      LAYER via ;
        RECT 2.120 1.740 2.380 2.000 ;
        RECT 5.200 1.750 5.460 2.010 ;
      LAYER met2 ;
        RECT 2.090 1.920 2.400 2.040 ;
        RECT 5.170 1.920 5.480 2.050 ;
        RECT -0.360 1.720 5.480 1.920 ;
        RECT 2.090 1.710 2.400 1.720 ;
    END
  END INPUT1_2
  PIN SELECT3
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER li1 ;
        RECT -0.100 0.640 0.070 0.660 ;
        RECT -0.120 0.210 0.090 0.640 ;
      LAYER mcon ;
        RECT -0.100 0.490 0.070 0.660 ;
      LAYER met1 ;
        RECT -0.130 0.530 0.100 0.720 ;
        RECT -0.130 0.430 0.220 0.530 ;
        RECT -0.120 0.210 0.220 0.430 ;
      LAYER via ;
        RECT -0.040 0.240 0.220 0.500 ;
      LAYER met2 ;
        RECT -0.360 0.330 0.250 0.530 ;
        RECT -0.070 0.240 0.250 0.330 ;
    END
  END SELECT3
  PIN INPUT2_3
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER li1 ;
        RECT 0.580 1.150 0.930 1.320 ;
        RECT 0.750 1.120 0.930 1.150 ;
        RECT 3.780 1.120 3.950 1.400 ;
        RECT 0.750 1.090 1.070 1.120 ;
        RECT 3.670 1.090 3.990 1.120 ;
        RECT 0.750 0.900 1.080 1.090 ;
        RECT 3.670 0.900 4.000 1.090 ;
        RECT 0.750 0.860 1.070 0.900 ;
        RECT 3.670 0.860 3.990 0.900 ;
      LAYER mcon ;
        RECT 0.810 0.910 0.980 1.080 ;
        RECT 3.730 0.910 3.900 1.080 ;
      LAYER met1 ;
        RECT 0.740 0.830 1.060 1.150 ;
        RECT 3.660 0.830 3.980 1.150 ;
      LAYER via ;
        RECT 0.770 0.860 1.030 1.120 ;
        RECT 3.690 0.860 3.950 1.120 ;
      LAYER met2 ;
        RECT 0.740 1.030 1.050 1.150 ;
        RECT 3.660 1.030 3.970 1.150 ;
        RECT -0.360 0.830 4.010 1.030 ;
        RECT 0.740 0.820 1.050 0.830 ;
        RECT 3.660 0.820 3.970 0.830 ;
    END
  END INPUT2_3
  PIN SELECT4
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER li1 ;
        RECT -0.120 -0.430 0.090 0.000 ;
        RECT -0.100 -0.450 0.070 -0.430 ;
      LAYER met1 ;
        RECT -0.120 -0.220 0.220 0.000 ;
        RECT -0.130 -0.320 0.220 -0.220 ;
        RECT -0.130 -0.510 0.100 -0.320 ;
      LAYER via ;
        RECT -0.040 -0.290 0.220 -0.030 ;
      LAYER met2 ;
        RECT -0.070 -0.120 0.250 -0.030 ;
        RECT -0.360 -0.320 0.250 -0.120 ;
    END
  END SELECT4
  PIN INPUT2_4
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER li1 ;
        RECT 0.750 -0.690 1.070 -0.650 ;
        RECT 3.670 -0.690 3.990 -0.650 ;
        RECT 0.750 -0.880 1.080 -0.690 ;
        RECT 3.670 -0.880 4.000 -0.690 ;
        RECT 0.750 -0.910 1.070 -0.880 ;
        RECT 3.670 -0.910 3.990 -0.880 ;
        RECT 0.750 -0.940 0.930 -0.910 ;
        RECT 0.580 -1.110 0.930 -0.940 ;
        RECT 3.780 -1.190 3.950 -0.910 ;
      LAYER mcon ;
        RECT 0.810 -0.870 0.980 -0.700 ;
        RECT 3.730 -0.870 3.900 -0.700 ;
      LAYER met1 ;
        RECT 0.740 -0.940 1.060 -0.620 ;
        RECT 3.660 -0.940 3.980 -0.620 ;
      LAYER via ;
        RECT 0.770 -0.910 1.030 -0.650 ;
        RECT 3.690 -0.910 3.950 -0.650 ;
      LAYER met2 ;
        RECT 0.740 -0.620 1.050 -0.610 ;
        RECT 3.660 -0.620 3.970 -0.610 ;
        RECT -0.360 -0.820 4.010 -0.620 ;
        RECT 0.740 -0.940 1.050 -0.820 ;
        RECT 3.660 -0.940 3.970 -0.820 ;
    END
  END INPUT2_4
  PIN INPUT1_4
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER li1 ;
        RECT 2.130 -1.020 2.300 -0.850 ;
        RECT 5.240 -1.010 5.410 -0.850 ;
        RECT 2.100 -1.060 2.420 -1.020 ;
        RECT 5.180 -1.050 5.500 -1.010 ;
        RECT 2.100 -1.250 2.430 -1.060 ;
        RECT 5.180 -1.240 5.510 -1.050 ;
        RECT 2.100 -1.280 2.420 -1.250 ;
        RECT 5.180 -1.270 5.500 -1.240 ;
      LAYER mcon ;
        RECT 2.160 -1.240 2.330 -1.070 ;
        RECT 5.240 -1.230 5.410 -1.060 ;
      LAYER met1 ;
        RECT 2.090 -1.310 2.410 -0.990 ;
        RECT 5.170 -1.300 5.490 -0.980 ;
      LAYER via ;
        RECT 2.120 -1.280 2.380 -1.020 ;
        RECT 5.200 -1.270 5.460 -1.010 ;
      LAYER met2 ;
        RECT 2.090 -1.100 2.400 -0.980 ;
        RECT 5.170 -1.100 5.480 -0.970 ;
        RECT -0.360 -1.300 5.480 -1.100 ;
        RECT 2.090 -1.310 2.400 -1.300 ;
    END
  END INPUT1_4
  PIN OUTPUT4
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER li1 ;
        RECT 1.360 -0.700 1.550 -0.690 ;
        RECT 1.350 -0.920 1.550 -0.700 ;
        RECT 2.810 -0.900 3.000 -0.670 ;
        RECT 1.350 -1.190 1.520 -0.920 ;
        RECT 2.820 -1.190 2.990 -0.900 ;
        RECT 4.520 -0.910 4.710 -0.680 ;
        RECT 4.520 -1.200 4.690 -0.910 ;
        RECT 5.750 -0.930 5.940 -0.900 ;
        RECT 5.750 -1.100 6.190 -0.930 ;
        RECT 5.750 -1.130 5.940 -1.100 ;
      LAYER mcon ;
        RECT 1.370 -0.890 1.540 -0.720 ;
        RECT 2.820 -0.870 2.990 -0.700 ;
        RECT 4.530 -0.880 4.700 -0.710 ;
        RECT 5.760 -1.100 5.930 -0.930 ;
      LAYER met1 ;
        RECT 1.350 -0.400 1.610 -0.080 ;
        RECT 2.770 -0.390 3.030 -0.070 ;
        RECT 4.520 -0.370 4.780 -0.050 ;
        RECT 5.560 -0.130 5.820 -0.060 ;
        RECT 1.360 -0.660 1.530 -0.400 ;
        RECT 2.810 -0.640 2.980 -0.390 ;
        RECT 1.340 -0.950 1.570 -0.660 ;
        RECT 2.790 -0.930 3.020 -0.640 ;
        RECT 4.530 -0.650 4.700 -0.370 ;
        RECT 5.560 -0.380 5.920 -0.130 ;
        RECT 4.500 -0.940 4.730 -0.650 ;
        RECT 5.730 -0.870 5.920 -0.380 ;
        RECT 5.730 -1.160 5.960 -0.870 ;
      LAYER via ;
        RECT 1.350 -0.370 1.610 -0.110 ;
        RECT 2.770 -0.360 3.030 -0.100 ;
        RECT 4.520 -0.340 4.780 -0.080 ;
        RECT 5.560 -0.350 5.820 -0.090 ;
      LAYER met2 ;
        RECT 1.320 -0.120 1.640 -0.110 ;
        RECT 2.740 -0.120 3.060 -0.100 ;
        RECT 4.490 -0.120 4.810 -0.080 ;
        RECT 5.530 -0.120 5.850 -0.090 ;
        RECT 1.320 -0.320 6.720 -0.120 ;
        RECT 1.320 -0.370 1.640 -0.320 ;
        RECT 2.740 -0.360 3.060 -0.320 ;
        RECT 4.490 -0.340 4.810 -0.320 ;
        RECT 5.530 -0.350 5.850 -0.320 ;
    END
  END OUTPUT4
  PIN OUTPUT3
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER li1 ;
        RECT 1.350 1.130 1.520 1.400 ;
        RECT 1.350 0.910 1.550 1.130 ;
        RECT 2.820 1.110 2.990 1.400 ;
        RECT 4.520 1.120 4.690 1.410 ;
        RECT 5.750 1.310 5.940 1.340 ;
        RECT 5.750 1.140 6.190 1.310 ;
        RECT 1.360 0.900 1.550 0.910 ;
        RECT 2.810 0.880 3.000 1.110 ;
        RECT 4.520 0.890 4.710 1.120 ;
        RECT 5.750 1.110 5.940 1.140 ;
      LAYER mcon ;
        RECT 5.760 1.140 5.930 1.310 ;
        RECT 1.370 0.930 1.540 1.100 ;
        RECT 2.820 0.910 2.990 1.080 ;
        RECT 4.530 0.920 4.700 1.090 ;
      LAYER met1 ;
        RECT 1.340 0.870 1.570 1.160 ;
        RECT 1.360 0.610 1.530 0.870 ;
        RECT 2.790 0.850 3.020 1.140 ;
        RECT 4.500 0.860 4.730 1.150 ;
        RECT 5.730 1.080 5.960 1.370 ;
        RECT 1.350 0.290 1.610 0.610 ;
        RECT 2.810 0.600 2.980 0.850 ;
        RECT 2.770 0.280 3.030 0.600 ;
        RECT 4.530 0.580 4.700 0.860 ;
        RECT 5.730 0.590 5.920 1.080 ;
        RECT 4.520 0.260 4.780 0.580 ;
        RECT 5.560 0.340 5.920 0.590 ;
        RECT 5.560 0.270 5.820 0.340 ;
      LAYER via ;
        RECT 1.350 0.320 1.610 0.580 ;
        RECT 2.770 0.310 3.030 0.570 ;
        RECT 4.520 0.290 4.780 0.550 ;
        RECT 5.560 0.300 5.820 0.560 ;
      LAYER met2 ;
        RECT 1.320 0.530 1.640 0.580 ;
        RECT 2.740 0.530 3.060 0.570 ;
        RECT 4.490 0.530 4.810 0.550 ;
        RECT 5.530 0.530 5.850 0.560 ;
        RECT 1.320 0.330 6.720 0.530 ;
        RECT 1.320 0.320 1.640 0.330 ;
        RECT 2.740 0.310 3.060 0.330 ;
        RECT 4.490 0.290 4.810 0.330 ;
        RECT 5.530 0.300 5.850 0.330 ;
    END
  END OUTPUT3
  PIN OUTPUT2
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER li1 ;
        RECT 1.360 2.320 1.550 2.330 ;
        RECT 1.350 2.100 1.550 2.320 ;
        RECT 2.810 2.120 3.000 2.350 ;
        RECT 1.350 1.830 1.520 2.100 ;
        RECT 2.820 1.830 2.990 2.120 ;
        RECT 4.520 2.110 4.710 2.340 ;
        RECT 4.520 1.820 4.690 2.110 ;
        RECT 5.750 2.090 5.940 2.120 ;
        RECT 5.750 1.920 6.190 2.090 ;
        RECT 5.750 1.890 5.940 1.920 ;
      LAYER mcon ;
        RECT 1.370 2.130 1.540 2.300 ;
        RECT 2.820 2.150 2.990 2.320 ;
        RECT 4.530 2.140 4.700 2.310 ;
        RECT 5.760 1.920 5.930 2.090 ;
      LAYER met1 ;
        RECT 1.350 2.620 1.610 2.940 ;
        RECT 2.770 2.630 3.030 2.950 ;
        RECT 4.520 2.650 4.780 2.970 ;
        RECT 5.560 2.890 5.820 2.960 ;
        RECT 1.360 2.360 1.530 2.620 ;
        RECT 2.810 2.380 2.980 2.630 ;
        RECT 1.340 2.070 1.570 2.360 ;
        RECT 2.790 2.090 3.020 2.380 ;
        RECT 4.530 2.370 4.700 2.650 ;
        RECT 5.560 2.640 5.920 2.890 ;
        RECT 4.500 2.080 4.730 2.370 ;
        RECT 5.730 2.150 5.920 2.640 ;
        RECT 5.730 1.860 5.960 2.150 ;
      LAYER via ;
        RECT 1.350 2.650 1.610 2.910 ;
        RECT 2.770 2.660 3.030 2.920 ;
        RECT 4.520 2.680 4.780 2.940 ;
        RECT 5.560 2.670 5.820 2.930 ;
      LAYER met2 ;
        RECT 1.320 2.900 1.640 2.910 ;
        RECT 2.740 2.900 3.060 2.920 ;
        RECT 4.490 2.900 4.810 2.940 ;
        RECT 5.530 2.900 5.850 2.930 ;
        RECT 1.320 2.700 6.720 2.900 ;
        RECT 1.320 2.650 1.640 2.700 ;
        RECT 2.740 2.660 3.060 2.700 ;
        RECT 4.490 2.680 4.810 2.700 ;
        RECT 5.530 2.670 5.850 2.700 ;
    END
  END OUTPUT2
  PIN OUTPUT1
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER li1 ;
        RECT 1.350 4.150 1.520 4.420 ;
        RECT 1.350 3.930 1.550 4.150 ;
        RECT 2.820 4.130 2.990 4.420 ;
        RECT 4.520 4.140 4.690 4.430 ;
        RECT 5.750 4.330 5.940 4.360 ;
        RECT 5.750 4.160 6.190 4.330 ;
        RECT 1.360 3.920 1.550 3.930 ;
        RECT 2.810 3.900 3.000 4.130 ;
        RECT 4.520 3.910 4.710 4.140 ;
        RECT 5.750 4.130 5.940 4.160 ;
      LAYER mcon ;
        RECT 5.760 4.160 5.930 4.330 ;
        RECT 1.370 3.950 1.540 4.120 ;
        RECT 2.820 3.930 2.990 4.100 ;
        RECT 4.530 3.940 4.700 4.110 ;
      LAYER met1 ;
        RECT 1.340 3.890 1.570 4.180 ;
        RECT 1.360 3.630 1.530 3.890 ;
        RECT 2.790 3.870 3.020 4.160 ;
        RECT 4.500 3.880 4.730 4.170 ;
        RECT 5.730 4.100 5.960 4.390 ;
        RECT 1.350 3.310 1.610 3.630 ;
        RECT 2.810 3.620 2.980 3.870 ;
        RECT 2.770 3.300 3.030 3.620 ;
        RECT 4.530 3.600 4.700 3.880 ;
        RECT 5.730 3.610 5.920 4.100 ;
        RECT 4.520 3.280 4.780 3.600 ;
        RECT 5.560 3.360 5.920 3.610 ;
        RECT 5.560 3.290 5.820 3.360 ;
      LAYER via ;
        RECT 1.350 3.340 1.610 3.600 ;
        RECT 2.770 3.330 3.030 3.590 ;
        RECT 4.520 3.310 4.780 3.570 ;
        RECT 5.560 3.320 5.820 3.580 ;
      LAYER met2 ;
        RECT 1.320 3.550 1.640 3.600 ;
        RECT 2.740 3.550 3.060 3.590 ;
        RECT 4.490 3.550 4.810 3.570 ;
        RECT 5.530 3.550 5.850 3.580 ;
        RECT 1.320 3.350 6.720 3.550 ;
        RECT 1.320 3.340 1.640 3.350 ;
        RECT 2.740 3.330 3.060 3.350 ;
        RECT 4.490 3.310 4.810 3.350 ;
        RECT 5.530 3.320 5.850 3.350 ;
    END
  END OUTPUT1
  OBS
      LAYER li1 ;
        RECT 1.750 3.710 2.080 3.830 ;
        RECT 1.260 3.530 5.480 3.710 ;
        RECT 1.260 2.540 5.480 2.720 ;
        RECT 1.750 2.420 2.080 2.540 ;
        RECT 2.100 1.460 2.420 1.490 ;
        RECT 2.100 1.270 2.430 1.460 ;
        RECT 5.180 1.450 5.500 1.480 ;
        RECT 2.100 1.230 2.420 1.270 ;
        RECT 5.180 1.260 5.510 1.450 ;
        RECT 2.130 1.060 2.300 1.230 ;
        RECT 5.180 1.220 5.500 1.260 ;
        RECT 5.240 1.060 5.410 1.220 ;
        RECT 1.750 0.690 2.080 0.810 ;
        RECT 1.260 0.510 5.480 0.690 ;
        RECT 1.260 -0.480 5.480 -0.300 ;
        RECT 1.750 -0.600 2.080 -0.480 ;
      LAYER mcon ;
        RECT 2.160 1.280 2.330 1.450 ;
        RECT 5.240 1.270 5.410 1.440 ;
      LAYER met1 ;
        RECT 2.090 1.200 2.410 1.520 ;
        RECT 5.170 1.190 5.490 1.510 ;
      LAYER via ;
        RECT 2.120 1.230 2.380 1.490 ;
        RECT 5.200 1.220 5.460 1.480 ;
      LAYER met2 ;
        RECT 2.090 1.510 2.400 1.520 ;
        RECT -0.360 1.310 5.480 1.510 ;
        RECT 2.090 1.190 2.400 1.310 ;
        RECT 5.170 1.180 5.480 1.310 ;
  END
END sky130_hilas_Tgate4Double01

MACRO sky130_hilas_FGVaractorTunnelCap01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_FGVaractorTunnelCap01 ;
  ORIGIN 10.050 3.800 ;
  SIZE 2.220 BY 1.690 ;
  OBS
      LAYER nwell ;
        RECT -10.050 -3.800 -7.830 -2.110 ;
      LAYER li1 ;
        RECT -9.750 -3.280 -9.520 -2.590 ;
      LAYER mcon ;
        RECT -9.720 -2.800 -9.550 -2.630 ;
        RECT -9.720 -3.250 -9.550 -3.080 ;
      LAYER met1 ;
        RECT -9.770 -3.330 -9.510 -2.540 ;
  END
END sky130_hilas_FGVaractorTunnelCap01

MACRO sky130_hilas_WTAblockSample01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_WTAblockSample01 ;
  ORIGIN 20.050 0.050 ;
  SIZE 33.420 BY 12.030 ;
  OBS
      LAYER nwell ;
        RECT -20.040 11.970 -17.490 11.980 ;
        RECT -20.050 6.000 -17.490 11.970 ;
        RECT -20.050 5.950 -17.460 6.000 ;
        RECT -20.040 5.940 -17.460 5.950 ;
        RECT -15.960 5.990 -13.730 11.970 ;
        RECT -11.710 6.000 -8.270 11.980 ;
        RECT -2.490 11.970 0.060 11.980 ;
        RECT -15.960 5.940 -13.700 5.990 ;
        RECT -20.020 -0.030 -17.460 5.940 ;
        RECT -20.010 -0.040 -17.460 -0.030 ;
        RECT -15.930 -0.040 -13.700 5.940 ;
        RECT -11.710 5.930 -8.240 6.000 ;
        RECT -6.250 5.990 -4.020 11.970 ;
        RECT -2.490 6.000 0.070 11.970 ;
        RECT -2.490 5.990 0.090 6.000 ;
        RECT -6.250 5.940 -3.990 5.990 ;
        RECT -2.490 5.940 0.100 5.990 ;
        RECT -11.680 -0.050 -8.240 5.930 ;
        RECT -6.220 -0.040 -3.990 5.940 ;
        RECT -2.460 -0.030 0.100 5.940 ;
        RECT -2.460 -0.040 0.090 -0.030 ;
      LAYER li1 ;
        RECT 10.630 11.650 10.950 11.680 ;
        RECT -19.650 11.300 -19.450 11.650 ;
        RECT -17.910 11.570 -17.590 11.580 ;
        RECT -18.170 11.400 -17.590 11.570 ;
        RECT -17.920 11.350 -17.590 11.400 ;
        RECT -17.910 11.320 -17.590 11.350 ;
        RECT -2.390 11.570 -2.070 11.580 ;
        RECT -2.390 11.400 -1.810 11.570 ;
        RECT -2.390 11.350 -2.060 11.400 ;
        RECT -2.390 11.320 -2.070 11.350 ;
        RECT -19.660 11.270 -19.450 11.300 ;
        RECT -0.530 11.300 -0.330 11.650 ;
        RECT 10.630 11.480 12.420 11.650 ;
        RECT 10.630 11.460 10.960 11.480 ;
        RECT 10.630 11.420 10.950 11.460 ;
        RECT -19.660 10.680 -19.440 11.270 ;
        RECT -18.920 10.710 -18.720 11.280 ;
        RECT -17.910 10.990 -17.590 11.030 ;
        RECT -17.920 10.950 -17.590 10.990 ;
        RECT -18.170 10.780 -17.590 10.950 ;
        RECT -17.910 10.770 -17.590 10.780 ;
        RECT -2.390 10.990 -2.070 11.030 ;
        RECT -2.390 10.950 -2.060 10.990 ;
        RECT -2.390 10.780 -1.810 10.950 ;
        RECT -2.390 10.770 -2.070 10.780 ;
        RECT -1.260 10.710 -1.060 11.280 ;
        RECT -0.530 11.270 -0.320 11.300 ;
        RECT -0.540 10.680 -0.320 11.270 ;
        RECT 12.250 11.250 12.420 11.480 ;
        RECT 11.100 11.000 11.440 11.250 ;
        RECT 11.610 11.080 11.940 11.250 ;
        RECT 12.160 11.080 12.500 11.250 ;
        RECT 10.780 10.740 11.440 11.000 ;
        RECT 11.690 10.910 11.860 11.080 ;
        RECT 12.250 10.910 12.420 11.080 ;
        RECT 11.610 10.740 11.940 10.910 ;
        RECT 12.160 10.740 12.500 10.910 ;
        RECT 11.690 10.510 11.940 10.740 ;
        RECT 12.820 10.660 13.330 11.330 ;
        RECT 11.690 10.340 12.360 10.510 ;
        RECT -19.660 9.650 -19.440 10.240 ;
        RECT -19.660 9.620 -19.450 9.650 ;
        RECT -18.920 9.640 -18.720 10.210 ;
        RECT -17.910 10.140 -17.590 10.150 ;
        RECT -18.170 9.970 -17.590 10.140 ;
        RECT -17.920 9.930 -17.590 9.970 ;
        RECT -17.910 9.890 -17.590 9.930 ;
        RECT -2.390 10.140 -2.070 10.150 ;
        RECT -2.390 9.970 -1.810 10.140 ;
        RECT -2.390 9.930 -2.060 9.970 ;
        RECT -2.390 9.890 -2.070 9.930 ;
        RECT -1.260 9.640 -1.060 10.210 ;
        RECT -0.540 9.650 -0.320 10.240 ;
        RECT 11.690 10.110 11.940 10.340 ;
        RECT 10.780 9.850 11.440 10.110 ;
        RECT 11.610 9.940 11.940 10.110 ;
        RECT 12.160 9.940 12.500 10.110 ;
        RECT -19.650 9.270 -19.450 9.620 ;
        RECT -0.530 9.620 -0.320 9.650 ;
        RECT -17.910 9.570 -17.590 9.600 ;
        RECT -17.920 9.520 -17.590 9.570 ;
        RECT -18.170 9.350 -17.590 9.520 ;
        RECT -17.910 9.340 -17.590 9.350 ;
        RECT -2.390 9.570 -2.070 9.600 ;
        RECT -2.390 9.520 -2.060 9.570 ;
        RECT -2.390 9.350 -1.810 9.520 ;
        RECT -2.390 9.340 -2.070 9.350 ;
        RECT -0.530 9.270 -0.330 9.620 ;
        RECT 11.100 9.600 11.440 9.850 ;
        RECT 11.690 9.770 11.860 9.940 ;
        RECT 12.250 9.770 12.420 9.940 ;
        RECT 11.610 9.600 11.940 9.770 ;
        RECT 12.160 9.600 12.500 9.770 ;
        RECT 10.630 9.390 10.950 9.430 ;
        RECT 10.630 9.370 10.960 9.390 ;
        RECT 12.250 9.370 12.420 9.600 ;
        RECT 12.820 9.520 13.330 10.190 ;
        RECT 10.630 9.200 12.420 9.370 ;
        RECT 10.630 9.170 10.950 9.200 ;
        RECT -19.280 8.870 -18.840 9.040 ;
        RECT -14.980 8.660 -14.430 9.090 ;
        RECT -10.950 8.730 -10.400 9.160 ;
        RECT -9.580 8.730 -9.030 9.160 ;
        RECT -5.550 8.660 -5.000 9.090 ;
        RECT -1.140 8.870 -0.700 9.040 ;
        RECT 10.630 8.880 10.950 8.910 ;
        RECT 10.630 8.710 12.420 8.880 ;
        RECT 10.630 8.690 10.960 8.710 ;
        RECT 10.630 8.650 10.950 8.690 ;
        RECT -19.650 8.290 -19.450 8.640 ;
        RECT -17.910 8.560 -17.590 8.570 ;
        RECT -18.170 8.390 -17.590 8.560 ;
        RECT -17.920 8.340 -17.590 8.390 ;
        RECT -17.910 8.310 -17.590 8.340 ;
        RECT -2.390 8.560 -2.070 8.570 ;
        RECT -2.390 8.390 -1.810 8.560 ;
        RECT -2.390 8.340 -2.060 8.390 ;
        RECT -2.390 8.310 -2.070 8.340 ;
        RECT -19.660 8.260 -19.450 8.290 ;
        RECT -0.530 8.290 -0.330 8.640 ;
        RECT 12.250 8.480 12.420 8.710 ;
        RECT -19.660 7.670 -19.440 8.260 ;
        RECT -18.920 7.700 -18.720 8.270 ;
        RECT -17.910 7.980 -17.590 8.020 ;
        RECT -17.920 7.940 -17.590 7.980 ;
        RECT -18.170 7.770 -17.590 7.940 ;
        RECT -17.910 7.760 -17.590 7.770 ;
        RECT -2.390 7.980 -2.070 8.020 ;
        RECT -2.390 7.940 -2.060 7.980 ;
        RECT -2.390 7.770 -1.810 7.940 ;
        RECT -2.390 7.760 -2.070 7.770 ;
        RECT -1.260 7.700 -1.060 8.270 ;
        RECT -0.530 8.260 -0.320 8.290 ;
        RECT -0.540 7.670 -0.320 8.260 ;
        RECT 11.100 8.230 11.440 8.480 ;
        RECT 11.610 8.310 11.940 8.480 ;
        RECT 12.160 8.310 12.500 8.480 ;
        RECT 10.780 7.970 11.440 8.230 ;
        RECT 11.690 8.140 11.860 8.310 ;
        RECT 12.250 8.140 12.420 8.310 ;
        RECT 11.610 7.970 11.940 8.140 ;
        RECT 12.160 7.970 12.500 8.140 ;
        RECT 11.690 7.740 11.940 7.970 ;
        RECT 12.820 7.890 13.330 8.560 ;
        RECT 11.690 7.570 12.360 7.740 ;
        RECT 11.690 7.340 11.940 7.570 ;
        RECT -19.660 6.650 -19.440 7.240 ;
        RECT -19.660 6.620 -19.450 6.650 ;
        RECT -18.920 6.640 -18.720 7.210 ;
        RECT -17.910 7.140 -17.590 7.150 ;
        RECT -18.170 6.970 -17.590 7.140 ;
        RECT -17.920 6.930 -17.590 6.970 ;
        RECT -17.910 6.890 -17.590 6.930 ;
        RECT -2.390 7.140 -2.070 7.150 ;
        RECT -2.390 6.970 -1.810 7.140 ;
        RECT -2.390 6.930 -2.060 6.970 ;
        RECT -2.390 6.890 -2.070 6.930 ;
        RECT -1.260 6.640 -1.060 7.210 ;
        RECT -0.540 6.650 -0.320 7.240 ;
        RECT 10.780 7.080 11.440 7.340 ;
        RECT 11.610 7.170 11.940 7.340 ;
        RECT 12.160 7.170 12.500 7.340 ;
        RECT 11.100 6.830 11.440 7.080 ;
        RECT 11.690 7.000 11.860 7.170 ;
        RECT 12.250 7.000 12.420 7.170 ;
        RECT 11.610 6.830 11.940 7.000 ;
        RECT 12.160 6.830 12.500 7.000 ;
        RECT -19.650 6.270 -19.450 6.620 ;
        RECT -0.530 6.620 -0.320 6.650 ;
        RECT 10.630 6.620 10.950 6.660 ;
        RECT -17.910 6.570 -17.590 6.600 ;
        RECT -17.920 6.520 -17.590 6.570 ;
        RECT -18.170 6.350 -17.590 6.520 ;
        RECT -17.910 6.340 -17.590 6.350 ;
        RECT -2.390 6.570 -2.070 6.600 ;
        RECT -2.390 6.520 -2.060 6.570 ;
        RECT -2.390 6.350 -1.810 6.520 ;
        RECT -2.390 6.340 -2.070 6.350 ;
        RECT -0.530 6.270 -0.330 6.620 ;
        RECT 10.630 6.600 10.960 6.620 ;
        RECT 12.250 6.600 12.420 6.830 ;
        RECT 12.820 6.750 13.330 7.420 ;
        RECT 10.630 6.430 12.420 6.600 ;
        RECT 10.630 6.400 10.950 6.430 ;
        RECT 10.650 5.670 10.970 5.700 ;
        RECT -19.620 5.320 -19.420 5.670 ;
        RECT -17.880 5.590 -17.560 5.600 ;
        RECT -18.140 5.420 -17.560 5.590 ;
        RECT -17.890 5.370 -17.560 5.420 ;
        RECT -17.880 5.340 -17.560 5.370 ;
        RECT -2.360 5.590 -2.040 5.600 ;
        RECT -2.360 5.420 -1.780 5.590 ;
        RECT -2.360 5.370 -2.030 5.420 ;
        RECT -2.360 5.340 -2.040 5.370 ;
        RECT -19.630 5.290 -19.420 5.320 ;
        RECT -0.500 5.320 -0.300 5.670 ;
        RECT 10.650 5.500 12.440 5.670 ;
        RECT 10.650 5.480 10.980 5.500 ;
        RECT 10.650 5.440 10.970 5.480 ;
        RECT -19.630 4.700 -19.410 5.290 ;
        RECT -18.890 4.730 -18.690 5.300 ;
        RECT -17.880 5.010 -17.560 5.050 ;
        RECT -17.890 4.970 -17.560 5.010 ;
        RECT -18.140 4.800 -17.560 4.970 ;
        RECT -17.880 4.790 -17.560 4.800 ;
        RECT -2.360 5.010 -2.040 5.050 ;
        RECT -2.360 4.970 -2.030 5.010 ;
        RECT -2.360 4.800 -1.780 4.970 ;
        RECT -2.360 4.790 -2.040 4.800 ;
        RECT -1.230 4.730 -1.030 5.300 ;
        RECT -0.500 5.290 -0.290 5.320 ;
        RECT -0.510 4.700 -0.290 5.290 ;
        RECT 12.270 5.270 12.440 5.500 ;
        RECT 11.120 5.020 11.460 5.270 ;
        RECT 11.630 5.100 11.960 5.270 ;
        RECT 12.180 5.100 12.520 5.270 ;
        RECT 10.800 4.760 11.460 5.020 ;
        RECT 11.710 4.930 11.880 5.100 ;
        RECT 12.270 4.930 12.440 5.100 ;
        RECT 11.630 4.760 11.960 4.930 ;
        RECT 12.180 4.760 12.520 4.930 ;
        RECT 11.710 4.530 11.960 4.760 ;
        RECT 12.840 4.680 13.350 5.350 ;
        RECT 11.710 4.360 12.380 4.530 ;
        RECT -19.630 3.670 -19.410 4.260 ;
        RECT -19.630 3.640 -19.420 3.670 ;
        RECT -18.890 3.660 -18.690 4.230 ;
        RECT -17.880 4.160 -17.560 4.170 ;
        RECT -18.140 3.990 -17.560 4.160 ;
        RECT -17.890 3.950 -17.560 3.990 ;
        RECT -17.880 3.910 -17.560 3.950 ;
        RECT -2.360 4.160 -2.040 4.170 ;
        RECT -2.360 3.990 -1.780 4.160 ;
        RECT -2.360 3.950 -2.030 3.990 ;
        RECT -2.360 3.910 -2.040 3.950 ;
        RECT -1.230 3.660 -1.030 4.230 ;
        RECT -0.510 3.670 -0.290 4.260 ;
        RECT 11.710 4.130 11.960 4.360 ;
        RECT 10.800 3.870 11.460 4.130 ;
        RECT 11.630 3.960 11.960 4.130 ;
        RECT 12.180 3.960 12.520 4.130 ;
        RECT -19.620 3.290 -19.420 3.640 ;
        RECT -0.500 3.640 -0.290 3.670 ;
        RECT -17.880 3.590 -17.560 3.620 ;
        RECT -17.890 3.540 -17.560 3.590 ;
        RECT -18.140 3.370 -17.560 3.540 ;
        RECT -17.880 3.360 -17.560 3.370 ;
        RECT -2.360 3.590 -2.040 3.620 ;
        RECT -2.360 3.540 -2.030 3.590 ;
        RECT -2.360 3.370 -1.780 3.540 ;
        RECT -2.360 3.360 -2.040 3.370 ;
        RECT -0.500 3.290 -0.300 3.640 ;
        RECT 11.120 3.620 11.460 3.870 ;
        RECT 11.710 3.790 11.880 3.960 ;
        RECT 12.270 3.790 12.440 3.960 ;
        RECT 11.630 3.620 11.960 3.790 ;
        RECT 12.180 3.620 12.520 3.790 ;
        RECT 10.650 3.410 10.970 3.450 ;
        RECT 10.650 3.390 10.980 3.410 ;
        RECT 12.270 3.390 12.440 3.620 ;
        RECT 12.840 3.540 13.350 4.210 ;
        RECT 10.650 3.220 12.440 3.390 ;
        RECT 10.650 3.190 10.970 3.220 ;
        RECT -19.250 2.890 -18.810 3.060 ;
        RECT -14.950 2.680 -14.400 3.110 ;
        RECT -10.920 2.750 -10.370 3.180 ;
        RECT -9.550 2.750 -9.000 3.180 ;
        RECT -5.520 2.680 -4.970 3.110 ;
        RECT -1.110 2.890 -0.670 3.060 ;
        RECT 10.650 2.900 10.970 2.930 ;
        RECT 10.650 2.730 12.440 2.900 ;
        RECT 10.650 2.710 10.980 2.730 ;
        RECT 10.650 2.670 10.970 2.710 ;
        RECT -19.620 2.310 -19.420 2.660 ;
        RECT -17.880 2.580 -17.560 2.590 ;
        RECT -18.140 2.410 -17.560 2.580 ;
        RECT -17.890 2.360 -17.560 2.410 ;
        RECT -17.880 2.330 -17.560 2.360 ;
        RECT -2.360 2.580 -2.040 2.590 ;
        RECT -2.360 2.410 -1.780 2.580 ;
        RECT -2.360 2.360 -2.030 2.410 ;
        RECT -2.360 2.330 -2.040 2.360 ;
        RECT -19.630 2.280 -19.420 2.310 ;
        RECT -0.500 2.310 -0.300 2.660 ;
        RECT 12.270 2.500 12.440 2.730 ;
        RECT -19.630 1.690 -19.410 2.280 ;
        RECT -18.890 1.720 -18.690 2.290 ;
        RECT -17.880 2.000 -17.560 2.040 ;
        RECT -17.890 1.960 -17.560 2.000 ;
        RECT -18.140 1.790 -17.560 1.960 ;
        RECT -17.880 1.780 -17.560 1.790 ;
        RECT -2.360 2.000 -2.040 2.040 ;
        RECT -2.360 1.960 -2.030 2.000 ;
        RECT -2.360 1.790 -1.780 1.960 ;
        RECT -2.360 1.780 -2.040 1.790 ;
        RECT -1.230 1.720 -1.030 2.290 ;
        RECT -0.500 2.280 -0.290 2.310 ;
        RECT -0.510 1.690 -0.290 2.280 ;
        RECT 11.120 2.250 11.460 2.500 ;
        RECT 11.630 2.330 11.960 2.500 ;
        RECT 12.180 2.330 12.520 2.500 ;
        RECT 10.800 1.990 11.460 2.250 ;
        RECT 11.710 2.160 11.880 2.330 ;
        RECT 12.270 2.160 12.440 2.330 ;
        RECT 11.630 1.990 11.960 2.160 ;
        RECT 12.180 1.990 12.520 2.160 ;
        RECT 11.710 1.760 11.960 1.990 ;
        RECT 12.840 1.910 13.350 2.580 ;
        RECT 11.710 1.590 12.380 1.760 ;
        RECT 11.710 1.360 11.960 1.590 ;
        RECT -19.630 0.670 -19.410 1.260 ;
        RECT -19.630 0.640 -19.420 0.670 ;
        RECT -18.890 0.660 -18.690 1.230 ;
        RECT -17.880 1.160 -17.560 1.170 ;
        RECT -18.140 0.990 -17.560 1.160 ;
        RECT -17.890 0.950 -17.560 0.990 ;
        RECT -17.880 0.910 -17.560 0.950 ;
        RECT -2.360 1.160 -2.040 1.170 ;
        RECT -2.360 0.990 -1.780 1.160 ;
        RECT -2.360 0.950 -2.030 0.990 ;
        RECT -2.360 0.910 -2.040 0.950 ;
        RECT -1.230 0.660 -1.030 1.230 ;
        RECT -0.510 0.670 -0.290 1.260 ;
        RECT 10.800 1.100 11.460 1.360 ;
        RECT 11.630 1.190 11.960 1.360 ;
        RECT 12.180 1.190 12.520 1.360 ;
        RECT 11.120 0.850 11.460 1.100 ;
        RECT 11.710 1.020 11.880 1.190 ;
        RECT 12.270 1.020 12.440 1.190 ;
        RECT 11.630 0.850 11.960 1.020 ;
        RECT 12.180 0.850 12.520 1.020 ;
        RECT -19.620 0.290 -19.420 0.640 ;
        RECT -0.500 0.640 -0.290 0.670 ;
        RECT 10.650 0.640 10.970 0.680 ;
        RECT -17.880 0.590 -17.560 0.620 ;
        RECT -17.890 0.540 -17.560 0.590 ;
        RECT -18.140 0.370 -17.560 0.540 ;
        RECT -17.880 0.360 -17.560 0.370 ;
        RECT -2.360 0.590 -2.040 0.620 ;
        RECT -2.360 0.540 -2.030 0.590 ;
        RECT -2.360 0.370 -1.780 0.540 ;
        RECT -2.360 0.360 -2.040 0.370 ;
        RECT -0.500 0.290 -0.300 0.640 ;
        RECT 10.650 0.620 10.980 0.640 ;
        RECT 12.270 0.620 12.440 0.850 ;
        RECT 12.840 0.770 13.350 1.440 ;
        RECT 10.650 0.450 12.440 0.620 ;
        RECT 10.650 0.420 10.970 0.450 ;
      LAYER mcon ;
        RECT -17.820 11.360 -17.650 11.530 ;
        RECT -2.330 11.360 -2.160 11.530 ;
        RECT 10.690 11.470 10.860 11.640 ;
        RECT -19.630 11.100 -19.460 11.270 ;
        RECT -18.900 11.070 -18.730 11.240 ;
        RECT -1.250 11.070 -1.080 11.240 ;
        RECT -17.820 10.810 -17.650 10.980 ;
        RECT -2.330 10.810 -2.160 10.980 ;
        RECT -0.520 11.100 -0.350 11.270 ;
        RECT 10.840 10.790 11.010 10.960 ;
        RECT 12.990 10.910 13.160 11.080 ;
        RECT 11.730 10.340 11.900 10.510 ;
        RECT -19.630 9.650 -19.460 9.820 ;
        RECT -17.820 9.940 -17.650 10.110 ;
        RECT -2.330 9.940 -2.160 10.110 ;
        RECT -18.900 9.680 -18.730 9.850 ;
        RECT -1.250 9.680 -1.080 9.850 ;
        RECT 10.840 9.890 11.010 10.060 ;
        RECT -0.520 9.650 -0.350 9.820 ;
        RECT -17.820 9.390 -17.650 9.560 ;
        RECT -2.330 9.390 -2.160 9.560 ;
        RECT 12.990 9.770 13.160 9.940 ;
        RECT 10.690 9.210 10.860 9.380 ;
        RECT -14.700 8.740 -14.430 9.010 ;
        RECT -10.670 8.810 -10.400 9.080 ;
        RECT -9.580 8.810 -9.310 9.080 ;
        RECT -5.550 8.740 -5.280 9.010 ;
        RECT -0.880 8.870 -0.700 9.040 ;
        RECT 10.690 8.700 10.860 8.870 ;
        RECT -17.820 8.350 -17.650 8.520 ;
        RECT -2.330 8.350 -2.160 8.520 ;
        RECT -19.630 8.090 -19.460 8.260 ;
        RECT -18.900 8.060 -18.730 8.230 ;
        RECT -1.250 8.060 -1.080 8.230 ;
        RECT -17.820 7.800 -17.650 7.970 ;
        RECT -2.330 7.800 -2.160 7.970 ;
        RECT -0.520 8.090 -0.350 8.260 ;
        RECT 10.840 8.020 11.010 8.190 ;
        RECT 12.990 8.140 13.160 8.310 ;
        RECT 11.730 7.570 11.900 7.740 ;
        RECT -19.630 6.650 -19.460 6.820 ;
        RECT -17.820 6.940 -17.650 7.110 ;
        RECT -2.330 6.940 -2.160 7.110 ;
        RECT -18.900 6.680 -18.730 6.850 ;
        RECT -1.250 6.680 -1.080 6.850 ;
        RECT 10.840 7.120 11.010 7.290 ;
        RECT 12.990 7.000 13.160 7.170 ;
        RECT -0.520 6.650 -0.350 6.820 ;
        RECT -17.820 6.390 -17.650 6.560 ;
        RECT -2.330 6.390 -2.160 6.560 ;
        RECT 10.690 6.440 10.860 6.610 ;
        RECT -17.790 5.380 -17.620 5.550 ;
        RECT -2.300 5.380 -2.130 5.550 ;
        RECT 10.710 5.490 10.880 5.660 ;
        RECT -19.600 5.120 -19.430 5.290 ;
        RECT -18.870 5.090 -18.700 5.260 ;
        RECT -1.220 5.090 -1.050 5.260 ;
        RECT -17.790 4.830 -17.620 5.000 ;
        RECT -2.300 4.830 -2.130 5.000 ;
        RECT -0.490 5.120 -0.320 5.290 ;
        RECT 10.860 4.810 11.030 4.980 ;
        RECT 13.010 4.930 13.180 5.100 ;
        RECT 11.750 4.360 11.920 4.530 ;
        RECT -19.600 3.670 -19.430 3.840 ;
        RECT -17.790 3.960 -17.620 4.130 ;
        RECT -2.300 3.960 -2.130 4.130 ;
        RECT -18.870 3.700 -18.700 3.870 ;
        RECT -1.220 3.700 -1.050 3.870 ;
        RECT 10.860 3.910 11.030 4.080 ;
        RECT -0.490 3.670 -0.320 3.840 ;
        RECT -17.790 3.410 -17.620 3.580 ;
        RECT -2.300 3.410 -2.130 3.580 ;
        RECT 13.010 3.790 13.180 3.960 ;
        RECT 10.710 3.230 10.880 3.400 ;
        RECT -14.670 2.760 -14.400 3.030 ;
        RECT -10.640 2.830 -10.370 3.100 ;
        RECT -9.550 2.830 -9.280 3.100 ;
        RECT -5.520 2.760 -5.250 3.030 ;
        RECT -0.850 2.890 -0.670 3.060 ;
        RECT 10.710 2.720 10.880 2.890 ;
        RECT -17.790 2.370 -17.620 2.540 ;
        RECT -2.300 2.370 -2.130 2.540 ;
        RECT -19.600 2.110 -19.430 2.280 ;
        RECT -18.870 2.080 -18.700 2.250 ;
        RECT -1.220 2.080 -1.050 2.250 ;
        RECT -17.790 1.820 -17.620 1.990 ;
        RECT -2.300 1.820 -2.130 1.990 ;
        RECT -0.490 2.110 -0.320 2.280 ;
        RECT 10.860 2.040 11.030 2.210 ;
        RECT 13.010 2.160 13.180 2.330 ;
        RECT 11.750 1.590 11.920 1.760 ;
        RECT -19.600 0.670 -19.430 0.840 ;
        RECT -17.790 0.960 -17.620 1.130 ;
        RECT -2.300 0.960 -2.130 1.130 ;
        RECT -18.870 0.700 -18.700 0.870 ;
        RECT -1.220 0.700 -1.050 0.870 ;
        RECT 10.860 1.140 11.030 1.310 ;
        RECT 13.010 1.020 13.180 1.190 ;
        RECT -0.490 0.670 -0.320 0.840 ;
        RECT -17.790 0.410 -17.620 0.580 ;
        RECT -2.300 0.410 -2.130 0.580 ;
        RECT 10.710 0.460 10.880 0.630 ;
      LAYER met1 ;
        RECT -19.690 11.330 -19.530 11.980 ;
        RECT -19.690 10.780 -19.420 11.330 ;
        RECT -19.700 10.730 -19.420 10.780 ;
        RECT -19.280 10.990 -19.090 11.980 ;
        RECT -18.880 11.300 -18.720 11.980 ;
        RECT -18.920 11.280 -18.720 11.300 ;
        RECT -17.900 11.290 -17.580 11.610 ;
        RECT -18.930 11.040 -18.700 11.280 ;
        RECT -19.280 10.870 -19.110 10.990 ;
        RECT -19.700 10.640 -19.530 10.730 ;
        RECT -19.690 10.280 -19.530 10.640 ;
        RECT -19.700 10.190 -19.530 10.280 ;
        RECT -19.700 10.140 -19.420 10.190 ;
        RECT -19.690 9.590 -19.420 10.140 ;
        RECT -19.280 10.050 -19.120 10.870 ;
        RECT -18.920 10.820 -18.720 11.040 ;
        RECT -18.880 10.100 -18.720 10.820 ;
        RECT -17.900 10.740 -17.580 11.060 ;
        RECT -19.280 9.930 -19.110 10.050 ;
        RECT -19.690 8.320 -19.530 9.590 ;
        RECT -19.280 9.070 -19.090 9.930 ;
        RECT -18.920 9.880 -18.720 10.100 ;
        RECT -18.930 9.640 -18.700 9.880 ;
        RECT -17.900 9.860 -17.580 10.180 ;
        RECT -14.760 10.060 -14.380 11.980 ;
        RECT -18.920 9.620 -18.720 9.640 ;
        RECT -19.310 8.840 -19.070 9.070 ;
        RECT -19.690 7.770 -19.420 8.320 ;
        RECT -19.700 7.720 -19.420 7.770 ;
        RECT -19.280 7.980 -19.090 8.840 ;
        RECT -18.880 8.290 -18.720 9.620 ;
        RECT -17.900 9.310 -17.580 9.630 ;
        RECT -18.920 8.270 -18.720 8.290 ;
        RECT -17.900 8.280 -17.580 8.600 ;
        RECT -18.930 8.030 -18.700 8.270 ;
        RECT -14.760 8.200 -14.370 10.060 ;
        RECT -19.280 7.860 -19.110 7.980 ;
        RECT -19.700 7.630 -19.530 7.720 ;
        RECT -19.690 7.280 -19.530 7.630 ;
        RECT -19.700 7.190 -19.530 7.280 ;
        RECT -19.700 7.140 -19.420 7.190 ;
        RECT -19.690 6.590 -19.420 7.140 ;
        RECT -19.280 7.050 -19.120 7.860 ;
        RECT -18.920 7.810 -18.720 8.030 ;
        RECT -18.880 7.100 -18.720 7.810 ;
        RECT -17.900 7.730 -17.580 8.050 ;
        RECT -19.280 6.930 -19.110 7.050 ;
        RECT -19.690 6.000 -19.530 6.590 ;
        RECT -19.280 6.000 -19.090 6.930 ;
        RECT -18.920 6.880 -18.720 7.100 ;
        RECT -18.930 6.640 -18.700 6.880 ;
        RECT -17.900 6.860 -17.580 7.180 ;
        RECT -18.920 6.620 -18.720 6.640 ;
        RECT -18.880 6.000 -18.720 6.620 ;
        RECT -17.900 6.310 -17.580 6.630 ;
        RECT -14.760 6.000 -14.380 8.200 ;
        RECT -10.730 6.000 -10.330 11.980 ;
        RECT -9.650 6.000 -9.250 11.980 ;
        RECT -5.600 10.060 -5.220 11.980 ;
        RECT -2.400 11.290 -2.080 11.610 ;
        RECT -1.260 11.300 -1.100 11.980 ;
        RECT -1.260 11.280 -1.060 11.300 ;
        RECT -2.400 10.740 -2.080 11.060 ;
        RECT -1.280 11.040 -1.050 11.280 ;
        RECT -1.260 10.820 -1.060 11.040 ;
        RECT -0.890 10.990 -0.700 11.980 ;
        RECT -0.450 11.330 -0.290 11.980 ;
        RECT 10.620 11.390 10.940 11.710 ;
        RECT -0.870 10.870 -0.700 10.990 ;
        RECT -5.610 8.200 -5.220 10.060 ;
        RECT -2.400 9.860 -2.080 10.180 ;
        RECT -1.260 10.100 -1.100 10.820 ;
        RECT -1.260 9.880 -1.060 10.100 ;
        RECT -0.860 10.050 -0.700 10.870 ;
        RECT -0.560 10.780 -0.290 11.330 ;
        RECT -0.560 10.730 -0.280 10.780 ;
        RECT -0.450 10.640 -0.280 10.730 ;
        RECT 10.770 10.710 11.090 11.030 ;
        RECT -0.450 10.280 -0.290 10.640 ;
        RECT -0.450 10.190 -0.280 10.280 ;
        RECT -0.870 9.930 -0.700 10.050 ;
        RECT -1.280 9.640 -1.050 9.880 ;
        RECT -2.400 9.310 -2.080 9.630 ;
        RECT -1.260 9.620 -1.060 9.640 ;
        RECT -2.400 8.280 -2.080 8.600 ;
        RECT -1.260 8.290 -1.100 9.620 ;
        RECT -0.890 9.070 -0.700 9.930 ;
        RECT -0.560 10.140 -0.280 10.190 ;
        RECT -0.560 9.590 -0.290 10.140 ;
        RECT 10.770 9.820 11.090 10.140 ;
        RECT -0.910 8.840 -0.670 9.070 ;
        RECT -1.260 8.270 -1.060 8.290 ;
        RECT -5.600 6.000 -5.220 8.200 ;
        RECT -2.400 7.730 -2.080 8.050 ;
        RECT -1.280 8.030 -1.050 8.270 ;
        RECT -1.260 7.810 -1.060 8.030 ;
        RECT -0.890 7.980 -0.700 8.840 ;
        RECT -0.450 8.320 -0.290 9.590 ;
        RECT 10.620 9.140 10.940 9.460 ;
        RECT 10.620 8.620 10.940 8.940 ;
        RECT -0.870 7.860 -0.700 7.980 ;
        RECT -2.400 6.860 -2.080 7.180 ;
        RECT -1.260 7.100 -1.100 7.810 ;
        RECT -1.260 6.880 -1.060 7.100 ;
        RECT -0.860 7.050 -0.700 7.860 ;
        RECT -0.560 7.770 -0.290 8.320 ;
        RECT 10.770 7.940 11.090 8.260 ;
        RECT -0.560 7.720 -0.280 7.770 ;
        RECT -0.450 7.630 -0.280 7.720 ;
        RECT -0.450 7.280 -0.290 7.630 ;
        RECT -0.450 7.190 -0.280 7.280 ;
        RECT -0.870 6.930 -0.700 7.050 ;
        RECT -1.280 6.640 -1.050 6.880 ;
        RECT -2.400 6.310 -2.080 6.630 ;
        RECT -1.260 6.620 -1.060 6.640 ;
        RECT -1.260 6.000 -1.100 6.620 ;
        RECT -0.890 6.000 -0.700 6.930 ;
        RECT -0.560 7.140 -0.280 7.190 ;
        RECT -0.560 6.590 -0.290 7.140 ;
        RECT 10.770 7.050 11.090 7.370 ;
        RECT -0.450 6.000 -0.290 6.590 ;
        RECT 10.620 6.370 10.940 6.690 ;
        RECT 11.700 6.370 11.930 11.710 ;
        RECT 12.960 6.370 13.190 11.710 ;
        RECT -19.690 5.930 -19.500 6.000 ;
        RECT -19.280 5.940 -19.060 6.000 ;
        RECT -18.880 5.940 -18.690 6.000 ;
        RECT -19.660 5.350 -19.500 5.930 ;
        RECT -19.660 4.800 -19.390 5.350 ;
        RECT -19.670 4.750 -19.390 4.800 ;
        RECT -19.250 5.010 -19.060 5.940 ;
        RECT -18.850 5.320 -18.690 5.940 ;
        RECT -14.760 5.930 -14.350 6.000 ;
        RECT -10.730 5.930 -10.300 6.000 ;
        RECT -9.650 5.930 -9.220 6.000 ;
        RECT -5.600 5.930 -5.190 6.000 ;
        RECT -1.260 5.940 -1.070 6.000 ;
        RECT -0.890 5.940 -0.670 6.000 ;
        RECT -0.450 5.940 -0.260 6.000 ;
        RECT -18.890 5.300 -18.690 5.320 ;
        RECT -17.870 5.310 -17.550 5.630 ;
        RECT -18.900 5.060 -18.670 5.300 ;
        RECT -19.250 4.890 -19.080 5.010 ;
        RECT -19.670 4.660 -19.500 4.750 ;
        RECT -19.660 4.300 -19.500 4.660 ;
        RECT -19.670 4.210 -19.500 4.300 ;
        RECT -19.670 4.160 -19.390 4.210 ;
        RECT -19.660 3.610 -19.390 4.160 ;
        RECT -19.250 4.070 -19.090 4.890 ;
        RECT -18.890 4.840 -18.690 5.060 ;
        RECT -18.850 4.120 -18.690 4.840 ;
        RECT -17.870 4.760 -17.550 5.080 ;
        RECT -19.250 3.950 -19.080 4.070 ;
        RECT -19.660 2.340 -19.500 3.610 ;
        RECT -19.250 3.090 -19.060 3.950 ;
        RECT -18.890 3.900 -18.690 4.120 ;
        RECT -18.900 3.660 -18.670 3.900 ;
        RECT -17.870 3.880 -17.550 4.200 ;
        RECT -14.730 4.080 -14.350 5.930 ;
        RECT -18.890 3.640 -18.690 3.660 ;
        RECT -19.280 2.860 -19.040 3.090 ;
        RECT -19.660 1.790 -19.390 2.340 ;
        RECT -19.670 1.740 -19.390 1.790 ;
        RECT -19.250 2.000 -19.060 2.860 ;
        RECT -18.850 2.310 -18.690 3.640 ;
        RECT -17.870 3.330 -17.550 3.650 ;
        RECT -18.890 2.290 -18.690 2.310 ;
        RECT -17.870 2.300 -17.550 2.620 ;
        RECT -18.900 2.050 -18.670 2.290 ;
        RECT -14.730 2.220 -14.340 4.080 ;
        RECT -19.250 1.880 -19.080 2.000 ;
        RECT -19.670 1.650 -19.500 1.740 ;
        RECT -19.660 1.300 -19.500 1.650 ;
        RECT -19.670 1.210 -19.500 1.300 ;
        RECT -19.670 1.160 -19.390 1.210 ;
        RECT -19.660 0.610 -19.390 1.160 ;
        RECT -19.250 1.070 -19.090 1.880 ;
        RECT -18.890 1.830 -18.690 2.050 ;
        RECT -18.850 1.120 -18.690 1.830 ;
        RECT -17.870 1.750 -17.550 2.070 ;
        RECT -19.250 0.950 -19.080 1.070 ;
        RECT -19.660 -0.050 -19.500 0.610 ;
        RECT -19.250 -0.040 -19.060 0.950 ;
        RECT -18.890 0.900 -18.690 1.120 ;
        RECT -18.900 0.660 -18.670 0.900 ;
        RECT -17.870 0.880 -17.550 1.200 ;
        RECT -18.890 0.640 -18.690 0.660 ;
        RECT -18.850 -0.040 -18.690 0.640 ;
        RECT -17.870 0.330 -17.550 0.650 ;
        RECT -14.730 -0.050 -14.350 2.220 ;
        RECT -10.700 -0.050 -10.300 5.930 ;
        RECT -9.620 -0.050 -9.220 5.930 ;
        RECT -5.570 4.080 -5.190 5.930 ;
        RECT -2.370 5.310 -2.050 5.630 ;
        RECT -1.230 5.320 -1.070 5.940 ;
        RECT -1.230 5.300 -1.030 5.320 ;
        RECT -2.370 4.760 -2.050 5.080 ;
        RECT -1.250 5.060 -1.020 5.300 ;
        RECT -1.230 4.840 -1.030 5.060 ;
        RECT -0.860 5.010 -0.670 5.940 ;
        RECT -0.420 5.350 -0.260 5.940 ;
        RECT 10.640 5.410 10.960 5.730 ;
        RECT -0.840 4.890 -0.670 5.010 ;
        RECT -5.580 2.220 -5.190 4.080 ;
        RECT -2.370 3.880 -2.050 4.200 ;
        RECT -1.230 4.120 -1.070 4.840 ;
        RECT -1.230 3.900 -1.030 4.120 ;
        RECT -0.830 4.070 -0.670 4.890 ;
        RECT -0.530 4.800 -0.260 5.350 ;
        RECT -0.530 4.750 -0.250 4.800 ;
        RECT -0.420 4.660 -0.250 4.750 ;
        RECT 10.790 4.730 11.110 5.050 ;
        RECT -0.420 4.300 -0.260 4.660 ;
        RECT -0.420 4.210 -0.250 4.300 ;
        RECT -0.840 3.950 -0.670 4.070 ;
        RECT -1.250 3.660 -1.020 3.900 ;
        RECT -2.370 3.330 -2.050 3.650 ;
        RECT -1.230 3.640 -1.030 3.660 ;
        RECT -2.370 2.300 -2.050 2.620 ;
        RECT -1.230 2.310 -1.070 3.640 ;
        RECT -0.860 3.090 -0.670 3.950 ;
        RECT -0.530 4.160 -0.250 4.210 ;
        RECT -0.530 3.610 -0.260 4.160 ;
        RECT 10.790 3.840 11.110 4.160 ;
        RECT -0.880 2.860 -0.640 3.090 ;
        RECT -1.230 2.290 -1.030 2.310 ;
        RECT -5.570 -0.050 -5.190 2.220 ;
        RECT -2.370 1.750 -2.050 2.070 ;
        RECT -1.250 2.050 -1.020 2.290 ;
        RECT -1.230 1.830 -1.030 2.050 ;
        RECT -0.860 2.000 -0.670 2.860 ;
        RECT -0.420 2.340 -0.260 3.610 ;
        RECT 10.640 3.160 10.960 3.480 ;
        RECT 10.640 2.640 10.960 2.960 ;
        RECT -0.840 1.880 -0.670 2.000 ;
        RECT -2.370 0.880 -2.050 1.200 ;
        RECT -1.230 1.120 -1.070 1.830 ;
        RECT -1.230 0.900 -1.030 1.120 ;
        RECT -0.830 1.070 -0.670 1.880 ;
        RECT -0.530 1.790 -0.260 2.340 ;
        RECT 10.790 1.960 11.110 2.280 ;
        RECT -0.530 1.740 -0.250 1.790 ;
        RECT -0.420 1.650 -0.250 1.740 ;
        RECT -0.420 1.300 -0.260 1.650 ;
        RECT -0.420 1.210 -0.250 1.300 ;
        RECT -0.840 0.950 -0.670 1.070 ;
        RECT -1.250 0.660 -1.020 0.900 ;
        RECT -2.370 0.330 -2.050 0.650 ;
        RECT -1.230 0.640 -1.030 0.660 ;
        RECT -1.230 -0.040 -1.070 0.640 ;
        RECT -0.860 -0.040 -0.670 0.950 ;
        RECT -0.530 1.160 -0.250 1.210 ;
        RECT -0.530 0.610 -0.260 1.160 ;
        RECT 10.790 1.070 11.110 1.390 ;
        RECT -0.420 -0.040 -0.260 0.610 ;
        RECT 10.640 0.390 10.960 0.710 ;
        RECT 11.720 0.390 11.950 5.730 ;
        RECT 12.980 0.390 13.210 5.730 ;
      LAYER via ;
        RECT -17.870 11.320 -17.610 11.580 ;
        RECT -17.870 10.770 -17.610 11.030 ;
        RECT -17.870 9.890 -17.610 10.150 ;
        RECT -17.870 9.340 -17.610 9.600 ;
        RECT -17.870 8.310 -17.610 8.570 ;
        RECT -17.870 7.760 -17.610 8.020 ;
        RECT -17.870 6.890 -17.610 7.150 ;
        RECT -17.870 6.340 -17.610 6.600 ;
        RECT -2.370 11.320 -2.110 11.580 ;
        RECT -2.370 10.770 -2.110 11.030 ;
        RECT 10.650 11.420 10.910 11.680 ;
        RECT -2.370 9.890 -2.110 10.150 ;
        RECT 10.800 10.740 11.060 11.000 ;
        RECT -2.370 9.340 -2.110 9.600 ;
        RECT -2.370 8.310 -2.110 8.570 ;
        RECT 10.800 9.850 11.060 10.110 ;
        RECT -2.370 7.760 -2.110 8.020 ;
        RECT 10.650 9.170 10.910 9.430 ;
        RECT 10.650 8.650 10.910 8.910 ;
        RECT -2.370 6.890 -2.110 7.150 ;
        RECT 10.800 7.970 11.060 8.230 ;
        RECT -2.370 6.340 -2.110 6.600 ;
        RECT 10.800 7.080 11.060 7.340 ;
        RECT 10.650 6.400 10.910 6.660 ;
        RECT -17.840 5.340 -17.580 5.600 ;
        RECT -17.840 4.790 -17.580 5.050 ;
        RECT -17.840 3.910 -17.580 4.170 ;
        RECT -17.840 3.360 -17.580 3.620 ;
        RECT -17.840 2.330 -17.580 2.590 ;
        RECT -17.840 1.780 -17.580 2.040 ;
        RECT -17.840 0.910 -17.580 1.170 ;
        RECT -17.840 0.360 -17.580 0.620 ;
        RECT -2.340 5.340 -2.080 5.600 ;
        RECT -2.340 4.790 -2.080 5.050 ;
        RECT 10.670 5.440 10.930 5.700 ;
        RECT -2.340 3.910 -2.080 4.170 ;
        RECT 10.820 4.760 11.080 5.020 ;
        RECT -2.340 3.360 -2.080 3.620 ;
        RECT -2.340 2.330 -2.080 2.590 ;
        RECT 10.820 3.870 11.080 4.130 ;
        RECT -2.340 1.780 -2.080 2.040 ;
        RECT 10.670 3.190 10.930 3.450 ;
        RECT 10.670 2.670 10.930 2.930 ;
        RECT -2.340 0.910 -2.080 1.170 ;
        RECT 10.820 1.990 11.080 2.250 ;
        RECT -2.340 0.360 -2.080 0.620 ;
        RECT 10.820 1.100 11.080 1.360 ;
        RECT 10.670 0.420 10.930 0.680 ;
      LAYER met2 ;
        RECT 10.620 11.670 10.930 11.710 ;
        RECT -20.050 11.480 -19.910 11.490 ;
        RECT -17.890 11.480 -17.580 11.620 ;
        RECT -2.400 11.480 -2.090 11.620 ;
        RECT -20.050 11.300 0.070 11.480 ;
        RECT 10.520 11.460 10.930 11.670 ;
        RECT 10.620 11.380 10.930 11.460 ;
        RECT -17.890 11.290 -17.580 11.300 ;
        RECT -2.400 11.290 -2.090 11.300 ;
        RECT -17.890 11.050 -17.580 11.070 ;
        RECT -2.400 11.050 -2.090 11.070 ;
        RECT -20.050 10.870 0.070 11.050 ;
        RECT 10.770 10.970 11.080 11.030 ;
        RECT -17.890 10.740 -17.580 10.870 ;
        RECT -2.400 10.740 -2.090 10.870 ;
        RECT 10.770 10.810 13.350 10.970 ;
        RECT 10.770 10.700 11.080 10.810 ;
        RECT -20.050 10.050 -19.980 10.060 ;
        RECT -17.890 10.050 -17.580 10.180 ;
        RECT -2.400 10.050 -2.090 10.180 ;
        RECT -20.050 9.870 0.080 10.050 ;
        RECT 10.770 10.040 11.080 10.150 ;
        RECT 10.770 9.880 13.350 10.040 ;
        RECT -17.890 9.850 -17.580 9.870 ;
        RECT -2.400 9.850 -2.090 9.870 ;
        RECT 10.770 9.820 11.080 9.880 ;
        RECT -17.890 9.620 -17.580 9.630 ;
        RECT -2.400 9.620 -2.090 9.630 ;
        RECT -20.050 9.440 0.080 9.620 ;
        RECT -17.890 9.300 -17.580 9.440 ;
        RECT -2.400 9.300 -2.090 9.440 ;
        RECT 10.620 9.390 10.930 9.470 ;
        RECT 10.520 9.180 10.930 9.390 ;
        RECT 10.620 9.140 10.930 9.180 ;
        RECT 10.620 8.900 10.930 8.940 ;
        RECT 10.520 8.690 10.930 8.900 ;
        RECT 10.620 8.610 10.930 8.690 ;
        RECT -17.890 8.470 -17.580 8.610 ;
        RECT -20.050 8.460 -17.580 8.470 ;
        RECT -2.400 8.470 -2.090 8.610 ;
        RECT -2.400 8.460 0.080 8.470 ;
        RECT -20.050 8.290 0.080 8.460 ;
        RECT -17.890 8.280 -17.580 8.290 ;
        RECT -2.400 8.280 -2.090 8.290 ;
        RECT 10.770 8.200 11.080 8.260 ;
        RECT -17.890 8.040 -17.580 8.060 ;
        RECT -2.400 8.040 -2.090 8.060 ;
        RECT 10.770 8.040 13.350 8.200 ;
        RECT -20.050 7.870 0.080 8.040 ;
        RECT 10.770 7.930 11.080 8.040 ;
        RECT -20.050 7.860 -17.490 7.870 ;
        RECT -2.490 7.860 0.080 7.870 ;
        RECT -17.890 7.730 -17.580 7.860 ;
        RECT -2.400 7.730 -2.090 7.860 ;
        RECT 10.770 7.270 11.080 7.380 ;
        RECT -17.890 7.060 -17.580 7.180 ;
        RECT -2.400 7.060 -2.090 7.180 ;
        RECT -17.890 7.050 -2.090 7.060 ;
        RECT 10.770 7.110 13.350 7.270 ;
        RECT 10.770 7.050 11.080 7.110 ;
        RECT -20.050 6.890 0.080 7.050 ;
        RECT -20.050 6.870 -17.490 6.890 ;
        RECT -17.890 6.850 -17.580 6.870 ;
        RECT -12.310 6.800 -10.770 6.890 ;
        RECT -9.210 6.800 -7.670 6.890 ;
        RECT -2.490 6.870 0.080 6.890 ;
        RECT -2.400 6.850 -2.090 6.870 ;
        RECT -17.890 6.620 -17.580 6.630 ;
        RECT -2.400 6.620 -2.090 6.630 ;
        RECT 10.620 6.620 10.930 6.700 ;
        RECT -20.050 6.450 0.080 6.620 ;
        RECT -20.050 6.440 -17.580 6.450 ;
        RECT -17.890 6.300 -17.580 6.440 ;
        RECT -2.400 6.440 0.080 6.450 ;
        RECT -2.400 6.300 -2.090 6.440 ;
        RECT 10.520 6.410 10.930 6.620 ;
        RECT 10.620 6.370 10.930 6.410 ;
        RECT 10.640 5.690 10.950 5.730 ;
        RECT -20.020 5.500 -19.880 5.510 ;
        RECT -17.860 5.500 -17.550 5.640 ;
        RECT -2.370 5.500 -2.060 5.640 ;
        RECT -20.020 5.320 0.100 5.500 ;
        RECT 10.540 5.480 10.950 5.690 ;
        RECT 10.640 5.400 10.950 5.480 ;
        RECT -17.860 5.310 -17.550 5.320 ;
        RECT -2.370 5.310 -2.060 5.320 ;
        RECT -17.860 5.070 -17.550 5.090 ;
        RECT -2.370 5.070 -2.060 5.090 ;
        RECT -20.020 4.890 0.100 5.070 ;
        RECT 10.790 4.990 11.100 5.050 ;
        RECT -17.860 4.760 -17.550 4.890 ;
        RECT -2.370 4.760 -2.060 4.890 ;
        RECT 10.790 4.830 13.370 4.990 ;
        RECT 10.790 4.720 11.100 4.830 ;
        RECT -20.020 4.070 -19.950 4.080 ;
        RECT -17.860 4.070 -17.550 4.200 ;
        RECT -2.370 4.070 -2.060 4.200 ;
        RECT -20.020 3.890 0.110 4.070 ;
        RECT 10.790 4.060 11.100 4.170 ;
        RECT 10.790 3.900 13.370 4.060 ;
        RECT -17.860 3.870 -17.550 3.890 ;
        RECT -2.370 3.870 -2.060 3.890 ;
        RECT 10.790 3.840 11.100 3.900 ;
        RECT -17.860 3.640 -17.550 3.650 ;
        RECT -2.370 3.640 -2.060 3.650 ;
        RECT -20.020 3.460 0.110 3.640 ;
        RECT -17.860 3.320 -17.550 3.460 ;
        RECT -2.370 3.320 -2.060 3.460 ;
        RECT 10.640 3.410 10.950 3.490 ;
        RECT 10.540 3.200 10.950 3.410 ;
        RECT 10.640 3.160 10.950 3.200 ;
        RECT 10.640 2.920 10.950 2.960 ;
        RECT 10.540 2.710 10.950 2.920 ;
        RECT 10.640 2.630 10.950 2.710 ;
        RECT -17.860 2.490 -17.550 2.630 ;
        RECT -20.020 2.480 -17.550 2.490 ;
        RECT -2.370 2.490 -2.060 2.630 ;
        RECT -2.370 2.480 0.110 2.490 ;
        RECT -20.020 2.310 0.110 2.480 ;
        RECT -17.860 2.300 -17.550 2.310 ;
        RECT -2.370 2.300 -2.060 2.310 ;
        RECT 10.790 2.220 11.100 2.280 ;
        RECT -17.860 2.060 -17.550 2.080 ;
        RECT -2.370 2.060 -2.060 2.080 ;
        RECT 10.790 2.060 13.370 2.220 ;
        RECT -20.020 1.890 0.110 2.060 ;
        RECT 10.790 1.950 11.100 2.060 ;
        RECT -20.020 1.880 -17.460 1.890 ;
        RECT -2.460 1.880 0.110 1.890 ;
        RECT -17.860 1.750 -17.550 1.880 ;
        RECT -2.370 1.750 -2.060 1.880 ;
        RECT 10.790 1.290 11.100 1.400 ;
        RECT -17.860 1.080 -17.550 1.200 ;
        RECT -2.370 1.080 -2.060 1.200 ;
        RECT -17.860 1.070 -2.060 1.080 ;
        RECT 10.790 1.130 13.370 1.290 ;
        RECT 10.790 1.070 11.100 1.130 ;
        RECT -20.020 0.910 0.110 1.070 ;
        RECT -20.020 0.890 -17.460 0.910 ;
        RECT -17.860 0.870 -17.550 0.890 ;
        RECT -12.280 0.820 -10.740 0.910 ;
        RECT -9.180 0.820 -7.640 0.910 ;
        RECT -2.460 0.890 0.110 0.910 ;
        RECT -2.370 0.870 -2.060 0.890 ;
        RECT -17.860 0.640 -17.550 0.650 ;
        RECT -2.370 0.640 -2.060 0.650 ;
        RECT 10.640 0.640 10.950 0.720 ;
        RECT -20.020 0.470 0.110 0.640 ;
        RECT -20.020 0.460 -17.550 0.470 ;
        RECT -17.860 0.320 -17.550 0.460 ;
        RECT -2.370 0.460 0.110 0.470 ;
        RECT -2.370 0.320 -2.060 0.460 ;
        RECT 10.540 0.430 10.950 0.640 ;
        RECT 10.640 0.390 10.950 0.430 ;
  END
END sky130_hilas_WTAblockSample01

MACRO sky130_hilas_li2m2
  CLASS BLOCK ;
  FOREIGN sky130_hilas_li2m2 ;
  ORIGIN 0.140 0.150 ;
  SIZE 0.340 BY 0.330 ;
  OBS
      LAYER li1 ;
        RECT -0.130 0.100 0.190 0.140 ;
        RECT -0.130 -0.090 0.200 0.100 ;
        RECT -0.130 -0.120 0.190 -0.090 ;
      LAYER mcon ;
        RECT -0.070 -0.080 0.100 0.090 ;
      LAYER met1 ;
        RECT -0.140 -0.150 0.180 0.170 ;
      LAYER via ;
        RECT -0.110 -0.120 0.150 0.140 ;
      LAYER met2 ;
        RECT -0.140 -0.150 0.170 0.180 ;
  END
END sky130_hilas_li2m2

MACRO sky130_hilas_DAC_bit6_01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_DAC_bit6_01 ;
  ORIGIN -4.020 -5.240 ;
  SIZE 16.380 BY 13.680 ;
  OBS
      LAYER nwell ;
        RECT 5.760 18.660 7.370 18.920 ;
        RECT 5.630 13.270 7.370 18.660 ;
        RECT 5.630 13.010 7.240 13.270 ;
        RECT 4.190 5.270 5.800 10.920 ;
        RECT 7.520 10.200 17.620 10.270 ;
        RECT 18.680 5.270 20.290 10.920 ;
      LAYER li1 ;
        RECT 6.140 17.440 6.310 17.700 ;
        RECT 6.820 17.440 6.990 17.700 ;
        RECT 6.010 17.370 6.310 17.440 ;
        RECT 6.690 17.370 6.990 17.440 ;
        RECT 6.010 17.110 6.180 17.370 ;
        RECT 6.690 17.110 6.860 17.370 ;
        RECT 6.140 16.480 6.310 16.740 ;
        RECT 6.820 16.480 6.990 16.740 ;
        RECT 6.010 16.410 6.310 16.480 ;
        RECT 6.690 16.410 6.990 16.480 ;
        RECT 6.010 16.150 6.180 16.410 ;
        RECT 6.690 16.150 6.860 16.410 ;
        RECT 6.140 15.520 6.310 15.780 ;
        RECT 6.820 15.520 6.990 15.780 ;
        RECT 6.010 15.450 6.310 15.520 ;
        RECT 6.690 15.450 6.990 15.520 ;
        RECT 6.010 15.190 6.180 15.450 ;
        RECT 6.690 15.190 6.860 15.450 ;
        RECT 6.140 14.560 6.310 14.820 ;
        RECT 6.820 14.560 6.990 14.820 ;
        RECT 6.010 14.490 6.310 14.560 ;
        RECT 6.690 14.490 6.990 14.560 ;
        RECT 6.010 14.230 6.180 14.490 ;
        RECT 6.690 14.230 6.860 14.490 ;
        RECT 4.220 10.710 4.430 11.140 ;
        RECT 5.810 10.720 6.020 11.150 ;
        RECT 7.210 10.740 7.640 10.760 ;
        RECT 4.240 10.690 4.410 10.710 ;
        RECT 5.830 10.700 6.000 10.720 ;
        RECT 7.190 10.570 7.640 10.740 ;
        RECT 9.010 10.710 9.220 11.140 ;
        RECT 10.620 10.710 10.830 11.140 ;
        RECT 12.240 10.710 12.450 11.140 ;
        RECT 13.850 10.720 14.060 11.150 ;
        RECT 15.460 10.720 15.670 11.150 ;
        RECT 16.770 11.040 16.980 11.050 ;
        RECT 16.660 11.000 16.980 11.040 ;
        RECT 17.330 11.000 17.650 11.040 ;
        RECT 16.660 10.810 16.990 11.000 ;
        RECT 17.330 10.810 17.660 11.000 ;
        RECT 16.660 10.780 16.980 10.810 ;
        RECT 17.330 10.780 17.650 10.810 ;
        RECT 9.030 10.690 9.200 10.710 ;
        RECT 10.640 10.690 10.810 10.710 ;
        RECT 12.260 10.690 12.430 10.710 ;
        RECT 13.870 10.700 14.040 10.720 ;
        RECT 15.480 10.700 15.650 10.720 ;
        RECT 7.210 10.550 7.640 10.570 ;
        RECT 7.800 10.270 7.970 10.280 ;
        RECT 16.770 10.270 16.980 10.780 ;
        RECT 17.440 10.270 17.610 10.780 ;
        RECT 6.190 10.040 17.620 10.270 ;
        RECT 4.080 9.400 4.290 9.830 ;
        RECT 4.100 9.380 4.270 9.400 ;
        RECT 4.140 8.450 4.350 8.880 ;
        RECT 4.160 8.430 4.330 8.450 ;
        RECT 4.140 7.510 4.350 7.940 ;
        RECT 4.160 7.490 4.330 7.510 ;
        RECT 6.190 6.480 6.360 10.040 ;
        RECT 6.850 5.500 7.020 9.710 ;
        RECT 7.800 6.480 7.970 10.040 ;
        RECT 8.480 5.500 8.650 9.670 ;
        RECT 9.390 6.480 9.560 10.040 ;
        RECT 10.080 5.500 10.250 9.750 ;
        RECT 11.010 6.480 11.180 10.040 ;
        RECT 11.700 5.500 11.870 9.700 ;
        RECT 12.630 6.500 12.800 10.040 ;
        RECT 13.300 5.500 13.470 9.750 ;
        RECT 14.230 6.510 14.400 10.040 ;
        RECT 14.920 5.500 15.090 9.750 ;
        RECT 15.840 6.500 16.010 10.040 ;
        RECT 16.520 5.500 16.690 9.730 ;
        RECT 17.450 6.470 17.620 10.040 ;
        RECT 18.130 5.500 18.300 9.910 ;
        RECT 6.850 5.270 7.040 5.500 ;
        RECT 8.470 5.270 8.660 5.500 ;
        RECT 10.070 5.270 10.260 5.500 ;
        RECT 11.690 5.270 11.880 5.500 ;
        RECT 13.290 5.270 13.480 5.500 ;
        RECT 14.910 5.270 15.100 5.500 ;
        RECT 16.510 5.270 16.700 5.500 ;
        RECT 18.120 5.270 18.310 5.500 ;
        RECT 6.850 5.250 7.020 5.270 ;
        RECT 8.480 5.250 8.650 5.270 ;
        RECT 10.080 5.250 10.250 5.270 ;
        RECT 11.700 5.250 11.870 5.270 ;
        RECT 13.300 5.250 13.470 5.270 ;
        RECT 14.920 5.250 15.090 5.270 ;
        RECT 16.520 5.250 16.690 5.270 ;
        RECT 18.130 5.250 18.300 5.270 ;
      LAYER mcon ;
        RECT 16.720 10.820 16.890 10.990 ;
        RECT 17.390 10.820 17.560 10.990 ;
        RECT 6.860 5.300 7.030 5.470 ;
        RECT 8.480 5.300 8.650 5.470 ;
        RECT 10.080 5.300 10.250 5.470 ;
        RECT 11.700 5.300 11.870 5.470 ;
        RECT 13.300 5.300 13.470 5.470 ;
        RECT 14.920 5.300 15.090 5.470 ;
        RECT 16.520 5.300 16.690 5.470 ;
        RECT 18.130 5.300 18.300 5.470 ;
      LAYER met1 ;
        RECT 4.170 10.860 4.490 11.180 ;
        RECT 5.760 10.870 6.080 11.190 ;
        RECT 4.210 10.630 4.440 10.860 ;
        RECT 5.800 10.640 6.030 10.870 ;
        RECT 8.960 10.860 9.280 11.180 ;
        RECT 10.570 10.860 10.890 11.180 ;
        RECT 12.190 10.860 12.510 11.180 ;
        RECT 13.800 10.870 14.120 11.190 ;
        RECT 15.410 10.870 15.730 11.190 ;
        RECT 7.360 10.770 7.680 10.810 ;
        RECT 7.130 10.540 7.680 10.770 ;
        RECT 9.000 10.630 9.230 10.860 ;
        RECT 10.610 10.630 10.840 10.860 ;
        RECT 12.230 10.630 12.460 10.860 ;
        RECT 13.840 10.640 14.070 10.870 ;
        RECT 15.450 10.640 15.680 10.870 ;
        RECT 16.650 10.750 16.970 11.070 ;
        RECT 17.320 10.750 17.640 11.070 ;
        RECT 7.360 10.490 7.680 10.540 ;
        RECT 4.030 9.550 4.350 9.870 ;
        RECT 4.070 9.320 4.300 9.550 ;
        RECT 4.090 8.600 4.410 8.920 ;
        RECT 10.560 8.800 14.010 8.970 ;
        RECT 4.130 8.370 4.360 8.600 ;
        RECT 4.090 7.660 4.410 7.980 ;
        RECT 4.130 7.430 4.360 7.660 ;
        RECT 12.110 6.290 12.290 7.810 ;
        RECT 13.810 6.960 14.010 8.800 ;
        RECT 12.110 5.970 12.370 6.290 ;
        RECT 6.830 5.480 7.060 5.530 ;
        RECT 8.450 5.480 8.680 5.530 ;
        RECT 10.050 5.480 10.280 5.530 ;
        RECT 11.670 5.480 11.900 5.530 ;
        RECT 13.270 5.480 13.500 5.530 ;
        RECT 14.890 5.480 15.120 5.530 ;
        RECT 16.490 5.480 16.720 5.530 ;
        RECT 18.100 5.480 18.330 5.530 ;
        RECT 6.830 5.250 20.300 5.480 ;
        RECT 6.830 5.240 7.060 5.250 ;
        RECT 8.450 5.240 8.680 5.250 ;
        RECT 10.050 5.240 10.280 5.250 ;
        RECT 11.670 5.240 11.900 5.250 ;
        RECT 13.270 5.240 13.500 5.250 ;
        RECT 14.890 5.240 15.120 5.250 ;
        RECT 16.490 5.240 16.720 5.250 ;
        RECT 18.100 5.240 18.330 5.250 ;
      LAYER via ;
        RECT 4.200 10.890 4.460 11.150 ;
        RECT 5.790 10.900 6.050 11.160 ;
        RECT 8.990 10.890 9.250 11.150 ;
        RECT 10.600 10.890 10.860 11.150 ;
        RECT 12.220 10.890 12.480 11.150 ;
        RECT 13.830 10.900 14.090 11.160 ;
        RECT 15.440 10.900 15.700 11.160 ;
        RECT 7.390 10.520 7.650 10.780 ;
        RECT 16.680 10.780 16.940 11.040 ;
        RECT 17.350 10.780 17.610 11.040 ;
        RECT 4.060 9.580 4.320 9.840 ;
        RECT 4.120 8.630 4.380 8.890 ;
        RECT 4.120 7.690 4.380 7.950 ;
        RECT 12.110 6.000 12.370 6.260 ;
      LAYER met2 ;
        RECT 4.180 11.180 10.870 11.210 ;
        RECT 4.170 11.020 10.890 11.180 ;
        RECT 4.170 10.860 4.490 11.020 ;
        RECT 5.760 10.870 6.080 11.020 ;
        RECT 8.960 10.860 9.280 11.020 ;
        RECT 10.570 10.860 10.890 11.020 ;
        RECT 12.190 10.860 12.510 11.180 ;
        RECT 13.800 10.890 14.120 11.190 ;
        RECT 13.800 10.870 14.130 10.890 ;
        RECT 15.410 10.870 15.730 11.190 ;
        RECT 16.530 10.930 17.690 11.210 ;
        RECT 7.360 10.660 7.680 10.810 ;
        RECT 7.300 10.490 7.680 10.660 ;
        RECT 4.180 10.200 5.880 10.260 ;
        RECT 7.300 10.200 7.520 10.490 ;
        RECT 12.220 10.210 12.470 10.860 ;
        RECT 12.220 10.200 12.500 10.210 ;
        RECT 4.180 10.050 12.500 10.200 ;
        RECT 4.180 9.870 4.280 10.050 ;
        RECT 5.720 9.900 12.500 10.050 ;
        RECT 4.030 9.550 4.350 9.870 ;
        RECT 4.090 8.600 4.410 8.920 ;
        RECT 13.930 8.330 14.130 10.870 ;
        RECT 4.180 8.120 14.130 8.330 ;
        RECT 4.090 7.660 4.410 7.980 ;
        RECT 15.530 7.350 15.680 10.870 ;
        RECT 16.650 10.750 16.960 10.930 ;
        RECT 17.280 10.920 17.690 10.930 ;
        RECT 17.320 10.750 17.630 10.920 ;
        RECT 4.180 7.150 15.690 7.350 ;
        RECT 12.080 6.230 12.400 6.260 ;
        RECT 4.180 6.030 12.400 6.230 ;
        RECT 12.080 6.000 12.400 6.030 ;
  END
END sky130_hilas_DAC_bit6_01

MACRO sky130_hilas_WTAsinglestage01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_WTAsinglestage01 ;
  ORIGIN 1.080 0.760 ;
  SIZE 2.830 BY 1.430 ;
  OBS
      LAYER li1 ;
        RECT 0.110 0.610 0.320 0.630 ;
        RECT 0.090 0.440 0.760 0.610 ;
        RECT 0.090 0.210 0.340 0.440 ;
        RECT -0.820 -0.050 -0.160 0.210 ;
        RECT 0.010 0.040 0.340 0.210 ;
        RECT 0.560 0.040 0.900 0.210 ;
        RECT -0.500 -0.300 -0.160 -0.050 ;
        RECT 0.090 -0.130 0.260 0.040 ;
        RECT 0.650 -0.130 0.820 0.040 ;
        RECT 0.010 -0.300 0.340 -0.130 ;
        RECT 0.560 -0.300 0.900 -0.130 ;
        RECT -0.970 -0.510 -0.650 -0.470 ;
        RECT -0.970 -0.530 -0.640 -0.510 ;
        RECT 0.650 -0.530 0.820 -0.300 ;
        RECT 1.220 -0.380 1.730 0.290 ;
        RECT -0.970 -0.700 0.820 -0.530 ;
        RECT -0.970 -0.730 -0.650 -0.700 ;
      LAYER mcon ;
        RECT 0.130 0.440 0.300 0.610 ;
        RECT -0.760 -0.010 -0.590 0.160 ;
        RECT 1.390 -0.130 1.560 0.040 ;
        RECT -0.910 -0.690 -0.740 -0.520 ;
      LAYER met1 ;
        RECT -0.830 -0.080 -0.510 0.240 ;
        RECT -0.980 -0.760 -0.660 -0.440 ;
        RECT 0.100 -0.760 0.330 0.670 ;
        RECT 1.360 -0.760 1.590 0.530 ;
      LAYER via ;
        RECT -0.800 -0.050 -0.540 0.210 ;
        RECT -0.950 -0.730 -0.690 -0.470 ;
      LAYER met2 ;
        RECT -0.830 0.140 -0.520 0.250 ;
        RECT -0.830 -0.020 1.750 0.140 ;
        RECT -0.830 -0.080 -0.520 -0.020 ;
        RECT -0.980 -0.510 -0.670 -0.430 ;
        RECT -1.080 -0.720 -0.670 -0.510 ;
        RECT -0.980 -0.760 -0.670 -0.720 ;
  END
END sky130_hilas_WTAsinglestage01

MACRO sky130_hilas_TACoreBlock
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TACoreBlock ;
  ORIGIN 4.570 0.970 ;
  SIZE 9.540 BY 5.020 ;
  OBS
      LAYER nwell ;
        RECT -4.570 2.190 -2.340 4.040 ;
        RECT 2.410 2.130 4.970 3.970 ;
        RECT 2.410 2.120 4.960 2.130 ;
        RECT -4.310 -0.970 -2.580 0.930 ;
      LAYER li1 ;
        RECT 2.510 3.320 2.830 3.330 ;
        RECT 2.510 3.150 3.090 3.320 ;
        RECT 2.510 3.110 2.840 3.150 ;
        RECT 2.510 3.070 2.830 3.110 ;
        RECT 3.640 2.820 3.840 3.390 ;
        RECT 4.360 2.830 4.580 3.420 ;
        RECT 4.370 2.800 4.580 2.830 ;
        RECT 2.510 2.750 2.830 2.780 ;
        RECT 2.510 2.700 2.840 2.750 ;
        RECT 2.510 2.530 3.090 2.700 ;
        RECT 2.510 2.520 2.830 2.530 ;
        RECT 4.370 2.450 4.570 2.800 ;
        RECT -0.080 -0.130 0.250 0.040 ;
      LAYER mcon ;
        RECT 2.570 3.120 2.740 3.290 ;
        RECT 3.650 2.860 3.820 3.030 ;
        RECT 4.380 2.830 4.550 3.000 ;
        RECT 2.570 2.570 2.740 2.740 ;
      LAYER met1 ;
        RECT -3.920 2.190 -3.540 4.050 ;
        RECT 2.500 3.040 2.820 3.360 ;
        RECT 3.640 3.280 3.800 3.970 ;
        RECT 3.640 3.060 3.840 3.280 ;
        RECT 4.040 3.230 4.200 3.970 ;
        RECT 4.450 3.460 4.610 3.970 ;
        RECT 4.450 3.370 4.620 3.460 ;
        RECT 4.030 3.110 4.200 3.230 ;
        RECT 3.620 2.820 3.850 3.060 ;
        RECT 2.500 2.490 2.820 2.810 ;
        RECT 3.640 2.800 3.840 2.820 ;
        RECT 3.640 2.120 3.800 2.800 ;
        RECT 4.010 2.120 4.200 3.110 ;
        RECT 4.340 3.320 4.620 3.370 ;
        RECT 4.340 2.770 4.610 3.320 ;
        RECT 4.450 2.120 4.610 2.770 ;
      LAYER via ;
        RECT 2.530 3.070 2.790 3.330 ;
        RECT 2.530 2.520 2.790 2.780 ;
      LAYER met2 ;
        RECT 2.500 3.230 2.810 3.360 ;
        RECT 2.410 3.050 4.970 3.230 ;
        RECT 2.500 3.030 2.810 3.050 ;
        RECT 2.500 2.800 2.810 2.810 ;
        RECT 2.500 2.620 4.970 2.800 ;
        RECT 2.500 2.480 2.810 2.620 ;
  END
END sky130_hilas_TACoreBlock

MACRO sky130_hilas_pFETdevice01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pFETdevice01 ;
  ORIGIN 0.790 0.780 ;
  SIZE 1.610 BY 1.210 ;
  OBS
      LAYER nwell ;
        RECT -0.790 -0.780 0.820 0.430 ;
      LAYER li1 ;
        RECT -0.410 -0.160 -0.240 0.170 ;
        RECT 0.270 -0.160 0.440 0.170 ;
  END
END sky130_hilas_pFETdevice01

MACRO sky130_hilas_pFETdevice01ba
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pFETdevice01ba ;
  ORIGIN 0.790 1.140 ;
  SIZE 1.870 BY 1.570 ;
  OBS
      LAYER nwell ;
        RECT -0.790 -0.780 0.820 0.430 ;
      LAYER li1 ;
        RECT 0.780 -1.060 0.990 -0.630 ;
        RECT 0.800 -1.080 0.970 -1.060 ;
      LAYER met1 ;
        RECT 0.780 -0.850 1.000 -0.630 ;
        RECT 0.770 -1.140 1.000 -0.850 ;
  END
END sky130_hilas_pFETdevice01ba

MACRO sky130_hilas_overlapCap01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_overlapCap01 ;
  ORIGIN 2.870 0.710 ;
  SIZE 2.870 BY 2.080 ;
  OBS
      LAYER nwell ;
        RECT -2.810 -0.650 -0.090 1.310 ;
      LAYER li1 ;
        RECT -2.410 -0.260 -0.460 0.910 ;
      LAYER mcon ;
        RECT -1.930 0.570 -1.760 0.740 ;
        RECT -1.930 0.230 -1.760 0.400 ;
        RECT -1.930 -0.110 -1.760 0.060 ;
      LAYER met1 ;
        RECT -1.970 0.320 -1.710 0.800 ;
        RECT -1.980 -0.200 -1.710 0.320 ;
        RECT -1.980 -0.650 -1.720 -0.200 ;
  END
END sky130_hilas_overlapCap01

MACRO sky130_hilas_swc4x1cellOverlap
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc4x1cellOverlap ;
  ORIGIN 2.640 4.130 ;
  SIZE 10.080 BY 6.710 ;
  OBS
      LAYER nwell ;
        RECT 2.230 2.230 4.950 2.520 ;
        RECT -2.630 0.370 -0.900 2.230 ;
        RECT -2.640 -1.470 -0.900 0.370 ;
        RECT 2.230 2.220 7.430 2.230 ;
        RECT 2.230 -0.570 7.440 2.220 ;
        RECT -2.630 -3.820 -0.900 -1.470 ;
        RECT 2.220 -3.800 7.440 -0.570 ;
        RECT 2.220 -3.810 7.430 -3.800 ;
        RECT 2.220 -4.070 4.940 -3.810 ;
      LAYER li1 ;
        RECT 2.630 0.950 4.580 2.120 ;
        RECT 4.980 1.820 5.300 1.830 ;
        RECT 4.980 1.650 5.560 1.820 ;
        RECT 4.980 1.600 5.310 1.650 ;
        RECT 4.980 1.570 5.300 1.600 ;
        RECT 6.840 1.550 7.040 1.900 ;
        RECT 4.980 1.240 5.300 1.280 ;
        RECT 4.980 1.200 5.310 1.240 ;
        RECT 4.980 1.030 5.560 1.200 ;
        RECT 4.980 1.020 5.300 1.030 ;
        RECT 6.110 0.960 6.310 1.530 ;
        RECT 6.840 1.520 7.050 1.550 ;
        RECT 6.830 0.930 7.050 1.520 ;
        RECT 2.630 -0.580 4.580 0.590 ;
        RECT 4.980 0.390 5.300 0.400 ;
        RECT 4.980 0.220 5.560 0.390 ;
        RECT 4.980 0.180 5.310 0.220 ;
        RECT 4.980 0.140 5.300 0.180 ;
        RECT 6.110 -0.110 6.310 0.460 ;
        RECT 6.830 -0.100 7.050 0.490 ;
        RECT 6.840 -0.130 7.050 -0.100 ;
        RECT 4.980 -0.180 5.300 -0.150 ;
        RECT 4.980 -0.230 5.310 -0.180 ;
        RECT 4.980 -0.400 5.560 -0.230 ;
        RECT 4.980 -0.410 5.300 -0.400 ;
        RECT 6.840 -0.480 7.040 -0.130 ;
        RECT -2.210 -1.020 -1.660 -0.590 ;
        RECT 6.230 -0.880 6.670 -0.710 ;
        RECT 2.620 -2.140 4.570 -0.970 ;
        RECT 4.980 -1.190 5.300 -1.180 ;
        RECT 4.980 -1.360 5.560 -1.190 ;
        RECT 4.980 -1.410 5.310 -1.360 ;
        RECT 4.980 -1.440 5.300 -1.410 ;
        RECT 6.840 -1.460 7.040 -1.110 ;
        RECT 4.980 -1.770 5.300 -1.730 ;
        RECT 4.980 -1.810 5.310 -1.770 ;
        RECT 4.980 -1.980 5.560 -1.810 ;
        RECT 4.980 -1.990 5.300 -1.980 ;
        RECT 6.110 -2.050 6.310 -1.480 ;
        RECT 6.840 -1.490 7.050 -1.460 ;
        RECT 6.830 -2.080 7.050 -1.490 ;
        RECT 2.620 -3.680 4.570 -2.510 ;
        RECT 4.980 -2.610 5.300 -2.600 ;
        RECT 4.980 -2.780 5.560 -2.610 ;
        RECT 4.980 -2.820 5.310 -2.780 ;
        RECT 4.980 -2.860 5.300 -2.820 ;
        RECT 6.110 -3.110 6.310 -2.540 ;
        RECT 6.830 -3.100 7.050 -2.510 ;
        RECT 6.840 -3.130 7.050 -3.100 ;
        RECT 4.980 -3.180 5.300 -3.150 ;
        RECT 4.980 -3.230 5.310 -3.180 ;
        RECT 4.980 -3.400 5.560 -3.230 ;
        RECT 4.980 -3.410 5.300 -3.400 ;
        RECT 6.840 -3.480 7.040 -3.130 ;
      LAYER mcon ;
        RECT 3.110 1.780 3.280 1.950 ;
        RECT 3.110 1.440 3.280 1.610 ;
        RECT 5.040 1.610 5.210 1.780 ;
        RECT 6.120 1.320 6.290 1.490 ;
        RECT 3.110 1.100 3.280 1.270 ;
        RECT 5.040 1.060 5.210 1.230 ;
        RECT 6.850 1.350 7.020 1.520 ;
        RECT 3.110 0.250 3.280 0.420 ;
        RECT 5.040 0.190 5.210 0.360 ;
        RECT 3.110 -0.090 3.280 0.080 ;
        RECT 6.120 -0.070 6.290 0.100 ;
        RECT 6.850 -0.100 7.020 0.070 ;
        RECT 3.110 -0.430 3.280 -0.260 ;
        RECT 5.040 -0.360 5.210 -0.190 ;
        RECT -2.210 -0.940 -1.940 -0.670 ;
        RECT 6.490 -0.880 6.670 -0.710 ;
        RECT 3.100 -1.310 3.270 -1.140 ;
        RECT 5.040 -1.400 5.210 -1.230 ;
        RECT 3.100 -1.650 3.270 -1.480 ;
        RECT 6.120 -1.690 6.290 -1.520 ;
        RECT 3.100 -1.990 3.270 -1.820 ;
        RECT 5.040 -1.950 5.210 -1.780 ;
        RECT 6.850 -1.660 7.020 -1.490 ;
        RECT 3.100 -2.850 3.270 -2.680 ;
        RECT 5.040 -2.810 5.210 -2.640 ;
        RECT 3.100 -3.190 3.270 -3.020 ;
        RECT 6.120 -3.070 6.290 -2.900 ;
        RECT 6.850 -3.100 7.020 -2.930 ;
        RECT 3.100 -3.530 3.270 -3.360 ;
        RECT 5.040 -3.360 5.210 -3.190 ;
      LAYER met1 ;
        RECT -2.280 -3.820 -1.880 2.170 ;
        RECT 3.070 1.530 3.330 2.010 ;
        RECT 4.970 1.540 5.290 1.860 ;
        RECT 6.110 1.550 6.270 2.230 ;
        RECT 6.110 1.530 6.310 1.550 ;
        RECT 3.060 1.010 3.330 1.530 ;
        RECT 3.060 0.560 3.320 1.010 ;
        RECT 4.970 0.990 5.290 1.310 ;
        RECT 6.090 1.290 6.320 1.530 ;
        RECT 6.110 1.070 6.310 1.290 ;
        RECT 6.480 1.240 6.670 2.230 ;
        RECT 6.920 1.580 7.080 2.230 ;
        RECT 6.500 1.120 6.670 1.240 ;
        RECT 3.070 0.000 3.330 0.480 ;
        RECT 4.970 0.110 5.290 0.430 ;
        RECT 6.110 0.350 6.270 1.070 ;
        RECT 6.110 0.130 6.310 0.350 ;
        RECT 6.510 0.300 6.670 1.120 ;
        RECT 6.810 1.030 7.080 1.580 ;
        RECT 6.810 0.980 7.090 1.030 ;
        RECT 6.920 0.890 7.090 0.980 ;
        RECT 6.920 0.530 7.080 0.890 ;
        RECT 6.920 0.440 7.090 0.530 ;
        RECT 6.500 0.180 6.670 0.300 ;
        RECT 3.060 -0.520 3.330 0.000 ;
        RECT 6.090 -0.110 6.320 0.130 ;
        RECT 4.970 -0.440 5.290 -0.120 ;
        RECT 6.110 -0.130 6.310 -0.110 ;
        RECT 3.060 -0.970 3.320 -0.520 ;
        RECT 3.060 -1.560 3.320 -1.080 ;
        RECT 4.970 -1.470 5.290 -1.150 ;
        RECT 6.110 -1.460 6.270 -0.130 ;
        RECT 6.480 -0.680 6.670 0.180 ;
        RECT 6.810 0.390 7.090 0.440 ;
        RECT 6.810 -0.160 7.080 0.390 ;
        RECT 6.460 -0.910 6.700 -0.680 ;
        RECT 6.110 -1.480 6.310 -1.460 ;
        RECT 3.050 -2.080 3.320 -1.560 ;
        RECT 4.970 -2.020 5.290 -1.700 ;
        RECT 6.090 -1.720 6.320 -1.480 ;
        RECT 6.110 -1.940 6.310 -1.720 ;
        RECT 6.480 -1.770 6.670 -0.910 ;
        RECT 6.920 -1.430 7.080 -0.160 ;
        RECT 6.500 -1.890 6.670 -1.770 ;
        RECT 3.050 -2.530 3.310 -2.080 ;
        RECT 3.060 -3.100 3.320 -2.620 ;
        RECT 4.970 -2.890 5.290 -2.570 ;
        RECT 6.110 -2.650 6.270 -1.940 ;
        RECT 6.110 -2.870 6.310 -2.650 ;
        RECT 6.510 -2.700 6.670 -1.890 ;
        RECT 6.810 -1.980 7.080 -1.430 ;
        RECT 6.810 -2.030 7.090 -1.980 ;
        RECT 6.920 -2.120 7.090 -2.030 ;
        RECT 6.920 -2.470 7.080 -2.120 ;
        RECT 6.920 -2.560 7.090 -2.470 ;
        RECT 6.500 -2.820 6.670 -2.700 ;
        RECT 3.050 -3.620 3.320 -3.100 ;
        RECT 6.090 -3.110 6.320 -2.870 ;
        RECT 4.970 -3.440 5.290 -3.120 ;
        RECT 6.110 -3.130 6.310 -3.110 ;
        RECT 3.050 -4.070 3.310 -3.620 ;
        RECT 6.110 -3.810 6.270 -3.130 ;
        RECT 6.480 -3.810 6.670 -2.820 ;
        RECT 6.810 -2.610 7.090 -2.560 ;
        RECT 6.810 -3.160 7.080 -2.610 ;
        RECT 6.920 -3.810 7.080 -3.160 ;
      LAYER via ;
        RECT 5.000 1.570 5.260 1.830 ;
        RECT 5.000 1.020 5.260 1.280 ;
        RECT 5.000 0.140 5.260 0.400 ;
        RECT 5.000 -0.410 5.260 -0.150 ;
        RECT 5.000 -1.440 5.260 -1.180 ;
        RECT 5.000 -1.990 5.260 -1.730 ;
        RECT 5.000 -2.860 5.260 -2.600 ;
        RECT 5.000 -3.410 5.260 -3.150 ;
      LAYER met2 ;
        RECT 4.970 1.730 5.280 1.870 ;
        RECT -2.640 1.550 7.440 1.730 ;
        RECT 4.970 1.540 5.280 1.550 ;
        RECT 4.970 1.300 5.280 1.320 ;
        RECT -2.640 1.120 7.440 1.300 ;
        RECT 4.970 0.990 5.280 1.120 ;
        RECT 4.970 0.300 5.280 0.430 ;
        RECT -2.640 0.120 7.440 0.300 ;
        RECT 4.970 0.100 5.280 0.120 ;
        RECT 4.970 -0.130 5.280 -0.120 ;
        RECT -2.640 -0.200 4.960 -0.130 ;
        RECT 4.970 -0.200 7.440 -0.130 ;
        RECT -2.640 -0.310 7.440 -0.200 ;
        RECT 4.970 -0.450 5.280 -0.310 ;
        RECT 4.970 -1.280 5.280 -1.140 ;
        RECT 4.970 -1.290 7.440 -1.280 ;
        RECT -2.620 -1.460 7.440 -1.290 ;
        RECT 4.970 -1.470 5.280 -1.460 ;
        RECT 4.970 -1.710 5.280 -1.690 ;
        RECT -2.620 -1.880 7.440 -1.710 ;
        RECT 4.880 -1.890 7.440 -1.880 ;
        RECT 4.970 -2.020 5.280 -1.890 ;
        RECT 4.970 -2.690 5.280 -2.570 ;
        RECT -2.620 -2.700 5.280 -2.690 ;
        RECT -2.620 -2.860 7.440 -2.700 ;
        RECT -1.840 -2.950 -0.300 -2.860 ;
        RECT 4.880 -2.880 7.440 -2.860 ;
        RECT 4.970 -2.900 5.280 -2.880 ;
        RECT 4.970 -3.130 5.280 -3.120 ;
        RECT -2.620 -3.300 7.440 -3.130 ;
        RECT 4.970 -3.310 7.440 -3.300 ;
        RECT 4.970 -3.450 5.280 -3.310 ;
  END
END sky130_hilas_swc4x1cellOverlap

MACRO sky130_hilas_Tgate4Single01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_Tgate4Single01 ;
  ORIGIN 0.360 1.410 ;
  SIZE 4.760 BY 6.050 ;
  PIN INPUT1_4
    USE ANALOG ;
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER li1 ;
        RECT 1.420 -1.010 1.590 -0.850 ;
        RECT 2.920 -1.010 3.090 -0.850 ;
        RECT 1.290 -1.050 1.610 -1.010 ;
        RECT 2.860 -1.050 3.180 -1.010 ;
        RECT 1.290 -1.240 1.620 -1.050 ;
        RECT 2.860 -1.240 3.190 -1.050 ;
        RECT 1.290 -1.270 1.610 -1.240 ;
        RECT 2.860 -1.270 3.180 -1.240 ;
      LAYER mcon ;
        RECT 1.350 -1.230 1.520 -1.060 ;
        RECT 2.920 -1.230 3.090 -1.060 ;
      LAYER met1 ;
        RECT 1.280 -1.300 1.600 -0.980 ;
        RECT 2.850 -1.300 3.170 -0.980 ;
      LAYER via ;
        RECT 1.310 -1.270 1.570 -1.010 ;
        RECT 2.880 -1.270 3.140 -1.010 ;
      LAYER met2 ;
        RECT 1.280 -1.090 1.590 -0.970 ;
        RECT 0.510 -1.100 1.630 -1.090 ;
        RECT 2.850 -1.100 3.160 -0.970 ;
        RECT -0.360 -1.300 3.160 -1.100 ;
        RECT 0.510 -1.310 1.630 -1.300 ;
    END
  END INPUT1_4
  PIN VPWR
    USE ANALOG ;
    ANTENNADIFFAREA 0.908800 ;
    PORT
      LAYER nwell ;
        RECT -0.240 -1.410 2.520 4.640 ;
      LAYER li1 ;
        RECT 0.070 4.130 0.240 4.410 ;
        RECT 0.070 4.090 0.280 4.130 ;
        RECT 0.070 4.070 0.300 4.090 ;
        RECT 0.070 4.050 0.330 4.070 ;
        RECT 0.070 4.000 0.410 4.050 ;
        RECT 0.070 3.940 0.560 4.000 ;
        RECT 0.070 3.910 0.580 3.940 ;
        RECT 0.110 3.880 0.580 3.910 ;
        RECT 0.240 3.830 0.580 3.880 ;
        RECT 0.360 3.820 0.580 3.830 ;
        RECT 0.370 3.790 0.580 3.820 ;
        RECT 0.390 3.710 0.580 3.790 ;
        RECT 0.390 3.540 0.910 3.710 ;
        RECT 0.390 3.510 0.580 3.540 ;
        RECT 0.390 2.710 0.580 2.740 ;
        RECT 0.390 2.540 0.910 2.710 ;
        RECT 0.390 2.460 0.580 2.540 ;
        RECT 0.370 2.430 0.580 2.460 ;
        RECT 0.360 2.420 0.580 2.430 ;
        RECT 0.240 2.370 0.580 2.420 ;
        RECT 0.110 2.340 0.580 2.370 ;
        RECT 0.070 2.310 0.580 2.340 ;
        RECT 0.070 2.250 0.560 2.310 ;
        RECT 0.070 2.200 0.410 2.250 ;
        RECT 0.070 2.180 0.330 2.200 ;
        RECT 0.070 2.160 0.300 2.180 ;
        RECT 0.070 2.120 0.280 2.160 ;
        RECT 0.070 1.840 0.240 2.120 ;
        RECT 0.070 1.110 0.240 1.390 ;
        RECT 0.070 1.070 0.280 1.110 ;
        RECT 0.070 1.050 0.300 1.070 ;
        RECT 0.070 1.030 0.330 1.050 ;
        RECT 0.070 0.980 0.410 1.030 ;
        RECT 0.070 0.920 0.560 0.980 ;
        RECT 0.070 0.890 0.580 0.920 ;
        RECT 0.110 0.860 0.580 0.890 ;
        RECT 0.240 0.810 0.580 0.860 ;
        RECT 0.360 0.800 0.580 0.810 ;
        RECT 0.370 0.770 0.580 0.800 ;
        RECT 0.390 0.690 0.580 0.770 ;
        RECT 0.390 0.520 0.910 0.690 ;
        RECT 0.390 0.490 0.580 0.520 ;
        RECT 0.390 -0.310 0.580 -0.280 ;
        RECT 0.390 -0.480 0.910 -0.310 ;
        RECT 0.390 -0.560 0.580 -0.480 ;
        RECT 0.370 -0.590 0.580 -0.560 ;
        RECT 0.360 -0.600 0.580 -0.590 ;
        RECT 0.240 -0.650 0.580 -0.600 ;
        RECT 0.110 -0.680 0.580 -0.650 ;
        RECT 0.070 -0.710 0.580 -0.680 ;
        RECT 0.070 -0.770 0.560 -0.710 ;
        RECT 0.070 -0.820 0.410 -0.770 ;
        RECT 0.070 -0.840 0.330 -0.820 ;
        RECT 0.070 -0.860 0.300 -0.840 ;
        RECT 0.070 -0.900 0.280 -0.860 ;
        RECT 0.070 -1.180 0.240 -0.900 ;
      LAYER mcon ;
        RECT 0.400 3.540 0.570 3.710 ;
        RECT 0.400 2.540 0.570 2.710 ;
        RECT 0.400 0.520 0.570 0.690 ;
        RECT 0.400 -0.480 0.570 -0.310 ;
      LAYER met1 ;
        RECT 0.380 3.770 0.580 4.640 ;
        RECT 0.370 3.480 0.600 3.770 ;
        RECT 0.380 2.770 0.580 3.480 ;
        RECT 0.370 2.480 0.600 2.770 ;
        RECT 0.380 0.750 0.580 2.480 ;
        RECT 0.370 0.460 0.600 0.750 ;
        RECT 0.380 -0.250 0.580 0.460 ;
        RECT 0.370 -0.540 0.600 -0.250 ;
        RECT 0.380 -1.410 0.580 -0.540 ;
    END
  END VPWR
  PIN SELECT4
    USE ANALOG ;
    ANTENNAGATEAREA 0.372000 ;
    PORT
      LAYER li1 ;
        RECT -0.120 -0.430 0.090 0.000 ;
        RECT -0.100 -0.450 0.070 -0.430 ;
      LAYER met1 ;
        RECT -0.120 -0.220 0.220 0.000 ;
        RECT -0.130 -0.320 0.220 -0.220 ;
        RECT -0.130 -0.510 0.100 -0.320 ;
      LAYER via ;
        RECT -0.040 -0.290 0.220 -0.030 ;
      LAYER met2 ;
        RECT -0.070 -0.120 0.250 -0.030 ;
        RECT -0.360 -0.320 0.250 -0.120 ;
    END
  END SELECT4
  PIN SELECT3
    USE ANALOG ;
    ANTENNAGATEAREA 0.372000 ;
    PORT
      LAYER li1 ;
        RECT -0.100 0.640 0.070 0.660 ;
        RECT -0.120 0.210 0.090 0.640 ;
      LAYER mcon ;
        RECT -0.100 0.490 0.070 0.660 ;
      LAYER met1 ;
        RECT -0.130 0.530 0.100 0.720 ;
        RECT -0.130 0.430 0.220 0.530 ;
        RECT -0.120 0.210 0.220 0.430 ;
      LAYER via ;
        RECT -0.040 0.240 0.220 0.500 ;
      LAYER met2 ;
        RECT -0.360 0.330 0.250 0.530 ;
        RECT -0.070 0.240 0.250 0.330 ;
    END
  END SELECT3
  PIN INPUT1_3
    USE ANALOG ;
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER li1 ;
        RECT 1.290 1.450 1.610 1.480 ;
        RECT 2.860 1.450 3.180 1.480 ;
        RECT 1.290 1.260 1.620 1.450 ;
        RECT 2.860 1.260 3.190 1.450 ;
        RECT 1.290 1.220 1.610 1.260 ;
        RECT 2.860 1.220 3.180 1.260 ;
        RECT 1.420 1.060 1.590 1.220 ;
        RECT 2.920 1.060 3.090 1.220 ;
      LAYER mcon ;
        RECT 1.350 1.270 1.520 1.440 ;
        RECT 2.920 1.270 3.090 1.440 ;
      LAYER met1 ;
        RECT 1.280 1.190 1.600 1.510 ;
        RECT 2.850 1.190 3.170 1.510 ;
      LAYER via ;
        RECT 1.310 1.220 1.570 1.480 ;
        RECT 2.880 1.220 3.140 1.480 ;
      LAYER met2 ;
        RECT 0.510 1.510 1.630 1.520 ;
        RECT -0.360 1.310 3.160 1.510 ;
        RECT 0.510 1.300 1.630 1.310 ;
        RECT 1.280 1.180 1.590 1.300 ;
        RECT 2.850 1.180 3.160 1.310 ;
    END
  END INPUT1_3
  PIN INPUT1_2
    USE ANALOG ;
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER li1 ;
        RECT 1.420 2.010 1.590 2.170 ;
        RECT 2.920 2.010 3.090 2.170 ;
        RECT 1.290 1.970 1.610 2.010 ;
        RECT 2.860 1.970 3.180 2.010 ;
        RECT 1.290 1.780 1.620 1.970 ;
        RECT 2.860 1.780 3.190 1.970 ;
        RECT 1.290 1.750 1.610 1.780 ;
        RECT 2.860 1.750 3.180 1.780 ;
      LAYER mcon ;
        RECT 1.350 1.790 1.520 1.960 ;
        RECT 2.920 1.790 3.090 1.960 ;
      LAYER met1 ;
        RECT 1.280 1.720 1.600 2.040 ;
        RECT 2.850 1.720 3.170 2.040 ;
      LAYER via ;
        RECT 1.310 1.750 1.570 2.010 ;
        RECT 2.880 1.750 3.140 2.010 ;
      LAYER met2 ;
        RECT 1.280 1.930 1.590 2.050 ;
        RECT 0.510 1.920 1.630 1.930 ;
        RECT 2.850 1.920 3.160 2.050 ;
        RECT -0.360 1.720 3.160 1.920 ;
        RECT 0.510 1.710 1.630 1.720 ;
    END
  END INPUT1_2
  PIN SELECT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.372000 ;
    PORT
      LAYER li1 ;
        RECT -0.120 2.590 0.090 3.020 ;
        RECT -0.100 2.570 0.070 2.590 ;
      LAYER met1 ;
        RECT -0.120 2.800 0.220 3.020 ;
        RECT -0.130 2.700 0.220 2.800 ;
        RECT -0.130 2.510 0.100 2.700 ;
      LAYER via ;
        RECT -0.040 2.730 0.220 2.990 ;
      LAYER met2 ;
        RECT -0.070 2.900 0.250 2.990 ;
        RECT -0.360 2.700 0.250 2.900 ;
    END
  END SELECT2
  PIN SELECT1
    USE ANALOG ;
    ANTENNAGATEAREA 0.372000 ;
    PORT
      LAYER li1 ;
        RECT -0.100 3.660 0.070 3.680 ;
        RECT -0.120 3.230 0.090 3.660 ;
      LAYER mcon ;
        RECT -0.100 3.510 0.070 3.680 ;
      LAYER met1 ;
        RECT -0.130 3.550 0.100 3.740 ;
        RECT -0.130 3.450 0.220 3.550 ;
        RECT -0.120 3.230 0.220 3.450 ;
      LAYER via ;
        RECT -0.040 3.260 0.220 3.520 ;
      LAYER met2 ;
        RECT -0.360 3.350 0.250 3.550 ;
        RECT -0.070 3.260 0.250 3.350 ;
    END
  END SELECT1
  PIN INPUT1_1
    USE ANALOG ;
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER li1 ;
        RECT 1.290 4.470 1.610 4.500 ;
        RECT 2.860 4.470 3.180 4.500 ;
        RECT 1.290 4.280 1.620 4.470 ;
        RECT 2.860 4.280 3.190 4.470 ;
        RECT 1.290 4.240 1.610 4.280 ;
        RECT 2.860 4.240 3.180 4.280 ;
        RECT 1.420 4.080 1.590 4.240 ;
        RECT 2.920 4.080 3.090 4.240 ;
      LAYER mcon ;
        RECT 1.350 4.290 1.520 4.460 ;
        RECT 2.920 4.290 3.090 4.460 ;
      LAYER met1 ;
        RECT 1.280 4.210 1.600 4.530 ;
        RECT 2.850 4.210 3.170 4.530 ;
      LAYER via ;
        RECT 1.310 4.240 1.570 4.500 ;
        RECT 2.880 4.240 3.140 4.500 ;
      LAYER met2 ;
        RECT 0.510 4.530 1.630 4.540 ;
        RECT -0.360 4.330 3.160 4.530 ;
        RECT 0.510 4.320 1.630 4.330 ;
        RECT 1.280 4.200 1.590 4.320 ;
        RECT 2.850 4.200 3.160 4.330 ;
    END
  END INPUT1_1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 4.150 3.740 4.320 4.420 ;
        RECT 3.890 3.700 4.320 3.740 ;
        RECT 3.540 3.540 4.320 3.700 ;
        RECT 3.540 3.530 4.080 3.540 ;
        RECT 3.890 3.510 4.080 3.530 ;
        RECT 3.890 2.720 4.080 2.740 ;
        RECT 3.540 2.710 4.080 2.720 ;
        RECT 3.540 2.550 4.320 2.710 ;
        RECT 3.890 2.510 4.320 2.550 ;
        RECT 4.150 1.830 4.320 2.510 ;
        RECT 4.150 0.720 4.320 1.400 ;
        RECT 3.890 0.680 4.320 0.720 ;
        RECT 3.540 0.520 4.320 0.680 ;
        RECT 3.540 0.510 4.080 0.520 ;
        RECT 3.890 0.490 4.080 0.510 ;
        RECT 3.890 -0.300 4.080 -0.280 ;
        RECT 3.540 -0.310 4.080 -0.300 ;
        RECT 3.540 -0.470 4.320 -0.310 ;
        RECT 3.890 -0.510 4.320 -0.470 ;
        RECT 4.150 -1.190 4.320 -0.510 ;
      LAYER mcon ;
        RECT 3.900 3.540 4.070 3.710 ;
        RECT 3.900 2.540 4.070 2.710 ;
        RECT 3.900 0.520 4.070 0.690 ;
        RECT 3.900 -0.480 4.070 -0.310 ;
      LAYER met1 ;
        RECT 3.890 3.770 4.080 4.640 ;
        RECT 3.870 3.480 4.100 3.770 ;
        RECT 3.890 2.770 4.080 3.480 ;
        RECT 3.870 2.480 4.100 2.770 ;
        RECT 3.890 0.750 4.080 2.480 ;
        RECT 3.870 0.460 4.100 0.750 ;
        RECT 3.890 -0.250 4.080 0.460 ;
        RECT 3.870 -0.540 4.100 -0.250 ;
        RECT 3.890 -1.410 4.080 -0.540 ;
    END
  END VGND
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.182900 ;
    PORT
      LAYER li1 ;
        RECT 2.300 4.330 2.490 4.350 ;
        RECT 2.030 4.160 2.490 4.330 ;
        RECT 2.280 4.150 2.490 4.160 ;
        RECT 2.300 4.120 2.490 4.150 ;
        RECT 3.430 4.330 3.620 4.360 ;
        RECT 3.430 4.160 3.870 4.330 ;
        RECT 3.430 4.130 3.620 4.160 ;
      LAYER mcon ;
        RECT 2.310 4.150 2.480 4.320 ;
        RECT 3.440 4.160 3.610 4.330 ;
      LAYER met1 ;
        RECT 2.280 4.090 2.510 4.380 ;
        RECT 3.410 4.100 3.640 4.390 ;
        RECT 2.300 3.620 2.490 4.090 ;
        RECT 2.230 3.300 2.490 3.620 ;
        RECT 3.410 3.610 3.600 4.100 ;
        RECT 3.240 3.360 3.600 3.610 ;
        RECT 3.240 3.290 3.500 3.360 ;
      LAYER via ;
        RECT 2.230 3.330 2.490 3.590 ;
        RECT 3.240 3.320 3.500 3.580 ;
      LAYER met2 ;
        RECT 2.200 3.550 2.520 3.590 ;
        RECT 3.210 3.550 3.530 3.580 ;
        RECT 2.150 3.350 4.400 3.550 ;
        RECT 2.200 3.330 2.520 3.350 ;
        RECT 3.210 3.320 3.530 3.350 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.182900 ;
    PORT
      LAYER li1 ;
        RECT 2.300 2.100 2.490 2.130 ;
        RECT 2.280 2.090 2.490 2.100 ;
        RECT 2.030 1.920 2.490 2.090 ;
        RECT 2.300 1.900 2.490 1.920 ;
        RECT 3.430 2.090 3.620 2.120 ;
        RECT 3.430 1.920 3.870 2.090 ;
        RECT 3.430 1.890 3.620 1.920 ;
      LAYER mcon ;
        RECT 2.310 1.930 2.480 2.100 ;
        RECT 3.440 1.920 3.610 2.090 ;
      LAYER met1 ;
        RECT 2.230 2.630 2.490 2.950 ;
        RECT 3.240 2.890 3.500 2.960 ;
        RECT 3.240 2.640 3.600 2.890 ;
        RECT 2.300 2.160 2.490 2.630 ;
        RECT 2.280 1.870 2.510 2.160 ;
        RECT 3.410 2.150 3.600 2.640 ;
        RECT 3.410 1.860 3.640 2.150 ;
      LAYER via ;
        RECT 2.230 2.660 2.490 2.920 ;
        RECT 3.240 2.670 3.500 2.930 ;
      LAYER met2 ;
        RECT 2.200 2.900 2.520 2.920 ;
        RECT 3.210 2.900 3.530 2.930 ;
        RECT 2.150 2.700 4.400 2.900 ;
        RECT 2.200 2.660 2.520 2.700 ;
        RECT 3.210 2.670 3.530 2.700 ;
    END
  END OUTPUT2
  PIN OUTPUT3
    USE ANALOG ;
    ANTENNADIFFAREA 0.182900 ;
    PORT
      LAYER li1 ;
        RECT 2.300 1.310 2.490 1.330 ;
        RECT 2.030 1.140 2.490 1.310 ;
        RECT 2.280 1.130 2.490 1.140 ;
        RECT 2.300 1.100 2.490 1.130 ;
        RECT 3.430 1.310 3.620 1.340 ;
        RECT 3.430 1.140 3.870 1.310 ;
        RECT 3.430 1.110 3.620 1.140 ;
      LAYER mcon ;
        RECT 2.310 1.130 2.480 1.300 ;
        RECT 3.440 1.140 3.610 1.310 ;
      LAYER met1 ;
        RECT 2.280 1.070 2.510 1.360 ;
        RECT 3.410 1.080 3.640 1.370 ;
        RECT 2.300 0.600 2.490 1.070 ;
        RECT 2.230 0.280 2.490 0.600 ;
        RECT 3.410 0.590 3.600 1.080 ;
        RECT 3.240 0.340 3.600 0.590 ;
        RECT 3.240 0.270 3.500 0.340 ;
      LAYER via ;
        RECT 2.230 0.310 2.490 0.570 ;
        RECT 3.240 0.300 3.500 0.560 ;
      LAYER met2 ;
        RECT 2.200 0.530 2.520 0.570 ;
        RECT 3.210 0.530 3.530 0.560 ;
        RECT 2.150 0.330 4.400 0.530 ;
        RECT 2.200 0.310 2.520 0.330 ;
        RECT 3.210 0.300 3.530 0.330 ;
    END
  END OUTPUT3
  PIN OUTPUT4
    USE ANALOG ;
    ANTENNADIFFAREA 0.182900 ;
    PORT
      LAYER li1 ;
        RECT 2.300 -0.920 2.490 -0.890 ;
        RECT 2.280 -0.930 2.490 -0.920 ;
        RECT 2.030 -1.100 2.490 -0.930 ;
        RECT 2.300 -1.120 2.490 -1.100 ;
        RECT 3.430 -0.930 3.620 -0.900 ;
        RECT 3.430 -1.100 3.870 -0.930 ;
        RECT 3.430 -1.130 3.620 -1.100 ;
      LAYER mcon ;
        RECT 2.310 -1.090 2.480 -0.920 ;
        RECT 3.440 -1.100 3.610 -0.930 ;
      LAYER met1 ;
        RECT 2.230 -0.390 2.490 -0.070 ;
        RECT 3.240 -0.130 3.500 -0.060 ;
        RECT 3.240 -0.380 3.600 -0.130 ;
        RECT 2.300 -0.860 2.490 -0.390 ;
        RECT 2.280 -1.150 2.510 -0.860 ;
        RECT 3.410 -0.870 3.600 -0.380 ;
        RECT 3.410 -1.160 3.640 -0.870 ;
      LAYER via ;
        RECT 2.230 -0.360 2.490 -0.100 ;
        RECT 3.240 -0.350 3.500 -0.090 ;
      LAYER met2 ;
        RECT 2.200 -0.120 2.520 -0.100 ;
        RECT 3.210 -0.120 3.530 -0.090 ;
        RECT 2.150 -0.320 4.400 -0.120 ;
        RECT 2.200 -0.360 2.520 -0.320 ;
        RECT 3.210 -0.350 3.530 -0.320 ;
    END
  END OUTPUT4
  OBS
      LAYER li1 ;
        RECT 1.750 3.710 2.080 3.830 ;
        RECT 1.260 3.530 3.160 3.710 ;
        RECT 1.260 2.540 3.160 2.720 ;
        RECT 1.750 2.420 2.080 2.540 ;
        RECT 1.750 0.690 2.080 0.810 ;
        RECT 1.260 0.510 3.160 0.690 ;
        RECT 1.260 -0.480 3.160 -0.300 ;
        RECT 1.750 -0.600 2.080 -0.480 ;
  END
END sky130_hilas_Tgate4Single01

MACRO sky130_hilas_nFETLargePart1
  CLASS BLOCK ;
  FOREIGN sky130_hilas_nFETLargePart1 ;
  ORIGIN 1.650 0.310 ;
  SIZE 3.020 BY 2.720 ;
  OBS
      LAYER li1 ;
        RECT -1.600 -0.130 -1.430 2.270 ;
        RECT -1.050 -0.130 -0.880 2.270 ;
        RECT -0.500 -0.130 -0.330 2.270 ;
        RECT 0.050 -0.130 0.220 2.270 ;
        RECT 0.600 -0.130 0.770 2.270 ;
        RECT 1.150 -0.130 1.320 2.270 ;
  END
END sky130_hilas_nFETLargePart1

MACRO sky130_hilas_TA2Cell_1FG
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TA2Cell_1FG ;
  ORIGIN 26.160 -1.400 ;
  SIZE 28.090 BY 6.050 ;
  PIN VINP_AMP1
    USE ANALOG ;
    PORT
      LAYER li1 ;
        RECT -21.560 6.440 -16.500 7.270 ;
        RECT -17.050 6.360 -16.570 6.440 ;
        RECT -17.050 6.110 -16.580 6.360 ;
      LAYER mcon ;
        RECT -16.810 6.150 -16.640 6.320 ;
      LAYER met1 ;
        RECT -16.890 6.080 -16.570 6.400 ;
      LAYER via ;
        RECT -16.860 6.110 -16.600 6.370 ;
      LAYER met2 ;
        RECT -16.880 6.370 -16.570 6.410 ;
        RECT -17.260 6.350 -16.420 6.370 ;
        RECT -17.260 6.170 -14.630 6.350 ;
        RECT -16.880 6.080 -16.570 6.170 ;
    END
  END VINP_AMP1
  PIN VINP_AMP2
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER li1 ;
        RECT -2.190 4.730 -1.870 4.760 ;
        RECT -2.190 4.540 -1.860 4.730 ;
        RECT -2.190 4.500 -1.870 4.540 ;
        RECT -2.190 4.420 -2.020 4.500 ;
        RECT -2.240 4.250 -2.020 4.420 ;
        RECT -2.240 4.090 -2.070 4.250 ;
      LAYER mcon ;
        RECT -2.130 4.550 -1.960 4.720 ;
      LAYER met1 ;
        RECT -2.200 4.470 -1.880 4.790 ;
      LAYER via ;
        RECT -2.170 4.500 -1.910 4.760 ;
      LAYER met2 ;
        RECT -2.200 4.750 -1.890 4.790 ;
        RECT -2.520 4.740 -1.860 4.750 ;
        RECT -2.520 4.510 -1.420 4.740 ;
        RECT -2.200 4.460 -1.890 4.510 ;
    END
  END VINP_AMP2
  PIN VINN_AMP2
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER li1 ;
        RECT -2.220 7.400 -2.050 7.450 ;
        RECT -2.220 7.140 -1.660 7.400 ;
        RECT -2.220 7.120 -2.050 7.140 ;
      LAYER mcon ;
        RECT -1.890 7.180 -1.720 7.350 ;
      LAYER met1 ;
        RECT -1.970 7.110 -1.650 7.430 ;
      LAYER via ;
        RECT -1.940 7.140 -1.680 7.400 ;
      LAYER met2 ;
        RECT -1.960 7.430 -1.650 7.440 ;
        RECT -2.530 7.420 -1.650 7.430 ;
        RECT -2.600 7.180 -1.650 7.420 ;
        RECT -1.960 7.110 -1.650 7.180 ;
    END
  END VINN_AMP2
  PIN GATECOLSELECT
    USE ANALOG ;
    ANTENNAGATEAREA 0.310000 ;
    PORT
      LAYER li1 ;
        RECT -4.160 5.980 -3.970 5.990 ;
        RECT -4.160 5.690 -3.960 5.980 ;
        RECT -4.170 5.360 -3.930 5.690 ;
        RECT -4.170 3.160 -3.930 3.490 ;
        RECT -4.160 2.870 -3.960 3.160 ;
        RECT -4.160 2.860 -3.970 2.870 ;
      LAYER mcon ;
        RECT -4.150 5.730 -3.970 5.920 ;
        RECT -4.150 2.930 -3.970 3.120 ;
      LAYER met1 ;
        RECT -4.160 5.990 -3.970 7.450 ;
        RECT -4.160 5.960 -3.940 5.990 ;
        RECT -4.180 5.690 -3.930 5.960 ;
        RECT -4.170 5.680 -3.930 5.690 ;
        RECT -4.170 5.440 -3.940 5.680 ;
        RECT -4.130 3.410 -3.970 5.440 ;
        RECT -4.170 3.170 -3.940 3.410 ;
        RECT -4.170 3.160 -3.930 3.170 ;
        RECT -4.180 2.890 -3.930 3.160 ;
        RECT -4.160 2.860 -3.940 2.890 ;
        RECT -4.160 1.400 -3.970 2.860 ;
    END
  END GATECOLSELECT
  PIN VPWR
    USE ANALOG ;
    ANTENNADIFFAREA 1.373600 ;
    PORT
      LAYER nwell ;
        RECT 0.650 1.400 1.930 7.450 ;
      LAYER li1 ;
        RECT 0.860 5.840 1.560 6.150 ;
        RECT 0.710 5.610 1.560 5.840 ;
        RECT 0.860 5.270 1.560 5.610 ;
        RECT 0.860 3.250 1.560 3.590 ;
        RECT 0.710 3.020 1.560 3.250 ;
        RECT 0.860 2.710 1.560 3.020 ;
      LAYER mcon ;
        RECT 0.720 5.640 0.890 5.810 ;
        RECT 0.720 3.050 0.890 3.220 ;
      LAYER met1 ;
        RECT 0.630 7.300 0.910 7.450 ;
        RECT 0.640 5.870 0.910 7.300 ;
        RECT 0.640 5.580 0.920 5.870 ;
        RECT 0.640 3.280 0.910 5.580 ;
        RECT 0.640 2.990 0.920 3.280 ;
        RECT 0.640 1.400 0.910 2.990 ;
    END
  END VPWR
  PIN VGND
    USE ANALOG ;
    ANTENNADIFFAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT -0.160 6.170 0.390 7.160 ;
        RECT -0.160 4.690 0.390 5.680 ;
        RECT -0.160 3.210 0.390 4.200 ;
        RECT -0.160 1.730 0.390 2.720 ;
      LAYER mcon ;
        RECT 0.060 6.580 0.230 6.750 ;
        RECT 0.060 5.100 0.230 5.270 ;
        RECT 0.060 3.620 0.230 3.790 ;
        RECT 0.060 2.140 0.230 2.310 ;
      LAYER met1 ;
        RECT -0.030 1.400 0.310 7.450 ;
    END
  END VGND
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -6.510 7.440 -3.200 7.450 ;
        RECT -6.510 1.410 -1.350 7.440 ;
        RECT -3.210 1.400 -1.350 1.410 ;
      LAYER li1 ;
        RECT -3.800 6.770 -3.600 7.120 ;
        RECT -3.800 6.740 -3.590 6.770 ;
        RECT -4.530 4.880 -4.360 6.490 ;
        RECT -3.810 6.160 -3.590 6.740 ;
        RECT -3.800 6.150 -3.590 6.160 ;
        RECT -4.530 4.690 -4.350 4.880 ;
        RECT -4.530 3.970 -4.350 4.160 ;
        RECT -4.530 2.360 -4.360 3.970 ;
        RECT -3.800 2.690 -3.590 2.700 ;
        RECT -3.810 2.110 -3.590 2.690 ;
        RECT -3.800 2.080 -3.590 2.110 ;
        RECT -3.800 1.730 -3.600 2.080 ;
      LAYER mcon ;
        RECT -3.790 6.570 -3.620 6.740 ;
        RECT -3.790 2.110 -3.620 2.280 ;
      LAYER met1 ;
        RECT -3.720 6.800 -3.440 7.450 ;
        RECT -3.830 6.200 -3.440 6.800 ;
        RECT -4.560 4.880 -4.320 5.010 ;
        RECT -4.560 4.560 -4.300 4.880 ;
        RECT -3.720 4.600 -3.440 6.200 ;
        RECT -3.720 4.280 -3.360 4.600 ;
        RECT -4.560 3.960 -4.300 4.280 ;
        RECT -4.560 3.840 -4.320 3.960 ;
        RECT -3.720 2.650 -3.440 4.280 ;
        RECT -3.830 2.050 -3.440 2.650 ;
        RECT -3.720 1.400 -3.440 2.050 ;
      LAYER via ;
        RECT -4.560 4.590 -4.300 4.850 ;
        RECT -3.620 4.310 -3.360 4.570 ;
        RECT -4.560 3.990 -4.300 4.250 ;
      LAYER met2 ;
        RECT -4.590 4.590 -4.270 4.850 ;
        RECT -4.550 4.570 -3.370 4.590 ;
        RECT -4.550 4.310 -3.330 4.570 ;
        RECT -4.550 4.250 -3.370 4.310 ;
        RECT -4.590 4.240 -3.370 4.250 ;
        RECT -4.590 3.990 -4.270 4.240 ;
    END
  END VINJ
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER li1 ;
        RECT -0.750 4.990 -0.550 5.020 ;
        RECT -0.980 4.730 -0.550 4.990 ;
        RECT 1.320 4.910 1.640 4.950 ;
        RECT 1.320 4.850 1.650 4.910 ;
        RECT -0.750 4.690 -0.550 4.730 ;
        RECT 0.850 4.720 1.650 4.850 ;
        RECT 0.850 4.690 1.640 4.720 ;
        RECT 0.850 4.670 1.550 4.690 ;
      LAYER mcon ;
        RECT -0.920 4.780 -0.750 4.950 ;
        RECT 1.380 4.730 1.550 4.900 ;
      LAYER met1 ;
        RECT -0.990 4.700 -0.670 5.020 ;
        RECT 1.310 4.660 1.630 4.980 ;
      LAYER via ;
        RECT -0.960 4.730 -0.700 4.990 ;
        RECT 1.340 4.690 1.600 4.950 ;
      LAYER met2 ;
        RECT -0.990 4.970 -0.680 5.020 ;
        RECT 1.310 4.970 1.620 4.990 ;
        RECT -0.990 4.740 1.930 4.970 ;
        RECT -0.990 4.690 -0.680 4.740 ;
        RECT 1.310 4.660 1.620 4.740 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER li1 ;
        RECT -0.750 4.160 -0.550 4.200 ;
        RECT 1.310 4.190 1.630 4.230 ;
        RECT -0.980 3.900 -0.550 4.160 ;
        RECT 0.850 4.010 1.640 4.190 ;
        RECT 1.310 4.000 1.640 4.010 ;
        RECT 1.310 3.970 1.630 4.000 ;
        RECT -0.750 3.870 -0.550 3.900 ;
      LAYER mcon ;
        RECT -0.920 3.940 -0.750 4.110 ;
        RECT 1.370 4.010 1.540 4.180 ;
      LAYER met1 ;
        RECT -0.990 3.870 -0.670 4.190 ;
        RECT 1.300 3.940 1.620 4.260 ;
      LAYER via ;
        RECT -0.960 3.900 -0.700 4.160 ;
        RECT 1.330 3.970 1.590 4.230 ;
      LAYER met2 ;
        RECT -0.990 4.140 -0.680 4.200 ;
        RECT 1.300 4.140 1.610 4.270 ;
        RECT -0.990 3.920 1.930 4.140 ;
        RECT -0.990 3.870 -0.680 3.920 ;
    END
  END OUTPUT2
  OBS
      LAYER nwell ;
        RECT -26.160 1.410 -22.850 7.440 ;
        RECT -21.120 5.060 -18.400 6.710 ;
        RECT -16.370 6.700 -12.990 7.450 ;
        RECT -21.110 5.020 -18.400 5.060 ;
        RECT -21.110 3.690 -18.400 3.730 ;
        RECT -21.120 2.040 -18.400 3.690 ;
        RECT -16.380 3.130 -12.980 6.700 ;
        RECT -10.960 5.060 -8.240 6.710 ;
        RECT -10.960 5.020 -8.250 5.060 ;
        RECT -10.960 3.690 -8.250 3.730 ;
        RECT -16.370 1.410 -12.990 3.130 ;
        RECT -10.960 2.040 -8.240 3.690 ;
      LAYER li1 ;
        RECT -0.750 7.120 -0.550 7.160 ;
        RECT -25.760 6.770 -25.560 7.120 ;
        RECT -24.280 6.870 -23.750 7.040 ;
        RECT -5.610 6.870 -5.080 7.040 ;
        RECT -25.770 6.740 -25.560 6.770 ;
        RECT -25.770 6.160 -25.550 6.740 ;
        RECT -25.770 6.150 -25.560 6.160 ;
        RECT -25.390 5.980 -25.200 5.990 ;
        RECT -25.400 5.690 -25.200 5.980 ;
        RECT -25.430 5.360 -25.190 5.690 ;
        RECT -25.000 4.880 -24.830 6.490 ;
        RECT -25.010 4.690 -24.830 4.880 ;
        RECT -24.170 5.960 -24.000 6.480 ;
        RECT -23.580 6.290 -23.250 6.460 ;
        RECT -22.230 6.290 -21.880 6.460 ;
        RECT -7.480 6.290 -7.130 6.460 ;
        RECT -6.110 6.290 -5.780 6.460 ;
        RECT -24.170 5.700 -23.840 5.960 ;
        RECT -24.170 4.790 -24.000 5.700 ;
        RECT -23.580 5.500 -23.250 5.670 ;
        RECT -22.230 5.500 -21.880 5.670 ;
        RECT -18.930 5.500 -18.700 6.190 ;
        RECT -15.620 5.310 -15.070 5.740 ;
        RECT -14.290 5.310 -13.740 5.740 ;
        RECT -10.660 5.500 -10.430 6.190 ;
        RECT -5.360 5.960 -5.190 6.480 ;
        RECT -2.800 6.040 -2.620 6.970 ;
        RECT -2.070 6.710 -1.740 6.880 ;
        RECT -0.980 6.860 -0.550 7.120 ;
        RECT -0.750 6.830 -0.550 6.860 ;
        RECT 1.210 7.040 1.790 7.210 ;
        RECT 1.210 6.940 1.600 7.040 ;
        RECT 1.210 6.910 1.590 6.940 ;
        RECT 1.210 6.760 1.570 6.910 ;
        RECT -1.990 6.570 -1.740 6.710 ;
        RECT 0.860 6.590 1.570 6.760 ;
        RECT -1.990 6.310 -1.510 6.570 ;
        RECT -1.160 6.470 -0.990 6.510 ;
        RECT -0.750 6.470 -0.550 6.500 ;
        RECT -5.520 5.700 -5.190 5.960 ;
        RECT -2.920 6.010 -2.600 6.040 ;
        RECT -2.920 5.820 -2.590 6.010 ;
        RECT -2.920 5.780 -2.600 5.820 ;
        RECT -7.480 5.500 -7.130 5.670 ;
        RECT -6.110 5.500 -5.780 5.670 ;
        RECT -23.580 4.710 -23.250 4.880 ;
        RECT -22.230 4.710 -21.890 4.880 ;
        RECT -25.010 3.970 -24.830 4.160 ;
        RECT -23.500 4.140 -23.330 4.710 ;
        RECT -17.860 4.480 -17.670 4.880 ;
        RECT -11.690 4.480 -11.500 4.880 ;
        RECT -7.470 4.710 -7.130 4.880 ;
        RECT -6.110 4.710 -5.780 4.880 ;
        RECT -5.360 4.790 -5.190 5.700 ;
        RECT -17.860 4.470 -17.480 4.480 ;
        RECT -21.220 4.290 -17.480 4.470 ;
        RECT -17.860 4.250 -17.480 4.290 ;
        RECT -11.880 4.470 -11.500 4.480 ;
        RECT -11.880 4.290 -8.140 4.470 ;
        RECT -11.880 4.250 -11.500 4.290 ;
        RECT -25.430 3.160 -25.190 3.490 ;
        RECT -25.400 2.870 -25.200 3.160 ;
        RECT -25.390 2.860 -25.200 2.870 ;
        RECT -25.770 2.690 -25.560 2.700 ;
        RECT -25.770 2.110 -25.550 2.690 ;
        RECT -25.000 2.360 -24.830 3.970 ;
        RECT -24.170 3.200 -24.000 4.060 ;
        RECT -23.580 3.970 -23.250 4.140 ;
        RECT -22.230 3.970 -21.890 4.140 ;
        RECT -17.860 3.870 -17.670 4.250 ;
        RECT -15.620 3.580 -15.070 4.010 ;
        RECT -14.290 3.580 -13.740 4.010 ;
        RECT -11.690 3.870 -11.500 4.250 ;
        RECT -6.030 4.140 -5.860 4.710 ;
        RECT -7.470 3.970 -7.130 4.140 ;
        RECT -6.110 3.970 -5.780 4.140 ;
        RECT -24.170 2.940 -23.840 3.200 ;
        RECT -23.580 3.180 -23.250 3.350 ;
        RECT -22.230 3.180 -21.880 3.350 ;
        RECT -24.170 2.370 -24.000 2.940 ;
        RECT -18.930 2.560 -18.700 3.290 ;
        RECT -23.580 2.390 -23.250 2.560 ;
        RECT -22.230 2.390 -21.880 2.560 ;
        RECT -16.890 2.430 -16.550 2.680 ;
        RECT -10.660 2.560 -10.430 3.290 ;
        RECT -7.480 3.180 -7.130 3.350 ;
        RECT -6.110 3.180 -5.780 3.350 ;
        RECT -5.360 3.200 -5.190 4.060 ;
        RECT -5.520 2.940 -5.190 3.200 ;
        RECT -16.890 2.350 -16.540 2.430 ;
        RECT -7.480 2.390 -7.130 2.560 ;
        RECT -6.110 2.390 -5.780 2.560 ;
        RECT -5.360 2.370 -5.190 2.940 ;
        RECT -25.770 2.080 -25.560 2.110 ;
        RECT -25.760 1.730 -25.560 2.080 ;
        RECT -24.280 1.810 -23.750 1.980 ;
        RECT -21.590 1.500 -16.540 2.350 ;
        RECT -5.610 1.810 -5.080 1.980 ;
        RECT -2.800 1.870 -2.620 5.780 ;
        RECT -1.990 4.930 -1.820 6.310 ;
        RECT -1.160 6.210 -0.550 6.470 ;
        RECT -1.160 6.180 -0.990 6.210 ;
        RECT -0.750 6.170 -0.550 6.210 ;
        RECT -1.160 5.640 -0.990 5.670 ;
        RECT -0.750 5.640 -0.550 5.680 ;
        RECT -1.160 5.380 -0.550 5.640 ;
        RECT -1.160 5.340 -0.990 5.380 ;
        RECT -0.750 5.350 -0.550 5.380 ;
        RECT -1.710 3.830 -1.520 3.950 ;
        RECT -2.070 3.720 -1.520 3.830 ;
        RECT -2.070 3.660 -1.530 3.720 ;
        RECT -1.990 1.880 -1.820 3.660 ;
        RECT -1.160 3.510 -0.990 3.550 ;
        RECT -0.750 3.510 -0.550 3.540 ;
        RECT -1.160 3.250 -0.550 3.510 ;
        RECT -1.160 3.220 -0.990 3.250 ;
        RECT -0.750 3.210 -0.550 3.250 ;
        RECT -1.160 2.680 -0.990 2.710 ;
        RECT -0.750 2.680 -0.550 2.720 ;
        RECT -1.160 2.420 -0.550 2.680 ;
        RECT -1.160 2.380 -0.990 2.420 ;
        RECT -0.750 2.390 -0.550 2.420 ;
        RECT 0.860 2.100 1.570 2.270 ;
        RECT -0.750 2.030 -0.550 2.060 ;
        RECT -0.980 1.770 -0.550 2.030 ;
        RECT -0.750 1.730 -0.550 1.770 ;
        RECT 1.210 1.820 1.570 2.100 ;
        RECT 1.210 1.650 1.790 1.820 ;
      LAYER mcon ;
        RECT -23.930 6.870 -23.750 7.040 ;
        RECT -25.740 6.570 -25.570 6.740 ;
        RECT -25.390 5.730 -25.210 5.920 ;
        RECT -18.900 5.990 -18.730 6.160 ;
        RECT -24.070 5.740 -23.900 5.910 ;
        RECT -10.630 5.990 -10.460 6.160 ;
        RECT -18.900 5.540 -18.730 5.710 ;
        RECT -15.340 5.390 -15.070 5.660 ;
        RECT -14.290 5.390 -14.020 5.660 ;
        RECT -0.920 6.900 -0.750 7.070 ;
        RECT 1.330 6.950 1.500 7.120 ;
        RECT -1.740 6.350 -1.570 6.520 ;
        RECT -10.630 5.540 -10.460 5.710 ;
        RECT -5.460 5.740 -5.290 5.910 ;
        RECT -2.860 5.830 -2.690 6.000 ;
        RECT -17.660 4.280 -17.490 4.450 ;
        RECT -11.870 4.280 -11.700 4.450 ;
        RECT -25.390 2.930 -25.210 3.120 ;
        RECT -15.340 3.660 -15.070 3.930 ;
        RECT -14.290 3.660 -14.020 3.930 ;
        RECT -24.070 2.980 -23.900 3.150 ;
        RECT -18.900 3.040 -18.730 3.210 ;
        RECT -18.900 2.590 -18.730 2.760 ;
        RECT -10.630 3.040 -10.460 3.210 ;
        RECT -5.460 2.980 -5.290 3.150 ;
        RECT -16.780 2.460 -16.610 2.630 ;
        RECT -10.630 2.590 -10.460 2.760 ;
        RECT -25.740 2.110 -25.570 2.280 ;
        RECT -23.930 1.810 -23.750 1.980 ;
        RECT -0.970 6.250 -0.800 6.420 ;
        RECT -0.970 5.430 -0.800 5.600 ;
        RECT -1.700 3.750 -1.530 3.920 ;
        RECT -0.970 3.290 -0.800 3.460 ;
        RECT -0.970 2.470 -0.800 2.640 ;
        RECT -0.920 1.820 -0.750 1.990 ;
        RECT 1.290 1.760 1.460 1.930 ;
      LAYER met1 ;
        RECT -25.920 6.800 -25.640 7.450 ;
        RECT -25.920 6.200 -25.530 6.800 ;
        RECT -25.920 2.650 -25.640 6.200 ;
        RECT -25.390 5.990 -25.200 7.450 ;
        RECT -23.980 6.770 -23.680 7.150 ;
        RECT -18.910 6.240 -18.680 7.450 ;
        RECT -17.690 6.480 -17.460 7.450 ;
        RECT -25.420 5.960 -25.200 5.990 ;
        RECT -25.430 5.690 -25.180 5.960 ;
        RECT -25.430 5.680 -25.190 5.690 ;
        RECT -25.420 5.440 -25.190 5.680 ;
        RECT -24.150 5.670 -23.830 5.990 ;
        RECT -18.940 5.450 -18.680 6.240 ;
        RECT -17.700 6.230 -17.460 6.480 ;
        RECT -25.390 3.410 -25.230 5.440 ;
        RECT -25.040 4.880 -24.800 5.010 ;
        RECT -25.060 4.560 -24.800 4.880 ;
        RECT -25.060 3.960 -24.800 4.280 ;
        RECT -25.040 3.840 -24.800 3.960 ;
        RECT -25.420 3.170 -25.190 3.410 ;
        RECT -18.910 3.300 -18.680 5.450 ;
        RECT -25.430 3.160 -25.190 3.170 ;
        RECT -25.430 2.890 -25.180 3.160 ;
        RECT -24.150 2.910 -23.830 3.230 ;
        RECT -25.420 2.860 -25.200 2.890 ;
        RECT -25.920 2.050 -25.530 2.650 ;
        RECT -25.920 1.400 -25.640 2.050 ;
        RECT -25.390 1.400 -25.200 2.860 ;
        RECT -18.940 2.510 -18.680 3.300 ;
        RECT -23.980 1.700 -23.680 2.080 ;
        RECT -18.910 1.400 -18.680 2.510 ;
        RECT -17.690 1.400 -17.460 6.230 ;
        RECT -16.860 2.390 -16.540 2.710 ;
        RECT -15.400 1.410 -14.980 7.450 ;
        RECT -14.380 1.400 -13.960 7.450 ;
        RECT -11.900 1.400 -11.670 7.450 ;
        RECT -10.680 6.240 -10.450 7.450 ;
        RECT -5.680 6.770 -5.380 7.150 ;
        RECT -0.990 6.830 -0.670 7.150 ;
        RECT 1.260 6.880 1.580 7.200 ;
        RECT -1.820 6.280 -1.500 6.600 ;
        RECT -10.680 5.450 -10.420 6.240 ;
        RECT -1.040 6.180 -0.720 6.500 ;
        RECT -5.530 5.670 -5.210 5.990 ;
        RECT -2.930 5.750 -2.610 6.070 ;
        RECT -1.710 5.590 -1.500 5.700 ;
        RECT -10.680 3.300 -10.450 5.450 ;
        RECT -1.730 5.270 -1.470 5.590 ;
        RECT -1.040 5.350 -0.720 5.670 ;
        RECT -1.710 3.980 -1.500 5.270 ;
        RECT -1.730 3.690 -1.500 3.980 ;
        RECT -10.680 2.510 -10.420 3.300 ;
        RECT -5.530 2.910 -5.210 3.230 ;
        RECT -1.040 3.220 -0.720 3.540 ;
        RECT -10.680 1.400 -10.450 2.510 ;
        RECT -1.040 2.390 -0.720 2.710 ;
        RECT -5.680 1.700 -5.380 2.080 ;
        RECT -0.990 1.740 -0.670 2.060 ;
        RECT 1.220 1.690 1.540 2.010 ;
      LAYER via ;
        RECT -23.960 6.830 -23.700 7.100 ;
        RECT -24.120 5.700 -23.860 5.960 ;
        RECT -25.060 4.590 -24.800 4.850 ;
        RECT -25.060 3.990 -24.800 4.250 ;
        RECT -24.120 2.940 -23.860 3.200 ;
        RECT -23.960 1.750 -23.700 2.020 ;
        RECT -16.830 2.420 -16.570 2.680 ;
        RECT -5.660 6.830 -5.400 7.100 ;
        RECT -0.960 6.860 -0.700 7.120 ;
        RECT 1.290 6.910 1.550 7.170 ;
        RECT -1.790 6.310 -1.530 6.570 ;
        RECT -1.010 6.210 -0.750 6.470 ;
        RECT -5.500 5.700 -5.240 5.960 ;
        RECT -2.900 5.780 -2.640 6.040 ;
        RECT -1.730 5.300 -1.470 5.560 ;
        RECT -1.010 5.380 -0.750 5.640 ;
        RECT -1.010 3.250 -0.750 3.510 ;
        RECT -5.500 2.940 -5.240 3.200 ;
        RECT -1.010 2.420 -0.750 2.680 ;
        RECT -5.660 1.750 -5.400 2.020 ;
        RECT -0.960 1.770 -0.700 2.030 ;
        RECT 1.250 1.720 1.510 1.980 ;
      LAYER met2 ;
        RECT -23.980 6.970 -23.680 7.150 ;
        RECT -5.680 6.970 -5.380 7.150 ;
        RECT -23.980 6.950 -23.430 6.970 ;
        RECT -5.930 6.950 -5.380 6.970 ;
        RECT -0.990 7.110 -0.680 7.160 ;
        RECT 1.260 7.110 1.570 7.210 ;
        RECT -26.160 6.770 -3.200 6.950 ;
        RECT -0.990 6.880 1.570 7.110 ;
        RECT -0.990 6.830 -0.680 6.880 ;
        RECT -1.810 6.570 -1.500 6.610 ;
        RECT -1.990 6.430 -1.270 6.570 ;
        RECT -1.040 6.430 -0.730 6.510 ;
        RECT -1.990 6.320 -0.730 6.430 ;
        RECT -1.810 6.280 -0.730 6.320 ;
        RECT -1.540 6.220 -0.730 6.280 ;
        RECT -1.540 6.210 -1.270 6.220 ;
        RECT -1.040 6.180 -0.730 6.220 ;
        RECT -24.140 5.930 -23.830 6.000 ;
        RECT -26.160 5.920 -23.830 5.930 ;
        RECT -5.530 5.930 -5.220 6.000 ;
        RECT -2.930 5.930 -2.620 6.070 ;
        RECT -26.160 5.710 -6.670 5.920 ;
        RECT -24.850 5.700 -6.670 5.710 ;
        RECT -24.140 5.670 -23.830 5.700 ;
        RECT -25.090 4.730 -7.850 4.950 ;
        RECT -25.090 4.590 -24.770 4.730 ;
        RECT -25.070 4.250 -24.810 4.590 ;
        RECT -25.090 3.990 -24.770 4.250 ;
        RECT -24.140 3.170 -23.830 3.240 ;
        RECT -26.160 2.960 -11.150 3.170 ;
        RECT -24.850 2.950 -11.150 2.960 ;
        RECT -24.140 2.910 -23.830 2.950 ;
        RECT -16.850 2.650 -16.540 2.720 ;
        RECT -17.310 2.640 -16.420 2.650 ;
        RECT -17.310 2.430 -14.630 2.640 ;
        RECT -11.370 2.620 -11.150 2.950 ;
        RECT -8.070 3.120 -7.850 4.730 ;
        RECT -6.890 4.500 -6.670 5.700 ;
        RECT -5.530 5.740 -2.620 5.930 ;
        RECT -5.530 5.710 -2.930 5.740 ;
        RECT -5.530 5.670 -5.220 5.710 ;
        RECT -1.470 5.640 -1.270 5.650 ;
        RECT -1.470 5.630 -1.250 5.640 ;
        RECT -1.040 5.630 -0.730 5.670 ;
        RECT -1.470 5.560 -0.730 5.630 ;
        RECT -1.760 5.540 -0.730 5.560 ;
        RECT -1.810 5.420 -0.730 5.540 ;
        RECT -1.810 5.300 -1.250 5.420 ;
        RECT -1.040 5.340 -0.730 5.420 ;
        RECT -1.810 5.290 -1.340 5.300 ;
        RECT -6.920 4.460 -6.670 4.500 ;
        RECT -6.920 3.820 -6.660 4.460 ;
        RECT -6.920 3.610 -2.790 3.820 ;
        RECT -3.000 3.470 -2.790 3.610 ;
        RECT -1.040 3.470 -0.730 3.550 ;
        RECT -3.000 3.260 -0.730 3.470 ;
        RECT -5.530 3.170 -5.220 3.240 ;
        RECT -1.040 3.220 -0.730 3.260 ;
        RECT -5.530 3.120 -3.200 3.170 ;
        RECT -8.070 2.960 -3.200 3.120 ;
        RECT -8.070 2.900 -5.220 2.960 ;
        RECT -1.040 2.670 -0.730 2.710 ;
        RECT -7.000 2.620 -0.730 2.670 ;
        RECT -11.370 2.460 -0.730 2.620 ;
        RECT -17.310 2.410 -16.420 2.430 ;
        RECT -16.850 2.390 -16.540 2.410 ;
        RECT -11.370 2.400 -6.610 2.460 ;
        RECT -1.040 2.380 -0.730 2.460 ;
        RECT -23.850 2.080 -23.690 2.090 ;
        RECT -5.670 2.080 -5.510 2.090 ;
        RECT -26.160 2.070 -23.600 2.080 ;
        RECT -5.760 2.070 -3.200 2.080 ;
        RECT -26.160 1.920 -3.200 2.070 ;
        RECT -26.160 1.900 -23.600 1.920 ;
        RECT -5.760 1.900 -3.200 1.920 ;
        RECT -0.990 1.980 -0.680 2.060 ;
        RECT 1.220 1.980 1.530 2.020 ;
        RECT -23.980 1.700 -23.680 1.900 ;
        RECT -5.680 1.700 -5.380 1.900 ;
        RECT -0.990 1.750 1.720 1.980 ;
        RECT -0.990 1.730 -0.680 1.750 ;
        RECT 1.220 1.690 1.530 1.750 ;
  END
END sky130_hilas_TA2Cell_1FG

MACRO sky130_hilas_swc2x2varactor
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc2x2varactor ;
  ORIGIN 14.660 4.420 ;
  SIZE 14.680 BY 7.010 ;
  OBS
      LAYER nwell ;
        RECT -14.660 1.750 -12.750 2.270 ;
        RECT -14.650 -4.400 -12.750 1.750 ;
        RECT -9.920 0.260 -7.130 2.240 ;
        RECT -9.940 -2.530 -7.120 0.260 ;
        RECT -9.900 -4.400 -7.120 -2.530 ;
        RECT -5.720 -4.400 -4.250 2.260 ;
        RECT -3.240 0.170 0.020 2.380 ;
        RECT -3.240 0.160 -0.020 0.170 ;
        RECT -5.070 -4.420 -4.250 -4.400 ;
      LAYER li1 ;
        RECT -5.230 1.720 -4.890 1.890 ;
        RECT -2.560 1.500 -2.210 1.670 ;
        RECT -1.660 1.410 -1.460 1.750 ;
        RECT -5.230 0.930 -4.890 1.100 ;
        RECT -2.560 0.880 -2.210 1.050 ;
        RECT -0.930 0.800 -0.730 1.800 ;
        RECT -5.230 0.360 -4.890 0.530 ;
        RECT -5.240 -1.170 -4.890 -1.000 ;
        RECT -5.230 -2.690 -4.890 -2.520 ;
        RECT -5.230 -3.250 -4.890 -3.080 ;
        RECT -13.790 -3.950 -13.510 -3.520 ;
        RECT -6.600 -3.780 -6.260 -3.610 ;
        RECT -5.230 -4.040 -4.890 -3.870 ;
  END
END sky130_hilas_swc2x2varactor

MACRO sky130_hilas_drainSelect01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_drainSelect01 ;
  ORIGIN -10.720 -0.050 ;
  SIZE 5.420 BY 6.050 ;
  PIN DRAIN4
    ANTENNADIFFAREA 0.275800 ;
    PORT
      LAYER li1 ;
        RECT 12.100 0.620 12.270 0.630 ;
        RECT 14.810 0.620 15.050 0.660 ;
        RECT 11.820 0.450 12.780 0.620 ;
        RECT 14.810 0.450 15.380 0.620 ;
        RECT 14.810 0.420 15.050 0.450 ;
      LAYER mcon ;
        RECT 12.100 0.460 12.270 0.630 ;
        RECT 14.850 0.450 15.020 0.620 ;
      LAYER met1 ;
        RECT 12.230 0.660 12.570 0.700 ;
        RECT 12.010 0.620 12.570 0.660 ;
        RECT 14.660 0.670 15.030 0.680 ;
        RECT 12.010 0.450 12.690 0.620 ;
        RECT 12.010 0.430 12.570 0.450 ;
        RECT 12.230 0.380 12.570 0.430 ;
        RECT 14.660 0.410 15.080 0.670 ;
        RECT 14.660 0.390 15.030 0.410 ;
      LAYER via ;
        RECT 12.280 0.410 12.540 0.670 ;
        RECT 14.690 0.410 14.950 0.670 ;
      LAYER met2 ;
        RECT 11.070 0.670 12.530 0.740 ;
        RECT 11.070 0.620 12.570 0.670 ;
        RECT 14.660 0.620 14.980 0.700 ;
        RECT 11.070 0.570 14.980 0.620 ;
        RECT 12.250 0.430 14.980 0.570 ;
        RECT 12.250 0.410 12.570 0.430 ;
        RECT 14.660 0.380 14.980 0.430 ;
    END
  END DRAIN4
  PIN DRAIN3
    ANTENNADIFFAREA 0.275800 ;
    PORT
      LAYER li1 ;
        RECT 14.810 2.770 15.050 2.800 ;
        RECT 11.820 2.600 12.780 2.770 ;
        RECT 14.810 2.600 15.380 2.770 ;
        RECT 12.100 2.590 12.270 2.600 ;
        RECT 14.810 2.560 15.050 2.600 ;
      LAYER mcon ;
        RECT 14.850 2.600 15.020 2.770 ;
      LAYER met1 ;
        RECT 12.230 2.790 12.570 2.840 ;
        RECT 12.010 2.770 12.570 2.790 ;
        RECT 14.660 2.810 15.030 2.830 ;
        RECT 12.010 2.600 12.690 2.770 ;
        RECT 12.010 2.560 12.570 2.600 ;
        RECT 12.230 2.520 12.570 2.560 ;
        RECT 14.660 2.550 15.080 2.810 ;
        RECT 14.660 2.540 15.030 2.550 ;
      LAYER via ;
        RECT 12.280 2.550 12.540 2.810 ;
        RECT 14.690 2.550 14.950 2.810 ;
      LAYER met2 ;
        RECT 12.250 2.790 12.570 2.810 ;
        RECT 14.660 2.790 14.980 2.840 ;
        RECT 12.250 2.600 14.980 2.790 ;
        RECT 11.070 2.570 11.770 2.580 ;
        RECT 12.250 2.570 12.570 2.600 ;
        RECT 11.070 2.550 12.570 2.570 ;
        RECT 11.070 2.410 12.500 2.550 ;
        RECT 14.660 2.520 14.980 2.600 ;
    END
  END DRAIN3
  PIN DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.275800 ;
    PORT
      LAYER li1 ;
        RECT 12.100 3.550 12.270 3.560 ;
        RECT 14.810 3.550 15.050 3.590 ;
        RECT 11.820 3.380 12.780 3.550 ;
        RECT 14.810 3.380 15.380 3.550 ;
        RECT 14.810 3.350 15.050 3.380 ;
      LAYER mcon ;
        RECT 12.100 3.390 12.270 3.560 ;
        RECT 14.850 3.380 15.020 3.550 ;
      LAYER met1 ;
        RECT 12.230 3.590 12.570 3.630 ;
        RECT 12.010 3.550 12.570 3.590 ;
        RECT 14.660 3.600 15.030 3.610 ;
        RECT 12.010 3.380 12.690 3.550 ;
        RECT 12.010 3.360 12.570 3.380 ;
        RECT 12.230 3.310 12.570 3.360 ;
        RECT 14.660 3.340 15.080 3.600 ;
        RECT 14.660 3.320 15.030 3.340 ;
      LAYER via ;
        RECT 12.280 3.340 12.540 3.600 ;
        RECT 14.690 3.340 14.950 3.600 ;
      LAYER met2 ;
        RECT 11.070 3.720 11.740 3.740 ;
        RECT 11.070 3.600 12.460 3.720 ;
        RECT 11.070 3.560 12.570 3.600 ;
        RECT 12.250 3.550 12.570 3.560 ;
        RECT 14.660 3.550 14.980 3.630 ;
        RECT 12.250 3.360 14.980 3.550 ;
        RECT 12.250 3.340 12.570 3.360 ;
        RECT 14.660 3.310 14.980 3.360 ;
    END
  END DRAIN2
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.275800 ;
    PORT
      LAYER li1 ;
        RECT 14.810 5.700 15.050 5.730 ;
        RECT 11.820 5.530 12.780 5.700 ;
        RECT 14.810 5.530 15.380 5.700 ;
        RECT 12.100 5.520 12.270 5.530 ;
        RECT 14.810 5.490 15.050 5.530 ;
      LAYER mcon ;
        RECT 14.850 5.530 15.020 5.700 ;
      LAYER met1 ;
        RECT 12.230 5.720 12.570 5.770 ;
        RECT 12.010 5.700 12.570 5.720 ;
        RECT 14.660 5.740 15.030 5.760 ;
        RECT 12.010 5.530 12.690 5.700 ;
        RECT 12.010 5.490 12.570 5.530 ;
        RECT 12.230 5.450 12.570 5.490 ;
        RECT 14.660 5.480 15.080 5.740 ;
        RECT 14.660 5.470 15.030 5.480 ;
      LAYER via ;
        RECT 12.280 5.480 12.540 5.740 ;
        RECT 14.690 5.480 14.950 5.740 ;
      LAYER met2 ;
        RECT 12.250 5.720 12.570 5.740 ;
        RECT 14.660 5.720 14.980 5.770 ;
        RECT 11.070 5.590 11.800 5.600 ;
        RECT 12.250 5.590 14.980 5.720 ;
        RECT 11.070 5.530 14.980 5.590 ;
        RECT 11.070 5.480 12.570 5.530 ;
        RECT 11.070 5.430 12.490 5.480 ;
        RECT 14.660 5.450 14.980 5.530 ;
        RECT 11.070 5.420 11.800 5.430 ;
    END
  END DRAIN1
  PIN DRAINSELECT1
    USE ANALOG ;
    ANTENNAGATEAREA 0.625000 ;
    PORT
      LAYER li1 ;
        RECT 15.760 5.180 15.930 5.220 ;
        RECT 15.760 5.010 15.990 5.180 ;
        RECT 15.760 4.660 15.930 5.010 ;
      LAYER mcon ;
        RECT 15.820 5.010 15.990 5.180 ;
      LAYER met1 ;
        RECT 15.760 4.980 16.140 5.220 ;
    END
  END DRAINSELECT1
  PIN DRAINSELECT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.625000 ;
    PORT
      LAYER li1 ;
        RECT 15.760 4.070 15.930 4.420 ;
        RECT 15.760 3.900 15.990 4.070 ;
        RECT 15.760 3.860 15.930 3.900 ;
      LAYER mcon ;
        RECT 15.820 3.900 15.990 4.070 ;
      LAYER met1 ;
        RECT 15.760 3.860 16.140 4.100 ;
    END
  END DRAINSELECT2
  PIN DRAINSELECT3
    USE ANALOG ;
    ANTENNAGATEAREA 0.625000 ;
    PORT
      LAYER li1 ;
        RECT 15.760 2.250 15.930 2.290 ;
        RECT 15.760 2.080 15.990 2.250 ;
        RECT 15.760 1.730 15.930 2.080 ;
      LAYER mcon ;
        RECT 15.820 2.080 15.990 2.250 ;
      LAYER met1 ;
        RECT 15.760 2.050 16.140 2.290 ;
    END
  END DRAINSELECT3
  PIN DRAINSELECT4
    USE ANALOG ;
    ANTENNAGATEAREA 0.625000 ;
    PORT
      LAYER li1 ;
        RECT 15.760 1.140 15.930 1.490 ;
        RECT 15.760 0.970 15.990 1.140 ;
        RECT 15.760 0.930 15.930 0.970 ;
      LAYER mcon ;
        RECT 15.820 0.970 15.990 1.140 ;
      LAYER met1 ;
        RECT 15.760 0.930 16.140 1.170 ;
    END
  END DRAINSELECT4
  PIN VINJ
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 11.120 4.840 11.290 5.770 ;
        RECT 11.120 3.310 11.290 4.240 ;
        RECT 11.120 1.910 11.290 2.840 ;
        RECT 11.120 0.380 11.290 1.310 ;
      LAYER mcon ;
        RECT 11.120 5.200 11.290 5.370 ;
        RECT 11.120 3.710 11.290 3.880 ;
        RECT 11.120 2.270 11.290 2.440 ;
        RECT 11.120 0.780 11.290 0.950 ;
      LAYER met1 ;
        RECT 11.080 0.050 11.330 6.100 ;
    END
  END VINJ
  PIN DRAIN_MUX
    USE ANALOG ;
    ANTENNADIFFAREA 0.719200 ;
    PORT
      LAYER li1 ;
        RECT 13.230 5.530 14.570 5.700 ;
        RECT 13.230 3.380 14.570 3.550 ;
        RECT 13.230 2.600 14.570 2.770 ;
        RECT 13.230 0.450 14.570 0.620 ;
      LAYER mcon ;
        RECT 14.100 5.530 14.270 5.700 ;
        RECT 14.100 3.380 14.270 3.550 ;
        RECT 14.100 2.600 14.270 2.770 ;
        RECT 14.100 0.450 14.270 0.620 ;
      LAYER met1 ;
        RECT 14.070 0.050 14.300 6.100 ;
    END
  END DRAIN_MUX
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 15.400 5.080 15.590 5.100 ;
        RECT 15.030 4.910 15.590 5.080 ;
        RECT 15.400 4.870 15.590 4.910 ;
        RECT 15.400 4.170 15.590 4.210 ;
        RECT 15.030 4.000 15.590 4.170 ;
        RECT 15.400 3.980 15.590 4.000 ;
        RECT 15.400 2.150 15.590 2.170 ;
        RECT 15.030 1.980 15.590 2.150 ;
        RECT 15.400 1.940 15.590 1.980 ;
        RECT 15.400 1.240 15.590 1.280 ;
        RECT 15.030 1.070 15.590 1.240 ;
        RECT 15.400 1.050 15.590 1.070 ;
      LAYER mcon ;
        RECT 15.410 4.900 15.580 5.070 ;
        RECT 15.410 4.010 15.580 4.180 ;
        RECT 15.410 1.970 15.580 2.140 ;
        RECT 15.410 1.080 15.580 1.250 ;
      LAYER met1 ;
        RECT 15.420 5.130 15.610 6.100 ;
        RECT 15.380 4.840 15.610 5.130 ;
        RECT 15.420 4.240 15.610 4.840 ;
        RECT 15.380 3.950 15.610 4.240 ;
        RECT 15.420 2.200 15.610 3.950 ;
        RECT 15.380 1.910 15.610 2.200 ;
        RECT 15.420 1.310 15.610 1.910 ;
        RECT 15.380 1.020 15.610 1.310 ;
        RECT 15.420 0.050 15.610 1.020 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 10.720 0.050 13.920 6.100 ;
      LAYER li1 ;
        RECT 12.260 5.080 12.590 5.260 ;
        RECT 11.820 4.910 14.570 5.080 ;
        RECT 11.820 4.000 14.570 4.170 ;
        RECT 12.260 3.820 12.590 4.000 ;
        RECT 12.260 2.150 12.590 2.330 ;
        RECT 11.820 1.980 14.570 2.150 ;
        RECT 11.820 1.070 14.570 1.240 ;
        RECT 12.260 0.890 12.590 1.070 ;
  END
END sky130_hilas_drainSelect01

MACRO sky130_hilas_TunVaractorCapcitor
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TunVaractorCapcitor ;
  ORIGIN 14.660 4.420 ;
  SIZE 10.430 BY 7.010 ;
  OBS
      LAYER nwell ;
        RECT -14.660 1.750 -12.750 2.260 ;
        RECT -14.650 -4.400 -12.750 1.750 ;
        RECT -9.920 0.260 -7.130 2.240 ;
        RECT -9.940 -2.530 -7.120 0.260 ;
        RECT -9.900 -4.400 -7.120 -2.530 ;
        RECT -5.720 -4.400 -4.250 2.260 ;
        RECT -5.070 -4.420 -4.250 -4.400 ;
      LAYER li1 ;
        RECT -5.230 1.720 -4.890 1.890 ;
        RECT -5.230 0.930 -4.890 1.100 ;
        RECT -5.230 0.360 -4.890 0.530 ;
        RECT -5.240 -1.170 -4.890 -1.000 ;
        RECT -5.230 -2.690 -4.890 -2.520 ;
        RECT -5.230 -3.250 -4.890 -3.080 ;
        RECT -13.790 -3.950 -13.510 -3.520 ;
        RECT -6.600 -3.780 -6.260 -3.610 ;
        RECT -5.230 -4.040 -4.890 -3.870 ;
  END
END sky130_hilas_TunVaractorCapcitor

MACRO sky130_hilas_pFETmirror
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pFETmirror ;
  ORIGIN 0.610 -0.820 ;
  SIZE 2.190 BY 2.030 ;
  OBS
      LAYER nwell ;
        RECT -0.610 1.120 1.580 2.850 ;
      LAYER li1 ;
        RECT -0.400 2.010 1.360 2.530 ;
        RECT -0.400 1.400 0.310 1.570 ;
        RECT 0.620 1.400 1.320 1.570 ;
        RECT -0.050 1.230 0.310 1.400 ;
        RECT -0.050 0.870 0.600 1.230 ;
        RECT -0.050 0.820 0.220 0.870 ;
        RECT 0.850 0.820 1.100 1.400 ;
  END
END sky130_hilas_pFETmirror

MACRO sky130_hilas_pFETdevice01c
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pFETdevice01c ;
  ORIGIN 0.790 1.140 ;
  SIZE 1.870 BY 1.570 ;
  OBS
      LAYER nwell ;
        RECT -0.790 -0.780 0.820 0.430 ;
      LAYER li1 ;
        RECT 0.780 -1.060 0.990 -0.630 ;
        RECT 0.800 -1.080 0.970 -1.060 ;
      LAYER met1 ;
        RECT 0.780 -0.850 1.000 -0.630 ;
        RECT 0.770 -1.140 1.000 -0.850 ;
  END
END sky130_hilas_pFETdevice01c

MACRO sky130_hilas_swc4x1BiasCell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc4x1BiasCell ;
  ORIGIN 2.660 3.820 ;
  SIZE 10.110 BY 6.050 ;
  PIN BIAS1
    USE ANALOG ;
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER li1 ;
        RECT 4.980 1.240 5.300 1.280 ;
        RECT 4.980 1.200 5.310 1.240 ;
        RECT 4.980 1.030 5.560 1.200 ;
        RECT 4.980 1.020 5.300 1.030 ;
      LAYER mcon ;
        RECT 5.040 1.060 5.210 1.230 ;
      LAYER met1 ;
        RECT 4.970 0.990 5.290 1.310 ;
      LAYER via ;
        RECT 5.000 1.020 5.260 1.280 ;
      LAYER met2 ;
        RECT 4.970 1.300 5.280 1.320 ;
        RECT -2.640 1.120 7.440 1.300 ;
        RECT -2.640 1.110 -2.490 1.120 ;
        RECT 4.970 0.990 5.280 1.120 ;
    END
  END BIAS1
  PIN BIAS2
    USE ANALOG ;
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER li1 ;
        RECT 4.980 0.390 5.300 0.400 ;
        RECT 4.980 0.220 5.560 0.390 ;
        RECT 4.980 0.180 5.310 0.220 ;
        RECT 4.980 0.140 5.300 0.180 ;
      LAYER mcon ;
        RECT 5.040 0.190 5.210 0.360 ;
      LAYER met1 ;
        RECT 4.970 0.110 5.290 0.430 ;
      LAYER via ;
        RECT 5.000 0.140 5.260 0.400 ;
      LAYER met2 ;
        RECT -2.660 0.300 -2.520 0.320 ;
        RECT 4.970 0.300 5.280 0.430 ;
        RECT -2.660 0.120 7.450 0.300 ;
        RECT 4.970 0.100 5.280 0.120 ;
    END
  END BIAS2
  PIN BIAS3
    USE ANALOG ;
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER li1 ;
        RECT 4.980 -1.770 5.300 -1.730 ;
        RECT 4.980 -1.810 5.310 -1.770 ;
        RECT 4.980 -1.980 5.560 -1.810 ;
        RECT 4.980 -1.990 5.300 -1.980 ;
      LAYER mcon ;
        RECT 5.040 -1.950 5.210 -1.780 ;
      LAYER met1 ;
        RECT 4.970 -2.020 5.290 -1.700 ;
      LAYER via ;
        RECT 5.000 -1.990 5.260 -1.730 ;
      LAYER met2 ;
        RECT 4.970 -1.710 5.280 -1.690 ;
        RECT -2.630 -1.870 7.440 -1.710 ;
        RECT -2.620 -1.880 7.440 -1.870 ;
        RECT 4.880 -1.890 7.440 -1.880 ;
        RECT 4.970 -2.020 5.280 -1.890 ;
    END
  END BIAS3
  PIN BIAS4
    USE ANALOG ;
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER li1 ;
        RECT 4.980 -2.610 5.300 -2.600 ;
        RECT 4.980 -2.780 5.560 -2.610 ;
        RECT 4.980 -2.820 5.310 -2.780 ;
        RECT 4.980 -2.860 5.300 -2.820 ;
      LAYER mcon ;
        RECT 5.040 -2.810 5.210 -2.640 ;
      LAYER met1 ;
        RECT 4.970 -2.890 5.290 -2.570 ;
      LAYER via ;
        RECT 5.000 -2.860 5.260 -2.600 ;
      LAYER met2 ;
        RECT 4.970 -2.690 5.280 -2.570 ;
        RECT -2.630 -2.700 5.280 -2.690 ;
        RECT -2.630 -2.860 7.440 -2.700 ;
        RECT -1.840 -2.950 -0.300 -2.860 ;
        RECT 4.880 -2.880 7.440 -2.860 ;
        RECT 4.970 -2.900 5.280 -2.880 ;
    END
  END BIAS4
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 1.978000 ;
    PORT
      LAYER nwell ;
        RECT -2.630 1.600 -0.900 2.230 ;
        RECT -2.640 -1.470 -0.900 1.600 ;
        RECT -2.630 -3.820 -0.900 -1.470 ;
      LAYER li1 ;
        RECT -2.210 -1.020 -1.660 -0.590 ;
      LAYER mcon ;
        RECT -2.210 -0.940 -1.940 -0.670 ;
      LAYER met1 ;
        RECT -2.280 -3.820 -1.880 2.230 ;
    END
  END VTUN
  PIN GATE
    USE ANALOG ;
    ANTENNADIFFAREA 2.743300 ;
    PORT
      LAYER nwell ;
        RECT 1.120 -3.820 3.350 2.230 ;
      LAYER li1 ;
        RECT 1.820 -1.090 2.370 -0.660 ;
      LAYER mcon ;
        RECT 1.820 -1.010 2.090 -0.740 ;
      LAYER met1 ;
        RECT 1.770 0.310 2.150 2.230 ;
        RECT 1.760 -1.550 2.150 0.310 ;
        RECT 1.770 -3.820 2.150 -1.550 ;
    END
  END GATE
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 4.880 2.220 7.430 2.230 ;
        RECT 4.880 -3.800 7.440 2.220 ;
        RECT 4.880 -3.810 7.430 -3.800 ;
      LAYER li1 ;
        RECT 6.840 1.550 7.040 1.900 ;
        RECT 6.840 1.520 7.050 1.550 ;
        RECT 6.830 0.930 7.050 1.520 ;
        RECT 6.830 -0.100 7.050 0.490 ;
        RECT 6.840 -0.130 7.050 -0.100 ;
        RECT 6.840 -0.480 7.040 -0.130 ;
        RECT 6.840 -1.460 7.040 -1.110 ;
        RECT 6.840 -1.490 7.050 -1.460 ;
        RECT 6.830 -2.080 7.050 -1.490 ;
        RECT 6.830 -3.100 7.050 -2.510 ;
        RECT 6.840 -3.130 7.050 -3.100 ;
        RECT 6.840 -3.480 7.040 -3.130 ;
      LAYER mcon ;
        RECT 6.850 1.350 7.020 1.520 ;
        RECT 6.850 -0.100 7.020 0.070 ;
        RECT 6.850 -1.660 7.020 -1.490 ;
        RECT 6.850 -3.100 7.020 -2.930 ;
      LAYER met1 ;
        RECT 6.920 1.580 7.080 2.230 ;
        RECT 6.810 1.030 7.080 1.580 ;
        RECT 6.810 0.980 7.090 1.030 ;
        RECT 6.920 0.890 7.090 0.980 ;
        RECT 6.920 0.530 7.080 0.890 ;
        RECT 6.920 0.440 7.090 0.530 ;
        RECT 6.810 0.390 7.090 0.440 ;
        RECT 6.810 -0.160 7.080 0.390 ;
        RECT 6.920 -1.430 7.080 -0.160 ;
        RECT 6.810 -1.980 7.080 -1.430 ;
        RECT 6.810 -2.030 7.090 -1.980 ;
        RECT 6.920 -2.120 7.090 -2.030 ;
        RECT 6.920 -2.470 7.080 -2.120 ;
        RECT 6.920 -2.560 7.090 -2.470 ;
        RECT 6.810 -2.610 7.090 -2.560 ;
        RECT 6.810 -3.160 7.080 -2.610 ;
        RECT 6.920 -3.810 7.080 -3.160 ;
    END
  END VINJ
  PIN VPWR
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 6.110 0.960 6.310 1.530 ;
        RECT 6.110 -0.110 6.310 0.460 ;
        RECT 6.110 -2.050 6.310 -1.480 ;
        RECT 6.110 -3.110 6.310 -2.540 ;
      LAYER mcon ;
        RECT 6.120 1.320 6.290 1.490 ;
        RECT 6.120 -0.070 6.290 0.100 ;
        RECT 6.120 -1.690 6.290 -1.520 ;
        RECT 6.120 -3.070 6.290 -2.900 ;
      LAYER met1 ;
        RECT 6.110 1.550 6.270 2.230 ;
        RECT 6.110 1.530 6.310 1.550 ;
        RECT 6.090 1.290 6.320 1.530 ;
        RECT 6.110 1.070 6.310 1.290 ;
        RECT 6.110 0.350 6.270 1.070 ;
        RECT 6.110 0.130 6.310 0.350 ;
        RECT 6.090 -0.110 6.320 0.130 ;
        RECT 6.110 -0.130 6.310 -0.110 ;
        RECT 6.110 -1.460 6.270 -0.130 ;
        RECT 6.110 -1.480 6.310 -1.460 ;
        RECT 6.090 -1.720 6.320 -1.480 ;
        RECT 6.110 -1.940 6.310 -1.720 ;
        RECT 6.110 -2.650 6.270 -1.940 ;
        RECT 6.110 -2.870 6.310 -2.650 ;
        RECT 6.090 -3.110 6.320 -2.870 ;
        RECT 6.110 -3.130 6.310 -3.110 ;
        RECT 6.110 -3.810 6.270 -3.130 ;
    END
  END VPWR
  PIN GATESELECT
    USE ANALOG ;
    ANTENNAGATEAREA 0.620000 ;
    PORT
      LAYER li1 ;
        RECT 6.230 -0.880 6.670 -0.710 ;
      LAYER mcon ;
        RECT 6.490 -0.880 6.670 -0.710 ;
      LAYER met1 ;
        RECT 6.480 1.240 6.670 2.230 ;
        RECT 6.500 1.120 6.670 1.240 ;
        RECT 6.510 0.300 6.670 1.120 ;
        RECT 6.500 0.180 6.670 0.300 ;
        RECT 6.480 -0.680 6.670 0.180 ;
        RECT 6.460 -0.910 6.700 -0.680 ;
        RECT 6.480 -1.770 6.670 -0.910 ;
        RECT 6.500 -1.890 6.670 -1.770 ;
        RECT 6.510 -2.700 6.670 -1.890 ;
        RECT 6.500 -2.820 6.670 -2.700 ;
        RECT 6.480 -3.810 6.670 -2.820 ;
    END
  END GATESELECT
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER li1 ;
        RECT 4.980 1.820 5.300 1.830 ;
        RECT 4.980 1.650 5.560 1.820 ;
        RECT 4.980 1.600 5.310 1.650 ;
        RECT 4.980 1.570 5.300 1.600 ;
      LAYER mcon ;
        RECT 5.040 1.610 5.210 1.780 ;
      LAYER met1 ;
        RECT 4.970 1.540 5.290 1.860 ;
      LAYER via ;
        RECT 5.000 1.570 5.260 1.830 ;
      LAYER met2 ;
        RECT 4.970 1.730 5.280 1.870 ;
        RECT 4.870 1.550 7.440 1.730 ;
        RECT 4.970 1.540 5.280 1.550 ;
    END
  END DRAIN1
  PIN DRAIN2
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER li1 ;
        RECT 4.980 -0.180 5.300 -0.150 ;
        RECT 4.980 -0.230 5.310 -0.180 ;
        RECT 4.980 -0.400 5.560 -0.230 ;
        RECT 4.980 -0.410 5.300 -0.400 ;
      LAYER mcon ;
        RECT 5.040 -0.360 5.210 -0.190 ;
      LAYER met1 ;
        RECT 4.970 -0.440 5.290 -0.120 ;
      LAYER via ;
        RECT 5.000 -0.410 5.260 -0.150 ;
      LAYER met2 ;
        RECT 4.970 -0.130 5.280 -0.120 ;
        RECT 4.970 -0.170 7.440 -0.130 ;
        RECT 4.880 -0.310 7.440 -0.170 ;
        RECT 4.970 -0.450 5.280 -0.310 ;
    END
  END DRAIN2
  PIN DRAIN3
    USE ANALOG ;
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER li1 ;
        RECT 4.980 -1.190 5.300 -1.180 ;
        RECT 4.980 -1.360 5.560 -1.190 ;
        RECT 4.980 -1.410 5.310 -1.360 ;
        RECT 4.980 -1.440 5.300 -1.410 ;
      LAYER mcon ;
        RECT 5.040 -1.400 5.210 -1.230 ;
      LAYER met1 ;
        RECT 4.970 -1.470 5.290 -1.150 ;
      LAYER via ;
        RECT 5.000 -1.440 5.260 -1.180 ;
      LAYER met2 ;
        RECT 4.970 -1.280 5.280 -1.140 ;
        RECT 4.970 -1.290 7.450 -1.280 ;
        RECT 4.850 -1.460 7.450 -1.290 ;
        RECT 4.970 -1.470 5.280 -1.460 ;
    END
  END DRAIN3
  PIN DRAIN4
    USE ANALOG ;
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER li1 ;
        RECT 4.980 -3.180 5.300 -3.150 ;
        RECT 4.980 -3.230 5.310 -3.180 ;
        RECT 4.980 -3.400 5.560 -3.230 ;
        RECT 4.980 -3.410 5.300 -3.400 ;
      LAYER mcon ;
        RECT 5.040 -3.360 5.210 -3.190 ;
      LAYER met1 ;
        RECT 4.970 -3.440 5.290 -3.120 ;
      LAYER via ;
        RECT 5.000 -3.410 5.260 -3.150 ;
      LAYER met2 ;
        RECT 4.970 -3.130 5.280 -3.120 ;
        RECT 4.870 -3.300 7.440 -3.130 ;
        RECT 4.970 -3.310 7.440 -3.300 ;
        RECT 4.970 -3.450 5.280 -3.310 ;
    END
  END DRAIN4
END sky130_hilas_swc4x1BiasCell

MACRO sky130_hilas_nMirror03
  CLASS BLOCK ;
  FOREIGN sky130_hilas_nMirror03 ;
  ORIGIN 0.590 0.050 ;
  SIZE 1.840 BY 1.270 ;
  OBS
      LAYER li1 ;
        RECT 0.000 1.040 0.200 1.080 ;
        RECT -0.230 0.780 0.200 1.040 ;
        RECT 0.000 0.750 0.200 0.780 ;
        RECT -0.410 0.390 -0.240 0.430 ;
        RECT 0.000 0.390 0.200 0.420 ;
        RECT -0.410 0.130 0.200 0.390 ;
        RECT -0.410 0.100 -0.240 0.130 ;
        RECT 0.000 0.090 0.200 0.130 ;
        RECT 0.590 0.090 1.140 1.080 ;
      LAYER mcon ;
        RECT -0.170 0.820 0.000 0.990 ;
        RECT 0.810 0.500 0.980 0.670 ;
        RECT -0.220 0.170 -0.050 0.340 ;
      LAYER met1 ;
        RECT -0.240 0.750 0.080 1.070 ;
        RECT 0.780 0.440 1.010 0.730 ;
        RECT -0.290 0.100 0.030 0.420 ;
      LAYER via ;
        RECT -0.210 0.780 0.050 1.040 ;
        RECT -0.260 0.130 0.000 0.390 ;
      LAYER met2 ;
        RECT -0.240 0.750 0.070 1.080 ;
        RECT -0.290 0.350 0.020 0.430 ;
        RECT -0.590 0.140 0.020 0.350 ;
        RECT -0.290 0.100 0.020 0.140 ;
  END
END sky130_hilas_nMirror03

MACRO sky130_hilas_FGHugeVaractorCapacitor01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_FGHugeVaractorCapacitor01 ;
  ORIGIN 5.560 8.160 ;
  SIZE 10.290 BY 5.990 ;
  OBS
      LAYER nwell ;
        RECT -5.560 -6.770 4.130 -2.170 ;
        RECT -5.560 -8.160 4.730 -6.770 ;
      LAYER li1 ;
        RECT 4.100 -7.860 4.270 -7.190 ;
      LAYER mcon ;
        RECT 4.100 -7.610 4.270 -7.440 ;
      LAYER met1 ;
        RECT 4.070 -7.700 4.310 -7.340 ;
  END
END sky130_hilas_FGHugeVaractorCapacitor01

MACRO sky130_hilas_nFETmirrorPairs
  CLASS BLOCK ;
  FOREIGN sky130_hilas_nFETmirrorPairs ;
  ORIGIN 0.330 1.920 ;
  SIZE 1.660 BY 2.750 ;
  OBS
      LAYER li1 ;
        RECT -0.050 0.640 0.220 0.830 ;
        RECT 0.850 0.650 1.100 0.830 ;
        RECT -0.080 0.470 0.250 0.640 ;
        RECT 0.770 0.470 1.100 0.650 ;
        RECT -0.120 -0.200 0.290 0.040 ;
        RECT 0.730 -0.200 1.140 0.040 ;
        RECT -0.120 -0.580 1.140 -0.200 ;
        RECT -0.120 -0.840 0.290 -0.580 ;
        RECT 0.730 -0.830 1.140 -0.580 ;
        RECT -0.090 -1.430 0.250 -1.260 ;
        RECT 0.760 -1.430 1.120 -1.250 ;
        RECT -0.010 -1.920 0.170 -1.430 ;
        RECT 0.840 -1.920 1.030 -1.430 ;
  END
END sky130_hilas_nFETmirrorPairs

MACRO sky130_hilas_DAC6TransistorStack01a
  CLASS BLOCK ;
  FOREIGN sky130_hilas_DAC6TransistorStack01a ;
  ORIGIN -0.280 1.740 ;
  SIZE 1.720 BY 5.650 ;
  OBS
      LAYER nwell ;
        RECT 0.280 -1.740 1.890 3.910 ;
  END
END sky130_hilas_DAC6TransistorStack01a

MACRO sky130_hilas_TgateSingle01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TgateSingle01 ;
  ORIGIN 2.630 1.810 ;
  SIZE 4.760 BY 1.520 ;
  OBS
      LAYER nwell ;
        RECT -2.510 -1.810 0.250 -0.290 ;
      LAYER li1 ;
        RECT -2.390 -0.830 -2.180 -0.400 ;
        RECT -1.880 -0.710 -1.690 -0.680 ;
        RECT 1.620 -0.700 1.810 -0.680 ;
        RECT -2.370 -0.850 -2.200 -0.830 ;
        RECT -1.880 -0.880 -1.360 -0.710 ;
        RECT -1.010 -0.880 0.890 -0.700 ;
        RECT 1.270 -0.710 1.810 -0.700 ;
        RECT 1.270 -0.870 2.050 -0.710 ;
        RECT -1.880 -0.960 -1.690 -0.880 ;
        RECT -1.900 -0.990 -1.690 -0.960 ;
        RECT -1.910 -1.000 -1.690 -0.990 ;
        RECT -0.520 -1.000 -0.190 -0.880 ;
        RECT 1.620 -0.910 2.050 -0.870 ;
        RECT -2.030 -1.050 -1.690 -1.000 ;
        RECT -2.160 -1.080 -1.690 -1.050 ;
        RECT -2.200 -1.110 -1.690 -1.080 ;
        RECT -2.200 -1.170 -1.710 -1.110 ;
        RECT -2.200 -1.220 -1.860 -1.170 ;
        RECT -2.200 -1.240 -1.940 -1.220 ;
        RECT -2.200 -1.260 -1.970 -1.240 ;
        RECT -2.200 -1.300 -1.990 -1.260 ;
        RECT -2.200 -1.580 -2.030 -1.300 ;
        RECT -0.850 -1.410 -0.680 -1.250 ;
        RECT 0.030 -1.320 0.220 -1.290 ;
        RECT 0.010 -1.330 0.220 -1.320 ;
        RECT -0.980 -1.450 -0.660 -1.410 ;
        RECT -0.980 -1.640 -0.650 -1.450 ;
        RECT -0.240 -1.500 0.220 -1.330 ;
        RECT 0.650 -1.410 0.820 -1.250 ;
        RECT 1.160 -1.330 1.350 -1.300 ;
        RECT 0.030 -1.520 0.220 -1.500 ;
        RECT 0.590 -1.450 0.910 -1.410 ;
        RECT 0.590 -1.640 0.920 -1.450 ;
        RECT 1.160 -1.500 1.600 -1.330 ;
        RECT 1.160 -1.530 1.350 -1.500 ;
        RECT 1.880 -1.590 2.050 -0.910 ;
        RECT -0.980 -1.670 -0.660 -1.640 ;
        RECT 0.590 -1.670 0.910 -1.640 ;
      LAYER mcon ;
        RECT -1.870 -0.880 -1.700 -0.710 ;
        RECT 1.630 -0.880 1.800 -0.710 ;
        RECT -0.920 -1.630 -0.750 -1.460 ;
        RECT 0.040 -1.490 0.210 -1.320 ;
        RECT 0.650 -1.630 0.820 -1.460 ;
        RECT 1.170 -1.500 1.340 -1.330 ;
      LAYER met1 ;
        RECT -2.390 -0.620 -2.050 -0.400 ;
        RECT -2.400 -0.720 -2.050 -0.620 ;
        RECT -1.890 -0.650 -1.690 -0.290 ;
        RECT -2.400 -0.910 -2.170 -0.720 ;
        RECT -1.900 -0.940 -1.670 -0.650 ;
        RECT -0.040 -0.790 0.220 -0.470 ;
        RECT 0.970 -0.530 1.230 -0.460 ;
        RECT 0.970 -0.780 1.330 -0.530 ;
        RECT 1.620 -0.650 1.810 -0.290 ;
        RECT -1.890 -1.810 -1.690 -0.940 ;
        RECT 0.030 -1.260 0.220 -0.790 ;
        RECT -0.990 -1.700 -0.670 -1.380 ;
        RECT 0.010 -1.550 0.240 -1.260 ;
        RECT 1.140 -1.270 1.330 -0.780 ;
        RECT 1.600 -0.940 1.830 -0.650 ;
        RECT 0.580 -1.700 0.900 -1.380 ;
        RECT 1.140 -1.560 1.370 -1.270 ;
        RECT 1.620 -1.810 1.810 -0.940 ;
      LAYER via ;
        RECT -2.310 -0.690 -2.050 -0.430 ;
        RECT -0.040 -0.760 0.220 -0.500 ;
        RECT 0.970 -0.750 1.230 -0.490 ;
        RECT -0.960 -1.670 -0.700 -1.410 ;
        RECT 0.610 -1.670 0.870 -1.410 ;
      LAYER met2 ;
        RECT -2.340 -0.520 -2.020 -0.430 ;
        RECT -0.070 -0.520 0.250 -0.500 ;
        RECT 0.940 -0.520 1.260 -0.490 ;
        RECT -2.630 -0.720 -2.020 -0.520 ;
        RECT -0.120 -0.720 2.130 -0.520 ;
        RECT -0.070 -0.760 0.250 -0.720 ;
        RECT 0.940 -0.750 1.260 -0.720 ;
        RECT -0.990 -1.490 -0.680 -1.370 ;
        RECT -1.760 -1.500 -0.640 -1.490 ;
        RECT 0.580 -1.500 0.890 -1.370 ;
        RECT -2.630 -1.700 0.890 -1.500 ;
        RECT -1.760 -1.710 -0.640 -1.700 ;
  END
END sky130_hilas_TgateSingle01

MACRO sky130_hilas_cellAttempt01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_cellAttempt01 ;
  ORIGIN 2.640 3.820 ;
  SIZE 10.080 BY 6.050 ;
  OBS
      LAYER nwell ;
        RECT -2.630 0.370 -0.900 2.230 ;
        RECT 4.880 2.220 7.430 2.230 ;
        RECT -2.640 -1.470 -0.900 0.370 ;
        RECT -2.630 -3.820 -0.900 -1.470 ;
        RECT 1.120 -3.810 3.350 2.220 ;
        RECT 4.880 -3.800 7.440 2.220 ;
        RECT 4.880 -3.810 7.430 -3.800 ;
      LAYER li1 ;
        RECT 4.980 1.820 5.300 1.830 ;
        RECT 4.980 1.650 5.560 1.820 ;
        RECT 4.980 1.600 5.310 1.650 ;
        RECT 4.980 1.570 5.300 1.600 ;
        RECT 6.840 1.550 7.040 1.900 ;
        RECT 4.980 1.240 5.300 1.280 ;
        RECT 4.980 1.200 5.310 1.240 ;
        RECT 4.980 1.030 5.560 1.200 ;
        RECT 4.980 1.020 5.300 1.030 ;
        RECT 6.110 0.960 6.310 1.530 ;
        RECT 6.840 1.520 7.050 1.550 ;
        RECT 6.830 0.930 7.050 1.520 ;
        RECT 4.980 0.390 5.300 0.400 ;
        RECT 4.980 0.220 5.560 0.390 ;
        RECT 4.980 0.180 5.310 0.220 ;
        RECT 4.980 0.140 5.300 0.180 ;
        RECT 6.110 -0.110 6.310 0.460 ;
        RECT 6.830 -0.100 7.050 0.490 ;
        RECT 6.840 -0.130 7.050 -0.100 ;
        RECT 4.980 -0.180 5.300 -0.150 ;
        RECT 4.980 -0.230 5.310 -0.180 ;
        RECT 4.980 -0.400 5.560 -0.230 ;
        RECT 4.980 -0.410 5.300 -0.400 ;
        RECT 6.840 -0.480 7.040 -0.130 ;
        RECT -2.210 -1.020 -1.660 -0.590 ;
        RECT 1.820 -1.090 2.370 -0.660 ;
        RECT 6.230 -0.880 6.670 -0.710 ;
        RECT 4.980 -1.190 5.300 -1.180 ;
        RECT 4.980 -1.360 5.560 -1.190 ;
        RECT 4.980 -1.410 5.310 -1.360 ;
        RECT 4.980 -1.440 5.300 -1.410 ;
        RECT 6.840 -1.460 7.040 -1.110 ;
        RECT 4.980 -1.770 5.300 -1.730 ;
        RECT 4.980 -1.810 5.310 -1.770 ;
        RECT 4.980 -1.980 5.560 -1.810 ;
        RECT 4.980 -1.990 5.300 -1.980 ;
        RECT 6.110 -2.050 6.310 -1.480 ;
        RECT 6.840 -1.490 7.050 -1.460 ;
        RECT 6.830 -2.080 7.050 -1.490 ;
        RECT 4.980 -2.610 5.300 -2.600 ;
        RECT 4.980 -2.780 5.560 -2.610 ;
        RECT 4.980 -2.820 5.310 -2.780 ;
        RECT 4.980 -2.860 5.300 -2.820 ;
        RECT 6.110 -3.110 6.310 -2.540 ;
        RECT 6.830 -3.100 7.050 -2.510 ;
        RECT 6.840 -3.130 7.050 -3.100 ;
        RECT 4.980 -3.180 5.300 -3.150 ;
        RECT 4.980 -3.230 5.310 -3.180 ;
        RECT 4.980 -3.400 5.560 -3.230 ;
        RECT 4.980 -3.410 5.300 -3.400 ;
        RECT 6.840 -3.480 7.040 -3.130 ;
      LAYER mcon ;
        RECT 5.040 1.610 5.210 1.780 ;
        RECT 6.120 1.320 6.290 1.490 ;
        RECT 5.040 1.060 5.210 1.230 ;
        RECT 6.850 1.350 7.020 1.520 ;
        RECT 5.040 0.190 5.210 0.360 ;
        RECT 6.120 -0.070 6.290 0.100 ;
        RECT 6.850 -0.100 7.020 0.070 ;
        RECT 5.040 -0.360 5.210 -0.190 ;
        RECT -2.210 -0.940 -1.940 -0.670 ;
        RECT 1.820 -1.010 2.090 -0.740 ;
        RECT 6.490 -0.880 6.670 -0.710 ;
        RECT 5.040 -1.400 5.210 -1.230 ;
        RECT 6.120 -1.690 6.290 -1.520 ;
        RECT 5.040 -1.950 5.210 -1.780 ;
        RECT 6.850 -1.660 7.020 -1.490 ;
        RECT 5.040 -2.810 5.210 -2.640 ;
        RECT 6.120 -3.070 6.290 -2.900 ;
        RECT 6.850 -3.100 7.020 -2.930 ;
        RECT 5.040 -3.360 5.210 -3.190 ;
      LAYER met1 ;
        RECT -2.280 -3.820 -1.880 2.170 ;
        RECT 1.770 0.310 2.150 2.230 ;
        RECT 4.970 1.540 5.290 1.860 ;
        RECT 6.110 1.550 6.270 2.230 ;
        RECT 6.110 1.530 6.310 1.550 ;
        RECT 4.970 0.990 5.290 1.310 ;
        RECT 6.090 1.290 6.320 1.530 ;
        RECT 6.110 1.070 6.310 1.290 ;
        RECT 6.480 1.240 6.670 2.230 ;
        RECT 6.920 1.580 7.080 2.230 ;
        RECT 6.500 1.120 6.670 1.240 ;
        RECT 1.760 -1.550 2.150 0.310 ;
        RECT 4.970 0.110 5.290 0.430 ;
        RECT 6.110 0.350 6.270 1.070 ;
        RECT 6.110 0.130 6.310 0.350 ;
        RECT 6.510 0.300 6.670 1.120 ;
        RECT 6.810 1.030 7.080 1.580 ;
        RECT 6.810 0.980 7.090 1.030 ;
        RECT 6.920 0.890 7.090 0.980 ;
        RECT 6.920 0.530 7.080 0.890 ;
        RECT 6.920 0.440 7.090 0.530 ;
        RECT 6.500 0.180 6.670 0.300 ;
        RECT 6.090 -0.110 6.320 0.130 ;
        RECT 4.970 -0.440 5.290 -0.120 ;
        RECT 6.110 -0.130 6.310 -0.110 ;
        RECT 4.970 -1.470 5.290 -1.150 ;
        RECT 6.110 -1.460 6.270 -0.130 ;
        RECT 6.480 -0.680 6.670 0.180 ;
        RECT 6.810 0.390 7.090 0.440 ;
        RECT 6.810 -0.160 7.080 0.390 ;
        RECT 6.460 -0.910 6.700 -0.680 ;
        RECT 6.110 -1.480 6.310 -1.460 ;
        RECT 1.770 -3.810 2.150 -1.550 ;
        RECT 4.970 -2.020 5.290 -1.700 ;
        RECT 6.090 -1.720 6.320 -1.480 ;
        RECT 6.110 -1.940 6.310 -1.720 ;
        RECT 6.480 -1.770 6.670 -0.910 ;
        RECT 6.920 -1.430 7.080 -0.160 ;
        RECT 6.500 -1.890 6.670 -1.770 ;
        RECT 4.970 -2.890 5.290 -2.570 ;
        RECT 6.110 -2.650 6.270 -1.940 ;
        RECT 6.110 -2.870 6.310 -2.650 ;
        RECT 6.510 -2.700 6.670 -1.890 ;
        RECT 6.810 -1.980 7.080 -1.430 ;
        RECT 6.810 -2.030 7.090 -1.980 ;
        RECT 6.920 -2.120 7.090 -2.030 ;
        RECT 6.920 -2.470 7.080 -2.120 ;
        RECT 6.920 -2.560 7.090 -2.470 ;
        RECT 6.500 -2.820 6.670 -2.700 ;
        RECT 6.090 -3.110 6.320 -2.870 ;
        RECT 4.970 -3.440 5.290 -3.120 ;
        RECT 6.110 -3.130 6.310 -3.110 ;
        RECT 6.110 -3.810 6.270 -3.130 ;
        RECT 6.480 -3.810 6.670 -2.820 ;
        RECT 6.810 -2.610 7.090 -2.560 ;
        RECT 6.810 -3.160 7.080 -2.610 ;
        RECT 6.920 -3.810 7.080 -3.160 ;
      LAYER via ;
        RECT 5.000 1.570 5.260 1.830 ;
        RECT 5.000 1.020 5.260 1.280 ;
        RECT 5.000 0.140 5.260 0.400 ;
        RECT 5.000 -0.410 5.260 -0.150 ;
        RECT 5.000 -1.440 5.260 -1.180 ;
        RECT 5.000 -1.990 5.260 -1.730 ;
        RECT 5.000 -2.860 5.260 -2.600 ;
        RECT 5.000 -3.410 5.260 -3.150 ;
      LAYER met2 ;
        RECT 4.970 1.730 5.280 1.870 ;
        RECT -2.640 1.550 7.440 1.730 ;
        RECT 4.970 1.540 5.280 1.550 ;
        RECT 4.970 1.300 5.280 1.320 ;
        RECT -2.640 1.120 7.440 1.300 ;
        RECT 4.970 0.990 5.280 1.120 ;
        RECT 4.970 0.300 5.280 0.430 ;
        RECT -2.640 0.120 7.440 0.300 ;
        RECT 4.970 0.100 5.280 0.120 ;
        RECT 4.970 -0.130 5.280 -0.120 ;
        RECT -2.640 -0.310 7.440 -0.130 ;
        RECT 4.970 -0.450 5.280 -0.310 ;
        RECT 4.970 -1.280 5.280 -1.140 ;
        RECT 4.970 -1.290 7.440 -1.280 ;
        RECT -2.620 -1.460 7.440 -1.290 ;
        RECT 4.970 -1.470 5.280 -1.460 ;
        RECT 4.970 -1.710 5.280 -1.690 ;
        RECT -2.620 -1.880 7.440 -1.710 ;
        RECT 4.880 -1.890 7.440 -1.880 ;
        RECT 4.970 -2.020 5.280 -1.890 ;
        RECT 4.970 -2.690 5.280 -2.570 ;
        RECT -2.620 -2.700 5.280 -2.690 ;
        RECT -2.620 -2.860 7.440 -2.700 ;
        RECT -1.840 -2.950 -0.300 -2.860 ;
        RECT 4.880 -2.880 7.440 -2.860 ;
        RECT 4.970 -2.900 5.280 -2.880 ;
        RECT 4.970 -3.130 5.280 -3.120 ;
        RECT -2.620 -3.300 7.440 -3.130 ;
        RECT 4.970 -3.310 7.440 -3.300 ;
        RECT 4.970 -3.450 5.280 -3.310 ;
  END
END sky130_hilas_cellAttempt01

MACRO sky130_hilas_TA2SignalBiasCell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TA2SignalBiasCell ;
  ORIGIN 5.260 -1.400 ;
  SIZE 8.450 BY 6.050 ;
  PIN VOUT_AMP2
    USE ANALOG ;
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER li1 ;
        RECT 0.510 4.990 0.710 5.020 ;
        RECT 0.280 4.730 0.710 4.990 ;
        RECT 2.580 4.910 2.900 4.950 ;
        RECT 2.580 4.850 2.910 4.910 ;
        RECT 0.510 4.690 0.710 4.730 ;
        RECT 2.110 4.720 2.910 4.850 ;
        RECT 2.110 4.690 2.900 4.720 ;
        RECT 2.110 4.670 2.810 4.690 ;
      LAYER mcon ;
        RECT 0.340 4.780 0.510 4.950 ;
        RECT 2.640 4.730 2.810 4.900 ;
      LAYER met1 ;
        RECT 0.270 4.700 0.590 5.020 ;
        RECT 2.570 4.660 2.890 4.980 ;
      LAYER via ;
        RECT 0.300 4.730 0.560 4.990 ;
        RECT 2.600 4.690 2.860 4.950 ;
      LAYER met2 ;
        RECT 0.270 4.970 0.580 5.020 ;
        RECT 2.570 4.970 2.880 4.990 ;
        RECT 0.270 4.740 3.190 4.970 ;
        RECT 0.270 4.690 0.580 4.740 ;
        RECT 2.570 4.660 2.880 4.740 ;
    END
  END VOUT_AMP2
  PIN VOUT_AMP1
    USE ANALOG ;
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER li1 ;
        RECT 0.510 4.160 0.710 4.200 ;
        RECT 2.570 4.190 2.890 4.230 ;
        RECT 0.280 3.900 0.710 4.160 ;
        RECT 2.110 4.010 2.900 4.190 ;
        RECT 2.570 4.000 2.900 4.010 ;
        RECT 2.570 3.970 2.890 4.000 ;
        RECT 0.510 3.870 0.710 3.900 ;
      LAYER mcon ;
        RECT 0.340 3.940 0.510 4.110 ;
        RECT 2.630 4.010 2.800 4.180 ;
      LAYER met1 ;
        RECT 0.270 3.870 0.590 4.190 ;
        RECT 2.560 3.940 2.880 4.260 ;
      LAYER via ;
        RECT 0.300 3.900 0.560 4.160 ;
        RECT 2.590 3.970 2.850 4.230 ;
      LAYER met2 ;
        RECT 0.270 4.140 0.580 4.200 ;
        RECT 2.560 4.140 2.870 4.270 ;
        RECT 0.270 3.920 3.190 4.140 ;
        RECT 0.270 3.870 0.580 3.920 ;
    END
  END VOUT_AMP1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 1.100 6.170 1.650 7.160 ;
        RECT 1.100 4.690 1.650 5.680 ;
        RECT 1.100 3.210 1.650 4.200 ;
        RECT 1.100 1.730 1.650 2.720 ;
      LAYER mcon ;
        RECT 1.320 6.580 1.490 6.750 ;
        RECT 1.320 5.100 1.490 5.270 ;
        RECT 1.320 3.620 1.490 3.790 ;
        RECT 1.320 2.140 1.490 2.310 ;
      LAYER met1 ;
        RECT 1.230 1.400 1.570 7.450 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 1.920 7.270 3.190 7.450 ;
        RECT 1.910 1.400 3.190 7.270 ;
      LAYER li1 ;
        RECT 2.120 5.840 2.820 6.150 ;
        RECT 1.970 5.610 2.820 5.840 ;
        RECT 2.120 5.270 2.820 5.610 ;
        RECT 2.120 3.250 2.820 3.590 ;
        RECT 1.970 3.020 2.820 3.250 ;
        RECT 2.120 2.710 2.820 3.020 ;
      LAYER mcon ;
        RECT 1.980 5.640 2.150 5.810 ;
        RECT 1.980 3.050 2.150 3.220 ;
      LAYER met1 ;
        RECT 1.900 5.870 2.170 7.450 ;
        RECT 1.900 5.580 2.180 5.870 ;
        RECT 1.900 3.280 2.170 5.580 ;
        RECT 1.900 2.990 2.180 3.280 ;
        RECT 1.900 1.400 2.170 2.990 ;
    END
    PORT
      LAYER li1 ;
        RECT -4.850 6.960 -4.670 6.980 ;
        RECT -4.930 6.920 -4.610 6.960 ;
        RECT -4.930 6.730 -4.600 6.920 ;
        RECT -4.930 6.700 -4.610 6.730 ;
        RECT -4.850 3.070 -4.670 6.700 ;
        RECT -4.970 3.030 -4.650 3.070 ;
        RECT -4.970 2.840 -4.640 3.030 ;
        RECT -4.970 2.810 -4.650 2.840 ;
        RECT -4.850 1.880 -4.670 2.810 ;
      LAYER mcon ;
        RECT -4.870 6.740 -4.700 6.910 ;
        RECT -4.910 2.850 -4.740 3.020 ;
      LAYER met1 ;
        RECT -4.940 6.670 -4.620 6.990 ;
        RECT -4.980 2.780 -4.660 3.100 ;
      LAYER via ;
        RECT -4.910 6.700 -4.650 6.960 ;
        RECT -4.950 2.810 -4.690 3.070 ;
      LAYER met2 ;
        RECT -4.900 7.000 -4.660 7.450 ;
        RECT -4.940 6.670 -4.630 7.000 ;
        RECT -4.980 2.780 -4.670 3.110 ;
    END
  END VPWR
  PIN VINN_AMP2
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER li1 ;
        RECT -0.960 7.400 -0.790 7.450 ;
        RECT -0.960 7.140 -0.400 7.400 ;
        RECT -0.960 7.120 -0.790 7.140 ;
      LAYER mcon ;
        RECT -0.630 7.180 -0.460 7.350 ;
      LAYER met1 ;
        RECT -0.710 7.110 -0.390 7.430 ;
      LAYER via ;
        RECT -0.680 7.140 -0.420 7.400 ;
      LAYER met2 ;
        RECT -1.300 7.430 -1.050 7.440 ;
        RECT -0.700 7.430 -0.390 7.440 ;
        RECT -1.300 7.180 -0.390 7.430 ;
        RECT -0.700 7.110 -0.390 7.180 ;
    END
  END VINN_AMP2
  PIN VINP_AMP2
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER li1 ;
        RECT -0.930 4.730 -0.610 4.760 ;
        RECT -0.930 4.540 -0.600 4.730 ;
        RECT -0.930 4.500 -0.610 4.540 ;
        RECT -0.930 4.420 -0.760 4.500 ;
        RECT -0.980 4.250 -0.760 4.420 ;
        RECT -0.980 4.090 -0.810 4.250 ;
      LAYER mcon ;
        RECT -0.870 4.550 -0.700 4.720 ;
      LAYER met1 ;
        RECT -0.940 4.470 -0.620 4.790 ;
      LAYER via ;
        RECT -0.910 4.500 -0.650 4.760 ;
      LAYER met2 ;
        RECT -0.940 4.750 -0.630 4.790 ;
        RECT -1.030 4.740 -0.600 4.750 ;
        RECT -1.260 4.510 -0.160 4.740 ;
        RECT -0.940 4.460 -0.630 4.510 ;
    END
  END VINP_AMP2
  PIN VINP_AMP1
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER li1 ;
        RECT -2.540 4.600 -2.370 4.760 ;
        RECT -2.540 4.430 -2.320 4.600 ;
        RECT -2.490 4.350 -2.320 4.430 ;
        RECT -2.490 4.310 -2.170 4.350 ;
        RECT -2.490 4.120 -2.160 4.310 ;
        RECT -2.490 4.090 -2.170 4.120 ;
      LAYER mcon ;
        RECT -2.430 4.130 -2.260 4.300 ;
      LAYER met1 ;
        RECT -2.500 4.060 -2.180 4.380 ;
      LAYER via ;
        RECT -2.470 4.090 -2.210 4.350 ;
      LAYER met2 ;
        RECT -2.500 4.340 -2.190 4.390 ;
        RECT -2.820 4.110 -1.720 4.340 ;
        RECT -2.820 4.100 -2.160 4.110 ;
        RECT -2.500 4.060 -2.190 4.100 ;
    END
  END VINP_AMP1
  PIN VINN_AMP1
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER li1 ;
        RECT -2.520 1.710 -2.350 1.730 ;
        RECT -2.520 1.450 -1.960 1.710 ;
        RECT -2.520 1.400 -2.350 1.450 ;
      LAYER mcon ;
        RECT -2.190 1.500 -2.020 1.670 ;
      LAYER met1 ;
        RECT -2.270 1.420 -1.950 1.740 ;
      LAYER via ;
        RECT -2.240 1.450 -1.980 1.710 ;
      LAYER met2 ;
        RECT -2.260 1.670 -1.950 1.740 ;
        RECT -2.860 1.420 -1.950 1.670 ;
        RECT -2.260 1.410 -1.950 1.420 ;
    END
  END VINN_AMP1
  PIN VBIAS2
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER li1 ;
        RECT -4.270 1.710 -4.100 1.730 ;
        RECT -4.270 1.450 -3.710 1.710 ;
        RECT -4.270 1.400 -4.100 1.450 ;
      LAYER mcon ;
        RECT -3.940 1.500 -3.770 1.670 ;
      LAYER met1 ;
        RECT -4.020 1.420 -3.700 1.740 ;
      LAYER via ;
        RECT -3.990 1.450 -3.730 1.710 ;
      LAYER met2 ;
        RECT -4.010 1.670 -3.700 1.740 ;
        RECT -4.580 1.660 -3.700 1.670 ;
        RECT -5.260 1.430 -3.700 1.660 ;
        RECT -4.580 1.420 -3.700 1.430 ;
        RECT -4.010 1.410 -3.700 1.420 ;
    END
  END VBIAS2
  PIN VBIAS1
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER li1 ;
        RECT -4.290 4.600 -4.120 4.760 ;
        RECT -4.290 4.430 -4.070 4.600 ;
        RECT -4.240 4.350 -4.070 4.430 ;
        RECT -4.240 4.310 -3.920 4.350 ;
        RECT -4.240 4.120 -3.910 4.310 ;
        RECT -4.240 4.090 -3.920 4.120 ;
      LAYER mcon ;
        RECT -4.180 4.130 -4.010 4.300 ;
      LAYER met1 ;
        RECT -4.250 4.060 -3.930 4.380 ;
      LAYER via ;
        RECT -4.220 4.090 -3.960 4.350 ;
      LAYER met2 ;
        RECT -4.250 4.340 -3.940 4.390 ;
        RECT -5.260 4.110 -3.470 4.340 ;
        RECT -5.260 4.100 -3.910 4.110 ;
        RECT -4.250 4.060 -3.940 4.100 ;
    END
  END VBIAS1
  OBS
      LAYER nwell ;
        RECT -5.260 7.440 -1.650 7.450 ;
        RECT -5.260 1.410 -0.090 7.440 ;
        RECT -1.950 1.400 -0.090 1.410 ;
      LAYER li1 ;
        RECT 0.510 7.120 0.710 7.160 ;
        RECT -4.040 5.950 -3.870 6.970 ;
        RECT -4.090 5.910 -3.770 5.950 ;
        RECT -4.090 5.720 -3.760 5.910 ;
        RECT -4.090 5.690 -3.770 5.720 ;
        RECT -4.040 5.190 -3.870 5.690 ;
        RECT -4.120 5.130 -3.580 5.190 ;
        RECT -4.120 5.020 -3.570 5.130 ;
        RECT -3.760 4.900 -3.570 5.020 ;
        RECT -4.040 2.540 -3.870 3.920 ;
        RECT -3.100 3.070 -2.920 6.980 ;
        RECT -2.290 5.190 -2.120 6.970 ;
        RECT -1.540 6.040 -1.360 6.970 ;
        RECT -0.810 6.710 -0.480 6.880 ;
        RECT 0.280 6.860 0.710 7.120 ;
        RECT 0.510 6.830 0.710 6.860 ;
        RECT 2.470 7.040 3.050 7.210 ;
        RECT 2.470 6.940 2.860 7.040 ;
        RECT 2.470 6.910 2.850 6.940 ;
        RECT 2.470 6.760 2.830 6.910 ;
        RECT -0.730 6.570 -0.480 6.710 ;
        RECT 2.120 6.590 2.830 6.760 ;
        RECT -0.730 6.310 -0.250 6.570 ;
        RECT 0.100 6.470 0.270 6.510 ;
        RECT 0.510 6.470 0.710 6.500 ;
        RECT -1.660 6.010 -1.340 6.040 ;
        RECT -1.660 5.820 -1.330 6.010 ;
        RECT -1.660 5.780 -1.340 5.820 ;
        RECT -2.370 5.130 -1.830 5.190 ;
        RECT -2.370 5.020 -1.820 5.130 ;
        RECT -2.010 4.900 -1.820 5.020 ;
        RECT -3.220 3.030 -2.900 3.070 ;
        RECT -3.220 2.840 -2.890 3.030 ;
        RECT -3.220 2.810 -2.900 2.840 ;
        RECT -4.040 2.280 -3.560 2.540 ;
        RECT -4.040 2.140 -3.790 2.280 ;
        RECT -4.120 1.970 -3.790 2.140 ;
        RECT -3.100 1.880 -2.920 2.810 ;
        RECT -2.290 2.540 -2.120 3.920 ;
        RECT -2.290 2.280 -1.810 2.540 ;
        RECT -2.290 2.140 -2.040 2.280 ;
        RECT -2.370 1.970 -2.040 2.140 ;
        RECT -1.540 1.870 -1.360 5.780 ;
        RECT -0.730 4.930 -0.560 6.310 ;
        RECT 0.100 6.210 0.710 6.470 ;
        RECT 0.100 6.180 0.270 6.210 ;
        RECT 0.510 6.170 0.710 6.210 ;
        RECT 0.100 5.640 0.270 5.670 ;
        RECT 0.510 5.640 0.710 5.680 ;
        RECT 0.100 5.380 0.710 5.640 ;
        RECT 0.100 5.340 0.270 5.380 ;
        RECT 0.510 5.350 0.710 5.380 ;
        RECT -0.450 3.830 -0.260 3.950 ;
        RECT -0.810 3.720 -0.260 3.830 ;
        RECT -0.810 3.660 -0.270 3.720 ;
        RECT -0.730 1.880 -0.560 3.660 ;
        RECT 0.100 3.510 0.270 3.550 ;
        RECT 0.510 3.510 0.710 3.540 ;
        RECT 0.100 3.250 0.710 3.510 ;
        RECT 0.100 3.220 0.270 3.250 ;
        RECT 0.510 3.210 0.710 3.250 ;
        RECT 0.100 2.680 0.270 2.710 ;
        RECT 0.510 2.680 0.710 2.720 ;
        RECT 0.100 2.420 0.710 2.680 ;
        RECT 0.100 2.380 0.270 2.420 ;
        RECT 0.510 2.390 0.710 2.420 ;
        RECT 2.120 2.100 2.830 2.270 ;
        RECT 0.510 2.030 0.710 2.060 ;
        RECT 0.280 1.770 0.710 2.030 ;
        RECT 0.510 1.730 0.710 1.770 ;
        RECT 2.470 1.820 2.830 2.100 ;
        RECT 2.470 1.650 3.050 1.820 ;
      LAYER mcon ;
        RECT -4.030 5.730 -3.860 5.900 ;
        RECT -3.750 4.930 -3.580 5.100 ;
        RECT 0.340 6.900 0.510 7.070 ;
        RECT 2.590 6.950 2.760 7.120 ;
        RECT -0.480 6.350 -0.310 6.520 ;
        RECT -1.600 5.830 -1.430 6.000 ;
        RECT -2.000 4.930 -1.830 5.100 ;
        RECT -3.160 2.850 -2.990 3.020 ;
        RECT -3.790 2.330 -3.620 2.500 ;
        RECT -2.040 2.330 -1.870 2.500 ;
        RECT 0.290 6.250 0.460 6.420 ;
        RECT 0.290 5.430 0.460 5.600 ;
        RECT -0.440 3.750 -0.270 3.920 ;
        RECT 0.290 3.290 0.460 3.460 ;
        RECT 0.290 2.470 0.460 2.640 ;
        RECT 0.340 1.820 0.510 1.990 ;
        RECT 2.550 1.760 2.720 1.930 ;
      LAYER met1 ;
        RECT 0.270 6.830 0.590 7.150 ;
        RECT 2.520 6.880 2.840 7.200 ;
        RECT -0.560 6.280 -0.240 6.600 ;
        RECT 0.220 6.180 0.540 6.500 ;
        RECT -4.100 5.660 -3.780 5.980 ;
        RECT -1.670 5.750 -1.350 6.070 ;
        RECT -0.450 5.590 -0.240 5.700 ;
        RECT -0.470 5.270 -0.210 5.590 ;
        RECT 0.220 5.350 0.540 5.670 ;
        RECT -3.780 4.870 -3.550 5.160 ;
        RECT -2.030 4.870 -1.800 5.160 ;
        RECT -3.760 3.580 -3.550 4.870 ;
        RECT -2.010 3.580 -1.800 4.870 ;
        RECT -0.450 3.980 -0.240 5.270 ;
        RECT -0.470 3.690 -0.240 3.980 ;
        RECT -3.780 3.260 -3.520 3.580 ;
        RECT -2.030 3.260 -1.770 3.580 ;
        RECT -3.760 3.150 -3.550 3.260 ;
        RECT -2.010 3.150 -1.800 3.260 ;
        RECT 0.220 3.220 0.540 3.540 ;
        RECT -3.230 2.780 -2.910 3.100 ;
        RECT -3.870 2.250 -3.550 2.570 ;
        RECT -2.120 2.250 -1.800 2.570 ;
        RECT 0.220 2.390 0.540 2.710 ;
        RECT 0.270 1.740 0.590 2.060 ;
        RECT 2.480 1.690 2.800 2.010 ;
      LAYER via ;
        RECT 0.300 6.860 0.560 7.120 ;
        RECT 2.550 6.910 2.810 7.170 ;
        RECT -0.530 6.310 -0.270 6.570 ;
        RECT 0.250 6.210 0.510 6.470 ;
        RECT -4.070 5.690 -3.810 5.950 ;
        RECT -1.640 5.780 -1.380 6.040 ;
        RECT -0.470 5.300 -0.210 5.560 ;
        RECT 0.250 5.380 0.510 5.640 ;
        RECT -3.780 3.290 -3.520 3.550 ;
        RECT -2.030 3.290 -1.770 3.550 ;
        RECT 0.250 3.250 0.510 3.510 ;
        RECT -3.200 2.810 -2.940 3.070 ;
        RECT -3.840 2.280 -3.580 2.540 ;
        RECT -2.090 2.280 -1.830 2.540 ;
        RECT 0.250 2.420 0.510 2.680 ;
        RECT 0.300 1.770 0.560 2.030 ;
        RECT 2.510 1.720 2.770 1.980 ;
      LAYER met2 ;
        RECT 0.270 7.110 0.580 7.160 ;
        RECT 2.520 7.110 2.830 7.210 ;
        RECT 0.270 6.880 2.830 7.110 ;
        RECT 0.270 6.830 0.580 6.880 ;
        RECT -0.550 6.570 -0.240 6.610 ;
        RECT -0.730 6.430 0.010 6.570 ;
        RECT 0.220 6.430 0.530 6.510 ;
        RECT -0.730 6.320 0.530 6.430 ;
        RECT -0.550 6.280 0.530 6.320 ;
        RECT -0.240 6.220 0.530 6.280 ;
        RECT -0.240 6.200 0.010 6.220 ;
        RECT 0.220 6.180 0.530 6.220 ;
        RECT -4.100 5.930 -3.790 5.990 ;
        RECT -1.670 5.930 -1.360 6.070 ;
        RECT -4.100 5.740 -1.360 5.930 ;
        RECT -4.100 5.710 -1.620 5.740 ;
        RECT -4.100 5.660 -3.790 5.710 ;
        RECT -0.210 5.630 0.000 5.640 ;
        RECT 0.220 5.630 0.530 5.670 ;
        RECT -0.210 5.560 0.530 5.630 ;
        RECT -0.500 5.540 0.530 5.560 ;
        RECT -0.550 5.420 0.530 5.540 ;
        RECT -0.550 5.350 0.000 5.420 ;
        RECT -0.550 5.290 -0.080 5.350 ;
        RECT 0.220 5.340 0.530 5.420 ;
        RECT -3.860 3.310 -3.390 3.560 ;
        RECT -2.110 3.470 -1.640 3.560 ;
        RECT 0.220 3.470 0.530 3.550 ;
        RECT -2.110 3.310 0.530 3.470 ;
        RECT -3.810 3.290 -3.490 3.310 ;
        RECT -2.060 3.290 0.530 3.310 ;
        RECT -1.770 3.270 0.530 3.290 ;
        RECT -0.080 3.260 0.530 3.270 ;
        RECT 0.220 3.220 0.530 3.260 ;
        RECT -3.230 3.100 -2.920 3.110 ;
        RECT -3.340 2.920 -2.920 3.100 ;
        RECT -3.360 2.910 -2.920 2.920 ;
        RECT -3.580 2.780 -2.920 2.910 ;
        RECT -3.580 2.570 -3.220 2.780 ;
        RECT 0.220 2.670 0.530 2.710 ;
        RECT -2.060 2.570 0.530 2.670 ;
        RECT -3.860 2.530 -3.220 2.570 ;
        RECT -2.110 2.530 0.530 2.570 ;
        RECT -4.040 2.290 -3.220 2.530 ;
        RECT -2.290 2.460 0.530 2.530 ;
        RECT -4.040 2.280 -3.490 2.290 ;
        RECT -2.290 2.280 -1.740 2.460 ;
        RECT 0.220 2.380 0.530 2.460 ;
        RECT -3.860 2.240 -3.550 2.280 ;
        RECT -2.110 2.240 -1.800 2.280 ;
        RECT 0.270 1.980 0.580 2.060 ;
        RECT 2.480 1.980 2.790 2.020 ;
        RECT 0.270 1.750 2.980 1.980 ;
        RECT 0.270 1.730 0.580 1.750 ;
        RECT 2.480 1.690 2.790 1.750 ;
  END
END sky130_hilas_TA2SignalBiasCell

MACRO sky130_hilas_WTA4stage01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_WTA4stage01 ;
  ORIGIN 0.540 -0.010 ;
  SIZE 2.830 BY 5.340 ;
  OBS
      LAYER li1 ;
        RECT -0.430 5.290 -0.110 5.320 ;
        RECT -0.430 5.120 1.360 5.290 ;
        RECT -0.430 5.100 -0.100 5.120 ;
        RECT -0.430 5.060 -0.110 5.100 ;
        RECT 1.190 4.890 1.360 5.120 ;
        RECT 0.040 4.640 0.380 4.890 ;
        RECT 0.550 4.720 0.880 4.890 ;
        RECT 1.100 4.720 1.440 4.890 ;
        RECT -0.280 4.380 0.380 4.640 ;
        RECT 0.630 4.550 0.800 4.720 ;
        RECT 1.190 4.550 1.360 4.720 ;
        RECT 0.550 4.380 0.880 4.550 ;
        RECT 1.100 4.380 1.440 4.550 ;
        RECT 0.630 4.150 0.880 4.380 ;
        RECT 1.760 4.300 2.270 4.970 ;
        RECT 0.630 3.980 1.300 4.150 ;
        RECT 0.630 3.750 0.880 3.980 ;
        RECT -0.280 3.490 0.380 3.750 ;
        RECT 0.550 3.580 0.880 3.750 ;
        RECT 1.100 3.580 1.440 3.750 ;
        RECT 0.040 3.240 0.380 3.490 ;
        RECT 0.630 3.410 0.800 3.580 ;
        RECT 1.190 3.410 1.360 3.580 ;
        RECT 0.550 3.240 0.880 3.410 ;
        RECT 1.100 3.240 1.440 3.410 ;
        RECT -0.430 3.030 -0.110 3.070 ;
        RECT -0.430 3.010 -0.100 3.030 ;
        RECT 1.190 3.010 1.360 3.240 ;
        RECT 1.760 3.160 2.270 3.830 ;
        RECT -0.430 2.840 1.360 3.010 ;
        RECT -0.430 2.810 -0.110 2.840 ;
        RECT -0.430 2.520 -0.110 2.550 ;
        RECT -0.430 2.350 1.360 2.520 ;
        RECT -0.430 2.330 -0.100 2.350 ;
        RECT -0.430 2.290 -0.110 2.330 ;
        RECT 1.190 2.120 1.360 2.350 ;
        RECT 0.040 1.870 0.380 2.120 ;
        RECT 0.550 1.950 0.880 2.120 ;
        RECT 1.100 1.950 1.440 2.120 ;
        RECT -0.280 1.610 0.380 1.870 ;
        RECT 0.630 1.780 0.800 1.950 ;
        RECT 1.190 1.780 1.360 1.950 ;
        RECT 0.550 1.610 0.880 1.780 ;
        RECT 1.100 1.610 1.440 1.780 ;
        RECT 0.630 1.380 0.880 1.610 ;
        RECT 1.760 1.530 2.270 2.200 ;
        RECT 0.630 1.210 1.300 1.380 ;
        RECT 0.630 0.980 0.880 1.210 ;
        RECT -0.280 0.720 0.380 0.980 ;
        RECT 0.550 0.810 0.880 0.980 ;
        RECT 1.100 0.810 1.440 0.980 ;
        RECT 0.040 0.470 0.380 0.720 ;
        RECT 0.630 0.640 0.800 0.810 ;
        RECT 1.190 0.640 1.360 0.810 ;
        RECT 0.550 0.470 0.880 0.640 ;
        RECT 1.100 0.470 1.440 0.640 ;
        RECT -0.430 0.260 -0.110 0.300 ;
        RECT -0.430 0.240 -0.100 0.260 ;
        RECT 1.190 0.240 1.360 0.470 ;
        RECT 1.760 0.390 2.270 1.060 ;
        RECT -0.430 0.070 1.360 0.240 ;
        RECT -0.430 0.040 -0.110 0.070 ;
      LAYER mcon ;
        RECT -0.370 5.110 -0.200 5.280 ;
        RECT -0.220 4.430 -0.050 4.600 ;
        RECT 1.930 4.550 2.100 4.720 ;
        RECT 0.670 3.980 0.840 4.150 ;
        RECT -0.220 3.530 -0.050 3.700 ;
        RECT 1.930 3.410 2.100 3.580 ;
        RECT -0.370 2.850 -0.200 3.020 ;
        RECT -0.370 2.340 -0.200 2.510 ;
        RECT -0.220 1.660 -0.050 1.830 ;
        RECT 1.930 1.780 2.100 1.950 ;
        RECT 0.670 1.210 0.840 1.380 ;
        RECT -0.220 0.760 -0.050 0.930 ;
        RECT 1.930 0.640 2.100 0.810 ;
        RECT -0.370 0.080 -0.200 0.250 ;
      LAYER met1 ;
        RECT -0.440 5.030 -0.120 5.350 ;
        RECT -0.290 4.350 0.030 4.670 ;
        RECT -0.290 3.460 0.030 3.780 ;
        RECT -0.440 2.780 -0.120 3.100 ;
        RECT -0.440 2.260 -0.120 2.580 ;
        RECT -0.290 1.580 0.030 1.900 ;
        RECT -0.290 0.690 0.030 1.010 ;
        RECT -0.440 0.010 -0.120 0.330 ;
        RECT 0.640 0.010 0.870 5.350 ;
        RECT 1.900 0.010 2.130 5.350 ;
      LAYER via ;
        RECT -0.410 5.060 -0.150 5.320 ;
        RECT -0.260 4.380 0.000 4.640 ;
        RECT -0.260 3.490 0.000 3.750 ;
        RECT -0.410 2.810 -0.150 3.070 ;
        RECT -0.410 2.290 -0.150 2.550 ;
        RECT -0.260 1.610 0.000 1.870 ;
        RECT -0.260 0.720 0.000 0.980 ;
        RECT -0.410 0.040 -0.150 0.300 ;
      LAYER met2 ;
        RECT -0.440 5.310 -0.130 5.350 ;
        RECT -0.540 5.100 -0.130 5.310 ;
        RECT -0.440 5.020 -0.130 5.100 ;
        RECT -0.290 4.610 0.020 4.670 ;
        RECT -0.290 4.450 2.290 4.610 ;
        RECT -0.290 4.340 0.020 4.450 ;
        RECT -0.290 3.680 0.020 3.790 ;
        RECT -0.290 3.520 2.290 3.680 ;
        RECT -0.290 3.460 0.020 3.520 ;
        RECT -0.440 3.030 -0.130 3.110 ;
        RECT -0.540 2.820 -0.130 3.030 ;
        RECT -0.440 2.780 -0.130 2.820 ;
        RECT -0.440 2.540 -0.130 2.580 ;
        RECT -0.540 2.330 -0.130 2.540 ;
        RECT -0.440 2.250 -0.130 2.330 ;
        RECT -0.290 1.840 0.020 1.900 ;
        RECT -0.290 1.680 2.290 1.840 ;
        RECT -0.290 1.570 0.020 1.680 ;
        RECT -0.290 0.910 0.020 1.020 ;
        RECT -0.290 0.750 2.290 0.910 ;
        RECT -0.290 0.690 0.020 0.750 ;
        RECT -0.440 0.260 -0.130 0.340 ;
        RECT -0.540 0.050 -0.130 0.260 ;
        RECT -0.440 0.010 -0.130 0.050 ;
  END
END sky130_hilas_WTA4stage01

MACRO sky130_hilas_TgateVinj01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TgateVinj01 ;
  ORIGIN 2.100 0.400 ;
  SIZE 5.420 BY 1.590 ;
  OBS
      LAYER nwell ;
        RECT -2.100 -0.400 1.100 1.190 ;
      LAYER li1 ;
        RECT -1.700 -0.070 -1.530 0.860 ;
        RECT 2.580 0.790 2.770 0.830 ;
        RECT -1.000 0.620 1.750 0.790 ;
        RECT 2.210 0.620 2.770 0.790 ;
        RECT -0.560 0.440 -0.230 0.620 ;
        RECT 2.580 0.600 2.770 0.620 ;
        RECT 2.940 0.690 3.110 1.040 ;
        RECT 2.940 0.520 3.170 0.690 ;
        RECT 2.940 0.480 3.110 0.520 ;
        RECT -0.720 0.170 -0.550 0.180 ;
        RECT 1.990 0.170 2.230 0.210 ;
        RECT -1.000 0.000 -0.040 0.170 ;
        RECT 0.410 0.000 1.750 0.170 ;
        RECT 1.990 0.000 2.560 0.170 ;
        RECT 1.990 -0.030 2.230 0.000 ;
      LAYER mcon ;
        RECT 2.590 0.630 2.760 0.800 ;
        RECT -1.700 0.330 -1.530 0.500 ;
        RECT 3.000 0.520 3.170 0.690 ;
        RECT -0.720 0.010 -0.550 0.180 ;
        RECT 1.280 0.000 1.450 0.170 ;
        RECT 2.030 0.000 2.200 0.170 ;
      LAYER met1 ;
        RECT -1.740 -0.400 -1.490 1.190 ;
        RECT -0.590 0.210 -0.250 0.250 ;
        RECT -0.810 0.170 -0.250 0.210 ;
        RECT -0.810 0.000 -0.130 0.170 ;
        RECT -0.810 -0.020 -0.250 0.000 ;
        RECT -0.590 -0.070 -0.250 -0.020 ;
        RECT 1.250 -0.400 1.480 1.190 ;
        RECT 2.600 0.860 2.790 1.190 ;
        RECT 2.560 0.570 2.790 0.860 ;
        RECT 1.840 0.220 2.210 0.230 ;
        RECT 1.840 -0.040 2.260 0.220 ;
        RECT 1.840 -0.060 2.210 -0.040 ;
        RECT 2.600 -0.400 2.790 0.570 ;
        RECT 2.940 0.480 3.320 0.720 ;
      LAYER via ;
        RECT -0.540 -0.040 -0.280 0.220 ;
        RECT 1.870 -0.040 2.130 0.220 ;
      LAYER met2 ;
        RECT -0.570 0.170 -0.250 0.220 ;
        RECT 1.840 0.170 2.160 0.250 ;
        RECT -0.570 -0.020 2.160 0.170 ;
        RECT -0.570 -0.040 -0.250 -0.020 ;
        RECT 1.840 -0.070 2.160 -0.020 ;
  END
END sky130_hilas_TgateVinj01

MACRO sky130_hilas_capacitorSize04
  CLASS BLOCK ;
  FOREIGN sky130_hilas_capacitorSize04 ;
  ORIGIN -14.150 0.180 ;
  SIZE 5.780 BY 5.290 ;
  PIN CAP1TERM02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 19.240 4.130 19.610 4.190 ;
        RECT 19.240 3.850 19.920 4.130 ;
        RECT 19.240 3.790 19.610 3.850 ;
      LAYER via2 ;
        RECT 19.290 3.850 19.570 4.130 ;
      LAYER met3 ;
        RECT 15.860 4.340 18.160 5.110 ;
        RECT 15.860 3.590 19.810 4.340 ;
        RECT 15.860 2.830 18.160 3.590 ;
      LAYER via3 ;
        RECT 19.210 3.740 19.640 4.220 ;
      LAYER met4 ;
        RECT 19.110 3.650 19.770 4.310 ;
    END
  END CAP1TERM02
  PIN CAP2TERM02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 19.240 1.130 19.610 1.190 ;
        RECT 19.240 0.850 19.930 1.130 ;
        RECT 19.240 0.790 19.610 0.850 ;
      LAYER via2 ;
        RECT 19.290 0.850 19.570 1.130 ;
      LAYER met3 ;
        RECT 15.860 1.330 18.160 2.100 ;
        RECT 19.020 1.330 19.810 1.340 ;
        RECT 15.860 0.600 19.810 1.330 ;
        RECT 15.860 -0.180 18.160 0.600 ;
        RECT 19.020 0.590 19.810 0.600 ;
      LAYER via3 ;
        RECT 19.210 0.740 19.640 1.220 ;
      LAYER met4 ;
        RECT 19.110 0.650 19.770 1.310 ;
    END
  END CAP2TERM02
  PIN CAP2TERM01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 14.400 1.130 14.770 1.190 ;
        RECT 14.170 0.850 14.770 1.130 ;
        RECT 14.400 0.790 14.770 0.850 ;
      LAYER via2 ;
        RECT 14.450 0.850 14.730 1.130 ;
      LAYER met3 ;
        RECT 14.180 0.590 14.970 1.340 ;
      LAYER via3 ;
        RECT 14.370 0.740 14.800 1.220 ;
      LAYER met4 ;
        RECT 14.270 1.050 14.930 1.310 ;
        RECT 16.710 1.050 17.160 1.060 ;
        RECT 14.270 0.650 17.210 1.050 ;
        RECT 14.720 0.640 17.210 0.650 ;
        RECT 16.690 0.560 17.210 0.640 ;
    END
  END CAP2TERM01
  PIN CAP1TERM01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 14.370 4.130 14.740 4.190 ;
        RECT 14.170 3.850 14.740 4.130 ;
        RECT 14.370 3.790 14.740 3.850 ;
      LAYER via2 ;
        RECT 14.420 3.850 14.700 4.130 ;
      LAYER met3 ;
        RECT 14.150 3.590 14.940 4.340 ;
      LAYER via3 ;
        RECT 14.340 3.740 14.770 4.220 ;
      LAYER met4 ;
        RECT 14.240 4.060 14.900 4.310 ;
        RECT 16.710 4.060 17.160 4.070 ;
        RECT 14.240 3.650 17.210 4.060 ;
        RECT 16.690 3.570 17.210 3.650 ;
    END
  END CAP1TERM01
  OBS
      LAYER met2 ;
        RECT 14.170 4.800 19.920 4.980 ;
        RECT 14.170 4.370 19.920 4.550 ;
        RECT 14.170 3.370 19.920 3.550 ;
        RECT 14.170 2.940 19.920 3.120 ;
        RECT 14.170 1.790 19.920 1.960 ;
        RECT 14.170 1.370 19.920 1.540 ;
        RECT 14.170 0.390 19.920 0.560 ;
        RECT 14.170 -0.050 19.920 0.120 ;
  END
END sky130_hilas_capacitorSize04

MACRO sky130_hilas_TAcoreblock
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TAcoreblock ;
  ORIGIN -4.630 -1.990 ;
  SIZE 2.190 BY 4.770 ;
  OBS
      LAYER nwell ;
        RECT 4.630 5.030 6.820 6.760 ;
      LAYER li1 ;
        RECT 4.840 5.920 6.600 6.440 ;
        RECT 4.840 5.310 5.550 5.480 ;
        RECT 5.860 5.310 6.560 5.480 ;
        RECT 5.190 5.140 5.550 5.310 ;
        RECT 5.190 4.780 5.840 5.140 ;
        RECT 5.190 4.550 5.460 4.780 ;
        RECT 6.090 4.560 6.340 5.310 ;
        RECT 5.160 4.380 5.490 4.550 ;
        RECT 6.010 4.380 6.340 4.560 ;
        RECT 5.120 3.710 5.530 3.950 ;
        RECT 5.970 3.710 6.380 3.950 ;
        RECT 5.120 3.330 6.380 3.710 ;
        RECT 5.120 3.070 5.530 3.330 ;
        RECT 5.970 3.080 6.380 3.330 ;
        RECT 5.150 2.480 5.490 2.650 ;
        RECT 6.000 2.480 6.360 2.660 ;
        RECT 5.230 1.990 5.410 2.480 ;
        RECT 6.080 1.990 6.270 2.480 ;
  END
END sky130_hilas_TAcoreblock

MACRO sky130_hilas_nFETLarge
  CLASS BLOCK ;
  FOREIGN sky130_hilas_nFETLarge ;
  ORIGIN -0.640 -4.200 ;
  SIZE 4.370 BY 5.830 ;
  PIN GATE
    USE ANALOG ;
    ANTENNAGATEAREA 6.396000 ;
    PORT
      LAYER li1 ;
        RECT 0.830 4.950 1.340 5.210 ;
        RECT 0.830 4.880 1.350 4.950 ;
        RECT 0.840 4.200 1.350 4.880 ;
      LAYER mcon ;
        RECT 1.000 4.740 1.170 4.910 ;
        RECT 1.010 4.270 1.180 4.440 ;
      LAYER met1 ;
        RECT 0.930 4.670 1.250 4.990 ;
        RECT 0.940 4.200 1.260 4.520 ;
      LAYER via ;
        RECT 0.960 4.700 1.220 4.960 ;
        RECT 0.970 4.230 1.230 4.490 ;
      LAYER met2 ;
        RECT 0.640 4.530 1.240 5.020 ;
        RECT 0.640 4.200 1.250 4.530 ;
    END
  END GATE
  PIN SOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 4.231200 ;
    PORT
      LAYER li1 ;
        RECT 1.590 9.750 1.760 9.780 ;
        RECT 2.690 9.750 2.860 9.780 ;
        RECT 1.520 9.710 1.840 9.750 ;
        RECT 2.610 9.710 2.930 9.750 ;
        RECT 3.790 9.740 3.960 9.780 ;
        RECT 1.520 9.520 1.850 9.710 ;
        RECT 2.610 9.520 2.940 9.710 ;
        RECT 3.710 9.700 4.030 9.740 ;
        RECT 1.520 9.490 1.840 9.520 ;
        RECT 2.610 9.490 2.930 9.520 ;
        RECT 3.710 9.510 4.040 9.700 ;
        RECT 1.590 6.970 1.760 9.490 ;
        RECT 2.690 6.970 2.860 9.490 ;
        RECT 3.710 9.480 4.030 9.510 ;
        RECT 3.790 6.970 3.960 9.480 ;
        RECT 1.510 6.930 1.830 6.970 ;
        RECT 2.610 6.930 2.930 6.970 ;
        RECT 3.710 6.930 4.030 6.970 ;
        RECT 1.510 6.740 1.840 6.930 ;
        RECT 2.610 6.740 2.940 6.930 ;
        RECT 3.710 6.740 4.040 6.930 ;
        RECT 1.510 6.710 1.830 6.740 ;
        RECT 2.610 6.710 2.930 6.740 ;
        RECT 3.710 6.710 4.030 6.740 ;
        RECT 1.590 5.600 1.760 6.710 ;
        RECT 2.690 5.600 2.860 6.710 ;
        RECT 3.790 5.600 3.960 6.710 ;
        RECT 1.510 5.560 1.830 5.600 ;
        RECT 2.610 5.560 2.930 5.600 ;
        RECT 3.710 5.560 4.030 5.600 ;
        RECT 1.510 5.370 1.840 5.560 ;
        RECT 2.610 5.370 2.940 5.560 ;
        RECT 3.710 5.370 4.040 5.560 ;
        RECT 1.510 5.340 1.830 5.370 ;
        RECT 2.610 5.340 2.930 5.370 ;
        RECT 3.710 5.340 4.030 5.370 ;
        RECT 1.590 4.600 1.760 5.340 ;
        RECT 2.690 4.600 2.860 5.340 ;
        RECT 3.790 4.600 3.960 5.340 ;
      LAYER mcon ;
        RECT 1.580 9.530 1.750 9.700 ;
        RECT 2.670 9.530 2.840 9.700 ;
        RECT 3.770 9.520 3.940 9.690 ;
        RECT 1.570 6.750 1.740 6.920 ;
        RECT 2.670 6.750 2.840 6.920 ;
        RECT 3.770 6.750 3.940 6.920 ;
        RECT 1.570 5.380 1.740 5.550 ;
        RECT 2.670 5.380 2.840 5.550 ;
        RECT 3.770 5.380 3.940 5.550 ;
      LAYER met1 ;
        RECT 1.510 9.460 1.830 9.780 ;
        RECT 2.600 9.460 2.920 9.780 ;
        RECT 3.700 9.450 4.020 9.770 ;
        RECT 1.500 6.680 1.820 7.000 ;
        RECT 2.600 6.680 2.920 7.000 ;
        RECT 3.700 6.680 4.020 7.000 ;
        RECT 1.500 5.310 1.820 5.630 ;
        RECT 2.600 5.310 2.920 5.630 ;
        RECT 3.700 5.310 4.020 5.630 ;
      LAYER via ;
        RECT 1.540 9.490 1.800 9.750 ;
        RECT 2.630 9.490 2.890 9.750 ;
        RECT 3.730 9.480 3.990 9.740 ;
        RECT 1.530 6.710 1.790 6.970 ;
        RECT 2.630 6.710 2.890 6.970 ;
        RECT 3.730 6.710 3.990 6.970 ;
        RECT 1.530 5.340 1.790 5.600 ;
        RECT 2.630 5.340 2.890 5.600 ;
        RECT 3.730 5.340 3.990 5.600 ;
      LAYER met2 ;
        RECT 0.970 9.790 4.030 9.800 ;
        RECT 0.880 9.460 4.030 9.790 ;
        RECT 0.880 7.010 1.200 9.460 ;
        RECT 3.700 9.450 4.010 9.460 ;
        RECT 0.880 6.680 4.040 7.010 ;
        RECT 0.880 5.640 1.200 6.680 ;
        RECT 0.880 5.320 4.040 5.640 ;
        RECT 1.500 5.310 1.810 5.320 ;
        RECT 2.600 5.310 2.910 5.320 ;
        RECT 3.700 5.310 4.010 5.320 ;
    END
  END SOURCE
  PIN DRAIN
    USE ANALOG ;
    ANTENNADIFFAREA 4.231200 ;
    PORT
      LAYER li1 ;
        RECT 2.140 9.070 2.310 9.780 ;
        RECT 2.070 9.030 2.390 9.070 ;
        RECT 3.240 9.050 3.410 9.780 ;
        RECT 2.070 8.840 2.400 9.030 ;
        RECT 3.160 9.010 3.480 9.050 ;
        RECT 4.340 9.040 4.510 9.780 ;
        RECT 2.070 8.810 2.390 8.840 ;
        RECT 3.160 8.820 3.490 9.010 ;
        RECT 4.270 9.000 4.590 9.040 ;
        RECT 2.140 7.700 2.310 8.810 ;
        RECT 3.160 8.790 3.480 8.820 ;
        RECT 4.270 8.810 4.600 9.000 ;
        RECT 3.240 7.700 3.410 8.790 ;
        RECT 4.270 8.780 4.590 8.810 ;
        RECT 4.340 7.700 4.510 8.780 ;
        RECT 2.070 7.660 2.390 7.700 ;
        RECT 3.160 7.660 3.480 7.700 ;
        RECT 4.260 7.660 4.580 7.700 ;
        RECT 2.070 7.470 2.400 7.660 ;
        RECT 3.160 7.470 3.490 7.660 ;
        RECT 4.260 7.470 4.590 7.660 ;
        RECT 2.070 7.440 2.390 7.470 ;
        RECT 3.160 7.440 3.480 7.470 ;
        RECT 4.260 7.440 4.580 7.470 ;
        RECT 2.140 4.920 2.310 7.440 ;
        RECT 3.240 4.920 3.410 7.440 ;
        RECT 4.340 4.930 4.510 7.440 ;
        RECT 2.070 4.880 2.390 4.920 ;
        RECT 3.160 4.880 3.480 4.920 ;
        RECT 4.260 4.890 4.580 4.930 ;
        RECT 2.070 4.690 2.400 4.880 ;
        RECT 3.160 4.690 3.490 4.880 ;
        RECT 4.260 4.700 4.590 4.890 ;
        RECT 2.070 4.660 2.390 4.690 ;
        RECT 3.160 4.660 3.480 4.690 ;
        RECT 4.260 4.670 4.580 4.700 ;
        RECT 2.140 4.600 2.310 4.660 ;
        RECT 3.240 4.600 3.410 4.660 ;
        RECT 4.340 4.600 4.510 4.670 ;
      LAYER mcon ;
        RECT 2.130 8.850 2.300 9.020 ;
        RECT 3.220 8.830 3.390 9.000 ;
        RECT 4.330 8.820 4.500 8.990 ;
        RECT 2.130 7.480 2.300 7.650 ;
        RECT 3.220 7.480 3.390 7.650 ;
        RECT 4.320 7.480 4.490 7.650 ;
        RECT 2.130 4.700 2.300 4.870 ;
        RECT 3.220 4.700 3.390 4.870 ;
        RECT 4.320 4.710 4.490 4.880 ;
      LAYER met1 ;
        RECT 2.060 8.780 2.380 9.100 ;
        RECT 3.150 8.760 3.470 9.080 ;
        RECT 4.260 8.750 4.580 9.070 ;
        RECT 2.060 7.410 2.380 7.730 ;
        RECT 3.150 7.410 3.470 7.730 ;
        RECT 4.250 7.410 4.570 7.730 ;
        RECT 2.060 4.630 2.380 4.950 ;
        RECT 3.150 4.630 3.470 4.950 ;
        RECT 4.250 4.640 4.570 4.960 ;
      LAYER via ;
        RECT 2.090 8.810 2.350 9.070 ;
        RECT 3.180 8.790 3.440 9.050 ;
        RECT 4.290 8.780 4.550 9.040 ;
        RECT 2.090 7.440 2.350 7.700 ;
        RECT 3.180 7.440 3.440 7.700 ;
        RECT 4.280 7.440 4.540 7.700 ;
        RECT 2.090 4.660 2.350 4.920 ;
        RECT 3.180 4.660 3.440 4.920 ;
        RECT 4.280 4.670 4.540 4.930 ;
      LAYER met2 ;
        RECT 2.060 9.080 2.370 9.110 ;
        RECT 3.150 9.080 3.460 9.090 ;
        RECT 2.060 8.780 5.010 9.080 ;
        RECT 3.150 8.760 3.460 8.780 ;
        RECT 4.260 8.740 5.010 8.780 ;
        RECT 4.630 8.610 5.010 8.740 ;
        RECT 4.660 7.740 5.010 8.610 ;
        RECT 2.060 7.410 5.010 7.740 ;
        RECT 4.660 4.970 5.010 7.410 ;
        RECT 2.070 4.960 5.010 4.970 ;
        RECT 2.060 4.650 5.010 4.960 ;
        RECT 2.060 4.640 4.780 4.650 ;
        RECT 2.060 4.630 2.370 4.640 ;
        RECT 3.150 4.630 3.460 4.640 ;
    END
  END DRAIN
END sky130_hilas_nFETLarge

MACRO sky130_hilas_mcap2m4
  CLASS BLOCK ;
  FOREIGN sky130_hilas_mcap2m4 ;
  ORIGIN 0.360 0.360 ;
  SIZE 0.790 BY 0.750 ;
  OBS
      LAYER met2 ;
        RECT -0.140 -0.160 0.230 0.240 ;
      LAYER via2 ;
        RECT -0.090 -0.100 0.190 0.180 ;
      LAYER met3 ;
        RECT -0.360 -0.360 0.430 0.390 ;
      LAYER via3 ;
        RECT -0.170 -0.210 0.260 0.270 ;
      LAYER met4 ;
        RECT -0.270 -0.300 0.390 0.360 ;
  END
END sky130_hilas_mcap2m4

MACRO sky130_hilas_all
  CLASS BLOCK ;
  FOREIGN sky130_hilas_all ;
  ORIGIN 6.020 4.410 ;
  SIZE 1.770 BY 6.670 ;
  OBS
      LAYER nwell ;
        RECT -5.720 -0.430 -4.250 2.260 ;
        RECT -6.010 -0.670 -4.250 -0.430 ;
        RECT -6.020 -1.500 -4.250 -0.670 ;
        RECT -5.720 -4.410 -4.250 -1.500 ;
      LAYER li1 ;
        RECT -5.400 1.720 -4.900 1.890 ;
        RECT -5.230 0.930 -4.890 1.100 ;
        RECT -5.230 0.360 -4.890 0.530 ;
        RECT -5.690 -1.170 -4.890 -1.000 ;
        RECT -5.230 -2.690 -4.890 -2.520 ;
        RECT -5.230 -3.250 -4.890 -3.080 ;
        RECT -5.230 -4.040 -4.890 -3.870 ;
      LAYER mcon ;
        RECT -5.400 -1.170 -5.220 -1.000 ;
      LAYER met1 ;
        RECT -5.360 1.950 -5.020 2.000 ;
        RECT -5.460 1.700 -4.900 1.950 ;
        RECT -5.360 1.670 -5.020 1.700 ;
        RECT -5.200 -0.960 -4.950 -0.950 ;
        RECT -5.690 -1.170 -5.540 -1.000 ;
        RECT -5.460 -1.210 -4.920 -0.960 ;
      LAYER via ;
        RECT -5.320 1.700 -5.060 1.960 ;
        RECT -5.200 -1.210 -4.950 -0.950 ;
      LAYER met2 ;
        RECT -5.360 1.960 -5.020 2.000 ;
        RECT -5.720 1.700 -4.530 1.960 ;
        RECT -5.360 1.670 -5.020 1.700 ;
        RECT -5.220 -0.940 -4.920 -0.930 ;
        RECT -5.220 -0.950 -4.910 -0.940 ;
        RECT -5.420 -1.220 -4.890 -0.950 ;
        RECT -5.220 -1.240 -4.920 -1.220 ;
  END
END sky130_hilas_all

MACRO sky130_hilas_nOverlapCap01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_nOverlapCap01 ;
  ORIGIN 0.620 0.430 ;
  SIZE 1.290 BY 1.290 ;
  OBS
      LAYER li1 ;
        RECT -0.060 -0.220 0.110 0.670 ;
      LAYER mcon ;
        RECT -0.060 0.470 0.110 0.640 ;
      LAYER met1 ;
        RECT -0.090 -0.430 0.140 0.860 ;
  END
END sky130_hilas_nOverlapCap01

MACRO sky130_hilas_pFETmed
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pFETmed ;
  ORIGIN -1.470 0.220 ;
  SIZE 1.190 BY 2.870 ;
  OBS
      LAYER nwell ;
        RECT 1.470 -0.220 2.660 2.650 ;
      LAYER li1 ;
        RECT 1.710 -0.070 1.880 2.420 ;
        RECT 2.260 -0.080 2.430 2.420 ;
  END
END sky130_hilas_pFETmed

MACRO sky130_hilas_poly2li
  CLASS BLOCK ;
  FOREIGN sky130_hilas_poly2li ;
  ORIGIN 0.090 0.140 ;
  SIZE 0.270 BY 0.330 ;
  OBS
      LAYER li1 ;
        RECT -0.040 -0.140 0.130 0.190 ;
  END
END sky130_hilas_poly2li

MACRO sky130_hilas_nFETmed
  CLASS BLOCK ;
  FOREIGN sky130_hilas_nFETmed ;
  ORIGIN 0.120 0.440 ;
  SIZE 0.820 BY 2.720 ;
  OBS
      LAYER li1 ;
        RECT -0.070 -0.260 0.100 2.140 ;
        RECT 0.480 -0.260 0.650 2.140 ;
  END
END sky130_hilas_nFETmed

MACRO sky130_hilas_DAC6TransistorStack01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_DAC6TransistorStack01 ;
  ORIGIN -0.280 1.740 ;
  SIZE 1.720 BY 5.650 ;
  OBS
      LAYER nwell ;
        RECT 0.280 -1.740 1.890 3.910 ;
      LAYER li1 ;
        RECT 0.660 2.360 0.830 2.690 ;
        RECT 1.340 2.360 1.510 2.690 ;
        RECT 0.660 1.400 0.830 1.730 ;
        RECT 1.340 1.400 1.510 1.730 ;
        RECT 0.660 0.440 0.830 0.770 ;
        RECT 1.340 0.440 1.510 0.770 ;
        RECT 0.660 -0.520 0.830 -0.190 ;
        RECT 1.340 -0.520 1.510 -0.190 ;
  END
END sky130_hilas_DAC6TransistorStack01

MACRO sky130_hilas_DoubleTGate01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_DoubleTGate01 ;
  ORIGIN -10.720 -0.050 ;
  SIZE 5.420 BY 6.050 ;
  OBS
      LAYER nwell ;
        RECT 10.720 0.050 13.920 6.100 ;
      LAYER li1 ;
        RECT 11.120 4.840 11.290 5.770 ;
        RECT 14.810 5.700 15.050 5.730 ;
        RECT 11.820 5.530 12.780 5.700 ;
        RECT 13.230 5.530 14.570 5.700 ;
        RECT 14.810 5.530 15.380 5.700 ;
        RECT 12.100 5.520 12.270 5.530 ;
        RECT 14.810 5.490 15.050 5.530 ;
        RECT 12.260 5.080 12.590 5.260 ;
        RECT 15.760 5.180 15.930 5.220 ;
        RECT 15.400 5.080 15.590 5.100 ;
        RECT 11.820 4.910 14.570 5.080 ;
        RECT 15.030 4.910 15.590 5.080 ;
        RECT 15.400 4.870 15.590 4.910 ;
        RECT 15.760 5.010 15.990 5.180 ;
        RECT 15.760 4.660 15.930 5.010 ;
        RECT 11.120 3.310 11.290 4.240 ;
        RECT 15.400 4.170 15.590 4.210 ;
        RECT 11.820 4.000 14.570 4.170 ;
        RECT 15.030 4.000 15.590 4.170 ;
        RECT 12.260 3.820 12.590 4.000 ;
        RECT 15.400 3.980 15.590 4.000 ;
        RECT 15.760 4.070 15.930 4.420 ;
        RECT 15.760 3.900 15.990 4.070 ;
        RECT 15.760 3.860 15.930 3.900 ;
        RECT 12.100 3.550 12.270 3.560 ;
        RECT 14.810 3.550 15.050 3.590 ;
        RECT 11.820 3.380 12.780 3.550 ;
        RECT 13.230 3.380 14.570 3.550 ;
        RECT 14.810 3.380 15.380 3.550 ;
        RECT 14.810 3.350 15.050 3.380 ;
        RECT 11.120 1.910 11.290 2.840 ;
        RECT 14.810 2.770 15.050 2.800 ;
        RECT 11.820 2.600 12.780 2.770 ;
        RECT 13.230 2.600 14.570 2.770 ;
        RECT 14.810 2.600 15.380 2.770 ;
        RECT 12.100 2.590 12.270 2.600 ;
        RECT 14.810 2.560 15.050 2.600 ;
        RECT 12.260 2.150 12.590 2.330 ;
        RECT 15.760 2.250 15.930 2.290 ;
        RECT 15.400 2.150 15.590 2.170 ;
        RECT 11.820 1.980 14.570 2.150 ;
        RECT 15.030 1.980 15.590 2.150 ;
        RECT 15.400 1.940 15.590 1.980 ;
        RECT 15.760 2.080 15.990 2.250 ;
        RECT 15.760 1.730 15.930 2.080 ;
        RECT 11.120 0.380 11.290 1.310 ;
        RECT 15.400 1.240 15.590 1.280 ;
        RECT 11.820 1.070 14.570 1.240 ;
        RECT 15.030 1.070 15.590 1.240 ;
        RECT 12.260 0.890 12.590 1.070 ;
        RECT 15.400 1.050 15.590 1.070 ;
        RECT 15.760 1.140 15.930 1.490 ;
        RECT 15.760 0.970 15.990 1.140 ;
        RECT 15.760 0.930 15.930 0.970 ;
        RECT 12.100 0.620 12.270 0.630 ;
        RECT 14.810 0.620 15.050 0.660 ;
        RECT 11.820 0.450 12.780 0.620 ;
        RECT 13.230 0.450 14.570 0.620 ;
        RECT 14.810 0.450 15.380 0.620 ;
        RECT 14.810 0.420 15.050 0.450 ;
      LAYER mcon ;
        RECT 14.100 5.530 14.270 5.700 ;
        RECT 14.850 5.530 15.020 5.700 ;
        RECT 11.120 5.200 11.290 5.370 ;
        RECT 15.410 4.900 15.580 5.070 ;
        RECT 15.820 5.010 15.990 5.180 ;
        RECT 15.410 4.010 15.580 4.180 ;
        RECT 11.120 3.710 11.290 3.880 ;
        RECT 15.820 3.900 15.990 4.070 ;
        RECT 12.100 3.390 12.270 3.560 ;
        RECT 14.100 3.380 14.270 3.550 ;
        RECT 14.850 3.380 15.020 3.550 ;
        RECT 14.100 2.600 14.270 2.770 ;
        RECT 14.850 2.600 15.020 2.770 ;
        RECT 11.120 2.270 11.290 2.440 ;
        RECT 15.410 1.970 15.580 2.140 ;
        RECT 15.820 2.080 15.990 2.250 ;
        RECT 15.410 1.080 15.580 1.250 ;
        RECT 11.120 0.780 11.290 0.950 ;
        RECT 15.820 0.970 15.990 1.140 ;
        RECT 12.100 0.460 12.270 0.630 ;
        RECT 14.100 0.450 14.270 0.620 ;
        RECT 14.850 0.450 15.020 0.620 ;
      LAYER met1 ;
        RECT 11.080 0.050 11.330 6.100 ;
        RECT 12.230 5.720 12.570 5.770 ;
        RECT 12.010 5.700 12.570 5.720 ;
        RECT 12.010 5.530 12.690 5.700 ;
        RECT 12.010 5.490 12.570 5.530 ;
        RECT 12.230 5.450 12.570 5.490 ;
        RECT 12.230 3.590 12.570 3.630 ;
        RECT 12.010 3.550 12.570 3.590 ;
        RECT 12.010 3.380 12.690 3.550 ;
        RECT 12.010 3.360 12.570 3.380 ;
        RECT 12.230 3.310 12.570 3.360 ;
        RECT 12.230 2.790 12.570 2.840 ;
        RECT 12.010 2.770 12.570 2.790 ;
        RECT 12.010 2.600 12.690 2.770 ;
        RECT 12.010 2.560 12.570 2.600 ;
        RECT 12.230 2.520 12.570 2.560 ;
        RECT 12.230 0.660 12.570 0.700 ;
        RECT 12.010 0.620 12.570 0.660 ;
        RECT 12.010 0.450 12.690 0.620 ;
        RECT 12.010 0.430 12.570 0.450 ;
        RECT 12.230 0.380 12.570 0.430 ;
        RECT 14.070 0.050 14.300 6.100 ;
        RECT 14.660 5.740 15.030 5.760 ;
        RECT 14.660 5.480 15.080 5.740 ;
        RECT 14.660 5.470 15.030 5.480 ;
        RECT 15.420 5.130 15.610 6.100 ;
        RECT 15.380 4.840 15.610 5.130 ;
        RECT 15.760 4.980 16.140 5.220 ;
        RECT 15.420 4.240 15.610 4.840 ;
        RECT 15.380 3.950 15.610 4.240 ;
        RECT 14.660 3.600 15.030 3.610 ;
        RECT 14.660 3.340 15.080 3.600 ;
        RECT 14.660 3.320 15.030 3.340 ;
        RECT 14.660 2.810 15.030 2.830 ;
        RECT 14.660 2.550 15.080 2.810 ;
        RECT 14.660 2.540 15.030 2.550 ;
        RECT 15.420 2.200 15.610 3.950 ;
        RECT 15.760 3.860 16.140 4.100 ;
        RECT 15.380 1.910 15.610 2.200 ;
        RECT 15.760 2.050 16.140 2.290 ;
        RECT 15.420 1.310 15.610 1.910 ;
        RECT 15.380 1.020 15.610 1.310 ;
        RECT 14.660 0.670 15.030 0.680 ;
        RECT 14.660 0.410 15.080 0.670 ;
        RECT 14.660 0.390 15.030 0.410 ;
        RECT 15.420 0.050 15.610 1.020 ;
        RECT 15.760 0.930 16.140 1.170 ;
      LAYER via ;
        RECT 12.280 5.480 12.540 5.740 ;
        RECT 12.280 3.340 12.540 3.600 ;
        RECT 12.280 2.550 12.540 2.810 ;
        RECT 12.280 0.410 12.540 0.670 ;
        RECT 14.690 5.480 14.950 5.740 ;
        RECT 14.690 3.340 14.950 3.600 ;
        RECT 14.690 2.550 14.950 2.810 ;
        RECT 14.690 0.410 14.950 0.670 ;
      LAYER met2 ;
        RECT 12.250 5.720 12.570 5.740 ;
        RECT 14.660 5.720 14.980 5.770 ;
        RECT 11.070 5.590 11.800 5.600 ;
        RECT 12.250 5.590 14.980 5.720 ;
        RECT 11.070 5.530 14.980 5.590 ;
        RECT 11.070 5.480 12.570 5.530 ;
        RECT 11.070 5.430 12.490 5.480 ;
        RECT 14.660 5.450 14.980 5.530 ;
        RECT 11.070 5.420 11.800 5.430 ;
        RECT 11.070 3.720 11.740 3.740 ;
        RECT 11.070 3.600 12.460 3.720 ;
        RECT 11.070 3.560 12.570 3.600 ;
        RECT 12.250 3.550 12.570 3.560 ;
        RECT 14.660 3.550 14.980 3.630 ;
        RECT 12.250 3.360 14.980 3.550 ;
        RECT 12.250 3.340 12.570 3.360 ;
        RECT 14.660 3.310 14.980 3.360 ;
        RECT 12.250 2.790 12.570 2.810 ;
        RECT 14.660 2.790 14.980 2.840 ;
        RECT 12.250 2.600 14.980 2.790 ;
        RECT 11.070 2.570 11.770 2.580 ;
        RECT 12.250 2.570 12.570 2.600 ;
        RECT 11.070 2.550 12.570 2.570 ;
        RECT 11.070 2.410 12.500 2.550 ;
        RECT 14.660 2.520 14.980 2.600 ;
        RECT 11.070 0.670 12.530 0.740 ;
        RECT 11.070 0.620 12.570 0.670 ;
        RECT 14.660 0.620 14.980 0.700 ;
        RECT 11.070 0.570 14.980 0.620 ;
        RECT 12.250 0.430 14.980 0.570 ;
        RECT 12.250 0.410 12.570 0.430 ;
        RECT 14.660 0.380 14.980 0.430 ;
  END
END sky130_hilas_DoubleTGate01

MACRO sky130_hilas_DAC6TransistorStack01c
  CLASS BLOCK ;
  FOREIGN sky130_hilas_DAC6TransistorStack01c ;
  ORIGIN -0.280 1.740 ;
  SIZE 1.870 BY 5.650 ;
  OBS
      LAYER nwell ;
        RECT 0.280 -1.740 1.890 3.910 ;
      LAYER li1 ;
        RECT 0.660 2.360 0.830 2.690 ;
        RECT 1.340 2.360 1.510 2.690 ;
        RECT 0.660 1.400 0.830 1.730 ;
        RECT 1.340 1.400 1.510 1.730 ;
        RECT 0.660 -0.520 0.830 -0.190 ;
        RECT 1.340 -0.520 1.510 -0.190 ;
        RECT 1.850 -0.460 2.060 -0.030 ;
        RECT 1.870 -0.480 2.040 -0.460 ;
      LAYER met1 ;
        RECT 1.850 -0.250 2.070 -0.030 ;
        RECT 1.840 -0.540 2.070 -0.250 ;
  END
END sky130_hilas_DAC6TransistorStack01c

MACRO sky130_hilas_TgateSingle01Part1
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TgateSingle01Part1 ;
  ORIGIN -2.570 1.810 ;
  SIZE 1.880 BY 1.520 ;
  OBS
      LAYER li1 ;
        RECT 3.940 -0.700 4.130 -0.680 ;
        RECT 2.570 -0.880 3.210 -0.700 ;
        RECT 3.590 -0.710 4.130 -0.700 ;
        RECT 3.590 -0.870 4.370 -0.710 ;
        RECT 3.940 -0.910 4.370 -0.870 ;
        RECT 2.970 -1.410 3.140 -1.250 ;
        RECT 3.480 -1.330 3.670 -1.300 ;
        RECT 2.910 -1.450 3.230 -1.410 ;
        RECT 2.910 -1.640 3.240 -1.450 ;
        RECT 3.480 -1.500 3.920 -1.330 ;
        RECT 3.480 -1.530 3.670 -1.500 ;
        RECT 4.200 -1.590 4.370 -0.910 ;
        RECT 2.910 -1.670 3.230 -1.640 ;
      LAYER mcon ;
        RECT 3.950 -0.880 4.120 -0.710 ;
        RECT 2.970 -1.630 3.140 -1.460 ;
        RECT 3.490 -1.500 3.660 -1.330 ;
      LAYER met1 ;
        RECT 3.290 -0.530 3.550 -0.460 ;
        RECT 3.290 -0.780 3.650 -0.530 ;
        RECT 3.940 -0.650 4.130 -0.290 ;
        RECT 3.460 -1.270 3.650 -0.780 ;
        RECT 3.920 -0.940 4.150 -0.650 ;
        RECT 2.900 -1.700 3.220 -1.380 ;
        RECT 3.460 -1.560 3.690 -1.270 ;
        RECT 3.940 -1.810 4.130 -0.940 ;
      LAYER via ;
        RECT 3.290 -0.750 3.550 -0.490 ;
        RECT 2.930 -1.670 3.190 -1.410 ;
      LAYER met2 ;
        RECT 3.260 -0.520 3.580 -0.490 ;
        RECT 2.570 -0.720 4.450 -0.520 ;
        RECT 3.260 -0.750 3.580 -0.720 ;
        RECT 2.900 -1.500 3.210 -1.370 ;
        RECT 2.570 -1.700 3.210 -1.500 ;
  END
END sky130_hilas_TgateSingle01Part1

MACRO sky130_hilas_pFETLarge
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pFETLarge ;
  ORIGIN -0.640 -4.190 ;
  SIZE 4.640 BY 5.990 ;
  PIN GATE
    ANTENNAGATEAREA 6.526000 ;
    PORT
      LAYER li1 ;
        RECT 0.830 4.950 1.340 5.210 ;
        RECT 0.830 4.880 1.350 4.950 ;
        RECT 0.840 4.200 1.350 4.880 ;
      LAYER mcon ;
        RECT 1.000 4.740 1.170 4.910 ;
        RECT 1.010 4.270 1.180 4.440 ;
      LAYER met1 ;
        RECT 0.930 4.670 1.250 4.990 ;
        RECT 0.940 4.200 1.260 4.520 ;
      LAYER via ;
        RECT 0.960 4.700 1.220 4.960 ;
        RECT 0.970 4.230 1.230 4.490 ;
      LAYER met2 ;
        RECT 0.640 4.530 1.240 5.020 ;
        RECT 0.640 4.200 1.250 4.530 ;
    END
  END GATE
  PIN SOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 4.367400 ;
    PORT
      LAYER li1 ;
        RECT 1.600 9.750 1.770 9.840 ;
        RECT 2.700 9.750 2.870 9.840 ;
        RECT 1.520 9.710 1.840 9.750 ;
        RECT 2.610 9.710 2.930 9.750 ;
        RECT 3.800 9.740 3.970 9.840 ;
        RECT 1.520 9.520 1.850 9.710 ;
        RECT 2.610 9.520 2.940 9.710 ;
        RECT 3.710 9.700 4.030 9.740 ;
        RECT 1.520 9.490 1.840 9.520 ;
        RECT 2.610 9.490 2.930 9.520 ;
        RECT 3.710 9.510 4.040 9.700 ;
        RECT 1.600 6.970 1.770 9.490 ;
        RECT 2.700 6.970 2.870 9.490 ;
        RECT 3.710 9.480 4.030 9.510 ;
        RECT 3.800 6.970 3.970 9.480 ;
        RECT 1.510 6.930 1.830 6.970 ;
        RECT 2.610 6.930 2.930 6.970 ;
        RECT 3.710 6.930 4.030 6.970 ;
        RECT 1.510 6.740 1.840 6.930 ;
        RECT 2.610 6.740 2.940 6.930 ;
        RECT 3.710 6.740 4.040 6.930 ;
        RECT 1.510 6.710 1.830 6.740 ;
        RECT 2.610 6.710 2.930 6.740 ;
        RECT 3.710 6.710 4.030 6.740 ;
        RECT 1.600 5.600 1.770 6.710 ;
        RECT 2.700 5.600 2.870 6.710 ;
        RECT 3.800 5.600 3.970 6.710 ;
        RECT 1.510 5.560 1.830 5.600 ;
        RECT 2.610 5.560 2.930 5.600 ;
        RECT 3.710 5.560 4.030 5.600 ;
        RECT 1.510 5.370 1.840 5.560 ;
        RECT 2.610 5.370 2.940 5.560 ;
        RECT 3.710 5.370 4.040 5.560 ;
        RECT 1.510 5.340 1.830 5.370 ;
        RECT 2.610 5.340 2.930 5.370 ;
        RECT 3.710 5.340 4.030 5.370 ;
        RECT 1.600 4.520 1.770 5.340 ;
        RECT 2.700 4.510 2.870 5.340 ;
        RECT 3.800 4.510 3.970 5.340 ;
      LAYER mcon ;
        RECT 1.580 9.530 1.750 9.700 ;
        RECT 2.670 9.530 2.840 9.700 ;
        RECT 3.770 9.520 3.940 9.690 ;
        RECT 1.570 6.750 1.740 6.920 ;
        RECT 2.670 6.750 2.840 6.920 ;
        RECT 3.770 6.750 3.940 6.920 ;
        RECT 1.570 5.380 1.740 5.550 ;
        RECT 2.670 5.380 2.840 5.550 ;
        RECT 3.770 5.380 3.940 5.550 ;
      LAYER met1 ;
        RECT 1.510 9.460 1.830 9.780 ;
        RECT 2.600 9.460 2.920 9.780 ;
        RECT 3.700 9.450 4.020 9.770 ;
        RECT 1.500 6.680 1.820 7.000 ;
        RECT 2.600 6.680 2.920 7.000 ;
        RECT 3.700 6.680 4.020 7.000 ;
        RECT 1.500 5.310 1.820 5.630 ;
        RECT 2.600 5.310 2.920 5.630 ;
        RECT 3.700 5.310 4.020 5.630 ;
      LAYER via ;
        RECT 1.540 9.490 1.800 9.750 ;
        RECT 2.630 9.490 2.890 9.750 ;
        RECT 3.730 9.480 3.990 9.740 ;
        RECT 1.530 6.710 1.790 6.970 ;
        RECT 2.630 6.710 2.890 6.970 ;
        RECT 3.730 6.710 3.990 6.970 ;
        RECT 1.530 5.340 1.790 5.600 ;
        RECT 2.630 5.340 2.890 5.600 ;
        RECT 3.730 5.340 3.990 5.600 ;
      LAYER met2 ;
        RECT 0.970 9.790 4.030 9.800 ;
        RECT 0.880 9.460 4.030 9.790 ;
        RECT 0.880 7.010 1.200 9.460 ;
        RECT 3.700 9.450 4.010 9.460 ;
        RECT 0.880 6.680 4.040 7.010 ;
        RECT 0.880 5.640 1.200 6.680 ;
        RECT 0.880 5.320 4.040 5.640 ;
        RECT 1.500 5.310 1.810 5.320 ;
        RECT 2.600 5.310 2.910 5.320 ;
        RECT 3.700 5.310 4.010 5.320 ;
    END
  END SOURCE
  PIN DRAIN
    USE ANALOG ;
    ANTENNADIFFAREA 4.317200 ;
    PORT
      LAYER li1 ;
        RECT 2.150 9.070 2.320 9.840 ;
        RECT 2.070 9.030 2.390 9.070 ;
        RECT 3.250 9.050 3.420 9.840 ;
        RECT 2.070 8.840 2.400 9.030 ;
        RECT 3.160 9.010 3.480 9.050 ;
        RECT 4.350 9.040 4.520 9.840 ;
        RECT 2.070 8.810 2.390 8.840 ;
        RECT 3.160 8.820 3.490 9.010 ;
        RECT 4.270 9.000 4.590 9.040 ;
        RECT 2.150 7.700 2.320 8.810 ;
        RECT 3.160 8.790 3.480 8.820 ;
        RECT 4.270 8.810 4.600 9.000 ;
        RECT 3.250 7.700 3.420 8.790 ;
        RECT 4.270 8.780 4.590 8.810 ;
        RECT 4.350 7.700 4.520 8.780 ;
        RECT 2.070 7.660 2.390 7.700 ;
        RECT 3.160 7.660 3.480 7.700 ;
        RECT 4.260 7.660 4.580 7.700 ;
        RECT 2.070 7.470 2.400 7.660 ;
        RECT 3.160 7.470 3.490 7.660 ;
        RECT 4.260 7.470 4.590 7.660 ;
        RECT 2.070 7.440 2.390 7.470 ;
        RECT 3.160 7.440 3.480 7.470 ;
        RECT 4.260 7.440 4.580 7.470 ;
        RECT 2.150 4.920 2.320 7.440 ;
        RECT 3.250 4.920 3.420 7.440 ;
        RECT 4.350 4.930 4.520 7.440 ;
        RECT 2.070 4.880 2.390 4.920 ;
        RECT 3.160 4.880 3.480 4.920 ;
        RECT 4.260 4.890 4.580 4.930 ;
        RECT 2.070 4.690 2.400 4.880 ;
        RECT 3.160 4.690 3.490 4.880 ;
        RECT 4.260 4.700 4.590 4.890 ;
        RECT 2.070 4.660 2.390 4.690 ;
        RECT 3.160 4.660 3.480 4.690 ;
        RECT 4.260 4.670 4.580 4.700 ;
        RECT 2.150 4.510 2.320 4.660 ;
        RECT 3.250 4.510 3.420 4.660 ;
        RECT 4.350 4.510 4.520 4.670 ;
      LAYER mcon ;
        RECT 2.130 8.850 2.300 9.020 ;
        RECT 3.220 8.830 3.390 9.000 ;
        RECT 4.330 8.820 4.500 8.990 ;
        RECT 2.130 7.480 2.300 7.650 ;
        RECT 3.220 7.480 3.390 7.650 ;
        RECT 4.320 7.480 4.490 7.650 ;
        RECT 2.130 4.700 2.300 4.870 ;
        RECT 3.220 4.700 3.390 4.870 ;
        RECT 4.320 4.710 4.490 4.880 ;
      LAYER met1 ;
        RECT 2.060 8.780 2.380 9.100 ;
        RECT 3.150 8.760 3.470 9.080 ;
        RECT 4.260 8.750 4.580 9.070 ;
        RECT 2.060 7.410 2.380 7.730 ;
        RECT 3.150 7.410 3.470 7.730 ;
        RECT 4.250 7.410 4.570 7.730 ;
        RECT 2.060 4.630 2.380 4.950 ;
        RECT 3.150 4.630 3.470 4.950 ;
        RECT 4.250 4.640 4.570 4.960 ;
      LAYER via ;
        RECT 2.090 8.810 2.350 9.070 ;
        RECT 3.180 8.790 3.440 9.050 ;
        RECT 4.290 8.780 4.550 9.040 ;
        RECT 2.090 7.440 2.350 7.700 ;
        RECT 3.180 7.440 3.440 7.700 ;
        RECT 4.280 7.440 4.540 7.700 ;
        RECT 2.090 4.660 2.350 4.920 ;
        RECT 3.180 4.660 3.440 4.920 ;
        RECT 4.280 4.670 4.540 4.930 ;
      LAYER met2 ;
        RECT 2.060 9.080 2.370 9.110 ;
        RECT 3.150 9.080 3.460 9.090 ;
        RECT 2.060 8.780 5.010 9.080 ;
        RECT 3.150 8.760 3.460 8.780 ;
        RECT 4.260 8.740 5.010 8.780 ;
        RECT 4.630 8.610 5.010 8.740 ;
        RECT 4.660 7.740 5.010 8.610 ;
        RECT 2.060 7.410 5.010 7.740 ;
        RECT 4.660 4.970 5.010 7.410 ;
        RECT 2.070 4.960 5.010 4.970 ;
        RECT 2.060 4.650 5.010 4.960 ;
        RECT 2.060 4.640 4.780 4.650 ;
        RECT 2.060 4.630 2.370 4.640 ;
        RECT 3.150 4.630 3.460 4.640 ;
    END
  END DRAIN
  PIN WELL
    USE ANALOG ;
    ANTENNADIFFAREA 0.213200 ;
    PORT
      LAYER nwell ;
        RECT 1.360 4.370 5.280 10.070 ;
      LAYER li1 ;
        RECT 4.890 9.110 5.060 9.870 ;
      LAYER mcon ;
        RECT 4.890 9.700 5.060 9.870 ;
        RECT 4.890 9.360 5.060 9.530 ;
      LAYER met1 ;
        RECT 4.780 9.980 5.040 10.180 ;
        RECT 4.780 9.170 5.090 9.980 ;
        RECT 4.780 4.190 5.040 9.170 ;
    END
  END WELL
END sky130_hilas_pFETLarge

MACRO sky130_hilas_FGBias2x1cell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_FGBias2x1cell ;
  ORIGIN 3.960 3.820 ;
  SIZE 11.530 BY 6.050 ;
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 2.516100 ;
    PORT
      LAYER nwell ;
        RECT -3.950 1.480 -2.220 2.230 ;
        RECT -3.950 -2.090 -2.210 1.480 ;
        RECT -3.950 -3.810 -2.220 -2.090 ;
      LAYER li1 ;
        RECT -3.520 0.090 -2.970 0.520 ;
        RECT -3.520 -1.640 -2.970 -1.210 ;
      LAYER mcon ;
        RECT -3.520 0.170 -3.250 0.440 ;
        RECT -3.520 -1.560 -3.250 -1.290 ;
      LAYER met1 ;
        RECT -3.610 -3.820 -3.190 2.230 ;
    END
  END VTUN
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT -0.920 -0.740 -0.730 -0.340 ;
        RECT -1.110 -0.750 -0.730 -0.740 ;
        RECT -1.110 -0.930 2.630 -0.750 ;
        RECT -1.110 -0.970 -0.730 -0.930 ;
        RECT -0.920 -1.350 -0.730 -0.970 ;
      LAYER mcon ;
        RECT -1.100 -0.940 -0.930 -0.770 ;
      LAYER met1 ;
        RECT -1.130 -3.820 -0.900 2.230 ;
    END
  END VGND
  PIN GATE_CONTROL
    USE ANALOG ;
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT -0.190 -0.160 2.530 1.490 ;
        RECT -0.190 -0.200 2.520 -0.160 ;
        RECT -0.190 -1.530 2.520 -1.490 ;
        RECT -0.190 -3.180 2.530 -1.530 ;
      LAYER li1 ;
        RECT 0.110 0.280 0.340 0.970 ;
        RECT 0.110 -2.660 0.340 -1.930 ;
      LAYER mcon ;
        RECT 0.140 0.770 0.310 0.940 ;
        RECT 0.140 0.320 0.310 0.490 ;
        RECT 0.140 -2.180 0.310 -2.010 ;
        RECT 0.140 -2.630 0.310 -2.460 ;
      LAYER met1 ;
        RECT 0.090 1.020 0.320 2.230 ;
        RECT 0.090 0.230 0.350 1.020 ;
        RECT 0.090 -1.920 0.320 0.230 ;
        RECT 0.090 -2.710 0.350 -1.920 ;
        RECT 0.090 -3.820 0.320 -2.710 ;
    END
  END GATE_CONTROL
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.105400 ;
    PORT
      LAYER li1 ;
        RECT 5.160 1.650 5.690 1.820 ;
      LAYER met1 ;
        RECT 5.090 1.550 5.390 1.930 ;
      LAYER via ;
        RECT 5.110 1.610 5.370 1.880 ;
      LAYER met2 ;
        RECT 5.090 1.750 5.390 1.930 ;
        RECT 4.840 1.730 5.390 1.750 ;
        RECT -3.960 1.550 7.570 1.730 ;
    END
  END DRAIN1
  PIN DRAIN4
    USE ANALOG ;
    ANTENNADIFFAREA 0.105400 ;
    PORT
      LAYER li1 ;
        RECT 5.160 -3.410 5.690 -3.240 ;
      LAYER met1 ;
        RECT 5.090 -3.520 5.390 -3.140 ;
      LAYER via ;
        RECT 5.110 -3.470 5.370 -3.200 ;
      LAYER met2 ;
        RECT 5.100 -3.140 5.260 -3.130 ;
        RECT 5.010 -3.150 7.570 -3.140 ;
        RECT -3.960 -3.300 7.570 -3.150 ;
        RECT 5.010 -3.320 7.570 -3.300 ;
        RECT 5.090 -3.520 5.390 -3.320 ;
    END
  END DRAIN4
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 4.260 -3.810 7.570 2.230 ;
      LAYER li1 ;
        RECT 6.970 1.550 7.170 1.900 ;
        RECT 6.970 1.520 7.180 1.550 ;
        RECT 6.240 -0.340 6.410 1.270 ;
        RECT 6.960 0.940 7.180 1.520 ;
        RECT 6.970 0.930 7.180 0.940 ;
        RECT 6.240 -0.530 6.420 -0.340 ;
        RECT 6.240 -1.250 6.420 -1.060 ;
        RECT 6.240 -2.860 6.410 -1.250 ;
        RECT 6.970 -2.530 7.180 -2.520 ;
        RECT 6.960 -3.110 7.180 -2.530 ;
        RECT 6.970 -3.140 7.180 -3.110 ;
        RECT 6.970 -3.490 7.170 -3.140 ;
      LAYER mcon ;
        RECT 6.980 1.350 7.150 1.520 ;
        RECT 6.980 -3.110 7.150 -2.940 ;
      LAYER met1 ;
        RECT 7.050 1.580 7.330 2.230 ;
        RECT 6.940 0.980 7.330 1.580 ;
        RECT 6.210 -0.340 6.450 -0.210 ;
        RECT 6.210 -0.660 6.470 -0.340 ;
        RECT 7.050 -0.620 7.330 0.980 ;
        RECT 7.050 -0.940 7.410 -0.620 ;
        RECT 6.210 -1.260 6.470 -0.940 ;
        RECT 6.210 -1.380 6.450 -1.260 ;
        RECT 7.050 -2.570 7.330 -0.940 ;
        RECT 6.940 -3.170 7.330 -2.570 ;
        RECT 7.050 -3.820 7.330 -3.170 ;
      LAYER via ;
        RECT 6.210 -0.630 6.470 -0.370 ;
        RECT 7.150 -0.910 7.410 -0.650 ;
        RECT 6.210 -1.230 6.470 -0.970 ;
      LAYER met2 ;
        RECT 6.180 -0.630 6.500 -0.370 ;
        RECT 6.220 -0.650 7.400 -0.630 ;
        RECT 6.220 -0.910 7.440 -0.650 ;
        RECT 6.220 -0.970 7.400 -0.910 ;
        RECT 6.180 -0.980 7.400 -0.970 ;
        RECT 6.180 -1.230 6.500 -0.980 ;
    END
  END VINJ
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER li1 ;
        RECT 5.410 0.740 5.580 1.260 ;
        RECT 5.250 0.480 5.580 0.740 ;
        RECT 5.410 -0.430 5.580 0.480 ;
      LAYER mcon ;
        RECT 5.310 0.520 5.480 0.690 ;
      LAYER met1 ;
        RECT 5.240 0.450 5.560 0.770 ;
      LAYER via ;
        RECT 5.270 0.480 5.530 0.740 ;
      LAYER met2 ;
        RECT 5.240 0.710 5.550 0.780 ;
        RECT 5.240 0.490 7.570 0.710 ;
        RECT 5.240 0.450 5.550 0.490 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER li1 ;
        RECT 5.410 -2.020 5.580 -1.160 ;
        RECT 5.250 -2.280 5.580 -2.020 ;
        RECT 5.410 -2.850 5.580 -2.280 ;
      LAYER mcon ;
        RECT 5.310 -2.240 5.480 -2.070 ;
      LAYER met1 ;
        RECT 5.240 -2.310 5.560 -1.990 ;
      LAYER via ;
        RECT 5.270 -2.280 5.530 -2.020 ;
      LAYER met2 ;
        RECT 5.240 -2.050 5.550 -1.980 ;
        RECT 5.240 -2.260 7.570 -2.050 ;
        RECT 5.240 -2.310 5.550 -2.260 ;
    END
  END OUTPUT2
  OBS
      LAYER li1 ;
        RECT 3.290 1.070 3.640 1.240 ;
        RECT 4.660 1.070 4.990 1.240 ;
        RECT 6.610 0.760 6.800 0.770 ;
        RECT 6.610 0.470 6.810 0.760 ;
        RECT 3.290 0.280 3.640 0.450 ;
        RECT 4.660 0.280 4.990 0.450 ;
        RECT 6.600 0.140 6.840 0.470 ;
        RECT 3.300 -0.510 3.640 -0.340 ;
        RECT 4.660 -0.510 4.990 -0.340 ;
        RECT 4.740 -1.080 4.910 -0.510 ;
        RECT 3.300 -1.250 3.640 -1.080 ;
        RECT 4.660 -1.250 4.990 -1.080 ;
        RECT 3.290 -2.040 3.640 -1.870 ;
        RECT 4.660 -2.040 4.990 -1.870 ;
        RECT 6.600 -2.060 6.840 -1.730 ;
        RECT 6.610 -2.350 6.810 -2.060 ;
        RECT 6.610 -2.360 6.800 -2.350 ;
        RECT 3.290 -2.830 3.640 -2.660 ;
        RECT 4.660 -2.830 4.990 -2.660 ;
      LAYER mcon ;
        RECT 6.620 0.510 6.800 0.700 ;
        RECT 6.620 -2.290 6.800 -2.100 ;
      LAYER met1 ;
        RECT 6.610 0.770 6.800 2.230 ;
        RECT 6.610 0.740 6.830 0.770 ;
        RECT 6.590 0.470 6.840 0.740 ;
        RECT 6.600 0.460 6.840 0.470 ;
        RECT 6.600 0.220 6.830 0.460 ;
        RECT 6.640 -1.810 6.800 0.220 ;
        RECT 6.600 -2.050 6.830 -1.810 ;
        RECT 6.600 -2.060 6.840 -2.050 ;
        RECT 6.590 -2.330 6.840 -2.060 ;
        RECT 6.610 -2.360 6.830 -2.330 ;
        RECT 6.610 -3.820 6.800 -2.360 ;
  END
END sky130_hilas_FGBias2x1cell

MACRO sky130_hilas_TgateSingle01Part2
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TgateSingle01Part2 ;
  ORIGIN 0.670 1.810 ;
  SIZE 1.630 BY 1.430 ;
  OBS
      LAYER nwell ;
        RECT -0.180 -0.970 0.960 -0.380 ;
        RECT -0.670 -1.810 0.960 -0.970 ;
      LAYER li1 ;
        RECT -0.180 -0.880 0.960 -0.700 ;
        RECT -0.140 -1.410 0.030 -1.250 ;
        RECT 0.740 -1.320 0.930 -1.290 ;
        RECT 0.720 -1.330 0.930 -1.320 ;
        RECT -0.270 -1.450 0.050 -1.410 ;
        RECT -0.270 -1.640 0.060 -1.450 ;
        RECT 0.470 -1.500 0.930 -1.330 ;
        RECT 0.740 -1.520 0.930 -1.500 ;
        RECT -0.270 -1.670 0.050 -1.640 ;
      LAYER mcon ;
        RECT -0.210 -1.630 -0.040 -1.460 ;
        RECT 0.750 -1.490 0.920 -1.320 ;
      LAYER met1 ;
        RECT 0.670 -0.790 0.930 -0.470 ;
        RECT 0.740 -1.260 0.930 -0.790 ;
        RECT -0.280 -1.700 0.040 -1.380 ;
        RECT 0.720 -1.550 0.950 -1.260 ;
      LAYER via ;
        RECT 0.670 -0.760 0.930 -0.500 ;
        RECT -0.250 -1.670 0.010 -1.410 ;
      LAYER met2 ;
        RECT 0.640 -0.520 0.960 -0.500 ;
        RECT 0.590 -0.720 0.960 -0.520 ;
        RECT 0.640 -0.760 0.960 -0.720 ;
        RECT -0.670 -1.500 -0.450 -1.490 ;
        RECT -0.280 -1.500 0.030 -1.370 ;
        RECT -0.670 -1.700 0.960 -1.500 ;
        RECT -0.670 -1.710 -0.450 -1.700 ;
  END
END sky130_hilas_TgateSingle01Part2

MACRO sky130_hilas_DAC5bit01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_DAC5bit01 ;
  ORIGIN -3.820 -5.240 ;
  SIZE 16.580 BY 5.970 ;
  PIN A0
    USE ANALOG ;
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER li1 ;
        RECT 12.090 7.980 12.260 8.000 ;
        RECT 12.070 7.550 12.280 7.980 ;
      LAYER mcon ;
        RECT 12.090 7.830 12.260 8.000 ;
      LAYER met1 ;
        RECT 12.060 7.770 12.290 8.060 ;
        RECT 12.070 7.550 12.290 7.770 ;
        RECT 12.110 6.290 12.290 7.550 ;
        RECT 12.110 5.970 12.370 6.290 ;
      LAYER via ;
        RECT 12.110 6.000 12.370 6.260 ;
      LAYER met2 ;
        RECT 12.080 6.230 12.400 6.260 ;
        RECT 3.820 6.030 12.400 6.230 ;
        RECT 12.080 6.000 12.400 6.030 ;
    END
  END A0
  PIN A2
    USE ANALOG ;
    ANTENNAGATEAREA 0.608400 ;
    PORT
      LAYER li1 ;
        RECT 13.850 10.720 14.060 11.150 ;
        RECT 13.870 10.700 14.040 10.720 ;
      LAYER met1 ;
        RECT 13.800 10.870 14.120 11.190 ;
        RECT 13.840 10.640 14.070 10.870 ;
      LAYER via ;
        RECT 13.830 10.900 14.090 11.160 ;
      LAYER met2 ;
        RECT 13.800 10.890 14.120 11.190 ;
        RECT 13.800 10.870 14.130 10.890 ;
        RECT 13.930 8.330 14.130 10.870 ;
        RECT 3.820 8.120 14.130 8.330 ;
    END
  END A2
  PIN A3
    USE ANALOG ;
    ANTENNAGATEAREA 2.281500 ;
    PORT
      LAYER li1 ;
        RECT 7.210 10.740 7.640 10.760 ;
        RECT 7.190 10.570 7.640 10.740 ;
        RECT 12.240 10.710 12.450 11.140 ;
        RECT 12.260 10.690 12.430 10.710 ;
        RECT 7.210 10.550 7.640 10.570 ;
        RECT 4.080 9.400 4.290 9.830 ;
        RECT 4.100 9.380 4.270 9.400 ;
        RECT 10.560 8.460 10.770 8.890 ;
        RECT 10.580 8.440 10.750 8.460 ;
        RECT 13.810 6.550 14.020 6.980 ;
        RECT 13.830 6.530 14.000 6.550 ;
      LAYER met1 ;
        RECT 12.190 10.860 12.510 11.180 ;
        RECT 7.360 10.770 7.680 10.810 ;
        RECT 7.130 10.540 7.680 10.770 ;
        RECT 12.230 10.630 12.460 10.860 ;
        RECT 7.360 10.490 7.680 10.540 ;
        RECT 4.030 9.550 4.350 9.870 ;
        RECT 4.070 9.320 4.300 9.550 ;
        RECT 10.560 8.800 14.010 8.970 ;
        RECT 10.560 8.670 10.780 8.800 ;
        RECT 10.550 8.380 10.780 8.670 ;
        RECT 13.810 6.980 14.010 8.800 ;
        RECT 13.810 6.760 14.030 6.980 ;
        RECT 13.800 6.470 14.030 6.760 ;
      LAYER via ;
        RECT 12.220 10.890 12.480 11.150 ;
        RECT 7.390 10.520 7.650 10.780 ;
        RECT 4.060 9.580 4.320 9.840 ;
      LAYER met2 ;
        RECT 12.190 10.860 12.510 11.180 ;
        RECT 7.360 10.660 7.680 10.810 ;
        RECT 7.300 10.490 7.680 10.660 ;
        RECT 3.820 10.200 5.880 10.260 ;
        RECT 7.300 10.200 7.520 10.490 ;
        RECT 12.220 10.210 12.470 10.860 ;
        RECT 12.220 10.200 12.500 10.210 ;
        RECT 3.820 10.050 12.500 10.200 ;
        RECT 4.080 9.870 4.280 10.050 ;
        RECT 5.720 9.900 12.500 10.050 ;
        RECT 4.030 9.550 4.350 9.870 ;
    END
  END A3
  PIN A4
    USE ANALOG ;
    ANTENNAGATEAREA 3.650400 ;
    PORT
      LAYER li1 ;
        RECT 4.220 10.710 4.430 11.140 ;
        RECT 5.810 10.720 6.020 11.150 ;
        RECT 4.240 10.690 4.410 10.710 ;
        RECT 5.830 10.700 6.000 10.720 ;
        RECT 9.010 10.710 9.220 11.140 ;
        RECT 10.620 10.710 10.830 11.140 ;
        RECT 9.030 10.690 9.200 10.710 ;
        RECT 10.640 10.690 10.810 10.710 ;
      LAYER met1 ;
        RECT 4.170 10.860 4.490 11.180 ;
        RECT 5.760 10.870 6.080 11.190 ;
        RECT 4.210 10.630 4.440 10.860 ;
        RECT 5.800 10.640 6.030 10.870 ;
        RECT 8.960 10.860 9.280 11.180 ;
        RECT 10.570 10.860 10.890 11.180 ;
        RECT 9.000 10.630 9.230 10.860 ;
        RECT 10.610 10.630 10.840 10.860 ;
      LAYER via ;
        RECT 4.200 10.890 4.460 11.150 ;
        RECT 5.790 10.900 6.050 11.160 ;
        RECT 8.990 10.890 9.250 11.150 ;
        RECT 10.600 10.890 10.860 11.150 ;
      LAYER met2 ;
        RECT 3.820 11.180 10.870 11.210 ;
        RECT 3.820 11.020 10.890 11.180 ;
        RECT 3.820 11.000 3.970 11.020 ;
        RECT 4.170 10.860 4.490 11.020 ;
        RECT 5.760 10.870 6.080 11.020 ;
        RECT 8.960 10.860 9.280 11.020 ;
        RECT 10.570 10.860 10.890 11.020 ;
    END
  END A4
  PIN VPWR
    USE ANALOG ;
    ANTENNADIFFAREA 3.264300 ;
    PORT
      LAYER li1 ;
        RECT 16.770 11.040 16.980 11.050 ;
        RECT 16.660 11.000 16.980 11.040 ;
        RECT 17.330 11.000 17.650 11.040 ;
        RECT 16.660 10.810 16.990 11.000 ;
        RECT 17.330 10.810 17.660 11.000 ;
        RECT 16.660 10.780 16.980 10.810 ;
        RECT 17.330 10.780 17.650 10.810 ;
        RECT 7.800 10.270 7.970 10.280 ;
        RECT 16.770 10.270 16.980 10.780 ;
        RECT 17.440 10.270 17.610 10.780 ;
        RECT 6.190 10.040 17.620 10.270 ;
        RECT 6.190 9.700 6.360 10.040 ;
        RECT 7.800 9.700 7.970 10.040 ;
        RECT 6.180 9.370 6.360 9.700 ;
        RECT 7.790 9.370 7.970 9.700 ;
        RECT 6.190 8.740 6.360 9.370 ;
        RECT 7.800 8.740 7.970 9.370 ;
        RECT 6.180 8.410 6.360 8.740 ;
        RECT 7.790 8.410 7.970 8.740 ;
        RECT 6.190 7.780 6.360 8.410 ;
        RECT 7.800 7.780 7.970 8.410 ;
        RECT 6.180 7.450 6.360 7.780 ;
        RECT 7.790 7.450 7.970 7.780 ;
        RECT 6.190 6.820 6.360 7.450 ;
        RECT 7.800 6.820 7.970 7.450 ;
        RECT 6.180 6.490 6.360 6.820 ;
        RECT 7.790 6.490 7.970 6.820 ;
        RECT 6.190 6.480 6.360 6.490 ;
        RECT 7.800 6.480 7.970 6.490 ;
        RECT 9.390 9.700 9.560 10.040 ;
        RECT 9.390 9.370 9.570 9.700 ;
        RECT 9.390 8.740 9.560 9.370 ;
        RECT 9.390 8.410 9.570 8.740 ;
        RECT 9.390 7.780 9.560 8.410 ;
        RECT 9.390 7.450 9.570 7.780 ;
        RECT 9.390 6.820 9.560 7.450 ;
        RECT 9.390 6.490 9.570 6.820 ;
        RECT 9.390 6.480 9.560 6.490 ;
        RECT 11.010 6.480 11.180 10.040 ;
        RECT 12.630 9.700 12.800 10.040 ;
        RECT 12.620 9.370 12.800 9.700 ;
        RECT 12.630 8.740 12.800 9.370 ;
        RECT 12.620 8.410 12.800 8.740 ;
        RECT 12.630 6.820 12.800 8.410 ;
        RECT 12.620 6.500 12.800 6.820 ;
        RECT 12.620 6.490 12.790 6.500 ;
        RECT 14.230 6.490 14.400 10.040 ;
        RECT 15.840 6.490 16.010 10.040 ;
        RECT 17.450 6.470 17.620 10.040 ;
      LAYER mcon ;
        RECT 16.720 10.820 16.890 10.990 ;
        RECT 17.390 10.820 17.560 10.990 ;
      LAYER met1 ;
        RECT 16.650 10.750 16.970 11.070 ;
        RECT 17.320 10.750 17.640 11.070 ;
      LAYER via ;
        RECT 16.680 10.780 16.940 11.040 ;
        RECT 17.350 10.780 17.610 11.040 ;
      LAYER met2 ;
        RECT 16.530 10.930 17.690 11.210 ;
        RECT 16.650 10.750 16.960 10.930 ;
        RECT 17.280 10.920 17.690 10.930 ;
        RECT 17.320 10.750 17.630 10.920 ;
    END
  END VPWR
  PIN DRAIN
    USE ANALOG ;
    ANTENNADIFFAREA 3.264300 ;
    PORT
      LAYER li1 ;
        RECT 6.850 9.700 7.020 9.710 ;
        RECT 6.850 9.370 7.030 9.700 ;
        RECT 8.470 9.670 8.640 9.700 ;
        RECT 8.470 9.370 8.650 9.670 ;
        RECT 6.850 8.740 7.020 9.370 ;
        RECT 8.480 8.740 8.650 9.370 ;
        RECT 6.850 8.410 7.030 8.740 ;
        RECT 8.470 8.410 8.650 8.740 ;
        RECT 6.850 7.780 7.020 8.410 ;
        RECT 8.480 7.780 8.650 8.410 ;
        RECT 6.850 7.450 7.030 7.780 ;
        RECT 8.470 7.450 8.650 7.780 ;
        RECT 6.850 6.820 7.020 7.450 ;
        RECT 8.480 6.820 8.650 7.450 ;
        RECT 6.850 6.490 7.030 6.820 ;
        RECT 8.470 6.490 8.650 6.820 ;
        RECT 6.850 5.500 7.020 6.490 ;
        RECT 8.480 5.500 8.650 6.490 ;
        RECT 10.080 5.500 10.250 9.750 ;
        RECT 11.690 9.370 11.870 9.700 ;
        RECT 11.700 8.740 11.870 9.370 ;
        RECT 11.690 8.410 11.870 8.740 ;
        RECT 11.700 7.780 11.870 8.410 ;
        RECT 11.690 7.450 11.870 7.780 ;
        RECT 11.700 6.820 11.870 7.450 ;
        RECT 11.690 6.490 11.870 6.820 ;
        RECT 11.700 5.500 11.870 6.490 ;
        RECT 13.300 5.500 13.470 9.750 ;
        RECT 14.920 9.700 15.090 9.750 ;
        RECT 14.910 9.370 15.090 9.700 ;
        RECT 14.920 8.740 15.090 9.370 ;
        RECT 14.910 8.410 15.090 8.740 ;
        RECT 14.920 7.780 15.090 8.410 ;
        RECT 14.910 7.450 15.090 7.780 ;
        RECT 14.920 6.820 15.090 7.450 ;
        RECT 14.910 6.490 15.090 6.820 ;
        RECT 14.920 5.500 15.090 6.490 ;
        RECT 16.520 5.500 16.690 9.730 ;
        RECT 18.130 5.500 18.300 9.910 ;
        RECT 6.850 5.270 7.040 5.500 ;
        RECT 8.470 5.270 8.660 5.500 ;
        RECT 10.070 5.270 10.260 5.500 ;
        RECT 11.690 5.270 11.880 5.500 ;
        RECT 13.290 5.270 13.480 5.500 ;
        RECT 14.910 5.270 15.100 5.500 ;
        RECT 16.510 5.270 16.700 5.500 ;
        RECT 18.120 5.270 18.310 5.500 ;
        RECT 6.850 5.250 7.020 5.270 ;
        RECT 8.480 5.250 8.650 5.270 ;
        RECT 10.080 5.250 10.250 5.270 ;
        RECT 11.700 5.250 11.870 5.270 ;
        RECT 13.300 5.250 13.470 5.270 ;
        RECT 14.920 5.250 15.090 5.270 ;
        RECT 16.520 5.250 16.690 5.270 ;
        RECT 18.130 5.250 18.300 5.270 ;
      LAYER mcon ;
        RECT 6.860 5.300 7.030 5.470 ;
        RECT 8.480 5.300 8.650 5.470 ;
        RECT 10.080 5.300 10.250 5.470 ;
        RECT 11.700 5.300 11.870 5.470 ;
        RECT 13.300 5.300 13.470 5.470 ;
        RECT 14.920 5.300 15.090 5.470 ;
        RECT 16.520 5.300 16.690 5.470 ;
        RECT 18.130 5.300 18.300 5.470 ;
      LAYER met1 ;
        RECT 6.830 5.480 7.060 5.530 ;
        RECT 8.450 5.480 8.680 5.530 ;
        RECT 10.050 5.480 10.280 5.530 ;
        RECT 11.670 5.480 11.900 5.530 ;
        RECT 13.270 5.480 13.500 5.530 ;
        RECT 14.890 5.480 15.120 5.530 ;
        RECT 16.490 5.480 16.720 5.530 ;
        RECT 18.100 5.480 18.330 5.530 ;
        RECT 6.830 5.250 20.400 5.480 ;
        RECT 6.830 5.240 7.060 5.250 ;
        RECT 8.450 5.240 8.680 5.250 ;
        RECT 10.050 5.240 10.280 5.250 ;
        RECT 11.670 5.240 11.900 5.250 ;
        RECT 13.270 5.240 13.500 5.250 ;
        RECT 14.890 5.240 15.120 5.250 ;
        RECT 16.490 5.240 16.720 5.250 ;
        RECT 18.100 5.240 18.330 5.250 ;
    END
  END DRAIN
  OBS
      LAYER nwell ;
        RECT 4.190 5.270 20.290 10.920 ;
      LAYER li1 ;
        RECT 15.460 10.720 15.670 11.150 ;
        RECT 15.480 10.700 15.650 10.720 ;
        RECT 4.140 8.450 4.350 8.880 ;
        RECT 4.160 8.430 4.330 8.450 ;
        RECT 4.140 7.510 4.350 7.940 ;
        RECT 4.160 7.490 4.330 7.510 ;
      LAYER met1 ;
        RECT 15.410 10.870 15.730 11.190 ;
        RECT 15.450 10.640 15.680 10.870 ;
        RECT 4.090 8.600 4.410 8.920 ;
        RECT 4.130 8.370 4.360 8.600 ;
        RECT 4.090 7.660 4.410 7.980 ;
        RECT 4.130 7.430 4.360 7.660 ;
      LAYER via ;
        RECT 15.440 10.900 15.700 11.160 ;
        RECT 4.120 8.630 4.380 8.890 ;
        RECT 4.120 7.690 4.380 7.950 ;
      LAYER met2 ;
        RECT 15.410 10.870 15.730 11.190 ;
        RECT 4.090 8.600 4.410 8.920 ;
        RECT 4.090 7.660 4.410 7.980 ;
        RECT 15.530 7.350 15.680 10.870 ;
        RECT 3.820 7.150 15.690 7.350 ;
  END
END sky130_hilas_DAC5bit01

MACRO sky130_hilas_swc4x1cellOverlap2
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc4x1cellOverlap2 ;
  ORIGIN 1.910 3.820 ;
  SIZE 9.350 BY 6.050 ;
  OBS
      LAYER nwell ;
        RECT 0.880 2.220 7.430 2.230 ;
        RECT 0.880 -3.800 7.440 2.220 ;
        RECT 0.880 -3.810 7.430 -3.800 ;
        RECT 0.880 -3.820 4.880 -3.810 ;
      LAYER li1 ;
        RECT -0.850 1.020 -0.680 1.910 ;
        RECT 1.230 0.920 4.540 1.900 ;
        RECT 4.980 1.820 5.300 1.830 ;
        RECT 4.980 1.650 5.560 1.820 ;
        RECT 4.980 1.600 5.310 1.650 ;
        RECT 4.980 1.570 5.300 1.600 ;
        RECT 6.840 1.550 7.040 1.900 ;
        RECT 4.980 1.240 5.300 1.280 ;
        RECT 4.980 1.200 5.310 1.240 ;
        RECT 4.980 1.030 5.560 1.200 ;
        RECT 4.980 1.020 5.300 1.030 ;
        RECT 6.110 0.960 6.310 1.530 ;
        RECT 6.840 1.520 7.050 1.550 ;
        RECT 6.830 0.930 7.050 1.520 ;
        RECT -0.850 -0.500 -0.680 0.390 ;
        RECT 1.230 -0.550 4.540 0.430 ;
        RECT 4.980 0.390 5.300 0.400 ;
        RECT 4.980 0.220 5.560 0.390 ;
        RECT 4.980 0.180 5.310 0.220 ;
        RECT 4.980 0.140 5.300 0.180 ;
        RECT 6.110 -0.110 6.310 0.460 ;
        RECT 6.830 -0.100 7.050 0.490 ;
        RECT 6.840 -0.130 7.050 -0.100 ;
        RECT 4.980 -0.180 5.300 -0.150 ;
        RECT 4.980 -0.230 5.310 -0.180 ;
        RECT 4.980 -0.400 5.560 -0.230 ;
        RECT 4.980 -0.410 5.300 -0.400 ;
        RECT 6.840 -0.480 7.040 -0.130 ;
        RECT 6.230 -0.880 6.670 -0.710 ;
        RECT -0.850 -1.950 -0.680 -1.060 ;
        RECT 1.230 -2.020 4.540 -1.040 ;
        RECT 4.980 -1.190 5.300 -1.180 ;
        RECT 4.980 -1.360 5.560 -1.190 ;
        RECT 4.980 -1.410 5.310 -1.360 ;
        RECT 4.980 -1.440 5.300 -1.410 ;
        RECT 6.840 -1.460 7.040 -1.110 ;
        RECT 4.980 -1.770 5.300 -1.730 ;
        RECT 4.980 -1.810 5.310 -1.770 ;
        RECT 4.980 -1.980 5.560 -1.810 ;
        RECT 4.980 -1.990 5.300 -1.980 ;
        RECT 6.110 -2.050 6.310 -1.480 ;
        RECT 6.840 -1.490 7.050 -1.460 ;
        RECT 6.830 -2.080 7.050 -1.490 ;
        RECT -0.850 -3.490 -0.680 -2.600 ;
        RECT 1.230 -3.490 4.540 -2.510 ;
        RECT 4.980 -2.610 5.300 -2.600 ;
        RECT 4.980 -2.780 5.560 -2.610 ;
        RECT 4.980 -2.820 5.310 -2.780 ;
        RECT 4.980 -2.860 5.300 -2.820 ;
        RECT 6.110 -3.110 6.310 -2.540 ;
        RECT 6.830 -3.100 7.050 -2.510 ;
        RECT 6.840 -3.130 7.050 -3.100 ;
        RECT 4.980 -3.180 5.300 -3.150 ;
        RECT 4.980 -3.230 5.310 -3.180 ;
        RECT 4.980 -3.400 5.560 -3.230 ;
        RECT 4.980 -3.410 5.300 -3.400 ;
        RECT 6.840 -3.480 7.040 -3.130 ;
      LAYER mcon ;
        RECT -0.850 1.710 -0.680 1.880 ;
        RECT 2.800 1.670 2.970 1.840 ;
        RECT 5.040 1.610 5.210 1.780 ;
        RECT 2.800 1.320 2.970 1.490 ;
        RECT 6.120 1.320 6.290 1.490 ;
        RECT 2.800 0.980 2.970 1.150 ;
        RECT 5.040 1.060 5.210 1.230 ;
        RECT 6.850 1.350 7.020 1.520 ;
        RECT -0.850 0.190 -0.680 0.360 ;
        RECT 2.800 0.200 2.970 0.370 ;
        RECT 5.040 0.190 5.210 0.360 ;
        RECT 2.800 -0.150 2.970 0.020 ;
        RECT 6.120 -0.070 6.290 0.100 ;
        RECT 6.850 -0.100 7.020 0.070 ;
        RECT 2.800 -0.490 2.970 -0.320 ;
        RECT 5.040 -0.360 5.210 -0.190 ;
        RECT 6.490 -0.880 6.670 -0.710 ;
        RECT -0.850 -1.260 -0.680 -1.090 ;
        RECT 2.800 -1.270 2.970 -1.100 ;
        RECT 5.040 -1.400 5.210 -1.230 ;
        RECT 2.800 -1.620 2.970 -1.450 ;
        RECT 6.120 -1.690 6.290 -1.520 ;
        RECT 2.800 -1.960 2.970 -1.790 ;
        RECT 5.040 -1.950 5.210 -1.780 ;
        RECT 6.850 -1.660 7.020 -1.490 ;
        RECT -0.850 -2.800 -0.680 -2.630 ;
        RECT 2.800 -2.740 2.970 -2.570 ;
        RECT 5.040 -2.810 5.210 -2.640 ;
        RECT 2.800 -3.090 2.970 -2.920 ;
        RECT 6.120 -3.070 6.290 -2.900 ;
        RECT 6.850 -3.100 7.020 -2.930 ;
        RECT 2.800 -3.430 2.970 -3.260 ;
        RECT 5.040 -3.360 5.210 -3.190 ;
      LAYER met1 ;
        RECT -0.900 -3.820 -0.630 2.230 ;
        RECT 2.760 1.260 3.000 1.900 ;
        RECT 4.970 1.540 5.290 1.860 ;
        RECT 6.110 1.550 6.270 2.230 ;
        RECT 6.110 1.530 6.310 1.550 ;
        RECT 2.770 1.000 3.000 1.260 ;
        RECT 2.770 0.780 3.010 1.000 ;
        RECT 4.970 0.990 5.290 1.310 ;
        RECT 6.090 1.290 6.320 1.530 ;
        RECT 6.110 1.070 6.310 1.290 ;
        RECT 6.480 1.240 6.670 2.230 ;
        RECT 6.920 1.580 7.080 2.230 ;
        RECT 6.500 1.120 6.670 1.240 ;
        RECT 2.760 -0.210 3.000 0.430 ;
        RECT 4.970 0.110 5.290 0.430 ;
        RECT 6.110 0.350 6.270 1.070 ;
        RECT 6.110 0.130 6.310 0.350 ;
        RECT 6.510 0.300 6.670 1.120 ;
        RECT 6.810 1.030 7.080 1.580 ;
        RECT 6.810 0.980 7.090 1.030 ;
        RECT 6.920 0.890 7.090 0.980 ;
        RECT 6.920 0.530 7.080 0.890 ;
        RECT 6.920 0.440 7.090 0.530 ;
        RECT 6.500 0.180 6.670 0.300 ;
        RECT 6.090 -0.110 6.320 0.130 ;
        RECT 2.770 -0.470 3.000 -0.210 ;
        RECT 4.970 -0.440 5.290 -0.120 ;
        RECT 6.110 -0.130 6.310 -0.110 ;
        RECT 2.770 -0.690 3.010 -0.470 ;
        RECT 2.760 -1.680 3.000 -1.040 ;
        RECT 4.970 -1.470 5.290 -1.150 ;
        RECT 6.110 -1.460 6.270 -0.130 ;
        RECT 6.480 -0.680 6.670 0.180 ;
        RECT 6.810 0.390 7.090 0.440 ;
        RECT 6.810 -0.160 7.080 0.390 ;
        RECT 6.460 -0.910 6.700 -0.680 ;
        RECT 6.110 -1.480 6.310 -1.460 ;
        RECT 2.770 -1.940 3.000 -1.680 ;
        RECT 2.770 -2.160 3.010 -1.940 ;
        RECT 4.970 -2.020 5.290 -1.700 ;
        RECT 6.090 -1.720 6.320 -1.480 ;
        RECT 6.110 -1.940 6.310 -1.720 ;
        RECT 6.480 -1.770 6.670 -0.910 ;
        RECT 6.920 -1.430 7.080 -0.160 ;
        RECT 6.500 -1.890 6.670 -1.770 ;
        RECT 2.760 -3.150 3.000 -2.510 ;
        RECT 4.970 -2.890 5.290 -2.570 ;
        RECT 6.110 -2.650 6.270 -1.940 ;
        RECT 6.110 -2.870 6.310 -2.650 ;
        RECT 6.510 -2.700 6.670 -1.890 ;
        RECT 6.810 -1.980 7.080 -1.430 ;
        RECT 6.810 -2.030 7.090 -1.980 ;
        RECT 6.920 -2.120 7.090 -2.030 ;
        RECT 6.920 -2.470 7.080 -2.120 ;
        RECT 6.920 -2.560 7.090 -2.470 ;
        RECT 6.500 -2.820 6.670 -2.700 ;
        RECT 6.090 -3.110 6.320 -2.870 ;
        RECT 2.770 -3.410 3.000 -3.150 ;
        RECT 2.770 -3.630 3.010 -3.410 ;
        RECT 4.970 -3.440 5.290 -3.120 ;
        RECT 6.110 -3.130 6.310 -3.110 ;
        RECT 6.110 -3.810 6.270 -3.130 ;
        RECT 6.480 -3.810 6.670 -2.820 ;
        RECT 6.810 -2.610 7.090 -2.560 ;
        RECT 6.810 -3.160 7.080 -2.610 ;
        RECT 6.920 -3.810 7.080 -3.160 ;
      LAYER via ;
        RECT 5.000 1.570 5.260 1.830 ;
        RECT 5.000 1.020 5.260 1.280 ;
        RECT 5.000 0.140 5.260 0.400 ;
        RECT 5.000 -0.410 5.260 -0.150 ;
        RECT 5.000 -1.440 5.260 -1.180 ;
        RECT 5.000 -1.990 5.260 -1.730 ;
        RECT 5.000 -2.860 5.260 -2.600 ;
        RECT 5.000 -3.410 5.260 -3.150 ;
      LAYER met2 ;
        RECT 4.970 1.730 5.280 1.870 ;
        RECT -1.910 1.550 7.440 1.730 ;
        RECT 4.970 1.540 5.280 1.550 ;
        RECT 4.970 1.300 5.280 1.320 ;
        RECT -1.910 1.120 7.440 1.300 ;
        RECT 4.970 0.990 5.280 1.120 ;
        RECT 4.970 0.300 5.280 0.430 ;
        RECT -1.910 0.120 7.440 0.300 ;
        RECT 4.970 0.100 5.280 0.120 ;
        RECT 4.970 -0.130 5.280 -0.120 ;
        RECT -1.910 -0.200 4.960 -0.130 ;
        RECT 4.970 -0.200 7.440 -0.130 ;
        RECT -1.910 -0.310 7.440 -0.200 ;
        RECT 4.970 -0.450 5.280 -0.310 ;
        RECT 4.970 -1.280 5.280 -1.140 ;
        RECT 4.970 -1.290 7.440 -1.280 ;
        RECT -1.910 -1.460 7.440 -1.290 ;
        RECT 4.970 -1.470 5.280 -1.460 ;
        RECT 4.970 -1.710 5.280 -1.690 ;
        RECT -1.910 -1.880 7.440 -1.710 ;
        RECT 4.880 -1.890 7.440 -1.880 ;
        RECT 4.970 -2.020 5.280 -1.890 ;
        RECT 4.970 -2.690 5.280 -2.570 ;
        RECT -1.910 -2.700 5.280 -2.690 ;
        RECT -1.910 -2.860 7.440 -2.700 ;
        RECT 4.880 -2.880 7.440 -2.860 ;
        RECT 4.970 -2.900 5.280 -2.880 ;
        RECT 4.970 -3.130 5.280 -3.120 ;
        RECT -1.910 -3.300 7.440 -3.130 ;
        RECT 4.970 -3.310 7.440 -3.300 ;
        RECT 4.970 -3.450 5.280 -3.310 ;
  END
END sky130_hilas_swc4x1cellOverlap2

MACRO sky130_hilas_pFETdevice01d
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pFETdevice01d ;
  ORIGIN 0.920 1.020 ;
  SIZE 1.840 BY 1.450 ;
  OBS
      LAYER nwell ;
        RECT -0.790 -0.780 0.820 0.430 ;
      LAYER li1 ;
        RECT -0.860 -0.110 -0.650 0.320 ;
        RECT -0.840 -0.130 -0.670 -0.110 ;
        RECT -0.410 -0.160 -0.240 0.170 ;
        RECT 0.270 -0.160 0.440 0.170 ;
        RECT 0.670 -0.590 0.840 -0.570 ;
        RECT 0.650 -1.020 0.860 -0.590 ;
      LAYER mcon ;
        RECT 0.670 -0.740 0.840 -0.570 ;
      LAYER met1 ;
        RECT -0.860 0.100 -0.640 0.320 ;
        RECT -0.870 -0.190 -0.640 0.100 ;
        RECT 0.640 -0.800 0.870 -0.510 ;
        RECT 0.650 -1.020 0.870 -0.800 ;
  END
END sky130_hilas_pFETdevice01d

MACRO sky130_hilas_pTransistorPair
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pTransistorPair ;
  ORIGIN -1.330 4.400 ;
  SIZE 1.870 BY 6.050 ;
  OBS
      LAYER nwell ;
        RECT 1.330 -4.390 3.190 1.650 ;
      LAYER li1 ;
        RECT 1.740 -2.730 1.920 1.180 ;
        RECT 2.550 -0.610 2.720 1.170 ;
        RECT 2.470 -0.670 3.010 -0.610 ;
        RECT 2.470 -0.780 3.020 -0.670 ;
        RECT 2.830 -0.900 3.020 -0.780 ;
        RECT 2.300 -1.200 2.470 -1.040 ;
        RECT 2.300 -1.370 2.520 -1.200 ;
        RECT 2.350 -1.450 2.520 -1.370 ;
        RECT 2.350 -1.490 2.670 -1.450 ;
        RECT 2.350 -1.680 2.680 -1.490 ;
        RECT 2.350 -1.710 2.670 -1.680 ;
        RECT 1.620 -2.770 1.940 -2.730 ;
        RECT 1.620 -2.960 1.950 -2.770 ;
        RECT 1.620 -2.990 1.940 -2.960 ;
        RECT 1.740 -3.920 1.920 -2.990 ;
        RECT 2.550 -3.260 2.720 -1.880 ;
        RECT 2.550 -3.520 3.030 -3.260 ;
        RECT 2.550 -3.660 2.800 -3.520 ;
        RECT 2.470 -3.830 2.800 -3.660 ;
        RECT 2.320 -4.090 2.490 -4.070 ;
        RECT 2.320 -4.350 2.880 -4.090 ;
        RECT 2.320 -4.400 2.490 -4.350 ;
      LAYER mcon ;
        RECT 2.840 -0.870 3.010 -0.700 ;
        RECT 2.410 -1.670 2.580 -1.500 ;
        RECT 1.680 -2.950 1.850 -2.780 ;
        RECT 2.800 -3.470 2.970 -3.300 ;
        RECT 2.650 -4.300 2.820 -4.130 ;
      LAYER met1 ;
        RECT 2.810 -0.930 3.040 -0.640 ;
        RECT 2.340 -1.740 2.660 -1.420 ;
        RECT 2.830 -2.220 3.040 -0.930 ;
        RECT 2.810 -2.540 3.070 -2.220 ;
        RECT 2.830 -2.650 3.040 -2.540 ;
        RECT 1.610 -3.020 1.930 -2.700 ;
        RECT 2.720 -3.550 3.040 -3.230 ;
        RECT 2.570 -4.380 2.890 -4.060 ;
      LAYER via ;
        RECT 2.370 -1.710 2.630 -1.450 ;
        RECT 2.810 -2.510 3.070 -2.250 ;
        RECT 1.640 -2.990 1.900 -2.730 ;
        RECT 2.750 -3.520 3.010 -3.260 ;
        RECT 2.600 -4.350 2.860 -4.090 ;
      LAYER met2 ;
        RECT 2.340 -1.460 2.650 -1.410 ;
        RECT 2.250 -1.690 3.120 -1.460 ;
        RECT 2.250 -1.700 2.680 -1.690 ;
        RECT 2.340 -1.740 2.650 -1.700 ;
        RECT 2.730 -2.490 3.200 -2.240 ;
        RECT 2.780 -2.510 3.100 -2.490 ;
        RECT 1.610 -3.020 1.920 -2.690 ;
        RECT 2.730 -3.270 3.040 -3.230 ;
        RECT 2.550 -3.520 3.100 -3.270 ;
        RECT 2.730 -3.560 3.040 -3.520 ;
        RECT 2.580 -4.130 2.890 -4.060 ;
        RECT 2.010 -4.380 2.890 -4.130 ;
        RECT 2.580 -4.390 2.890 -4.380 ;
  END
END sky130_hilas_pTransistorPair

MACRO sky130_hilas_TA2Cell_1FG_Strong
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TA2Cell_1FG_Strong ;
  ORIGIN 26.170 -1.400 ;
  SIZE 28.100 BY 6.050 ;
  PIN VINP_AMP2
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER li1 ;
        RECT -2.190 4.730 -1.870 4.760 ;
        RECT -2.190 4.540 -1.860 4.730 ;
        RECT -2.190 4.500 -1.870 4.540 ;
        RECT -2.190 4.420 -2.020 4.500 ;
        RECT -2.240 4.250 -2.020 4.420 ;
        RECT -2.240 4.090 -2.070 4.250 ;
      LAYER mcon ;
        RECT -2.130 4.550 -1.960 4.720 ;
      LAYER met1 ;
        RECT -2.200 4.470 -1.880 4.790 ;
      LAYER via ;
        RECT -2.170 4.500 -1.910 4.760 ;
      LAYER met2 ;
        RECT -2.200 4.750 -1.890 4.790 ;
        RECT -2.520 4.740 -1.860 4.750 ;
        RECT -2.520 4.510 -1.420 4.740 ;
        RECT -2.200 4.460 -1.890 4.510 ;
    END
  END VINP_AMP2
  PIN VINN_AMP2
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER li1 ;
        RECT -2.220 7.400 -2.050 7.450 ;
        RECT -2.220 7.140 -1.660 7.400 ;
        RECT -2.220 7.120 -2.050 7.140 ;
      LAYER mcon ;
        RECT -1.890 7.180 -1.720 7.350 ;
      LAYER met1 ;
        RECT -1.970 7.110 -1.650 7.430 ;
      LAYER via ;
        RECT -1.940 7.140 -1.680 7.400 ;
      LAYER met2 ;
        RECT -1.960 7.430 -1.650 7.440 ;
        RECT -2.530 7.420 -1.650 7.430 ;
        RECT -2.600 7.180 -1.650 7.420 ;
        RECT -1.960 7.110 -1.650 7.180 ;
    END
  END VINN_AMP2
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.650 1.400 1.930 7.450 ;
      LAYER li1 ;
        RECT 0.860 5.840 1.560 6.150 ;
        RECT 0.710 5.610 1.560 5.840 ;
        RECT 0.860 5.270 1.560 5.610 ;
        RECT 0.860 3.250 1.560 3.590 ;
        RECT 0.710 3.020 1.560 3.250 ;
        RECT 0.860 2.710 1.560 3.020 ;
      LAYER mcon ;
        RECT 0.720 5.640 0.890 5.810 ;
        RECT 0.720 3.050 0.890 3.220 ;
      LAYER met1 ;
        RECT 0.630 7.300 0.910 7.450 ;
        RECT 0.640 5.870 0.910 7.300 ;
        RECT 0.640 5.580 0.920 5.870 ;
        RECT 0.640 3.280 0.910 5.580 ;
        RECT 0.640 2.990 0.920 3.280 ;
        RECT 0.640 1.400 0.910 2.990 ;
    END
  END VPWR
  PIN GATECOLSELECT
    USE ANALOG ;
    ANTENNAGATEAREA 0.310000 ;
    PORT
      LAYER li1 ;
        RECT -4.160 5.980 -3.970 5.990 ;
        RECT -4.160 5.690 -3.960 5.980 ;
        RECT -4.170 5.360 -3.930 5.690 ;
        RECT -4.170 3.160 -3.930 3.490 ;
        RECT -4.160 2.870 -3.960 3.160 ;
        RECT -4.160 2.860 -3.970 2.870 ;
      LAYER mcon ;
        RECT -4.150 5.730 -3.970 5.920 ;
        RECT -4.150 2.930 -3.970 3.120 ;
      LAYER met1 ;
        RECT -4.160 5.990 -3.970 7.450 ;
        RECT -4.160 5.960 -3.940 5.990 ;
        RECT -4.180 5.690 -3.930 5.960 ;
        RECT -4.170 5.680 -3.930 5.690 ;
        RECT -4.170 5.440 -3.940 5.680 ;
        RECT -4.130 3.410 -3.970 5.440 ;
        RECT -4.170 3.170 -3.940 3.410 ;
        RECT -4.170 3.160 -3.930 3.170 ;
        RECT -4.180 2.890 -3.930 3.160 ;
        RECT -4.160 2.860 -3.940 2.890 ;
        RECT -4.160 1.400 -3.970 2.860 ;
    END
  END GATECOLSELECT
  PIN VINP_AMP1
    USE ANALOG ;
    ANTENNADIFFAREA 0.217200 ;
    PORT
      LAYER li1 ;
        RECT -23.520 7.020 -23.330 7.050 ;
        RECT -23.520 6.850 -22.460 7.020 ;
        RECT -23.520 6.820 -23.330 6.850 ;
        RECT -22.630 6.460 -22.460 6.850 ;
        RECT -22.630 6.290 -21.890 6.460 ;
        RECT -23.520 4.880 -23.330 5.060 ;
        RECT -23.590 4.710 -23.240 4.880 ;
      LAYER mcon ;
        RECT -23.510 6.850 -23.340 7.020 ;
        RECT -23.510 4.860 -23.340 5.030 ;
      LAYER met1 ;
        RECT -23.530 7.080 -23.320 7.450 ;
        RECT -23.540 6.790 -23.310 7.080 ;
        RECT -23.530 5.090 -23.320 6.790 ;
        RECT -23.540 4.800 -23.310 5.090 ;
        RECT -23.530 4.660 -23.320 4.800 ;
    END
  END VINP_AMP1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT -0.160 6.170 0.390 7.160 ;
        RECT -0.160 4.690 0.390 5.680 ;
        RECT -0.160 3.210 0.390 4.200 ;
        RECT -0.160 1.730 0.390 2.720 ;
      LAYER mcon ;
        RECT 0.060 6.580 0.230 6.750 ;
        RECT 0.060 5.100 0.230 5.270 ;
        RECT 0.060 3.620 0.230 3.790 ;
        RECT 0.060 2.140 0.230 2.310 ;
      LAYER met1 ;
        RECT -0.030 1.400 0.310 7.450 ;
    END
  END VGND
  PIN OUTPUT2
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER li1 ;
        RECT -0.750 4.160 -0.550 4.200 ;
        RECT 1.310 4.190 1.630 4.230 ;
        RECT -0.980 3.900 -0.550 4.160 ;
        RECT 0.850 4.010 1.640 4.190 ;
        RECT 1.310 4.000 1.640 4.010 ;
        RECT 1.310 3.970 1.630 4.000 ;
        RECT -0.750 3.870 -0.550 3.900 ;
      LAYER mcon ;
        RECT -0.920 3.940 -0.750 4.110 ;
        RECT 1.370 4.010 1.540 4.180 ;
      LAYER met1 ;
        RECT -0.990 3.870 -0.670 4.190 ;
        RECT 1.300 3.940 1.620 4.260 ;
      LAYER via ;
        RECT -0.960 3.900 -0.700 4.160 ;
        RECT 1.330 3.970 1.590 4.230 ;
      LAYER met2 ;
        RECT -0.990 4.140 -0.680 4.200 ;
        RECT 1.300 4.140 1.610 4.270 ;
        RECT 1.750 4.140 1.930 4.150 ;
        RECT -0.990 3.920 1.930 4.140 ;
        RECT -0.990 3.870 -0.680 3.920 ;
    END
  END OUTPUT2
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER li1 ;
        RECT -0.750 4.990 -0.550 5.020 ;
        RECT -0.980 4.730 -0.550 4.990 ;
        RECT 1.320 4.910 1.640 4.950 ;
        RECT 1.320 4.850 1.650 4.910 ;
        RECT -0.750 4.690 -0.550 4.730 ;
        RECT 0.850 4.720 1.650 4.850 ;
        RECT 0.850 4.690 1.640 4.720 ;
        RECT 0.850 4.670 1.550 4.690 ;
      LAYER mcon ;
        RECT -0.920 4.780 -0.750 4.950 ;
        RECT 1.380 4.730 1.550 4.900 ;
      LAYER met1 ;
        RECT -0.990 4.700 -0.670 5.020 ;
        RECT 1.310 4.660 1.630 4.980 ;
      LAYER via ;
        RECT -0.960 4.730 -0.700 4.990 ;
        RECT 1.340 4.690 1.600 4.950 ;
      LAYER met2 ;
        RECT -0.990 4.970 -0.680 5.020 ;
        RECT 1.310 4.970 1.620 4.990 ;
        RECT -0.990 4.740 1.930 4.970 ;
        RECT -0.990 4.690 -0.680 4.740 ;
        RECT 1.310 4.660 1.620 4.740 ;
    END
  END OUTPUT1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -6.510 7.440 -3.200 7.450 ;
        RECT -6.510 1.410 -1.350 7.440 ;
        RECT -3.210 1.400 -1.350 1.410 ;
      LAYER li1 ;
        RECT -3.800 6.770 -3.600 7.120 ;
        RECT -3.800 6.740 -3.590 6.770 ;
        RECT -4.530 4.880 -4.360 6.490 ;
        RECT -3.810 6.160 -3.590 6.740 ;
        RECT -3.800 6.150 -3.590 6.160 ;
        RECT -4.530 4.690 -4.350 4.880 ;
        RECT -4.530 3.970 -4.350 4.160 ;
        RECT -4.530 2.360 -4.360 3.970 ;
        RECT -3.800 2.690 -3.590 2.700 ;
        RECT -3.810 2.110 -3.590 2.690 ;
        RECT -3.800 2.080 -3.590 2.110 ;
        RECT -3.800 1.730 -3.600 2.080 ;
      LAYER mcon ;
        RECT -3.790 6.570 -3.620 6.740 ;
        RECT -3.790 2.110 -3.620 2.280 ;
      LAYER met1 ;
        RECT -3.720 6.800 -3.440 7.450 ;
        RECT -3.830 6.200 -3.440 6.800 ;
        RECT -4.560 4.880 -4.320 5.010 ;
        RECT -4.560 4.560 -4.300 4.880 ;
        RECT -3.720 4.600 -3.440 6.200 ;
        RECT -3.720 4.280 -3.360 4.600 ;
        RECT -4.560 3.960 -4.300 4.280 ;
        RECT -4.560 3.840 -4.320 3.960 ;
        RECT -3.720 2.650 -3.440 4.280 ;
        RECT -3.830 2.050 -3.440 2.650 ;
        RECT -3.720 1.400 -3.440 2.050 ;
      LAYER via ;
        RECT -4.560 4.590 -4.300 4.850 ;
        RECT -3.620 4.310 -3.360 4.570 ;
        RECT -4.560 3.990 -4.300 4.250 ;
      LAYER met2 ;
        RECT -4.590 4.590 -4.270 4.850 ;
        RECT -4.550 4.570 -3.370 4.590 ;
        RECT -4.550 4.310 -3.330 4.570 ;
        RECT -4.550 4.250 -3.370 4.310 ;
        RECT -4.590 4.240 -3.370 4.250 ;
        RECT -4.590 3.990 -4.270 4.240 ;
    END
  END VINJ
  OBS
      LAYER nwell ;
        RECT -26.170 1.410 -22.860 7.440 ;
        RECT -21.130 5.060 -18.410 6.710 ;
        RECT -16.380 6.700 -12.990 7.450 ;
        RECT -21.130 5.020 -18.420 5.060 ;
        RECT -21.130 3.690 -18.420 3.730 ;
        RECT -21.130 2.040 -18.410 3.690 ;
        RECT -16.390 3.130 -12.980 6.700 ;
        RECT -10.960 5.060 -8.240 6.710 ;
        RECT -10.960 5.020 -8.250 5.060 ;
        RECT -10.960 3.690 -8.250 3.730 ;
        RECT -16.380 1.410 -12.990 3.130 ;
        RECT -10.960 2.040 -8.240 3.690 ;
      LAYER li1 ;
        RECT -0.750 7.120 -0.550 7.160 ;
        RECT -25.770 6.770 -25.570 7.120 ;
        RECT -24.290 6.870 -23.760 7.040 ;
        RECT -5.610 6.870 -5.080 7.040 ;
        RECT -25.780 6.740 -25.570 6.770 ;
        RECT -25.780 6.160 -25.560 6.740 ;
        RECT -25.780 6.150 -25.570 6.160 ;
        RECT -25.400 5.980 -25.210 5.990 ;
        RECT -25.410 5.690 -25.210 5.980 ;
        RECT -25.440 5.360 -25.200 5.690 ;
        RECT -25.010 4.880 -24.840 6.490 ;
        RECT -24.180 5.390 -24.010 6.480 ;
        RECT -23.050 6.460 -22.860 6.490 ;
        RECT -23.590 6.290 -22.860 6.460 ;
        RECT -7.480 6.290 -7.130 6.460 ;
        RECT -6.110 6.290 -5.780 6.460 ;
        RECT -23.050 6.260 -22.860 6.290 ;
        RECT -20.830 5.670 -20.600 6.190 ;
        RECT -23.590 5.500 -20.600 5.670 ;
        RECT -24.410 5.350 -24.010 5.390 ;
        RECT -24.420 5.160 -24.010 5.350 ;
        RECT -15.630 5.310 -15.080 5.740 ;
        RECT -14.290 5.310 -13.740 5.740 ;
        RECT -10.660 5.500 -10.430 6.190 ;
        RECT -5.360 5.960 -5.190 6.480 ;
        RECT -2.800 6.040 -2.620 6.970 ;
        RECT -2.070 6.710 -1.740 6.880 ;
        RECT -0.980 6.860 -0.550 7.120 ;
        RECT -0.750 6.830 -0.550 6.860 ;
        RECT 1.210 7.040 1.790 7.210 ;
        RECT 1.210 6.940 1.600 7.040 ;
        RECT 1.210 6.910 1.590 6.940 ;
        RECT 1.210 6.760 1.570 6.910 ;
        RECT -1.990 6.570 -1.740 6.710 ;
        RECT 0.860 6.590 1.570 6.760 ;
        RECT -1.990 6.310 -1.510 6.570 ;
        RECT -1.160 6.470 -0.990 6.510 ;
        RECT -0.750 6.470 -0.550 6.500 ;
        RECT -5.520 5.700 -5.190 5.960 ;
        RECT -2.920 6.010 -2.600 6.040 ;
        RECT -2.920 5.820 -2.590 6.010 ;
        RECT -2.920 5.780 -2.600 5.820 ;
        RECT -7.480 5.500 -7.130 5.670 ;
        RECT -6.110 5.500 -5.780 5.670 ;
        RECT -24.410 5.130 -24.010 5.160 ;
        RECT -25.020 4.690 -24.840 4.880 ;
        RECT -24.180 4.790 -24.010 5.130 ;
        RECT -22.670 4.300 -22.460 4.730 ;
        RECT -22.240 4.710 -21.900 4.880 ;
        RECT -22.650 4.280 -22.480 4.300 ;
        RECT -25.020 3.970 -24.840 4.160 ;
        RECT -25.440 3.160 -25.200 3.490 ;
        RECT -25.410 2.870 -25.210 3.160 ;
        RECT -25.400 2.860 -25.210 2.870 ;
        RECT -25.780 2.690 -25.570 2.700 ;
        RECT -25.780 2.110 -25.560 2.690 ;
        RECT -25.010 2.360 -24.840 3.970 ;
        RECT -24.180 3.700 -24.010 4.060 ;
        RECT -23.590 3.970 -23.240 4.140 ;
        RECT -23.050 4.120 -22.860 4.170 ;
        RECT -22.150 4.140 -21.980 4.710 ;
        RECT -17.870 4.480 -17.680 4.880 ;
        RECT -11.690 4.480 -11.500 4.880 ;
        RECT -7.470 4.710 -7.130 4.880 ;
        RECT -6.110 4.710 -5.780 4.880 ;
        RECT -5.360 4.790 -5.190 5.700 ;
        RECT -17.870 4.470 -17.490 4.480 ;
        RECT -21.230 4.290 -17.490 4.470 ;
        RECT -17.870 4.250 -17.490 4.290 ;
        RECT -11.880 4.470 -11.500 4.480 ;
        RECT -11.880 4.290 -8.140 4.470 ;
        RECT -11.880 4.250 -11.500 4.290 ;
        RECT -23.050 4.110 -22.820 4.120 ;
        RECT -22.240 4.110 -21.900 4.140 ;
        RECT -23.050 3.970 -21.900 4.110 ;
        RECT -23.510 3.760 -23.320 3.970 ;
        RECT -23.050 3.940 -22.070 3.970 ;
        RECT -22.910 3.910 -22.070 3.940 ;
        RECT -17.870 3.870 -17.680 4.250 ;
        RECT -24.420 3.660 -24.010 3.700 ;
        RECT -24.430 3.470 -24.010 3.660 ;
        RECT -15.630 3.580 -15.080 4.010 ;
        RECT -14.290 3.580 -13.740 4.010 ;
        RECT -11.690 3.870 -11.500 4.250 ;
        RECT -6.030 4.140 -5.860 4.710 ;
        RECT -7.470 3.970 -7.130 4.140 ;
        RECT -6.110 3.970 -5.780 4.140 ;
        RECT -24.420 3.440 -24.010 3.470 ;
        RECT -24.180 2.370 -24.010 3.440 ;
        RECT -23.590 3.250 -20.660 3.350 ;
        RECT -23.590 3.180 -20.600 3.250 ;
        RECT -21.570 2.860 -21.400 2.920 ;
        RECT -21.590 2.650 -21.380 2.860 ;
        RECT -23.060 2.560 -22.870 2.590 ;
        RECT -21.570 2.580 -21.400 2.650 ;
        RECT -20.830 2.560 -20.600 3.180 ;
        RECT -10.660 2.560 -10.430 3.290 ;
        RECT -7.480 3.180 -7.130 3.350 ;
        RECT -6.110 3.180 -5.780 3.350 ;
        RECT -5.360 3.200 -5.190 4.060 ;
        RECT -5.520 2.940 -5.190 3.200 ;
        RECT -23.590 2.390 -22.870 2.560 ;
        RECT -23.060 2.360 -22.870 2.390 ;
        RECT -22.700 2.390 -21.890 2.560 ;
        RECT -7.480 2.390 -7.130 2.560 ;
        RECT -6.110 2.390 -5.780 2.560 ;
        RECT -25.780 2.080 -25.570 2.110 ;
        RECT -25.770 1.730 -25.570 2.080 ;
        RECT -23.490 2.050 -23.300 2.080 ;
        RECT -22.700 2.050 -22.510 2.390 ;
        RECT -5.360 2.370 -5.190 2.940 ;
        RECT -24.290 1.810 -23.760 1.980 ;
        RECT -23.490 1.870 -22.510 2.050 ;
        RECT -23.490 1.850 -23.300 1.870 ;
        RECT -5.610 1.810 -5.080 1.980 ;
        RECT -2.800 1.870 -2.620 5.780 ;
        RECT -1.990 4.930 -1.820 6.310 ;
        RECT -1.160 6.210 -0.550 6.470 ;
        RECT -1.160 6.180 -0.990 6.210 ;
        RECT -0.750 6.170 -0.550 6.210 ;
        RECT -1.160 5.640 -0.990 5.670 ;
        RECT -0.750 5.640 -0.550 5.680 ;
        RECT -1.160 5.380 -0.550 5.640 ;
        RECT -1.160 5.340 -0.990 5.380 ;
        RECT -0.750 5.350 -0.550 5.380 ;
        RECT -1.710 3.830 -1.520 3.950 ;
        RECT -2.070 3.720 -1.520 3.830 ;
        RECT -2.070 3.660 -1.530 3.720 ;
        RECT -1.990 1.880 -1.820 3.660 ;
        RECT -1.160 3.510 -0.990 3.550 ;
        RECT -0.750 3.510 -0.550 3.540 ;
        RECT -1.160 3.250 -0.550 3.510 ;
        RECT -1.160 3.220 -0.990 3.250 ;
        RECT -0.750 3.210 -0.550 3.250 ;
        RECT -1.160 2.680 -0.990 2.710 ;
        RECT -0.750 2.680 -0.550 2.720 ;
        RECT -1.160 2.420 -0.550 2.680 ;
        RECT -1.160 2.380 -0.990 2.420 ;
        RECT -0.750 2.390 -0.550 2.420 ;
        RECT 0.860 2.100 1.570 2.270 ;
        RECT -0.750 2.030 -0.550 2.060 ;
        RECT -0.980 1.770 -0.550 2.030 ;
        RECT -0.750 1.730 -0.550 1.770 ;
        RECT 1.210 1.820 1.570 2.100 ;
        RECT 1.210 1.650 1.790 1.820 ;
      LAYER mcon ;
        RECT -23.940 6.870 -23.760 7.040 ;
        RECT -25.750 6.570 -25.580 6.740 ;
        RECT -25.400 5.730 -25.220 5.920 ;
        RECT -23.040 6.290 -22.870 6.460 ;
        RECT -20.800 5.990 -20.630 6.160 ;
        RECT -10.630 5.990 -10.460 6.160 ;
        RECT -20.800 5.540 -20.630 5.710 ;
        RECT -24.320 5.170 -24.150 5.340 ;
        RECT -15.350 5.390 -15.080 5.660 ;
        RECT -14.290 5.390 -14.020 5.660 ;
        RECT -0.920 6.900 -0.750 7.070 ;
        RECT 1.330 6.950 1.500 7.120 ;
        RECT -1.740 6.350 -1.570 6.520 ;
        RECT -10.630 5.540 -10.460 5.710 ;
        RECT -5.460 5.740 -5.290 5.910 ;
        RECT -2.860 5.830 -2.690 6.000 ;
        RECT -17.670 4.280 -17.500 4.450 ;
        RECT -11.870 4.280 -11.700 4.450 ;
        RECT -25.400 2.930 -25.220 3.120 ;
        RECT -23.040 3.970 -22.870 4.140 ;
        RECT -23.500 3.790 -23.330 3.960 ;
        RECT -24.330 3.480 -24.160 3.650 ;
        RECT -15.350 3.660 -15.080 3.930 ;
        RECT -14.290 3.660 -14.020 3.930 ;
        RECT -20.800 3.040 -20.630 3.210 ;
        RECT -20.800 2.590 -20.630 2.760 ;
        RECT -10.630 3.040 -10.460 3.210 ;
        RECT -5.460 2.980 -5.290 3.150 ;
        RECT -10.630 2.590 -10.460 2.760 ;
        RECT -23.050 2.390 -22.880 2.560 ;
        RECT -25.750 2.110 -25.580 2.280 ;
        RECT -23.940 1.810 -23.760 1.980 ;
        RECT -23.480 1.880 -23.310 2.050 ;
        RECT -0.970 6.250 -0.800 6.420 ;
        RECT -0.970 5.430 -0.800 5.600 ;
        RECT -1.700 3.750 -1.530 3.920 ;
        RECT -0.970 3.290 -0.800 3.460 ;
        RECT -0.970 2.470 -0.800 2.640 ;
        RECT -0.920 1.820 -0.750 1.990 ;
        RECT 1.290 1.760 1.460 1.930 ;
      LAYER met1 ;
        RECT -25.810 6.800 -25.650 7.450 ;
        RECT -25.810 6.250 -25.540 6.800 ;
        RECT -25.820 6.200 -25.540 6.250 ;
        RECT -25.820 6.110 -25.650 6.200 ;
        RECT -25.810 2.740 -25.650 6.110 ;
        RECT -25.400 5.990 -25.210 7.450 ;
        RECT -23.990 6.770 -23.690 7.150 ;
        RECT -23.060 6.520 -22.870 7.450 ;
        RECT -23.070 6.230 -22.840 6.520 ;
        RECT -25.430 5.960 -25.210 5.990 ;
        RECT -25.440 5.690 -25.190 5.960 ;
        RECT -25.440 5.680 -25.200 5.690 ;
        RECT -25.430 5.440 -25.200 5.680 ;
        RECT -25.400 3.410 -25.240 5.440 ;
        RECT -24.400 5.100 -24.080 5.420 ;
        RECT -25.050 4.590 -24.810 5.010 ;
        RECT -25.080 4.270 -24.810 4.590 ;
        RECT -25.050 3.840 -24.810 4.270 ;
        RECT -23.060 4.200 -22.870 6.230 ;
        RECT -22.650 4.730 -22.440 7.450 ;
        RECT -22.680 4.220 -22.440 4.730 ;
        RECT -23.510 4.020 -23.320 4.150 ;
        RECT -23.530 3.730 -23.300 4.020 ;
        RECT -23.070 3.910 -22.840 4.200 ;
        RECT -24.410 3.410 -24.090 3.730 ;
        RECT -25.430 3.170 -25.200 3.410 ;
        RECT -25.440 3.160 -25.200 3.170 ;
        RECT -25.440 2.890 -25.190 3.160 ;
        RECT -25.430 2.860 -25.210 2.890 ;
        RECT -25.820 2.650 -25.650 2.740 ;
        RECT -25.820 2.600 -25.540 2.650 ;
        RECT -25.810 2.050 -25.540 2.600 ;
        RECT -25.810 1.400 -25.650 2.050 ;
        RECT -25.400 1.400 -25.210 2.860 ;
        RECT -23.510 2.110 -23.320 3.730 ;
        RECT -23.060 2.620 -22.870 3.910 ;
        RECT -23.080 2.330 -22.850 2.620 ;
        RECT -23.990 1.700 -23.690 2.080 ;
        RECT -23.510 1.900 -23.280 2.110 ;
        RECT -23.520 1.820 -23.280 1.900 ;
        RECT -23.520 1.400 -23.290 1.820 ;
        RECT -23.060 1.400 -22.870 2.330 ;
        RECT -22.650 1.400 -22.440 4.220 ;
        RECT -21.570 2.920 -21.390 7.450 ;
        RECT -20.850 5.450 -20.590 6.240 ;
        RECT -21.630 2.580 -21.340 2.920 ;
        RECT -21.570 1.400 -21.390 2.580 ;
        RECT -20.850 2.510 -20.590 3.300 ;
        RECT -17.700 1.400 -17.470 7.450 ;
        RECT -15.410 1.400 -14.990 7.450 ;
        RECT -14.380 1.400 -13.960 7.450 ;
        RECT -11.900 1.400 -11.670 7.450 ;
        RECT -10.680 6.240 -10.450 7.450 ;
        RECT -5.680 6.770 -5.380 7.150 ;
        RECT -0.990 6.830 -0.670 7.150 ;
        RECT 1.260 6.880 1.580 7.200 ;
        RECT -1.820 6.280 -1.500 6.600 ;
        RECT -10.680 5.450 -10.420 6.240 ;
        RECT -1.040 6.180 -0.720 6.500 ;
        RECT -5.530 5.670 -5.210 5.990 ;
        RECT -2.930 5.750 -2.610 6.070 ;
        RECT -1.710 5.590 -1.500 5.700 ;
        RECT -10.680 3.300 -10.450 5.450 ;
        RECT -1.730 5.270 -1.470 5.590 ;
        RECT -1.040 5.350 -0.720 5.670 ;
        RECT -1.710 3.980 -1.500 5.270 ;
        RECT -1.730 3.690 -1.500 3.980 ;
        RECT -10.680 2.510 -10.420 3.300 ;
        RECT -5.530 2.910 -5.210 3.230 ;
        RECT -1.040 3.220 -0.720 3.540 ;
        RECT -10.680 1.400 -10.450 2.510 ;
        RECT -1.040 2.390 -0.720 2.710 ;
        RECT -5.680 1.700 -5.380 2.080 ;
        RECT -0.990 1.740 -0.670 2.060 ;
        RECT 1.220 1.690 1.540 2.010 ;
      LAYER via ;
        RECT -23.970 6.830 -23.710 7.100 ;
        RECT -24.370 5.130 -24.110 5.390 ;
        RECT -25.080 4.300 -24.820 4.560 ;
        RECT -24.380 3.440 -24.120 3.700 ;
        RECT -23.970 1.750 -23.710 2.020 ;
        RECT -5.660 6.830 -5.400 7.100 ;
        RECT -0.960 6.860 -0.700 7.120 ;
        RECT 1.290 6.910 1.550 7.170 ;
        RECT -1.790 6.310 -1.530 6.570 ;
        RECT -1.010 6.210 -0.750 6.470 ;
        RECT -5.500 5.700 -5.240 5.960 ;
        RECT -2.900 5.780 -2.640 6.040 ;
        RECT -1.730 5.300 -1.470 5.560 ;
        RECT -1.010 5.380 -0.750 5.640 ;
        RECT -1.010 3.250 -0.750 3.510 ;
        RECT -5.500 2.940 -5.240 3.200 ;
        RECT -1.010 2.420 -0.750 2.680 ;
        RECT -5.660 1.750 -5.400 2.020 ;
        RECT -0.960 1.770 -0.700 2.030 ;
        RECT 1.250 1.720 1.510 1.980 ;
      LAYER met2 ;
        RECT -23.990 6.970 -23.690 7.150 ;
        RECT -5.680 6.970 -5.380 7.150 ;
        RECT -23.990 6.950 -23.440 6.970 ;
        RECT -5.930 6.950 -5.380 6.970 ;
        RECT -0.990 7.110 -0.680 7.160 ;
        RECT 1.260 7.110 1.570 7.210 ;
        RECT -26.170 6.770 -3.200 6.950 ;
        RECT -0.990 6.880 1.570 7.110 ;
        RECT -0.990 6.830 -0.680 6.880 ;
        RECT -1.810 6.570 -1.500 6.610 ;
        RECT -1.990 6.430 -1.270 6.570 ;
        RECT -1.040 6.430 -0.730 6.510 ;
        RECT -1.990 6.320 -0.730 6.430 ;
        RECT -1.810 6.280 -0.730 6.320 ;
        RECT -1.540 6.220 -0.730 6.280 ;
        RECT -1.540 6.210 -1.270 6.220 ;
        RECT -1.040 6.180 -0.730 6.220 ;
        RECT -5.530 5.930 -5.220 6.000 ;
        RECT -2.930 5.930 -2.620 6.070 ;
        RECT -5.530 5.740 -2.620 5.930 ;
        RECT -5.530 5.710 -2.930 5.740 ;
        RECT -5.530 5.670 -5.220 5.710 ;
        RECT -1.470 5.640 -1.270 5.650 ;
        RECT -1.470 5.630 -1.250 5.640 ;
        RECT -1.040 5.630 -0.730 5.670 ;
        RECT -1.470 5.560 -0.730 5.630 ;
        RECT -1.760 5.540 -0.730 5.560 ;
        RECT -24.390 5.410 -24.080 5.430 ;
        RECT -1.810 5.420 -0.730 5.540 ;
        RECT -14.660 5.410 -6.670 5.420 ;
        RECT -24.390 5.220 -6.670 5.410 ;
        RECT -1.810 5.300 -1.250 5.420 ;
        RECT -1.040 5.340 -0.730 5.420 ;
        RECT -1.810 5.290 -1.340 5.300 ;
        RECT -24.390 5.100 -24.080 5.220 ;
        RECT -25.110 4.530 -24.790 4.560 ;
        RECT -8.070 4.540 -7.850 4.550 ;
        RECT -14.650 4.530 -7.820 4.540 ;
        RECT -25.110 4.300 -7.820 4.530 ;
        RECT -6.890 4.500 -6.670 5.220 ;
        RECT -14.650 4.290 -7.820 4.300 ;
        RECT -24.400 3.550 -24.090 3.740 ;
        RECT -14.650 3.550 -11.140 3.560 ;
        RECT -24.400 3.410 -11.140 3.550 ;
        RECT -24.370 3.370 -11.140 3.410 ;
        RECT -24.370 3.360 -14.650 3.370 ;
        RECT -11.370 2.770 -11.140 3.370 ;
        RECT -8.110 3.120 -7.820 4.290 ;
        RECT -6.920 4.460 -6.670 4.500 ;
        RECT -6.920 3.820 -6.660 4.460 ;
        RECT -6.920 3.610 -2.790 3.820 ;
        RECT -3.000 3.470 -2.790 3.610 ;
        RECT -1.040 3.470 -0.730 3.550 ;
        RECT -3.000 3.260 -0.730 3.470 ;
        RECT -5.530 3.170 -5.220 3.240 ;
        RECT -1.040 3.220 -0.730 3.260 ;
        RECT -5.530 3.120 -3.200 3.170 ;
        RECT -8.110 2.960 -3.200 3.120 ;
        RECT -8.110 2.900 -5.220 2.960 ;
        RECT -8.110 2.890 -7.820 2.900 ;
        RECT -11.370 2.620 -11.150 2.770 ;
        RECT -1.040 2.670 -0.730 2.710 ;
        RECT -7.000 2.620 -0.730 2.670 ;
        RECT -11.370 2.460 -0.730 2.620 ;
        RECT -11.370 2.400 -6.610 2.460 ;
        RECT -1.040 2.380 -0.730 2.460 ;
        RECT -23.860 2.080 -23.700 2.090 ;
        RECT -5.670 2.080 -5.510 2.090 ;
        RECT -26.170 2.070 -23.610 2.080 ;
        RECT -5.760 2.070 -3.200 2.080 ;
        RECT -26.170 1.920 -3.200 2.070 ;
        RECT -26.170 1.900 -23.610 1.920 ;
        RECT -5.760 1.900 -3.200 1.920 ;
        RECT -0.990 1.980 -0.680 2.060 ;
        RECT 1.220 1.980 1.530 2.020 ;
        RECT -23.990 1.700 -23.690 1.900 ;
        RECT -5.680 1.700 -5.380 1.900 ;
        RECT -0.990 1.750 1.720 1.980 ;
        RECT -0.990 1.730 -0.680 1.750 ;
        RECT 1.220 1.690 1.530 1.750 ;
  END
END sky130_hilas_TA2Cell_1FG_Strong

MACRO sky130_hilas_FGcharacterization01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_FGcharacterization01 ;
  ORIGIN 9.120 -2.590 ;
  SIZE 29.950 BY 6.050 ;
  PIN VTUNVARACTOR01
    USE ANALOG ;
    ANTENNADIFFAREA 0.604400 ;
    PORT
      LAYER nwell ;
        RECT -9.120 6.880 -6.900 8.570 ;
      LAYER li1 ;
        RECT -8.820 7.400 -8.590 8.090 ;
      LAYER mcon ;
        RECT -8.790 7.880 -8.620 8.050 ;
        RECT -8.790 7.430 -8.620 7.600 ;
      LAYER met1 ;
        RECT -8.840 7.350 -8.580 8.640 ;
    END
  END VTUNVARACTOR01
  PIN VARACTORCAP01
    USE ANALOG ;
    ANTENNADIFFAREA 0.859400 ;
    PORT
      LAYER nwell ;
        RECT -4.420 8.580 -1.710 8.620 ;
        RECT -4.420 6.930 -1.700 8.580 ;
      LAYER li1 ;
        RECT -4.120 7.450 -3.890 8.140 ;
      LAYER mcon ;
        RECT -4.090 7.930 -3.920 8.100 ;
        RECT -4.090 7.480 -3.920 7.650 ;
      LAYER met1 ;
        RECT -4.140 7.390 -3.870 8.640 ;
    END
  END VARACTORCAP01
  PIN OVERLAPCAP01
    USE ANALOG ;
    ANTENNADIFFAREA 0.336400 ;
    PORT
      LAYER li1 ;
        RECT 0.200 7.270 3.510 8.250 ;
      LAYER mcon ;
        RECT 1.770 8.020 1.940 8.190 ;
        RECT 1.770 7.670 1.940 7.840 ;
        RECT 1.770 7.330 1.940 7.500 ;
      LAYER met1 ;
        RECT 1.730 7.610 1.970 8.640 ;
        RECT 1.740 7.350 1.970 7.610 ;
        RECT 1.740 7.130 1.980 7.350 ;
    END
  END OVERLAPCAP01
  PIN VARACTORCAP02
    USE ANALOG ;
    ANTENNADIFFAREA 1.740800 ;
    PORT
      LAYER nwell ;
        RECT -4.420 5.590 -1.710 5.630 ;
        RECT -4.420 2.930 -1.700 5.590 ;
      LAYER li1 ;
        RECT -4.120 4.460 -3.890 5.150 ;
        RECT -4.120 3.450 -3.890 4.140 ;
      LAYER mcon ;
        RECT -4.090 4.940 -3.920 5.110 ;
        RECT -4.090 4.490 -3.920 4.660 ;
        RECT -4.090 3.930 -3.920 4.100 ;
        RECT -4.090 3.480 -3.920 3.650 ;
      LAYER met1 ;
        RECT -4.140 5.180 -3.880 5.200 ;
        RECT -4.150 2.590 -3.840 5.180 ;
    END
  END VARACTORCAP02
  PIN OVERLAPCAP02
    USE ANALOG ;
    ANTENNADIFFAREA 0.672800 ;
    PORT
      LAYER li1 ;
        RECT 0.200 4.470 3.510 5.450 ;
        RECT 0.200 2.920 3.510 3.900 ;
      LAYER mcon ;
        RECT 1.770 5.220 1.940 5.390 ;
        RECT 1.770 4.870 1.940 5.040 ;
        RECT 1.770 4.530 1.940 4.700 ;
        RECT 1.770 3.670 1.940 3.840 ;
        RECT 1.770 3.320 1.940 3.490 ;
        RECT 1.770 2.980 1.940 3.150 ;
      LAYER met1 ;
        RECT 1.730 4.810 1.970 5.450 ;
        RECT 1.740 4.550 1.970 4.810 ;
        RECT 1.740 3.900 1.980 4.550 ;
        RECT 1.730 3.260 1.980 3.900 ;
        RECT 1.740 2.590 1.980 3.260 ;
    END
  END OVERLAPCAP02
  PIN LARGECAPACITOR
    USE ANALOG ;
    ANTENNADIFFAREA 6.082200 ;
    PORT
      LAYER nwell ;
        RECT 5.430 4.000 15.120 8.600 ;
        RECT 5.430 2.610 15.720 4.000 ;
      LAYER li1 ;
        RECT 15.090 2.910 15.260 3.580 ;
      LAYER mcon ;
        RECT 15.090 3.160 15.260 3.330 ;
      LAYER met1 ;
        RECT 15.050 2.590 15.340 3.650 ;
    END
  END LARGECAPACITOR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT -5.270 6.370 -5.100 6.390 ;
        RECT -5.270 6.200 -2.210 6.370 ;
        RECT -5.270 5.550 -5.100 6.200 ;
        RECT -6.370 5.380 -5.100 5.550 ;
        RECT -5.270 2.970 -5.100 5.380 ;
        RECT 4.600 3.490 4.770 6.140 ;
        RECT 17.790 3.690 18.110 3.730 ;
        RECT 19.220 3.690 19.540 3.710 ;
        RECT 16.830 3.520 20.410 3.690 ;
        RECT -5.330 2.930 -5.010 2.970 ;
        RECT 4.590 2.950 4.770 3.490 ;
        RECT 17.790 3.500 18.120 3.520 ;
        RECT 17.790 3.470 18.110 3.500 ;
        RECT 19.220 3.480 19.550 3.520 ;
        RECT 19.220 3.450 19.540 3.480 ;
        RECT 16.930 3.080 17.250 3.120 ;
        RECT 17.640 3.090 17.960 3.130 ;
        RECT 18.380 3.090 18.700 3.130 ;
        RECT 19.080 3.090 19.400 3.130 ;
        RECT 20.010 3.090 20.330 3.130 ;
        RECT 16.930 3.070 17.260 3.080 ;
        RECT 17.640 3.070 17.970 3.090 ;
        RECT 16.930 3.020 17.970 3.070 ;
        RECT 18.380 3.020 18.710 3.090 ;
        RECT 19.080 3.020 19.410 3.090 ;
        RECT 20.010 3.020 20.340 3.090 ;
        RECT -5.330 2.740 -5.000 2.930 ;
        RECT 4.530 2.910 4.850 2.950 ;
        RECT -5.330 2.710 -5.010 2.740 ;
        RECT 4.530 2.720 4.860 2.910 ;
        RECT 16.930 2.850 20.360 3.020 ;
        RECT 16.930 2.840 17.780 2.850 ;
        RECT 4.530 2.690 4.850 2.720 ;
      LAYER mcon ;
        RECT 17.850 3.510 18.020 3.680 ;
        RECT 19.280 3.490 19.450 3.660 ;
        RECT -5.270 2.750 -5.100 2.920 ;
        RECT 4.590 2.730 4.760 2.900 ;
        RECT 16.990 2.900 17.160 3.070 ;
        RECT 17.700 2.910 17.870 3.080 ;
        RECT 18.440 2.910 18.610 3.080 ;
        RECT 19.140 2.910 19.310 3.080 ;
        RECT 20.070 2.910 20.240 3.080 ;
      LAYER met1 ;
        RECT 17.780 3.440 18.100 3.760 ;
        RECT 19.210 3.420 19.530 3.740 ;
        RECT -5.340 2.680 -5.020 3.000 ;
        RECT 4.520 2.660 4.840 2.980 ;
        RECT 16.920 2.830 17.240 3.150 ;
        RECT 17.630 2.840 17.950 3.160 ;
        RECT 18.370 2.840 18.690 3.160 ;
        RECT 19.070 2.840 19.390 3.160 ;
        RECT 20.000 2.840 20.320 3.160 ;
      LAYER via ;
        RECT 17.810 3.470 18.070 3.730 ;
        RECT 19.240 3.450 19.500 3.710 ;
        RECT -5.310 2.710 -5.050 2.970 ;
        RECT 4.550 2.690 4.810 2.950 ;
        RECT 16.950 2.860 17.210 3.120 ;
        RECT 17.660 2.870 17.920 3.130 ;
        RECT 18.400 2.870 18.660 3.130 ;
        RECT 19.100 2.870 19.360 3.130 ;
        RECT 20.030 2.870 20.290 3.130 ;
      LAYER met2 ;
        RECT 17.780 3.540 18.090 3.770 ;
        RECT 19.210 3.540 19.520 3.750 ;
        RECT 16.950 3.210 20.830 3.540 ;
        RECT 16.940 3.160 20.830 3.210 ;
        RECT 16.920 3.050 20.830 3.160 ;
        RECT -5.340 2.870 -5.030 3.010 ;
        RECT 4.520 2.870 4.830 2.990 ;
        RECT 16.920 2.870 17.940 3.050 ;
        RECT -5.340 2.840 17.940 2.870 ;
        RECT 18.370 2.840 18.680 3.050 ;
        RECT 19.070 2.840 19.380 3.050 ;
        RECT 20.000 2.840 20.310 3.050 ;
        RECT -5.340 2.680 17.920 2.840 ;
        RECT -5.310 2.660 17.920 2.680 ;
    END
  END VGND
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.150 2.590 3.850 8.580 ;
        RECT 17.990 5.090 20.730 8.590 ;
      LAYER li1 ;
        RECT 19.200 7.310 19.520 7.350 ;
        RECT 18.320 7.140 20.400 7.310 ;
        RECT 19.200 7.120 19.530 7.140 ;
        RECT 19.200 7.090 19.520 7.120 ;
        RECT 3.230 6.610 3.400 6.960 ;
        RECT 18.400 6.730 20.220 6.900 ;
        RECT 3.230 6.570 4.130 6.610 ;
        RECT 3.230 6.380 4.140 6.570 ;
        RECT 19.200 6.490 19.520 6.510 ;
        RECT 3.230 6.350 4.130 6.380 ;
        RECT 3.230 5.950 3.400 6.350 ;
        RECT 18.320 6.320 20.400 6.490 ;
        RECT 19.200 6.280 19.530 6.320 ;
        RECT 19.200 6.250 19.520 6.280 ;
      LAYER mcon ;
        RECT 18.570 7.140 18.740 7.310 ;
        RECT 19.260 7.130 19.430 7.300 ;
        RECT 19.980 7.140 20.150 7.310 ;
        RECT 18.740 6.730 18.910 6.900 ;
        RECT 19.800 6.730 19.970 6.900 ;
        RECT 3.870 6.390 4.040 6.560 ;
        RECT 18.570 6.320 18.740 6.490 ;
        RECT 19.260 6.290 19.430 6.460 ;
        RECT 19.980 6.320 20.150 6.490 ;
      LAYER met1 ;
        RECT 18.530 7.140 18.790 7.420 ;
        RECT 19.190 7.140 19.510 7.380 ;
        RECT 19.940 7.140 20.200 7.410 ;
        RECT 3.800 6.320 4.120 6.640 ;
        RECT 18.490 6.480 20.240 7.140 ;
        RECT 18.510 6.240 18.770 6.480 ;
        RECT 19.190 6.220 19.510 6.480 ;
        RECT 19.940 6.220 20.200 6.480 ;
      LAYER via ;
        RECT 18.530 7.130 18.790 7.390 ;
        RECT 19.220 7.090 19.480 7.350 ;
        RECT 19.940 7.120 20.200 7.380 ;
        RECT 18.530 6.690 18.790 6.950 ;
        RECT 19.940 6.670 20.200 6.930 ;
        RECT 3.830 6.350 4.090 6.610 ;
        RECT 18.510 6.270 18.770 6.530 ;
        RECT 19.220 6.250 19.480 6.510 ;
        RECT 19.940 6.250 20.200 6.510 ;
      LAYER met2 ;
        RECT 3.510 7.180 18.160 7.310 ;
        RECT 18.500 7.180 18.820 7.390 ;
        RECT 19.190 7.180 19.500 7.390 ;
        RECT 19.910 7.180 20.230 7.380 ;
        RECT 3.510 7.100 20.830 7.180 ;
        RECT 3.850 6.650 4.090 7.100 ;
        RECT 18.020 6.930 20.830 7.100 ;
        RECT 3.800 6.320 4.110 6.650 ;
        RECT 18.160 6.420 20.830 6.930 ;
        RECT 18.480 6.270 18.800 6.420 ;
        RECT 19.190 6.220 19.500 6.420 ;
        RECT 19.910 6.250 20.230 6.420 ;
    END
  END VINJ
  PIN OUTPUT
    USE ANALOG ;
    ANTENNADIFFAREA 0.359600 ;
    PORT
      LAYER li1 ;
        RECT 19.730 5.480 20.400 5.650 ;
        RECT 19.730 4.360 20.400 4.530 ;
      LAYER mcon ;
        RECT 19.980 5.480 20.150 5.650 ;
        RECT 19.980 4.360 20.150 4.530 ;
      LAYER met1 ;
        RECT 19.950 5.190 20.180 5.710 ;
        RECT 19.940 4.870 20.200 5.190 ;
        RECT 19.950 4.300 20.180 4.870 ;
      LAYER via ;
        RECT 19.940 4.900 20.200 5.160 ;
      LAYER met2 ;
        RECT 20.210 5.160 20.830 5.190 ;
        RECT 19.910 4.900 20.830 5.160 ;
        RECT 20.210 4.870 20.830 4.900 ;
    END
  END OUTPUT
  PIN VREF
    USE ANALOG ;
    ANTENNAGATEAREA 0.315000 ;
    PORT
      LAYER li1 ;
        RECT 17.400 6.480 17.610 6.910 ;
        RECT 17.420 6.460 17.590 6.480 ;
      LAYER met1 ;
        RECT 17.350 6.630 17.670 6.950 ;
        RECT 17.390 6.400 17.620 6.630 ;
      LAYER via ;
        RECT 17.380 6.660 17.640 6.920 ;
      LAYER met2 ;
        RECT 17.350 6.630 17.670 6.950 ;
        RECT 17.380 5.590 17.650 6.630 ;
        RECT 17.380 5.580 20.170 5.590 ;
        RECT 17.380 5.360 20.830 5.580 ;
        RECT 17.900 5.350 20.830 5.360 ;
    END
  END VREF
  PIN AMPLIFIERBIAS
    USE ANALOG ;
    ANTENNAGATEAREA 0.477400 ;
    PORT
      LAYER li1 ;
        RECT 17.920 4.910 18.090 4.940 ;
        RECT 17.760 4.880 18.090 4.910 ;
        RECT 17.750 4.690 18.090 4.880 ;
        RECT 17.760 4.650 18.090 4.690 ;
        RECT 17.920 4.610 18.090 4.650 ;
      LAYER mcon ;
        RECT 17.850 4.700 18.020 4.870 ;
      LAYER met1 ;
        RECT 17.770 4.620 18.090 4.940 ;
      LAYER via ;
        RECT 17.800 4.650 18.060 4.910 ;
      LAYER met2 ;
        RECT 17.780 4.710 18.090 4.940 ;
        RECT 17.780 4.610 20.830 4.710 ;
        RECT 17.800 4.480 20.830 4.610 ;
    END
  END AMPLIFIERBIAS
  OBS
      LAYER li1 ;
        RECT 16.860 8.200 17.530 8.370 ;
        RECT 19.160 8.160 19.330 8.470 ;
        RECT 20.560 8.170 20.730 8.470 ;
        RECT 18.320 7.990 19.330 8.160 ;
        RECT 19.730 7.990 20.730 8.170 ;
        RECT 16.860 7.410 17.530 7.580 ;
        RECT 1.830 6.680 2.000 6.720 ;
        RECT 2.510 6.690 2.680 6.720 ;
        RECT 1.760 6.640 2.080 6.680 ;
        RECT 2.450 6.650 2.770 6.690 ;
        RECT 1.760 6.450 2.090 6.640 ;
        RECT 2.450 6.460 2.780 6.650 ;
        RECT 1.760 6.420 2.080 6.450 ;
        RECT 2.450 6.430 2.770 6.460 ;
        RECT 1.830 6.390 2.000 6.420 ;
        RECT 2.510 6.390 2.680 6.430 ;
        RECT 16.860 5.980 17.530 6.150 ;
        RECT 18.320 5.480 19.000 5.650 ;
        RECT 17.830 5.360 18.020 5.420 ;
        RECT 16.850 5.190 18.020 5.360 ;
        RECT -8.010 3.730 -7.840 4.620 ;
        RECT 16.850 4.580 17.520 4.750 ;
        RECT 19.170 4.530 19.340 4.590 ;
        RECT 18.320 4.360 19.340 4.530 ;
        RECT 19.170 4.260 19.340 4.360 ;
      LAYER mcon ;
        RECT 17.110 8.200 17.280 8.370 ;
        RECT 18.570 7.990 18.740 8.160 ;
        RECT 19.980 7.990 20.150 8.160 ;
        RECT 17.110 7.410 17.280 7.580 ;
        RECT 1.820 6.460 1.990 6.630 ;
        RECT 2.510 6.470 2.680 6.640 ;
        RECT 17.110 5.980 17.280 6.150 ;
        RECT 18.570 5.480 18.740 5.650 ;
        RECT 17.840 5.220 18.010 5.390 ;
        RECT -8.010 4.420 -7.840 4.590 ;
        RECT 17.100 4.580 17.270 4.750 ;
        RECT 18.570 4.360 18.740 4.530 ;
      LAYER met1 ;
        RECT 17.070 8.400 17.330 8.490 ;
        RECT 17.050 8.170 17.340 8.400 ;
        RECT 19.930 8.240 20.190 8.440 ;
        RECT 17.810 7.930 18.840 8.240 ;
        RECT 19.870 7.930 20.250 8.240 ;
        RECT 17.000 7.480 17.390 7.610 ;
        RECT 16.970 7.190 17.390 7.480 ;
        RECT 1.750 6.390 2.070 6.710 ;
        RECT 2.440 6.400 2.760 6.720 ;
        RECT 16.970 6.250 17.200 7.190 ;
        RECT 16.970 6.180 17.330 6.250 ;
        RECT 16.970 6.070 17.390 6.180 ;
        RECT 17.000 5.950 17.390 6.070 ;
        RECT -8.040 4.640 -7.810 4.810 ;
        RECT 17.060 4.780 17.330 5.950 ;
        RECT 17.810 5.160 18.050 7.930 ;
        RECT -8.050 2.590 -7.800 4.640 ;
        RECT 17.000 4.550 17.330 4.780 ;
        RECT 18.540 4.300 18.770 5.710 ;
      LAYER via ;
        RECT 17.070 8.200 17.330 8.460 ;
        RECT 19.930 8.150 20.190 8.410 ;
        RECT 1.780 6.420 2.040 6.680 ;
        RECT 2.470 6.430 2.730 6.690 ;
      LAYER met2 ;
        RECT 17.040 8.410 17.360 8.460 ;
        RECT 17.040 8.170 20.220 8.410 ;
        RECT 19.900 8.150 20.220 8.170 ;
        RECT 1.750 6.390 2.060 6.720 ;
        RECT 2.440 6.400 2.750 6.730 ;
  END
END sky130_hilas_FGcharacterization01

MACRO sky130_hilas_m22m4
  CLASS BLOCK ;
  FOREIGN sky130_hilas_m22m4 ;
  ORIGIN 0.360 0.360 ;
  SIZE 0.790 BY 0.750 ;
  OBS
      LAYER met2 ;
        RECT -0.140 -0.160 0.230 0.240 ;
      LAYER via2 ;
        RECT -0.090 -0.100 0.190 0.180 ;
      LAYER met3 ;
        RECT -0.360 -0.360 0.430 0.390 ;
      LAYER via3 ;
        RECT -0.170 -0.210 0.260 0.270 ;
      LAYER met4 ;
        RECT -0.270 -0.300 0.390 0.360 ;
  END
END sky130_hilas_m22m4

MACRO sky130_hilas_DAC6bit01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_DAC6bit01 ;
  ORIGIN -0.230 0.060 ;
  SIZE 33.400 BY 13.680 ;
  OBS
      LAYER nwell ;
        RECT 18.990 13.360 20.600 13.620 ;
        RECT 18.860 7.970 20.600 13.360 ;
        RECT 18.860 7.710 20.470 7.970 ;
        RECT 0.600 -0.030 16.700 5.620 ;
        RECT 17.420 -0.030 19.030 5.620 ;
        RECT 20.750 4.900 30.850 4.970 ;
        RECT 31.910 -0.030 33.520 5.620 ;
      LAYER li1 ;
        RECT 19.370 12.140 19.540 12.400 ;
        RECT 20.050 12.140 20.220 12.400 ;
        RECT 19.240 12.070 19.540 12.140 ;
        RECT 19.920 12.070 20.220 12.140 ;
        RECT 19.240 11.810 19.410 12.070 ;
        RECT 19.920 11.810 20.090 12.070 ;
        RECT 19.370 11.180 19.540 11.440 ;
        RECT 20.050 11.180 20.220 11.440 ;
        RECT 19.240 11.110 19.540 11.180 ;
        RECT 19.920 11.110 20.220 11.180 ;
        RECT 19.240 10.850 19.410 11.110 ;
        RECT 19.920 10.850 20.090 11.110 ;
        RECT 19.370 10.220 19.540 10.480 ;
        RECT 20.050 10.220 20.220 10.480 ;
        RECT 19.240 10.150 19.540 10.220 ;
        RECT 19.920 10.150 20.220 10.220 ;
        RECT 19.240 9.890 19.410 10.150 ;
        RECT 19.920 9.890 20.090 10.150 ;
        RECT 19.370 9.260 19.540 9.520 ;
        RECT 20.050 9.260 20.220 9.520 ;
        RECT 19.240 9.190 19.540 9.260 ;
        RECT 19.920 9.190 20.220 9.260 ;
        RECT 19.240 8.930 19.410 9.190 ;
        RECT 19.920 8.930 20.090 9.190 ;
        RECT 0.630 5.410 0.840 5.840 ;
        RECT 2.220 5.420 2.430 5.850 ;
        RECT 3.620 5.440 4.050 5.460 ;
        RECT 0.650 5.390 0.820 5.410 ;
        RECT 2.240 5.400 2.410 5.420 ;
        RECT 3.600 5.270 4.050 5.440 ;
        RECT 5.420 5.410 5.630 5.840 ;
        RECT 7.030 5.410 7.240 5.840 ;
        RECT 8.650 5.410 8.860 5.840 ;
        RECT 10.260 5.420 10.470 5.850 ;
        RECT 11.870 5.420 12.080 5.850 ;
        RECT 13.180 5.740 13.390 5.750 ;
        RECT 13.070 5.700 13.390 5.740 ;
        RECT 13.740 5.700 14.060 5.740 ;
        RECT 13.070 5.510 13.400 5.700 ;
        RECT 13.740 5.510 14.070 5.700 ;
        RECT 13.070 5.480 13.390 5.510 ;
        RECT 13.740 5.480 14.060 5.510 ;
        RECT 5.440 5.390 5.610 5.410 ;
        RECT 7.050 5.390 7.220 5.410 ;
        RECT 8.670 5.390 8.840 5.410 ;
        RECT 10.280 5.400 10.450 5.420 ;
        RECT 11.890 5.400 12.060 5.420 ;
        RECT 3.620 5.250 4.050 5.270 ;
        RECT 4.210 4.970 4.380 4.980 ;
        RECT 13.180 4.970 13.390 5.480 ;
        RECT 13.850 4.970 14.020 5.480 ;
        RECT 17.450 5.410 17.660 5.840 ;
        RECT 19.040 5.420 19.250 5.850 ;
        RECT 20.440 5.440 20.870 5.460 ;
        RECT 17.470 5.390 17.640 5.410 ;
        RECT 19.060 5.400 19.230 5.420 ;
        RECT 20.420 5.270 20.870 5.440 ;
        RECT 22.240 5.410 22.450 5.840 ;
        RECT 23.850 5.410 24.060 5.840 ;
        RECT 25.470 5.410 25.680 5.840 ;
        RECT 27.080 5.420 27.290 5.850 ;
        RECT 28.690 5.420 28.900 5.850 ;
        RECT 30.000 5.740 30.210 5.750 ;
        RECT 29.890 5.700 30.210 5.740 ;
        RECT 30.560 5.700 30.880 5.740 ;
        RECT 29.890 5.510 30.220 5.700 ;
        RECT 30.560 5.510 30.890 5.700 ;
        RECT 29.890 5.480 30.210 5.510 ;
        RECT 30.560 5.480 30.880 5.510 ;
        RECT 22.260 5.390 22.430 5.410 ;
        RECT 23.870 5.390 24.040 5.410 ;
        RECT 25.490 5.390 25.660 5.410 ;
        RECT 27.100 5.400 27.270 5.420 ;
        RECT 28.710 5.400 28.880 5.420 ;
        RECT 20.440 5.250 20.870 5.270 ;
        RECT 21.030 4.970 21.200 4.980 ;
        RECT 30.000 4.970 30.210 5.480 ;
        RECT 30.670 4.970 30.840 5.480 ;
        RECT 2.600 4.740 14.030 4.970 ;
        RECT 0.490 4.100 0.700 4.530 ;
        RECT 2.600 4.400 2.770 4.740 ;
        RECT 0.510 4.080 0.680 4.100 ;
        RECT 2.590 4.070 2.770 4.400 ;
        RECT 0.550 3.150 0.760 3.580 ;
        RECT 2.600 3.440 2.770 4.070 ;
        RECT 0.570 3.130 0.740 3.150 ;
        RECT 2.590 3.110 2.770 3.440 ;
        RECT 0.550 2.210 0.760 2.640 ;
        RECT 2.600 2.480 2.770 3.110 ;
        RECT 0.570 2.190 0.740 2.210 ;
        RECT 2.590 2.150 2.770 2.480 ;
        RECT 2.600 1.520 2.770 2.150 ;
        RECT 2.590 1.190 2.770 1.520 ;
        RECT 2.600 1.180 2.770 1.190 ;
        RECT 3.260 4.400 3.430 4.410 ;
        RECT 4.210 4.400 4.380 4.740 ;
        RECT 5.800 4.400 5.970 4.740 ;
        RECT 3.260 4.070 3.440 4.400 ;
        RECT 4.200 4.070 4.380 4.400 ;
        RECT 4.880 4.370 5.050 4.400 ;
        RECT 4.880 4.070 5.060 4.370 ;
        RECT 3.260 3.440 3.430 4.070 ;
        RECT 4.210 3.440 4.380 4.070 ;
        RECT 4.890 3.440 5.060 4.070 ;
        RECT 3.260 3.110 3.440 3.440 ;
        RECT 4.200 3.110 4.380 3.440 ;
        RECT 4.880 3.110 5.060 3.440 ;
        RECT 3.260 2.480 3.430 3.110 ;
        RECT 4.210 2.480 4.380 3.110 ;
        RECT 4.890 2.480 5.060 3.110 ;
        RECT 3.260 2.150 3.440 2.480 ;
        RECT 4.200 2.150 4.380 2.480 ;
        RECT 4.880 2.150 5.060 2.480 ;
        RECT 3.260 1.520 3.430 2.150 ;
        RECT 4.210 1.520 4.380 2.150 ;
        RECT 4.890 1.520 5.060 2.150 ;
        RECT 3.260 1.190 3.440 1.520 ;
        RECT 4.200 1.190 4.380 1.520 ;
        RECT 4.880 1.190 5.060 1.520 ;
        RECT 3.260 0.200 3.430 1.190 ;
        RECT 4.210 1.180 4.380 1.190 ;
        RECT 4.890 0.200 5.060 1.190 ;
        RECT 5.800 4.070 5.980 4.400 ;
        RECT 5.800 3.440 5.970 4.070 ;
        RECT 5.800 3.110 5.980 3.440 ;
        RECT 5.800 2.480 5.970 3.110 ;
        RECT 5.800 2.150 5.980 2.480 ;
        RECT 5.800 1.520 5.970 2.150 ;
        RECT 5.800 1.190 5.980 1.520 ;
        RECT 5.800 1.180 5.970 1.190 ;
        RECT 6.490 0.200 6.660 4.450 ;
        RECT 6.970 3.160 7.180 3.590 ;
        RECT 6.990 3.140 7.160 3.160 ;
        RECT 7.420 1.180 7.590 4.740 ;
        RECT 9.040 4.400 9.210 4.740 ;
        RECT 8.100 4.070 8.280 4.400 ;
        RECT 9.030 4.070 9.210 4.400 ;
        RECT 8.110 3.440 8.280 4.070 ;
        RECT 9.040 3.440 9.210 4.070 ;
        RECT 8.100 3.110 8.280 3.440 ;
        RECT 9.030 3.110 9.210 3.440 ;
        RECT 8.110 2.480 8.280 3.110 ;
        RECT 8.500 2.680 8.670 2.700 ;
        RECT 8.100 2.150 8.280 2.480 ;
        RECT 8.480 2.250 8.690 2.680 ;
        RECT 8.110 1.520 8.280 2.150 ;
        RECT 9.040 1.520 9.210 3.110 ;
        RECT 8.100 1.190 8.280 1.520 ;
        RECT 9.030 1.200 9.210 1.520 ;
        RECT 9.030 1.190 9.200 1.200 ;
        RECT 8.110 0.200 8.280 1.190 ;
        RECT 9.710 0.200 9.880 4.450 ;
        RECT 10.220 1.250 10.430 1.680 ;
        RECT 10.240 1.230 10.410 1.250 ;
        RECT 10.640 1.190 10.810 4.740 ;
        RECT 11.330 4.400 11.500 4.450 ;
        RECT 11.320 4.070 11.500 4.400 ;
        RECT 11.330 3.440 11.500 4.070 ;
        RECT 11.320 3.110 11.500 3.440 ;
        RECT 11.330 2.480 11.500 3.110 ;
        RECT 11.320 2.150 11.500 2.480 ;
        RECT 11.330 1.520 11.500 2.150 ;
        RECT 11.320 1.190 11.500 1.520 ;
        RECT 12.250 1.190 12.420 4.740 ;
        RECT 11.330 0.200 11.500 1.190 ;
        RECT 12.930 0.200 13.100 4.430 ;
        RECT 13.860 1.170 14.030 4.740 ;
        RECT 19.420 4.740 30.850 4.970 ;
        RECT 14.540 0.200 14.710 4.610 ;
        RECT 17.310 4.100 17.520 4.530 ;
        RECT 17.330 4.080 17.500 4.100 ;
        RECT 17.370 3.150 17.580 3.580 ;
        RECT 17.390 3.130 17.560 3.150 ;
        RECT 17.370 2.210 17.580 2.640 ;
        RECT 17.390 2.190 17.560 2.210 ;
        RECT 19.420 1.180 19.590 4.740 ;
        RECT 20.080 0.200 20.250 4.410 ;
        RECT 21.030 1.180 21.200 4.740 ;
        RECT 21.710 0.200 21.880 4.370 ;
        RECT 22.620 1.180 22.790 4.740 ;
        RECT 23.310 0.200 23.480 4.450 ;
        RECT 24.240 1.180 24.410 4.740 ;
        RECT 24.930 0.200 25.100 4.400 ;
        RECT 25.860 1.200 26.030 4.740 ;
        RECT 26.530 0.200 26.700 4.450 ;
        RECT 27.460 1.210 27.630 4.740 ;
        RECT 28.150 0.200 28.320 4.450 ;
        RECT 29.070 1.200 29.240 4.740 ;
        RECT 29.750 0.200 29.920 4.430 ;
        RECT 30.680 1.170 30.850 4.740 ;
        RECT 31.360 0.200 31.530 4.610 ;
        RECT 3.260 -0.030 3.450 0.200 ;
        RECT 4.880 -0.030 5.070 0.200 ;
        RECT 6.480 -0.030 6.670 0.200 ;
        RECT 8.100 -0.030 8.290 0.200 ;
        RECT 9.700 -0.030 9.890 0.200 ;
        RECT 11.320 -0.030 11.510 0.200 ;
        RECT 12.920 -0.030 13.110 0.200 ;
        RECT 14.530 -0.030 14.720 0.200 ;
        RECT 20.080 -0.030 20.270 0.200 ;
        RECT 21.700 -0.030 21.890 0.200 ;
        RECT 23.300 -0.030 23.490 0.200 ;
        RECT 24.920 -0.030 25.110 0.200 ;
        RECT 26.520 -0.030 26.710 0.200 ;
        RECT 28.140 -0.030 28.330 0.200 ;
        RECT 29.740 -0.030 29.930 0.200 ;
        RECT 31.350 -0.030 31.540 0.200 ;
        RECT 3.260 -0.050 3.430 -0.030 ;
        RECT 4.890 -0.050 5.060 -0.030 ;
        RECT 6.490 -0.050 6.660 -0.030 ;
        RECT 8.110 -0.050 8.280 -0.030 ;
        RECT 9.710 -0.050 9.880 -0.030 ;
        RECT 11.330 -0.050 11.500 -0.030 ;
        RECT 12.930 -0.050 13.100 -0.030 ;
        RECT 14.540 -0.050 14.710 -0.030 ;
        RECT 20.080 -0.050 20.250 -0.030 ;
        RECT 21.710 -0.050 21.880 -0.030 ;
        RECT 23.310 -0.050 23.480 -0.030 ;
        RECT 24.930 -0.050 25.100 -0.030 ;
        RECT 26.530 -0.050 26.700 -0.030 ;
        RECT 28.150 -0.050 28.320 -0.030 ;
        RECT 29.750 -0.050 29.920 -0.030 ;
        RECT 31.360 -0.050 31.530 -0.030 ;
      LAYER mcon ;
        RECT 13.130 5.520 13.300 5.690 ;
        RECT 13.800 5.520 13.970 5.690 ;
        RECT 29.950 5.520 30.120 5.690 ;
        RECT 30.620 5.520 30.790 5.690 ;
        RECT 8.500 2.530 8.670 2.700 ;
        RECT 3.270 0.000 3.440 0.170 ;
        RECT 4.890 0.000 5.060 0.170 ;
        RECT 6.490 0.000 6.660 0.170 ;
        RECT 8.110 0.000 8.280 0.170 ;
        RECT 9.710 0.000 9.880 0.170 ;
        RECT 11.330 0.000 11.500 0.170 ;
        RECT 12.930 0.000 13.100 0.170 ;
        RECT 14.540 0.000 14.710 0.170 ;
        RECT 20.090 0.000 20.260 0.170 ;
        RECT 21.710 0.000 21.880 0.170 ;
        RECT 23.310 0.000 23.480 0.170 ;
        RECT 24.930 0.000 25.100 0.170 ;
        RECT 26.530 0.000 26.700 0.170 ;
        RECT 28.150 0.000 28.320 0.170 ;
        RECT 29.750 0.000 29.920 0.170 ;
        RECT 31.360 0.000 31.530 0.170 ;
      LAYER met1 ;
        RECT 0.580 5.560 0.900 5.880 ;
        RECT 2.170 5.570 2.490 5.890 ;
        RECT 0.620 5.330 0.850 5.560 ;
        RECT 2.210 5.340 2.440 5.570 ;
        RECT 5.370 5.560 5.690 5.880 ;
        RECT 6.980 5.560 7.300 5.880 ;
        RECT 8.600 5.560 8.920 5.880 ;
        RECT 10.210 5.570 10.530 5.890 ;
        RECT 11.820 5.570 12.140 5.890 ;
        RECT 3.770 5.470 4.090 5.510 ;
        RECT 3.540 5.240 4.090 5.470 ;
        RECT 5.410 5.330 5.640 5.560 ;
        RECT 7.020 5.330 7.250 5.560 ;
        RECT 8.640 5.330 8.870 5.560 ;
        RECT 10.250 5.340 10.480 5.570 ;
        RECT 11.860 5.340 12.090 5.570 ;
        RECT 13.060 5.450 13.380 5.770 ;
        RECT 13.730 5.450 14.050 5.770 ;
        RECT 17.400 5.560 17.720 5.880 ;
        RECT 18.990 5.570 19.310 5.890 ;
        RECT 17.440 5.330 17.670 5.560 ;
        RECT 19.030 5.340 19.260 5.570 ;
        RECT 22.190 5.560 22.510 5.880 ;
        RECT 23.800 5.560 24.120 5.880 ;
        RECT 25.420 5.560 25.740 5.880 ;
        RECT 27.030 5.570 27.350 5.890 ;
        RECT 28.640 5.570 28.960 5.890 ;
        RECT 20.590 5.470 20.910 5.510 ;
        RECT 20.360 5.240 20.910 5.470 ;
        RECT 22.230 5.330 22.460 5.560 ;
        RECT 23.840 5.330 24.070 5.560 ;
        RECT 25.460 5.330 25.690 5.560 ;
        RECT 27.070 5.340 27.300 5.570 ;
        RECT 28.680 5.340 28.910 5.570 ;
        RECT 29.880 5.450 30.200 5.770 ;
        RECT 30.550 5.450 30.870 5.770 ;
        RECT 3.770 5.190 4.090 5.240 ;
        RECT 20.590 5.190 20.910 5.240 ;
        RECT 0.440 4.250 0.760 4.570 ;
        RECT 17.260 4.250 17.580 4.570 ;
        RECT 0.480 4.020 0.710 4.250 ;
        RECT 17.300 4.020 17.530 4.250 ;
        RECT 0.500 3.300 0.820 3.620 ;
        RECT 6.970 3.500 10.420 3.670 ;
        RECT 6.970 3.370 7.190 3.500 ;
        RECT 0.540 3.070 0.770 3.300 ;
        RECT 6.960 3.080 7.190 3.370 ;
        RECT 0.500 2.360 0.820 2.680 ;
        RECT 8.470 2.470 8.700 2.760 ;
        RECT 0.540 2.130 0.770 2.360 ;
        RECT 8.480 2.250 8.700 2.470 ;
        RECT 8.520 0.990 8.700 2.250 ;
        RECT 10.220 1.680 10.420 3.500 ;
        RECT 17.320 3.300 17.640 3.620 ;
        RECT 23.790 3.500 27.240 3.670 ;
        RECT 17.360 3.070 17.590 3.300 ;
        RECT 17.320 2.360 17.640 2.680 ;
        RECT 17.360 2.130 17.590 2.360 ;
        RECT 10.220 1.460 10.440 1.680 ;
        RECT 10.210 1.170 10.440 1.460 ;
        RECT 25.340 0.990 25.520 2.510 ;
        RECT 27.040 1.660 27.240 3.500 ;
        RECT 8.520 0.670 8.780 0.990 ;
        RECT 25.340 0.670 25.600 0.990 ;
        RECT 3.240 0.180 3.470 0.230 ;
        RECT 4.860 0.180 5.090 0.230 ;
        RECT 6.460 0.180 6.690 0.230 ;
        RECT 8.080 0.180 8.310 0.230 ;
        RECT 9.680 0.180 9.910 0.230 ;
        RECT 11.300 0.180 11.530 0.230 ;
        RECT 12.900 0.180 13.130 0.230 ;
        RECT 14.510 0.180 14.740 0.230 ;
        RECT 20.060 0.180 20.290 0.230 ;
        RECT 21.680 0.180 21.910 0.230 ;
        RECT 23.280 0.180 23.510 0.230 ;
        RECT 24.900 0.180 25.130 0.230 ;
        RECT 26.500 0.180 26.730 0.230 ;
        RECT 28.120 0.180 28.350 0.230 ;
        RECT 29.720 0.180 29.950 0.230 ;
        RECT 31.330 0.180 31.560 0.230 ;
        RECT 3.240 -0.050 16.810 0.180 ;
        RECT 20.060 -0.050 33.530 0.180 ;
        RECT 3.240 -0.060 3.470 -0.050 ;
        RECT 4.860 -0.060 5.090 -0.050 ;
        RECT 6.460 -0.060 6.690 -0.050 ;
        RECT 8.080 -0.060 8.310 -0.050 ;
        RECT 9.680 -0.060 9.910 -0.050 ;
        RECT 11.300 -0.060 11.530 -0.050 ;
        RECT 12.900 -0.060 13.130 -0.050 ;
        RECT 14.510 -0.060 14.740 -0.050 ;
        RECT 20.060 -0.060 20.290 -0.050 ;
        RECT 21.680 -0.060 21.910 -0.050 ;
        RECT 23.280 -0.060 23.510 -0.050 ;
        RECT 24.900 -0.060 25.130 -0.050 ;
        RECT 26.500 -0.060 26.730 -0.050 ;
        RECT 28.120 -0.060 28.350 -0.050 ;
        RECT 29.720 -0.060 29.950 -0.050 ;
        RECT 31.330 -0.060 31.560 -0.050 ;
      LAYER via ;
        RECT 0.610 5.590 0.870 5.850 ;
        RECT 2.200 5.600 2.460 5.860 ;
        RECT 5.400 5.590 5.660 5.850 ;
        RECT 7.010 5.590 7.270 5.850 ;
        RECT 8.630 5.590 8.890 5.850 ;
        RECT 10.240 5.600 10.500 5.860 ;
        RECT 11.850 5.600 12.110 5.860 ;
        RECT 3.800 5.220 4.060 5.480 ;
        RECT 13.090 5.480 13.350 5.740 ;
        RECT 13.760 5.480 14.020 5.740 ;
        RECT 17.430 5.590 17.690 5.850 ;
        RECT 19.020 5.600 19.280 5.860 ;
        RECT 22.220 5.590 22.480 5.850 ;
        RECT 23.830 5.590 24.090 5.850 ;
        RECT 25.450 5.590 25.710 5.850 ;
        RECT 27.060 5.600 27.320 5.860 ;
        RECT 28.670 5.600 28.930 5.860 ;
        RECT 20.620 5.220 20.880 5.480 ;
        RECT 29.910 5.480 30.170 5.740 ;
        RECT 30.580 5.480 30.840 5.740 ;
        RECT 0.470 4.280 0.730 4.540 ;
        RECT 17.290 4.280 17.550 4.540 ;
        RECT 0.530 3.330 0.790 3.590 ;
        RECT 0.530 2.390 0.790 2.650 ;
        RECT 17.350 3.330 17.610 3.590 ;
        RECT 17.350 2.390 17.610 2.650 ;
        RECT 8.520 0.700 8.780 0.960 ;
        RECT 25.340 0.700 25.600 0.960 ;
      LAYER met2 ;
        RECT 0.230 5.880 7.280 5.910 ;
        RECT 0.230 5.720 7.300 5.880 ;
        RECT 0.230 5.700 0.380 5.720 ;
        RECT 0.580 5.560 0.900 5.720 ;
        RECT 2.170 5.570 2.490 5.720 ;
        RECT 5.370 5.560 5.690 5.720 ;
        RECT 6.980 5.560 7.300 5.720 ;
        RECT 8.600 5.560 8.920 5.880 ;
        RECT 10.210 5.590 10.530 5.890 ;
        RECT 10.210 5.570 10.540 5.590 ;
        RECT 11.820 5.570 12.140 5.890 ;
        RECT 12.940 5.630 14.100 5.910 ;
        RECT 17.410 5.880 24.100 5.910 ;
        RECT 3.770 5.360 4.090 5.510 ;
        RECT 3.710 5.190 4.090 5.360 ;
        RECT 0.230 4.900 2.290 4.960 ;
        RECT 3.710 4.900 3.930 5.190 ;
        RECT 8.630 4.910 8.880 5.560 ;
        RECT 8.630 4.900 8.910 4.910 ;
        RECT 0.230 4.750 8.910 4.900 ;
        RECT 0.490 4.570 0.690 4.750 ;
        RECT 2.130 4.600 8.910 4.750 ;
        RECT 0.440 4.250 0.760 4.570 ;
        RECT 0.500 3.300 0.820 3.620 ;
        RECT 10.340 3.030 10.540 5.570 ;
        RECT 0.230 2.820 10.540 3.030 ;
        RECT 0.500 2.360 0.820 2.680 ;
        RECT 11.940 2.050 12.090 5.570 ;
        RECT 13.060 5.450 13.370 5.630 ;
        RECT 13.690 5.620 14.100 5.630 ;
        RECT 17.400 5.720 24.120 5.880 ;
        RECT 13.730 5.450 14.040 5.620 ;
        RECT 17.400 5.560 17.720 5.720 ;
        RECT 18.990 5.570 19.310 5.720 ;
        RECT 22.190 5.560 22.510 5.720 ;
        RECT 23.800 5.560 24.120 5.720 ;
        RECT 25.420 5.560 25.740 5.880 ;
        RECT 27.030 5.590 27.350 5.890 ;
        RECT 27.030 5.570 27.360 5.590 ;
        RECT 28.640 5.570 28.960 5.890 ;
        RECT 29.760 5.630 30.920 5.910 ;
        RECT 20.590 5.360 20.910 5.510 ;
        RECT 20.530 5.190 20.910 5.360 ;
        RECT 17.410 4.900 19.110 4.960 ;
        RECT 20.530 4.900 20.750 5.190 ;
        RECT 25.450 4.910 25.700 5.560 ;
        RECT 25.450 4.900 25.730 4.910 ;
        RECT 17.410 4.750 25.730 4.900 ;
        RECT 17.410 4.570 17.510 4.750 ;
        RECT 18.950 4.600 25.730 4.750 ;
        RECT 17.260 4.250 17.580 4.570 ;
        RECT 17.320 3.300 17.640 3.620 ;
        RECT 27.160 3.030 27.360 5.570 ;
        RECT 17.410 2.820 27.360 3.030 ;
        RECT 17.320 2.360 17.640 2.680 ;
        RECT 28.760 2.050 28.910 5.570 ;
        RECT 29.880 5.450 30.190 5.630 ;
        RECT 30.510 5.620 30.920 5.630 ;
        RECT 30.550 5.450 30.860 5.620 ;
        RECT 0.230 1.850 12.100 2.050 ;
        RECT 17.410 1.850 28.920 2.050 ;
        RECT 8.490 0.930 8.810 0.960 ;
        RECT 25.310 0.930 25.630 0.960 ;
        RECT 0.230 0.730 8.810 0.930 ;
        RECT 17.410 0.730 25.630 0.930 ;
        RECT 8.490 0.700 8.810 0.730 ;
        RECT 25.310 0.700 25.630 0.730 ;
  END
END sky130_hilas_DAC6bit01

MACRO sky130_hilas_swc4x2cellOverlap
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc4x2cellOverlap ;
  ORIGIN 10.010 -7.280 ;
  SIZE 17.980 BY 6.050 ;
  PIN VERT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.372000 ;
    PORT
      LAYER li1 ;
        RECT -8.880 12.060 -8.680 12.630 ;
        RECT -8.880 10.990 -8.680 11.560 ;
        RECT -8.880 9.050 -8.680 9.620 ;
        RECT -8.880 7.990 -8.680 8.560 ;
      LAYER mcon ;
        RECT -8.860 12.420 -8.690 12.590 ;
        RECT -8.860 11.030 -8.690 11.200 ;
        RECT -8.860 9.410 -8.690 9.580 ;
        RECT -8.860 8.030 -8.690 8.200 ;
      LAYER met1 ;
        RECT -8.840 12.650 -8.680 13.330 ;
        RECT -8.880 12.630 -8.680 12.650 ;
        RECT -8.890 12.390 -8.660 12.630 ;
        RECT -8.880 12.170 -8.680 12.390 ;
        RECT -8.840 11.450 -8.680 12.170 ;
        RECT -8.880 11.230 -8.680 11.450 ;
        RECT -8.890 10.990 -8.660 11.230 ;
        RECT -8.880 10.970 -8.680 10.990 ;
        RECT -8.840 9.640 -8.680 10.970 ;
        RECT -8.880 9.620 -8.680 9.640 ;
        RECT -8.890 9.380 -8.660 9.620 ;
        RECT -8.880 9.160 -8.680 9.380 ;
        RECT -8.840 8.450 -8.680 9.160 ;
        RECT -8.880 8.230 -8.680 8.450 ;
        RECT -8.890 7.990 -8.660 8.230 ;
        RECT -8.880 7.970 -8.680 7.990 ;
        RECT -8.840 7.290 -8.680 7.970 ;
    END
  END VERT1
  PIN HORIZ1
    USE ANALOG ;
    ANTENNADIFFAREA 0.174000 ;
    PORT
      LAYER li1 ;
        RECT -7.870 12.340 -7.550 12.380 ;
        RECT -7.880 12.300 -7.550 12.340 ;
        RECT -8.130 12.130 -7.550 12.300 ;
        RECT -7.870 12.120 -7.550 12.130 ;
        RECT 5.500 12.340 5.820 12.380 ;
        RECT 5.500 12.300 5.830 12.340 ;
        RECT 5.500 12.130 6.080 12.300 ;
        RECT 5.500 12.120 5.820 12.130 ;
      LAYER mcon ;
        RECT -7.780 12.160 -7.610 12.330 ;
        RECT 5.560 12.160 5.730 12.330 ;
      LAYER met1 ;
        RECT -7.860 12.090 -7.540 12.410 ;
        RECT 5.490 12.090 5.810 12.410 ;
      LAYER via ;
        RECT -7.830 12.120 -7.570 12.380 ;
        RECT 5.520 12.120 5.780 12.380 ;
      LAYER met2 ;
        RECT -7.850 12.400 -7.540 12.420 ;
        RECT 5.490 12.400 5.800 12.420 ;
        RECT -10.010 12.220 7.970 12.400 ;
        RECT -7.850 12.090 -7.540 12.220 ;
        RECT 5.490 12.090 5.800 12.220 ;
    END
  END HORIZ1
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.198400 ;
    PORT
      LAYER li1 ;
        RECT -7.870 12.920 -7.550 12.930 ;
        RECT -8.130 12.750 -7.550 12.920 ;
        RECT -7.880 12.700 -7.550 12.750 ;
        RECT -7.870 12.670 -7.550 12.700 ;
        RECT 5.500 12.920 5.820 12.930 ;
        RECT 5.500 12.750 6.080 12.920 ;
        RECT 5.500 12.700 5.830 12.750 ;
        RECT 5.500 12.670 5.820 12.700 ;
      LAYER mcon ;
        RECT -7.780 12.710 -7.610 12.880 ;
        RECT 5.560 12.710 5.730 12.880 ;
      LAYER met1 ;
        RECT -7.860 12.640 -7.540 12.960 ;
        RECT 5.490 12.640 5.810 12.960 ;
      LAYER via ;
        RECT -7.830 12.670 -7.570 12.930 ;
        RECT 5.520 12.670 5.780 12.930 ;
      LAYER met2 ;
        RECT -7.850 12.830 -7.540 12.970 ;
        RECT 5.490 12.830 5.800 12.970 ;
        RECT -10.010 12.650 7.960 12.830 ;
        RECT -7.850 12.640 -7.540 12.650 ;
        RECT 5.490 12.640 5.800 12.650 ;
    END
  END DRAIN1
  PIN HORIZ2
    USE ANALOG ;
    ANTENNADIFFAREA 0.174000 ;
    PORT
      LAYER li1 ;
        RECT -7.870 11.490 -7.550 11.500 ;
        RECT -8.130 11.320 -7.550 11.490 ;
        RECT -7.880 11.280 -7.550 11.320 ;
        RECT -7.870 11.240 -7.550 11.280 ;
        RECT 5.500 11.490 5.820 11.500 ;
        RECT 5.500 11.320 6.080 11.490 ;
        RECT 5.500 11.280 5.830 11.320 ;
        RECT 5.500 11.240 5.820 11.280 ;
      LAYER mcon ;
        RECT -7.780 11.290 -7.610 11.460 ;
        RECT 5.560 11.290 5.730 11.460 ;
      LAYER met1 ;
        RECT -7.860 11.210 -7.540 11.530 ;
        RECT 5.490 11.210 5.810 11.530 ;
      LAYER via ;
        RECT -7.830 11.240 -7.570 11.500 ;
        RECT 5.520 11.240 5.780 11.500 ;
      LAYER met2 ;
        RECT -7.850 11.400 -7.540 11.530 ;
        RECT 5.490 11.400 5.800 11.530 ;
        RECT -10.010 11.220 7.970 11.400 ;
        RECT -7.850 11.200 -7.540 11.220 ;
        RECT 5.490 11.200 5.800 11.220 ;
    END
  END HORIZ2
  PIN DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.198400 ;
    PORT
      LAYER li1 ;
        RECT -7.870 10.920 -7.550 10.950 ;
        RECT -7.880 10.870 -7.550 10.920 ;
        RECT -8.130 10.700 -7.550 10.870 ;
        RECT -7.870 10.690 -7.550 10.700 ;
        RECT 5.500 10.920 5.820 10.950 ;
        RECT 5.500 10.870 5.830 10.920 ;
        RECT 5.500 10.700 6.080 10.870 ;
        RECT 5.500 10.690 5.820 10.700 ;
      LAYER mcon ;
        RECT -7.780 10.740 -7.610 10.910 ;
        RECT 5.560 10.740 5.730 10.910 ;
      LAYER met1 ;
        RECT -7.860 10.660 -7.540 10.980 ;
        RECT 5.490 10.660 5.810 10.980 ;
      LAYER via ;
        RECT -7.830 10.690 -7.570 10.950 ;
        RECT 5.520 10.690 5.780 10.950 ;
      LAYER met2 ;
        RECT -7.850 10.970 -7.540 10.980 ;
        RECT 5.490 10.970 5.800 10.980 ;
        RECT -10.010 10.790 7.970 10.970 ;
        RECT -7.850 10.650 -7.540 10.790 ;
        RECT 5.490 10.650 5.800 10.790 ;
    END
  END DRAIN2
  PIN DRAIN3
    USE ANALOG ;
    ANTENNADIFFAREA 0.198400 ;
    PORT
      LAYER li1 ;
        RECT -7.870 9.910 -7.550 9.920 ;
        RECT -8.130 9.740 -7.550 9.910 ;
        RECT -7.880 9.690 -7.550 9.740 ;
        RECT -7.870 9.660 -7.550 9.690 ;
        RECT 5.500 9.910 5.820 9.920 ;
        RECT 5.500 9.740 6.080 9.910 ;
        RECT 5.500 9.690 5.830 9.740 ;
        RECT 5.500 9.660 5.820 9.690 ;
      LAYER mcon ;
        RECT -7.780 9.700 -7.610 9.870 ;
        RECT 5.560 9.700 5.730 9.870 ;
      LAYER met1 ;
        RECT -7.860 9.630 -7.540 9.950 ;
        RECT 5.490 9.630 5.810 9.950 ;
      LAYER via ;
        RECT -7.830 9.660 -7.570 9.920 ;
        RECT 5.520 9.660 5.780 9.920 ;
      LAYER met2 ;
        RECT -7.850 9.820 -7.540 9.960 ;
        RECT -10.010 9.810 -7.540 9.820 ;
        RECT 5.490 9.820 5.800 9.960 ;
        RECT 5.490 9.810 7.960 9.820 ;
        RECT -10.010 9.640 7.960 9.810 ;
        RECT -7.850 9.630 -7.540 9.640 ;
        RECT 5.490 9.630 5.800 9.640 ;
    END
  END DRAIN3
  PIN HORIZ3
    USE ANALOG ;
    ANTENNADIFFAREA 0.174000 ;
    PORT
      LAYER li1 ;
        RECT -7.870 9.330 -7.550 9.370 ;
        RECT -7.880 9.290 -7.550 9.330 ;
        RECT -8.130 9.120 -7.550 9.290 ;
        RECT -7.870 9.110 -7.550 9.120 ;
        RECT 5.500 9.330 5.820 9.370 ;
        RECT 5.500 9.290 5.830 9.330 ;
        RECT 5.500 9.120 6.080 9.290 ;
        RECT 5.500 9.110 5.820 9.120 ;
      LAYER mcon ;
        RECT -7.780 9.150 -7.610 9.320 ;
        RECT 5.560 9.150 5.730 9.320 ;
      LAYER met1 ;
        RECT -7.860 9.080 -7.540 9.400 ;
        RECT 5.490 9.080 5.810 9.400 ;
      LAYER via ;
        RECT -7.830 9.110 -7.570 9.370 ;
        RECT 5.520 9.110 5.780 9.370 ;
      LAYER met2 ;
        RECT -7.850 9.390 -7.540 9.410 ;
        RECT 5.490 9.390 5.800 9.410 ;
        RECT -10.010 9.220 7.960 9.390 ;
        RECT -10.010 9.210 -7.450 9.220 ;
        RECT 5.400 9.210 7.960 9.220 ;
        RECT -7.850 9.080 -7.540 9.210 ;
        RECT 5.490 9.080 5.800 9.210 ;
    END
  END HORIZ3
  PIN HORIZ4
    USE ANALOG ;
    ANTENNADIFFAREA 0.174000 ;
    PORT
      LAYER li1 ;
        RECT -7.870 8.490 -7.550 8.500 ;
        RECT -8.130 8.320 -7.550 8.490 ;
        RECT -7.880 8.280 -7.550 8.320 ;
        RECT -7.870 8.240 -7.550 8.280 ;
        RECT 5.500 8.490 5.820 8.500 ;
        RECT 5.500 8.320 6.080 8.490 ;
        RECT 5.500 8.280 5.830 8.320 ;
        RECT 5.500 8.240 5.820 8.280 ;
      LAYER mcon ;
        RECT -7.780 8.290 -7.610 8.460 ;
        RECT 5.560 8.290 5.730 8.460 ;
      LAYER met1 ;
        RECT -7.860 8.210 -7.540 8.530 ;
        RECT 5.490 8.210 5.810 8.530 ;
      LAYER via ;
        RECT -7.830 8.240 -7.570 8.500 ;
        RECT 5.520 8.240 5.780 8.500 ;
      LAYER met2 ;
        RECT -7.850 8.410 -7.540 8.530 ;
        RECT 5.490 8.410 5.800 8.530 ;
        RECT -7.850 8.400 5.800 8.410 ;
        RECT -10.010 8.240 7.960 8.400 ;
        RECT -10.010 8.220 -7.450 8.240 ;
        RECT 5.400 8.220 7.960 8.240 ;
        RECT -7.850 8.200 -7.540 8.220 ;
        RECT 5.490 8.200 5.800 8.220 ;
    END
  END HORIZ4
  PIN DRAIN4
    USE ANALOG ;
    ANTENNADIFFAREA 0.198400 ;
    PORT
      LAYER li1 ;
        RECT -7.870 7.920 -7.550 7.950 ;
        RECT -7.880 7.870 -7.550 7.920 ;
        RECT -8.130 7.700 -7.550 7.870 ;
        RECT -7.870 7.690 -7.550 7.700 ;
        RECT 5.500 7.920 5.820 7.950 ;
        RECT 5.500 7.870 5.830 7.920 ;
        RECT 5.500 7.700 6.080 7.870 ;
        RECT 5.500 7.690 5.820 7.700 ;
      LAYER mcon ;
        RECT -7.780 7.740 -7.610 7.910 ;
        RECT 5.560 7.740 5.730 7.910 ;
      LAYER met1 ;
        RECT -7.860 7.660 -7.540 7.980 ;
        RECT 5.490 7.660 5.810 7.980 ;
      LAYER via ;
        RECT -7.830 7.690 -7.570 7.950 ;
        RECT 5.520 7.690 5.780 7.950 ;
      LAYER met2 ;
        RECT -7.850 7.970 -7.540 7.980 ;
        RECT 5.490 7.970 5.800 7.980 ;
        RECT -10.010 7.800 7.960 7.970 ;
        RECT -10.010 7.790 -7.540 7.800 ;
        RECT -7.850 7.650 -7.540 7.790 ;
        RECT 5.490 7.790 7.960 7.800 ;
        RECT 5.490 7.650 5.800 7.790 ;
    END
  END DRAIN4
  PIN VINJ
    ANTENNADIFFAREA 1.020000 ;
    PORT
      LAYER nwell ;
        RECT -10.000 13.320 -3.450 13.330 ;
        RECT -10.010 7.300 -3.450 13.320 ;
        RECT -10.000 7.290 -3.450 7.300 ;
        RECT -7.450 7.280 -3.450 7.290 ;
      LAYER li1 ;
        RECT -9.610 12.650 -9.410 13.000 ;
        RECT -9.620 12.620 -9.410 12.650 ;
        RECT -9.620 12.030 -9.400 12.620 ;
        RECT -9.620 11.000 -9.400 11.590 ;
        RECT -9.620 10.970 -9.410 11.000 ;
        RECT -9.610 10.620 -9.410 10.970 ;
        RECT -9.610 9.640 -9.410 9.990 ;
        RECT -9.620 9.610 -9.410 9.640 ;
        RECT -9.620 9.020 -9.400 9.610 ;
        RECT -9.620 8.000 -9.400 8.590 ;
        RECT -9.620 7.970 -9.410 8.000 ;
        RECT -9.610 7.620 -9.410 7.970 ;
      LAYER mcon ;
        RECT -9.590 12.450 -9.420 12.620 ;
        RECT -9.590 11.000 -9.420 11.170 ;
        RECT -9.590 9.440 -9.420 9.610 ;
        RECT -9.590 8.000 -9.420 8.170 ;
      LAYER met1 ;
        RECT -9.650 12.680 -9.490 13.330 ;
        RECT -9.650 12.130 -9.380 12.680 ;
        RECT -9.660 12.080 -9.380 12.130 ;
        RECT -9.660 11.990 -9.490 12.080 ;
        RECT -9.650 11.630 -9.490 11.990 ;
        RECT -9.660 11.540 -9.490 11.630 ;
        RECT -9.660 11.490 -9.380 11.540 ;
        RECT -9.650 10.940 -9.380 11.490 ;
        RECT -9.650 9.670 -9.490 10.940 ;
        RECT -9.650 9.120 -9.380 9.670 ;
        RECT -9.660 9.070 -9.380 9.120 ;
        RECT -9.660 8.980 -9.490 9.070 ;
        RECT -9.650 8.630 -9.490 8.980 ;
        RECT -9.660 8.540 -9.490 8.630 ;
        RECT -9.660 8.490 -9.380 8.540 ;
        RECT -9.650 7.940 -9.380 8.490 ;
        RECT -9.650 7.290 -9.490 7.940 ;
    END
    PORT
      LAYER nwell ;
        RECT 1.400 13.320 7.950 13.330 ;
        RECT 1.400 7.300 7.960 13.320 ;
        RECT 1.400 7.290 7.950 7.300 ;
        RECT 1.400 7.280 5.400 7.290 ;
      LAYER li1 ;
        RECT 7.360 12.650 7.560 13.000 ;
        RECT 7.360 12.620 7.570 12.650 ;
        RECT 7.350 12.030 7.570 12.620 ;
        RECT 7.350 11.000 7.570 11.590 ;
        RECT 7.360 10.970 7.570 11.000 ;
        RECT 7.360 10.620 7.560 10.970 ;
        RECT 7.360 9.640 7.560 9.990 ;
        RECT 7.360 9.610 7.570 9.640 ;
        RECT 7.350 9.020 7.570 9.610 ;
        RECT 7.350 8.000 7.570 8.590 ;
        RECT 7.360 7.970 7.570 8.000 ;
        RECT 7.360 7.620 7.560 7.970 ;
      LAYER mcon ;
        RECT 7.370 12.450 7.540 12.620 ;
        RECT 7.370 11.000 7.540 11.170 ;
        RECT 7.370 9.440 7.540 9.610 ;
        RECT 7.370 8.000 7.540 8.170 ;
      LAYER met1 ;
        RECT 7.440 12.680 7.600 13.330 ;
        RECT 7.330 12.130 7.600 12.680 ;
        RECT 7.330 12.080 7.610 12.130 ;
        RECT 7.440 11.990 7.610 12.080 ;
        RECT 7.440 11.630 7.600 11.990 ;
        RECT 7.440 11.540 7.610 11.630 ;
        RECT 7.330 11.490 7.610 11.540 ;
        RECT 7.330 10.940 7.600 11.490 ;
        RECT 7.440 9.670 7.600 10.940 ;
        RECT 7.330 9.120 7.600 9.670 ;
        RECT 7.330 9.070 7.610 9.120 ;
        RECT 7.440 8.980 7.610 9.070 ;
        RECT 7.440 8.630 7.600 8.980 ;
        RECT 7.440 8.540 7.610 8.630 ;
        RECT 7.330 8.490 7.610 8.540 ;
        RECT 7.330 7.940 7.600 8.490 ;
        RECT 7.440 7.290 7.600 7.940 ;
    END
  END VINJ
  PIN GATESELECT1
    USE ANALOG ;
    ANTENNAGATEAREA 0.620000 ;
    PORT
      LAYER li1 ;
        RECT -9.240 10.220 -8.800 10.390 ;
      LAYER met1 ;
        RECT -9.240 12.340 -9.050 13.330 ;
        RECT -9.240 12.220 -9.070 12.340 ;
        RECT -9.240 11.400 -9.080 12.220 ;
        RECT -9.240 11.280 -9.070 11.400 ;
        RECT -9.240 10.420 -9.050 11.280 ;
        RECT -9.270 10.190 -9.030 10.420 ;
        RECT -9.240 9.330 -9.050 10.190 ;
        RECT -9.240 9.210 -9.070 9.330 ;
        RECT -9.240 8.400 -9.080 9.210 ;
        RECT -9.240 8.280 -9.070 8.400 ;
        RECT -9.240 7.290 -9.050 8.280 ;
    END
  END GATESELECT1
  PIN VERT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.372000 ;
    PORT
      LAYER li1 ;
        RECT 6.630 12.060 6.830 12.630 ;
        RECT 6.630 10.990 6.830 11.560 ;
        RECT 6.630 9.050 6.830 9.620 ;
        RECT 6.630 7.990 6.830 8.560 ;
      LAYER mcon ;
        RECT 6.640 12.420 6.810 12.590 ;
        RECT 6.640 11.030 6.810 11.200 ;
        RECT 6.640 9.410 6.810 9.580 ;
        RECT 6.640 8.030 6.810 8.200 ;
      LAYER met1 ;
        RECT 6.630 12.650 6.790 13.330 ;
        RECT 6.630 12.630 6.830 12.650 ;
        RECT 6.610 12.390 6.840 12.630 ;
        RECT 6.630 12.170 6.830 12.390 ;
        RECT 6.630 11.450 6.790 12.170 ;
        RECT 6.630 11.230 6.830 11.450 ;
        RECT 6.610 10.990 6.840 11.230 ;
        RECT 6.630 10.970 6.830 10.990 ;
        RECT 6.630 9.640 6.790 10.970 ;
        RECT 6.630 9.620 6.830 9.640 ;
        RECT 6.610 9.380 6.840 9.620 ;
        RECT 6.630 9.160 6.830 9.380 ;
        RECT 6.630 8.450 6.790 9.160 ;
        RECT 6.630 8.230 6.830 8.450 ;
        RECT 6.610 7.990 6.840 8.230 ;
        RECT 6.630 7.970 6.830 7.990 ;
        RECT 6.630 7.290 6.790 7.970 ;
    END
  END VERT2
  PIN GATESELECT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.620000 ;
    PORT
      LAYER li1 ;
        RECT 6.750 10.220 7.190 10.390 ;
      LAYER mcon ;
        RECT 7.010 10.220 7.190 10.390 ;
      LAYER met1 ;
        RECT 7.000 12.340 7.190 13.330 ;
        RECT 7.020 12.220 7.190 12.340 ;
        RECT 7.030 11.400 7.190 12.220 ;
        RECT 7.020 11.280 7.190 11.400 ;
        RECT 7.000 10.420 7.190 11.280 ;
        RECT 6.980 10.190 7.220 10.420 ;
        RECT 7.000 9.330 7.190 10.190 ;
        RECT 7.020 9.210 7.190 9.330 ;
        RECT 7.030 8.400 7.190 9.210 ;
        RECT 7.020 8.280 7.190 8.400 ;
        RECT 7.000 7.290 7.190 8.280 ;
    END
  END GATESELECT2
  PIN GATE2
    USE ANALOG ;
    ANTENNADIFFAREA 1.345600 ;
    PORT
      LAYER li1 ;
        RECT 1.750 12.020 5.060 13.000 ;
        RECT 1.750 10.550 5.060 11.530 ;
        RECT 1.750 9.080 5.060 10.060 ;
        RECT 1.750 7.610 5.060 8.590 ;
      LAYER mcon ;
        RECT 3.320 12.770 3.490 12.940 ;
        RECT 3.320 12.420 3.490 12.590 ;
        RECT 3.320 12.080 3.490 12.250 ;
        RECT 3.320 11.300 3.490 11.470 ;
        RECT 3.320 10.950 3.490 11.120 ;
        RECT 3.320 10.610 3.490 10.780 ;
        RECT 3.320 9.830 3.490 10.000 ;
        RECT 3.320 9.480 3.490 9.650 ;
        RECT 3.320 9.140 3.490 9.310 ;
        RECT 3.320 8.360 3.490 8.530 ;
        RECT 3.320 8.010 3.490 8.180 ;
        RECT 3.320 7.670 3.490 7.840 ;
      LAYER met1 ;
        RECT 3.280 12.100 3.520 13.330 ;
        RECT 3.280 11.880 3.530 12.100 ;
        RECT 3.280 10.630 3.520 11.880 ;
        RECT 3.280 10.410 3.530 10.630 ;
        RECT 3.280 9.160 3.520 10.410 ;
        RECT 3.280 8.940 3.530 9.160 ;
        RECT 3.280 7.690 3.520 8.940 ;
        RECT 3.280 7.470 3.530 7.690 ;
        RECT 3.280 7.280 3.520 7.470 ;
    END
  END GATE2
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 1.345600 ;
    PORT
      LAYER li1 ;
        RECT -7.110 12.020 -3.800 13.000 ;
        RECT -7.110 10.550 -3.800 11.530 ;
        RECT -7.110 9.080 -3.800 10.060 ;
        RECT -7.110 7.610 -3.800 8.590 ;
      LAYER mcon ;
        RECT -5.540 12.770 -5.370 12.940 ;
        RECT -5.540 12.420 -5.370 12.590 ;
        RECT -5.540 12.080 -5.370 12.250 ;
        RECT -5.540 11.300 -5.370 11.470 ;
        RECT -5.540 10.950 -5.370 11.120 ;
        RECT -5.540 10.610 -5.370 10.780 ;
        RECT -5.540 9.830 -5.370 10.000 ;
        RECT -5.540 9.480 -5.370 9.650 ;
        RECT -5.540 9.140 -5.370 9.310 ;
        RECT -5.540 8.360 -5.370 8.530 ;
        RECT -5.540 8.010 -5.370 8.180 ;
        RECT -5.540 7.670 -5.370 7.840 ;
      LAYER met1 ;
        RECT -5.570 12.100 -5.320 13.330 ;
        RECT -5.580 11.880 -5.320 12.100 ;
        RECT -5.570 10.630 -5.320 11.880 ;
        RECT -5.580 10.410 -5.320 10.630 ;
        RECT -5.570 9.160 -5.320 10.410 ;
        RECT -5.580 8.940 -5.320 9.160 ;
        RECT -5.570 7.690 -5.320 8.940 ;
        RECT -5.580 7.470 -5.320 7.690 ;
        RECT -5.570 7.280 -5.320 7.470 ;
    END
  END GATE1
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 0.336400 ;
    PORT
      LAYER li1 ;
        RECT -1.890 12.120 -1.720 13.010 ;
        RECT -1.890 10.600 -1.720 11.490 ;
        RECT -1.890 9.150 -1.720 10.040 ;
        RECT -1.890 7.610 -1.720 8.500 ;
      LAYER mcon ;
        RECT -1.890 12.810 -1.720 12.980 ;
        RECT -1.890 11.290 -1.720 11.460 ;
        RECT -1.890 9.840 -1.720 10.010 ;
        RECT -1.890 8.300 -1.720 8.470 ;
      LAYER met1 ;
        RECT -1.960 7.280 -1.660 13.330 ;
    END
    PORT
      LAYER li1 ;
        RECT -0.330 12.120 -0.160 13.010 ;
        RECT -0.330 10.600 -0.160 11.490 ;
        RECT -0.330 9.150 -0.160 10.040 ;
        RECT -0.330 7.610 -0.160 8.500 ;
      LAYER mcon ;
        RECT -0.330 12.810 -0.160 12.980 ;
        RECT -0.330 11.290 -0.160 11.460 ;
        RECT -0.330 9.840 -0.160 10.010 ;
        RECT -0.330 8.300 -0.160 8.470 ;
      LAYER met1 ;
        RECT -0.380 7.280 -0.080 13.330 ;
    END
  END VTUN
END sky130_hilas_swc4x2cellOverlap

MACRO sky130_hilas_swc4x2cell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc4x2cell ;
  ORIGIN 10.040 0.040 ;
  SIZE 20.130 BY 6.050 ;
  PIN GATE2
    USE ANALOG ;
    ANTENNADIFFAREA 2.743300 ;
    PORT
      LAYER nwell ;
        RECT 3.760 -0.030 5.990 6.000 ;
      LAYER li1 ;
        RECT 4.460 2.690 5.010 3.120 ;
      LAYER mcon ;
        RECT 4.460 2.770 4.730 3.040 ;
      LAYER met1 ;
        RECT 4.410 4.090 4.790 6.010 ;
        RECT 4.400 2.230 4.790 4.090 ;
        RECT 4.410 -0.040 4.790 2.230 ;
    END
  END GATE2
  PIN VTUN
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -1.700 -0.040 1.740 6.010 ;
      LAYER li1 ;
        RECT -0.940 2.760 -0.390 3.190 ;
        RECT 0.430 2.760 0.980 3.190 ;
      LAYER mcon ;
        RECT -0.660 2.840 -0.390 3.110 ;
        RECT 0.430 2.840 0.700 3.110 ;
      LAYER met1 ;
        RECT -0.720 -0.040 -0.320 6.010 ;
        RECT 0.360 -0.040 0.760 6.010 ;
    END
  END VTUN
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 2.743300 ;
    PORT
      LAYER nwell ;
        RECT -5.950 -0.030 -3.720 6.000 ;
      LAYER li1 ;
        RECT -4.970 2.690 -4.420 3.120 ;
      LAYER mcon ;
        RECT -4.690 2.770 -4.420 3.040 ;
      LAYER met1 ;
        RECT -4.750 4.090 -4.370 6.010 ;
        RECT -4.750 2.230 -4.360 4.090 ;
        RECT -4.750 -0.040 -4.370 2.230 ;
    END
  END GATE1
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 7.520 6.000 10.070 6.010 ;
        RECT 7.520 -0.020 10.080 6.000 ;
        RECT 7.520 -0.030 10.070 -0.020 ;
      LAYER li1 ;
        RECT 9.480 5.330 9.680 5.680 ;
        RECT 9.480 5.300 9.690 5.330 ;
        RECT 9.470 4.710 9.690 5.300 ;
        RECT 9.470 3.680 9.690 4.270 ;
        RECT 9.480 3.650 9.690 3.680 ;
        RECT 9.480 3.300 9.680 3.650 ;
        RECT 9.480 2.320 9.680 2.670 ;
        RECT 9.480 2.290 9.690 2.320 ;
        RECT 9.470 1.700 9.690 2.290 ;
        RECT 9.470 0.680 9.690 1.270 ;
        RECT 9.480 0.650 9.690 0.680 ;
        RECT 9.480 0.300 9.680 0.650 ;
      LAYER mcon ;
        RECT 9.490 5.130 9.660 5.300 ;
        RECT 9.490 3.680 9.660 3.850 ;
        RECT 9.490 2.120 9.660 2.290 ;
        RECT 9.490 0.680 9.660 0.850 ;
      LAYER met1 ;
        RECT 9.560 5.360 9.720 6.010 ;
        RECT 9.450 4.810 9.720 5.360 ;
        RECT 9.450 4.760 9.730 4.810 ;
        RECT 9.560 4.670 9.730 4.760 ;
        RECT 9.560 4.310 9.720 4.670 ;
        RECT 9.560 4.220 9.730 4.310 ;
        RECT 9.450 4.170 9.730 4.220 ;
        RECT 9.450 3.620 9.720 4.170 ;
        RECT 9.560 2.350 9.720 3.620 ;
        RECT 9.450 1.800 9.720 2.350 ;
        RECT 9.450 1.750 9.730 1.800 ;
        RECT 9.560 1.660 9.730 1.750 ;
        RECT 9.560 1.310 9.720 1.660 ;
        RECT 9.560 1.220 9.730 1.310 ;
        RECT 9.450 1.170 9.730 1.220 ;
        RECT 9.450 0.620 9.720 1.170 ;
        RECT 9.560 -0.030 9.720 0.620 ;
    END
  END VPWR
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -10.030 6.000 -7.480 6.010 ;
        RECT -10.040 -0.020 -7.480 6.000 ;
        RECT -10.030 -0.030 -7.480 -0.020 ;
      LAYER li1 ;
        RECT -9.640 5.330 -9.440 5.680 ;
        RECT -9.650 5.300 -9.440 5.330 ;
        RECT -9.650 4.710 -9.430 5.300 ;
        RECT -9.650 3.680 -9.430 4.270 ;
        RECT -9.650 3.650 -9.440 3.680 ;
        RECT -9.640 3.300 -9.440 3.650 ;
        RECT -9.640 2.320 -9.440 2.670 ;
        RECT -9.650 2.290 -9.440 2.320 ;
        RECT -9.650 1.700 -9.430 2.290 ;
        RECT -9.650 0.680 -9.430 1.270 ;
        RECT -9.650 0.650 -9.440 0.680 ;
        RECT -9.640 0.300 -9.440 0.650 ;
      LAYER mcon ;
        RECT -9.620 5.130 -9.450 5.300 ;
        RECT -9.620 3.680 -9.450 3.850 ;
        RECT -9.620 2.120 -9.450 2.290 ;
        RECT -9.620 0.680 -9.450 0.850 ;
      LAYER met1 ;
        RECT -9.680 5.360 -9.520 6.010 ;
        RECT -9.680 4.810 -9.410 5.360 ;
        RECT -9.690 4.760 -9.410 4.810 ;
        RECT -9.690 4.670 -9.520 4.760 ;
        RECT -9.680 4.310 -9.520 4.670 ;
        RECT -9.690 4.220 -9.520 4.310 ;
        RECT -9.690 4.170 -9.410 4.220 ;
        RECT -9.680 3.620 -9.410 4.170 ;
        RECT -9.680 2.350 -9.520 3.620 ;
        RECT -9.680 1.800 -9.410 2.350 ;
        RECT -9.690 1.750 -9.410 1.800 ;
        RECT -9.690 1.660 -9.520 1.750 ;
        RECT -9.680 1.310 -9.520 1.660 ;
        RECT -9.690 1.220 -9.520 1.310 ;
        RECT -9.690 1.170 -9.410 1.220 ;
        RECT -9.680 0.620 -9.410 1.170 ;
        RECT -9.680 -0.040 -9.520 0.620 ;
    END
  END VINJ
  PIN GATESELECT1
    USE ANALOG ;
    ANTENNAGATEAREA 0.620000 ;
    PORT
      LAYER li1 ;
        RECT -9.270 2.900 -8.830 3.070 ;
      LAYER met1 ;
        RECT -9.270 5.020 -9.080 6.010 ;
        RECT -9.270 4.900 -9.100 5.020 ;
        RECT -9.270 4.080 -9.110 4.900 ;
        RECT -9.270 3.960 -9.100 4.080 ;
        RECT -9.270 3.100 -9.080 3.960 ;
        RECT -9.300 2.870 -9.060 3.100 ;
        RECT -9.270 2.010 -9.080 2.870 ;
        RECT -9.270 1.890 -9.100 2.010 ;
        RECT -9.270 1.080 -9.110 1.890 ;
        RECT -9.270 0.960 -9.100 1.080 ;
        RECT -9.270 -0.030 -9.080 0.960 ;
    END
  END GATESELECT1
  PIN GATESELECT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.620000 ;
    PORT
      LAYER li1 ;
        RECT 8.870 2.900 9.310 3.070 ;
      LAYER mcon ;
        RECT 9.130 2.900 9.310 3.070 ;
      LAYER met1 ;
        RECT 9.120 5.020 9.310 6.010 ;
        RECT 9.140 4.900 9.310 5.020 ;
        RECT 9.150 4.080 9.310 4.900 ;
        RECT 9.140 3.960 9.310 4.080 ;
        RECT 9.120 3.100 9.310 3.960 ;
        RECT 9.100 2.870 9.340 3.100 ;
        RECT 9.120 2.010 9.310 2.870 ;
        RECT 9.140 1.890 9.310 2.010 ;
        RECT 9.150 1.080 9.310 1.890 ;
        RECT 9.140 0.960 9.310 1.080 ;
        RECT 9.120 -0.030 9.310 0.960 ;
    END
  END GATESELECT2
  PIN VERT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.372000 ;
    PORT
      LAYER li1 ;
        RECT -8.910 4.740 -8.710 5.310 ;
        RECT -8.910 3.670 -8.710 4.240 ;
        RECT -8.910 1.730 -8.710 2.300 ;
        RECT -8.910 0.670 -8.710 1.240 ;
      LAYER mcon ;
        RECT -8.890 5.100 -8.720 5.270 ;
        RECT -8.890 3.710 -8.720 3.880 ;
        RECT -8.890 2.090 -8.720 2.260 ;
        RECT -8.890 0.710 -8.720 0.880 ;
      LAYER met1 ;
        RECT -8.870 5.330 -8.710 6.010 ;
        RECT -8.910 5.310 -8.710 5.330 ;
        RECT -8.920 5.070 -8.690 5.310 ;
        RECT -8.910 4.850 -8.710 5.070 ;
        RECT -8.870 4.130 -8.710 4.850 ;
        RECT -8.910 3.910 -8.710 4.130 ;
        RECT -8.920 3.670 -8.690 3.910 ;
        RECT -8.910 3.650 -8.710 3.670 ;
        RECT -8.870 2.320 -8.710 3.650 ;
        RECT -8.910 2.300 -8.710 2.320 ;
        RECT -8.920 2.060 -8.690 2.300 ;
        RECT -8.910 1.840 -8.710 2.060 ;
        RECT -8.870 1.130 -8.710 1.840 ;
        RECT -8.910 0.910 -8.710 1.130 ;
        RECT -8.920 0.670 -8.690 0.910 ;
        RECT -8.910 0.650 -8.710 0.670 ;
        RECT -8.870 -0.030 -8.710 0.650 ;
    END
  END VERT1
  PIN VERT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.372000 ;
    PORT
      LAYER li1 ;
        RECT 8.750 4.740 8.950 5.310 ;
        RECT 8.750 3.670 8.950 4.240 ;
        RECT 8.750 1.730 8.950 2.300 ;
        RECT 8.750 0.670 8.950 1.240 ;
      LAYER mcon ;
        RECT 8.760 5.100 8.930 5.270 ;
        RECT 8.760 3.710 8.930 3.880 ;
        RECT 8.760 2.090 8.930 2.260 ;
        RECT 8.760 0.710 8.930 0.880 ;
      LAYER met1 ;
        RECT 8.750 5.330 8.910 6.010 ;
        RECT 8.750 5.310 8.950 5.330 ;
        RECT 8.730 5.070 8.960 5.310 ;
        RECT 8.750 4.850 8.950 5.070 ;
        RECT 8.750 4.130 8.910 4.850 ;
        RECT 8.750 3.910 8.950 4.130 ;
        RECT 8.730 3.670 8.960 3.910 ;
        RECT 8.750 3.650 8.950 3.670 ;
        RECT 8.750 2.320 8.910 3.650 ;
        RECT 8.750 2.300 8.950 2.320 ;
        RECT 8.730 2.060 8.960 2.300 ;
        RECT 8.750 1.840 8.950 2.060 ;
        RECT 8.750 1.130 8.910 1.840 ;
        RECT 8.750 0.910 8.950 1.130 ;
        RECT 8.730 0.670 8.960 0.910 ;
        RECT 8.750 0.650 8.950 0.670 ;
        RECT 8.750 -0.030 8.910 0.650 ;
    END
  END VERT2
  PIN HORIZ1
    USE ANALOG ;
    ANTENNADIFFAREA 0.174000 ;
    PORT
      LAYER li1 ;
        RECT -7.900 5.020 -7.580 5.060 ;
        RECT -7.910 4.980 -7.580 5.020 ;
        RECT -8.160 4.810 -7.580 4.980 ;
        RECT -7.900 4.800 -7.580 4.810 ;
        RECT 7.620 5.020 7.940 5.060 ;
        RECT 7.620 4.980 7.950 5.020 ;
        RECT 7.620 4.810 8.200 4.980 ;
        RECT 7.620 4.800 7.940 4.810 ;
      LAYER mcon ;
        RECT -7.810 4.840 -7.640 5.010 ;
        RECT 7.680 4.840 7.850 5.010 ;
      LAYER met1 ;
        RECT -7.890 4.770 -7.570 5.090 ;
        RECT 7.610 4.770 7.930 5.090 ;
      LAYER via ;
        RECT -7.860 4.800 -7.600 5.060 ;
        RECT 7.640 4.800 7.900 5.060 ;
      LAYER met2 ;
        RECT -7.880 5.080 -7.570 5.100 ;
        RECT 7.610 5.080 7.920 5.100 ;
        RECT -10.040 4.900 10.080 5.080 ;
        RECT -7.880 4.770 -7.570 4.900 ;
        RECT 7.610 4.770 7.920 4.900 ;
    END
  END HORIZ1
  PIN HORIZ2
    USE ANALOG ;
    ANTENNADIFFAREA 0.174000 ;
    PORT
      LAYER li1 ;
        RECT -7.900 4.170 -7.580 4.180 ;
        RECT -8.160 4.000 -7.580 4.170 ;
        RECT -7.910 3.960 -7.580 4.000 ;
        RECT -7.900 3.920 -7.580 3.960 ;
        RECT 7.620 4.170 7.940 4.180 ;
        RECT 7.620 4.000 8.200 4.170 ;
        RECT 7.620 3.960 7.950 4.000 ;
        RECT 7.620 3.920 7.940 3.960 ;
      LAYER mcon ;
        RECT -7.810 3.970 -7.640 4.140 ;
        RECT 7.680 3.970 7.850 4.140 ;
      LAYER met1 ;
        RECT -7.890 3.890 -7.570 4.210 ;
        RECT 7.610 3.890 7.930 4.210 ;
      LAYER via ;
        RECT -7.860 3.920 -7.600 4.180 ;
        RECT 7.640 3.920 7.900 4.180 ;
      LAYER met2 ;
        RECT -10.040 4.080 -9.970 4.090 ;
        RECT -7.880 4.080 -7.570 4.210 ;
        RECT 7.610 4.080 7.920 4.210 ;
        RECT -10.040 3.900 10.090 4.080 ;
        RECT -7.880 3.880 -7.570 3.900 ;
        RECT 7.610 3.880 7.920 3.900 ;
    END
  END HORIZ2
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.198400 ;
    PORT
      LAYER li1 ;
        RECT -7.900 5.600 -7.580 5.610 ;
        RECT -8.160 5.430 -7.580 5.600 ;
        RECT -7.910 5.380 -7.580 5.430 ;
        RECT -7.900 5.350 -7.580 5.380 ;
        RECT 7.620 5.600 7.940 5.610 ;
        RECT 7.620 5.430 8.200 5.600 ;
        RECT 7.620 5.380 7.950 5.430 ;
        RECT 7.620 5.350 7.940 5.380 ;
      LAYER mcon ;
        RECT -7.810 5.390 -7.640 5.560 ;
        RECT 7.680 5.390 7.850 5.560 ;
      LAYER met1 ;
        RECT -7.890 5.320 -7.570 5.640 ;
        RECT 7.610 5.320 7.930 5.640 ;
      LAYER via ;
        RECT -7.860 5.350 -7.600 5.610 ;
        RECT 7.640 5.350 7.900 5.610 ;
      LAYER met2 ;
        RECT -10.040 5.510 -9.900 5.520 ;
        RECT -7.880 5.510 -7.570 5.650 ;
        RECT 7.610 5.510 7.920 5.650 ;
        RECT -10.040 5.330 10.080 5.510 ;
        RECT -7.880 5.320 -7.570 5.330 ;
        RECT 7.610 5.320 7.920 5.330 ;
    END
  END DRAIN1
  PIN DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.198400 ;
    PORT
      LAYER li1 ;
        RECT -7.900 3.600 -7.580 3.630 ;
        RECT -7.910 3.550 -7.580 3.600 ;
        RECT -8.160 3.380 -7.580 3.550 ;
        RECT -7.900 3.370 -7.580 3.380 ;
        RECT 7.620 3.600 7.940 3.630 ;
        RECT 7.620 3.550 7.950 3.600 ;
        RECT 7.620 3.380 8.200 3.550 ;
        RECT 7.620 3.370 7.940 3.380 ;
      LAYER mcon ;
        RECT -7.810 3.420 -7.640 3.590 ;
        RECT 7.680 3.420 7.850 3.590 ;
      LAYER met1 ;
        RECT -7.890 3.340 -7.570 3.660 ;
        RECT 7.610 3.340 7.930 3.660 ;
      LAYER via ;
        RECT -7.860 3.370 -7.600 3.630 ;
        RECT 7.640 3.370 7.900 3.630 ;
      LAYER met2 ;
        RECT -7.880 3.650 -7.570 3.660 ;
        RECT 7.610 3.650 7.920 3.660 ;
        RECT -10.040 3.470 10.090 3.650 ;
        RECT -7.880 3.330 -7.570 3.470 ;
        RECT 7.610 3.330 7.920 3.470 ;
    END
    PORT
      LAYER li1 ;
        RECT -7.900 0.600 -7.580 0.630 ;
        RECT -7.910 0.550 -7.580 0.600 ;
        RECT -8.160 0.380 -7.580 0.550 ;
        RECT -7.900 0.370 -7.580 0.380 ;
        RECT 7.620 0.600 7.940 0.630 ;
        RECT 7.620 0.550 7.950 0.600 ;
        RECT 7.620 0.380 8.200 0.550 ;
        RECT 7.620 0.370 7.940 0.380 ;
      LAYER mcon ;
        RECT -7.810 0.420 -7.640 0.590 ;
        RECT 7.680 0.420 7.850 0.590 ;
      LAYER met1 ;
        RECT -7.890 0.340 -7.570 0.660 ;
        RECT 7.610 0.340 7.930 0.660 ;
      LAYER via ;
        RECT -7.860 0.370 -7.600 0.630 ;
        RECT 7.640 0.370 7.900 0.630 ;
      LAYER met2 ;
        RECT -7.880 0.650 -7.570 0.660 ;
        RECT 7.610 0.650 7.920 0.660 ;
        RECT -10.040 0.480 10.090 0.650 ;
        RECT -10.040 0.470 -7.570 0.480 ;
        RECT -7.880 0.330 -7.570 0.470 ;
        RECT 7.610 0.470 10.090 0.480 ;
        RECT 7.610 0.330 7.920 0.470 ;
    END
  END DRAIN2
  PIN DRAIN3
    USE ANALOG ;
    ANTENNADIFFAREA 0.198400 ;
    PORT
      LAYER li1 ;
        RECT -7.900 2.590 -7.580 2.600 ;
        RECT -8.160 2.420 -7.580 2.590 ;
        RECT -7.910 2.370 -7.580 2.420 ;
        RECT -7.900 2.340 -7.580 2.370 ;
        RECT 7.620 2.590 7.940 2.600 ;
        RECT 7.620 2.420 8.200 2.590 ;
        RECT 7.620 2.370 7.950 2.420 ;
        RECT 7.620 2.340 7.940 2.370 ;
      LAYER mcon ;
        RECT -7.810 2.380 -7.640 2.550 ;
        RECT 7.680 2.380 7.850 2.550 ;
      LAYER met1 ;
        RECT -7.890 2.310 -7.570 2.630 ;
        RECT 7.610 2.310 7.930 2.630 ;
      LAYER via ;
        RECT -7.860 2.340 -7.600 2.600 ;
        RECT 7.640 2.340 7.900 2.600 ;
      LAYER met2 ;
        RECT -7.880 2.500 -7.570 2.640 ;
        RECT -10.040 2.490 -7.570 2.500 ;
        RECT 7.610 2.500 7.920 2.640 ;
        RECT 7.610 2.490 10.090 2.500 ;
        RECT -10.040 2.320 10.090 2.490 ;
        RECT -7.880 2.310 -7.570 2.320 ;
        RECT 7.610 2.310 7.920 2.320 ;
    END
  END DRAIN3
  PIN HORIZ3
    USE ANALOG ;
    ANTENNADIFFAREA 0.174000 ;
    PORT
      LAYER li1 ;
        RECT -7.900 2.010 -7.580 2.050 ;
        RECT -7.910 1.970 -7.580 2.010 ;
        RECT -8.160 1.800 -7.580 1.970 ;
        RECT -7.900 1.790 -7.580 1.800 ;
        RECT 7.620 2.010 7.940 2.050 ;
        RECT 7.620 1.970 7.950 2.010 ;
        RECT 7.620 1.800 8.200 1.970 ;
        RECT 7.620 1.790 7.940 1.800 ;
      LAYER mcon ;
        RECT -7.810 1.830 -7.640 2.000 ;
        RECT 7.680 1.830 7.850 2.000 ;
      LAYER met1 ;
        RECT -7.890 1.760 -7.570 2.080 ;
        RECT 7.610 1.760 7.930 2.080 ;
      LAYER via ;
        RECT -7.860 1.790 -7.600 2.050 ;
        RECT 7.640 1.790 7.900 2.050 ;
      LAYER met2 ;
        RECT -7.880 2.070 -7.570 2.090 ;
        RECT 7.610 2.070 7.920 2.090 ;
        RECT -10.040 1.900 10.090 2.070 ;
        RECT -10.040 1.890 -7.480 1.900 ;
        RECT 7.520 1.890 10.090 1.900 ;
        RECT -7.880 1.760 -7.570 1.890 ;
        RECT 7.610 1.760 7.920 1.890 ;
    END
  END HORIZ3
  PIN HORIZ4
    USE ANALOG ;
    ANTENNADIFFAREA 0.174000 ;
    PORT
      LAYER li1 ;
        RECT -7.900 1.170 -7.580 1.180 ;
        RECT -8.160 1.000 -7.580 1.170 ;
        RECT -7.910 0.960 -7.580 1.000 ;
        RECT -7.900 0.920 -7.580 0.960 ;
        RECT 7.620 1.170 7.940 1.180 ;
        RECT 7.620 1.000 8.200 1.170 ;
        RECT 7.620 0.960 7.950 1.000 ;
        RECT 7.620 0.920 7.940 0.960 ;
      LAYER mcon ;
        RECT -7.810 0.970 -7.640 1.140 ;
        RECT 7.680 0.970 7.850 1.140 ;
      LAYER met1 ;
        RECT -7.890 0.890 -7.570 1.210 ;
        RECT 7.610 0.890 7.930 1.210 ;
      LAYER via ;
        RECT -7.860 0.920 -7.600 1.180 ;
        RECT 7.640 0.920 7.900 1.180 ;
      LAYER met2 ;
        RECT -7.880 1.090 -7.570 1.210 ;
        RECT 7.610 1.090 7.920 1.210 ;
        RECT -7.880 1.080 7.920 1.090 ;
        RECT -10.040 0.920 10.090 1.080 ;
        RECT -10.040 0.900 -7.480 0.920 ;
        RECT -7.880 0.880 -7.570 0.900 ;
        RECT -2.300 0.830 -0.760 0.920 ;
        RECT 0.800 0.830 2.340 0.920 ;
        RECT 7.520 0.900 10.090 0.920 ;
        RECT 7.610 0.880 7.920 0.900 ;
    END
  END HORIZ4
END sky130_hilas_swc4x2cell

MACRO sky130_hilas_TACoreBlock2
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TACoreBlock2 ;
  ORIGIN 0.610 1.920 ;
  SIZE 2.190 BY 4.770 ;
  OBS
      LAYER nwell ;
        RECT -0.610 1.120 1.580 2.850 ;
      LAYER li1 ;
        RECT -0.400 2.010 1.360 2.530 ;
        RECT -0.400 1.400 0.310 1.570 ;
        RECT 0.620 1.400 1.320 1.570 ;
        RECT -0.050 1.230 0.310 1.400 ;
        RECT -0.050 0.870 0.600 1.230 ;
        RECT -0.050 0.640 0.220 0.870 ;
        RECT 0.850 0.650 1.100 1.400 ;
        RECT -0.080 0.470 0.250 0.640 ;
        RECT 0.770 0.470 1.100 0.650 ;
        RECT -0.120 -0.200 0.290 0.040 ;
        RECT 0.730 -0.200 1.140 0.040 ;
        RECT -0.120 -0.580 1.140 -0.200 ;
        RECT -0.120 -0.840 0.290 -0.580 ;
        RECT 0.730 -0.830 1.140 -0.580 ;
        RECT -0.090 -1.430 0.250 -1.260 ;
        RECT 0.760 -1.430 1.120 -1.250 ;
        RECT -0.010 -1.920 0.170 -1.430 ;
        RECT 0.840 -1.920 1.030 -1.430 ;
  END
END sky130_hilas_TACoreBlock2

MACRO sky130_hilas_nDiffThOxContact
  CLASS BLOCK ;
  FOREIGN sky130_hilas_nDiffThOxContact ;
  ORIGIN 0.260 -0.130 ;
  SIZE 0.670 BY 0.290 ;
  OBS
      LAYER li1 ;
        RECT -0.260 0.180 0.410 0.350 ;
      LAYER mcon ;
        RECT -0.010 0.180 0.160 0.350 ;
      LAYER met1 ;
        RECT -0.120 0.150 0.270 0.380 ;
  END
END sky130_hilas_nDiffThOxContact

MACRO sky130_hilas_capacitorSize01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_capacitorSize01 ;
  ORIGIN -14.140 0.480 ;
  SIZE 10.420 BY 5.830 ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 23.870 2.610 24.240 2.670 ;
        RECT 23.870 2.330 24.560 2.610 ;
        RECT 23.870 2.270 24.240 2.330 ;
      LAYER via2 ;
        RECT 23.920 2.330 24.200 2.610 ;
      LAYER met3 ;
        RECT 15.600 5.320 18.420 5.350 ;
        RECT 15.600 2.820 22.800 5.320 ;
        RECT 15.600 2.070 24.440 2.820 ;
        RECT 15.600 -0.460 22.800 2.070 ;
        RECT 18.390 -0.480 22.800 -0.460 ;
      LAYER via3 ;
        RECT 23.840 2.220 24.270 2.700 ;
      LAYER met4 ;
        RECT 23.740 2.130 24.400 2.790 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 14.380 2.600 14.750 2.660 ;
        RECT 14.160 2.320 14.750 2.600 ;
        RECT 14.380 2.260 14.750 2.320 ;
      LAYER via2 ;
        RECT 14.430 2.320 14.710 2.600 ;
      LAYER met3 ;
        RECT 14.160 2.060 14.950 2.810 ;
      LAYER via3 ;
        RECT 14.350 2.210 14.780 2.690 ;
      LAYER met4 ;
        RECT 14.250 2.720 14.910 2.780 ;
        RECT 15.300 2.720 16.310 2.730 ;
        RECT 14.250 2.220 17.940 2.720 ;
        RECT 14.250 2.210 15.660 2.220 ;
        RECT 14.250 2.120 14.910 2.210 ;
        RECT 17.300 1.100 17.930 2.220 ;
        RECT 17.300 1.090 19.450 1.100 ;
        RECT 16.490 0.620 19.530 1.090 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 14.140 4.800 24.560 4.980 ;
        RECT 14.140 4.370 24.560 4.550 ;
        RECT 14.170 3.370 24.560 3.550 ;
        RECT 22.650 3.120 24.560 3.130 ;
        RECT 14.170 2.940 24.560 3.120 ;
        RECT 14.170 1.790 24.560 1.960 ;
        RECT 14.170 1.370 24.560 1.540 ;
        RECT 14.170 0.390 24.560 0.560 ;
        RECT 14.170 -0.050 24.560 0.120 ;
  END
END sky130_hilas_capacitorSize01

MACRO sky130_hilas_FGtrans2x1cell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_FGtrans2x1cell ;
  ORIGIN 3.950 3.820 ;
  SIZE 11.520 BY 6.050 ;
  PIN GATESELECT
    USE ANALOG ;
    ANTENNAGATEAREA 0.310000 ;
    PORT
      LAYER li1 ;
        RECT 6.610 0.760 6.800 0.770 ;
        RECT 6.610 0.470 6.810 0.760 ;
        RECT 6.600 0.140 6.840 0.470 ;
        RECT 6.600 -2.060 6.840 -1.730 ;
        RECT 6.610 -2.350 6.810 -2.060 ;
        RECT 6.610 -2.360 6.800 -2.350 ;
      LAYER mcon ;
        RECT 6.620 0.510 6.800 0.700 ;
        RECT 6.620 -2.290 6.800 -2.100 ;
      LAYER met1 ;
        RECT 6.610 0.770 6.800 2.230 ;
        RECT 6.610 0.740 6.830 0.770 ;
        RECT 6.590 0.470 6.840 0.740 ;
        RECT 6.600 0.460 6.840 0.470 ;
        RECT 6.600 0.220 6.830 0.460 ;
        RECT 6.640 -1.810 6.800 0.220 ;
        RECT 6.600 -2.050 6.830 -1.810 ;
        RECT 6.600 -2.060 6.840 -2.050 ;
        RECT 6.590 -2.330 6.840 -2.060 ;
        RECT 6.610 -2.360 6.830 -2.330 ;
        RECT 6.610 -3.820 6.800 -2.360 ;
    END
  END GATESELECT
  PIN VINJ
    USE ANALOG ;
    ANTENNADIFFAREA 0.510000 ;
    PORT
      LAYER nwell ;
        RECT 4.260 -3.810 7.570 2.220 ;
      LAYER li1 ;
        RECT 6.970 1.550 7.170 1.900 ;
        RECT 6.970 1.520 7.180 1.550 ;
        RECT 6.960 0.940 7.180 1.520 ;
        RECT 6.970 0.930 7.180 0.940 ;
        RECT 6.970 -2.530 7.180 -2.520 ;
        RECT 6.960 -3.110 7.180 -2.530 ;
        RECT 6.970 -3.140 7.180 -3.110 ;
        RECT 6.970 -3.490 7.170 -3.140 ;
      LAYER mcon ;
        RECT 6.980 1.350 7.150 1.520 ;
        RECT 6.980 -3.110 7.150 -2.940 ;
      LAYER met1 ;
        RECT 7.050 1.580 7.210 2.230 ;
        RECT 6.940 1.030 7.210 1.580 ;
        RECT 6.940 0.980 7.220 1.030 ;
        RECT 7.050 0.890 7.220 0.980 ;
        RECT 7.050 -2.480 7.210 0.890 ;
        RECT 7.050 -2.570 7.220 -2.480 ;
        RECT 6.940 -2.620 7.220 -2.570 ;
        RECT 6.940 -3.170 7.210 -2.620 ;
        RECT 7.050 -3.820 7.210 -3.170 ;
    END
  END VINJ
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER li1 ;
        RECT 5.410 0.170 5.580 1.260 ;
        RECT 5.410 0.130 5.810 0.170 ;
        RECT 5.410 -0.060 5.820 0.130 ;
        RECT 5.410 -0.090 5.810 -0.060 ;
        RECT 5.410 -0.430 5.580 -0.090 ;
      LAYER mcon ;
        RECT 5.550 -0.050 5.720 0.120 ;
      LAYER met1 ;
        RECT 5.480 -0.120 5.800 0.200 ;
      LAYER via ;
        RECT 5.510 -0.090 5.770 0.170 ;
      LAYER met2 ;
        RECT 5.480 0.190 5.790 0.210 ;
        RECT -3.950 0.000 5.790 0.190 ;
        RECT 5.480 -0.120 5.790 0.000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.160 1.650 5.690 1.820 ;
      LAYER met1 ;
        RECT 5.090 1.550 5.390 1.930 ;
      LAYER via ;
        RECT 5.110 1.610 5.370 1.880 ;
      LAYER met2 ;
        RECT 5.090 1.750 5.390 1.930 ;
        RECT 4.840 1.730 5.390 1.750 ;
        RECT -3.950 1.550 7.570 1.730 ;
    END
  END DRAIN1
  PIN DRAIN4
    USE ANALOG ;
    ANTENNADIFFAREA 0.105400 ;
    PORT
      LAYER li1 ;
        RECT 5.160 -3.410 5.690 -3.240 ;
      LAYER met1 ;
        RECT 5.090 -3.520 5.390 -3.140 ;
      LAYER via ;
        RECT 5.110 -3.470 5.370 -3.200 ;
      LAYER met2 ;
        RECT 5.100 -3.140 5.260 -3.130 ;
        RECT 5.010 -3.150 7.570 -3.140 ;
        RECT -3.950 -3.300 7.570 -3.150 ;
        RECT 5.010 -3.320 7.570 -3.300 ;
        RECT 5.090 -3.520 5.390 -3.320 ;
    END
  END DRAIN4
  PIN PROG
    USE ANALOG ;
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER li1 ;
        RECT 3.860 -0.920 4.070 -0.490 ;
        RECT 3.880 -0.940 4.050 -0.920 ;
      LAYER met1 ;
        RECT 3.840 -0.490 4.050 2.230 ;
        RECT 3.840 -1.000 4.080 -0.490 ;
        RECT 3.840 -3.820 4.050 -1.000 ;
    END
  END PROG
  PIN RUN
    USE ANALOG ;
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER li1 ;
        RECT 2.800 -2.360 2.970 -2.300 ;
        RECT 2.780 -2.570 2.990 -2.360 ;
        RECT 2.800 -2.640 2.970 -2.570 ;
      LAYER met1 ;
        RECT 2.790 -2.300 2.970 2.230 ;
        RECT 2.740 -2.640 3.030 -2.300 ;
        RECT 2.790 -3.820 2.970 -2.640 ;
    END
  END RUN
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 0.217200 ;
    PORT
      LAYER li1 ;
        RECT 4.640 -1.250 4.990 -1.080 ;
        RECT 4.720 -1.460 4.910 -1.250 ;
        RECT 3.290 -2.830 4.100 -2.660 ;
        RECT 3.910 -3.170 4.100 -2.830 ;
        RECT 4.700 -3.170 4.890 -3.140 ;
        RECT 3.910 -3.350 4.890 -3.170 ;
        RECT 4.700 -3.370 4.890 -3.350 ;
      LAYER mcon ;
        RECT 4.730 -1.430 4.900 -1.260 ;
        RECT 4.710 -3.340 4.880 -3.170 ;
      LAYER met1 ;
        RECT 4.720 -1.200 4.910 -1.070 ;
        RECT 4.700 -1.490 4.930 -1.200 ;
        RECT 4.720 -3.110 4.910 -1.490 ;
        RECT 4.680 -3.320 4.910 -3.110 ;
        RECT 4.680 -3.400 4.920 -3.320 ;
        RECT 4.690 -3.820 4.920 -3.400 ;
    END
  END GATE1
  PIN GATE2
    USE ANALOG ;
    ANTENNADIFFAREA 0.217200 ;
    PORT
      LAYER li1 ;
        RECT 4.730 1.800 4.920 1.830 ;
        RECT 3.860 1.630 4.920 1.800 ;
        RECT 3.860 1.240 4.030 1.630 ;
        RECT 4.730 1.600 4.920 1.630 ;
        RECT 3.290 1.070 4.030 1.240 ;
        RECT 4.730 -0.340 4.920 -0.160 ;
        RECT 4.640 -0.510 4.990 -0.340 ;
      LAYER mcon ;
        RECT 4.740 1.630 4.910 1.800 ;
        RECT 4.740 -0.360 4.910 -0.190 ;
      LAYER met1 ;
        RECT 4.720 1.860 4.930 2.230 ;
        RECT 4.710 1.570 4.940 1.860 ;
        RECT 4.720 -0.130 4.930 1.570 ;
        RECT 4.710 -0.420 4.940 -0.130 ;
        RECT 4.720 -0.560 4.930 -0.420 ;
    END
  END GATE2
  PIN PROGGATE
    USE ANALOG ;
    ANTENNADIFFAREA 0.434600 ;
    PORT
      LAYER li1 ;
        RECT 4.260 1.240 4.450 1.270 ;
        RECT 4.260 1.070 4.990 1.240 ;
        RECT 4.260 1.040 4.450 1.070 ;
        RECT 3.300 -0.510 3.640 -0.340 ;
        RECT 3.380 -1.080 3.550 -0.510 ;
        RECT 3.300 -1.110 3.640 -1.080 ;
        RECT 4.260 -1.100 4.450 -1.050 ;
        RECT 4.220 -1.110 4.450 -1.100 ;
        RECT 3.300 -1.250 4.450 -1.110 ;
        RECT 3.470 -1.280 4.450 -1.250 ;
        RECT 3.470 -1.310 4.310 -1.280 ;
        RECT 4.270 -2.660 4.460 -2.630 ;
        RECT 4.270 -2.830 4.990 -2.660 ;
        RECT 4.270 -2.860 4.460 -2.830 ;
      LAYER mcon ;
        RECT 4.270 1.070 4.440 1.240 ;
        RECT 4.270 -1.250 4.440 -1.080 ;
        RECT 4.280 -2.830 4.450 -2.660 ;
      LAYER met1 ;
        RECT 4.270 1.300 4.460 2.230 ;
        RECT 4.240 1.010 4.470 1.300 ;
        RECT 4.270 -1.020 4.460 1.010 ;
        RECT 4.240 -1.310 4.470 -1.020 ;
        RECT 4.270 -2.600 4.460 -1.310 ;
        RECT 4.250 -2.890 4.480 -2.600 ;
        RECT 4.270 -3.820 4.460 -2.890 ;
    END
  END PROGGATE
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT -0.920 -0.740 -0.730 -0.340 ;
        RECT -1.110 -0.750 -0.730 -0.740 ;
        RECT -1.110 -0.930 2.630 -0.750 ;
        RECT -1.110 -0.970 -0.730 -0.930 ;
        RECT -0.920 -1.350 -0.730 -0.970 ;
      LAYER mcon ;
        RECT -1.100 -0.940 -0.930 -0.770 ;
      LAYER met1 ;
        RECT -1.130 -3.820 -0.900 2.230 ;
    END
  END VGND
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 2.516100 ;
    PORT
      LAYER nwell ;
        RECT -3.950 1.480 -2.220 2.230 ;
        RECT -3.950 -2.090 -2.210 1.480 ;
        RECT -3.950 -3.810 -2.220 -2.090 ;
      LAYER li1 ;
        RECT -3.520 0.090 -2.970 0.520 ;
        RECT -3.520 -1.640 -2.970 -1.210 ;
      LAYER mcon ;
        RECT -3.520 0.170 -3.250 0.440 ;
        RECT -3.520 -1.560 -3.250 -1.290 ;
      LAYER met1 ;
        RECT -3.610 -3.820 -3.190 2.230 ;
    END
  END VTUN
  PIN DRAIN
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER li1 ;
        RECT 5.410 -1.520 5.580 -1.160 ;
        RECT 5.410 -1.560 5.820 -1.520 ;
        RECT 5.410 -1.750 5.830 -1.560 ;
        RECT 5.410 -1.780 5.820 -1.750 ;
        RECT 5.410 -2.850 5.580 -1.780 ;
      LAYER mcon ;
        RECT 5.560 -1.740 5.730 -1.570 ;
      LAYER met1 ;
        RECT 5.490 -1.810 5.810 -1.490 ;
      LAYER via ;
        RECT 5.520 -1.780 5.780 -1.520 ;
      LAYER met2 ;
        RECT 5.490 -1.670 5.800 -1.480 ;
        RECT -3.950 -1.810 5.800 -1.670 ;
        RECT -3.950 -1.860 5.770 -1.810 ;
    END
  END DRAIN
  PIN VS
    USE ANALOG ;
    ANTENNADIFFAREA 1.030400 ;
    PORT
      LAYER li1 ;
        RECT 6.240 -0.340 6.410 1.270 ;
        RECT 6.240 -0.530 6.420 -0.340 ;
        RECT 6.240 -1.250 6.420 -1.060 ;
        RECT 6.240 -2.860 6.410 -1.250 ;
      LAYER met1 ;
        RECT 6.210 -0.630 6.450 -0.210 ;
        RECT 6.210 -0.950 6.480 -0.630 ;
        RECT 6.210 -1.380 6.450 -0.950 ;
      LAYER via ;
        RECT 6.220 -0.920 6.480 -0.660 ;
      LAYER met2 ;
        RECT 6.190 -0.690 6.510 -0.660 ;
        RECT -3.950 -0.920 6.510 -0.690 ;
    END
  END VS
  OBS
      LAYER nwell ;
        RECT -0.190 -0.160 2.530 1.490 ;
        RECT -0.180 -0.200 2.530 -0.160 ;
        RECT -0.180 -1.530 2.530 -1.490 ;
        RECT -0.190 -3.180 2.530 -1.530 ;
      LAYER li1 ;
        RECT 2.000 0.450 2.230 0.970 ;
        RECT 2.000 0.280 4.990 0.450 ;
        RECT 2.060 -1.970 4.990 -1.870 ;
        RECT 2.000 -2.040 4.990 -1.970 ;
        RECT 2.000 -2.660 2.230 -2.040 ;
      LAYER mcon ;
        RECT 2.030 0.770 2.200 0.940 ;
        RECT 2.030 0.320 2.200 0.490 ;
        RECT 2.030 -2.180 2.200 -2.010 ;
        RECT 2.030 -2.630 2.200 -2.460 ;
      LAYER met1 ;
        RECT 1.990 0.230 2.250 1.020 ;
        RECT 1.990 -2.710 2.250 -1.920 ;
  END
END sky130_hilas_FGtrans2x1cell

MACRO sky130_hilas_TgateDouble01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TgateDouble01 ;
  ORIGIN 2.630 1.810 ;
  SIZE 7.080 BY 1.520 ;
  OBS
      LAYER nwell ;
        RECT -2.510 -1.810 0.960 -0.290 ;
      LAYER li1 ;
        RECT -2.390 -0.830 -2.180 -0.400 ;
        RECT -1.880 -0.710 -1.690 -0.680 ;
        RECT 3.940 -0.700 4.130 -0.680 ;
        RECT -2.370 -0.850 -2.200 -0.830 ;
        RECT -1.880 -0.880 -1.360 -0.710 ;
        RECT -1.010 -0.880 3.210 -0.700 ;
        RECT 3.590 -0.710 4.130 -0.700 ;
        RECT 3.590 -0.870 4.370 -0.710 ;
        RECT -1.880 -0.960 -1.690 -0.880 ;
        RECT -1.900 -0.990 -1.690 -0.960 ;
        RECT -1.910 -1.000 -1.690 -0.990 ;
        RECT -0.520 -1.000 -0.190 -0.880 ;
        RECT 3.940 -0.910 4.370 -0.870 ;
        RECT -2.030 -1.050 -1.690 -1.000 ;
        RECT -2.160 -1.080 -1.690 -1.050 ;
        RECT -2.200 -1.110 -1.690 -1.080 ;
        RECT -1.520 -1.090 -1.200 -1.050 ;
        RECT -2.200 -1.170 -1.710 -1.110 ;
        RECT -2.200 -1.220 -1.860 -1.170 ;
        RECT -2.200 -1.240 -1.940 -1.220 ;
        RECT -2.200 -1.260 -1.970 -1.240 ;
        RECT -2.200 -1.300 -1.990 -1.260 ;
        RECT -1.520 -1.280 -1.190 -1.090 ;
        RECT -0.910 -1.100 -0.720 -1.090 ;
        RECT -2.200 -1.580 -2.030 -1.300 ;
        RECT -1.520 -1.310 -1.200 -1.280 ;
        RECT -1.520 -1.340 -1.340 -1.310 ;
        RECT -1.690 -1.510 -1.340 -1.340 ;
        RECT -0.920 -1.320 -0.720 -1.100 ;
        RECT -0.920 -1.590 -0.750 -1.320 ;
        RECT -0.140 -1.420 0.030 -1.250 ;
        RECT 0.540 -1.300 0.730 -1.070 ;
        RECT 1.400 -1.090 1.720 -1.050 ;
        RECT 1.400 -1.280 1.730 -1.090 ;
        RECT -0.170 -1.460 0.150 -1.420 ;
        RECT -0.170 -1.650 0.160 -1.460 ;
        RECT 0.550 -1.590 0.720 -1.300 ;
        RECT 1.400 -1.310 1.720 -1.280 ;
        RECT 2.250 -1.310 2.440 -1.080 ;
        RECT 1.510 -1.590 1.680 -1.310 ;
        RECT 2.250 -1.600 2.420 -1.310 ;
        RECT 2.970 -1.410 3.140 -1.250 ;
        RECT 3.480 -1.330 3.670 -1.300 ;
        RECT 2.910 -1.450 3.230 -1.410 ;
        RECT 2.910 -1.640 3.240 -1.450 ;
        RECT 3.480 -1.500 3.920 -1.330 ;
        RECT 3.480 -1.530 3.670 -1.500 ;
        RECT 4.200 -1.590 4.370 -0.910 ;
        RECT -0.170 -1.680 0.150 -1.650 ;
        RECT 2.910 -1.670 3.230 -1.640 ;
      LAYER mcon ;
        RECT -1.870 -0.880 -1.700 -0.710 ;
        RECT 3.950 -0.880 4.120 -0.710 ;
        RECT -1.460 -1.270 -1.290 -1.100 ;
        RECT -0.900 -1.290 -0.730 -1.120 ;
        RECT 0.550 -1.270 0.720 -1.100 ;
        RECT 1.460 -1.270 1.630 -1.100 ;
        RECT 2.260 -1.280 2.430 -1.110 ;
        RECT -0.110 -1.640 0.060 -1.470 ;
        RECT 2.970 -1.630 3.140 -1.460 ;
        RECT 3.490 -1.500 3.660 -1.330 ;
      LAYER met1 ;
        RECT -2.390 -0.620 -2.050 -0.400 ;
        RECT -2.400 -0.720 -2.050 -0.620 ;
        RECT -1.890 -0.650 -1.690 -0.290 ;
        RECT -2.400 -0.910 -2.170 -0.720 ;
        RECT -1.900 -0.940 -1.670 -0.650 ;
        RECT -0.920 -0.800 -0.660 -0.480 ;
        RECT 0.500 -0.790 0.760 -0.470 ;
        RECT 2.250 -0.770 2.510 -0.450 ;
        RECT 3.290 -0.530 3.550 -0.460 ;
        RECT -1.890 -1.810 -1.690 -0.940 ;
        RECT -1.530 -1.340 -1.210 -1.020 ;
        RECT -0.910 -1.060 -0.740 -0.800 ;
        RECT 0.540 -1.040 0.710 -0.790 ;
        RECT -0.930 -1.350 -0.700 -1.060 ;
        RECT 0.520 -1.330 0.750 -1.040 ;
        RECT 1.390 -1.340 1.710 -1.020 ;
        RECT 2.260 -1.050 2.430 -0.770 ;
        RECT 3.290 -0.780 3.650 -0.530 ;
        RECT 3.940 -0.650 4.130 -0.290 ;
        RECT 2.230 -1.340 2.460 -1.050 ;
        RECT 3.460 -1.270 3.650 -0.780 ;
        RECT 3.920 -0.940 4.150 -0.650 ;
        RECT -0.180 -1.710 0.140 -1.390 ;
        RECT 2.900 -1.700 3.220 -1.380 ;
        RECT 3.460 -1.560 3.690 -1.270 ;
        RECT 3.940 -1.810 4.130 -0.940 ;
      LAYER via ;
        RECT -2.310 -0.690 -2.050 -0.430 ;
        RECT -0.920 -0.770 -0.660 -0.510 ;
        RECT 0.500 -0.760 0.760 -0.500 ;
        RECT 2.250 -0.740 2.510 -0.480 ;
        RECT 3.290 -0.750 3.550 -0.490 ;
        RECT -1.500 -1.310 -1.240 -1.050 ;
        RECT 1.420 -1.310 1.680 -1.050 ;
        RECT -0.150 -1.680 0.110 -1.420 ;
        RECT 2.930 -1.670 3.190 -1.410 ;
      LAYER met2 ;
        RECT -2.340 -0.520 -2.020 -0.430 ;
        RECT -2.630 -0.720 -2.020 -0.520 ;
        RECT -0.950 -0.520 -0.630 -0.510 ;
        RECT 0.470 -0.520 0.790 -0.500 ;
        RECT 2.220 -0.520 2.540 -0.480 ;
        RECT 3.260 -0.520 3.580 -0.490 ;
        RECT -0.950 -0.720 4.450 -0.520 ;
        RECT -0.950 -0.770 -0.630 -0.720 ;
        RECT 0.470 -0.760 0.790 -0.720 ;
        RECT 2.220 -0.740 2.540 -0.720 ;
        RECT 3.260 -0.750 3.580 -0.720 ;
        RECT -1.530 -1.020 -1.220 -1.010 ;
        RECT 1.390 -1.020 1.700 -1.010 ;
        RECT -2.630 -1.220 1.740 -1.020 ;
        RECT -1.530 -1.340 -1.220 -1.220 ;
        RECT 1.390 -1.340 1.700 -1.220 ;
        RECT -0.180 -1.500 0.130 -1.380 ;
        RECT 2.900 -1.500 3.210 -1.370 ;
        RECT -2.630 -1.700 3.210 -1.500 ;
        RECT -0.180 -1.710 0.130 -1.700 ;
  END
END sky130_hilas_TgateDouble01

MACRO sky130_hilas_capacitorSize02
  CLASS BLOCK ;
  FOREIGN sky130_hilas_capacitorSize02 ;
  ORIGIN -14.140 0.480 ;
  SIZE 7.970 BY 5.830 ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 21.500 2.620 21.870 2.680 ;
        RECT 21.500 2.340 22.110 2.620 ;
        RECT 21.500 2.280 21.870 2.340 ;
      LAYER via2 ;
        RECT 21.550 2.340 21.830 2.620 ;
      LAYER met3 ;
        RECT 15.600 5.320 17.910 5.350 ;
        RECT 15.600 2.830 19.830 5.320 ;
        RECT 15.600 2.080 22.070 2.830 ;
        RECT 15.600 -0.460 19.830 2.080 ;
        RECT 17.880 -0.480 19.830 -0.460 ;
      LAYER via3 ;
        RECT 21.470 2.230 21.900 2.710 ;
      LAYER met4 ;
        RECT 21.370 2.140 22.030 2.800 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 14.380 2.600 14.750 2.660 ;
        RECT 14.160 2.320 14.750 2.600 ;
        RECT 14.380 2.260 14.750 2.320 ;
      LAYER via2 ;
        RECT 14.430 2.320 14.710 2.600 ;
      LAYER met3 ;
        RECT 14.160 2.060 14.950 2.810 ;
      LAYER via3 ;
        RECT 14.350 2.210 14.780 2.690 ;
      LAYER met4 ;
        RECT 14.250 2.720 14.910 2.780 ;
        RECT 15.300 2.720 16.310 2.730 ;
        RECT 14.250 2.220 17.940 2.720 ;
        RECT 14.250 2.210 15.660 2.220 ;
        RECT 14.250 2.120 14.910 2.210 ;
        RECT 17.300 1.100 17.930 2.220 ;
        RECT 17.300 1.090 19.450 1.100 ;
        RECT 15.980 0.790 19.450 1.090 ;
        RECT 15.980 0.620 18.990 0.790 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 14.140 4.800 22.110 4.980 ;
        RECT 14.140 4.370 22.110 4.550 ;
        RECT 14.170 3.370 22.110 3.550 ;
        RECT 14.170 2.940 22.110 3.120 ;
        RECT 14.170 1.790 22.110 1.960 ;
        RECT 14.170 1.370 22.110 1.540 ;
        RECT 14.170 0.390 22.110 0.560 ;
        RECT 14.170 -0.050 22.110 0.120 ;
  END
END sky130_hilas_capacitorSize02

MACRO sky130_hilas_pFETdevice01aa
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pFETdevice01aa ;
  ORIGIN 0.800 0.780 ;
  SIZE 1.720 BY 1.210 ;
  OBS
      LAYER nwell ;
        RECT -0.800 -0.780 0.810 0.430 ;
  END
END sky130_hilas_pFETdevice01aa

MACRO sky130_hilas_m12m2
  CLASS BLOCK ;
  FOREIGN sky130_hilas_m12m2 ;
  ORIGIN 0.090 0.100 ;
  SIZE 0.320 BY 0.320 ;
  OBS
      LAYER met1 ;
        RECT -0.060 -0.100 0.200 0.220 ;
      LAYER via ;
        RECT -0.060 -0.070 0.200 0.190 ;
      LAYER met2 ;
        RECT -0.090 -0.070 0.230 0.190 ;
  END
END sky130_hilas_m12m2

MACRO sky130_hilas_wellContact
  CLASS BLOCK ;
  FOREIGN sky130_hilas_wellContact ;
  ORIGIN 14.490 4.410 ;
  SIZE 1.740 BY 1.860 ;
  OBS
      LAYER nwell ;
        RECT -14.490 -4.400 -12.750 -2.560 ;
      LAYER li1 ;
        RECT -14.060 -3.950 -13.510 -3.520 ;
      LAYER mcon ;
        RECT -14.060 -3.870 -13.790 -3.600 ;
      LAYER met1 ;
        RECT -14.120 -4.410 -13.730 -2.550 ;
  END
END sky130_hilas_wellContact

MACRO sky130_hilas_DAC6TransistorStack01b
  CLASS BLOCK ;
  FOREIGN sky130_hilas_DAC6TransistorStack01b ;
  ORIGIN -0.150 1.740 ;
  SIZE 1.850 BY 5.650 ;
  OBS
      LAYER nwell ;
        RECT 0.280 -1.740 1.890 3.910 ;
      LAYER li1 ;
        RECT 0.660 2.360 0.830 2.690 ;
        RECT 1.340 2.360 1.510 2.690 ;
        RECT 0.210 1.450 0.420 1.880 ;
        RECT 0.230 1.430 0.400 1.450 ;
        RECT 0.660 1.400 0.830 1.730 ;
        RECT 1.340 1.400 1.510 1.730 ;
        RECT 1.740 0.970 1.910 0.990 ;
        RECT 0.660 0.440 0.830 0.770 ;
        RECT 1.340 0.440 1.510 0.770 ;
        RECT 1.720 0.540 1.930 0.970 ;
        RECT 0.660 -0.520 0.830 -0.190 ;
        RECT 1.340 -0.520 1.510 -0.190 ;
      LAYER mcon ;
        RECT 1.740 0.820 1.910 0.990 ;
      LAYER met1 ;
        RECT 0.210 1.660 0.430 1.880 ;
        RECT 0.200 1.370 0.430 1.660 ;
        RECT 1.710 0.760 1.940 1.050 ;
        RECT 1.720 0.540 1.940 0.760 ;
  END
END sky130_hilas_DAC6TransistorStack01b

MACRO sky130_hilas_WTA4Stage01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_WTA4Stage01 ;
  ORIGIN 11.210 0.430 ;
  SIZE 14.170 BY 6.050 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 2.430 4.110 2.940 4.780 ;
        RECT 2.430 2.970 2.940 3.640 ;
        RECT 2.430 1.340 2.940 2.010 ;
        RECT 2.430 0.200 2.940 0.870 ;
      LAYER mcon ;
        RECT 2.600 4.360 2.770 4.530 ;
        RECT 2.600 3.220 2.770 3.390 ;
        RECT 2.600 1.590 2.770 1.760 ;
        RECT 2.600 0.450 2.770 0.620 ;
      LAYER met1 ;
        RECT 2.570 -0.430 2.800 5.620 ;
    END
  END VGND
  PIN COMMONNODE
    USE ANALOG ;
    ANTENNAGATEAREA 0.472000 ;
    ANTENNADIFFAREA 0.708000 ;
    PORT
      LAYER li1 ;
        RECT 1.220 4.530 1.550 4.700 ;
        RECT 1.300 4.360 1.470 4.530 ;
        RECT 1.220 4.190 1.550 4.360 ;
        RECT 1.300 3.960 1.550 4.190 ;
        RECT 1.300 3.790 1.970 3.960 ;
        RECT 1.300 3.560 1.550 3.790 ;
        RECT 1.220 3.390 1.550 3.560 ;
        RECT 1.300 3.220 1.470 3.390 ;
        RECT 1.220 3.050 1.550 3.220 ;
        RECT 1.220 1.760 1.550 1.930 ;
        RECT 1.300 1.590 1.470 1.760 ;
        RECT 1.220 1.420 1.550 1.590 ;
        RECT 1.300 1.190 1.550 1.420 ;
        RECT 1.300 1.020 1.970 1.190 ;
        RECT 1.300 0.790 1.550 1.020 ;
        RECT 1.220 0.620 1.550 0.790 ;
        RECT 1.300 0.450 1.470 0.620 ;
        RECT 1.220 0.280 1.550 0.450 ;
      LAYER mcon ;
        RECT 1.340 3.790 1.510 3.960 ;
        RECT 1.340 1.020 1.510 1.190 ;
      LAYER met1 ;
        RECT 1.310 -0.430 1.540 5.620 ;
    END
  END COMMONNODE
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.258100 ;
    PORT
      LAYER li1 ;
        RECT -8.470 4.630 -8.150 4.670 ;
        RECT -8.480 4.590 -8.150 4.630 ;
        RECT -8.730 4.420 -8.150 4.590 ;
        RECT 0.710 4.450 1.050 4.700 ;
        RECT -8.470 4.410 -8.150 4.420 ;
        RECT 0.390 4.190 1.050 4.450 ;
      LAYER mcon ;
        RECT -8.380 4.450 -8.210 4.620 ;
        RECT 0.450 4.240 0.620 4.410 ;
      LAYER met1 ;
        RECT -8.460 4.380 -8.140 4.700 ;
        RECT 0.380 4.160 0.700 4.480 ;
      LAYER via ;
        RECT -8.430 4.410 -8.170 4.670 ;
        RECT 0.410 4.190 0.670 4.450 ;
      LAYER met2 ;
        RECT -8.450 4.690 -8.140 4.710 ;
        RECT -10.610 4.660 -0.530 4.690 ;
        RECT -10.610 4.570 -0.500 4.660 ;
        RECT -10.610 4.510 0.560 4.570 ;
        RECT -8.450 4.380 -8.140 4.510 ;
        RECT -0.680 4.500 0.560 4.510 ;
        RECT -0.650 4.480 0.560 4.500 ;
        RECT -0.650 4.420 0.690 4.480 ;
        RECT -0.650 4.370 2.960 4.420 ;
        RECT 0.380 4.260 2.960 4.370 ;
        RECT 0.380 4.150 0.690 4.260 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.258100 ;
    PORT
      LAYER li1 ;
        RECT -8.470 3.780 -8.150 3.790 ;
        RECT -8.730 3.610 -8.150 3.780 ;
        RECT -8.480 3.570 -8.150 3.610 ;
        RECT -8.470 3.530 -8.150 3.570 ;
        RECT 0.390 3.300 1.050 3.560 ;
        RECT 0.710 3.050 1.050 3.300 ;
      LAYER mcon ;
        RECT -8.380 3.580 -8.210 3.750 ;
        RECT 0.450 3.340 0.620 3.510 ;
      LAYER met1 ;
        RECT -8.460 3.500 -8.140 3.820 ;
        RECT 0.380 3.270 0.700 3.590 ;
      LAYER via ;
        RECT -8.430 3.530 -8.170 3.790 ;
        RECT 0.410 3.300 0.670 3.560 ;
      LAYER met2 ;
        RECT -8.450 3.690 -8.140 3.820 ;
        RECT -0.650 3.690 0.660 3.710 ;
        RECT -10.620 3.600 0.660 3.690 ;
        RECT -10.620 3.510 0.690 3.600 ;
        RECT -8.450 3.490 -8.140 3.510 ;
        RECT 0.380 3.490 0.690 3.510 ;
        RECT 0.380 3.330 2.960 3.490 ;
        RECT 0.380 3.270 0.690 3.330 ;
    END
  END OUTPUT2
  PIN OUTPUT3
    USE ANALOG ;
    ANTENNADIFFAREA 0.258100 ;
    PORT
      LAYER li1 ;
        RECT 0.710 1.680 1.050 1.930 ;
        RECT -8.470 1.620 -8.150 1.660 ;
        RECT -8.480 1.580 -8.150 1.620 ;
        RECT -8.730 1.410 -8.150 1.580 ;
        RECT 0.390 1.420 1.050 1.680 ;
        RECT -8.470 1.400 -8.150 1.410 ;
      LAYER mcon ;
        RECT -8.380 1.440 -8.210 1.610 ;
        RECT 0.450 1.470 0.620 1.640 ;
      LAYER met1 ;
        RECT -8.460 1.370 -8.140 1.690 ;
        RECT 0.380 1.390 0.700 1.710 ;
      LAYER via ;
        RECT -8.430 1.400 -8.170 1.660 ;
        RECT 0.410 1.420 0.670 1.680 ;
      LAYER met2 ;
        RECT -8.450 1.680 -8.140 1.700 ;
        RECT 0.380 1.680 0.690 1.710 ;
        RECT -10.610 1.650 0.690 1.680 ;
        RECT -10.610 1.520 2.960 1.650 ;
        RECT -10.610 1.510 -0.550 1.520 ;
        RECT -10.610 1.500 -8.050 1.510 ;
        RECT -8.450 1.370 -8.140 1.500 ;
        RECT 0.380 1.490 2.960 1.520 ;
        RECT 0.380 1.380 0.690 1.490 ;
    END
  END OUTPUT3
  PIN OUTPUT4
    USE ANALOG ;
    ANTENNADIFFAREA 0.258100 ;
    PORT
      LAYER li1 ;
        RECT -8.470 0.780 -8.150 0.790 ;
        RECT -8.730 0.610 -8.150 0.780 ;
        RECT -8.480 0.570 -8.150 0.610 ;
        RECT -8.470 0.530 -8.150 0.570 ;
        RECT 0.390 0.530 1.050 0.790 ;
        RECT 0.710 0.280 1.050 0.530 ;
      LAYER mcon ;
        RECT -8.380 0.580 -8.210 0.750 ;
        RECT 0.450 0.570 0.620 0.740 ;
      LAYER met1 ;
        RECT -8.460 0.500 -8.140 0.820 ;
        RECT 0.380 0.500 0.700 0.820 ;
      LAYER via ;
        RECT -8.430 0.530 -8.170 0.790 ;
        RECT 0.410 0.530 0.670 0.790 ;
      LAYER met2 ;
        RECT -8.450 0.700 -8.140 0.820 ;
        RECT 0.380 0.720 0.690 0.830 ;
        RECT 0.380 0.710 2.960 0.720 ;
        RECT -0.550 0.700 2.960 0.710 ;
        RECT -8.450 0.690 2.960 0.700 ;
        RECT -10.610 0.560 2.960 0.690 ;
        RECT -10.610 0.530 0.690 0.560 ;
        RECT -10.610 0.510 -8.050 0.530 ;
        RECT -8.450 0.490 -8.140 0.510 ;
        RECT -2.870 0.440 -1.330 0.530 ;
        RECT 0.380 0.500 0.690 0.530 ;
    END
  END OUTPUT4
  PIN INPUT1
    USE ANALOG ;
    ANTENNAGATEAREA 0.118000 ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER li1 ;
        RECT 0.240 5.100 0.560 5.130 ;
        RECT 0.240 4.930 2.030 5.100 ;
        RECT 0.240 4.910 0.570 4.930 ;
        RECT 0.240 4.870 0.560 4.910 ;
        RECT 1.860 4.700 2.030 4.930 ;
        RECT 1.770 4.530 2.110 4.700 ;
        RECT 1.860 4.360 2.030 4.530 ;
        RECT 1.770 4.190 2.110 4.360 ;
      LAYER mcon ;
        RECT 0.300 4.920 0.470 5.090 ;
      LAYER met1 ;
        RECT -7.620 5.050 -7.310 5.370 ;
        RECT -7.620 4.310 -7.400 5.050 ;
        RECT 0.230 4.840 0.550 5.160 ;
        RECT -7.720 3.990 -7.400 4.310 ;
      LAYER via ;
        RECT -7.570 5.080 -7.310 5.340 ;
        RECT 0.260 4.870 0.520 5.130 ;
        RECT -7.720 4.020 -7.460 4.280 ;
      LAYER met2 ;
        RECT -7.600 5.310 -7.280 5.340 ;
        RECT -7.600 5.120 0.070 5.310 ;
        RECT 0.230 5.120 0.540 5.160 ;
        RECT -7.600 5.100 0.540 5.120 ;
        RECT -7.600 5.080 -7.280 5.100 ;
        RECT -0.140 4.910 0.540 5.100 ;
        RECT 0.230 4.830 0.540 4.910 ;
        RECT -11.120 4.180 -10.970 4.690 ;
        RECT -7.750 4.180 -7.430 4.280 ;
        RECT -11.120 4.020 -7.430 4.180 ;
    END
  END INPUT1
  PIN INPUT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.118000 ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER li1 ;
        RECT 1.770 3.390 2.110 3.560 ;
        RECT 1.860 3.220 2.030 3.390 ;
        RECT 1.770 3.050 2.110 3.220 ;
        RECT 0.240 2.840 0.560 2.880 ;
        RECT 0.240 2.820 0.570 2.840 ;
        RECT 1.860 2.820 2.030 3.050 ;
        RECT 0.240 2.650 2.030 2.820 ;
        RECT 0.240 2.620 0.560 2.650 ;
      LAYER mcon ;
        RECT 0.300 2.660 0.470 2.830 ;
      LAYER met1 ;
        RECT -11.110 3.690 -10.850 3.810 ;
        RECT -11.120 3.490 -10.850 3.690 ;
        RECT -11.120 2.800 -10.910 3.490 ;
        RECT -11.130 2.480 -10.870 2.800 ;
        RECT 0.230 2.590 0.550 2.910 ;
      LAYER via ;
        RECT -11.110 3.520 -10.850 3.780 ;
        RECT -11.130 2.510 -10.870 2.770 ;
        RECT 0.260 2.620 0.520 2.880 ;
      LAYER met2 ;
        RECT -11.140 3.520 -10.820 3.780 ;
        RECT -11.070 3.510 -10.900 3.520 ;
        RECT -7.910 3.040 -7.680 3.050 ;
        RECT -7.910 3.010 -0.340 3.040 ;
        RECT -7.910 2.840 -0.280 3.010 ;
        RECT 0.230 2.840 0.540 2.920 ;
        RECT -11.160 2.740 -10.840 2.770 ;
        RECT -7.910 2.740 -7.670 2.840 ;
        RECT -11.160 2.560 -7.670 2.740 ;
        RECT -0.470 2.640 0.540 2.840 ;
        RECT 0.130 2.630 0.540 2.640 ;
        RECT 0.230 2.590 0.540 2.630 ;
        RECT -11.160 2.540 -7.750 2.560 ;
        RECT -11.160 2.510 -10.840 2.540 ;
    END
  END INPUT2
  PIN INPUT3
    USE ANALOG ;
    ANTENNAGATEAREA 0.118000 ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER li1 ;
        RECT 0.240 2.330 0.560 2.360 ;
        RECT 0.240 2.160 2.030 2.330 ;
        RECT 0.240 2.140 0.570 2.160 ;
        RECT 0.240 2.100 0.560 2.140 ;
        RECT 1.860 1.930 2.030 2.160 ;
        RECT 1.770 1.760 2.110 1.930 ;
        RECT 1.860 1.590 2.030 1.760 ;
        RECT 1.770 1.420 2.110 1.590 ;
      LAYER mcon ;
        RECT 0.300 2.150 0.470 2.320 ;
      LAYER met1 ;
        RECT -7.730 2.120 -7.470 2.420 ;
        RECT -7.730 2.100 -7.450 2.120 ;
        RECT -7.720 1.220 -7.450 2.100 ;
        RECT 0.230 2.070 0.550 2.390 ;
        RECT -7.710 0.930 -7.450 1.220 ;
      LAYER via ;
        RECT -7.730 2.130 -7.470 2.390 ;
        RECT 0.260 2.100 0.520 2.360 ;
        RECT -7.710 0.960 -7.450 1.220 ;
      LAYER met2 ;
        RECT -7.760 2.360 -7.440 2.390 ;
        RECT -7.760 2.340 -0.320 2.360 ;
        RECT 0.230 2.350 0.540 2.390 ;
        RECT 0.130 2.340 0.540 2.350 ;
        RECT -7.760 2.140 0.540 2.340 ;
        RECT -7.760 2.130 -7.440 2.140 ;
        RECT 0.230 2.060 0.540 2.140 ;
        RECT -11.180 1.180 -10.980 1.680 ;
        RECT -7.740 1.180 -7.420 1.220 ;
        RECT -11.180 0.980 -7.420 1.180 ;
        RECT -7.740 0.960 -7.420 0.980 ;
    END
  END INPUT3
  PIN INPUT4
    USE ANALOG ;
    ANTENNAGATEAREA 0.118000 ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER li1 ;
        RECT -11.200 0.690 -10.880 0.730 ;
        RECT -11.200 0.500 -10.870 0.690 ;
        RECT 1.770 0.620 2.110 0.790 ;
        RECT -11.200 0.470 -10.880 0.500 ;
        RECT -11.150 -0.120 -10.970 0.470 ;
        RECT 1.860 0.450 2.030 0.620 ;
        RECT 1.770 0.280 2.110 0.450 ;
        RECT 0.240 0.070 0.560 0.110 ;
        RECT 0.240 0.050 0.570 0.070 ;
        RECT 1.860 0.050 2.030 0.280 ;
        RECT 0.240 -0.120 2.030 0.050 ;
        RECT -11.150 -0.160 -10.830 -0.120 ;
        RECT 0.240 -0.150 0.560 -0.120 ;
        RECT -11.150 -0.350 -10.820 -0.160 ;
        RECT -11.150 -0.380 -10.830 -0.350 ;
      LAYER mcon ;
        RECT -11.140 0.510 -10.970 0.680 ;
        RECT 0.300 -0.110 0.470 0.060 ;
        RECT -11.090 -0.340 -10.920 -0.170 ;
      LAYER met1 ;
        RECT -11.210 0.440 -10.890 0.760 ;
        RECT -11.160 -0.410 -10.840 -0.090 ;
        RECT 0.230 -0.180 0.550 0.140 ;
      LAYER via ;
        RECT -11.180 0.470 -10.920 0.730 ;
        RECT -11.130 -0.380 -10.870 -0.120 ;
        RECT 0.260 -0.150 0.520 0.110 ;
      LAYER met2 ;
        RECT -11.210 0.440 -10.900 0.770 ;
        RECT 0.230 0.090 0.540 0.150 ;
        RECT -0.320 0.080 0.540 0.090 ;
        RECT -11.160 -0.200 -10.850 -0.080 ;
        RECT -7.900 -0.140 0.540 0.080 ;
        RECT -7.900 -0.150 -0.310 -0.140 ;
        RECT -7.900 -0.160 -7.130 -0.150 ;
        RECT -7.900 -0.200 -7.660 -0.160 ;
        RECT 0.230 -0.180 0.540 -0.140 ;
        RECT -11.160 -0.400 -7.660 -0.200 ;
        RECT -11.160 -0.410 -8.470 -0.400 ;
    END
  END INPUT4
  OBS
      LAYER nwell ;
        RECT -11.010 3.690 -8.050 5.620 ;
        RECT -11.120 2.540 -8.050 3.690 ;
        RECT -11.010 -0.420 -8.050 2.540 ;
        RECT -6.520 -0.430 -4.290 5.620 ;
        RECT -2.270 4.990 -0.540 5.620 ;
        RECT -2.270 1.920 -0.530 4.990 ;
        RECT -2.270 -0.430 -0.540 1.920 ;
      LAYER li1 ;
        RECT -10.210 4.940 -10.010 5.290 ;
        RECT -8.470 5.210 -8.150 5.220 ;
        RECT -8.730 5.040 -8.150 5.210 ;
        RECT -8.480 4.990 -8.150 5.040 ;
        RECT -8.470 4.960 -8.150 4.990 ;
        RECT -10.220 4.910 -10.010 4.940 ;
        RECT -10.220 4.320 -10.000 4.910 ;
        RECT -9.480 4.350 -9.280 4.920 ;
        RECT -10.220 3.290 -10.000 3.880 ;
        RECT -10.220 3.260 -10.010 3.290 ;
        RECT -9.480 3.280 -9.280 3.850 ;
        RECT -10.210 2.910 -10.010 3.260 ;
        RECT -8.470 3.210 -8.150 3.240 ;
        RECT -8.480 3.160 -8.150 3.210 ;
        RECT -8.730 2.990 -8.150 3.160 ;
        RECT -8.470 2.980 -8.150 2.990 ;
        RECT -9.840 2.510 -9.400 2.680 ;
        RECT -5.540 2.300 -4.990 2.730 ;
        RECT -1.510 2.370 -0.960 2.800 ;
        RECT -10.210 1.930 -10.010 2.280 ;
        RECT -8.470 2.200 -8.150 2.210 ;
        RECT -8.730 2.030 -8.150 2.200 ;
        RECT -8.480 1.980 -8.150 2.030 ;
        RECT -8.470 1.950 -8.150 1.980 ;
        RECT -10.220 1.900 -10.010 1.930 ;
        RECT -10.220 1.310 -10.000 1.900 ;
        RECT -9.480 1.340 -9.280 1.910 ;
        RECT -10.220 0.290 -10.000 0.880 ;
        RECT -10.220 0.260 -10.010 0.290 ;
        RECT -9.480 0.280 -9.280 0.850 ;
        RECT -10.210 -0.090 -10.010 0.260 ;
        RECT -8.470 0.210 -8.150 0.240 ;
        RECT -8.480 0.160 -8.150 0.210 ;
        RECT -8.730 -0.010 -8.150 0.160 ;
        RECT -8.470 -0.020 -8.150 -0.010 ;
      LAYER mcon ;
        RECT -8.380 5.000 -8.210 5.170 ;
        RECT -10.190 4.740 -10.020 4.910 ;
        RECT -9.460 4.710 -9.290 4.880 ;
        RECT -10.190 3.290 -10.020 3.460 ;
        RECT -9.460 3.320 -9.290 3.490 ;
        RECT -8.380 3.030 -8.210 3.200 ;
        RECT -5.260 2.380 -4.990 2.650 ;
        RECT -1.230 2.450 -0.960 2.720 ;
        RECT -8.380 1.990 -8.210 2.160 ;
        RECT -10.190 1.730 -10.020 1.900 ;
        RECT -9.460 1.700 -9.290 1.870 ;
        RECT -10.190 0.290 -10.020 0.460 ;
        RECT -9.460 0.320 -9.290 0.490 ;
        RECT -8.380 0.030 -8.210 0.200 ;
      LAYER met1 ;
        RECT -10.250 4.970 -10.090 5.620 ;
        RECT -10.250 4.420 -9.980 4.970 ;
        RECT -10.260 4.370 -9.980 4.420 ;
        RECT -9.840 4.630 -9.650 5.620 ;
        RECT -9.440 4.940 -9.280 5.620 ;
        RECT -9.480 4.920 -9.280 4.940 ;
        RECT -8.460 4.930 -8.140 5.250 ;
        RECT -9.490 4.680 -9.260 4.920 ;
        RECT -9.840 4.510 -9.670 4.630 ;
        RECT -10.260 4.280 -10.090 4.370 ;
        RECT -10.250 3.920 -10.090 4.280 ;
        RECT -10.260 3.830 -10.090 3.920 ;
        RECT -10.260 3.780 -9.980 3.830 ;
        RECT -10.250 3.230 -9.980 3.780 ;
        RECT -9.840 3.690 -9.680 4.510 ;
        RECT -9.480 4.460 -9.280 4.680 ;
        RECT -9.440 3.740 -9.280 4.460 ;
        RECT -9.840 3.570 -9.670 3.690 ;
        RECT -10.250 1.960 -10.090 3.230 ;
        RECT -9.840 2.710 -9.650 3.570 ;
        RECT -9.480 3.520 -9.280 3.740 ;
        RECT -5.320 3.700 -4.940 5.620 ;
        RECT -9.490 3.280 -9.260 3.520 ;
        RECT -9.480 3.260 -9.280 3.280 ;
        RECT -9.870 2.480 -9.630 2.710 ;
        RECT -10.250 1.410 -9.980 1.960 ;
        RECT -10.260 1.360 -9.980 1.410 ;
        RECT -9.840 1.620 -9.650 2.480 ;
        RECT -9.440 1.930 -9.280 3.260 ;
        RECT -8.460 2.950 -8.140 3.270 ;
        RECT -9.480 1.910 -9.280 1.930 ;
        RECT -8.460 1.920 -8.140 2.240 ;
        RECT -9.490 1.670 -9.260 1.910 ;
        RECT -5.320 1.840 -4.930 3.700 ;
        RECT -9.840 1.500 -9.670 1.620 ;
        RECT -10.260 1.270 -10.090 1.360 ;
        RECT -10.250 0.920 -10.090 1.270 ;
        RECT -10.260 0.830 -10.090 0.920 ;
        RECT -10.260 0.780 -9.980 0.830 ;
        RECT -10.250 0.230 -9.980 0.780 ;
        RECT -9.840 0.690 -9.680 1.500 ;
        RECT -9.480 1.450 -9.280 1.670 ;
        RECT -9.440 0.740 -9.280 1.450 ;
        RECT -9.840 0.570 -9.670 0.690 ;
        RECT -10.250 -0.420 -10.090 0.230 ;
        RECT -9.840 -0.420 -9.650 0.570 ;
        RECT -9.480 0.520 -9.280 0.740 ;
        RECT -9.490 0.280 -9.260 0.520 ;
        RECT -9.480 0.260 -9.280 0.280 ;
        RECT -9.440 -0.420 -9.280 0.260 ;
        RECT -8.460 -0.050 -8.140 0.270 ;
        RECT -5.320 -0.430 -4.940 1.840 ;
        RECT -1.290 -0.430 -0.890 5.620 ;
      LAYER via ;
        RECT -8.430 4.960 -8.170 5.220 ;
        RECT -8.430 2.980 -8.170 3.240 ;
        RECT -8.430 1.950 -8.170 2.210 ;
        RECT -8.430 -0.020 -8.170 0.240 ;
      LAYER met2 ;
        RECT -8.450 5.120 -8.140 5.260 ;
        RECT -11.000 4.940 -8.040 5.120 ;
        RECT -8.450 4.930 -8.140 4.940 ;
        RECT -8.450 3.260 -8.140 3.270 ;
        RECT -11.000 3.220 -8.140 3.260 ;
        RECT -11.000 3.080 -8.050 3.220 ;
        RECT -8.450 2.940 -8.140 3.080 ;
        RECT -8.450 2.110 -8.140 2.250 ;
        RECT -11.000 2.100 -8.140 2.110 ;
        RECT -11.000 1.930 -8.020 2.100 ;
        RECT -8.450 1.920 -8.140 1.930 ;
        RECT -8.450 0.260 -8.140 0.270 ;
        RECT -11.000 0.090 -8.040 0.260 ;
        RECT -11.000 0.080 -8.140 0.090 ;
        RECT -8.450 -0.060 -8.140 0.080 ;
  END
END sky130_hilas_WTA4Stage01

MACRO sky130_hilas_FGVaractorCapacitor
  CLASS BLOCK ;
  FOREIGN sky130_hilas_FGVaractorCapacitor ;
  ORIGIN 9.570 3.950 ;
  SIZE 2.230 BY 1.860 ;
  OBS
      LAYER nwell ;
        RECT -9.570 -3.950 -7.340 -2.100 ;
      LAYER met1 ;
        RECT -8.920 -3.950 -8.540 -2.090 ;
  END
END sky130_hilas_FGVaractorCapacitor

MACRO sky130_hilas_horizTransCell01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_horizTransCell01 ;
  ORIGIN 4.760 -0.480 ;
  SIZE 4.430 BY 3.110 ;
  OBS
      LAYER nwell ;
        RECT -3.640 0.480 -0.330 3.590 ;
      LAYER li1 ;
        RECT -4.600 3.040 -4.260 3.210 ;
        RECT -3.240 3.040 -2.910 3.210 ;
        RECT -4.610 2.250 -4.260 2.420 ;
        RECT -3.240 2.250 -2.910 2.420 ;
        RECT -4.610 1.460 -4.260 1.630 ;
        RECT -3.240 1.460 -2.910 1.630 ;
        RECT -2.490 1.440 -2.320 3.130 ;
        RECT -1.660 3.040 -1.480 3.230 ;
        RECT -1.660 1.430 -1.490 3.040 ;
        RECT -1.300 2.230 -1.060 2.560 ;
        RECT -1.290 1.940 -1.090 2.230 ;
        RECT -1.290 1.930 -1.100 1.940 ;
        RECT -0.930 1.760 -0.720 1.770 ;
        RECT -0.940 1.180 -0.720 1.760 ;
        RECT -0.930 1.150 -0.720 1.180 ;
        RECT -2.740 0.880 -2.210 1.050 ;
        RECT -0.930 0.800 -0.730 1.150 ;
      LAYER mcon ;
        RECT -1.280 2.000 -1.100 2.190 ;
        RECT -0.920 1.180 -0.750 1.350 ;
      LAYER met1 ;
        RECT -1.690 2.910 -1.450 3.290 ;
        RECT -1.260 2.480 -1.100 3.500 ;
        RECT -1.300 2.240 -1.070 2.480 ;
        RECT -1.300 2.230 -1.060 2.240 ;
        RECT -1.310 1.960 -1.060 2.230 ;
        RECT -1.290 1.930 -1.070 1.960 ;
        RECT -2.810 0.770 -2.510 1.150 ;
        RECT -1.290 0.480 -1.100 1.930 ;
        RECT -0.850 1.810 -0.690 3.500 ;
        RECT -0.850 1.720 -0.680 1.810 ;
        RECT -0.960 1.670 -0.680 1.720 ;
        RECT -0.960 1.120 -0.690 1.670 ;
        RECT -0.850 0.480 -0.690 1.120 ;
      LAYER via ;
        RECT -2.790 0.820 -2.530 1.090 ;
      LAYER met2 ;
        RECT -2.890 0.970 -0.330 1.150 ;
        RECT -2.810 0.770 -2.510 0.970 ;
  END
END sky130_hilas_horizTransCell01

MACRO sky130_hilas_CapModule01a
  CLASS BLOCK ;
  FOREIGN sky130_hilas_CapModule01a ;
  ORIGIN 4.160 2.160 ;
  SIZE 2.300 BY 2.280 ;
  OBS
      LAYER met3 ;
        RECT -4.160 -2.160 -1.860 0.120 ;
      LAYER met4 ;
        RECT -3.310 -0.930 -2.860 -0.920 ;
        RECT -3.330 -1.420 -2.810 -0.930 ;
  END
END sky130_hilas_CapModule01a

MACRO sky130_hilas_CapModule03
  CLASS BLOCK ;
  FOREIGN sky130_hilas_CapModule03 ;
  ORIGIN 3.920 2.470 ;
  SIZE 4.230 BY 5.830 ;
  OBS
      LAYER met3 ;
        RECT -3.920 3.330 -1.610 3.360 ;
        RECT -3.920 -2.450 0.310 3.330 ;
        RECT -1.640 -2.470 0.310 -2.450 ;
      LAYER met4 ;
        RECT -3.540 -1.370 -0.530 -0.900 ;
  END
END sky130_hilas_CapModule03

MACRO sky130_hilas_pFETmirror02
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pFETmirror02 ;
  ORIGIN 0.610 -0.890 ;
  SIZE 1.280 BY 2.840 ;
  OBS
      LAYER nwell ;
        RECT -0.610 0.890 0.670 3.730 ;
      LAYER li1 ;
        RECT -0.410 3.310 0.290 3.490 ;
        RECT -0.400 2.010 0.300 2.890 ;
        RECT -0.400 1.400 0.310 1.570 ;
        RECT -0.050 1.120 0.310 1.400 ;
        RECT -0.050 0.950 0.530 1.120 ;
  END
END sky130_hilas_pFETmirror02

MACRO sky130_hilas_overlapCap02a
  CLASS BLOCK ;
  FOREIGN sky130_hilas_overlapCap02a ;
  ORIGIN 5.210 0.540 ;
  SIZE 4.000 BY 1.640 ;
  OBS
      LAYER nwell ;
        RECT -5.210 -0.540 -1.210 1.100 ;
      LAYER li1 ;
        RECT -4.860 -0.210 -1.550 0.770 ;
      LAYER mcon ;
        RECT -3.290 0.540 -3.120 0.710 ;
        RECT -3.290 0.190 -3.120 0.360 ;
        RECT -3.290 -0.150 -3.120 0.020 ;
      LAYER met1 ;
        RECT -3.330 0.130 -3.090 0.770 ;
        RECT -3.320 -0.130 -3.090 0.130 ;
        RECT -3.320 -0.350 -3.080 -0.130 ;
  END
END sky130_hilas_overlapCap02a

MACRO sky130_hilas_DualTACore01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_DualTACore01 ;
  ORIGIN 1.720 0.220 ;
  SIZE 3.270 BY 5.720 ;
  OBS
      LAYER nwell ;
        RECT 0.270 -0.220 1.550 5.460 ;
      LAYER li1 ;
        RECT -1.130 5.310 -0.930 5.350 ;
        RECT -1.360 5.050 -0.930 5.310 ;
        RECT -1.130 5.020 -0.930 5.050 ;
        RECT -1.540 4.660 -1.370 4.700 ;
        RECT -1.130 4.660 -0.930 4.690 ;
        RECT -1.540 4.400 -0.930 4.660 ;
        RECT -1.540 4.370 -1.370 4.400 ;
        RECT -1.130 4.360 -0.930 4.400 ;
        RECT -0.540 4.360 0.010 5.350 ;
        RECT 0.830 5.230 1.410 5.400 ;
        RECT 0.830 5.130 1.220 5.230 ;
        RECT 0.830 5.100 1.210 5.130 ;
        RECT 0.830 4.950 1.190 5.100 ;
        RECT 0.480 4.780 1.190 4.950 ;
        RECT 0.480 4.030 1.180 4.340 ;
        RECT -1.540 3.830 -1.370 3.860 ;
        RECT -1.130 3.830 -0.930 3.870 ;
        RECT -1.540 3.570 -0.930 3.830 ;
        RECT -1.540 3.530 -1.370 3.570 ;
        RECT -1.130 3.540 -0.930 3.570 ;
        RECT -1.130 3.180 -0.930 3.210 ;
        RECT -1.360 2.920 -0.930 3.180 ;
        RECT -1.130 2.880 -0.930 2.920 ;
        RECT -0.540 2.880 0.010 3.870 ;
        RECT 0.330 3.800 1.180 4.030 ;
        RECT 0.480 3.460 1.180 3.800 ;
        RECT 0.940 3.100 1.260 3.140 ;
        RECT 0.940 3.040 1.270 3.100 ;
        RECT 0.470 2.910 1.270 3.040 ;
        RECT 0.470 2.880 1.260 2.910 ;
        RECT 0.470 2.860 1.170 2.880 ;
        RECT -1.130 2.350 -0.930 2.390 ;
        RECT -1.360 2.090 -0.930 2.350 ;
        RECT -1.130 2.060 -0.930 2.090 ;
        RECT -1.540 1.700 -1.370 1.740 ;
        RECT -1.130 1.700 -0.930 1.730 ;
        RECT -1.540 1.440 -0.930 1.700 ;
        RECT -1.540 1.410 -1.370 1.440 ;
        RECT -1.130 1.400 -0.930 1.440 ;
        RECT -0.540 1.400 0.010 2.390 ;
        RECT 0.930 2.380 1.250 2.420 ;
        RECT 0.470 2.200 1.260 2.380 ;
        RECT 0.930 2.190 1.260 2.200 ;
        RECT 0.930 2.160 1.250 2.190 ;
        RECT 0.480 1.440 1.180 1.780 ;
        RECT 0.330 1.210 1.180 1.440 ;
        RECT -1.540 0.870 -1.370 0.900 ;
        RECT -1.130 0.870 -0.930 0.910 ;
        RECT -1.540 0.610 -0.930 0.870 ;
        RECT -1.540 0.570 -1.370 0.610 ;
        RECT -1.130 0.580 -0.930 0.610 ;
        RECT -1.130 0.220 -0.930 0.250 ;
        RECT -1.360 -0.040 -0.930 0.220 ;
        RECT -1.130 -0.080 -0.930 -0.040 ;
        RECT -0.540 -0.080 0.010 0.910 ;
        RECT 0.480 0.900 1.180 1.210 ;
        RECT 0.480 0.290 1.190 0.460 ;
        RECT 0.830 0.010 1.190 0.290 ;
        RECT 0.830 -0.160 1.410 0.010 ;
      LAYER mcon ;
        RECT -1.300 5.090 -1.130 5.260 ;
        RECT 0.950 5.140 1.120 5.310 ;
        RECT -0.320 4.770 -0.150 4.940 ;
        RECT -1.350 4.440 -1.180 4.610 ;
        RECT -1.350 3.620 -1.180 3.790 ;
        RECT 0.340 3.830 0.510 4.000 ;
        RECT -0.320 3.290 -0.150 3.460 ;
        RECT -1.300 2.970 -1.130 3.140 ;
        RECT 1.000 2.920 1.170 3.090 ;
        RECT -1.300 2.130 -1.130 2.300 ;
        RECT 0.990 2.200 1.160 2.370 ;
        RECT -0.320 1.810 -0.150 1.980 ;
        RECT -1.350 1.480 -1.180 1.650 ;
        RECT 0.340 1.240 0.510 1.410 ;
        RECT -1.350 0.660 -1.180 0.830 ;
        RECT -0.320 0.330 -0.150 0.500 ;
        RECT -1.300 0.010 -1.130 0.180 ;
        RECT 0.910 -0.050 1.080 0.120 ;
      LAYER met1 ;
        RECT -1.370 5.020 -1.050 5.340 ;
        RECT -1.420 4.370 -1.100 4.690 ;
        RECT -1.420 3.540 -1.100 3.860 ;
        RECT -1.370 2.890 -1.050 3.210 ;
        RECT -1.370 2.060 -1.050 2.380 ;
        RECT -1.420 1.410 -1.100 1.730 ;
        RECT -1.420 0.580 -1.100 0.900 ;
        RECT -1.370 -0.070 -1.050 0.250 ;
        RECT -0.410 -0.220 -0.070 5.500 ;
        RECT 0.260 4.060 0.530 5.490 ;
        RECT 0.880 5.070 1.200 5.390 ;
        RECT 0.260 3.770 0.540 4.060 ;
        RECT 0.260 1.470 0.530 3.770 ;
        RECT 0.930 2.850 1.250 3.170 ;
        RECT 0.920 2.130 1.240 2.450 ;
        RECT 0.260 1.180 0.540 1.470 ;
        RECT 0.260 -0.210 0.530 1.180 ;
        RECT 0.840 -0.120 1.160 0.200 ;
      LAYER via ;
        RECT -1.340 5.050 -1.080 5.310 ;
        RECT -1.390 4.400 -1.130 4.660 ;
        RECT -1.390 3.570 -1.130 3.830 ;
        RECT -1.340 2.920 -1.080 3.180 ;
        RECT -1.340 2.090 -1.080 2.350 ;
        RECT -1.390 1.440 -1.130 1.700 ;
        RECT -1.390 0.610 -1.130 0.870 ;
        RECT -1.340 -0.040 -1.080 0.220 ;
        RECT 0.910 5.100 1.170 5.360 ;
        RECT 0.960 2.880 1.220 3.140 ;
        RECT 0.950 2.160 1.210 2.420 ;
        RECT 0.870 -0.090 1.130 0.170 ;
      LAYER met2 ;
        RECT -1.370 5.300 -1.060 5.350 ;
        RECT 0.880 5.300 1.190 5.400 ;
        RECT -1.370 5.070 1.190 5.300 ;
        RECT -1.370 5.020 -1.060 5.070 ;
        RECT -1.420 4.620 -1.110 4.700 ;
        RECT -1.720 4.410 -1.110 4.620 ;
        RECT -1.420 4.370 -1.110 4.410 ;
        RECT -1.420 3.820 -1.110 3.860 ;
        RECT -1.720 3.610 -1.110 3.820 ;
        RECT -1.420 3.530 -1.110 3.610 ;
        RECT -1.370 3.160 -1.060 3.210 ;
        RECT 0.930 3.160 1.240 3.180 ;
        RECT -1.370 2.930 1.550 3.160 ;
        RECT -1.370 2.880 -1.060 2.930 ;
        RECT 0.930 2.850 1.240 2.930 ;
        RECT -1.370 2.330 -1.060 2.390 ;
        RECT 0.920 2.330 1.230 2.460 ;
        RECT -1.370 2.110 1.550 2.330 ;
        RECT -1.370 2.060 -1.060 2.110 ;
        RECT -1.420 1.660 -1.110 1.740 ;
        RECT -1.720 1.450 -1.110 1.660 ;
        RECT -1.420 1.410 -1.110 1.450 ;
        RECT -1.420 0.860 -1.110 0.900 ;
        RECT -1.720 0.650 -1.110 0.860 ;
        RECT -1.420 0.570 -1.110 0.650 ;
        RECT -1.370 0.170 -1.060 0.250 ;
        RECT 0.840 0.170 1.150 0.210 ;
        RECT -1.370 -0.060 1.340 0.170 ;
        RECT -1.370 -0.080 -1.060 -0.060 ;
        RECT 0.840 -0.120 1.150 -0.060 ;
  END
END sky130_hilas_DualTACore01

MACRO sky130_hilas_TA2Cell_NoFG
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TA2Cell_NoFG ;
  ORIGIN 14.730 -1.400 ;
  SIZE 17.920 BY 6.050 ;
  PIN GATECOLSELECT
    ANTENNAGATEAREA 0.310000 ;
    PORT
      LAYER li1 ;
        RECT -4.160 5.980 -3.970 5.990 ;
        RECT -4.160 5.690 -3.960 5.980 ;
        RECT -4.170 5.360 -3.930 5.690 ;
        RECT -4.170 3.160 -3.930 3.490 ;
        RECT -4.160 2.870 -3.960 3.160 ;
        RECT -4.160 2.860 -3.970 2.870 ;
      LAYER mcon ;
        RECT -4.150 5.730 -3.970 5.920 ;
        RECT -4.150 2.930 -3.970 3.120 ;
      LAYER met1 ;
        RECT -4.160 5.990 -3.970 7.450 ;
        RECT -4.160 5.960 -3.940 5.990 ;
        RECT -4.180 5.690 -3.930 5.960 ;
        RECT -4.170 5.680 -3.930 5.690 ;
        RECT -4.170 5.440 -3.940 5.680 ;
        RECT -4.130 3.410 -3.970 5.440 ;
        RECT -4.170 3.170 -3.940 3.410 ;
        RECT -4.170 3.160 -3.930 3.170 ;
        RECT -4.180 2.890 -3.930 3.160 ;
        RECT -4.160 2.860 -3.940 2.890 ;
        RECT -4.160 1.400 -3.970 2.860 ;
    END
  END GATECOLSELECT
  PIN VINN_AMP1
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER li1 ;
        RECT -2.520 1.710 -2.350 1.730 ;
        RECT -2.520 1.450 -1.960 1.710 ;
        RECT -2.520 1.400 -2.350 1.450 ;
      LAYER mcon ;
        RECT -2.190 1.500 -2.020 1.670 ;
      LAYER met1 ;
        RECT -2.270 1.420 -1.950 1.740 ;
      LAYER via ;
        RECT -2.240 1.450 -1.980 1.710 ;
      LAYER met2 ;
        RECT -2.260 1.670 -1.950 1.740 ;
        RECT -2.860 1.420 -1.950 1.670 ;
        RECT -2.260 1.410 -1.950 1.420 ;
    END
  END VINN_AMP1
  PIN VINP_AMP2
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER li1 ;
        RECT -0.930 4.730 -0.610 4.760 ;
        RECT -0.930 4.540 -0.600 4.730 ;
        RECT -0.930 4.500 -0.610 4.540 ;
        RECT -0.930 4.420 -0.760 4.500 ;
        RECT -0.980 4.250 -0.760 4.420 ;
        RECT -0.980 4.090 -0.810 4.250 ;
      LAYER mcon ;
        RECT -0.870 4.550 -0.700 4.720 ;
      LAYER met1 ;
        RECT -0.940 4.470 -0.620 4.790 ;
      LAYER via ;
        RECT -0.910 4.500 -0.650 4.760 ;
      LAYER met2 ;
        RECT -0.940 4.750 -0.630 4.790 ;
        RECT -1.030 4.740 -0.600 4.750 ;
        RECT -1.260 4.510 -0.160 4.740 ;
        RECT -0.940 4.460 -0.630 4.510 ;
    END
  END VINP_AMP2
  PIN VINN_AMP2
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER li1 ;
        RECT -0.960 7.400 -0.790 7.450 ;
        RECT -0.960 7.140 -0.400 7.400 ;
        RECT -0.960 7.120 -0.790 7.140 ;
      LAYER mcon ;
        RECT -0.630 7.180 -0.460 7.350 ;
      LAYER met1 ;
        RECT -0.710 7.110 -0.390 7.430 ;
      LAYER via ;
        RECT -0.680 7.140 -0.420 7.400 ;
      LAYER met2 ;
        RECT -1.300 7.430 -1.050 7.440 ;
        RECT -0.700 7.430 -0.390 7.440 ;
        RECT -1.300 7.180 -0.390 7.430 ;
        RECT -0.700 7.110 -0.390 7.180 ;
    END
  END VINN_AMP2
  PIN VOUT_AMP1
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER li1 ;
        RECT 0.510 4.160 0.710 4.200 ;
        RECT 2.570 4.190 2.890 4.230 ;
        RECT 0.280 3.900 0.710 4.160 ;
        RECT 2.110 4.010 2.900 4.190 ;
        RECT 2.570 4.000 2.900 4.010 ;
        RECT 2.570 3.970 2.890 4.000 ;
        RECT 0.510 3.870 0.710 3.900 ;
      LAYER mcon ;
        RECT 0.340 3.940 0.510 4.110 ;
        RECT 2.630 4.010 2.800 4.180 ;
      LAYER met1 ;
        RECT 0.270 3.870 0.590 4.190 ;
        RECT 2.560 3.940 2.880 4.260 ;
      LAYER via ;
        RECT 0.300 3.900 0.560 4.160 ;
        RECT 2.590 3.970 2.850 4.230 ;
      LAYER met2 ;
        RECT 0.270 4.140 0.580 4.200 ;
        RECT 2.560 4.140 2.870 4.270 ;
        RECT 0.270 3.920 3.190 4.140 ;
        RECT 0.270 3.870 0.580 3.920 ;
    END
  END VOUT_AMP1
  PIN VOUT_AMP2
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER li1 ;
        RECT 0.510 4.990 0.710 5.020 ;
        RECT 0.280 4.730 0.710 4.990 ;
        RECT 2.580 4.910 2.900 4.950 ;
        RECT 2.580 4.850 2.910 4.910 ;
        RECT 0.510 4.690 0.710 4.730 ;
        RECT 2.110 4.720 2.910 4.850 ;
        RECT 2.110 4.690 2.900 4.720 ;
        RECT 2.110 4.670 2.810 4.690 ;
      LAYER mcon ;
        RECT 0.340 4.780 0.510 4.950 ;
        RECT 2.640 4.730 2.810 4.900 ;
      LAYER met1 ;
        RECT 0.270 4.700 0.590 5.020 ;
        RECT 2.570 4.660 2.890 4.980 ;
      LAYER via ;
        RECT 0.300 4.730 0.560 4.990 ;
        RECT 2.600 4.690 2.860 4.950 ;
      LAYER met2 ;
        RECT 0.270 4.970 0.580 5.020 ;
        RECT 2.570 4.970 2.880 4.990 ;
        RECT 0.270 4.740 3.190 4.970 ;
        RECT 0.270 4.690 0.580 4.740 ;
        RECT 2.570 4.660 2.880 4.740 ;
    END
  END VOUT_AMP2
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 1.100 6.170 1.650 7.160 ;
        RECT 1.100 4.690 1.650 5.680 ;
        RECT 1.100 3.210 1.650 4.200 ;
        RECT 1.100 1.730 1.650 2.720 ;
      LAYER mcon ;
        RECT 1.320 6.580 1.490 6.750 ;
        RECT 1.320 5.100 1.490 5.270 ;
        RECT 1.320 3.620 1.490 3.790 ;
        RECT 1.320 2.140 1.490 2.310 ;
      LAYER met1 ;
        RECT 1.230 1.400 1.570 7.450 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 1.920 7.270 3.190 7.450 ;
        RECT 1.910 1.400 3.190 7.270 ;
      LAYER li1 ;
        RECT 2.120 5.840 2.820 6.150 ;
        RECT 1.970 5.610 2.820 5.840 ;
        RECT 2.120 5.270 2.820 5.610 ;
        RECT 2.120 3.250 2.820 3.590 ;
        RECT 1.970 3.020 2.820 3.250 ;
        RECT 2.120 2.710 2.820 3.020 ;
      LAYER mcon ;
        RECT 1.980 5.640 2.150 5.810 ;
        RECT 1.980 3.050 2.150 3.220 ;
      LAYER met1 ;
        RECT 1.900 5.870 2.170 7.450 ;
        RECT 1.900 5.580 2.180 5.870 ;
        RECT 1.900 3.280 2.170 5.580 ;
        RECT 1.900 2.990 2.180 3.280 ;
        RECT 1.900 1.400 2.170 2.990 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT -14.720 6.700 -12.990 7.450 ;
        RECT -6.510 7.440 -1.650 7.450 ;
        RECT -14.720 3.130 -12.980 6.700 ;
        RECT -10.960 5.060 -8.240 6.710 ;
        RECT -10.960 5.020 -8.250 5.060 ;
        RECT -10.960 3.690 -8.250 3.730 ;
        RECT -14.720 1.410 -12.990 3.130 ;
        RECT -10.960 2.040 -8.240 3.690 ;
        RECT -6.510 1.410 -0.090 7.440 ;
        RECT -1.950 1.400 -0.090 1.410 ;
      LAYER li1 ;
        RECT 0.510 7.120 0.710 7.160 ;
        RECT -5.610 6.870 -5.080 7.040 ;
        RECT -3.800 6.770 -3.600 7.120 ;
        RECT -3.800 6.740 -3.590 6.770 ;
        RECT -7.480 6.290 -7.130 6.460 ;
        RECT -6.110 6.290 -5.780 6.460 ;
        RECT -14.290 5.310 -13.740 5.740 ;
        RECT -10.660 5.500 -10.430 6.190 ;
        RECT -5.360 5.960 -5.190 6.480 ;
        RECT -5.520 5.700 -5.190 5.960 ;
        RECT -7.480 5.500 -7.130 5.670 ;
        RECT -6.110 5.500 -5.780 5.670 ;
        RECT -11.690 4.480 -11.500 4.880 ;
        RECT -7.470 4.710 -7.130 4.880 ;
        RECT -6.110 4.710 -5.780 4.880 ;
        RECT -5.360 4.790 -5.190 5.700 ;
        RECT -4.530 4.880 -4.360 6.490 ;
        RECT -3.810 6.160 -3.590 6.740 ;
        RECT -3.800 6.150 -3.590 6.160 ;
        RECT -11.880 4.470 -11.500 4.480 ;
        RECT -11.880 4.290 -8.140 4.470 ;
        RECT -11.880 4.250 -11.500 4.290 ;
        RECT -14.290 3.580 -13.740 4.010 ;
        RECT -11.690 3.870 -11.500 4.250 ;
        RECT -6.030 4.140 -5.860 4.710 ;
        RECT -4.530 4.690 -4.350 4.880 ;
        RECT -7.470 3.970 -7.130 4.140 ;
        RECT -6.110 3.970 -5.780 4.140 ;
        RECT -10.660 2.560 -10.430 3.290 ;
        RECT -7.480 3.180 -7.130 3.350 ;
        RECT -6.110 3.180 -5.780 3.350 ;
        RECT -5.360 3.200 -5.190 4.060 ;
        RECT -5.520 2.940 -5.190 3.200 ;
        RECT -7.480 2.390 -7.130 2.560 ;
        RECT -6.110 2.390 -5.780 2.560 ;
        RECT -5.360 2.370 -5.190 2.940 ;
        RECT -4.530 3.970 -4.350 4.160 ;
        RECT -4.530 2.360 -4.360 3.970 ;
        RECT -3.100 3.070 -2.920 6.980 ;
        RECT -2.290 5.190 -2.120 6.970 ;
        RECT -1.540 6.040 -1.360 6.970 ;
        RECT -0.810 6.710 -0.480 6.880 ;
        RECT 0.280 6.860 0.710 7.120 ;
        RECT 0.510 6.830 0.710 6.860 ;
        RECT 2.470 7.040 3.050 7.210 ;
        RECT 2.470 6.940 2.860 7.040 ;
        RECT 2.470 6.910 2.850 6.940 ;
        RECT 2.470 6.760 2.830 6.910 ;
        RECT -0.730 6.570 -0.480 6.710 ;
        RECT 2.120 6.590 2.830 6.760 ;
        RECT -0.730 6.310 -0.250 6.570 ;
        RECT 0.100 6.470 0.270 6.510 ;
        RECT 0.510 6.470 0.710 6.500 ;
        RECT -1.660 6.010 -1.340 6.040 ;
        RECT -1.660 5.820 -1.330 6.010 ;
        RECT -1.660 5.780 -1.340 5.820 ;
        RECT -2.370 5.130 -1.830 5.190 ;
        RECT -2.370 5.020 -1.820 5.130 ;
        RECT -2.010 4.900 -1.820 5.020 ;
        RECT -2.540 4.600 -2.370 4.760 ;
        RECT -2.540 4.430 -2.320 4.600 ;
        RECT -2.490 4.350 -2.320 4.430 ;
        RECT -2.490 4.310 -2.170 4.350 ;
        RECT -2.490 4.120 -2.160 4.310 ;
        RECT -2.490 4.090 -2.170 4.120 ;
        RECT -3.220 3.030 -2.900 3.070 ;
        RECT -3.220 2.840 -2.890 3.030 ;
        RECT -3.220 2.810 -2.900 2.840 ;
        RECT -3.800 2.690 -3.590 2.700 ;
        RECT -3.810 2.110 -3.590 2.690 ;
        RECT -3.800 2.080 -3.590 2.110 ;
        RECT -5.610 1.810 -5.080 1.980 ;
        RECT -3.800 1.730 -3.600 2.080 ;
        RECT -3.100 1.880 -2.920 2.810 ;
        RECT -2.290 2.540 -2.120 3.920 ;
        RECT -2.290 2.280 -1.810 2.540 ;
        RECT -2.290 2.140 -2.040 2.280 ;
        RECT -2.370 1.970 -2.040 2.140 ;
        RECT -1.540 1.870 -1.360 5.780 ;
        RECT -0.730 4.930 -0.560 6.310 ;
        RECT 0.100 6.210 0.710 6.470 ;
        RECT 0.100 6.180 0.270 6.210 ;
        RECT 0.510 6.170 0.710 6.210 ;
        RECT 0.100 5.640 0.270 5.670 ;
        RECT 0.510 5.640 0.710 5.680 ;
        RECT 0.100 5.380 0.710 5.640 ;
        RECT 0.100 5.340 0.270 5.380 ;
        RECT 0.510 5.350 0.710 5.380 ;
        RECT -0.450 3.830 -0.260 3.950 ;
        RECT -0.810 3.720 -0.260 3.830 ;
        RECT -0.810 3.660 -0.270 3.720 ;
        RECT -0.730 1.880 -0.560 3.660 ;
        RECT 0.100 3.510 0.270 3.550 ;
        RECT 0.510 3.510 0.710 3.540 ;
        RECT 0.100 3.250 0.710 3.510 ;
        RECT 0.100 3.220 0.270 3.250 ;
        RECT 0.510 3.210 0.710 3.250 ;
        RECT 0.100 2.680 0.270 2.710 ;
        RECT 0.510 2.680 0.710 2.720 ;
        RECT 0.100 2.420 0.710 2.680 ;
        RECT 0.100 2.380 0.270 2.420 ;
        RECT 0.510 2.390 0.710 2.420 ;
        RECT 2.120 2.100 2.830 2.270 ;
        RECT 0.510 2.030 0.710 2.060 ;
        RECT 0.280 1.770 0.710 2.030 ;
        RECT 0.510 1.730 0.710 1.770 ;
        RECT 2.470 1.820 2.830 2.100 ;
        RECT 2.470 1.650 3.050 1.820 ;
      LAYER mcon ;
        RECT -3.790 6.570 -3.620 6.740 ;
        RECT -10.630 5.990 -10.460 6.160 ;
        RECT -14.290 5.390 -14.020 5.660 ;
        RECT -10.630 5.540 -10.460 5.710 ;
        RECT -5.460 5.740 -5.290 5.910 ;
        RECT -11.870 4.280 -11.700 4.450 ;
        RECT -14.290 3.660 -14.020 3.930 ;
        RECT -10.630 3.040 -10.460 3.210 ;
        RECT -5.460 2.980 -5.290 3.150 ;
        RECT -10.630 2.590 -10.460 2.760 ;
        RECT 0.340 6.900 0.510 7.070 ;
        RECT 2.590 6.950 2.760 7.120 ;
        RECT -0.480 6.350 -0.310 6.520 ;
        RECT -1.600 5.830 -1.430 6.000 ;
        RECT -2.000 4.930 -1.830 5.100 ;
        RECT -2.430 4.130 -2.260 4.300 ;
        RECT -3.160 2.850 -2.990 3.020 ;
        RECT -3.790 2.110 -3.620 2.280 ;
        RECT -2.040 2.330 -1.870 2.500 ;
        RECT 0.290 6.250 0.460 6.420 ;
        RECT 0.290 5.430 0.460 5.600 ;
        RECT -0.440 3.750 -0.270 3.920 ;
        RECT 0.290 3.290 0.460 3.460 ;
        RECT 0.290 2.470 0.460 2.640 ;
        RECT 0.340 1.820 0.510 1.990 ;
        RECT 2.550 1.760 2.720 1.930 ;
      LAYER met1 ;
        RECT -14.380 1.400 -13.960 7.450 ;
        RECT -11.900 1.400 -11.670 7.450 ;
        RECT -10.680 6.240 -10.450 7.450 ;
        RECT -5.680 6.770 -5.380 7.150 ;
        RECT -3.720 6.800 -3.440 7.450 ;
        RECT 0.270 6.830 0.590 7.150 ;
        RECT 2.520 6.880 2.840 7.200 ;
        RECT -10.680 5.450 -10.420 6.240 ;
        RECT -3.830 6.200 -3.440 6.800 ;
        RECT -0.560 6.280 -0.240 6.600 ;
        RECT -5.530 5.670 -5.210 5.990 ;
        RECT -10.680 3.300 -10.450 5.450 ;
        RECT -4.560 4.880 -4.320 5.010 ;
        RECT -4.560 4.560 -4.300 4.880 ;
        RECT -3.720 4.600 -3.440 6.200 ;
        RECT 0.220 6.180 0.540 6.500 ;
        RECT -1.670 5.750 -1.350 6.070 ;
        RECT -0.450 5.590 -0.240 5.700 ;
        RECT -0.470 5.270 -0.210 5.590 ;
        RECT 0.220 5.350 0.540 5.670 ;
        RECT -2.030 4.870 -1.800 5.160 ;
        RECT -3.720 4.280 -3.360 4.600 ;
        RECT -4.560 3.960 -4.300 4.280 ;
        RECT -4.560 3.840 -4.320 3.960 ;
        RECT -10.680 2.510 -10.420 3.300 ;
        RECT -5.530 2.910 -5.210 3.230 ;
        RECT -3.720 2.650 -3.440 4.280 ;
        RECT -2.500 4.060 -2.180 4.380 ;
        RECT -2.010 3.580 -1.800 4.870 ;
        RECT -0.450 3.980 -0.240 5.270 ;
        RECT -0.470 3.690 -0.240 3.980 ;
        RECT -2.030 3.260 -1.770 3.580 ;
        RECT -2.010 3.150 -1.800 3.260 ;
        RECT 0.220 3.220 0.540 3.540 ;
        RECT -3.230 2.780 -2.910 3.100 ;
        RECT -10.680 1.400 -10.450 2.510 ;
        RECT -5.680 1.700 -5.380 2.080 ;
        RECT -3.830 2.050 -3.440 2.650 ;
        RECT -2.120 2.250 -1.800 2.570 ;
        RECT 0.220 2.390 0.540 2.710 ;
        RECT -3.720 1.400 -3.440 2.050 ;
        RECT 0.270 1.740 0.590 2.060 ;
        RECT 2.480 1.690 2.800 2.010 ;
      LAYER via ;
        RECT -5.660 6.830 -5.400 7.100 ;
        RECT 0.300 6.860 0.560 7.120 ;
        RECT 2.550 6.910 2.810 7.170 ;
        RECT -0.530 6.310 -0.270 6.570 ;
        RECT -5.500 5.700 -5.240 5.960 ;
        RECT -4.560 4.590 -4.300 4.850 ;
        RECT 0.250 6.210 0.510 6.470 ;
        RECT -1.640 5.780 -1.380 6.040 ;
        RECT -0.470 5.300 -0.210 5.560 ;
        RECT 0.250 5.380 0.510 5.640 ;
        RECT -3.620 4.310 -3.360 4.570 ;
        RECT -4.560 3.990 -4.300 4.250 ;
        RECT -5.500 2.940 -5.240 3.200 ;
        RECT -2.470 4.090 -2.210 4.350 ;
        RECT -2.030 3.290 -1.770 3.550 ;
        RECT 0.250 3.250 0.510 3.510 ;
        RECT -3.200 2.810 -2.940 3.070 ;
        RECT -2.090 2.280 -1.830 2.540 ;
        RECT 0.250 2.420 0.510 2.680 ;
        RECT -5.660 1.750 -5.400 2.020 ;
        RECT 0.300 1.770 0.560 2.030 ;
        RECT 2.510 1.720 2.770 1.980 ;
      LAYER met2 ;
        RECT -5.680 6.970 -5.380 7.150 ;
        RECT -5.930 6.950 -5.380 6.970 ;
        RECT 0.270 7.110 0.580 7.160 ;
        RECT 2.520 7.110 2.830 7.210 ;
        RECT -14.730 6.770 -3.200 6.950 ;
        RECT 0.270 6.880 2.830 7.110 ;
        RECT 0.270 6.830 0.580 6.880 ;
        RECT -0.550 6.570 -0.240 6.610 ;
        RECT -0.730 6.430 0.010 6.570 ;
        RECT 0.220 6.430 0.530 6.510 ;
        RECT -0.730 6.320 0.530 6.430 ;
        RECT -0.550 6.280 0.530 6.320 ;
        RECT -0.240 6.220 0.530 6.280 ;
        RECT -0.240 6.200 0.010 6.220 ;
        RECT 0.220 6.180 0.530 6.220 ;
        RECT -5.530 5.930 -5.220 6.000 ;
        RECT -1.670 5.930 -1.360 6.070 ;
        RECT -5.530 5.740 -1.360 5.930 ;
        RECT -5.530 5.710 -1.620 5.740 ;
        RECT -5.530 5.670 -5.220 5.710 ;
        RECT -0.210 5.630 0.000 5.640 ;
        RECT 0.220 5.630 0.530 5.670 ;
        RECT -0.210 5.560 0.530 5.630 ;
        RECT -0.500 5.540 0.530 5.560 ;
        RECT -0.550 5.420 0.530 5.540 ;
        RECT -0.550 5.350 0.000 5.420 ;
        RECT -0.550 5.290 -0.080 5.350 ;
        RECT 0.220 5.340 0.530 5.420 ;
        RECT -4.590 4.590 -4.270 4.850 ;
        RECT -4.550 4.570 -3.370 4.590 ;
        RECT -4.550 4.310 -3.330 4.570 ;
        RECT -2.500 4.340 -2.190 4.390 ;
        RECT -4.550 4.250 -3.370 4.310 ;
        RECT -4.590 4.240 -3.370 4.250 ;
        RECT -4.590 3.990 -4.270 4.240 ;
        RECT -2.820 4.110 -1.720 4.340 ;
        RECT -2.820 4.100 -2.160 4.110 ;
        RECT -2.500 4.060 -2.190 4.100 ;
        RECT -2.110 3.470 -1.640 3.560 ;
        RECT 0.220 3.470 0.530 3.550 ;
        RECT -2.110 3.310 0.530 3.470 ;
        RECT -2.060 3.290 0.530 3.310 ;
        RECT -1.770 3.270 0.530 3.290 ;
        RECT -0.080 3.260 0.530 3.270 ;
        RECT -5.530 3.170 -5.220 3.240 ;
        RECT 0.220 3.220 0.530 3.260 ;
        RECT -3.340 3.170 -3.180 3.180 ;
        RECT -5.530 3.110 -3.180 3.170 ;
        RECT -5.530 2.960 -2.920 3.110 ;
        RECT -5.530 2.910 -5.220 2.960 ;
        RECT -3.340 2.780 -2.920 2.960 ;
        RECT 0.220 2.670 0.530 2.710 ;
        RECT -2.060 2.570 0.530 2.670 ;
        RECT -2.110 2.530 0.530 2.570 ;
        RECT -2.290 2.460 0.530 2.530 ;
        RECT -2.290 2.280 -1.740 2.460 ;
        RECT 0.220 2.380 0.530 2.460 ;
        RECT -2.110 2.240 -1.800 2.280 ;
        RECT -5.670 2.080 -5.510 2.090 ;
        RECT -5.760 2.070 -3.200 2.080 ;
        RECT -14.730 1.920 -3.200 2.070 ;
        RECT -5.760 1.900 -3.200 1.920 ;
        RECT 0.270 1.980 0.580 2.060 ;
        RECT 2.480 1.980 2.790 2.020 ;
        RECT -5.680 1.700 -5.380 1.900 ;
        RECT 0.270 1.750 2.980 1.980 ;
        RECT 0.270 1.730 0.580 1.750 ;
        RECT 2.480 1.690 2.790 1.750 ;
  END
END sky130_hilas_TA2Cell_NoFG

MACRO sky130_hilas_pFETdevice01b
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pFETdevice01b ;
  ORIGIN 0.790 1.140 ;
  SIZE 1.870 BY 1.570 ;
  OBS
      LAYER nwell ;
        RECT -0.790 -0.780 0.820 0.430 ;
      LAYER li1 ;
        RECT 0.780 -1.060 0.990 -0.630 ;
        RECT 0.800 -1.080 0.970 -1.060 ;
      LAYER met1 ;
        RECT 0.780 -0.850 1.000 -0.630 ;
        RECT 0.770 -1.140 1.000 -0.850 ;
  END
END sky130_hilas_pFETdevice01b

MACRO sky130_hilas_capacitorArray01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_capacitorArray01 ;
  ORIGIN 13.040 0.570 ;
  SIZE 36.700 BY 6.050 ;
  PIN CAPTERMINAL2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 22.970 2.220 23.660 2.630 ;
      LAYER via2 ;
        RECT 23.040 2.280 23.330 2.560 ;
      LAYER met3 ;
        RECT -0.530 3.270 22.190 5.320 ;
        RECT -0.530 1.630 23.340 3.270 ;
        RECT -0.530 -0.400 22.190 1.630 ;
        RECT 22.640 1.620 23.340 1.630 ;
    END
  END CAPTERMINAL2
  PIN CAPTERM01
    USE ANALOG ;
    ANTENNADIFFAREA 0.459000 ;
    PORT
      LAYER li1 ;
        RECT -5.420 4.490 -5.100 4.530 ;
        RECT -5.420 4.450 -5.090 4.490 ;
        RECT -5.420 4.280 -4.840 4.450 ;
        RECT -5.420 4.270 -5.100 4.280 ;
        RECT -4.290 4.210 -4.090 4.780 ;
        RECT -4.290 3.140 -4.090 3.710 ;
        RECT -4.290 1.200 -4.090 1.770 ;
        RECT -4.290 0.140 -4.090 0.710 ;
      LAYER mcon ;
        RECT -4.280 4.570 -4.110 4.740 ;
        RECT -5.360 4.310 -5.190 4.480 ;
        RECT -4.280 3.180 -4.110 3.350 ;
        RECT -4.280 1.560 -4.110 1.730 ;
        RECT -4.280 0.180 -4.110 0.350 ;
      LAYER met1 ;
        RECT -4.290 5.460 -4.130 5.480 ;
        RECT -4.340 5.140 -4.080 5.460 ;
        RECT -4.290 4.800 -4.130 5.140 ;
        RECT -4.290 4.780 -4.090 4.800 ;
        RECT -5.430 4.240 -5.110 4.560 ;
        RECT -4.310 4.540 -4.080 4.780 ;
        RECT -4.290 4.320 -4.090 4.540 ;
        RECT -4.290 3.600 -4.130 4.320 ;
        RECT -4.290 3.380 -4.090 3.600 ;
        RECT -4.310 3.140 -4.080 3.380 ;
        RECT -4.290 3.120 -4.090 3.140 ;
        RECT -4.290 1.790 -4.130 3.120 ;
        RECT -4.290 1.770 -4.090 1.790 ;
        RECT -4.310 1.530 -4.080 1.770 ;
        RECT -4.290 1.310 -4.090 1.530 ;
        RECT -4.290 0.600 -4.130 1.310 ;
        RECT -4.290 0.380 -4.090 0.600 ;
        RECT -4.310 0.140 -4.080 0.380 ;
        RECT -4.290 0.120 -4.090 0.140 ;
        RECT -4.290 -0.560 -4.130 0.120 ;
      LAYER via ;
        RECT -4.340 5.170 -4.080 5.430 ;
        RECT -5.400 4.270 -5.140 4.530 ;
      LAYER met2 ;
        RECT -2.300 5.450 -1.790 5.480 ;
        RECT -4.370 5.360 -4.050 5.430 ;
        RECT -2.300 5.360 -1.370 5.450 ;
        RECT -4.370 5.170 -1.370 5.360 ;
        RECT -1.870 5.150 -1.370 5.170 ;
        RECT -5.430 4.550 -5.120 4.570 ;
        RECT -13.040 4.370 23.660 4.550 ;
        RECT -5.430 4.240 -5.120 4.370 ;
        RECT -1.740 3.970 -1.370 4.370 ;
      LAYER via2 ;
        RECT -1.740 5.150 -1.460 5.430 ;
        RECT -1.690 4.030 -1.410 4.310 ;
      LAYER met3 ;
        RECT -1.790 5.170 -1.410 5.460 ;
        RECT -1.870 4.520 -1.330 5.170 ;
        RECT -1.960 3.770 -1.170 4.520 ;
      LAYER via3 ;
        RECT -1.770 3.920 -1.340 4.400 ;
      LAYER met4 ;
        RECT -1.870 4.310 -1.210 4.490 ;
        RECT -1.940 4.200 0.760 4.310 ;
        RECT -1.940 3.990 0.970 4.200 ;
        RECT -1.940 3.980 1.040 3.990 ;
        RECT -1.940 3.900 1.090 3.980 ;
        RECT -1.870 3.830 -1.210 3.900 ;
        RECT 0.460 3.560 1.090 3.900 ;
        RECT 0.570 3.490 1.090 3.560 ;
    END
  END CAPTERM01
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -5.520 -0.560 22.380 5.480 ;
        RECT -1.040 -0.570 22.380 -0.560 ;
      LAYER li1 ;
        RECT -3.560 4.800 -3.360 5.150 ;
        RECT -3.560 4.770 -3.350 4.800 ;
        RECT -3.570 4.180 -3.350 4.770 ;
        RECT -3.570 3.150 -3.350 3.740 ;
        RECT -3.560 3.120 -3.350 3.150 ;
        RECT -3.560 2.770 -3.360 3.120 ;
        RECT -3.560 1.790 -3.360 2.140 ;
        RECT -3.560 1.760 -3.350 1.790 ;
        RECT -3.570 1.170 -3.350 1.760 ;
        RECT -3.570 0.150 -3.350 0.740 ;
        RECT -3.560 0.120 -3.350 0.150 ;
        RECT -3.560 -0.230 -3.360 0.120 ;
      LAYER mcon ;
        RECT -3.550 4.600 -3.380 4.770 ;
        RECT -3.550 3.150 -3.380 3.320 ;
        RECT -3.550 1.590 -3.380 1.760 ;
        RECT -3.550 0.150 -3.380 0.320 ;
      LAYER met1 ;
        RECT -3.480 4.830 -3.320 5.480 ;
        RECT -3.590 4.280 -3.320 4.830 ;
        RECT -3.590 4.230 -3.310 4.280 ;
        RECT -3.480 4.140 -3.310 4.230 ;
        RECT -3.480 3.780 -3.320 4.140 ;
        RECT -3.480 3.690 -3.310 3.780 ;
        RECT -3.590 3.640 -3.310 3.690 ;
        RECT -3.590 3.090 -3.320 3.640 ;
        RECT -3.480 1.820 -3.320 3.090 ;
        RECT -3.590 1.270 -3.320 1.820 ;
        RECT -3.590 1.220 -3.310 1.270 ;
        RECT -3.480 1.130 -3.310 1.220 ;
        RECT -3.480 0.780 -3.320 1.130 ;
        RECT -3.480 0.690 -3.310 0.780 ;
        RECT -3.590 0.640 -3.310 0.690 ;
        RECT -3.590 0.090 -3.320 0.640 ;
        RECT -3.480 -0.560 -3.320 0.090 ;
    END
  END VINJ
  PIN GATESELECT
    ANTENNAGATEAREA 0.620000 ;
    PORT
      LAYER li1 ;
        RECT -4.170 2.370 -3.730 2.540 ;
      LAYER mcon ;
        RECT -3.910 2.370 -3.730 2.540 ;
      LAYER met1 ;
        RECT -3.920 4.490 -3.730 5.480 ;
        RECT -3.900 4.370 -3.730 4.490 ;
        RECT -3.890 3.550 -3.730 4.370 ;
        RECT -3.900 3.430 -3.730 3.550 ;
        RECT -3.920 2.570 -3.730 3.430 ;
        RECT -3.940 2.340 -3.700 2.570 ;
        RECT -3.920 1.480 -3.730 2.340 ;
        RECT -3.900 1.360 -3.730 1.480 ;
        RECT -3.890 0.550 -3.730 1.360 ;
        RECT -3.900 0.430 -3.730 0.550 ;
        RECT -3.920 -0.560 -3.730 0.430 ;
    END
  END GATESELECT
  PIN VTUN
    ANTENNADIFFAREA 1.978000 ;
    PORT
      LAYER nwell ;
        RECT -13.030 3.620 -11.300 5.480 ;
        RECT -13.040 1.780 -11.300 3.620 ;
        RECT -13.030 -0.570 -11.300 1.780 ;
      LAYER li1 ;
        RECT -12.610 2.230 -12.060 2.660 ;
      LAYER mcon ;
        RECT -12.610 2.310 -12.340 2.580 ;
      LAYER met1 ;
        RECT -12.680 -0.570 -12.280 5.480 ;
    END
  END VTUN
  PIN GATE
    USE ANALOG ;
    ANTENNADIFFAREA 2.743300 ;
    PORT
      LAYER nwell ;
        RECT -9.280 -0.560 -7.050 5.470 ;
      LAYER li1 ;
        RECT -8.580 2.160 -8.030 2.590 ;
      LAYER mcon ;
        RECT -8.580 2.240 -8.310 2.510 ;
      LAYER met1 ;
        RECT -8.630 3.560 -8.250 5.480 ;
        RECT -8.640 1.700 -8.250 3.560 ;
        RECT -8.630 -0.440 -8.250 1.700 ;
        RECT -8.640 -0.560 -8.250 -0.440 ;
    END
  END GATE
  OBS
      LAYER li1 ;
        RECT -5.420 5.070 -5.100 5.080 ;
        RECT -5.420 4.900 -4.840 5.070 ;
        RECT -5.420 4.850 -5.090 4.900 ;
        RECT -5.420 4.820 -5.100 4.850 ;
        RECT -5.420 3.640 -5.100 3.650 ;
        RECT -5.420 3.470 -4.840 3.640 ;
        RECT -5.420 3.430 -5.090 3.470 ;
        RECT -5.420 3.390 -5.100 3.430 ;
        RECT -5.420 3.070 -5.100 3.100 ;
        RECT -5.420 3.020 -5.090 3.070 ;
        RECT -5.420 2.850 -4.840 3.020 ;
        RECT -5.420 2.840 -5.100 2.850 ;
        RECT -5.420 2.060 -5.100 2.070 ;
        RECT -5.420 1.890 -4.840 2.060 ;
        RECT -5.420 1.840 -5.090 1.890 ;
        RECT -5.420 1.810 -5.100 1.840 ;
        RECT -5.420 1.480 -5.100 1.520 ;
        RECT -5.420 1.440 -5.090 1.480 ;
        RECT -5.420 1.270 -4.840 1.440 ;
        RECT -5.420 1.260 -5.100 1.270 ;
        RECT -5.420 0.640 -5.100 0.650 ;
        RECT -5.420 0.470 -4.840 0.640 ;
        RECT -5.420 0.430 -5.090 0.470 ;
        RECT -5.420 0.390 -5.100 0.430 ;
        RECT -5.420 0.070 -5.100 0.100 ;
        RECT -5.420 0.020 -5.090 0.070 ;
        RECT -5.420 -0.150 -4.840 0.020 ;
        RECT -5.420 -0.160 -5.100 -0.150 ;
      LAYER mcon ;
        RECT -5.360 4.860 -5.190 5.030 ;
        RECT -5.360 3.440 -5.190 3.610 ;
        RECT -5.360 2.890 -5.190 3.060 ;
        RECT -5.360 1.850 -5.190 2.020 ;
        RECT -5.360 1.300 -5.190 1.470 ;
        RECT -5.360 0.440 -5.190 0.610 ;
        RECT -5.360 -0.110 -5.190 0.060 ;
      LAYER met1 ;
        RECT -5.430 4.790 -5.110 5.110 ;
        RECT -5.430 3.360 -5.110 3.680 ;
        RECT -5.430 2.810 -5.110 3.130 ;
        RECT -5.430 1.780 -5.110 2.100 ;
        RECT -5.430 1.230 -5.110 1.550 ;
        RECT -5.430 0.360 -5.110 0.680 ;
        RECT -5.430 -0.190 -5.110 0.130 ;
      LAYER via ;
        RECT -5.400 4.820 -5.140 5.080 ;
        RECT -5.400 3.390 -5.140 3.650 ;
        RECT -5.400 2.840 -5.140 3.100 ;
        RECT -5.400 1.810 -5.140 2.070 ;
        RECT -5.400 1.260 -5.140 1.520 ;
        RECT -5.400 0.390 -5.140 0.650 ;
        RECT -5.400 -0.160 -5.140 0.100 ;
      LAYER met2 ;
        RECT -5.430 4.980 -5.120 5.120 ;
        RECT -13.040 4.800 23.660 4.980 ;
        RECT -5.430 4.790 -5.120 4.800 ;
        RECT -5.430 3.550 -5.120 3.680 ;
        RECT -3.160 3.550 -2.790 3.720 ;
        RECT -13.040 3.370 23.660 3.550 ;
        RECT -5.430 3.350 -5.120 3.370 ;
        RECT -3.160 3.320 -2.790 3.370 ;
        RECT -5.430 3.120 -5.120 3.130 ;
        RECT 22.650 3.120 23.660 3.130 ;
        RECT -13.040 2.940 23.660 3.120 ;
        RECT -5.430 2.800 -5.120 2.940 ;
        RECT -5.430 1.970 -5.120 2.110 ;
        RECT -5.430 1.960 -2.960 1.970 ;
        RECT -13.020 1.790 23.660 1.960 ;
        RECT -5.430 1.780 -5.120 1.790 ;
        RECT -5.430 1.540 -5.120 1.560 ;
        RECT -3.200 1.540 -2.830 1.630 ;
        RECT -13.020 1.370 23.660 1.540 ;
        RECT -5.520 1.360 -2.830 1.370 ;
        RECT -5.430 1.230 -5.120 1.360 ;
        RECT -3.200 1.230 -2.830 1.360 ;
        RECT -5.430 0.560 -5.120 0.680 ;
        RECT -2.110 0.560 -1.740 0.760 ;
        RECT -13.020 0.550 -5.120 0.560 ;
        RECT -4.190 0.550 23.660 0.560 ;
        RECT -13.020 0.390 23.660 0.550 ;
        RECT -12.240 0.300 -10.700 0.390 ;
        RECT -5.520 0.370 -2.960 0.390 ;
        RECT -5.430 0.350 -5.120 0.370 ;
        RECT -2.110 0.360 -1.740 0.390 ;
        RECT -5.430 0.120 -5.120 0.130 ;
        RECT -13.020 -0.050 23.660 0.120 ;
        RECT -5.430 -0.060 -2.960 -0.050 ;
        RECT -5.430 -0.200 -5.120 -0.060 ;
      LAYER via2 ;
        RECT -3.110 3.380 -2.830 3.660 ;
        RECT -3.150 1.290 -2.870 1.570 ;
        RECT -2.060 0.420 -1.780 0.700 ;
      LAYER met3 ;
        RECT -3.380 3.120 -2.590 3.870 ;
        RECT -3.420 1.730 -2.630 1.780 ;
        RECT -3.420 1.430 -2.490 1.730 ;
        RECT -3.420 1.030 -2.630 1.430 ;
        RECT -2.330 0.520 -1.540 0.910 ;
        RECT -2.330 0.220 -1.400 0.520 ;
        RECT -2.330 0.160 -1.540 0.220 ;
      LAYER via3 ;
        RECT -3.190 3.270 -2.760 3.750 ;
        RECT -3.230 1.180 -2.800 1.660 ;
        RECT -2.140 0.310 -1.710 0.790 ;
      LAYER met4 ;
        RECT -0.250 4.810 3.850 5.110 ;
        RECT 3.470 3.990 3.850 4.810 ;
        RECT 3.430 3.980 3.880 3.990 ;
        RECT 6.270 3.980 6.720 3.990 ;
        RECT 9.110 3.980 9.560 3.990 ;
        RECT 11.950 3.980 12.400 3.990 ;
        RECT 14.790 3.980 15.240 3.990 ;
        RECT 17.630 3.980 18.080 3.990 ;
        RECT 20.470 3.980 20.920 3.990 ;
        RECT -3.290 3.480 -2.630 3.840 ;
        RECT 3.410 3.490 3.930 3.980 ;
        RECT 6.250 3.940 6.770 3.980 ;
        RECT 9.090 3.940 9.610 3.980 ;
        RECT 6.250 3.640 9.610 3.940 ;
        RECT 6.250 3.490 6.770 3.640 ;
        RECT 9.090 3.490 9.610 3.640 ;
        RECT 11.930 3.920 12.450 3.980 ;
        RECT 14.770 3.920 15.290 3.980 ;
        RECT 17.610 3.920 18.130 3.980 ;
        RECT 20.450 3.920 20.970 3.980 ;
        RECT 11.930 3.620 20.970 3.920 ;
        RECT 11.930 3.490 12.450 3.620 ;
        RECT 14.770 3.590 18.130 3.620 ;
        RECT 14.770 3.490 15.290 3.590 ;
        RECT 17.610 3.490 18.130 3.590 ;
        RECT 20.450 3.490 20.970 3.620 ;
        RECT -3.290 3.180 -1.270 3.480 ;
        RECT -1.570 2.620 -1.270 3.180 ;
        RECT 6.310 2.620 6.610 3.490 ;
        RECT 9.290 2.620 9.590 3.490 ;
        RECT -1.570 2.320 9.590 2.620 ;
        RECT -3.330 1.730 -2.670 1.750 ;
        RECT 0.670 1.730 3.860 1.760 ;
        RECT 6.310 1.730 6.610 1.760 ;
        RECT -3.330 1.430 9.530 1.730 ;
        RECT -3.330 1.090 -2.670 1.430 ;
        RECT 0.670 1.130 0.970 1.430 ;
        RECT 3.560 1.130 3.860 1.430 ;
        RECT 6.310 1.130 6.610 1.430 ;
        RECT 9.230 1.130 9.530 1.430 ;
        RECT 11.990 1.130 12.290 3.490 ;
        RECT 14.820 1.130 15.120 3.490 ;
        RECT 17.630 1.130 17.930 3.490 ;
        RECT 20.580 1.130 20.880 3.490 ;
        RECT 0.590 1.120 1.040 1.130 ;
        RECT 3.430 1.120 3.880 1.130 ;
        RECT 6.270 1.120 6.720 1.130 ;
        RECT 9.110 1.120 9.560 1.130 ;
        RECT 11.950 1.120 12.400 1.130 ;
        RECT 14.790 1.120 15.240 1.130 ;
        RECT 17.630 1.120 18.080 1.130 ;
        RECT 20.470 1.120 20.920 1.130 ;
        RECT 0.570 1.060 1.090 1.120 ;
        RECT 3.410 1.090 3.930 1.120 ;
        RECT 6.250 1.090 6.770 1.120 ;
        RECT 3.410 1.060 6.770 1.090 ;
        RECT 9.090 1.060 9.610 1.120 ;
        RECT -2.240 0.520 -1.580 0.880 ;
        RECT 0.570 0.760 9.610 1.060 ;
        RECT 0.570 0.630 1.090 0.760 ;
        RECT 3.410 0.630 3.930 0.760 ;
        RECT 6.250 0.630 6.770 0.760 ;
        RECT 9.090 0.630 9.610 0.760 ;
        RECT 11.930 1.100 12.450 1.120 ;
        RECT 14.770 1.100 15.290 1.120 ;
        RECT 17.610 1.100 18.130 1.120 ;
        RECT 20.450 1.100 20.970 1.120 ;
        RECT 11.930 0.800 20.970 1.100 ;
        RECT 11.930 0.630 12.450 0.800 ;
        RECT 14.770 0.630 15.290 0.800 ;
        RECT 17.610 0.790 20.970 0.800 ;
        RECT 17.610 0.630 18.130 0.790 ;
        RECT 20.450 0.630 20.970 0.790 ;
        RECT -2.240 0.220 -1.190 0.520 ;
        RECT -1.490 -0.020 -1.190 0.220 ;
        RECT 20.640 -0.020 20.940 0.630 ;
        RECT -1.490 -0.320 20.940 -0.020 ;
  END
END sky130_hilas_capacitorArray01

MACRO sky130_hilas_li2m1
  CLASS BLOCK ;
  FOREIGN sky130_hilas_li2m1 ;
  ORIGIN 0.100 0.080 ;
  SIZE 0.230 BY 0.290 ;
  OBS
      LAYER li1 ;
        RECT -0.080 -0.050 0.110 0.180 ;
      LAYER mcon ;
        RECT -0.070 -0.020 0.100 0.150 ;
      LAYER met1 ;
        RECT -0.100 -0.080 0.130 0.210 ;
  END
END sky130_hilas_li2m1

MACRO sky130_hilas_capacitorSize03
  CLASS BLOCK ;
  FOREIGN sky130_hilas_capacitorSize03 ;
  ORIGIN -14.140 0.470 ;
  SIZE 5.790 BY 5.870 ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 19.230 2.640 19.600 2.700 ;
        RECT 19.230 2.360 19.930 2.640 ;
        RECT 19.230 2.300 19.600 2.360 ;
      LAYER via2 ;
        RECT 19.280 2.360 19.560 2.640 ;
      LAYER met3 ;
        RECT 15.590 2.850 18.430 5.400 ;
        RECT 15.590 2.100 19.800 2.850 ;
        RECT 15.590 -0.470 18.430 2.100 ;
      LAYER via3 ;
        RECT 19.200 2.250 19.630 2.730 ;
      LAYER met4 ;
        RECT 19.100 2.160 19.760 2.820 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 14.380 2.600 14.750 2.660 ;
        RECT 14.160 2.320 14.750 2.600 ;
        RECT 14.380 2.260 14.750 2.320 ;
      LAYER via2 ;
        RECT 14.430 2.320 14.710 2.600 ;
      LAYER met3 ;
        RECT 14.160 2.060 14.950 2.810 ;
      LAYER via3 ;
        RECT 14.350 2.210 14.780 2.690 ;
      LAYER met4 ;
        RECT 16.710 4.060 17.160 4.070 ;
        RECT 16.690 3.570 17.210 4.060 ;
        RECT 14.250 2.720 14.910 2.780 ;
        RECT 16.720 2.730 17.160 3.570 ;
        RECT 15.300 2.720 16.310 2.730 ;
        RECT 16.710 2.720 17.170 2.730 ;
        RECT 14.250 2.220 17.170 2.720 ;
        RECT 14.250 2.210 15.660 2.220 ;
        RECT 14.250 2.120 14.910 2.210 ;
        RECT 16.710 1.560 17.170 2.220 ;
        RECT 16.710 1.050 17.190 1.560 ;
        RECT 16.690 0.560 17.210 1.050 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 14.140 4.800 19.920 4.980 ;
        RECT 14.140 4.370 19.920 4.550 ;
        RECT 14.170 3.370 19.920 3.550 ;
        RECT 14.170 2.940 19.920 3.120 ;
        RECT 14.170 1.790 19.920 1.960 ;
        RECT 14.170 1.370 19.920 1.540 ;
        RECT 14.170 0.390 19.920 0.560 ;
        RECT 14.170 -0.050 19.920 0.120 ;
  END
END sky130_hilas_capacitorSize03

MACRO sky130_hilas_TunCap01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TunCap01 ;
  ORIGIN 14.510 4.000 ;
  SIZE 1.730 BY 1.900 ;
  OBS
      LAYER nwell ;
        RECT -14.510 -4.000 -12.780 -2.100 ;
  END
END sky130_hilas_TunCap01

MACRO sky130_hilas_pFETLargePart1
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pFETLargePart1 ;
  ORIGIN 0.060 0.090 ;
  SIZE 3.390 BY 2.870 ;
  OBS
      LAYER nwell ;
        RECT -0.060 -0.090 3.330 2.780 ;
      LAYER li1 ;
        RECT 0.180 0.060 0.350 2.550 ;
        RECT 0.730 0.050 0.900 2.550 ;
        RECT 1.280 0.050 1.450 2.550 ;
        RECT 1.830 0.050 2.000 2.550 ;
        RECT 2.380 0.050 2.550 2.550 ;
        RECT 2.930 0.050 3.100 2.550 ;
  END
END sky130_hilas_pFETLargePart1

MACRO sky130_hilas_pFETdevice01e
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pFETdevice01e ;
  ORIGIN 1.210 0.550 ;
  SIZE 2.030 BY 0.990 ;
  OBS
      LAYER nwell ;
        RECT -1.210 -0.550 0.820 0.440 ;
      LAYER li1 ;
        RECT -0.860 0.190 -0.540 0.230 ;
        RECT -0.860 0.170 -0.530 0.190 ;
        RECT -0.860 -0.030 -0.240 0.170 ;
        RECT -0.410 -0.160 -0.240 -0.030 ;
        RECT 0.270 0.130 0.440 0.170 ;
        RECT 0.270 0.090 0.760 0.130 ;
        RECT 0.270 -0.100 0.770 0.090 ;
        RECT 0.270 -0.130 0.760 -0.100 ;
        RECT 0.270 -0.160 0.440 -0.130 ;
        RECT -1.020 -0.270 -0.590 -0.250 ;
        RECT -1.040 -0.440 -0.590 -0.270 ;
        RECT -1.020 -0.460 -0.590 -0.440 ;
      LAYER mcon ;
        RECT -0.800 0.010 -0.630 0.180 ;
        RECT 0.500 -0.090 0.670 0.080 ;
      LAYER met1 ;
        RECT -0.870 -0.060 -0.550 0.260 ;
        RECT 0.430 -0.160 0.750 0.160 ;
        RECT -0.870 -0.240 -0.550 -0.200 ;
        RECT -1.100 -0.470 -0.550 -0.240 ;
        RECT -0.870 -0.520 -0.550 -0.470 ;
      LAYER via ;
        RECT -0.840 -0.030 -0.580 0.230 ;
        RECT 0.460 -0.130 0.720 0.130 ;
        RECT -0.840 -0.490 -0.580 -0.230 ;
      LAYER met2 ;
        RECT -0.870 0.160 -0.560 0.270 ;
        RECT -1.210 -0.030 -0.560 0.160 ;
        RECT -0.870 -0.060 -0.560 -0.030 ;
        RECT 0.430 -0.160 0.740 0.170 ;
        RECT -0.870 -0.260 -0.550 -0.200 ;
        RECT -1.210 -0.450 -0.550 -0.260 ;
        RECT -0.870 -0.520 -0.550 -0.450 ;
  END
END sky130_hilas_pFETdevice01e

MACRO sky130_hilas_nFET03
  CLASS BLOCK ;
  FOREIGN sky130_hilas_nFET03 ;
  ORIGIN 0.310 0.190 ;
  SIZE 0.890 BY 0.610 ;
  OBS
      LAYER li1 ;
        RECT -0.260 -0.050 -0.060 0.280 ;
        RECT 0.330 -0.050 0.530 0.280 ;
  END
END sky130_hilas_nFET03

MACRO sky130_hilas_nFETmirrorPairs2
  CLASS BLOCK ;
  FOREIGN sky130_hilas_nFETmirrorPairs2 ;
  ORIGIN 3.090 1.920 ;
  SIZE 4.670 BY 4.770 ;
  OBS
      LAYER nwell ;
        RECT -0.610 1.120 1.580 2.850 ;
      LAYER li1 ;
        RECT -0.400 2.010 1.360 2.530 ;
        RECT -0.400 1.400 0.310 1.570 ;
        RECT 0.620 1.400 1.320 1.570 ;
        RECT -0.050 1.230 0.310 1.400 ;
        RECT -0.050 0.870 0.600 1.230 ;
        RECT -3.040 0.410 -2.840 0.740 ;
        RECT -2.450 0.410 -2.250 0.740 ;
        RECT -0.050 0.640 0.220 0.870 ;
        RECT 0.850 0.650 1.100 1.400 ;
        RECT -0.080 0.470 0.250 0.640 ;
        RECT 0.770 0.470 1.100 0.650 ;
        RECT -3.040 -0.240 -2.840 0.090 ;
        RECT -2.450 -0.240 -2.250 0.090 ;
        RECT -0.120 -0.200 0.290 0.040 ;
        RECT 0.730 -0.200 1.140 0.040 ;
        RECT -0.120 -0.580 1.140 -0.200 ;
        RECT -3.040 -1.060 -2.840 -0.730 ;
        RECT -2.450 -1.060 -2.250 -0.730 ;
        RECT -0.120 -0.840 0.290 -0.580 ;
        RECT 0.730 -0.830 1.140 -0.580 ;
        RECT -3.040 -1.700 -2.840 -1.370 ;
        RECT -2.450 -1.700 -2.250 -1.370 ;
        RECT -0.090 -1.430 0.250 -1.260 ;
        RECT 0.760 -1.430 1.120 -1.250 ;
        RECT -0.010 -1.920 0.170 -1.430 ;
        RECT 0.840 -1.920 1.030 -1.430 ;
  END
END sky130_hilas_nFETmirrorPairs2

MACRO sky130_hilas_nFET03a
  CLASS BLOCK ;
  FOREIGN sky130_hilas_nFET03a ;
  ORIGIN 1.110 0.470 ;
  SIZE 2.080 BY 0.890 ;
  OBS
      LAYER li1 ;
        RECT -0.260 0.240 -0.060 0.280 ;
        RECT -0.570 -0.020 -0.060 0.240 ;
        RECT -0.260 -0.050 -0.060 -0.020 ;
        RECT 0.330 0.250 0.530 0.280 ;
        RECT 0.330 0.210 0.840 0.250 ;
        RECT 0.330 0.020 0.850 0.210 ;
        RECT 0.330 -0.010 0.840 0.020 ;
        RECT 0.330 -0.050 0.530 -0.010 ;
        RECT -1.010 -0.220 -0.580 -0.200 ;
        RECT -1.010 -0.390 -0.560 -0.220 ;
        RECT -1.010 -0.410 -0.580 -0.390 ;
      LAYER mcon ;
        RECT -0.510 0.020 -0.340 0.190 ;
        RECT 0.580 0.030 0.750 0.200 ;
        RECT -0.730 -0.390 -0.560 -0.220 ;
      LAYER met1 ;
        RECT -0.580 -0.050 -0.260 0.270 ;
        RECT 0.510 -0.040 0.830 0.280 ;
        RECT -1.050 -0.190 -0.730 -0.140 ;
        RECT -1.050 -0.420 -0.500 -0.190 ;
        RECT -1.050 -0.460 -0.730 -0.420 ;
      LAYER via ;
        RECT -0.550 -0.020 -0.290 0.240 ;
        RECT 0.540 -0.010 0.800 0.250 ;
        RECT -1.020 -0.430 -0.760 -0.170 ;
      LAYER met2 ;
        RECT -0.580 0.190 -0.270 0.280 ;
        RECT -1.110 0.020 -0.270 0.190 ;
        RECT -0.580 -0.050 -0.270 0.020 ;
        RECT 0.510 0.200 0.820 0.290 ;
        RECT 0.510 0.030 0.970 0.200 ;
        RECT 0.510 -0.040 0.820 0.030 ;
        RECT -1.050 -0.220 -0.730 -0.140 ;
        RECT -1.110 -0.390 -0.730 -0.220 ;
        RECT -1.050 -0.460 -0.730 -0.390 ;
  END
END sky130_hilas_nFET03a

END LIBRARY