VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_FGBiasWeakGate2x1cell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_FGBiasWeakGate2x1cell ;
  ORIGIN 3.960 3.820 ;
  SIZE 11.530 BY 6.050 ;
  PIN drain1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -3.960 1.550 5.110 1.730 ;
    END
  END drain1
  PIN Input1
    PORT
      LAYER met2 ;
        RECT -3.960 0.950 -1.990 1.130 ;
    END
  END Input1
  PIN output1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.530 0.490 7.570 0.710 ;
    END
  END output1
  PIN output2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.530 -2.260 7.570 -2.050 ;
    END
  END output2
  PIN Vinj
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 7.050 1.520 7.330 2.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 7.050 -3.820 7.330 -3.110 ;
    END
  END Vinj
  PIN GateSelect
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 6.610 0.700 6.800 2.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.610 -3.820 6.800 -2.290 ;
    END
  END GateSelect
  PIN GND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT -1.130 -0.770 -0.900 2.230 ;
    END
    PORT
      LAYER met1 ;
        RECT -1.130 -3.820 -0.900 -0.940 ;
    END
  END GND
  PIN gate_control
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 0.090 0.940 0.320 2.230 ;
    END
  END gate_control
  PIN Vtun
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT -3.610 0.440 -3.190 2.230 ;
    END
  END Vtun
  PIN gateControl
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 0.090 -3.820 0.320 -2.630 ;
    END
  END gateControl
  PIN drain4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -3.960 -3.300 5.110 -3.150 ;
    END
  END drain4
  PIN Input2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -3.960 -2.790 -2.020 -2.580 ;
    END
  END Input2
  PIN CommonSource
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -3.960 -0.490 6.210 -0.270 ;
    END
  END CommonSource
  OBS
      LAYER li1 ;
        RECT -3.520 -3.720 7.180 2.050 ;
      LAYER met1 ;
        RECT -2.910 0.160 -1.410 1.930 ;
        RECT -3.610 -3.810 -1.410 0.160 ;
        RECT -0.620 0.660 -0.190 1.930 ;
        RECT 0.600 0.660 6.330 1.930 ;
        RECT -0.620 0.420 6.330 0.660 ;
        RECT 7.080 0.420 7.330 1.240 ;
        RECT -0.620 -2.010 7.330 0.420 ;
        RECT -0.620 -2.350 6.330 -2.010 ;
        RECT -0.620 -3.810 -0.190 -2.350 ;
        RECT 0.600 -3.810 6.330 -2.350 ;
        RECT 7.080 -2.830 7.330 -2.010 ;
      LAYER met2 ;
        RECT 5.390 1.270 7.570 1.930 ;
        RECT -1.710 0.990 7.570 1.270 ;
        RECT -1.710 0.670 5.250 0.990 ;
        RECT -3.960 0.210 5.250 0.670 ;
        RECT -3.960 0.010 7.570 0.210 ;
        RECT 6.490 -0.770 7.570 0.010 ;
        RECT -3.960 -1.770 7.570 -0.770 ;
        RECT -3.960 -2.300 5.250 -1.770 ;
        RECT -1.740 -2.540 5.250 -2.300 ;
        RECT -1.740 -2.870 7.570 -2.540 ;
        RECT 5.390 -3.520 7.570 -2.870 ;
  END
END sky130_hilas_FGBiasWeakGate2x1cell
END LIBRARY

