magic
tech sky130A
timestamp 1637801776
<< error_p >>
rect -29 232 6 236
rect -252 210 -199 219
rect -279 204 -252 210
rect -199 204 -171 210
rect -73 209 -21 219
rect -101 204 -73 209
rect -279 185 -276 204
rect -252 168 -199 177
rect -73 167 -21 177
<< nwell >>
rect -336 144 -138 308
<< mvnmos >>
rect -73 177 -21 209
<< mvpmos >>
rect -252 177 -199 210
<< mvndiff >>
rect -101 202 -73 209
rect -101 185 -96 202
rect -79 185 -73 202
rect -101 177 -73 185
rect -21 201 7 209
rect -21 184 -15 201
rect 2 184 7 201
rect -21 177 7 184
<< mvpdiff >>
rect -279 202 -252 210
rect -279 185 -275 202
rect -258 185 -252 202
rect -279 177 -252 185
rect -199 202 -171 210
rect -199 185 -193 202
rect -176 185 -171 202
rect -199 177 -171 185
<< mvndiffc >>
rect -96 185 -79 202
rect -15 184 2 201
<< mvpdiffc >>
rect -275 185 -258 202
rect -193 185 -176 202
<< psubdiff >>
rect -29 256 15 264
rect -29 239 -15 256
rect 2 239 15 256
rect -29 232 15 239
<< mvnsubdiff >>
rect -286 267 -245 275
rect -286 250 -274 267
rect -257 250 -245 267
rect -286 241 -245 250
<< psubdiffcont >>
rect -15 239 2 256
<< mvnsubdiffcont >>
rect -274 250 -257 267
<< poly >>
rect -322 224 -36 227
rect -322 212 -21 224
rect -322 202 -295 212
rect -252 210 -199 212
rect -322 185 -317 202
rect -300 185 -295 202
rect -322 177 -295 185
rect -73 209 -21 212
rect -252 164 -199 177
rect -73 164 -21 177
<< polycont >>
rect -317 185 -300 202
<< locali >>
rect -274 267 -257 279
rect -274 248 -272 250
rect -15 256 2 264
rect -274 238 -257 248
rect -15 229 2 239
rect -317 202 -300 210
rect -302 183 -300 185
rect -317 177 -300 183
rect -275 204 -258 210
rect -275 202 -250 204
rect -258 197 -250 202
rect -275 180 -271 185
rect -254 180 -250 197
rect -201 202 -176 210
rect -201 185 -193 202
rect -176 185 -137 202
rect -120 185 -96 202
rect -79 185 -71 202
rect -15 201 2 212
rect -275 177 -250 180
rect -274 175 -250 177
rect -193 176 -176 185
rect -23 184 -15 201
rect 2 184 10 201
<< viali >>
rect -272 250 -257 265
rect -257 250 -255 265
rect -272 248 -255 250
rect -15 212 2 229
rect -319 185 -317 200
rect -317 185 -302 200
rect -319 183 -302 185
rect -271 185 -258 197
rect -258 185 -254 197
rect -271 180 -254 185
rect -137 185 -120 202
<< metal1 >>
rect -275 270 -253 304
rect -275 265 -252 270
rect -275 248 -272 265
rect -255 248 -252 265
rect -275 244 -252 248
rect -328 205 -297 211
rect -328 179 -325 205
rect -299 179 -297 205
rect -328 176 -297 179
rect -275 204 -253 244
rect -18 229 5 304
rect -18 212 -15 229
rect 2 212 5 229
rect -275 197 -250 204
rect -275 180 -271 197
rect -254 180 -250 197
rect -145 180 -142 206
rect -116 180 -113 206
rect -275 173 -250 180
rect -275 153 -253 173
rect -18 153 5 212
<< via1 >>
rect -325 200 -299 205
rect -325 183 -319 200
rect -319 183 -302 200
rect -302 183 -299 200
rect -325 179 -299 183
rect -142 202 -116 206
rect -142 185 -137 202
rect -137 185 -120 202
rect -120 185 -116 202
rect -142 180 -116 185
<< metal2 >>
rect -336 247 25 265
rect -328 195 -325 205
rect -329 179 -325 195
rect -299 179 -296 205
rect -145 180 -142 206
rect -116 198 -113 206
rect -116 180 25 198
<< labels >>
rlabel metal1 -275 153 -253 159 0 Vinj
rlabel metal1 -275 297 -253 304 0 Vinj
rlabel metal1 -18 295 5 304 0 GND
rlabel metal1 -18 153 5 159 0 GND
rlabel metal2 -336 247 -326 265 0 Input
rlabel metal2 16 247 25 265 0 Input
rlabel metal2 16 180 25 198 0 Output
<< end >>
