magic
tech sky130A
timestamp 1628707334
<< error_p >>
rect 62 613 69 614
rect 1 375 86 381
rect 0 347 86 375
rect 29 344 30 347
rect 42 344 48 347
rect 29 341 51 344
rect 52 341 86 347
rect 104 346 107 349
rect 27 338 86 341
rect 27 335 36 338
rect 29 319 30 335
rect 33 327 36 335
rect 42 335 86 338
rect 42 327 51 335
rect 33 324 51 327
rect 42 321 51 324
rect 42 319 48 321
rect 52 319 86 335
rect 107 345 110 346
rect 107 320 108 345
rect 29 318 86 319
<< nwell >>
rect 30 398 177 667
rect 1 374 177 398
rect 0 291 177 374
rect 30 0 177 291
<< mvpmos >>
rect 81 557 111 607
rect 81 420 111 471
rect 81 347 111 399
rect 81 266 111 318
rect 81 195 111 245
rect 81 60 111 110
<< mvndiff >>
rect 29 318 52 347
<< mvpdiff >>
rect 81 630 111 634
rect 81 613 87 630
rect 104 613 111 630
rect 81 607 111 613
rect 81 551 111 557
rect 81 534 87 551
rect 105 534 111 551
rect 81 529 111 534
rect 81 494 111 499
rect 81 477 87 494
rect 105 477 111 494
rect 81 471 111 477
rect 81 399 111 420
rect 81 341 111 347
rect 81 324 87 341
rect 105 324 111 341
rect 81 318 111 324
rect 81 245 111 266
rect 81 189 111 195
rect 81 172 87 189
rect 105 172 111 189
rect 81 168 111 172
rect 81 133 111 137
rect 81 116 87 133
rect 105 116 111 133
rect 81 110 111 116
rect 81 54 111 60
rect 81 37 87 54
rect 105 37 111 54
rect 81 33 111 37
<< mvpdiffc >>
rect 87 613 104 630
rect 87 534 105 551
rect 87 477 105 494
rect 87 324 105 341
rect 87 172 105 189
rect 87 116 105 133
rect 87 37 105 54
<< poly >>
rect 47 557 81 607
rect 111 557 124 607
rect 47 471 68 557
rect 47 420 81 471
rect 111 420 126 471
rect 68 347 81 399
rect 111 347 137 399
rect 114 318 137 347
rect 68 266 81 318
rect 111 266 137 318
rect 52 195 81 245
rect 111 195 124 245
rect 52 110 68 195
rect 52 60 81 110
rect 111 60 124 110
rect 52 59 68 60
<< locali >>
rect 80 613 87 630
rect 104 613 112 630
rect 79 534 87 551
rect 105 534 113 551
rect 79 477 87 494
rect 105 477 113 494
rect 48 324 62 341
rect 80 324 87 341
rect 105 324 113 341
rect 79 172 87 189
rect 105 172 113 189
rect 79 116 87 133
rect 105 116 113 133
rect 79 37 87 54
rect 105 37 113 54
<< viali >>
rect 62 613 80 630
rect 33 324 48 341
rect 62 324 80 341
<< metal1 >>
rect 66 637 100 641
rect 66 636 70 637
rect 56 630 70 636
rect 96 636 100 637
rect 56 613 62 630
rect 56 611 70 613
rect 96 611 112 636
rect 66 608 100 611
rect 56 341 82 345
rect 56 324 62 341
rect 80 324 82 341
rect 56 320 82 324
rect 107 320 110 345
<< via1 >>
rect 70 630 96 637
rect 70 613 80 630
rect 80 613 96 630
rect 70 611 96 613
rect 82 320 107 346
<< metal2 >>
rect 66 637 100 641
rect 30 611 70 637
rect 96 611 149 637
rect 66 608 100 611
rect 80 347 110 348
rect 80 346 111 347
rect 60 320 82 346
rect 107 320 113 346
rect 60 319 113 320
rect 80 317 110 319
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
