* NGSPICE file created from /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_pFETmed.ext - technology: sky130A


* Top level circuit /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_pFETmed

X0 a_440_n8# a_388_n34# a_330_n8# w_294_n44# sky130_fd_pr__pfet_01v8 w=2.51e+06u l=260000u
.end

