* Copyright 2020 The Hilas PDK Authors
* 
* This file is part of HILAS.
* 
* HILAS is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published by
* the Free Software Foundation, version 3 of the License.
* 
* HILAS is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
* 
* You should have received a copy of the GNU Lesser General Public License
* along with HILAS.  If not, see <https://www.gnu.org/licenses/>.
* 
* Licensed under the Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
* https://www.gnu.org/licenses/lgpl-3.0.en.html
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
* SPDX-License-Identifier: LGPL-3.0
* 
* 

* NGSPICE file created from sky130_hilas_drainSelect01.ext - technology: sky130A

.subckt sky130_hilas_TgateVinj01 a_n354_n14# $SUB a_86_n14# w_n420_n80# a_n194_n14#
+ a_446_110# DrainSelect
X0 a_n194_110# DrainSelect a_n354_n14# w_n420_n80# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
X1 a_446_110# DrainSelect a_n194_110# $SUB sky130_fd_pr__nfet_g5v0d10v5 w=310000u l=500000u
X2 a_86_n14# a_n194_110# a_n194_n14# w_n420_n80# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
X3 a_n194_n14# DrainSelect a_n354_n14# w_n420_n80# sky130_fd_pr__pfet_g5v0d10v5 w=320000u l=500000u
X4 a_n194_n14# DrainSelect a_86_n14# $SUB sky130_fd_pr__nfet_g5v0d10v5 w=310000u l=500000u
.ends

.subckt sky130_hilas_drainSelect01 DRAIN4 DRAIN3 DRAIN2 DRAIN1 DRAINSELECT1 DRAINSELECT2
+ DRAINSELECT3 DRAINSELECT4 VINJ DRAIN_MUX VGND
Xsky130_hilas_TgateVinj01_0 VINJ $SUB DRAIN_MUX sky130_hilas_TgateVinj01_3/w_n420_n80#
+ DRAIN2 VGND DRAINSELECT2 sky130_hilas_TgateVinj01
Xsky130_hilas_TgateVinj01_1 VINJ $SUB DRAIN_MUX sky130_hilas_TgateVinj01_3/w_n420_n80#
+ DRAIN1 VGND DRAINSELECT1 sky130_hilas_TgateVinj01
Xsky130_hilas_TgateVinj01_2 VINJ $SUB DRAIN_MUX sky130_hilas_TgateVinj01_3/w_n420_n80#
+ DRAIN4 VGND DRAINSELECT4 sky130_hilas_TgateVinj01
Xsky130_hilas_TgateVinj01_3 VINJ $SUB DRAIN_MUX sky130_hilas_TgateVinj01_3/w_n420_n80#
+ DRAIN3 VGND DRAINSELECT3 sky130_hilas_TgateVinj01
.ends

