**.subckt nFETLarge Gate1n Drain1n Source1n
*.ipin Gate1n
*.iopin Drain1n
*.iopin Source1n
XM3 Drain1n Gate1n Source1n GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
**.ends
.GLOBAL GND
** flattened .save nodes
.end
