magic
tech sky130A
timestamp 1627401235
<< error_s >>
rect 14865 37094 14894 37110
rect 14944 37094 14973 37110
rect 15023 37094 15052 37110
rect 15102 37094 15131 37110
rect 13727 37070 13734 37076
rect 14578 37070 14584 37076
rect 15410 37070 15416 37076
rect 15515 37070 15521 37076
rect 15930 37065 15936 37071
rect 15985 37065 15991 37071
rect 14865 37060 14866 37061
rect 14893 37060 14894 37061
rect 14944 37060 14945 37061
rect 14972 37060 14973 37061
rect 15023 37060 15024 37061
rect 15051 37060 15052 37061
rect 15102 37060 15103 37061
rect 15130 37060 15131 37061
rect 14815 37031 14832 37060
rect 14864 37059 14895 37060
rect 14943 37059 14974 37060
rect 15022 37059 15053 37060
rect 15101 37059 15132 37060
rect 14865 37052 14894 37059
rect 14944 37052 14973 37059
rect 15023 37052 15052 37059
rect 15102 37052 15131 37059
rect 14865 37038 14874 37052
rect 15121 37038 15131 37052
rect 14865 37032 14894 37038
rect 14944 37032 14973 37038
rect 15023 37032 15052 37038
rect 15102 37032 15131 37038
rect 14864 37031 14895 37032
rect 14943 37031 14974 37032
rect 15022 37031 15053 37032
rect 15101 37031 15132 37032
rect 15163 37031 15181 37060
rect 14865 37030 14866 37031
rect 14893 37030 14894 37031
rect 14944 37030 14945 37031
rect 14972 37030 14973 37031
rect 15023 37030 15024 37031
rect 15051 37030 15052 37031
rect 15102 37030 15103 37031
rect 15130 37030 15131 37031
rect 15404 37020 15410 37026
rect 15521 37020 15527 37026
rect 15924 37015 15930 37021
rect 15991 37015 15997 37021
rect 14865 36981 14894 36996
rect 14944 36981 14973 36996
rect 15023 36981 15052 36996
rect 15102 36981 15131 36996
rect 14865 36814 14894 36830
rect 14944 36814 14973 36830
rect 15023 36814 15052 36830
rect 15102 36814 15131 36830
rect 13419 36811 13424 36812
rect 14865 36780 14866 36781
rect 14893 36780 14894 36781
rect 14944 36780 14945 36781
rect 14972 36780 14973 36781
rect 15023 36780 15024 36781
rect 15051 36780 15052 36781
rect 15102 36780 15103 36781
rect 15130 36780 15131 36781
rect 14815 36751 14832 36780
rect 14864 36779 14895 36780
rect 14943 36779 14974 36780
rect 15022 36779 15053 36780
rect 15101 36779 15132 36780
rect 14865 36772 14894 36779
rect 14944 36772 14973 36779
rect 15023 36772 15052 36779
rect 15102 36772 15131 36779
rect 14865 36758 14874 36772
rect 15121 36758 15131 36772
rect 14865 36752 14894 36758
rect 14944 36752 14973 36758
rect 15023 36752 15052 36758
rect 15102 36752 15131 36758
rect 14864 36751 14895 36752
rect 14943 36751 14974 36752
rect 15022 36751 15053 36752
rect 15101 36751 15132 36752
rect 15163 36751 15181 36780
rect 15410 36771 15416 36777
rect 15515 36771 15521 36777
rect 14865 36750 14866 36751
rect 14893 36750 14894 36751
rect 14944 36750 14945 36751
rect 14972 36750 14973 36751
rect 15023 36750 15024 36751
rect 15051 36750 15052 36751
rect 15102 36750 15103 36751
rect 15130 36750 15131 36751
rect 15961 36732 15990 36750
rect 15404 36721 15410 36727
rect 15521 36721 15527 36727
rect 14865 36701 14894 36716
rect 14944 36701 14973 36716
rect 15023 36701 15052 36716
rect 15102 36701 15131 36716
rect 15961 36700 15962 36701
rect 15989 36700 15990 36701
rect 13131 36644 13132 36699
rect 14865 36659 14894 36675
rect 14944 36659 14973 36675
rect 15023 36659 15052 36675
rect 15102 36659 15131 36675
rect 15410 36670 15416 36676
rect 15515 36670 15521 36676
rect 15911 36671 15929 36700
rect 15960 36699 15991 36700
rect 15961 36690 15990 36699
rect 15961 36681 15971 36690
rect 15980 36681 15990 36690
rect 15961 36672 15990 36681
rect 15960 36671 15991 36672
rect 16022 36671 16040 36700
rect 15961 36670 15962 36671
rect 15989 36670 15990 36671
rect 14865 36625 14866 36626
rect 14893 36625 14894 36626
rect 14944 36625 14945 36626
rect 14972 36625 14973 36626
rect 15023 36625 15024 36626
rect 15051 36625 15052 36626
rect 15102 36625 15103 36626
rect 15130 36625 15131 36626
rect 13722 36604 13728 36610
rect 14584 36604 14590 36610
rect 14815 36596 14832 36625
rect 14864 36624 14895 36625
rect 14943 36624 14974 36625
rect 15022 36624 15053 36625
rect 15101 36624 15132 36625
rect 14865 36617 14894 36624
rect 14944 36617 14973 36624
rect 15023 36617 15052 36624
rect 15102 36617 15131 36624
rect 14865 36603 14874 36617
rect 15121 36603 15131 36617
rect 14865 36597 14894 36603
rect 14944 36597 14973 36603
rect 15023 36597 15052 36603
rect 15102 36597 15131 36603
rect 14864 36596 14895 36597
rect 14943 36596 14974 36597
rect 15022 36596 15053 36597
rect 15101 36596 15132 36597
rect 15163 36596 15181 36625
rect 15404 36620 15410 36626
rect 15521 36620 15527 36626
rect 15961 36621 15990 36639
rect 14865 36595 14866 36596
rect 14893 36595 14894 36596
rect 14944 36595 14945 36596
rect 14972 36595 14973 36596
rect 15023 36595 15024 36596
rect 15051 36595 15052 36596
rect 15102 36595 15103 36596
rect 15130 36595 15131 36596
rect 14865 36546 14894 36561
rect 14944 36546 14973 36561
rect 15023 36546 15052 36561
rect 15102 36546 15131 36561
rect 19537 35790 19550 35791
rect 19156 35569 19162 35575
rect 19209 35569 19215 35575
rect 19322 35569 19328 35575
rect 19375 35569 19381 35575
rect 19150 35519 19156 35525
rect 19215 35519 19221 35525
rect 19316 35519 19322 35525
rect 19381 35519 19387 35525
rect 18728 35510 18734 35516
rect 18833 35510 18839 35516
rect 19745 35510 19751 35516
rect 19850 35510 19856 35516
rect 18722 35460 18728 35466
rect 18839 35460 18845 35466
rect 19739 35460 19745 35466
rect 19856 35460 19862 35466
rect 16589 35330 16952 35331
rect 17009 35330 17132 35331
rect 17207 35324 17237 35443
rect 18728 35209 18734 35215
rect 18833 35209 18839 35215
rect 19745 35209 19751 35215
rect 19850 35209 19856 35215
rect 18722 35159 18728 35165
rect 18839 35159 18845 35165
rect 19156 35155 19162 35161
rect 19209 35155 19215 35161
rect 19322 35155 19328 35161
rect 19375 35155 19381 35161
rect 19739 35159 19745 35165
rect 19856 35159 19862 35165
rect 19150 35105 19156 35111
rect 19215 35105 19221 35111
rect 19316 35105 19322 35111
rect 19381 35105 19387 35111
rect 18990 35042 18994 35053
rect 18990 35028 18991 35039
rect 19099 35038 19100 35091
rect 19157 34966 19163 34972
rect 19210 34966 19216 34972
rect 19322 34966 19328 34972
rect 19375 34966 19381 34972
rect 19151 34916 19157 34922
rect 19216 34916 19222 34922
rect 19316 34916 19322 34922
rect 19381 34916 19387 34922
rect 18682 34907 18688 34913
rect 18787 34907 18793 34913
rect 19745 34907 19751 34913
rect 19850 34907 19856 34913
rect 18676 34857 18682 34863
rect 18793 34857 18799 34863
rect 19739 34857 19745 34863
rect 19856 34857 19862 34863
rect 19550 34722 19567 34723
rect 19550 34705 19567 34706
rect 18988 34688 18989 34701
rect 18682 34606 18688 34612
rect 18787 34606 18793 34612
rect 19745 34606 19751 34612
rect 19850 34606 19856 34612
rect 18676 34556 18682 34562
rect 18793 34556 18799 34562
rect 19157 34552 19163 34558
rect 19210 34552 19216 34558
rect 19322 34552 19328 34558
rect 19375 34552 19381 34558
rect 19739 34556 19745 34562
rect 19856 34556 19862 34562
rect 19151 34502 19157 34508
rect 19216 34502 19222 34508
rect 19316 34502 19322 34508
rect 19381 34502 19387 34508
rect 18730 34241 18736 34247
rect 18835 34241 18841 34247
rect 19701 34241 19707 34247
rect 19806 34241 19812 34247
rect 19156 34231 19162 34237
rect 19209 34231 19215 34237
rect 19327 34231 19333 34237
rect 19380 34231 19386 34237
rect 18724 34177 18730 34183
rect 18841 34177 18847 34183
rect 19150 34181 19156 34187
rect 19215 34181 19221 34187
rect 19321 34181 19327 34187
rect 19386 34181 19392 34187
rect 19695 34177 19701 34183
rect 19812 34177 19818 34183
rect 18730 34124 18736 34130
rect 18835 34124 18841 34130
rect 19156 34122 19162 34128
rect 19209 34122 19215 34128
rect 19327 34122 19333 34128
rect 19380 34122 19386 34128
rect 19701 34124 19707 34130
rect 19806 34124 19812 34130
rect 19150 34072 19156 34078
rect 19215 34072 19221 34078
rect 19321 34072 19327 34078
rect 19386 34072 19392 34078
rect 18724 34060 18730 34066
rect 18841 34060 18847 34066
rect 19695 34060 19701 34066
rect 19812 34060 19818 34066
rect 18730 33939 18736 33945
rect 18835 33939 18841 33945
rect 19701 33939 19707 33945
rect 19806 33939 19812 33945
rect 19156 33933 19162 33939
rect 19209 33933 19215 33939
rect 19327 33933 19333 33939
rect 19380 33933 19386 33939
rect 19150 33883 19156 33889
rect 19215 33883 19221 33889
rect 19321 33883 19327 33889
rect 19386 33883 19392 33889
rect 18724 33875 18730 33881
rect 18841 33875 18847 33881
rect 19695 33875 19701 33881
rect 19812 33875 19818 33881
rect 18730 33823 18736 33829
rect 18835 33823 18841 33829
rect 19701 33823 19707 33829
rect 19806 33823 19812 33829
rect 19156 33816 19162 33822
rect 19209 33816 19215 33822
rect 19327 33816 19333 33822
rect 19380 33816 19386 33822
rect 19150 33766 19156 33772
rect 19215 33766 19221 33772
rect 19321 33766 19327 33772
rect 19386 33766 19392 33772
rect 18724 33759 18730 33765
rect 18841 33759 18847 33765
rect 19695 33759 19701 33765
rect 19812 33759 19818 33765
rect 18730 33263 18736 33269
rect 18835 33263 18841 33269
rect 19156 33253 19162 33259
rect 19209 33253 19215 33259
rect 18724 33199 18730 33205
rect 18841 33199 18847 33205
rect 19150 33203 19156 33209
rect 19215 33203 19221 33209
rect 18730 33146 18736 33152
rect 18835 33146 18841 33152
rect 19156 33144 19162 33150
rect 19209 33144 19215 33150
rect 19150 33094 19156 33100
rect 19215 33094 19221 33100
rect 18724 33082 18730 33088
rect 18841 33082 18847 33088
rect 18730 32961 18736 32967
rect 18835 32961 18841 32967
rect 18993 32956 19010 32960
rect 19156 32955 19162 32961
rect 19209 32955 19215 32961
rect 19150 32905 19156 32911
rect 19215 32905 19221 32911
rect 18724 32897 18730 32903
rect 18841 32897 18847 32903
rect 18730 32845 18736 32851
rect 18835 32845 18841 32851
rect 19156 32838 19162 32844
rect 19209 32838 19215 32844
rect 19150 32788 19156 32794
rect 19215 32788 19221 32794
rect 18724 32781 18730 32787
rect 18841 32781 18847 32787
rect 24292 32042 24293 32055
rect 24292 32041 24306 32042
rect 13994 31883 14001 31921
rect 14008 31889 14015 31935
rect 14560 31499 14572 31502
rect 14548 31478 14553 31490
rect 18883 31450 18884 31468
rect 18897 31450 18898 31454
rect 14541 31138 14553 31146
rect 14772 31138 14774 31146
rect 23302 30993 23303 30995
rect 16235 30243 16402 30256
rect 16828 30246 16830 30259
rect 16232 30229 16402 30242
rect 16828 30232 16831 30245
rect 17238 30244 17239 30257
rect 17238 30230 17240 30243
<< metal1 >>
rect 2385 38791 2774 38908
rect 5244 38790 5633 38907
rect 8103 38790 8492 38907
rect 12293 38793 12682 38910
rect 16505 38791 16894 38908
rect 19364 38791 19753 38908
rect 22224 38791 22613 38908
rect 25083 38791 25472 38908
rect 27942 38791 28331 38908
rect 30801 38790 31190 38907
rect 33660 38790 34049 38907
rect 2937 36559 3260 37870
rect 5796 36900 6119 37870
rect 8655 37329 8978 37870
rect 9909 37649 9926 37661
rect 8612 37298 8995 37329
rect 8612 37073 8655 37298
rect 8978 37073 8995 37298
rect 8612 37055 8995 37073
rect 9874 36993 9926 37649
rect 9868 36982 9933 36993
rect 9868 36945 9874 36982
rect 9926 36945 9933 36982
rect 9868 36942 9933 36945
rect 5780 36849 6130 36900
rect 5780 36624 5796 36849
rect 6119 36624 6130 36849
rect 5780 36611 6130 36624
rect 2720 36520 3260 36559
rect 2720 36197 2754 36520
rect 2979 36197 3260 36520
rect 1476 36189 1815 36196
rect 1379 36180 1815 36189
rect 1056 35857 1601 36180
rect 1787 35857 1815 36180
rect 2720 36179 3014 36197
rect 9874 36174 9926 36942
rect 10214 36551 10255 37672
rect 12925 37472 13041 37663
rect 12925 37359 15661 37472
rect 12925 37339 15680 37359
rect 15528 37199 15661 37339
rect 17057 37248 17380 37871
rect 18221 37663 18282 37677
rect 18219 37467 18337 37663
rect 18139 37376 18337 37467
rect 18139 37358 18320 37376
rect 18663 37360 18735 37746
rect 18139 37289 18212 37358
rect 19916 37248 20239 37870
rect 22775 37248 23098 37870
rect 23668 37609 23687 37610
rect 24381 37609 24453 37746
rect 23668 37574 24453 37609
rect 23668 37361 23687 37574
rect 25634 37555 25957 37870
rect 25558 37527 25957 37555
rect 25556 37507 25957 37527
rect 25538 37410 25973 37507
rect 25538 37204 25634 37410
rect 25957 37204 25973 37410
rect 25538 37137 25973 37204
rect 28493 37089 28816 37870
rect 28463 37045 28818 37089
rect 28463 36715 28493 37045
rect 28699 36715 28818 37045
rect 28463 36684 28818 36715
rect 10202 36548 10255 36551
rect 10202 36507 10208 36548
rect 10249 36507 10255 36548
rect 31352 36526 31675 37870
rect 10202 36504 10255 36507
rect 9854 36165 9926 36174
rect 9854 36113 9860 36165
rect 9912 36113 9926 36165
rect 9854 36101 9926 36113
rect 1379 35789 1815 35857
rect 23 35305 148 35694
rect 2393 33321 2619 33325
rect 1056 32998 2406 33321
rect 2614 32998 2619 33321
rect 2393 32994 2619 32998
rect 24 32447 149 32836
rect 9874 32566 9926 36101
rect 10214 36079 10255 36504
rect 31332 36496 31691 36526
rect 31332 36290 31352 36496
rect 31675 36290 31691 36496
rect 31332 36273 31691 36290
rect 34211 36177 34534 37870
rect 10200 36069 10262 36079
rect 10200 36028 10213 36069
rect 10254 36028 10262 36069
rect 10200 36020 10262 36028
rect 34180 36054 34556 36177
rect 9866 32563 9929 32566
rect 9866 32511 9870 32563
rect 9922 32511 9929 32563
rect 9866 32506 9929 32511
rect 10214 32464 10255 36020
rect 34180 35849 34211 36054
rect 34534 35849 34556 36054
rect 34180 35815 34556 35849
rect 35615 36108 35956 36140
rect 35615 35785 35645 36108
rect 35844 35785 36279 36108
rect 26447 35719 26889 35780
rect 35615 35736 35956 35785
rect 26447 35687 26471 35719
rect 26693 35687 26889 35719
rect 26447 32769 26889 35687
rect 37183 35235 37308 35624
rect 34774 33249 35006 33257
rect 34774 32926 34790 33249
rect 34999 32926 36278 33249
rect 34774 32920 35006 32926
rect 26444 32757 26891 32769
rect 26444 32648 26455 32757
rect 26883 32648 26891 32757
rect 26444 32637 26891 32648
rect 10209 32461 10257 32464
rect 10209 32417 10213 32461
rect 10254 32417 10257 32461
rect 10209 32414 10257 32417
rect 2784 30462 3007 30470
rect 1057 30139 2796 30462
rect 3004 30139 3007 30462
rect 2784 30124 3007 30139
rect 23 29587 148 29976
rect 3235 27603 3476 27613
rect 1056 27280 3259 27603
rect 3467 27280 3476 27603
rect 3235 27270 3476 27280
rect 25 26728 150 27117
rect 3691 24744 3918 24751
rect 1057 24421 3700 24744
rect 3908 24421 3918 24744
rect 3691 24411 3918 24421
rect 24 23870 149 24259
rect 4127 21885 4352 21891
rect 1056 21562 4134 21885
rect 4342 21562 4352 21885
rect 4127 21554 4352 21562
rect 23 21010 148 21399
rect 4559 19026 4784 19037
rect 1056 18703 4799 19026
rect 4559 18692 4784 18703
rect 24 18152 149 18541
rect 26447 16507 26889 32637
rect 37182 32375 37307 32764
rect 34357 30390 34593 30403
rect 34357 30067 34365 30390
rect 34574 30067 36280 30390
rect 34357 30057 34593 30067
rect 37182 29515 37307 29904
rect 33956 27531 34184 27547
rect 33956 27208 33967 27531
rect 34176 27208 36278 27531
rect 33956 27197 34184 27208
rect 37183 26659 37308 27048
rect 33526 24672 33768 24684
rect 33526 24349 33542 24672
rect 33751 24349 36278 24672
rect 33526 24333 33768 24349
rect 37181 23798 37306 24187
rect 33137 21813 33364 21824
rect 33137 21490 33148 21813
rect 33357 21490 36279 21813
rect 33137 21477 33364 21490
rect 37183 20940 37308 21329
rect 32697 18954 32927 18962
rect 32697 18631 36279 18954
rect 32697 18621 32927 18631
rect 37183 18079 37308 18468
rect 26355 16496 26889 16507
rect 4965 16167 5206 16177
rect 1056 15844 4988 16167
rect 5196 15844 5206 16167
rect 26355 16054 26373 16496
rect 26815 16133 26889 16496
rect 26815 16054 26831 16133
rect 26355 16037 26831 16054
rect 4965 15826 5206 15844
rect 27 15294 152 15683
rect 5393 13308 5639 13315
rect 1056 12985 5639 13308
rect 5393 12980 5639 12985
rect 25 12433 150 12822
rect 5830 10449 6070 10463
rect 1055 10126 5850 10449
rect 6058 10126 6070 10449
rect 5830 10116 6070 10126
rect 24 9574 149 9963
rect 6224 7590 6473 7598
rect 1055 7267 6247 7590
rect 6455 7267 6473 7590
rect 6224 7248 6473 7267
rect 24 6715 149 7104
rect 6671 4731 6906 4741
rect 1057 4408 6691 4731
rect 6899 4408 6906 4731
rect 6671 4395 6906 4408
rect 25 3856 150 4245
rect 7071 1872 7342 1878
rect 1057 1549 7121 1872
rect 7329 1549 7342 1872
rect 7071 1537 7342 1549
rect 25 998 150 1387
<< via1 >>
rect 8655 37073 8978 37298
rect 9874 36945 9926 36982
rect 5796 36624 6119 36849
rect 2754 36197 2979 36520
rect 1601 35857 1787 36180
rect 25634 37204 25957 37410
rect 28493 36715 28699 37045
rect 10208 36507 10249 36548
rect 9860 36113 9912 36165
rect 2406 32998 2614 33321
rect 31352 36290 31675 36496
rect 10213 36028 10254 36069
rect 9870 32511 9922 32563
rect 34211 35849 34534 36054
rect 35645 35785 35844 36108
rect 26471 35687 26693 35719
rect 34790 32926 34999 33249
rect 26455 32648 26883 32757
rect 10213 32417 10254 32461
rect 2796 30139 3004 30462
rect 3259 27280 3467 27603
rect 3700 24421 3908 24744
rect 4134 21562 4342 21885
rect 34365 30067 34574 30390
rect 33967 27208 34176 27531
rect 33542 24349 33751 24672
rect 33148 21490 33357 21813
rect 4988 15844 5196 16167
rect 26373 16054 26815 16496
rect 5850 10126 6058 10449
rect 6247 7267 6455 7590
rect 6691 4408 6899 4731
rect 7121 1549 7329 1872
<< metal2 >>
rect 36872 38502 36991 38503
rect 365 38501 1658 38502
rect 352 38362 1658 38501
rect 35692 38450 36991 38502
rect 35671 38374 36991 38450
rect 352 38210 581 38362
rect 397 38206 581 38210
rect 441 37354 581 38206
rect 36775 38242 36991 38374
rect 1068 37725 1643 37865
rect 35607 37732 36274 37872
rect 1068 37253 1208 37725
rect 25519 37410 25999 37490
rect 8599 37324 9008 37349
rect 8599 37298 12796 37324
rect 8599 37073 8655 37298
rect 8978 37099 12796 37298
rect 25519 37281 25634 37410
rect 24349 37204 25634 37281
rect 25957 37281 25999 37410
rect 25957 37204 26004 37281
rect 8978 37073 9008 37099
rect 24349 37075 26004 37204
rect 36133 37181 36273 37732
rect 36775 37319 36903 38242
rect 36827 37245 36903 37319
rect 8599 37039 9008 37073
rect 28478 37045 28809 37074
rect 9869 36988 9931 36990
rect 9869 36982 12784 36988
rect 9869 36945 9874 36982
rect 9926 36951 12784 36982
rect 9926 36945 9931 36951
rect 9869 36944 9931 36945
rect 5787 36875 6125 36886
rect 5746 36849 12796 36875
rect 28478 36868 28493 37045
rect 5746 36650 5796 36849
rect 5787 36624 5796 36650
rect 6119 36650 12796 36849
rect 24349 36715 28493 36868
rect 28699 36868 28809 37045
rect 28699 36715 28841 36868
rect 24349 36662 28841 36715
rect 6119 36624 6125 36650
rect 5787 36618 6125 36624
rect 10204 36548 10252 36549
rect 2733 36520 2997 36544
rect 2733 36426 2754 36520
rect 2725 36201 2754 36426
rect 2733 36197 2754 36201
rect 2979 36426 2997 36520
rect 10204 36507 10208 36548
rect 10249 36546 10252 36548
rect 10249 36508 12783 36546
rect 10249 36507 10252 36508
rect 10204 36506 10252 36507
rect 31317 36496 31710 36505
rect 31317 36460 31352 36496
rect 2979 36201 12756 36426
rect 24349 36290 31352 36460
rect 31675 36290 31710 36496
rect 24349 36254 31710 36290
rect 31317 36253 31710 36254
rect 2979 36197 2997 36201
rect 1510 36180 1799 36188
rect 2733 36184 2997 36197
rect 1510 35992 1601 36180
rect 1507 35857 1601 35992
rect 1787 35992 1799 36180
rect 9857 36165 9919 36168
rect 9857 36113 9860 36165
rect 9912 36159 9919 36165
rect 9912 36118 12751 36159
rect 9912 36113 9919 36118
rect 9857 36109 9919 36113
rect 35367 36108 35938 36183
rect 10204 36069 10258 36072
rect 10204 36028 10213 36069
rect 10254 36028 12747 36069
rect 34197 36054 34547 36080
rect 10204 36024 10258 36028
rect 34197 36026 34211 36054
rect 1787 35857 12719 35992
rect 1507 35806 12719 35857
rect 24349 35849 34211 36026
rect 34534 36026 34547 36054
rect 34534 35849 34556 36026
rect 24349 35821 34556 35849
rect 35367 35785 35645 36108
rect 35844 35785 35938 36108
rect 24367 35719 26700 35724
rect 24367 35687 26471 35719
rect 26693 35687 26700 35719
rect 24367 35681 26700 35687
rect 35367 35619 35938 35785
rect 35323 35615 35938 35619
rect 24349 35569 35938 35615
rect 2396 35340 12748 35548
rect 24349 35379 35922 35569
rect 2396 33329 2604 35340
rect 34789 35141 34998 35159
rect 2812 34852 12796 35060
rect 24349 34932 34998 35141
rect 2389 33321 2623 33329
rect 2389 32998 2406 33321
rect 2614 32998 2623 33321
rect 2389 32992 2623 32998
rect 2396 32905 2604 32992
rect 2812 30469 3020 34852
rect 2790 30462 3020 30469
rect 2790 30139 2796 30462
rect 3004 30139 3020 30462
rect 2790 30128 3020 30139
rect 2812 30095 3020 30128
rect 3246 34370 12796 34578
rect 24349 34392 34584 34601
rect 3246 27621 3454 34370
rect 3700 33900 12796 34108
rect 24349 33904 34176 34113
rect 3225 27603 3482 27621
rect 3225 27280 3259 27603
rect 3467 27280 3482 27603
rect 3225 27261 3482 27280
rect 3246 27257 3454 27261
rect 3700 24759 3908 33900
rect 4135 33474 12796 33682
rect 3684 24744 3923 24759
rect 3684 24421 3700 24744
rect 3908 24421 3923 24744
rect 3684 24402 3923 24421
rect 3700 24349 3908 24402
rect 4135 21898 4343 33474
rect 24349 33384 33767 33593
rect 4569 33067 12796 33275
rect 4117 21885 4362 21898
rect 4117 21562 4134 21885
rect 4342 21562 4362 21885
rect 4117 21546 4362 21562
rect 4135 21534 4343 21546
rect 4569 19047 4777 33067
rect 24349 32880 33354 33089
rect 4985 32652 12796 32860
rect 26446 32758 26899 32766
rect 24377 32757 26906 32758
rect 4544 18674 4804 19047
rect 4569 18641 4777 18674
rect 4985 16184 5193 32652
rect 24377 32648 26455 32757
rect 26883 32648 26906 32757
rect 24377 32643 26906 32648
rect 26446 32641 26899 32643
rect 9867 32563 9927 32564
rect 9867 32511 9870 32563
rect 9922 32559 9927 32563
rect 9922 32515 12801 32559
rect 9922 32511 9927 32515
rect 9867 32508 9927 32511
rect 10210 32461 10256 32462
rect 10210 32417 10213 32461
rect 10254 32417 12797 32461
rect 10210 32415 10256 32417
rect 5410 32137 12796 32345
rect 24381 32329 32930 32538
rect 4943 16167 5214 16184
rect 4943 15844 4988 16167
rect 5196 15844 5214 16167
rect 4943 15817 5214 15844
rect 4985 15745 5193 15817
rect 5410 13322 5618 32137
rect 5836 31711 12796 31919
rect 5377 12974 5651 13322
rect 5410 12893 5618 12974
rect 5836 10493 6044 31711
rect 6251 31207 12796 31415
rect 5814 10449 6093 10493
rect 5814 10126 5850 10449
rect 6058 10126 6093 10449
rect 5814 10088 6093 10126
rect 5836 10060 6044 10088
rect 6251 7615 6459 31207
rect 6686 30646 12796 30854
rect 6202 7590 6485 7615
rect 6202 7267 6247 7590
rect 6455 7267 6485 7590
rect 6202 7237 6485 7267
rect 6251 7181 6459 7237
rect 6686 4757 6894 30646
rect 7102 30176 12796 30384
rect 6651 4731 6916 4757
rect 6651 4408 6691 4731
rect 6899 4408 6916 4731
rect 6651 4385 6916 4408
rect 6686 4384 6894 4385
rect 7102 1887 7310 30176
rect 7083 1872 7350 1887
rect 7083 1549 7121 1872
rect 7329 1549 7350 1872
rect 7083 1534 7350 1549
rect 13256 951 13590 30190
rect 14222 521 14424 30180
rect 14628 678 14830 30180
rect 14628 522 14831 678
rect 15025 677 15227 30180
rect 15425 677 15627 30180
rect 14628 521 14830 522
rect 15024 521 15227 677
rect 15424 521 15627 677
rect 15830 521 16032 30180
rect 16231 678 16433 30180
rect 16230 522 16433 678
rect 16231 521 16433 522
rect 16631 521 16833 30180
rect 17040 521 17242 30180
rect 17453 677 17655 30180
rect 17853 677 18055 30180
rect 18249 677 18451 30180
rect 17452 521 17655 677
rect 17852 521 18055 677
rect 18248 521 18451 677
rect 18654 678 18856 30180
rect 18654 522 18857 678
rect 18654 521 18856 522
rect 19063 521 19265 30180
rect 19464 676 19666 30180
rect 19868 677 20070 30180
rect 19464 521 19667 676
rect 19868 521 20071 677
rect 20277 675 20479 30180
rect 20277 521 20480 675
rect 20682 521 20884 30180
rect 21079 521 21281 30180
rect 21491 521 21693 30180
rect 19465 520 19667 521
rect 20278 519 20480 521
rect 21904 520 22106 30180
rect 22305 521 22507 30180
rect 22706 689 22908 30180
rect 22706 523 22910 689
rect 23115 687 23317 30180
rect 23115 521 23318 687
rect 23532 521 23734 30180
rect 23932 687 24134 30180
rect 24333 687 24535 30180
rect 24729 687 24931 30180
rect 23932 521 24135 687
rect 24330 521 24535 687
rect 24728 521 24931 687
rect 25134 687 25336 30180
rect 25540 687 25742 30180
rect 32721 19186 32930 32329
rect 33145 21833 33354 32880
rect 33558 24681 33767 33384
rect 33967 27558 34176 33904
rect 34375 30408 34584 34392
rect 34789 33264 34998 34932
rect 34769 33249 35012 33264
rect 34769 32926 34790 33249
rect 34999 32926 35012 33249
rect 34769 32910 35012 32926
rect 34789 32843 34998 32910
rect 34351 30390 34602 30408
rect 34351 30067 34365 30390
rect 34574 30067 34602 30390
rect 34351 30051 34602 30067
rect 33947 27531 34199 27558
rect 33947 27208 33967 27531
rect 34176 27208 34199 27531
rect 33947 27187 34199 27208
rect 33967 27184 34176 27187
rect 33531 24672 33767 24681
rect 33531 24349 33542 24672
rect 33751 24349 33767 24672
rect 33531 24339 33767 24349
rect 33558 24268 33767 24339
rect 33128 21813 33371 21833
rect 33128 21490 33148 21813
rect 33357 21490 33371 21813
rect 33128 21462 33371 21490
rect 32722 18996 32930 19186
rect 32722 18984 32931 18996
rect 32711 18978 32931 18984
rect 32685 18610 32938 18978
rect 32711 18608 32920 18610
rect 36829 17339 36903 17373
rect 36131 17236 36271 17314
rect 36763 17299 36904 17339
rect 36130 17224 36271 17236
rect 36765 17230 36903 17299
rect 36129 17209 36271 17224
rect 36129 17119 36270 17209
rect 36764 17113 36904 17230
rect 26362 16496 26822 16501
rect 26362 16054 26373 16496
rect 26815 16423 26822 16496
rect 26815 16255 36277 16423
rect 26815 16126 36290 16255
rect 26815 16054 26822 16126
rect 26362 16044 26822 16054
rect 25134 521 25338 687
rect 25540 521 25744 687
rect 438 33 578 230
rect 1068 0 1208 366
use sky130_hilas_TopProtection  sky130_hilas_TopProtection_0
timestamp 1626559870
transform 1 0 1616 0 1 37623
box -2 -76 34131 1170
use sky130_hilas_LeftProtection  sky130_hilas_LeftProtection_0
timestamp 1626559870
transform 1 0 2213 0 1 8665
box -2065 -8439 -833 28728
use sky130_hilas_RightProtection  sky130_hilas_RightProtection_0
timestamp 1626559870
transform 1 0 38009 0 1 8593
box -2054 8715 -826 28728
use sky130_hilas_TopLevelTextStructure  sky130_hilas_TopLevelTextStructure_0
timestamp 1626912190
transform 1 0 12501 0 1 30961
box 218 -793 13243 6785
<< labels >>
rlabel metal1 37183 18079 37308 18468 0 IO07
port 1 nsew
rlabel metal1 37183 20940 37308 21329 0 IO08
port 2 nsew
rlabel metal1 37181 23798 37306 24187 0 IO09
port 3 nsew
rlabel metal1 37183 26659 37308 27048 0 IO10
port 4 nsew
rlabel metal1 37182 29515 37307 29904 0 IO11
port 5 nsew
rlabel metal1 37182 32375 37307 32764 0 IO12
port 6 nsew
rlabel metal1 37183 35235 37308 35624 0 IO13
port 7 nsew
rlabel metal1 23 35305 148 35694 0 IO25
port 8 nsew
rlabel metal1 24 32447 149 32836 0 IO26
port 9 nsew
rlabel metal1 23 29587 148 29976 0 IO27
port 10 nsew
rlabel metal1 25 26728 150 27117 0 IO28
port 11 nsew
rlabel metal1 24 23870 149 24259 0 IO29
port 12 nsew
rlabel metal1 23 21010 148 21399 0 IO30
port 13 nsew
rlabel metal1 24 18152 149 18541 0 IO31
port 14 nsew
rlabel metal1 27 15294 152 15683 0 IO32
port 15 nsew
rlabel metal1 25 12433 150 12822 0 IO33
port 16 nsew
rlabel metal1 24 9574 149 9963 0 IO34
port 17 nsew
rlabel metal1 24 6715 149 7104 0 IO35
port 18 nsew
rlabel metal1 25 3856 150 4245 0 IO36
port 19 nsew
rlabel metal1 25 998 150 1387 0 IO37
port 20 nsew
rlabel metal2 352 38210 520 38501 0 VSSA1
port 21 nsew
rlabel metal1 2385 38791 2774 38908 0 ANALOG10
port 22 nsew
rlabel metal1 5244 38790 5633 38907 0 ANALOG09
port 23 nsew
rlabel metal1 8103 38790 8492 38907 0 ANALOG08
port 24 nsew
rlabel metal1 12293 38793 12682 38910 0 ANALOG07
port 25 nsew
rlabel metal1 16505 38791 16894 38908 0 ANALOG06
port 26 nsew
rlabel metal1 19364 38791 19753 38908 0 ANALOG05
port 27 nsew
rlabel metal1 22224 38791 22613 38908 0 ANALOG04
port 28 nsew
rlabel metal1 25083 38791 25472 38908 0 ANALOG03
port 29 nsew
rlabel metal1 27942 38791 28331 38908 0 ANALOG02
port 30 nsew
rlabel metal1 30801 38790 31190 38907 0 ANALOG01
port 31 nsew
rlabel metal1 33660 38790 34049 38907 0 ANALOG00
port 32 nsew
rlabel metal2 36872 38245 36991 38503 0 VSSA1
port 33 nsew
rlabel metal2 1068 0 1208 140 0 VDDA1
port 34 nsew
rlabel metal2 438 33 578 173 0 VSSA1
port 33 nsew
rlabel metal2 36130 17119 36270 17236 0 VDDA1
port 34 nsew
rlabel metal2 36764 17113 36904 17230 0 VSSA1
port 33 nsew
rlabel metal2 14222 521 14424 677 0 LADATAOUT00
port 36 nsew
rlabel metal2 14629 522 14831 678 0 LADATAOUT01
port 35 nsew
rlabel metal2 15024 521 15226 677 0 LADATAOUT02
port 37 nsew
rlabel metal2 15424 521 15626 677 0 LADATAOUT03
port 38 nsew
rlabel metal2 15830 521 16032 677 0 LADATAOUT04
port 39 nsew
rlabel metal2 16230 522 16432 678 0 LADATAOUT05
port 40 nsew
rlabel metal2 16631 521 16833 677 0 LADATAOUT06
port 41 nsew
rlabel metal2 17040 521 17242 677 0 LADATAOUT07
port 42 nsew
rlabel metal2 17452 521 17654 677 0 LADATAOUT08
port 43 nsew
rlabel metal2 17852 521 18054 677 0 LADATAOUT09
port 44 nsew
rlabel metal2 18248 521 18450 677 0 LADATAOUT10
port 45 nsew
rlabel metal2 18655 522 18857 678 0 LADATAOUT11
port 46 nsew
rlabel metal2 19063 521 19265 677 0 LADATAOUT12
port 47 nsew
rlabel metal2 19465 520 19667 676 0 LADATAOUT13
port 48 nsew
rlabel metal2 19869 521 20071 677 0 LADATAOUT14
port 49 nsew
rlabel metal2 20278 519 20480 675 0 LADATAOUT15
port 50 nsew
rlabel metal2 20682 521 20884 677 0 LADATA16
port 51 nsew
rlabel metal2 21079 521 21281 677 0 LADATAOUT17
port 52 nsew
rlabel metal2 21491 522 21693 678 0 LADATAOUT18
port 53 nsew
rlabel metal2 21904 520 22106 676 0 LADATAOUT19
port 54 nsew
rlabel metal2 22305 521 22507 677 0 LADATAOUT20
port 55 nsew
rlabel metal2 22706 523 22910 689 0 LADATAOUT21
port 56 nsew
rlabel metal2 23115 521 23318 687 0 LADATAOUT22
port 57 nsew
rlabel metal2 23530 521 23733 687 0 LADATAOUT23
port 58 nsew
rlabel metal2 23932 521 24135 687 0 LADATAOUT24
port 59 nsew
rlabel metal2 24330 521 24533 687 0 LADATAIN00
port 60 nsew
rlabel metal2 24728 521 24931 687 0 LADATAIN01
port 61 nsew
rlabel metal2 25135 521 25338 687 0 LADATAIN02
port 62 nsew
rlabel metal2 25541 521 25744 687 0 LADATAIN03
port 63 nsew
rlabel metal2 36174 16126 36290 16252 0 VCCA
port 64 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
