magic
tech sky130A
timestamp 1628704368
<< checkpaint >>
rect -107 994 1232 998
rect -592 -337 1232 994
rect -592 -341 747 -337
<< metal2 >>
rect 0 527 578 545
rect 0 484 578 502
rect 3 384 578 402
rect 3 341 578 359
rect 2 279 29 307
rect 542 283 579 311
rect 3 226 578 243
rect 3 184 578 201
rect 3 86 578 103
rect 3 42 578 59
<< metal3 >>
rect 145 332 172 333
rect 145 257 559 332
<< metal4 >>
rect 258 320 302 404
rect 116 319 217 320
rect 257 319 303 320
rect 45 269 303 319
rect 45 268 152 269
rect 257 203 303 269
rect 257 153 305 203
rect 302 123 305 153
use sky130_hilas_m22m4  sky130_hilas_m22m4_1
timestamp 1628704359
transform 1 0 523 0 1 293
box 0 0 79 75
use sky130_hilas_m22m4  sky130_hilas_m22m4_0
timestamp 1628704359
transform 1 0 38 0 1 289
box 0 0 79 75
use sky130_hilas_CapModule01  sky130_hilas_CapModule01_1
timestamp 1607800460
transform 1 0 588 0 1 546
box -443 -245 -159 41
use sky130_hilas_CapModule01  sky130_hilas_CapModule01_0
timestamp 1607800460
transform 1 0 588 0 1 245
box -443 -245 -159 41
<< labels >>
rlabel metal2 2 279 9 307 0 CAPTERM01
port 2 nsew analog default
rlabel metal2 571 283 579 311 0 CAPTERM02
port 1 nsew analog default
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
