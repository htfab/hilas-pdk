magic
tech sky130A
timestamp 1628178864
<< error_s >>
rect -138 -59 -98 -54
rect 88 -59 128 -52
rect -138 -101 -98 -96
rect 88 -101 128 -94
rect -62 -126 -22 -120
rect 88 -126 128 -120
rect -62 -168 -22 -162
rect 88 -168 128 -162
<< nwell >>
rect -251 -102 25 -25
rect -251 -119 -52 -102
rect -251 -181 -53 -119
rect -251 -186 25 -181
<< pmos >>
rect -138 -96 -98 -59
<< pdiff >>
rect -167 -71 -138 -59
rect -167 -88 -161 -71
rect -144 -88 -138 -71
rect -167 -96 -138 -88
rect -98 -71 -70 -59
rect -98 -88 -92 -71
rect -75 -88 -70 -71
rect -98 -96 -70 -88
<< pdiffc >>
rect -161 -88 -144 -71
rect -92 -88 -75 -71
<< nsubdiff >>
rect -227 -130 -195 -117
rect -227 -147 -220 -130
rect -203 -147 -195 -130
rect -227 -159 -195 -147
<< nsubdiffcont >>
rect -220 -147 -203 -130
<< poly >>
rect -234 -51 25 -36
rect -138 -59 -98 -51
rect -52 -83 -19 -77
rect -138 -118 -98 -96
rect -52 -100 -44 -83
rect -27 -100 -19 -83
rect -52 -112 -19 -100
<< polycont >>
rect -44 -100 -27 -83
<< locali >>
rect -101 -71 25 -70
rect -171 -83 -161 -71
rect -188 -88 -161 -83
rect -144 -88 -136 -71
rect -101 -88 -92 -71
rect -75 -83 25 -71
rect -75 -88 -44 -83
rect -188 -96 -169 -88
rect -190 -99 -169 -96
rect -191 -100 -169 -99
rect -52 -100 -44 -88
rect -27 -88 25 -83
rect -27 -100 -19 -88
rect -203 -105 -169 -100
rect -216 -108 -169 -105
rect -220 -111 -169 -108
rect -220 -117 -171 -111
rect -220 -122 -186 -117
rect -220 -124 -194 -122
rect -220 -126 -197 -124
rect -220 -130 -199 -126
rect -220 -158 -203 -147
<< metal1 >>
rect -189 -186 -169 -25
rect 162 -29 181 -25
rect 162 -186 181 -181
<< metal2 >>
rect -263 -72 -202 -52
rect 206 -72 213 -52
rect -176 -150 -64 -149
rect -263 -170 -64 -150
rect -176 -171 -64 -170
use sky130_hilas_poly2m1  sky130_hilas_poly2m1_0
timestamp 1628178864
transform 1 0 -236 0 1 -65
box -9 -26 24 25
use sky130_hilas_li2m1  sky130_hilas_li2m1_2
timestamp 1628178864
transform 1 0 -180 0 1 -86
box -10 -8 13 21
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1628178864
transform 1 0 -225 0 1 -62
box -9 -10 23 22
use sky130_hilas_TgateSingle01Part1  sky130_hilas_TgateSingle01Part1_0
timestamp 1628178864
transform 1 0 -232 0 1 0
box 257 -181 445 -29
use sky130_hilas_TgateSingle01Part2  sky130_hilas_TgateSingle01Part2_0
timestamp 1628178864
transform 1 0 -71 0 1 0
box -67 -181 96 -38
<< labels >>
rlabel metal2 -263 -72 -254 -52 0 Select
rlabel metal2 -263 -170 -254 -150 0 Input
<< end >>
