magic
tech sky130A
timestamp 1634057848
<< checkpaint >>
rect -367 -630 1369 1677
<< error_s >>
rect 201 820 241 826
rect 351 820 391 826
rect 201 778 241 784
rect 351 778 391 784
rect 125 754 165 759
rect 351 752 391 759
rect 125 712 165 717
rect 351 710 391 717
rect 125 650 165 655
rect 351 650 391 657
rect 125 608 165 613
rect 351 608 391 615
rect 201 583 241 589
rect 351 583 391 589
rect 201 541 241 547
rect 351 541 391 547
rect 201 500 241 506
rect 351 500 391 506
rect 201 458 241 464
rect 351 458 391 464
rect 125 434 165 439
rect 351 432 391 439
rect 125 392 165 397
rect 351 390 391 397
rect 125 330 165 335
rect 351 330 391 337
rect 125 288 165 293
rect 351 288 391 295
rect 201 263 241 269
rect 351 263 391 269
rect 201 221 241 227
rect 351 221 391 227
<< nwell >>
rect 12 752 13 790
<< metal1 >>
rect 74 827 94 831
rect 425 825 444 831
rect 74 226 94 230
rect 425 226 444 232
<< metal2 >>
rect 0 808 5 828
rect 0 710 6 730
rect 469 710 476 730
rect 0 637 6 657
rect 469 637 476 657
rect 0 539 5 559
rect 0 488 5 508
rect 0 390 6 410
rect 469 390 476 410
rect 0 317 6 337
rect 469 317 476 337
rect 0 219 5 239
use sky130_hilas_TgateSingle01  sky130_hilas_TgateSingle01_3
timestamp 1634057785
transform 1 0 263 0 1 709
box 0 0 476 338
use sky130_hilas_TgateSingle01  sky130_hilas_TgateSingle01_0
timestamp 1634057785
transform 1 0 263 0 -1 658
box 0 0 476 338
use sky130_hilas_TgateSingle01  sky130_hilas_TgateSingle01_2
timestamp 1634057785
transform 1 0 263 0 -1 338
box 0 0 476 338
use sky130_hilas_TgateSingle01  sky130_hilas_TgateSingle01_1
timestamp 1634057785
transform 1 0 263 0 1 389
box 0 0 476 338
<< labels >>
rlabel metal2 0 637 6 657 0 SELECT2
port 7 nsew analog default
rlabel metal1 74 226 94 230 0 VPWR
port 2 nsew analog default
rlabel metal2 0 539 5 559 0 INPUT1_2
port 6 nsew analog default
rlabel metal1 425 825 444 831 0 VGND
port 10 nsew ground default
rlabel metal1 425 226 444 232 0 VGND
port 10 nsew ground default
rlabel metal2 469 637 476 657 0 OUTPUT2
port 12 nsew analog default
rlabel metal1 74 827 94 831 0 VPWR
port 2 nsew power default
rlabel metal2 469 317 476 337 0 OUTPUT4
port 14 nsew
rlabel metal2 469 390 476 410 0 OUTPUT3
port 15 nsew
rlabel metal2 469 710 476 730 0 OUTPUT1
port 16 nsew
rlabel metal2 0 219 5 239 0 INPUT1_4
port 17 nsew
rlabel metal2 0 317 6 337 0 SELECT4
port 18 nsew
rlabel metal2 0 390 6 410 0 SELECT3
port 19 nsew
rlabel metal2 0 488 5 508 0 INPUT1_3
port 20 nsew
rlabel metal2 0 710 6 730 0 SELECT1
port 21 nsew
rlabel metal2 0 808 5 828 0 INPUT1_1
port 22 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
