magic
tech sky130A
timestamp 1628707293
<< checkpaint >>
rect 822 1537 2255 1681
rect 819 1387 2255 1537
rect 138 1316 2255 1387
rect -149 1096 2255 1316
rect -629 -184 2255 1096
rect -629 -350 1927 -184
rect -150 -615 1927 -350
rect 411 -630 1927 -615
<< error_s >>
rect 531 658 560 686
rect 610 658 639 686
rect 689 658 718 686
rect 509 651 739 658
rect 509 636 516 651
rect 531 645 560 651
rect 610 645 639 651
rect 689 645 718 651
rect 531 636 532 637
rect 559 636 560 637
rect 610 636 611 637
rect 638 636 639 637
rect 689 636 690 637
rect 717 636 718 637
rect 732 636 739 651
rect 481 607 522 636
rect 530 635 561 636
rect 609 635 640 636
rect 688 635 719 636
rect 531 608 560 635
rect 610 608 639 635
rect 689 608 718 635
rect 530 607 561 608
rect 609 607 640 608
rect 688 607 719 608
rect 726 607 768 636
rect 58 578 64 584
rect 111 578 117 584
rect 509 557 516 607
rect 531 606 532 607
rect 559 606 560 607
rect 610 606 611 607
rect 638 606 639 607
rect 689 606 690 607
rect 717 606 718 607
rect 732 579 739 607
rect 531 557 532 558
rect 559 557 560 558
rect 610 557 611 558
rect 638 557 639 558
rect 689 557 690 558
rect 717 557 718 558
rect 732 557 739 563
rect 752 562 753 563
rect 52 528 58 534
rect 117 528 123 534
rect 481 528 522 557
rect 530 556 561 557
rect 609 556 640 557
rect 688 556 719 557
rect 531 529 560 556
rect 610 529 639 556
rect 689 529 718 556
rect 530 528 561 529
rect 609 528 640 529
rect 688 528 719 529
rect 726 528 768 557
rect 509 519 516 528
rect 531 527 532 528
rect 559 527 560 528
rect 610 527 611 528
rect 638 527 639 528
rect 689 527 690 528
rect 717 527 718 528
rect 522 519 726 522
rect 732 519 739 528
rect 509 506 739 519
rect 531 505 560 506
rect 610 505 639 506
rect 689 505 718 506
rect 509 498 739 505
rect 509 483 516 498
rect 531 492 560 498
rect 610 492 639 498
rect 689 492 718 498
rect 570 484 596 490
rect 531 483 532 484
rect 559 483 560 484
rect 610 483 611 484
rect 638 483 639 484
rect 689 483 690 484
rect 717 483 718 484
rect 732 483 739 498
rect 58 469 64 475
rect 111 469 117 475
rect 481 454 522 483
rect 530 482 561 483
rect 609 482 640 483
rect 688 482 719 483
rect 531 455 560 482
rect 571 470 597 476
rect 610 455 639 482
rect 689 455 718 482
rect 530 454 561 455
rect 609 454 640 455
rect 688 454 719 455
rect 726 454 768 483
rect 52 419 58 425
rect 117 419 123 425
rect 509 404 516 454
rect 531 453 532 454
rect 559 453 560 454
rect 610 453 611 454
rect 638 453 639 454
rect 689 453 690 454
rect 717 453 718 454
rect 732 436 739 454
rect 531 404 532 405
rect 559 404 560 405
rect 610 404 611 405
rect 638 404 639 405
rect 689 404 690 405
rect 717 404 718 405
rect 732 404 739 419
rect 481 375 522 404
rect 530 403 561 404
rect 609 403 640 404
rect 688 403 719 404
rect 531 376 560 403
rect 610 376 639 403
rect 689 376 718 403
rect 530 375 561 376
rect 609 375 640 376
rect 688 375 719 376
rect 726 375 768 404
rect 509 363 516 375
rect 531 374 532 375
rect 559 374 560 375
rect 610 374 611 375
rect 638 374 639 375
rect 689 374 690 375
rect 717 374 718 375
rect 530 363 560 366
rect 609 363 639 366
rect 688 363 718 366
rect 732 363 739 375
rect 509 353 739 363
rect 530 349 560 353
rect 609 349 639 353
rect 688 349 718 353
rect 508 342 738 349
rect 508 327 515 342
rect 530 336 560 342
rect 609 336 639 342
rect 688 336 718 342
rect 570 331 596 334
rect 530 327 531 328
rect 558 327 559 328
rect 609 327 610 328
rect 637 327 638 328
rect 688 327 689 328
rect 716 327 717 328
rect 731 327 738 342
rect 480 298 521 327
rect 529 326 560 327
rect 608 326 639 327
rect 687 326 718 327
rect 530 299 559 326
rect 570 317 596 320
rect 609 299 638 326
rect 688 299 717 326
rect 529 298 560 299
rect 608 298 639 299
rect 687 298 718 299
rect 725 298 767 327
rect 58 280 64 286
rect 111 280 117 286
rect 508 248 515 298
rect 530 297 531 298
rect 558 297 559 298
rect 609 297 610 298
rect 637 297 638 298
rect 688 297 689 298
rect 716 297 717 298
rect 731 278 738 298
rect 530 248 531 249
rect 558 248 559 249
rect 609 248 610 249
rect 637 248 638 249
rect 688 248 689 249
rect 716 248 717 249
rect 731 248 738 261
rect 52 230 58 236
rect 117 230 123 236
rect 480 219 521 248
rect 529 247 560 248
rect 608 247 639 248
rect 687 247 718 248
rect 530 220 559 247
rect 609 220 638 247
rect 688 220 717 247
rect 529 219 560 220
rect 608 219 639 220
rect 687 219 718 220
rect 725 219 767 248
rect 508 209 515 219
rect 530 218 531 219
rect 558 218 559 219
rect 609 218 610 219
rect 637 218 638 219
rect 688 218 689 219
rect 716 218 717 219
rect 521 210 725 212
rect 530 209 559 210
rect 609 209 638 210
rect 688 209 717 210
rect 731 209 738 219
rect 508 197 738 209
rect 530 195 559 197
rect 609 195 638 197
rect 688 195 717 197
rect 508 188 738 195
rect 508 173 515 188
rect 530 182 559 188
rect 609 182 638 188
rect 688 182 717 188
rect 569 175 595 180
rect 530 173 531 174
rect 558 173 559 174
rect 609 173 610 174
rect 637 173 638 174
rect 688 173 689 174
rect 716 173 717 174
rect 731 173 738 188
rect 58 163 64 169
rect 111 163 117 169
rect 480 144 521 173
rect 529 172 560 173
rect 608 172 639 173
rect 687 172 718 173
rect 530 145 559 172
rect 570 161 596 166
rect 609 145 638 172
rect 688 145 717 172
rect 529 144 560 145
rect 608 144 639 145
rect 687 144 718 145
rect 725 144 767 173
rect 52 113 58 119
rect 117 113 123 119
rect 508 94 515 144
rect 530 143 531 144
rect 558 143 559 144
rect 609 143 610 144
rect 637 143 638 144
rect 688 143 689 144
rect 716 143 717 144
rect 731 136 738 144
rect 530 94 531 95
rect 558 94 559 95
rect 609 94 610 95
rect 637 94 638 95
rect 688 94 689 95
rect 716 94 717 95
rect 731 94 738 119
rect 480 65 521 94
rect 529 93 560 94
rect 608 93 639 94
rect 687 93 718 94
rect 530 66 559 93
rect 609 66 638 93
rect 688 66 717 93
rect 529 65 560 66
rect 608 65 639 66
rect 687 65 718 66
rect 725 65 767 94
rect 508 50 515 65
rect 530 64 531 65
rect 558 64 559 65
rect 609 64 610 65
rect 637 64 638 65
rect 688 64 689 65
rect 716 64 717 65
rect 530 50 559 56
rect 609 50 638 56
rect 688 50 717 56
rect 731 50 738 65
rect 508 43 738 50
rect 530 15 559 43
rect 609 15 638 43
rect 688 15 717 43
<< nwell >>
rect 896 356 931 357
rect 896 340 913 356
rect 930 340 931 356
<< poly >>
rect 717 575 753 579
rect 157 542 394 566
rect 717 563 752 575
rect 157 433 392 457
rect 717 419 752 436
rect 913 356 931 357
rect 929 340 931 356
rect 157 253 394 277
rect 584 261 752 278
rect 159 133 396 157
rect 584 119 752 136
<< polycont >>
rect 896 340 913 357
<< locali >>
rect 887 340 896 357
<< viali >>
rect 913 340 931 357
<< metal1 >>
rect 36 46 76 645
rect 918 360 931 362
rect 910 357 934 360
rect 910 340 913 357
rect 931 340 934 357
rect 910 337 934 340
rect 920 333 931 337
<< metal2 >>
rect 0 594 761 601
rect 0 583 764 594
rect 0 540 974 558
rect 0 452 761 458
rect 0 440 764 452
rect 0 408 760 415
rect 0 397 764 408
rect 2 282 764 299
rect 2 240 764 257
rect 2 142 764 159
rect 80 133 234 142
rect 2 98 764 115
use sky130_hilas_overlapCap01  sky130_hilas_overlapCap01_2
timestamp 1628705746
transform 1 0 767 0 1 240
box 0 0 287 208
use sky130_hilas_overlapCap01  sky130_hilas_overlapCap01_3
timestamp 1628705746
transform 1 0 767 0 1 86
box 0 0 287 208
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_1
timestamp 1628705728
transform 1 0 1041 0 1 0
box 0 0 256 191
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_2
timestamp 1628705728
transform 1 0 1041 0 -1 397
box 0 0 256 191
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_0
timestamp 1628705728
transform 1 0 1041 0 1 300
box 0 0 256 191
use sky130_hilas_overlapCap01  sky130_hilas_overlapCap01_1
timestamp 1628705746
transform 1 0 768 0 1 396
box 0 0 287 208
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_3
timestamp 1628705728
transform 1 0 1041 0 -1 698
box 0 0 256 191
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_1
timestamp 1628707260
transform 1 0 1452 0 1 446
box 0 0 173 190
use sky130_hilas_overlapCap01  sky130_hilas_overlapCap01_0
timestamp 1628705746
transform 1 0 768 0 1 549
box 0 0 287 208
use sky130_hilas_wellContact  sky130_hilas_wellContact_1
timestamp 1628705669
transform 1 0 1449 0 1 721
box 0 0 173 186
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_2
timestamp 1628707260
transform 1 0 1452 0 1 752
box 0 0 173 190
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_0
timestamp 1628707260
transform 1 0 1452 0 1 563
box 0 0 173 190
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_3
timestamp 1628707260
transform 1 0 1452 0 1 861
box 0 0 173 190
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
