magic
tech sky130A
timestamp 1629137245
<< checkpaint >>
rect 492 2079 2301 2123
rect -630 1750 2301 2079
rect -630 -233 2488 1750
rect 648 -256 2488 -233
rect 648 -630 2457 -256
<< error_s >>
rect 58 976 64 982
rect 111 976 117 982
rect 52 926 58 932
rect 117 926 123 932
rect 481 917 487 923
rect 586 917 592 923
rect 475 867 481 873
rect 592 867 598 873
rect 481 616 487 622
rect 586 616 592 622
rect 58 562 64 568
rect 111 562 117 568
rect 475 566 481 572
rect 592 566 598 572
rect 52 512 58 518
rect 117 512 123 518
<< nwell >>
rect 1665 1031 1792 1049
rect 1145 875 1311 897
rect 1191 714 1219 738
rect 1664 444 1792 463
<< locali >>
rect 283 783 329 792
rect 283 766 286 783
rect 303 766 329 783
rect 283 714 329 766
rect 283 697 286 714
rect 303 697 329 714
rect 283 691 329 697
<< viali >>
rect 286 766 303 783
rect 286 697 303 714
<< metal1 >>
rect 35 1042 77 1049
rect 405 1041 428 1049
rect 1057 1041 1076 1049
rect 1101 1041 1129 1049
rect 1596 1035 1630 1049
rect 1663 1034 1690 1049
rect 279 788 317 792
rect 279 695 283 788
rect 312 695 317 788
rect 279 691 317 695
rect 1596 444 1630 463
rect 1663 444 1690 465
<< via1 >>
rect 1600 883 1626 909
rect 283 783 312 788
rect 283 766 286 783
rect 286 766 303 783
rect 303 766 312 783
rect 283 714 312 766
rect 283 697 286 714
rect 286 697 303 714
rect 303 697 312 714
rect 283 695 312 697
<< metal2 >>
rect 1343 1022 1368 1048
rect 0 981 7 999
rect 1449 924 1474 961
rect 1596 909 1630 913
rect 1596 904 1600 909
rect 1145 875 1311 897
rect 1361 885 1600 904
rect 1361 828 1380 885
rect 1596 883 1600 885
rect 1626 883 1630 909
rect 1596 880 1630 883
rect 1452 839 1473 868
rect 282 809 1380 828
rect 282 791 301 809
rect 280 788 315 791
rect 280 695 283 788
rect 312 695 315 788
rect 1777 778 1792 800
rect 1347 755 1372 778
rect 1191 714 1219 738
rect 1777 696 1792 718
rect 280 692 315 695
rect 1296 631 1473 651
rect 1139 582 1155 622
rect 1267 550 1473 571
rect 0 496 8 511
rect 1187 446 1213 471
use sky130_hilas_FGBias2x1cell  sky130_hilas_FGBias2x1cell_0
timestamp 1628285143
transform 1 0 396 0 1 826
box -396 -429 1258 623
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_0
timestamp 1628285143
transform 1 0 989 0 1 884
box 133 -454 682 609
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1628285143
transform 1 0 1145 0 -1 609
box 133 -454 682 609
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1628285143
transform 1 0 1637 0 1 485
box -172 -111 221 635
<< labels >>
rlabel metal1 1596 444 1630 450 0 VGND
port 7 nsew ground default
rlabel metal1 1663 444 1690 450 0 VPWR
port 8 nsew power default
rlabel metal1 1596 1044 1630 1049 0 VGND
port 7 nsew ground default
rlabel metal1 1663 1044 1690 1049 0 VPWR
port 8 nsew power default
rlabel metal2 1347 755 1372 778 0 VIN21
port 3 nsew
rlabel metal2 1187 446 1210 471 0 VIN12
port 2 nsew analog default
rlabel metal2 1343 1022 1368 1048 0 VIN22
port 4 nsew
rlabel metal2 1777 696 1792 718 0 OUTPUT1
port 5 nsew
rlabel metal2 1777 778 1792 800 0 OUTPUT2
port 6 nsew
rlabel metal1 1057 1041 1076 1049 0 COLSEL1
port 1 nsew
rlabel metal2 0 981 7 999 0 DRAIN1
port 9 nsew
rlabel metal2 0 496 8 511 0 DRAIN2
port 10 nsew
rlabel metal1 35 1042 77 1049 0 VTUN
port 11 nsew
rlabel metal1 405 1041 428 1049 0 GATE1
port 12 nsew
rlabel metal1 1101 1041 1129 1049 0 VINJ
port 13 nsew
rlabel metal2 1191 714 1214 738 0 VIN11
port 14 nsew
<< end >>
