magic
tech sky130A
timestamp 1607392100
<< error_s >>
rect -678 1300 -649 1316
rect -599 1300 -570 1316
rect -520 1300 -491 1316
rect -441 1300 -412 1316
rect -195 1302 -166 1320
rect -39 1302 -10 1320
rect 207 1300 236 1316
rect 286 1300 315 1316
rect 365 1300 394 1316
rect 444 1300 473 1316
rect -195 1270 -194 1271
rect -167 1270 -166 1271
rect -39 1270 -38 1271
rect -11 1270 -10 1271
rect -678 1266 -677 1267
rect -650 1266 -649 1267
rect -599 1266 -598 1267
rect -571 1266 -570 1267
rect -520 1266 -519 1267
rect -492 1266 -491 1267
rect -441 1266 -440 1267
rect -413 1266 -412 1267
rect -728 1237 -711 1266
rect -679 1265 -648 1266
rect -600 1265 -569 1266
rect -521 1265 -490 1266
rect -442 1265 -411 1266
rect -678 1258 -649 1265
rect -599 1258 -570 1265
rect -520 1258 -491 1265
rect -441 1258 -412 1265
rect -678 1244 -669 1258
rect -422 1244 -412 1258
rect -678 1238 -649 1244
rect -599 1238 -570 1244
rect -520 1238 -491 1244
rect -441 1238 -412 1244
rect -679 1237 -648 1238
rect -600 1237 -569 1238
rect -521 1237 -490 1238
rect -442 1237 -411 1238
rect -380 1237 -362 1266
rect -245 1241 -227 1270
rect -196 1269 -165 1270
rect -195 1260 -166 1269
rect -195 1251 -185 1260
rect -176 1251 -166 1260
rect -195 1242 -166 1251
rect -196 1241 -165 1242
rect -134 1241 -116 1270
rect -89 1241 -71 1270
rect -40 1269 -9 1270
rect -39 1260 -10 1269
rect -39 1251 -29 1260
rect -20 1251 -10 1260
rect -39 1242 -10 1251
rect -40 1241 -9 1242
rect 22 1241 40 1270
rect 207 1266 208 1267
rect 235 1266 236 1267
rect 286 1266 287 1267
rect 314 1266 315 1267
rect 365 1266 366 1267
rect 393 1266 394 1267
rect 444 1266 445 1267
rect 472 1266 473 1267
rect -195 1240 -194 1241
rect -167 1240 -166 1241
rect -39 1240 -38 1241
rect -11 1240 -10 1241
rect 157 1237 175 1266
rect 206 1265 237 1266
rect 285 1265 316 1266
rect 364 1265 395 1266
rect 443 1265 474 1266
rect 207 1258 236 1265
rect 286 1258 315 1265
rect 365 1258 394 1265
rect 444 1258 473 1265
rect 207 1244 217 1258
rect 464 1244 473 1258
rect 207 1238 236 1244
rect 286 1238 315 1244
rect 365 1238 394 1244
rect 444 1238 473 1244
rect 206 1237 237 1238
rect 285 1237 316 1238
rect 364 1237 395 1238
rect 443 1237 474 1238
rect 506 1237 523 1266
rect 540 1244 542 1245
rect -678 1236 -677 1237
rect -650 1236 -649 1237
rect -599 1236 -598 1237
rect -571 1236 -570 1237
rect -520 1236 -519 1237
rect -492 1236 -491 1237
rect -441 1236 -440 1237
rect -413 1236 -412 1237
rect 207 1236 208 1237
rect 235 1236 236 1237
rect 286 1236 287 1237
rect 314 1236 315 1237
rect 365 1236 366 1237
rect 393 1236 394 1237
rect 444 1236 445 1237
rect 472 1236 473 1237
rect -678 1187 -649 1202
rect -599 1187 -570 1202
rect -520 1187 -491 1202
rect -441 1187 -412 1202
rect -195 1191 -166 1209
rect -39 1191 -10 1209
rect 207 1187 236 1202
rect 286 1187 315 1202
rect 365 1187 394 1202
rect 444 1187 473 1202
rect -678 1153 -649 1169
rect -599 1153 -570 1169
rect -520 1153 -491 1169
rect -441 1153 -412 1169
rect -195 1150 -166 1168
rect -39 1150 -10 1168
rect 207 1153 236 1169
rect 286 1153 315 1169
rect 365 1153 394 1169
rect 444 1153 473 1169
rect -678 1119 -677 1120
rect -650 1119 -649 1120
rect -599 1119 -598 1120
rect -571 1119 -570 1120
rect -520 1119 -519 1120
rect -492 1119 -491 1120
rect -441 1119 -440 1120
rect -413 1119 -412 1120
rect 207 1119 208 1120
rect 235 1119 236 1120
rect 286 1119 287 1120
rect 314 1119 315 1120
rect 365 1119 366 1120
rect 393 1119 394 1120
rect 444 1119 445 1120
rect 472 1119 473 1120
rect -767 1093 -754 1098
rect -753 1093 -740 1097
rect -767 1090 -740 1093
rect -728 1090 -711 1119
rect -679 1118 -648 1119
rect -600 1118 -569 1119
rect -521 1118 -490 1119
rect -442 1118 -411 1119
rect -678 1111 -649 1118
rect -599 1111 -570 1118
rect -520 1111 -491 1118
rect -441 1111 -412 1118
rect -678 1097 -669 1111
rect -422 1097 -412 1111
rect -678 1091 -649 1097
rect -599 1091 -570 1097
rect -520 1091 -491 1097
rect -441 1091 -412 1097
rect -679 1090 -648 1091
rect -600 1090 -569 1091
rect -521 1090 -490 1091
rect -442 1090 -411 1091
rect -380 1090 -362 1119
rect -195 1118 -194 1119
rect -167 1118 -166 1119
rect -39 1118 -38 1119
rect -11 1118 -10 1119
rect -678 1089 -677 1090
rect -650 1089 -649 1090
rect -599 1089 -598 1090
rect -571 1089 -570 1090
rect -520 1089 -519 1090
rect -492 1089 -491 1090
rect -441 1089 -440 1090
rect -413 1089 -412 1090
rect -245 1089 -227 1118
rect -196 1117 -165 1118
rect -195 1108 -166 1117
rect -195 1099 -185 1108
rect -176 1099 -166 1108
rect -195 1090 -166 1099
rect -196 1089 -165 1090
rect -134 1089 -116 1118
rect -89 1089 -71 1118
rect -40 1117 -9 1118
rect -39 1108 -10 1117
rect -39 1099 -29 1108
rect -20 1099 -10 1108
rect -39 1090 -10 1099
rect -40 1089 -9 1090
rect 22 1089 40 1118
rect 157 1090 175 1119
rect 206 1118 237 1119
rect 285 1118 316 1119
rect 364 1118 395 1119
rect 443 1118 474 1119
rect 207 1111 236 1118
rect 286 1111 315 1118
rect 365 1111 394 1118
rect 444 1111 473 1118
rect 207 1097 217 1111
rect 464 1097 473 1111
rect 207 1091 236 1097
rect 286 1091 315 1097
rect 365 1091 394 1097
rect 444 1091 473 1097
rect 206 1090 237 1091
rect 285 1090 316 1091
rect 364 1090 395 1091
rect 443 1090 474 1091
rect 506 1090 523 1119
rect 535 1093 548 1097
rect 549 1093 562 1098
rect 535 1090 562 1093
rect 207 1089 208 1090
rect 235 1089 236 1090
rect 286 1089 287 1090
rect 314 1089 315 1090
rect 365 1089 366 1090
rect 393 1089 394 1090
rect 444 1089 445 1090
rect 472 1089 473 1090
rect -195 1088 -194 1089
rect -167 1088 -166 1089
rect -39 1088 -38 1089
rect -11 1088 -10 1089
rect -678 1040 -649 1055
rect -599 1040 -570 1055
rect -520 1040 -491 1055
rect -441 1040 -412 1055
rect -195 1039 -166 1057
rect -39 1039 -10 1057
rect 207 1040 236 1055
rect 286 1040 315 1055
rect 365 1040 394 1055
rect 444 1040 473 1055
rect -678 1006 -649 1022
rect -599 1006 -570 1022
rect -520 1006 -491 1022
rect -441 1006 -412 1022
rect -195 1005 -166 1023
rect -39 1005 -10 1023
rect 207 1006 236 1022
rect 286 1006 315 1022
rect 365 1006 394 1022
rect 444 1006 473 1022
rect -195 973 -194 974
rect -167 973 -166 974
rect -39 973 -38 974
rect -11 973 -10 974
rect -678 972 -677 973
rect -650 972 -649 973
rect -599 972 -598 973
rect -571 972 -570 973
rect -520 972 -519 973
rect -492 972 -491 973
rect -441 972 -440 973
rect -413 972 -412 973
rect -728 943 -711 972
rect -679 971 -648 972
rect -600 971 -569 972
rect -521 971 -490 972
rect -442 971 -411 972
rect -678 964 -649 971
rect -599 964 -570 971
rect -520 964 -491 971
rect -441 964 -412 971
rect -678 950 -669 964
rect -422 950 -412 964
rect -678 944 -649 950
rect -599 944 -570 950
rect -520 944 -491 950
rect -441 944 -412 950
rect -679 943 -648 944
rect -600 943 -569 944
rect -521 943 -490 944
rect -442 943 -411 944
rect -380 943 -362 972
rect -245 944 -227 973
rect -196 972 -165 973
rect -195 963 -166 972
rect -195 954 -185 963
rect -176 954 -166 963
rect -195 945 -166 954
rect -196 944 -165 945
rect -134 944 -116 973
rect -89 944 -71 973
rect -40 972 -9 973
rect -39 963 -10 972
rect -39 954 -29 963
rect -20 954 -10 963
rect -39 945 -10 954
rect -40 944 -9 945
rect 22 944 40 973
rect 207 972 208 973
rect 235 972 236 973
rect 286 972 287 973
rect 314 972 315 973
rect 365 972 366 973
rect 393 972 394 973
rect 444 972 445 973
rect 472 972 473 973
rect -195 943 -194 944
rect -167 943 -166 944
rect -39 943 -38 944
rect -11 943 -10 944
rect 157 943 175 972
rect 206 971 237 972
rect 285 971 316 972
rect 364 971 395 972
rect 443 971 474 972
rect 207 964 236 971
rect 286 964 315 971
rect 365 964 394 971
rect 444 964 473 971
rect 207 950 217 964
rect 464 950 473 964
rect 207 944 236 950
rect 286 944 315 950
rect 365 944 394 950
rect 444 944 473 950
rect 206 943 237 944
rect 285 943 316 944
rect 364 943 395 944
rect 443 943 474 944
rect 506 943 523 972
rect -678 942 -677 943
rect -650 942 -649 943
rect -599 942 -598 943
rect -571 942 -570 943
rect -520 942 -519 943
rect -492 942 -491 943
rect -441 942 -440 943
rect -413 942 -412 943
rect 207 942 208 943
rect 235 942 236 943
rect 286 942 287 943
rect 314 942 315 943
rect 365 942 366 943
rect 393 942 394 943
rect 444 942 445 943
rect 472 942 473 943
rect -678 893 -649 908
rect -599 893 -570 908
rect -520 893 -491 908
rect -441 893 -412 908
rect -195 894 -166 912
rect -39 894 -10 912
rect 207 893 236 908
rect 286 893 315 908
rect 365 893 394 908
rect 444 893 473 908
rect -678 859 -649 875
rect -599 859 -570 875
rect -520 859 -491 875
rect -441 859 -412 875
rect -195 851 -166 869
rect -39 851 -10 869
rect 207 859 236 875
rect 286 859 315 875
rect 365 859 394 875
rect 444 859 473 875
rect -678 825 -677 826
rect -650 825 -649 826
rect -599 825 -598 826
rect -571 825 -570 826
rect -520 825 -519 826
rect -492 825 -491 826
rect -441 825 -440 826
rect -413 825 -412 826
rect 207 825 208 826
rect 235 825 236 826
rect 286 825 287 826
rect 314 825 315 826
rect 365 825 366 826
rect 393 825 394 826
rect 444 825 445 826
rect 472 825 473 826
rect -728 796 -711 825
rect -679 824 -648 825
rect -600 824 -569 825
rect -521 824 -490 825
rect -442 824 -411 825
rect -678 817 -649 824
rect -599 817 -570 824
rect -520 817 -491 824
rect -441 817 -412 824
rect -678 803 -669 817
rect -422 803 -412 817
rect -678 797 -649 803
rect -599 797 -570 803
rect -520 797 -491 803
rect -441 797 -412 803
rect -679 796 -648 797
rect -600 796 -569 797
rect -521 796 -490 797
rect -442 796 -411 797
rect -380 796 -362 825
rect -195 819 -194 820
rect -167 819 -166 820
rect -39 819 -38 820
rect -11 819 -10 820
rect -678 795 -677 796
rect -650 795 -649 796
rect -599 795 -598 796
rect -571 795 -570 796
rect -520 795 -519 796
rect -492 795 -491 796
rect -441 795 -440 796
rect -413 795 -412 796
rect -245 790 -227 819
rect -196 818 -165 819
rect -195 809 -166 818
rect -195 800 -185 809
rect -176 800 -166 809
rect -195 791 -166 800
rect -196 790 -165 791
rect -134 790 -116 819
rect -89 790 -71 819
rect -40 818 -9 819
rect -39 809 -10 818
rect -39 800 -29 809
rect -20 800 -10 809
rect -39 791 -10 800
rect -40 790 -9 791
rect 22 790 40 819
rect 157 796 175 825
rect 206 824 237 825
rect 285 824 316 825
rect 364 824 395 825
rect 443 824 474 825
rect 207 817 236 824
rect 286 817 315 824
rect 365 817 394 824
rect 444 817 473 824
rect 207 803 217 817
rect 464 803 473 817
rect 207 797 236 803
rect 286 797 315 803
rect 365 797 394 803
rect 444 797 473 803
rect 206 796 237 797
rect 285 796 316 797
rect 364 796 395 797
rect 443 796 474 797
rect 506 796 523 825
rect 207 795 208 796
rect 235 795 236 796
rect 286 795 287 796
rect 314 795 315 796
rect 365 795 366 796
rect 393 795 394 796
rect 444 795 445 796
rect 472 795 473 796
rect -195 789 -194 790
rect -167 789 -166 790
rect -39 789 -38 790
rect -11 789 -10 790
rect -678 746 -649 761
rect -599 746 -570 761
rect -520 746 -491 761
rect -441 746 -412 761
rect -195 740 -166 758
rect -39 740 -10 758
rect 207 746 236 761
rect 286 746 315 761
rect 365 746 394 761
rect 444 746 473 761
use swc4x1cellOverlap2  swc4x1cellOverlap2_1
timestamp 1607392100
transform -1 0 -257 0 1 1110
box -191 -382 744 223
use swc4x1cellOverlap2  swc4x1cellOverlap2_0
timestamp 1607392100
transform 1 0 52 0 1 1110
box -191 -382 744 223
<< end >>
