magic
tech sky130A
timestamp 1628704256
<< checkpaint >>
rect -630 1229 2255 1640
rect -630 -610 2422 1229
rect -630 -630 2255 -610
<< error_s >>
rect 58 537 64 543
rect 111 537 117 543
rect 52 487 58 493
rect 117 487 123 493
rect 481 478 487 484
rect 586 478 592 484
rect 475 428 481 434
rect 592 428 598 434
rect 481 177 487 183
rect 586 177 592 183
rect 58 123 64 129
rect 111 123 117 129
rect 475 127 481 133
rect 592 127 598 133
rect 52 73 58 79
rect 117 73 123 79
<< nwell >>
rect 1665 592 1792 610
rect 1145 436 1311 458
rect 1191 275 1219 299
rect 1664 5 1792 24
<< locali >>
rect 283 344 329 353
rect 283 327 286 344
rect 303 327 329 344
rect 283 275 329 327
rect 283 258 286 275
rect 303 258 329 275
rect 283 252 329 258
<< viali >>
rect 286 327 303 344
rect 286 258 303 275
<< metal1 >>
rect 35 603 77 610
rect 405 602 428 610
rect 1057 602 1076 610
rect 1101 602 1129 610
rect 1596 596 1630 610
rect 1663 595 1690 610
rect 279 349 317 353
rect 279 256 283 349
rect 312 256 317 349
rect 279 252 317 256
rect 1596 5 1630 24
rect 1663 5 1690 26
<< via1 >>
rect 1600 444 1626 470
rect 283 344 312 349
rect 283 327 286 344
rect 286 327 303 344
rect 303 327 312 344
rect 283 275 312 327
rect 283 258 286 275
rect 286 258 303 275
rect 303 258 312 275
rect 283 256 312 258
<< metal2 >>
rect 1343 583 1368 609
rect 0 542 7 560
rect 1449 485 1474 522
rect 1596 470 1630 474
rect 1596 465 1600 470
rect 1145 436 1311 458
rect 1361 446 1600 465
rect 1361 389 1380 446
rect 1596 444 1600 446
rect 1626 444 1630 470
rect 1596 441 1630 444
rect 1452 400 1473 429
rect 282 370 1380 389
rect 282 352 301 370
rect 280 349 315 352
rect 280 256 283 349
rect 312 256 315 349
rect 1777 339 1792 361
rect 1347 316 1372 339
rect 1191 275 1219 299
rect 1777 257 1792 279
rect 280 253 315 256
rect 1296 192 1473 212
rect 1139 143 1155 183
rect 1267 111 1473 132
rect 0 57 8 72
rect 1187 7 1213 32
use sky130_hilas_FGBias2x1cell  sky130_hilas_FGBias2x1cell_0
timestamp 1628285143
transform 1 0 396 0 1 387
box -396 -387 1229 623
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_0
timestamp 1628704233
transform 1 0 989 0 1 445
box 133 -440 320 165
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1628704233
transform 1 0 1145 0 -1 170
box 133 -440 320 165
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1628285143
transform 1 0 1637 0 1 46
box -172 -26 155 553
<< labels >>
rlabel metal1 1596 5 1630 11 0 VGND
port 7 nsew ground default
rlabel metal1 1663 5 1690 11 0 VPWR
port 8 nsew power default
rlabel metal1 1596 605 1630 610 0 VGND
port 7 nsew ground default
rlabel metal1 1663 605 1690 610 0 VPWR
port 8 nsew power default
rlabel metal2 1347 316 1372 339 0 VIN21
port 3 nsew
rlabel metal2 1187 7 1210 32 0 VIN12
port 2 nsew analog default
rlabel metal2 1343 583 1368 609 0 VIN22
port 4 nsew
rlabel metal2 1777 257 1792 279 0 OUTPUT1
port 5 nsew
rlabel metal2 1777 339 1792 361 0 OUTPUT2
port 6 nsew
rlabel metal1 1057 602 1076 610 0 COLSEL1
port 1 nsew
rlabel metal2 0 542 7 560 0 DRAIN1
port 9 nsew
rlabel metal2 0 57 8 72 0 DRAIN2
port 10 nsew
rlabel metal1 35 603 77 610 0 VTUN
port 11 nsew
rlabel metal1 405 602 428 610 0 GATE1
port 12 nsew
rlabel metal1 1101 602 1129 610 0 VINJ
port 13 nsew
rlabel metal2 1191 275 1214 299 0 VIN11
port 14 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
