magic
tech sky130A
timestamp 1634057745
<< checkpaint >>
rect -630 1202 2655 2117
rect -630 -234 3322 1202
rect 605 -514 3322 -234
rect 610 -592 3322 -514
rect 610 -610 1904 -592
<< error_s >>
rect 1348 612 1398 618
rect 1420 612 1470 618
rect 1348 570 1398 576
rect 1420 570 1470 576
rect 1420 543 1470 549
rect 1420 501 1470 507
rect 1420 460 1470 466
rect 1420 418 1470 424
rect 1348 391 1398 397
rect 1420 391 1470 397
rect 1348 349 1398 355
rect 1420 349 1470 355
rect 1348 288 1398 294
rect 1420 288 1470 294
rect 1348 246 1398 252
rect 1420 246 1470 252
rect 1420 219 1470 225
rect 1420 177 1470 183
rect 1420 135 1470 141
rect 1420 93 1470 99
rect 1348 66 1398 72
rect 1420 66 1470 72
rect 1348 24 1398 30
rect 1420 24 1470 30
<< nwell >>
rect 1241 618 1537 619
rect 1241 603 1282 618
rect 1810 609 1848 619
rect 2213 605 2253 619
rect 1241 602 1300 603
rect 1241 426 1282 602
rect 1230 384 1282 426
rect 1230 364 1281 384
rect 1230 311 1282 364
rect 1241 15 1282 311
<< poly >>
rect 2551 573 2571 619
rect 2551 14 2571 39
<< locali >>
rect 1227 32 1245 124
<< metal1 >>
rect 1317 612 1333 619
rect 1358 612 1377 619
rect 1398 612 1414 619
rect 1810 609 1848 619
rect 2213 591 2253 619
rect 2473 573 2496 619
rect 2599 573 2622 619
rect 1560 487 1581 561
rect 1230 311 1251 426
rect 1558 150 1574 300
rect 2599 184 2622 189
rect 2595 183 2623 184
rect 2595 181 2625 183
rect 2595 154 2596 181
rect 2623 154 2625 181
rect 2595 151 2625 154
rect 1810 14 1848 24
rect 2473 14 2496 39
rect 2599 14 2622 39
<< via1 >>
rect 2596 154 2623 181
<< metal2 >>
rect 1226 572 1299 590
rect 1584 569 2349 588
rect 1584 567 2366 569
rect 2328 548 2366 567
rect 2277 547 2291 548
rect 1230 484 1245 526
rect 2277 514 2292 547
rect 2277 494 2398 514
rect 1230 475 1557 484
rect 2512 483 2638 499
rect 1230 469 1573 475
rect 1543 459 1573 469
rect 1228 409 1260 436
rect 2288 428 2408 438
rect 2287 420 2408 428
rect 2380 408 2408 420
rect 2380 406 2383 408
rect 1223 377 1281 395
rect 2512 390 2638 406
rect 1551 361 1574 362
rect 1551 358 2308 361
rect 1551 341 2314 358
rect 1551 331 1575 341
rect 1230 313 1575 331
rect 2295 321 2366 341
rect 1230 311 1567 313
rect 1565 291 2310 293
rect 1565 271 2366 291
rect 1565 270 1597 271
rect 1226 248 1281 266
rect 1224 175 1244 225
rect 2286 209 2386 225
rect 2512 206 2638 222
rect 2593 181 2626 182
rect 1224 155 1579 175
rect 2593 173 2596 181
rect 1958 156 2596 173
rect 2593 154 2596 156
rect 2623 154 2626 181
rect 2593 153 2626 154
rect 1223 104 1251 131
rect 2287 111 2387 128
rect 2514 113 2638 129
rect 2287 110 2381 111
rect 1224 52 1281 70
rect 2310 65 2365 66
rect 1552 43 2365 65
rect 1552 42 2311 43
rect 1552 41 1629 42
rect 1228 24 1262 37
rect 1552 24 1576 41
rect 1228 16 1576 24
rect 1239 0 1576 16
use sky130_hilas_WTA4stage01  sky130_hilas_WTA4stage01_0
timestamp 1634057715
transform 1 0 2409 0 1 38
box 0 0 283 534
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1634057699
transform 1 0 1235 0 1 116
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1634057699
transform 1 0 1240 0 1 20
box 0 0 34 33
use sky130_hilas_m12m2  sky130_hilas_m12m2_4
timestamp 1634057711
transform 1 0 1564 0 1 278
box 0 0 32 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_2
timestamp 1634057711
transform 1 0 1564 0 1 466
box 0 0 32 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1634057711
transform 1 0 1566 0 1 571
box 0 0 32 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_3
timestamp 1634057711
transform 1 0 1237 0 1 416
box 0 0 32 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1634057711
transform 1 0 1235 0 1 315
box 0 0 32 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_5
timestamp 1634057711
transform 1 0 1551 0 1 160
box 0 0 32 32
use sky130_hilas_swc4x1BiasCell  sky130_hilas_swc4x1BiasCell_0
timestamp 1634057716
transform -1 0 2025 0 1 396
box 0 0 2025 1091
<< labels >>
rlabel metal2 2631 483 2638 499 0 OUTPUT1
port 4 nsew analog default
rlabel metal2 2633 390 2638 406 0 OUTPUT2
port 5 nsew analog default
rlabel metal2 2633 206 2638 222 0 OUTPUT3
port 6 nsew analog default
rlabel metal2 2633 113 2638 129 0 OUTPUT4
port 7 nsew analog default
rlabel metal1 2599 613 2622 619 0 VGND
port 1 nsew ground default
rlabel metal1 2599 14 2622 20 0 VGND
port 1 nsew ground default
rlabel metal2 1230 506 1245 526 0 INPUT1
port 8 nsew analog default
rlabel metal2 1230 409 1256 435 0 INPUT2
port 9 nsew analog default
rlabel metal2 1224 208 1244 225 0 INPUT3
port 10 nsew analog default
rlabel metal2 1223 104 1251 131 0 INPUT4
port 11 nsew analog default
rlabel metal1 1811 609 1847 619 0 GATE1
port 16 nsew
rlabel metal1 2213 605 2253 619 0 VTUN
port 17 nsew
rlabel metal1 2473 14 2496 20 0 WTAMIDDLENODE
port 18 nsew
rlabel metal1 2473 613 2496 619 0 WTAMIDDLENODE
port 18 nsew
rlabel metal1 1358 612 1377 619 0 COLSEL1
port 19 nsew
rlabel metal1 1317 612 1333 619 0 VINJ
port 21 nsew
rlabel metal1 1398 612 1414 619 0 VPWR
port 20 nsew
rlabel metal2 1226 572 1235 590 0 DRAIN1
port 12 nsew
rlabel metal2 1223 377 1232 395 0 DRAIN2
port 22 nsew
rlabel metal2 1226 248 1235 266 0 DRAIN3
port 23 nsew
rlabel metal2 1224 52 1233 70 0 DRAIN4
port 24 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
