magic
tech sky130A
timestamp 1632255311
<< error_s >>
rect 76 55 116 61
rect 135 49 151 54
rect 45 31 53 39
rect 53 23 61 26
rect 76 13 116 19
<< nwell >>
rect 49 84 163 143
rect 0 0 163 84
<< pmos >>
rect 76 19 116 55
<< pdiff >>
rect 47 48 76 55
rect 47 31 53 48
rect 70 31 76 48
rect 47 19 76 31
rect 116 48 145 55
rect 116 31 122 48
rect 139 31 145 48
rect 116 19 145 31
<< pdiffc >>
rect 53 31 70 48
rect 122 31 139 48
<< poly >>
rect 76 55 116 78
rect 76 6 116 19
<< locali >>
rect 49 93 163 111
rect 53 48 70 56
rect 114 31 122 48
rect 139 31 152 49
rect 53 26 70 31
<< metal1 >>
rect 141 55 160 114
rect 139 26 162 55
<< metal2 >>
rect 126 109 163 129
rect 0 31 22 32
rect 0 11 163 31
rect 0 10 22 11
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1632251356
transform 1 0 53 0 1 26
box 0 0 34 33
use sky130_hilas_li2m1  sky130_hilas_li2m1_3
timestamp 1632251332
transform 1 0 149 0 1 34
box 0 0 23 29
use sky130_hilas_m12m2  sky130_hilas_m12m2_2
timestamp 1632251372
transform 1 0 140 0 1 112
box 0 0 32 32
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
