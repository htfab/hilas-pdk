VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_cellattempt01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_cellattempt01 ;
  ORIGIN 2.640 3.820 ;
  SIZE 10.080 BY 6.050 ;
  OBS
      LAYER nwell ;
        RECT 6.320 -0.720 6.670 -0.710 ;
        RECT 6.320 -0.880 6.490 -0.720 ;
        RECT 6.660 -0.880 6.670 -0.720 ;
      LAYER li1 ;
        RECT 6.230 -0.880 6.670 -0.710 ;
      LAYER mcon ;
        RECT 6.490 -0.880 6.670 -0.710 ;
      LAYER met1 ;
        RECT -2.280 -3.820 -1.880 2.170 ;
        RECT 6.540 -0.680 6.670 -0.660 ;
        RECT 6.460 -0.910 6.700 -0.680 ;
        RECT 6.560 -0.950 6.670 -0.910 ;
      LAYER met2 ;
        RECT -2.640 1.660 4.970 1.730 ;
        RECT -2.640 1.550 5.000 1.660 ;
        RECT -2.640 1.120 7.100 1.300 ;
        RECT -2.640 0.240 4.970 0.300 ;
        RECT -2.640 0.120 5.000 0.240 ;
        RECT -2.640 -0.200 4.960 -0.130 ;
        RECT -2.640 -0.310 5.000 -0.200 ;
        RECT -2.620 -1.460 5.000 -1.290 ;
        RECT -2.620 -1.880 5.000 -1.710 ;
        RECT -2.620 -2.860 5.000 -2.690 ;
        RECT -1.840 -2.950 -0.300 -2.860 ;
        RECT -2.620 -3.300 5.000 -3.130 ;
  END
END sky130_hilas_cellattempt01
END LIBRARY

