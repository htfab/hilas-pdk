magic
tech sky130A
timestamp 1634057782
<< error_p >>
rect 2 28 65 29
<< mvndiff >>
rect 2 22 65 28
rect 2 5 8 22
rect 25 5 42 22
rect 59 5 65 22
rect 2 0 65 5
<< mvndiffc >>
rect 8 5 25 22
rect 42 5 59 22
<< locali >>
rect 0 5 8 22
rect 59 5 67 22
<< viali >>
rect 25 5 42 22
<< metal1 >>
rect 14 22 53 25
rect 14 5 25 22
rect 42 5 53 22
rect 14 2 53 5
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
