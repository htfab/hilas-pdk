magic
tech sky130A
timestamp 1627062638
<< metal1 >>
rect 34 619 63 624
rect 475 617 506 624
rect 776 619 800 624
rect 34 0 63 5
rect 475 0 506 6
rect 776 0 800 5
<< metal2 >>
rect 0 572 11 592
rect 871 474 880 506
rect 0 417 11 437
rect 871 319 880 351
rect 0 262 11 282
rect 871 164 880 196
rect 0 107 11 127
rect 871 9 880 41
use sky130_hilas_StepUpDigital  StepUpDigital_3
timestamp 1624113415
transform 1 0 -19 0 1 40
box 19 -40 899 119
use sky130_hilas_StepUpDigital  StepUpDigital_0
timestamp 1624113415
transform 1 0 -19 0 1 195
box 19 -40 899 119
use sky130_hilas_StepUpDigital  StepUpDigital_1
timestamp 1624113415
transform 1 0 -19 0 1 350
box 19 -40 899 119
use sky130_hilas_StepUpDigital  StepUpDigital_2
timestamp 1624113415
transform 1 0 -19 0 1 505
box 19 -40 899 119
<< labels >>
rlabel metal2 871 474 880 506 0 INPUT1
port 1 nsew
rlabel metal2 871 319 880 351 0 INPUT2
port 2 nsew
rlabel metal2 871 164 880 196 0 INPUT3
port 3 nsew
rlabel metal2 871 9 880 41 0 INPUT4
port 4 nsew
rlabel metal1 776 619 800 624 0 VPWR
port 5 nsew
rlabel metal1 776 0 800 5 0 VPWR
port 5 nsew
rlabel metal1 34 619 63 624 0 VINJ
port 6 nsew
rlabel metal1 34 0 63 5 0 VINJ
port 6 nsew
rlabel metal2 0 572 11 592 0 OUTPUT1
port 7 nsew
rlabel metal2 0 417 11 437 0 OUTPUT2
port 8 nsew
rlabel metal2 0 262 11 282 0 OUTPUT3
port 9 nsew
rlabel metal2 0 107 11 127 0 OUTPUT4
port 10 nsew
rlabel metal1 475 617 506 624 0 VGND
port 11 nsew
rlabel metal1 475 0 506 6 0 VGND
port 11 nsew
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
