magic
tech sky130A
timestamp 1628698502
<< checkpaint >>
rect -1156 1364 622 1375
rect -1156 -475 949 1364
rect -1156 -490 622 -475
<< error_s >>
rect 214 528 215 529
<< nwell >>
rect -569 744 -378 745
rect -569 184 -9 744
rect 191 727 319 745
rect -569 166 -526 184
rect -569 143 -498 166
rect -569 141 -526 143
rect 191 140 319 159
<< nsubdiff >>
rect -550 661 -519 698
rect -550 644 -544 661
rect -527 644 -519 661
rect -550 627 -519 644
rect -550 610 -544 627
rect -527 610 -519 627
rect -550 593 -519 610
rect -550 576 -544 593
rect -527 576 -519 593
rect -550 559 -519 576
rect -550 542 -544 559
rect -527 542 -519 559
rect -550 525 -519 542
rect -550 508 -544 525
rect -527 508 -519 525
rect -550 493 -519 508
rect -551 358 -519 391
rect -551 341 -543 358
rect -526 341 -519 358
rect -551 324 -519 341
rect -551 307 -543 324
rect -526 307 -519 324
rect -551 290 -519 307
rect -551 273 -543 290
rect -526 273 -519 290
rect -551 256 -519 273
rect -551 239 -543 256
rect -526 239 -519 256
rect -551 222 -519 239
rect -551 205 -543 222
rect -526 205 -519 222
rect -551 190 -519 205
<< nsubdiffcont >>
rect -544 644 -527 661
rect -544 610 -527 627
rect -544 576 -527 593
rect -544 542 -527 559
rect -544 508 -527 525
rect -543 341 -526 358
rect -543 307 -526 324
rect -543 273 -526 290
rect -543 239 -526 256
rect -543 205 -526 222
<< locali >>
rect -502 697 -468 698
rect -527 673 -468 697
rect -527 624 -485 673
rect 196 598 198 615
rect 215 598 221 615
rect 196 561 221 598
rect 196 545 217 561
rect 196 528 198 545
rect 215 528 217 545
rect 196 526 217 528
rect -544 491 -527 508
rect -543 197 -526 205
<< viali >>
rect -544 661 -527 678
rect -544 627 -527 644
rect -485 656 -468 673
rect -485 622 -468 639
rect -544 593 -527 610
rect -544 559 -527 576
rect -544 525 -527 542
rect 198 598 215 615
rect 198 528 215 545
rect -543 358 -526 375
rect -543 324 -526 341
rect -543 290 -526 307
rect -543 256 -526 273
rect -543 222 -526 239
<< metal1 >>
rect 123 731 157 745
rect 190 730 217 745
rect -547 698 -494 699
rect -547 697 -468 698
rect -547 691 -465 697
rect -547 678 -535 691
rect -547 661 -544 678
rect -476 673 -465 691
rect -547 644 -535 661
rect -468 667 -465 673
rect -468 656 -462 667
rect -547 627 -544 644
rect -476 639 -462 656
rect -547 619 -535 627
rect -468 638 -462 639
rect -468 622 -465 638
rect -476 619 -465 622
rect -547 613 -465 619
rect 193 615 225 619
rect -547 610 -483 613
rect -547 593 -544 610
rect -527 593 -483 610
rect -547 576 -483 593
rect -547 559 -544 576
rect -527 559 -483 576
rect -547 542 -483 559
rect -547 525 -544 542
rect -527 525 -483 542
rect 193 529 194 615
rect 220 529 225 615
rect 193 528 198 529
rect 215 528 225 529
rect 193 527 225 528
rect 196 526 225 527
rect -547 375 -483 525
rect -547 358 -543 375
rect -526 358 -483 375
rect -547 341 -483 358
rect -547 324 -543 341
rect -526 324 -483 341
rect -547 307 -483 324
rect -547 290 -543 307
rect -526 290 -483 307
rect -547 273 -483 290
rect -547 256 -543 273
rect -526 256 -483 273
rect -547 239 -483 256
rect -547 222 -543 239
rect -526 222 -483 239
rect -547 195 -483 222
rect -525 194 -483 195
rect 123 140 157 159
rect 190 140 217 161
<< via1 >>
rect -535 678 -476 691
rect -535 661 -527 678
rect -527 673 -476 678
rect -527 661 -485 673
rect -535 656 -485 661
rect -485 656 -476 673
rect -535 644 -476 656
rect -535 627 -527 644
rect -527 639 -476 644
rect -527 627 -485 639
rect -535 622 -485 627
rect -485 622 -476 639
rect -535 619 -476 622
rect 194 598 198 615
rect 198 598 215 615
rect 215 598 220 615
rect 194 545 220 598
rect 194 529 198 545
rect 198 529 215 545
rect 215 529 220 545
<< metal2 >>
rect -490 698 -466 745
rect -130 718 -105 744
rect -542 691 -466 698
rect -542 619 -535 691
rect -476 663 -466 691
rect -476 640 -88 663
rect -476 619 -466 640
rect -542 616 -466 619
rect -542 615 -497 616
rect -111 604 -88 640
rect -24 620 1 657
rect 191 615 224 619
rect 191 604 194 615
rect -381 571 -162 593
rect -111 584 194 604
rect -85 583 194 584
rect -21 535 0 564
rect 191 529 194 583
rect 220 529 224 615
rect 191 526 224 529
rect 304 474 319 496
rect -126 451 -101 474
rect -568 410 -422 434
rect -282 410 -254 434
rect -568 409 -504 410
rect 304 392 319 414
rect -177 327 0 347
rect -334 292 -318 310
rect -336 291 -318 292
rect -358 278 -318 291
rect -358 229 -322 278
rect -206 246 0 267
rect -564 143 -399 166
rect -286 142 -260 167
<< rmetal2 >>
rect -497 615 -466 616
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1628698494
transform 1 0 164 0 1 181
box -172 -26 155 553
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628698494
transform 1 0 -480 0 1 709
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628698494
transform 1 0 -396 0 1 581
box -14 -15 20 18
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_2
timestamp 1628698494
transform 1 0 -659 0 1 580
box 133 -440 320 165
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1628698494
transform 1 0 -328 0 -1 305
box 133 -440 320 165
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_0
timestamp 1628698494
transform 1 0 -484 0 1 580
box 133 -440 320 165
<< labels >>
rlabel metal1 123 140 157 146 0 VGND
port 3 nsew ground default
rlabel metal1 190 140 217 146 0 VPWR
port 4 nsew power default
rlabel metal1 123 740 157 745 0 VGND
port 3 nsew ground default
rlabel metal1 190 740 217 745 0 VPWR
port 4 nsew power default
rlabel metal2 -282 410 -259 434 0 VIN11
port 7 nsew analog default
rlabel metal2 -126 451 -101 474 0 VIN21
port 6 nsew analog default
rlabel metal2 -286 142 -263 167 0 VIN12
port 8 nsew analog default
rlabel metal2 -130 718 -105 744 0 VIN22
port 5 nsew analog default
rlabel metal2 304 392 319 414 0 VOUT_AMP1
port 2 nsew analog default
rlabel metal2 304 474 319 496 0 VOUT_AMP2
port 1 nsew analog default
rlabel metal2 -490 737 -466 745 0 VPWR
port 4 nsew power default
rlabel metal2 -526 410 -519 434 0 VBIAS1
port 10 nsew analog default
rlabel metal2 -526 143 -519 166 0 VBIAS2
port 9 nsew analog default
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
