VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_li2m1
  CLASS BLOCK ;
  FOREIGN /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_li2m1 ;
  ORIGIN 0.100 0.080 ;
  SIZE 0.230 BY 0.290 ;
  OBS
      LAYER li1 ;
        RECT -0.080 -0.050 0.110 0.180 ;
      LAYER met1 ;
        RECT -0.100 -0.080 0.130 0.210 ;
  END
END /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_li2m1
END LIBRARY

