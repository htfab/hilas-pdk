magic
tech sky130A
timestamp 1634057846
<< nwell >>
rect 1617 470 1845 633
rect 1617 218 1787 470
rect 1616 16 1787 218
<< nmos >>
rect 547 352 562 615
rect 547 21 562 284
rect 649 19 669 615
rect 702 19 722 615
rect 753 19 773 615
rect 804 19 824 615
rect 855 19 875 615
rect 906 19 926 615
rect 957 19 977 615
rect 1008 19 1028 615
rect 1059 19 1079 615
rect 1110 19 1130 615
rect 1161 19 1181 615
rect 1212 19 1232 615
rect 1263 19 1283 615
rect 1314 19 1334 615
rect 1365 19 1385 615
rect 1416 19 1436 615
rect 1525 415 1545 615
<< pmos >>
rect 1667 34 1687 615
rect 1719 34 1739 615
<< ndiff >>
rect 519 603 547 615
rect 519 360 523 603
rect 540 360 547 603
rect 519 352 547 360
rect 562 601 590 615
rect 562 358 568 601
rect 585 358 590 601
rect 562 352 590 358
rect 570 284 590 352
rect 518 273 547 284
rect 518 28 523 273
rect 540 28 547 273
rect 518 21 547 28
rect 562 272 590 284
rect 562 27 568 272
rect 585 27 590 272
rect 562 21 590 27
rect 620 607 649 615
rect 620 23 626 607
rect 643 23 649 607
rect 620 19 649 23
rect 669 607 702 615
rect 669 23 677 607
rect 694 23 702 607
rect 669 19 702 23
rect 722 607 753 615
rect 722 23 728 607
rect 745 23 753 607
rect 722 19 753 23
rect 773 607 804 615
rect 773 23 780 607
rect 797 23 804 607
rect 773 19 804 23
rect 824 607 855 615
rect 824 23 830 607
rect 847 23 855 607
rect 824 19 855 23
rect 875 607 906 615
rect 875 23 881 607
rect 898 23 906 607
rect 875 19 906 23
rect 926 607 957 615
rect 926 23 933 607
rect 950 23 957 607
rect 926 19 957 23
rect 977 607 1008 615
rect 977 23 984 607
rect 1001 23 1008 607
rect 977 19 1008 23
rect 1028 607 1059 615
rect 1028 23 1035 607
rect 1052 23 1059 607
rect 1028 19 1059 23
rect 1079 607 1110 615
rect 1079 23 1086 607
rect 1103 23 1110 607
rect 1079 19 1110 23
rect 1130 607 1161 615
rect 1130 23 1137 607
rect 1154 23 1161 607
rect 1130 19 1161 23
rect 1181 607 1212 615
rect 1181 23 1187 607
rect 1204 23 1212 607
rect 1181 19 1212 23
rect 1232 607 1263 615
rect 1232 23 1239 607
rect 1256 23 1263 607
rect 1232 19 1263 23
rect 1283 607 1314 615
rect 1283 23 1289 607
rect 1306 23 1314 607
rect 1283 19 1314 23
rect 1334 607 1365 615
rect 1334 23 1340 607
rect 1357 23 1365 607
rect 1334 19 1365 23
rect 1385 607 1416 615
rect 1385 23 1392 607
rect 1409 23 1416 607
rect 1385 19 1416 23
rect 1436 607 1467 615
rect 1436 23 1442 607
rect 1459 23 1467 607
rect 1494 606 1525 615
rect 1494 423 1501 606
rect 1518 423 1525 606
rect 1494 415 1525 423
rect 1545 606 1576 615
rect 1545 423 1552 606
rect 1569 423 1576 606
rect 1545 415 1576 423
rect 1436 19 1467 23
<< pdiff >>
rect 1637 594 1667 615
rect 1637 44 1644 594
rect 1661 44 1667 594
rect 1637 34 1667 44
rect 1687 594 1719 615
rect 1687 45 1694 594
rect 1711 45 1719 594
rect 1687 34 1719 45
rect 1739 593 1768 615
rect 1739 45 1745 593
rect 1762 45 1768 593
rect 1739 34 1768 45
<< ndiffc >>
rect 523 360 540 603
rect 568 358 585 601
rect 523 28 540 273
rect 568 27 585 272
rect 626 23 643 607
rect 677 23 694 607
rect 728 23 745 607
rect 780 23 797 607
rect 830 23 847 607
rect 881 23 898 607
rect 933 23 950 607
rect 984 23 1001 607
rect 1035 23 1052 607
rect 1086 23 1103 607
rect 1137 23 1154 607
rect 1187 23 1204 607
rect 1239 23 1256 607
rect 1289 23 1306 607
rect 1340 23 1357 607
rect 1392 23 1409 607
rect 1442 23 1459 607
rect 1501 423 1518 606
rect 1552 423 1569 606
<< pdiffc >>
rect 1644 44 1661 594
rect 1694 45 1711 594
rect 1745 45 1762 593
<< psubdiff >>
rect 1495 375 1571 387
rect 1495 30 1506 375
rect 1562 30 1571 375
rect 1495 18 1571 30
<< nsubdiff >>
rect 1795 594 1827 614
rect 1795 514 1802 594
rect 1819 514 1827 594
rect 1795 501 1827 514
<< psubdiffcont >>
rect 1506 30 1562 375
<< nsubdiffcont >>
rect 1802 514 1819 594
<< poly >>
rect 547 623 1617 638
rect 547 615 562 623
rect 649 615 669 623
rect 702 615 722 623
rect 753 615 773 623
rect 804 615 824 623
rect 855 615 875 623
rect 906 615 926 623
rect 957 615 977 623
rect 1008 615 1028 623
rect 1059 615 1079 623
rect 1110 615 1130 623
rect 1161 615 1181 623
rect 1212 615 1232 623
rect 1263 615 1283 623
rect 1314 615 1334 623
rect 1365 615 1385 623
rect 1416 615 1436 623
rect 1525 615 1545 623
rect 44 598 95 613
rect 44 92 59 598
rect 26 87 59 92
rect 26 70 34 87
rect 51 70 59 87
rect 26 65 59 70
rect 80 54 95 598
rect 116 598 167 613
rect 116 54 131 598
rect 80 38 131 54
rect 152 54 167 598
rect 188 598 239 613
rect 188 54 203 598
rect 152 38 203 54
rect 224 54 239 598
rect 260 598 311 613
rect 260 54 275 598
rect 224 38 275 54
rect 296 54 311 598
rect 332 598 383 613
rect 332 54 347 598
rect 296 38 347 54
rect 368 54 383 598
rect 404 598 455 613
rect 404 54 419 598
rect 368 38 419 54
rect 440 54 455 598
rect 547 339 562 352
rect 492 320 526 325
rect 492 303 500 320
rect 517 307 526 320
rect 517 303 562 307
rect 492 292 562 303
rect 547 284 562 292
rect 476 190 507 199
rect 476 173 481 190
rect 498 173 507 190
rect 476 164 507 173
rect 478 54 493 164
rect 440 38 493 54
rect 547 8 562 21
rect 1586 607 1617 623
rect 1667 615 1687 628
rect 1719 615 1739 628
rect 1586 424 1595 607
rect 1612 424 1617 607
rect 1586 416 1617 424
rect 1525 402 1545 415
rect 649 6 669 19
rect 702 6 722 19
rect 753 6 773 19
rect 804 6 824 19
rect 855 6 875 19
rect 906 6 926 19
rect 957 6 977 19
rect 1008 6 1028 19
rect 1059 6 1079 19
rect 1110 6 1130 19
rect 1161 6 1181 19
rect 1212 6 1232 19
rect 1263 6 1283 19
rect 1314 6 1334 19
rect 1365 6 1385 19
rect 1416 6 1436 19
rect 1591 269 1627 280
rect 1591 44 1596 269
rect 1613 44 1627 269
rect 1591 26 1627 44
rect 1667 26 1687 34
rect 1719 26 1739 34
rect 1591 11 1739 26
<< polycont >>
rect 34 70 51 87
rect 500 303 517 320
rect 481 173 498 190
rect 1595 424 1612 607
rect 1596 44 1613 269
<< locali >>
rect 523 603 540 611
rect 516 484 523 490
rect 516 474 522 484
rect 500 467 522 474
rect 500 448 523 467
rect 500 431 522 448
rect 500 412 523 431
rect 500 395 522 412
rect 500 380 523 395
rect 481 376 523 380
rect 481 359 484 376
rect 501 359 521 376
rect 538 359 540 360
rect 481 353 540 359
rect 568 601 585 617
rect 481 340 542 353
rect 481 337 484 340
rect 482 323 484 337
rect 501 323 522 340
rect 539 323 542 340
rect 482 322 542 323
rect 492 320 542 322
rect 492 303 500 320
rect 517 317 542 320
rect 517 303 525 317
rect 523 273 540 281
rect 481 191 498 198
rect 481 190 483 191
rect 481 165 498 173
rect 568 272 585 358
rect 24 87 60 90
rect 24 86 34 87
rect 24 69 33 86
rect 51 70 60 87
rect 50 69 60 70
rect 24 67 60 69
rect 523 20 540 28
rect 567 27 568 165
rect 624 607 645 615
rect 624 191 626 607
rect 624 174 625 191
rect 567 25 569 27
rect 567 16 585 25
rect 624 23 626 174
rect 643 23 645 607
rect 624 15 645 23
rect 675 607 696 615
rect 675 23 677 607
rect 694 89 696 607
rect 695 72 696 89
rect 694 23 696 72
rect 675 15 696 23
rect 726 607 747 615
rect 726 192 728 607
rect 726 175 727 192
rect 726 23 728 175
rect 745 23 747 607
rect 726 15 747 23
rect 778 607 799 615
rect 778 23 780 607
rect 797 89 799 607
rect 798 72 799 89
rect 797 23 799 72
rect 778 15 799 23
rect 828 607 849 615
rect 828 192 830 607
rect 828 175 829 192
rect 828 23 830 175
rect 847 23 849 607
rect 828 15 849 23
rect 879 607 900 617
rect 879 23 881 607
rect 898 89 900 607
rect 899 72 900 89
rect 898 23 900 72
rect 879 15 900 23
rect 931 607 952 617
rect 931 192 933 607
rect 931 175 932 192
rect 931 23 933 175
rect 950 23 952 607
rect 931 15 952 23
rect 982 607 1003 617
rect 982 23 984 607
rect 1001 599 1003 607
rect 1033 607 1054 617
rect 1001 89 1002 599
rect 1001 23 1002 72
rect 982 15 1002 23
rect 1033 192 1035 607
rect 1052 599 1054 607
rect 1084 607 1105 617
rect 1033 175 1034 192
rect 1033 23 1035 175
rect 1052 23 1053 599
rect 1033 15 1053 23
rect 1084 23 1086 607
rect 1103 599 1105 607
rect 1135 607 1156 617
rect 1103 89 1104 599
rect 1103 23 1104 72
rect 1084 15 1104 23
rect 1135 192 1137 607
rect 1135 175 1136 192
rect 1135 23 1137 175
rect 1154 23 1156 607
rect 1135 15 1156 23
rect 1185 607 1206 617
rect 1185 23 1187 607
rect 1204 89 1206 607
rect 1205 72 1206 89
rect 1204 23 1206 72
rect 1185 15 1206 23
rect 1237 607 1258 617
rect 1237 192 1239 607
rect 1237 175 1238 192
rect 1237 23 1239 175
rect 1256 23 1258 607
rect 1237 15 1258 23
rect 1287 607 1308 617
rect 1287 23 1289 607
rect 1306 89 1308 607
rect 1307 72 1308 89
rect 1306 23 1308 72
rect 1287 15 1308 23
rect 1338 607 1359 617
rect 1338 192 1340 607
rect 1338 175 1339 192
rect 1338 23 1340 175
rect 1357 23 1359 607
rect 1338 15 1359 23
rect 1390 607 1411 617
rect 1390 23 1392 607
rect 1409 90 1411 607
rect 1410 73 1411 90
rect 1409 23 1411 73
rect 1390 15 1411 23
rect 1440 607 1461 617
rect 1440 192 1442 607
rect 1440 175 1441 192
rect 1440 23 1442 175
rect 1459 23 1461 607
rect 1498 606 1522 617
rect 1498 423 1501 606
rect 1518 423 1522 606
rect 1498 388 1522 423
rect 1550 607 1616 616
rect 1550 606 1595 607
rect 1550 423 1552 606
rect 1569 515 1595 606
rect 1571 498 1595 515
rect 1612 514 1616 607
rect 1569 478 1595 498
rect 1614 497 1616 514
rect 1612 478 1616 497
rect 1571 461 1595 478
rect 1614 461 1616 478
rect 1569 440 1595 461
rect 1612 441 1616 461
rect 1570 424 1595 440
rect 1613 424 1616 441
rect 1570 423 1616 424
rect 1550 412 1616 423
rect 1642 594 1663 602
rect 1440 15 1461 23
rect 1496 382 1563 388
rect 1496 375 1524 382
rect 1541 375 1563 382
rect 1496 30 1506 375
rect 1562 30 1563 375
rect 1642 279 1644 594
rect 1594 269 1644 279
rect 1594 44 1596 269
rect 1613 93 1644 269
rect 1613 76 1623 93
rect 1640 76 1644 93
rect 1613 44 1644 76
rect 1661 44 1663 594
rect 1594 36 1663 44
rect 1692 594 1713 602
rect 1692 592 1694 594
rect 1692 575 1693 592
rect 1692 555 1694 575
rect 1692 538 1693 555
rect 1692 45 1694 538
rect 1711 45 1713 594
rect 1692 36 1713 45
rect 1743 593 1764 602
rect 1802 595 1819 602
rect 1743 515 1745 593
rect 1743 498 1744 515
rect 1743 478 1745 498
rect 1743 461 1744 478
rect 1743 442 1745 461
rect 1743 425 1744 442
rect 1743 45 1745 425
rect 1762 45 1764 593
rect 1818 594 1819 595
rect 1802 501 1819 514
rect 1743 36 1764 45
rect 1496 21 1563 30
<< viali >>
rect 522 467 523 484
rect 523 467 539 484
rect 522 431 523 448
rect 523 431 539 448
rect 522 395 523 412
rect 523 395 539 412
rect 484 359 501 376
rect 521 360 523 376
rect 523 360 538 376
rect 521 359 538 360
rect 484 323 501 340
rect 522 323 539 340
rect 483 190 500 191
rect 483 174 498 190
rect 498 174 500 190
rect 522 95 523 112
rect 523 95 539 112
rect 33 70 34 86
rect 34 70 50 86
rect 33 69 50 70
rect 522 58 523 75
rect 523 58 539 75
rect 625 174 626 191
rect 626 174 642 191
rect 570 97 585 114
rect 585 97 587 114
rect 569 61 585 78
rect 585 61 586 78
rect 569 27 585 42
rect 585 27 586 42
rect 569 25 586 27
rect 678 72 694 89
rect 694 72 695 89
rect 727 175 728 192
rect 728 175 744 192
rect 781 72 797 89
rect 797 72 798 89
rect 829 175 830 192
rect 830 175 846 192
rect 882 72 898 89
rect 898 72 899 89
rect 932 175 933 192
rect 933 175 949 192
rect 985 72 1001 89
rect 1001 72 1002 89
rect 1034 175 1035 192
rect 1035 175 1051 192
rect 1087 72 1103 89
rect 1103 72 1104 89
rect 1136 175 1137 192
rect 1137 175 1153 192
rect 1188 72 1204 89
rect 1204 72 1205 89
rect 1238 175 1239 192
rect 1239 175 1255 192
rect 1290 72 1306 89
rect 1306 72 1307 89
rect 1339 175 1340 192
rect 1340 175 1356 192
rect 1393 73 1409 90
rect 1409 73 1410 90
rect 1441 175 1442 192
rect 1442 175 1458 192
rect 1553 498 1569 515
rect 1569 498 1571 515
rect 1596 497 1612 514
rect 1612 497 1614 514
rect 1553 461 1569 478
rect 1569 461 1571 478
rect 1596 461 1612 478
rect 1612 461 1614 478
rect 1553 423 1569 440
rect 1569 423 1570 440
rect 1596 424 1612 441
rect 1612 424 1613 441
rect 1524 375 1541 382
rect 1524 365 1541 375
rect 1524 329 1541 346
rect 1524 293 1541 310
rect 1524 257 1541 274
rect 1524 221 1541 238
rect 1524 185 1541 202
rect 1524 149 1541 166
rect 1524 113 1541 130
rect 1524 77 1541 94
rect 1524 41 1541 58
rect 1623 76 1640 93
rect 1693 575 1694 592
rect 1694 575 1710 592
rect 1693 538 1694 555
rect 1694 538 1710 555
rect 1744 498 1745 515
rect 1745 498 1762 515
rect 1744 461 1745 478
rect 1745 461 1762 478
rect 1744 425 1745 442
rect 1745 425 1762 442
rect 1801 594 1818 595
rect 1801 578 1802 594
rect 1802 578 1818 594
rect 1801 539 1802 556
rect 1802 539 1818 556
<< metal1 >>
rect 1686 646 1718 647
rect 1686 620 1689 646
rect 1715 620 1718 646
rect 1686 615 1718 620
rect 1794 646 1827 647
rect 1794 620 1797 646
rect 1823 620 1827 646
rect 1690 592 1713 615
rect 1794 614 1827 620
rect 1690 575 1693 592
rect 1710 575 1713 592
rect 1690 555 1713 575
rect 1690 538 1693 555
rect 1710 538 1713 555
rect 1690 532 1713 538
rect 1798 595 1821 614
rect 1798 578 1801 595
rect 1818 578 1821 595
rect 1798 556 1821 578
rect 1798 539 1801 556
rect 1818 539 1821 556
rect 1798 533 1821 539
rect 1548 517 1579 521
rect 1733 517 1766 521
rect 1548 515 1766 517
rect 1548 498 1553 515
rect 1571 514 1744 515
rect 1571 498 1596 514
rect 1548 497 1596 498
rect 1614 498 1744 514
rect 1762 498 1766 515
rect 1614 497 1766 498
rect 518 484 542 490
rect 518 467 522 484
rect 539 467 542 484
rect 518 448 542 467
rect 518 431 522 448
rect 539 431 542 448
rect 518 412 542 431
rect 1548 478 1765 497
rect 1548 461 1553 478
rect 1571 461 1596 478
rect 1614 461 1744 478
rect 1762 461 1765 478
rect 1548 460 1765 461
rect 1548 440 1568 460
rect 1594 450 1765 460
rect 1594 442 1766 450
rect 1594 441 1744 442
rect 1548 423 1553 440
rect 1594 434 1596 441
rect 1570 424 1596 434
rect 1613 425 1744 441
rect 1762 425 1766 442
rect 1613 424 1766 425
rect 1570 423 1766 424
rect 1548 417 1766 423
rect 518 395 522 412
rect 539 395 542 412
rect 492 382 542 395
rect 481 376 542 382
rect 481 359 484 376
rect 501 359 521 376
rect 538 359 542 376
rect 481 352 542 359
rect 481 340 495 352
rect 521 340 542 352
rect 481 323 484 340
rect 521 326 522 340
rect 501 323 522 326
rect 539 323 542 340
rect 481 320 542 323
rect 481 317 504 320
rect 518 317 542 320
rect 1507 382 1555 389
rect 1507 365 1524 382
rect 1541 365 1555 382
rect 1507 346 1555 365
rect 1507 329 1524 346
rect 1541 329 1555 346
rect 1507 310 1555 329
rect 1507 293 1524 310
rect 1541 293 1555 310
rect 1507 274 1555 293
rect 1507 257 1524 274
rect 1541 257 1555 274
rect 1507 238 1555 257
rect 1507 221 1524 238
rect 1541 221 1555 238
rect 1507 202 1555 221
rect 478 196 1471 199
rect 478 195 826 196
rect 478 191 724 195
rect 478 174 483 191
rect 500 174 625 191
rect 642 174 724 191
rect 478 169 724 174
rect 750 170 826 195
rect 852 170 928 196
rect 954 170 1030 196
rect 1056 170 1133 196
rect 1159 170 1234 196
rect 1260 170 1336 196
rect 1362 170 1438 196
rect 1464 170 1471 196
rect 750 169 1471 170
rect 478 165 1471 169
rect 1507 185 1524 202
rect 1541 185 1555 202
rect 1507 166 1555 185
rect 1507 149 1524 166
rect 1541 149 1555 166
rect 1507 130 1555 149
rect 519 112 544 118
rect 519 97 522 112
rect 515 95 522 97
rect 539 97 544 112
rect 567 114 594 121
rect 567 97 570 114
rect 587 97 594 114
rect 1507 113 1524 130
rect 1541 113 1555 130
rect 805 97 1416 98
rect 539 95 545 97
rect 515 94 545 95
rect 22 92 60 94
rect 22 66 28 92
rect 54 66 60 92
rect 22 63 60 66
rect 515 68 518 94
rect 544 68 545 94
rect 567 86 594 97
rect 515 65 522 68
rect 519 58 522 65
rect 539 65 545 68
rect 561 78 594 86
rect 539 58 544 65
rect 519 52 544 58
rect 561 61 569 78
rect 586 61 594 78
rect 669 95 1416 97
rect 669 94 877 95
rect 669 68 672 94
rect 698 68 776 94
rect 802 69 877 94
rect 903 69 979 95
rect 1005 69 1082 95
rect 1108 69 1184 95
rect 1210 69 1286 95
rect 1312 69 1388 95
rect 1414 69 1416 95
rect 802 68 1416 69
rect 669 65 1416 68
rect 1507 94 1555 113
rect 1507 77 1524 94
rect 1541 77 1555 94
rect 1507 72 1555 77
rect 1611 98 1653 107
rect 1611 72 1619 98
rect 1645 72 1653 98
rect 669 64 702 65
rect 561 42 594 61
rect 561 37 569 42
rect 586 37 594 42
rect 561 11 565 37
rect 591 11 594 37
rect 561 7 594 11
rect 1507 58 1561 72
rect 1611 65 1653 72
rect 1507 41 1524 58
rect 1541 41 1561 58
rect 1507 34 1561 41
rect 1507 8 1519 34
rect 1545 8 1561 34
rect 1507 5 1561 8
<< via1 >>
rect 1689 620 1715 646
rect 1797 620 1823 646
rect 1568 440 1594 460
rect 1568 434 1570 440
rect 1570 434 1594 440
rect 495 340 521 352
rect 495 326 501 340
rect 501 326 521 340
rect 724 192 750 195
rect 724 175 727 192
rect 727 175 744 192
rect 744 175 750 192
rect 724 169 750 175
rect 826 192 852 196
rect 826 175 829 192
rect 829 175 846 192
rect 846 175 852 192
rect 826 170 852 175
rect 928 192 954 196
rect 928 175 932 192
rect 932 175 949 192
rect 949 175 954 192
rect 928 170 954 175
rect 1030 192 1056 196
rect 1030 175 1034 192
rect 1034 175 1051 192
rect 1051 175 1056 192
rect 1030 170 1056 175
rect 1133 192 1159 196
rect 1133 175 1136 192
rect 1136 175 1153 192
rect 1153 175 1159 192
rect 1133 170 1159 175
rect 1234 192 1260 196
rect 1234 175 1238 192
rect 1238 175 1255 192
rect 1255 175 1260 192
rect 1234 170 1260 175
rect 1336 192 1362 196
rect 1336 175 1339 192
rect 1339 175 1356 192
rect 1356 175 1362 192
rect 1336 170 1362 175
rect 1438 192 1464 196
rect 1438 175 1441 192
rect 1441 175 1458 192
rect 1458 175 1464 192
rect 1438 170 1464 175
rect 28 86 54 92
rect 28 69 33 86
rect 33 69 50 86
rect 50 69 54 86
rect 28 66 54 69
rect 518 75 544 94
rect 518 68 522 75
rect 522 68 539 75
rect 539 68 544 75
rect 672 89 698 94
rect 672 72 678 89
rect 678 72 695 89
rect 695 72 698 89
rect 672 68 698 72
rect 776 89 802 94
rect 776 72 781 89
rect 781 72 798 89
rect 798 72 802 89
rect 776 68 802 72
rect 877 89 903 95
rect 877 72 882 89
rect 882 72 899 89
rect 899 72 903 89
rect 877 69 903 72
rect 979 89 1005 95
rect 979 72 985 89
rect 985 72 1002 89
rect 1002 72 1005 89
rect 979 69 1005 72
rect 1082 89 1108 95
rect 1082 72 1087 89
rect 1087 72 1104 89
rect 1104 72 1108 89
rect 1082 69 1108 72
rect 1184 89 1210 95
rect 1184 72 1188 89
rect 1188 72 1205 89
rect 1205 72 1210 89
rect 1184 69 1210 72
rect 1286 89 1312 95
rect 1286 72 1290 89
rect 1290 72 1307 89
rect 1307 72 1312 89
rect 1286 69 1312 72
rect 1388 90 1414 95
rect 1388 73 1393 90
rect 1393 73 1410 90
rect 1410 73 1414 90
rect 1388 69 1414 73
rect 1619 93 1645 98
rect 1619 76 1623 93
rect 1623 76 1640 93
rect 1640 76 1645 93
rect 1619 72 1645 76
rect 565 25 569 37
rect 569 25 586 37
rect 586 25 591 37
rect 565 11 591 25
rect 1519 8 1545 34
<< metal2 >>
rect 0 646 1908 650
rect 0 642 1689 646
rect 0 613 69 642
rect 172 620 1689 642
rect 1715 620 1797 646
rect 1823 620 1908 646
rect 172 613 1908 620
rect 0 612 1908 613
rect 64 610 177 612
rect 1848 558 1908 584
rect 1848 494 1908 520
rect 1554 460 1608 467
rect 1554 434 1568 460
rect 1594 434 1908 460
rect 1554 427 1608 434
rect 1848 380 1908 406
rect 483 354 542 356
rect 483 324 491 354
rect 526 352 542 354
rect 526 326 550 352
rect 1845 326 1908 352
rect 526 324 542 326
rect 483 321 542 324
rect 1848 274 1908 300
rect 1848 222 1908 248
rect 822 196 856 200
rect 925 196 959 200
rect 1026 196 1060 200
rect 1129 196 1163 200
rect 1231 196 1265 200
rect 1332 196 1366 200
rect 1433 196 1467 200
rect 609 195 826 196
rect 609 170 724 195
rect 721 169 724 170
rect 750 170 826 195
rect 852 170 928 196
rect 954 170 1030 196
rect 1056 170 1133 196
rect 1159 170 1234 196
rect 1260 170 1336 196
rect 1362 170 1438 196
rect 1464 170 1467 196
rect 1845 170 1908 196
rect 750 169 752 170
rect 721 166 752 169
rect 822 164 856 170
rect 925 164 959 170
rect 1026 164 1060 170
rect 1129 164 1163 170
rect 1231 164 1265 170
rect 1332 164 1366 170
rect 1433 164 1467 170
rect 1848 118 1908 144
rect 1613 98 1651 106
rect 514 94 546 97
rect 23 92 59 93
rect 514 92 518 94
rect 0 66 28 92
rect 54 66 59 92
rect 512 68 518 92
rect 544 92 546 94
rect 669 94 701 97
rect 669 92 672 94
rect 544 68 672 92
rect 698 92 701 94
rect 773 94 805 97
rect 773 92 776 94
rect 698 68 776 92
rect 802 92 805 94
rect 875 95 906 98
rect 875 92 877 95
rect 802 69 877 92
rect 903 92 906 95
rect 977 95 1008 98
rect 977 92 979 95
rect 903 69 979 92
rect 1005 92 1008 95
rect 1079 95 1110 98
rect 1079 92 1082 95
rect 1005 69 1082 92
rect 1108 92 1110 95
rect 1181 95 1213 98
rect 1181 92 1184 95
rect 1108 69 1184 92
rect 1210 92 1213 95
rect 1283 95 1314 98
rect 1283 92 1286 95
rect 1210 69 1286 92
rect 1312 92 1314 95
rect 1385 95 1416 98
rect 1385 92 1388 95
rect 1312 69 1388 92
rect 1414 92 1416 95
rect 1613 92 1619 98
rect 1414 72 1619 92
rect 1645 92 1651 98
rect 1645 72 1908 92
rect 1414 69 1908 72
rect 802 68 1908 69
rect 512 66 1908 68
rect 23 65 59 66
rect 514 64 546 66
rect 669 65 701 66
rect 773 65 805 66
rect 875 65 906 66
rect 1385 65 1416 66
rect 0 37 1908 40
rect 0 11 565 37
rect 591 34 1908 37
rect 591 11 1519 34
rect 0 8 1519 11
rect 1545 8 1908 34
rect 0 0 1908 8
<< via2 >>
rect 69 613 172 642
rect 491 352 526 354
rect 491 326 495 352
rect 495 326 521 352
rect 521 326 526 352
rect 491 324 526 326
<< metal3 >>
rect 64 642 177 645
rect 64 613 69 642
rect 172 613 177 642
rect 64 609 70 613
rect 171 609 177 613
rect 64 608 177 609
rect 23 357 472 565
rect 23 354 529 357
rect 23 324 491 354
rect 526 324 529 354
rect 23 321 529 324
rect 23 48 472 321
<< via3 >>
rect 70 613 171 641
rect 70 609 171 613
<< mimcap >>
rect 55 522 440 538
rect 55 489 71 522
rect 176 489 440 522
rect 55 70 440 489
<< mimcapcontact >>
rect 71 489 176 522
<< metal4 >>
rect 68 641 180 643
rect 68 609 70 641
rect 171 609 180 641
rect 68 522 180 609
rect 68 489 71 522
rect 176 489 180 522
rect 68 484 180 489
<< labels >>
rlabel metal2 1896 612 1908 650 0 VPWR
port 2 nsew
rlabel metal2 1898 0 1908 40 0 VGND
port 3 nsew
rlabel metal2 1900 66 1908 92 0 PBIAS
port 4 nsew
rlabel metal2 1899 434 1908 460 0 NBIAS
port 5 nsew
rlabel metal2 0 612 9 650 0 VPWR
port 2 nsew
rlabel metal2 0 0 12 40 0 VGND
port 3 nsew
rlabel metal2 0 66 12 92 0 RESIST
port 6 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
