magic
tech sky130A
timestamp 1607392100
<< error_s >>
rect -1540 1135 -1534 1141
rect -1435 1135 -1429 1141
rect -569 1135 -563 1141
rect -464 1135 -458 1141
rect 510 1135 516 1141
rect 615 1135 621 1141
rect -1114 1125 -1108 1131
rect -1061 1125 -1055 1131
rect -943 1125 -937 1131
rect -890 1125 -884 1131
rect 936 1125 942 1131
rect 989 1125 995 1131
rect -1546 1071 -1540 1077
rect -1429 1071 -1423 1077
rect -1120 1075 -1114 1081
rect -1055 1075 -1049 1081
rect -949 1075 -943 1081
rect -884 1075 -878 1081
rect -575 1071 -569 1077
rect -458 1071 -452 1077
rect 504 1071 510 1077
rect 621 1071 627 1077
rect 930 1075 936 1081
rect 995 1075 1001 1081
rect -1540 1018 -1534 1024
rect -1435 1018 -1429 1024
rect -1114 1016 -1108 1022
rect -1061 1016 -1055 1022
rect -943 1016 -937 1022
rect -890 1016 -884 1022
rect -569 1018 -563 1024
rect -464 1018 -458 1024
rect 510 1018 516 1024
rect 615 1018 621 1024
rect 936 1016 942 1022
rect 989 1016 995 1022
rect -1120 966 -1114 972
rect -1055 966 -1049 972
rect -949 966 -943 972
rect -884 966 -878 972
rect 930 966 936 972
rect 995 966 1001 972
rect -1771 958 -1758 963
rect -1757 958 -1744 962
rect -1771 955 -1744 958
rect -1546 954 -1540 960
rect -1429 954 -1423 960
rect -575 954 -569 960
rect -458 954 -452 960
rect -254 958 -241 962
rect -240 958 -227 963
rect -254 955 -227 958
rect 504 954 510 960
rect 621 954 627 960
rect -1540 833 -1534 839
rect -1435 833 -1429 839
rect -569 833 -563 839
rect -464 833 -458 839
rect 510 833 516 839
rect 615 833 621 839
rect -1114 827 -1108 833
rect -1061 827 -1055 833
rect -943 827 -937 833
rect -890 827 -884 833
rect 936 827 942 833
rect 989 827 995 833
rect -1120 777 -1114 783
rect -1055 777 -1049 783
rect -949 777 -943 783
rect -884 777 -878 783
rect 930 777 936 783
rect 995 777 1001 783
rect -1546 769 -1540 775
rect -1429 769 -1423 775
rect -575 769 -569 775
rect -458 769 -452 775
rect 504 769 510 775
rect 621 769 627 775
rect -1540 717 -1534 723
rect -1435 717 -1429 723
rect -569 717 -563 723
rect -464 717 -458 723
rect -1114 710 -1108 716
rect -1061 710 -1055 716
rect -943 710 -937 716
rect -890 710 -884 716
rect -29 714 -28 726
rect 510 717 516 723
rect 615 717 621 723
rect -15 700 -14 712
rect 936 710 942 716
rect 989 710 995 716
rect -1120 660 -1114 666
rect -1055 660 -1049 666
rect -949 660 -943 666
rect -884 660 -878 666
rect 930 660 936 666
rect 995 660 1001 666
rect -1546 653 -1540 659
rect -1429 653 -1423 659
rect -575 653 -569 659
rect -458 653 -452 659
rect 504 653 510 659
rect 621 653 627 659
rect -1866 613 -1864 621
rect 184 613 185 621
rect -1953 600 -1952 608
rect -1872 600 -1871 608
rect -110 602 -109 608
rect -110 594 -108 602
rect -29 600 -28 608
rect -1537 537 -1531 543
rect -1432 537 -1426 543
rect -566 537 -560 543
rect -461 537 -455 543
rect 512 537 518 543
rect 617 537 623 543
rect -1111 527 -1105 533
rect -1058 527 -1052 533
rect -940 527 -934 533
rect -887 527 -881 533
rect 938 527 944 533
rect 991 527 997 533
rect -1543 473 -1537 479
rect -1426 473 -1420 479
rect -1117 477 -1111 483
rect -1052 477 -1046 483
rect -946 477 -940 483
rect -881 477 -875 483
rect -572 473 -566 479
rect -455 473 -449 479
rect 506 473 512 479
rect 623 473 629 479
rect 932 477 938 483
rect 997 477 1003 483
rect -1537 420 -1531 426
rect -1432 420 -1426 426
rect -1111 418 -1105 424
rect -1058 418 -1052 424
rect -940 418 -934 424
rect -887 418 -881 424
rect -566 420 -560 426
rect -461 420 -455 426
rect 512 420 518 426
rect 617 420 623 426
rect 938 418 944 424
rect 991 418 997 424
rect -1117 368 -1111 374
rect -1052 368 -1046 374
rect -946 368 -940 374
rect -881 368 -875 374
rect 932 368 938 374
rect 997 368 1003 374
rect -1768 360 -1755 365
rect -1754 360 -1741 364
rect -1768 357 -1741 360
rect -1543 356 -1537 362
rect -1426 356 -1420 362
rect -572 356 -566 362
rect -455 356 -449 362
rect -251 360 -238 364
rect -237 360 -224 365
rect -251 357 -224 360
rect 506 356 512 362
rect 623 356 629 362
rect -1537 235 -1531 241
rect -1432 235 -1426 241
rect -566 235 -560 241
rect -461 235 -455 241
rect 512 235 518 241
rect 617 235 623 241
rect -1111 229 -1105 235
rect -1058 229 -1052 235
rect -940 229 -934 235
rect -887 229 -881 235
rect 938 229 944 235
rect 991 229 997 235
rect -1117 179 -1111 185
rect -1052 179 -1046 185
rect -946 179 -940 185
rect -881 179 -875 185
rect 932 179 938 185
rect 997 179 1003 185
rect -1543 171 -1537 177
rect -1426 171 -1420 177
rect -572 171 -566 177
rect -455 171 -449 177
rect 506 171 512 177
rect 623 171 629 177
rect -1537 119 -1531 125
rect -1432 119 -1426 125
rect -566 119 -560 125
rect -461 119 -455 125
rect -1111 112 -1105 118
rect -1058 112 -1052 118
rect -940 112 -934 118
rect -887 112 -881 118
rect -27 116 -25 128
rect 512 119 518 125
rect 617 119 623 125
rect -27 68 -26 116
rect -13 102 -11 114
rect 938 112 944 118
rect 991 112 997 118
rect -13 82 -12 102
rect -1117 62 -1111 68
rect -1052 62 -1046 68
rect -946 62 -940 68
rect -881 62 -875 68
rect 932 62 938 68
rect 997 62 1003 68
rect -1543 55 -1537 61
rect -1426 55 -1420 61
rect -572 55 -566 61
rect -455 55 -449 61
rect 506 55 512 61
rect 623 55 629 61
use sky130_hilas_WTA4stage01  sky130_hilas_WTA4stage01_1
timestamp 1607392100
transform 1 0 1106 0 1 636
box -1121 -43 296 562
use sky130_hilas_WTA4stage01  sky130_hilas_WTA4stage01_0
timestamp 1607392100
transform 1 0 1108 0 1 38
box -1121 -43 296 562
use sky130_hilas_swc4x2cell  sky130_hilas_swc4x2cell_1
timestamp 1607392100
transform 1 0 -1001 0 1 597
box -1004 -4 1008 601
use sky130_hilas_swc4x2cell  sky130_hilas_swc4x2cell_0
timestamp 1607392100
transform 1 0 -998 0 1 -1
box -1004 -4 1008 601
<< end >>
