magic
tech sky130A
timestamp 1628617005
<< checkpaint >>
rect -630 608 4720 2962
rect 267 263 4574 608
rect 2429 216 4574 263
rect 2429 -176 4371 216
rect 2429 -630 4238 -176
<< error_s >>
rect 964 1475 1014 1481
rect 1036 1475 1086 1481
rect 3004 1475 3054 1481
rect 3076 1475 3126 1481
rect 3464 1479 3491 1485
rect 964 1433 1014 1439
rect 1036 1433 1086 1439
rect 3004 1433 3054 1439
rect 3076 1433 3126 1439
rect 3464 1437 3491 1443
rect 3464 1412 3491 1418
rect 3464 1370 3491 1376
rect 3464 1329 3491 1335
rect 3464 1287 3491 1293
rect 3464 1262 3491 1268
rect 3464 1220 3491 1226
rect 3464 1179 3491 1185
rect 3464 1137 3491 1143
rect 3464 1112 3491 1118
rect 3464 1070 3491 1076
rect 3464 1029 3491 1035
rect 3464 987 3491 993
rect 964 962 1014 968
rect 1036 962 1086 968
rect 3004 962 3054 968
rect 3076 962 3126 968
rect 3464 962 3491 968
rect 964 920 1014 926
rect 1036 920 1086 926
rect 3004 920 3054 926
rect 3076 920 3126 926
rect 3464 920 3491 926
<< nwell >>
rect 897 1502 1095 1503
rect 3193 1502 3340 1503
rect 3578 1485 3706 1503
rect 897 1435 904 1453
rect 897 948 905 966
rect 3578 898 3706 917
<< locali >>
rect 1746 1239 1766 1246
rect 1746 1222 1747 1239
rect 1764 1222 1766 1239
rect 1746 1167 1766 1222
rect 1746 1150 1748 1167
rect 1765 1150 1766 1167
rect 1746 1145 1766 1150
rect 2321 1239 2350 1246
rect 2321 1222 2326 1239
rect 2343 1222 2350 1239
rect 2321 1167 2350 1222
rect 2321 1150 2326 1167
rect 2343 1150 2350 1167
rect 2321 1145 2350 1150
<< viali >>
rect 1747 1222 1764 1239
rect 1748 1150 1765 1167
rect 2326 1222 2343 1239
rect 2326 1150 2343 1167
<< metal1 >>
rect 921 1498 949 1503
rect 921 1497 953 1498
rect 974 1497 993 1503
rect 921 1471 924 1497
rect 950 1471 953 1497
rect 1622 1494 1645 1502
rect 1744 1494 1767 1502
rect 1973 1487 2117 1503
rect 2323 1494 2346 1503
rect 2445 1495 2468 1503
rect 3097 1495 3116 1503
rect 3141 1498 3169 1503
rect 3141 1496 3173 1498
rect 921 1470 953 1471
rect 3141 1470 3144 1496
rect 3170 1470 3173 1496
rect 3510 1489 3544 1503
rect 3576 1488 3604 1503
rect 3141 1468 3173 1470
rect 1747 1221 1764 1222
rect 2326 1221 2343 1222
rect 1745 1190 1777 1192
rect 1745 1151 1748 1190
rect 1774 1164 1777 1190
rect 1765 1162 1777 1164
rect 2315 1184 2347 1187
rect 1765 1151 1769 1162
rect 2315 1158 2318 1184
rect 2344 1158 2347 1184
rect 2315 1155 2326 1158
rect 1767 1145 1769 1151
rect 2343 1155 2347 1158
rect 3359 945 3392 947
rect 2315 932 2347 934
rect 2315 906 2318 932
rect 2344 906 2347 932
rect 3359 919 3362 945
rect 3389 919 3392 945
rect 3359 918 3392 919
rect 2315 904 2347 906
rect 3358 915 3400 918
rect 3460 917 3510 918
rect 3460 915 3544 917
rect 3358 904 3544 915
rect 3097 898 3116 903
rect 3141 898 3169 903
rect 3386 901 3476 904
rect 3510 898 3544 904
rect 3577 898 3604 919
<< via1 >>
rect 924 1471 950 1497
rect 3144 1470 3170 1496
rect 1748 1167 1774 1190
rect 1748 1164 1765 1167
rect 1765 1164 1774 1167
rect 2318 1167 2344 1184
rect 2318 1158 2326 1167
rect 2326 1158 2343 1167
rect 2343 1158 2344 1167
rect 2318 906 2344 932
rect 3362 919 3389 945
<< metal2 >>
rect 921 1497 953 1498
rect 921 1471 924 1497
rect 950 1486 953 1497
rect 3141 1496 3173 1498
rect 3141 1486 3144 1496
rect 950 1471 3144 1486
rect 921 1470 3144 1471
rect 3170 1470 3173 1496
rect 3253 1476 3284 1500
rect 921 1468 3173 1470
rect 897 1435 904 1453
rect 3364 1413 3386 1415
rect 1787 1375 1871 1395
rect 3359 1379 3386 1413
rect 1832 1328 2846 1350
rect 3185 1329 3220 1351
rect 1827 1231 2728 1253
rect 1745 1190 1777 1192
rect 1745 1164 1748 1190
rect 1774 1187 1777 1190
rect 1774 1184 2347 1187
rect 1774 1164 2318 1184
rect 1745 1162 2318 1164
rect 2315 1158 2318 1162
rect 2344 1158 2347 1184
rect 2315 1155 2347 1158
rect 1832 1053 2398 1075
rect 1782 1023 1830 1024
rect 1782 999 1871 1023
rect 2376 1020 2398 1053
rect 2706 1070 2728 1231
rect 2824 1208 2846 1328
rect 3366 1322 3386 1323
rect 3366 1289 3388 1322
rect 3368 1288 3388 1289
rect 3261 1209 3293 1233
rect 3695 1232 3706 1255
rect 2821 1204 2846 1208
rect 2821 1140 2847 1204
rect 3695 1150 3706 1172
rect 2821 1119 3234 1140
rect 3213 1105 3234 1119
rect 3213 1084 3415 1105
rect 2706 1048 2991 1070
rect 2813 1020 3415 1025
rect 2376 1004 3415 1020
rect 2376 998 2852 1004
rect 897 948 905 966
rect 3359 945 3392 947
rect 2315 933 2347 934
rect 3359 933 3362 945
rect 2315 932 3362 933
rect 2315 906 2318 932
rect 2344 919 3362 932
rect 3389 919 3392 945
rect 2344 917 3392 919
rect 2344 916 2384 917
rect 2344 906 2347 916
rect 2315 904 2347 906
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1628616992
transform 1 0 3551 0 1 939
box 0 0 358 746
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1628616992
transform 1 0 3059 0 -1 1063
box 0 0 549 1063
use sky130_hilas_FGBias2x1cell  sky130_hilas_FGBias2x1cell_0
timestamp 1628616997
transform 1 0 2436 0 1 1280
box 0 0 1654 1052
use sky130_hilas_FGBiasWeakGate2x1cell  sky130_hilas_FGBiasWeakGate2x1cell_0
timestamp 1628616992
transform -1 0 1654 0 1 1280
box 0 0 1654 1052
<< labels >>
rlabel metal2 1787 1375 1823 1394 0 VIN11
port 2 nsew analog default
rlabel metal2 1782 999 1818 1024 0 VIN12
port 1 nsew analog default
rlabel metal1 3510 1497 3544 1503 0 VGND
port 7 nsew analog default
rlabel metal1 3576 1497 3604 1503 0 VPWR
port 6 nsew analog default
rlabel metal1 3577 898 3604 904 0 VPWR
port 6 nsew power default
rlabel metal1 3510 898 3544 904 0 VGND
port 7 nsew ground default
rlabel metal2 3261 1209 3293 1233 0 VIN21
port 3 nsew analog default
rlabel metal2 3253 1476 3284 1500 1 VIN22
port 4 n analog default
rlabel metal1 3141 1495 3169 1503 0 VINJ
port 8 nsew power default
rlabel metal1 3141 898 3169 903 0 VINJ
port 8 nsew power default
rlabel metal2 3695 1232 3706 1255 0 OUTPUT1
port 9 nsew analog default
rlabel metal2 3695 1150 3706 1172 0 OUTPUT2
port 10 nsew analog default
rlabel metal2 897 1435 904 1453 0 DRAIN1
port 11 nsew
rlabel metal2 897 948 905 966 0 DRAIN2
port 12 nsew
rlabel metal1 921 1496 949 1503 0 VINJ
port 8 nsew
rlabel metal1 974 1497 993 1503 0 COLSEL2
port 13 nsew
rlabel metal1 1622 1494 1645 1502 0 GATE2
port 14 nsew
rlabel metal1 1744 1494 1767 1502 0 VGND
port 7 nsew
rlabel metal1 2445 1495 2468 1503 0 GATE1
port 15 nsew
rlabel metal1 2323 1495 2346 1503 0 VGND
port 7 nsew
rlabel metal1 3097 1495 3116 1503 0 COLSEL1
port 16 nsew
rlabel metal1 3097 898 3116 903 0 COLSEL1
port 16 nsew
rlabel metal1 2015 1491 2075 1503 0 VTUN
port 17 nsew
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
