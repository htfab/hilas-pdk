magic
tech sky130A
timestamp 1628704380
<< nwell >>
rect 0 30 219 203
<< pmos >>
rect 21 82 89 112
rect 125 82 193 112
<< pdiff >>
rect 21 136 89 142
rect 21 119 29 136
rect 47 119 65 136
rect 83 119 89 136
rect 21 112 89 119
rect 125 136 193 142
rect 125 119 133 136
rect 151 119 170 136
rect 189 119 193 136
rect 125 112 193 119
rect 21 75 89 82
rect 21 58 29 75
rect 47 58 65 75
rect 83 58 89 75
rect 21 49 89 58
rect 125 75 193 82
rect 125 58 131 75
rect 149 58 167 75
rect 185 58 193 75
rect 125 54 193 58
rect 132 49 193 54
<< pdiffc >>
rect 29 119 47 136
rect 65 119 83 136
rect 133 119 151 136
rect 170 119 189 136
rect 29 58 47 75
rect 65 58 83 75
rect 131 58 149 75
rect 167 58 185 75
<< nsubdiff >>
rect 21 171 89 183
rect 21 154 29 171
rect 47 154 65 171
rect 83 154 89 171
rect 21 142 89 154
rect 125 171 193 183
rect 125 154 133 171
rect 151 154 170 171
rect 189 154 193 171
rect 125 142 193 154
<< nsubdiffcont >>
rect 29 154 47 171
rect 65 154 83 171
rect 133 154 151 171
rect 170 154 189 171
<< poly >>
rect 8 82 21 112
rect 89 82 125 112
rect 193 82 206 112
rect 97 38 114 82
rect 91 30 118 38
rect 91 13 96 30
rect 113 13 118 30
rect 91 5 118 13
<< polycont >>
rect 96 13 113 30
<< locali >>
rect 21 154 29 171
rect 47 154 65 171
rect 83 154 133 171
rect 151 154 170 171
rect 189 154 197 171
rect 21 136 197 154
rect 21 119 29 136
rect 47 119 65 136
rect 83 119 133 136
rect 151 119 170 136
rect 189 119 197 136
rect 21 58 29 75
rect 47 58 65 75
rect 83 58 92 75
rect 123 58 131 75
rect 149 58 167 75
rect 185 58 193 75
rect 56 41 92 58
rect 56 30 121 41
rect 56 13 96 30
rect 113 13 121 30
rect 56 5 121 13
rect 56 0 83 5
rect 146 0 171 58
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
