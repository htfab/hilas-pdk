magic
tech sky130A
timestamp 1628164971
<< nmos >>
rect 0 -6 27 36
<< ndiff >>
rect -31 20 0 36
rect -31 3 -26 20
rect -6 3 0 20
rect -31 -6 0 3
rect 27 20 58 36
rect 27 3 33 20
rect 53 3 58 20
rect 27 -6 58 3
<< ndiffc >>
rect -26 3 -6 20
rect 33 3 53 20
<< poly >>
rect 0 36 27 49
rect 0 -14 27 -6
rect -81 -19 27 -14
rect -81 -36 -73 -19
rect -56 -29 27 -19
rect -56 -36 -48 -29
rect -81 -41 -48 -36
<< polycont >>
rect -73 -36 -56 -19
<< locali >>
rect -26 20 -6 28
rect -26 -5 -6 3
rect 33 20 53 28
rect 33 -5 53 3
rect -81 -36 -73 -19
rect -56 -36 -48 -19
<< metal2 >>
rect -111 2 -51 19
rect 75 3 97 20
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628164971
transform 1 0 65 0 1 11
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628164971
transform 1 0 -44 0 1 10
box -14 -15 20 18
<< end >>
