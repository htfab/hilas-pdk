* NGSPICE file created from /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_swc4x2cellOverlap.ext - technology: sky130A

.subckt sky130_hilas_nOverlapCap01 VSUBS a_n114_n76# a_n24_14#
X0 a_n24_14# a_n114_n76# a_n24_14# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=580000u l=1.86e+06u
.ends

.subckt sky130_hilas_horizPcell01 VSUBS a_n502_286# a_n508_162# w_n578_94# a_n578_238#
+ m1_n258_94# a_n300_94# a_n344_286#
X0 w_n578_94# a_n300_94# a_n344_162# w_n578_94# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
X1 a_n344_286# a_n578_238# a_n502_286# w_n578_94# sky130_fd_pr__pfet_g5v0d10v5 w=300000u l=500000u
X2 a_n344_162# a_n578_238# a_n508_162# w_n578_94# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
.ends

.subckt sky130_hilas_overlapCap02a VSUBS a_n1004_n70# w_n1042_n108# a_n908_28#
X0 a_n908_28# a_n1004_n70# a_n908_28# w_n1042_n108# sky130_fd_pr__pfet_g5v0d10v5 w=465000u l=500000u
.ends

.subckt sky130_hilas_swc4x1cellOverlap2 VSUBS m2_n382_24# a_1264_n176# sky130_hilas_overlapCap02a_3/a_n908_28#
+ m2_n382_n572# m2_n382_n62# sky130_hilas_overlapCap02a_2/a_n908_28# m2_n382_310#
+ m2_n382_224# sky130_hilas_overlapCap02a_1/a_n908_28# sky130_hilas_horizPcell01_3/a_n344_286#
+ sky130_hilas_overlapCap02a_0/a_n908_28# m2_n382_n292# m2_n382_n660# m1_n180_n764#
+ w_1264_n176# m2_n382_n376#
Xsky130_hilas_nOverlapCap01_0 VSUBS a_n38_228# m1_n180_n764# sky130_hilas_nOverlapCap01
Xsky130_hilas_horizPcell01_0 VSUBS m2_n382_24# m2_n382_n62# w_1264_n176# a_n38_10#
+ a_1264_n176# a_1264_n176# sky130_hilas_horizPcell01_3/a_n344_286# sky130_hilas_horizPcell01
Xsky130_hilas_nOverlapCap01_1 VSUBS a_n38_10# m1_n180_n764# sky130_hilas_nOverlapCap01
Xsky130_hilas_horizPcell01_1 VSUBS m2_n382_n572# m2_n382_n660# w_1264_n176# a_n38_n590#
+ a_1264_n176# a_1264_n176# sky130_hilas_horizPcell01_3/a_n344_286# sky130_hilas_horizPcell01
Xsky130_hilas_horizPcell01_2 VSUBS m2_n382_n376# m2_n382_n292# w_1264_n176# a_n38_n350#
+ a_1264_n176# a_1264_n176# sky130_hilas_horizPcell01_3/a_n344_286# sky130_hilas_horizPcell01
Xsky130_hilas_nOverlapCap01_2 VSUBS a_n38_n350# m1_n180_n764# sky130_hilas_nOverlapCap01
Xsky130_hilas_horizPcell01_3 VSUBS m2_n382_224# m2_n382_310# w_1264_n176# a_n38_228#
+ a_1264_n176# a_1264_n176# sky130_hilas_horizPcell01_3/a_n344_286# sky130_hilas_horizPcell01
Xsky130_hilas_nOverlapCap01_3 VSUBS a_n38_n590# m1_n180_n764# sky130_hilas_nOverlapCap01
Xsky130_hilas_overlapCap02a_0 VSUBS a_n38_228# w_1264_n176# sky130_hilas_overlapCap02a_0/a_n908_28#
+ sky130_hilas_overlapCap02a
Xsky130_hilas_overlapCap02a_1 VSUBS a_n38_10# w_1264_n176# sky130_hilas_overlapCap02a_1/a_n908_28#
+ sky130_hilas_overlapCap02a
Xsky130_hilas_overlapCap02a_2 VSUBS a_n38_n350# w_1264_n176# sky130_hilas_overlapCap02a_2/a_n908_28#
+ sky130_hilas_overlapCap02a
Xsky130_hilas_overlapCap02a_3 VSUBS a_n38_n590# w_1264_n176# sky130_hilas_overlapCap02a_3/a_n908_28#
+ sky130_hilas_overlapCap02a
.ends

.subckt home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_swc4x2cellOverlap
+ Vert1 Horiz1 drain1 Horiz2 drain2 drain3 Horiz3 Horiz4 drain4 Vinj GateSelect1 Vert2
+ GateSelect2 Gate2 Gate1 Vtun
Xsky130_hilas_swc4x1cellOverlap2_0 VSUBS Horiz2 GateSelect2 Gate2 Horiz4 drain2 Gate2
+ drain1 Horiz1 Gate2 Vert2 Gate2 drain3 drain4 Vtun Vinj Horiz3 sky130_hilas_swc4x1cellOverlap2
Xsky130_hilas_swc4x1cellOverlap2_1 VSUBS Horiz2 GateSelect1 Gate1 Horiz4 drain2 Gate1
+ drain1 Horiz1 Gate1 Vert1 Gate1 drain3 drain4 Vtun Vinj Horiz3 sky130_hilas_swc4x1cellOverlap2
.ends

