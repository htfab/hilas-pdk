* NGSPICE file created from /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_capacitorSize02.ext - technology: sky130A

.subckt sky130_hilas_CapModule03 m3_n784_n490# $SUB c1_n664_n410#
X0 c1_n664_n410# m3_n784_n490# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=3.22e+06u
.ends

.subckt home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_capacitorSize02
+ CapTerm02 CapTerm01
Xsky130_hilas_CapModule03_0 CapTerm02 $SUB CapTerm01 sky130_hilas_CapModule03
.ends

