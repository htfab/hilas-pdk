magic
tech sky130A
timestamp 1634057795
<< checkpaint >>
rect -630 -630 2887 1682
<< mvnmos >>
rect 3184 1139 3234 1379
rect 3184 863 3234 1103
<< mvndiff >>
rect 3155 1374 3184 1379
rect 3155 1159 3161 1374
rect 3178 1159 3184 1374
rect 3155 1139 3184 1159
rect 3234 1373 3271 1379
rect 3234 1159 3240 1373
rect 3257 1168 3271 1373
rect 3257 1159 3283 1168
rect 3234 1141 3283 1159
rect 3234 1139 3260 1141
rect 3254 1103 3260 1139
rect 3155 1083 3184 1103
rect 3155 873 3161 1083
rect 3178 873 3184 1083
rect 3155 863 3184 873
rect 3234 1100 3260 1103
rect 3277 1100 3283 1141
rect 3234 1083 3283 1100
rect 3234 873 3240 1083
rect 3257 1074 3283 1083
rect 3257 873 3271 1074
rect 3234 863 3271 873
<< mvndiffc >>
rect 3161 1159 3178 1374
rect 3240 1159 3257 1373
rect 3161 873 3178 1083
rect 3260 1100 3277 1141
rect 3240 873 3257 1083
<< psubdiff >>
rect 3271 1360 3314 1379
rect 3271 1184 3284 1360
rect 3302 1184 3314 1360
rect 3271 1168 3314 1184
rect 3271 1067 3314 1074
rect 3271 875 3284 1067
rect 3302 875 3314 1067
rect 3271 863 3314 875
<< psubdiffcont >>
rect 3284 1184 3302 1360
rect 3284 875 3302 1067
<< poly >>
rect 2688 1398 2775 1420
rect 2688 852 2721 854
rect 2688 835 2696 852
rect 2713 835 2721 852
rect 2688 830 2721 835
rect 2797 1398 2885 1420
rect 2742 830 2830 854
rect 2907 1398 2995 1420
rect 2852 830 2940 854
rect 3017 1398 3105 1420
rect 2962 830 3050 854
rect 3184 1415 3234 1420
rect 3184 1398 3200 1415
rect 3217 1398 3234 1415
rect 3184 1379 3234 1398
rect 3184 1103 3234 1139
rect 3072 852 3105 854
rect 3072 835 3080 852
rect 3097 835 3105 852
rect 3072 830 3105 835
rect 3184 830 3234 863
<< polycont >>
rect 2696 835 2713 852
rect 3200 1398 3217 1415
rect 3080 835 3097 852
<< npolyres >>
rect 2688 854 2721 1398
rect 2742 854 2775 1398
rect 2797 854 2830 1398
rect 2852 854 2885 1398
rect 2907 854 2940 1398
rect 2962 854 2995 1398
rect 3017 854 3050 1398
rect 3072 854 3105 1398
<< locali >>
rect 3132 1398 3200 1415
rect 3217 1398 3225 1415
rect 3132 1374 3180 1398
rect 3132 1369 3161 1374
rect 3132 1159 3136 1369
rect 3154 1159 3161 1369
rect 3178 1159 3180 1374
rect 3132 1151 3180 1159
rect 3238 1373 3302 1381
rect 3238 1159 3240 1373
rect 3257 1360 3302 1373
rect 3257 1184 3284 1360
rect 3257 1159 3302 1184
rect 3238 1141 3302 1159
rect 3238 1100 3260 1141
rect 3277 1100 3302 1141
rect 3129 1083 3180 1091
rect 3042 899 3078 909
rect 3042 882 3053 899
rect 3070 882 3078 899
rect 3042 871 3078 882
rect 2667 852 2721 853
rect 2667 851 2696 852
rect 2667 834 2670 851
rect 2687 835 2696 851
rect 2713 835 2721 852
rect 3052 852 3078 871
rect 3129 873 3136 1083
rect 3154 873 3161 1083
rect 3178 873 3180 1083
rect 3129 866 3180 873
rect 3159 865 3180 866
rect 3238 1083 3302 1100
rect 3238 873 3240 1083
rect 3257 1067 3302 1083
rect 3257 930 3284 1067
rect 3257 913 3265 930
rect 3282 913 3284 930
rect 3257 893 3284 913
rect 3257 876 3265 893
rect 3282 876 3284 893
rect 3257 875 3284 876
rect 3257 873 3302 875
rect 3238 866 3302 873
rect 3238 865 3289 866
rect 3257 856 3289 865
rect 3052 835 3080 852
rect 3097 835 3105 852
rect 3257 839 3265 856
rect 3282 839 3289 856
rect 3257 836 3289 839
rect 2687 834 2721 835
rect 2667 831 2721 834
<< viali >>
rect 3136 1159 3154 1369
rect 3053 882 3070 899
rect 2670 834 2687 851
rect 3136 873 3154 1083
rect 3265 913 3282 930
rect 3265 876 3282 893
rect 3265 839 3282 856
<< metal1 >>
rect 3130 1369 3170 1376
rect 3130 1362 3136 1369
rect 3154 1362 3170 1369
rect 3130 1168 3135 1362
rect 3164 1168 3170 1362
rect 3130 1159 3136 1168
rect 3154 1159 3170 1168
rect 3130 1155 3170 1159
rect 2660 1146 2686 1149
rect 2660 1117 2686 1120
rect 2664 868 2685 1117
rect 3131 1084 3162 1089
rect 3131 1083 3174 1084
rect 3042 905 3078 909
rect 3042 879 3048 905
rect 3074 879 3078 905
rect 3042 871 3078 879
rect 3131 873 3136 1083
rect 3154 1077 3174 1083
rect 3168 967 3174 1077
rect 3154 873 3174 967
rect 3131 872 3174 873
rect 3255 930 3291 933
rect 3255 913 3265 930
rect 3282 913 3291 930
rect 3255 893 3291 913
rect 3255 876 3265 893
rect 3282 876 3291 893
rect 2664 862 2686 868
rect 3131 867 3162 872
rect 2664 854 2689 862
rect 3255 856 3291 876
rect 2664 851 2693 854
rect 2664 834 2670 851
rect 2687 834 2693 851
rect 2664 831 2693 834
rect 3255 844 3265 856
rect 3282 844 3291 856
rect 3255 818 3260 844
rect 3286 818 3291 844
rect 3255 813 3291 818
<< via1 >>
rect 3135 1168 3136 1362
rect 3136 1168 3154 1362
rect 3154 1168 3164 1362
rect 2660 1120 2686 1146
rect 3048 899 3074 905
rect 3048 882 3053 899
rect 3053 882 3070 899
rect 3070 882 3074 899
rect 3048 879 3074 882
rect 3142 967 3154 1077
rect 3154 967 3168 1077
rect 3260 839 3265 844
rect 3265 839 3282 844
rect 3282 839 3286 844
rect 3260 818 3286 839
<< metal2 >>
rect 3132 1362 3166 1367
rect 3132 1238 3135 1362
rect 2633 1219 3135 1238
rect 3132 1168 3135 1219
rect 3164 1218 3166 1362
rect 3164 1192 3338 1218
rect 3164 1168 3166 1192
rect 3132 1158 3166 1168
rect 2659 1146 2687 1150
rect 2657 1144 2660 1146
rect 2629 1121 2660 1144
rect 2657 1120 2660 1121
rect 2686 1120 2689 1146
rect 2659 1116 2687 1120
rect 3131 1077 3175 1091
rect 3131 1052 3142 1077
rect 2633 1033 3142 1052
rect 3131 967 3142 1033
rect 3168 1060 3175 1077
rect 3168 1034 3338 1060
rect 3168 1033 3217 1034
rect 3168 967 3175 1033
rect 3131 964 3175 967
rect 3044 905 3078 909
rect 3044 879 3048 905
rect 3074 904 3078 905
rect 3074 879 3338 904
rect 3044 878 3338 879
rect 3044 875 3078 878
rect 3147 844 3338 852
rect 3147 818 3260 844
rect 3286 818 3338 844
rect 3147 812 3338 818
use sky130_hilas_FGtrans2x1cell2  sky130_hilas_FGtrans2x1cell2_0
timestamp 1634057748
transform -1 0 2257 0 -1 1052
box 0 0 2257 1052
<< labels >>
rlabel metal2 3325 1192 3338 1218 0 NBIAS
port 1 nsew
rlabel metal2 3326 1034 3338 1060 0 PBIAS
port 2 nsew
rlabel metal2 3328 812 3338 852 0 VGND
port 3 nsew
rlabel metal2 3328 878 3338 904 0 RESIST
port 4 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
