magic
tech sky130A
timestamp 1627742263
<< error_p >>
rect 410 83 460 92
rect 460 77 491 83
rect 567 77 595 93
rect 709 77 737 93
rect 678 51 683 56
rect 410 41 460 50
rect 567 35 595 51
rect 709 35 737 51
rect 338 15 389 25
rect 306 10 325 15
rect 518 14 546 31
rect 758 14 786 31
rect 306 -17 311 10
rect 389 -17 420 -11
rect 338 -27 389 -17
rect 518 -28 546 -11
rect 758 -28 786 -11
<< nwell >>
rect 659 -40 836 119
<< nmos >>
rect 567 51 595 77
rect 518 -11 546 14
<< pmos >>
rect 709 51 737 77
rect 758 -11 786 14
<< mvnmos >>
rect 410 50 460 83
rect 338 -17 389 15
<< ndiff >>
rect 533 72 567 77
rect 533 55 544 72
rect 561 55 567 72
rect 533 51 567 55
rect 595 72 624 77
rect 595 55 601 72
rect 618 55 624 72
rect 595 51 624 55
rect 489 10 518 14
rect 489 -7 495 10
rect 512 -7 518 10
rect 489 -11 518 -7
rect 546 10 575 14
rect 546 -7 552 10
rect 569 -7 575 10
rect 546 -11 575 -7
<< pdiff >>
rect 678 72 709 77
rect 678 55 684 72
rect 702 55 709 72
rect 678 51 709 55
rect 737 72 773 77
rect 737 55 743 72
rect 760 55 773 72
rect 737 51 773 55
rect 729 10 758 14
rect 729 -7 735 10
rect 752 -7 758 10
rect 729 -11 758 -7
rect 786 10 817 14
rect 786 -7 793 10
rect 810 -7 817 10
rect 786 -11 817 -7
<< mvndiff >>
rect 382 75 410 83
rect 382 58 386 75
rect 404 58 410 75
rect 382 50 410 58
rect 460 75 491 83
rect 460 58 466 75
rect 484 58 491 75
rect 460 50 491 58
rect 306 7 338 15
rect 306 -10 313 7
rect 331 -10 338 7
rect 306 -17 338 -10
rect 389 5 420 15
rect 389 -12 395 5
rect 413 -12 420 5
rect 389 -17 420 -12
<< ndiffc >>
rect 544 55 561 72
rect 601 55 618 72
rect 495 -7 512 10
rect 552 -7 569 10
<< pdiffc >>
rect 684 55 702 72
rect 743 55 760 72
rect 735 -7 752 10
rect 793 -7 810 10
<< mvndiffc >>
rect 386 58 404 75
rect 466 58 484 75
rect 313 -10 331 7
rect 395 -12 413 5
<< psubdiff >>
rect 491 72 533 77
rect 491 55 503 72
rect 520 55 533 72
rect 491 51 533 55
<< nsubdiff >>
rect 773 72 818 77
rect 773 55 785 72
rect 802 55 818 72
rect 773 51 818 55
<< psubdiffcont >>
rect 503 55 520 72
<< nsubdiffcont >>
rect 785 55 802 72
<< poly >>
rect 410 85 595 100
rect 340 77 368 85
rect 410 83 460 85
rect 340 65 345 77
rect 302 60 345 65
rect 363 60 368 77
rect 302 50 368 60
rect 567 77 595 85
rect 709 77 737 93
rect 302 33 317 50
rect 410 37 460 50
rect 567 42 595 51
rect 709 42 737 51
rect 287 18 317 33
rect 287 -10 303 18
rect 338 15 389 29
rect 278 -25 303 -10
rect 518 14 546 33
rect 567 32 737 42
rect 567 27 642 32
rect 634 15 642 27
rect 659 27 737 32
rect 659 15 667 27
rect 434 -1 461 14
rect 338 -19 389 -17
rect 434 -18 439 -1
rect 456 -18 461 -1
rect 634 9 667 15
rect 758 14 786 31
rect 843 -6 881 4
rect 434 -19 461 -18
rect 338 -34 461 -19
rect 518 -19 546 -11
rect 758 -19 786 -11
rect 843 -19 853 -6
rect 518 -23 853 -19
rect 870 -23 881 -6
rect 518 -34 881 -23
<< polycont >>
rect 345 60 363 77
rect 642 15 659 32
rect 439 -18 456 -1
rect 853 -23 870 -6
<< locali >>
rect 345 77 363 85
rect 635 80 670 82
rect 363 75 409 77
rect 363 60 386 75
rect 345 58 386 60
rect 404 58 413 75
rect 458 58 466 75
rect 484 72 504 75
rect 635 72 641 80
rect 484 58 503 72
rect 345 52 363 58
rect 487 55 503 58
rect 520 55 544 72
rect 561 55 569 72
rect 593 55 601 72
rect 618 59 641 72
rect 662 72 670 80
rect 662 59 684 72
rect 618 55 684 59
rect 702 55 710 72
rect 735 55 743 72
rect 760 55 785 72
rect 802 55 811 72
rect 487 41 513 55
rect 395 24 513 41
rect 788 54 811 55
rect 788 39 815 54
rect 278 -10 313 7
rect 331 -10 340 7
rect 395 5 413 24
rect 487 10 513 24
rect 634 32 667 36
rect 634 15 642 32
rect 659 15 667 32
rect 634 10 667 15
rect 788 22 792 39
rect 809 22 815 39
rect 788 10 815 22
rect 395 -20 413 -12
rect 437 -1 458 7
rect 437 -18 439 -1
rect 456 -18 458 -1
rect 487 -7 495 10
rect 512 -7 520 10
rect 544 -7 552 10
rect 569 -7 735 10
rect 752 -7 760 10
rect 785 -7 793 10
rect 810 -7 818 10
rect 853 -4 870 2
rect 487 -12 504 -7
rect 785 -8 818 -7
rect 437 -26 458 -18
rect 853 -31 870 -26
<< viali >>
rect 641 59 662 80
rect 792 22 809 39
rect 851 -6 873 -4
rect 851 -23 853 -6
rect 853 -23 870 -6
rect 870 -23 873 -6
rect 851 -26 873 -23
<< metal1 >>
rect 434 10 462 13
rect 434 -16 435 10
rect 461 -16 462 10
rect 434 -20 462 -16
rect 487 -40 518 119
rect 635 82 670 84
rect 635 56 639 82
rect 665 56 670 82
rect 635 55 670 56
rect 650 53 670 55
rect 788 39 812 119
rect 788 22 792 39
rect 809 22 812 39
rect 788 -40 812 22
rect 845 -2 886 2
rect 845 -28 849 -2
rect 875 -28 886 -2
rect 845 -31 886 -28
<< via1 >>
rect 435 -16 461 10
rect 639 80 665 82
rect 639 59 641 80
rect 641 59 662 80
rect 662 59 665 80
rect 639 56 665 59
rect 849 -4 875 -2
rect 849 -26 851 -4
rect 851 -26 873 -4
rect 873 -26 875 -4
rect 849 -28 875 -26
<< metal2 >>
rect 639 82 665 85
rect 431 10 465 11
rect 431 -16 435 10
rect 461 5 465 10
rect 639 5 665 56
rect 461 -16 675 5
rect 431 -17 675 -16
rect 846 -2 892 1
rect 846 -28 849 -2
rect 875 -28 892 -2
rect 846 -31 892 -28
<< labels >>
rlabel metal2 885 -31 892 1 0 Input
rlabel metal1 788 115 812 119 0 Vdd
rlabel metal1 788 -40 812 -36 0 Vdd
rlabel metal1 487 115 518 119 0 GND
rlabel metal1 487 -40 518 -35 0 GND
<< end >>
