magic
tech sky130A
magscale 1 2
timestamp 1627063299
<< error_s >>
rect 1062 1286 1120 1342
rect 1220 1286 1278 1342
rect 1378 1286 1436 1342
rect 1018 1272 1478 1286
rect 1018 1242 1032 1272
rect 1062 1260 1120 1272
rect 1220 1260 1278 1272
rect 1378 1260 1436 1272
rect 1062 1242 1063 1243
rect 1119 1242 1120 1243
rect 1220 1242 1221 1243
rect 1277 1242 1278 1243
rect 1378 1242 1379 1243
rect 1435 1242 1436 1243
rect 1464 1242 1478 1272
rect 962 1184 1044 1242
rect 1061 1241 1121 1242
rect 1219 1241 1279 1242
rect 1377 1241 1437 1242
rect 1062 1185 1120 1241
rect 1061 1184 1121 1185
rect 1018 1084 1032 1184
rect 1062 1183 1063 1184
rect 1119 1183 1120 1184
rect 1150 1182 1184 1186
rect 1220 1185 1278 1241
rect 1378 1185 1436 1241
rect 1219 1184 1279 1185
rect 1377 1184 1437 1185
rect 1452 1184 1536 1242
rect 1638 1204 1738 1226
rect 1782 1204 1882 1226
rect 1220 1183 1221 1184
rect 1277 1183 1278 1184
rect 1378 1183 1379 1184
rect 1435 1183 1436 1184
rect 1150 1144 1184 1148
rect 1464 1128 1478 1184
rect 1574 1142 1638 1143
rect 1638 1120 1738 1142
rect 1782 1120 1882 1142
rect 1150 1114 1184 1118
rect 1062 1084 1063 1085
rect 1119 1084 1120 1085
rect 1220 1084 1221 1085
rect 1277 1084 1278 1085
rect 1378 1084 1379 1085
rect 1435 1084 1436 1085
rect 1464 1084 1478 1096
rect 1504 1094 1506 1096
rect 962 1026 1044 1084
rect 1061 1083 1121 1084
rect 1219 1083 1279 1084
rect 1377 1083 1437 1084
rect 1062 1027 1120 1083
rect 1150 1076 1184 1080
rect 1220 1027 1278 1083
rect 1378 1027 1436 1083
rect 1061 1026 1121 1027
rect 1219 1026 1279 1027
rect 1377 1026 1437 1027
rect 1452 1026 1536 1084
rect 1638 1080 1738 1104
rect 1580 1079 1638 1080
rect 1018 1008 1032 1026
rect 1062 1025 1063 1026
rect 1119 1025 1120 1026
rect 1220 1025 1221 1026
rect 1277 1025 1278 1026
rect 1378 1025 1379 1026
rect 1435 1025 1436 1026
rect 1044 1008 1452 1014
rect 1464 1008 1478 1026
rect 1793 1020 1800 1080
rect 1018 982 1478 1008
rect 1638 996 1738 1020
rect 1062 980 1120 982
rect 1220 980 1278 982
rect 1378 980 1436 982
rect 1018 966 1478 980
rect 1018 936 1032 966
rect 1062 954 1120 966
rect 1220 954 1278 966
rect 1378 954 1436 966
rect 1140 938 1192 950
rect 1062 936 1063 937
rect 1119 936 1120 937
rect 1220 936 1221 937
rect 1277 936 1278 937
rect 1378 936 1379 937
rect 1435 936 1436 937
rect 1464 936 1478 966
rect 962 878 1044 936
rect 1061 935 1121 936
rect 1219 935 1279 936
rect 1377 935 1437 936
rect 1062 879 1120 935
rect 1142 910 1194 922
rect 1061 878 1121 879
rect 1018 778 1032 878
rect 1062 877 1063 878
rect 1119 877 1120 878
rect 1150 876 1184 880
rect 1220 879 1278 935
rect 1378 879 1436 935
rect 1219 878 1279 879
rect 1377 878 1437 879
rect 1452 878 1536 936
rect 1638 916 1738 940
rect 1220 877 1221 878
rect 1277 877 1278 878
rect 1378 877 1379 878
rect 1435 877 1436 878
rect 1464 842 1478 878
rect 1580 856 1638 857
rect 1793 856 1800 916
rect 1150 838 1184 842
rect 1638 832 1738 856
rect 1150 808 1184 812
rect 1062 778 1063 779
rect 1119 778 1120 779
rect 1220 778 1221 779
rect 1277 778 1278 779
rect 1378 778 1379 779
rect 1435 778 1436 779
rect 1464 778 1478 808
rect 1494 792 1520 800
rect 1522 792 1548 802
rect 1638 794 1738 816
rect 1782 794 1882 816
rect 1574 793 1638 794
rect 1494 786 1548 792
rect 962 720 1044 778
rect 1061 777 1121 778
rect 1219 777 1279 778
rect 1377 777 1437 778
rect 1062 721 1120 777
rect 1150 770 1184 774
rect 1220 721 1278 777
rect 1378 721 1436 777
rect 1061 720 1121 721
rect 1219 720 1279 721
rect 1377 720 1437 721
rect 1452 720 1536 778
rect 1018 696 1032 720
rect 1062 719 1063 720
rect 1119 719 1120 720
rect 1220 719 1221 720
rect 1277 719 1278 720
rect 1378 719 1379 720
rect 1435 719 1436 720
rect 1060 696 1120 702
rect 1218 696 1278 702
rect 1376 696 1436 702
rect 1464 696 1478 720
rect 1638 710 1738 732
rect 1782 710 1882 732
rect 1018 676 1478 696
rect 1060 668 1120 676
rect 1218 668 1278 676
rect 1376 668 1436 676
rect 1016 654 1476 668
rect 1016 624 1030 654
rect 1060 642 1120 654
rect 1218 642 1278 654
rect 1376 642 1436 654
rect 1140 632 1192 638
rect 1060 624 1061 625
rect 1117 624 1118 625
rect 1218 624 1219 625
rect 1275 624 1276 625
rect 1376 624 1377 625
rect 1433 624 1434 625
rect 1462 624 1476 654
rect 960 566 1042 624
rect 1059 623 1119 624
rect 1217 623 1277 624
rect 1375 623 1435 624
rect 1060 567 1118 623
rect 1140 604 1192 610
rect 1059 566 1119 567
rect 1016 466 1030 566
rect 1060 565 1061 566
rect 1117 565 1118 566
rect 1148 564 1182 568
rect 1218 567 1276 623
rect 1376 567 1434 623
rect 1217 566 1277 567
rect 1375 566 1435 567
rect 1450 566 1534 624
rect 1638 602 1738 624
rect 1782 602 1882 624
rect 1218 565 1219 566
rect 1275 565 1276 566
rect 1376 565 1377 566
rect 1433 565 1434 566
rect 1148 526 1182 530
rect 1462 526 1476 566
rect 1574 540 1638 541
rect 1638 518 1738 540
rect 1782 518 1882 540
rect 1148 496 1182 500
rect 1060 466 1061 467
rect 1117 466 1118 467
rect 1218 466 1219 467
rect 1275 466 1276 467
rect 1376 466 1377 467
rect 1433 466 1434 467
rect 1462 466 1476 492
rect 1638 478 1738 502
rect 1580 477 1638 478
rect 960 408 1042 466
rect 1059 465 1119 466
rect 1217 465 1277 466
rect 1375 465 1435 466
rect 1060 409 1118 465
rect 1148 458 1182 462
rect 1218 409 1276 465
rect 1376 409 1434 465
rect 1059 408 1119 409
rect 1217 408 1277 409
rect 1375 408 1435 409
rect 1450 408 1534 466
rect 1793 418 1800 478
rect 1016 388 1030 408
rect 1060 407 1061 408
rect 1117 407 1118 408
rect 1218 407 1219 408
rect 1275 407 1276 408
rect 1376 407 1377 408
rect 1433 407 1434 408
rect 1042 390 1450 394
rect 1060 388 1118 390
rect 1218 388 1276 390
rect 1376 388 1434 390
rect 1462 388 1476 408
rect 1638 394 1738 418
rect 1016 364 1476 388
rect 1060 360 1118 364
rect 1218 360 1276 364
rect 1376 360 1434 364
rect 1016 346 1476 360
rect 1016 316 1030 346
rect 1060 334 1118 346
rect 1218 334 1276 346
rect 1376 334 1434 346
rect 1138 320 1190 330
rect 1060 316 1061 317
rect 1117 316 1118 317
rect 1218 316 1219 317
rect 1275 316 1276 317
rect 1376 316 1377 317
rect 1433 316 1434 317
rect 1462 316 1476 346
rect 1638 316 1738 340
rect 960 258 1042 316
rect 1059 315 1119 316
rect 1217 315 1277 316
rect 1375 315 1435 316
rect 1060 259 1118 315
rect 1140 292 1192 302
rect 1059 258 1119 259
rect 1016 158 1030 258
rect 1060 257 1061 258
rect 1117 257 1118 258
rect 1148 256 1182 260
rect 1218 259 1276 315
rect 1376 259 1434 315
rect 1217 258 1277 259
rect 1375 258 1435 259
rect 1450 258 1534 316
rect 1218 257 1219 258
rect 1275 257 1276 258
rect 1376 257 1377 258
rect 1433 257 1434 258
rect 1462 242 1476 258
rect 1580 256 1638 257
rect 1793 256 1800 316
rect 1638 232 1738 256
rect 1148 218 1182 222
rect 1148 188 1182 192
rect 1060 158 1061 159
rect 1117 158 1118 159
rect 1218 158 1219 159
rect 1275 158 1276 159
rect 1376 158 1377 159
rect 1433 158 1434 159
rect 1462 158 1476 208
rect 1638 194 1738 216
rect 1782 194 1882 216
rect 1574 193 1638 194
rect 960 100 1042 158
rect 1059 157 1119 158
rect 1217 157 1277 158
rect 1375 157 1435 158
rect 1060 101 1118 157
rect 1148 150 1182 154
rect 1218 101 1276 157
rect 1376 101 1434 157
rect 1059 100 1119 101
rect 1217 100 1277 101
rect 1375 100 1435 101
rect 1450 100 1534 158
rect 1638 110 1738 132
rect 1782 110 1882 132
rect 1016 70 1030 100
rect 1060 99 1061 100
rect 1117 99 1118 100
rect 1218 99 1219 100
rect 1275 99 1276 100
rect 1376 99 1377 100
rect 1433 99 1434 100
rect 1060 70 1118 82
rect 1218 70 1276 82
rect 1376 70 1434 82
rect 1462 70 1476 100
rect 1016 56 1476 70
rect 1060 0 1118 56
rect 1218 0 1276 56
rect 1376 0 1434 56
<< nwell >>
rect 1792 682 1862 684
rect 1792 650 1826 682
rect 1860 650 1862 682
<< poly >>
rect 1434 1120 1506 1128
rect 314 1054 788 1102
rect 1434 1096 1504 1120
rect 314 836 784 884
rect 1434 808 1504 842
rect 1826 682 1862 684
rect 1858 650 1862 682
rect 314 476 788 524
rect 1168 492 1504 526
rect 318 236 792 284
rect 1168 208 1504 242
<< polycont >>
rect 1792 650 1826 684
<< locali >>
rect 1774 650 1792 684
<< viali >>
rect 1826 650 1862 684
<< metal1 >>
rect 72 62 152 1260
rect 1836 690 1862 694
rect 1820 684 1868 690
rect 1820 650 1826 684
rect 1862 650 1868 684
rect 1820 644 1868 650
rect 1840 636 1862 644
<< metal2 >>
rect 0 1158 1522 1172
rect 0 1136 1528 1158
rect 0 1050 1948 1086
rect 0 874 1522 886
rect 0 850 1528 874
rect 0 786 1520 800
rect 0 764 1528 786
rect 4 534 1528 568
rect 4 450 1528 484
rect 4 254 1528 288
rect 160 236 468 254
rect 4 166 1528 200
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_1
timestamp 1608066871
transform 1 0 2904 0 1 862
box -2902 -800 -2556 -420
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_0
timestamp 1608066871
transform 1 0 2904 0 1 1096
box -2902 -800 -2556 -420
use sky130_hilas_overlapCap01  sky130_hilas_overlapCap01_2
timestamp 1607257541
transform 1 0 1534 0 1 450
box -574 -142 0 274
use sky130_hilas_overlapCap01  sky130_hilas_overlapCap01_3
timestamp 1607257541
transform 1 0 1534 0 1 142
box -574 -142 0 274
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_2
timestamp 1607386385
transform 1 0 2082 0 -1 764
box -578 94 -66 464
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_1
timestamp 1607386385
transform 1 0 2082 0 1 -30
box -578 94 -66 464
use sky130_hilas_wellContact  sky130_hilas_wellContact_1
timestamp 1606753443
transform 1 0 2898 0 1 1412
box -2898 -882 -2550 -510
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_3
timestamp 1608066871
transform 1 0 2904 0 1 1692
box -2902 -800 -2556 -420
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_2
timestamp 1608066871
transform 1 0 2904 0 1 1474
box -2902 -800 -2556 -420
use sky130_hilas_overlapCap01  sky130_hilas_overlapCap01_1
timestamp 1607257541
transform 1 0 1536 0 1 762
box -574 -142 0 274
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_0
timestamp 1607386385
transform 1 0 2082 0 1 570
box -578 94 -66 464
use sky130_hilas_overlapCap01  sky130_hilas_overlapCap01_0
timestamp 1607257541
transform 1 0 1536 0 1 1068
box -574 -142 0 274
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_3
timestamp 1607386385
transform 1 0 2082 0 -1 1366
box -578 94 -66 464
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
