magic
tech sky130A
timestamp 1629420194
<< error_s >>
rect -18 20 21 23
rect -18 -22 21 -19
<< nwell >>
rect -79 -78 82 43
<< pmos >>
rect -18 -19 21 20
<< pdiff >>
rect -45 9 -18 20
rect -45 -8 -41 9
rect -24 -8 -18 9
rect -45 -19 -18 -8
rect 21 9 48 20
rect 21 -8 27 9
rect 44 -8 48 9
rect 21 -19 48 -8
<< pdiffc >>
rect -41 -8 -24 9
rect 27 -8 44 9
<< poly >>
rect -18 20 21 33
rect -18 -27 21 -19
rect -18 -42 72 -27
rect 56 -59 72 -42
rect 56 -70 73 -59
rect 56 -74 72 -70
rect 58 -76 72 -74
rect 58 -84 64 -76
<< locali >>
rect -41 9 -24 17
rect -41 -16 -24 -8
rect 27 9 44 17
rect 27 -16 44 -8
use sky130_hilas_poly2m1  sky130_hilas_poly2m1_0
timestamp 1629420194
transform 1 0 -85 0 1 7
box -9 -26 24 25
use sky130_hilas_poly2m1  sky130_hilas_poly2m1_2
timestamp 1629420194
transform 1 0 73 0 -1 -77
box -9 -26 24 25
<< end >>
