magic
tech sky130A
timestamp 1629137164
<< metal2 >>
rect 22 54 59 60
rect 22 26 27 54
rect 55 26 59 54
rect 22 20 59 26
<< via2 >>
rect 27 26 55 54
<< metal3 >>
rect 0 63 79 75
rect 0 15 19 63
rect 62 15 79 63
rect 0 0 79 15
<< via3 >>
rect 19 54 62 63
rect 19 26 27 54
rect 27 26 55 54
rect 55 26 62 54
rect 19 15 62 26
<< metal4 >>
rect 9 63 75 72
rect 9 15 19 63
rect 62 15 75 63
rect 9 6 75 15
<< end >>
