magic
tech sky130A
timestamp 1628707349
<< checkpaint >>
rect -548 1121 1020 1234
rect -630 -517 1020 1121
rect -548 -630 1020 -517
<< nwell >>
rect 390 156 471 448
<< psubdiff >>
rect 397 562 441 586
rect 397 545 410 562
rect 427 545 441 562
rect 397 528 441 545
rect 397 511 410 528
rect 427 511 441 528
rect 397 494 441 511
rect 397 477 410 494
rect 427 477 441 494
rect 397 468 441 477
rect 398 104 441 130
rect 398 87 411 104
rect 428 87 441 104
rect 398 70 441 87
rect 398 53 411 70
rect 428 53 441 70
rect 398 36 441 53
rect 398 19 411 36
rect 428 19 441 36
rect 398 14 441 19
<< nsubdiff >>
rect 398 405 440 417
rect 398 387 409 405
rect 427 387 440 405
rect 398 368 440 387
rect 398 350 409 368
rect 427 350 440 368
rect 398 332 440 350
rect 398 314 409 332
rect 427 314 440 332
rect 398 296 440 314
rect 398 278 409 296
rect 427 278 440 296
rect 398 261 440 278
rect 398 243 410 261
rect 428 243 440 261
rect 398 225 440 243
rect 398 207 410 225
rect 428 207 440 225
rect 398 198 440 207
<< psubdiffcont >>
rect 410 545 427 562
rect 410 511 427 528
rect 410 477 427 494
rect 411 87 428 104
rect 411 53 428 70
rect 411 19 428 36
<< nsubdiffcont >>
rect 409 387 427 405
rect 409 350 427 368
rect 409 314 427 332
rect 409 278 427 296
rect 410 243 428 261
rect 410 207 428 225
<< locali >>
rect 373 562 435 579
rect 373 545 410 562
rect 427 545 435 562
rect 373 528 435 545
rect 373 511 410 528
rect 427 511 435 528
rect 373 494 435 511
rect 373 490 410 494
rect 399 477 410 490
rect 427 477 435 494
rect 399 475 435 477
rect 371 405 429 413
rect 371 387 409 405
rect 427 387 429 405
rect 371 374 429 387
rect 371 368 434 374
rect 371 350 409 368
rect 427 350 434 368
rect 371 332 434 350
rect 371 328 409 332
rect 371 311 374 328
rect 391 311 408 328
rect 427 314 434 332
rect 425 311 434 314
rect 371 296 434 311
rect 371 293 409 296
rect 371 276 374 293
rect 391 276 408 293
rect 427 278 434 296
rect 425 276 434 278
rect 371 261 434 276
rect 371 243 410 261
rect 428 243 434 261
rect 371 236 434 243
rect 371 225 429 236
rect 371 207 410 225
rect 428 207 429 225
rect 371 199 429 207
rect 373 104 428 114
rect 373 87 411 104
rect 373 70 428 87
rect 373 53 411 70
rect 373 36 428 53
rect 373 25 411 36
rect 411 11 428 19
<< viali >>
rect 374 311 391 328
rect 408 314 409 328
rect 409 314 425 328
rect 408 311 425 314
rect 374 276 391 293
rect 408 278 409 293
rect 409 278 425 293
rect 408 276 425 278
<< metal1 >>
rect 82 541 103 604
rect 82 525 330 541
rect 364 550 471 604
rect 364 541 383 550
rect 356 525 383 541
rect 82 524 383 525
rect 409 524 471 550
rect 82 510 471 524
rect 82 509 383 510
rect 82 483 328 509
rect 354 484 383 509
rect 409 484 471 510
rect 354 483 471 484
rect 82 473 471 483
rect 82 419 471 442
rect 82 392 119 419
rect 146 392 174 419
rect 201 392 471 419
rect 82 362 471 392
rect 82 361 174 362
rect 82 334 118 361
rect 145 335 174 361
rect 201 335 471 362
rect 145 334 471 335
rect 82 328 471 334
rect 82 311 374 328
rect 391 311 408 328
rect 425 311 471 328
rect 82 293 471 311
rect 82 278 374 293
rect 82 277 174 278
rect 82 258 119 277
rect 82 257 99 258
rect 82 250 119 257
rect 146 258 174 277
rect 146 251 174 257
rect 201 276 374 278
rect 391 276 408 293
rect 425 276 471 293
rect 201 258 471 276
rect 334 257 471 258
rect 201 251 471 257
rect 146 250 471 251
rect 82 227 471 250
rect 82 200 119 227
rect 146 225 471 227
rect 146 200 172 225
rect 82 198 172 200
rect 199 198 471 225
rect 82 163 471 198
rect 82 100 471 127
rect 82 74 344 100
rect 370 74 392 100
rect 418 74 471 100
rect 82 59 471 74
rect 82 33 342 59
rect 368 33 391 59
rect 417 33 471 59
rect 82 3 471 33
rect 82 0 99 3
rect 373 1 471 3
rect 372 0 471 1
<< via1 >>
rect 330 525 356 551
rect 383 524 409 550
rect 328 483 354 509
rect 383 484 409 510
rect 119 392 146 419
rect 174 392 201 419
rect 118 334 145 361
rect 174 335 201 362
rect 119 250 146 277
rect 174 251 201 278
rect 119 200 146 227
rect 172 198 199 225
rect 344 74 370 100
rect 392 74 418 100
rect 342 33 368 59
rect 391 33 417 59
<< metal2 >>
rect 104 419 234 604
rect 104 392 119 419
rect 146 392 174 419
rect 201 392 234 419
rect 104 362 234 392
rect 104 361 174 362
rect 104 334 118 361
rect 145 335 174 361
rect 201 335 234 362
rect 145 334 234 335
rect 104 278 234 334
rect 104 277 174 278
rect 104 250 119 277
rect 146 251 174 277
rect 201 251 234 278
rect 146 250 234 251
rect 104 227 234 250
rect 104 200 119 227
rect 146 225 234 227
rect 146 200 172 225
rect 104 198 172 200
rect 199 198 234 225
rect 104 0 234 198
rect 312 551 442 604
rect 312 525 330 551
rect 356 550 442 551
rect 356 525 383 550
rect 312 524 383 525
rect 409 524 442 550
rect 312 510 442 524
rect 312 509 383 510
rect 312 483 328 509
rect 354 484 383 509
rect 409 484 442 510
rect 354 483 442 484
rect 312 100 442 483
rect 312 74 344 100
rect 370 74 392 100
rect 418 74 442 100
rect 312 59 442 74
rect 312 33 342 59
rect 368 33 391 59
rect 417 33 442 59
rect 312 0 442 33
use sky130_hilas_decoup_cap_00  CapDeco_0
timestamp 1628705748
transform 1 0 0 0 -1 491
box 0 0 308 307
use sky130_hilas_decoup_cap_00  CapDeco_1
timestamp 1628705748
transform 1 0 0 0 1 113
box 0 0 308 307
<< labels >>
rlabel metal1 82 254 99 350 0 VPWR
port 1 nsew
rlabel metal1 454 256 471 350 0 VPWR
port 1 nsew
rlabel metal1 461 541 471 604 0 VGND
port 1 nsew
rlabel metal1 82 541 90 604 0 VGND
port 1 nsew
rlabel metal1 82 0 91 63 0 VGND
port 1 nsew
rlabel metal1 456 0 471 63 0 VGND
port 1 nsew
rlabel metal2 104 594 234 604 0 VPWR
port 1 nsew
rlabel metal2 312 596 442 604 0 VGND
port 2 nsew
rlabel metal2 104 0 234 12 0 VPWR
port 1 nsew
rlabel metal2 312 0 442 12 0 VGND
port 2 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
