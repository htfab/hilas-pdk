magic
tech sky130A
timestamp 1623107852
use sky130_hilas_decoup_cap_00  CapDeco_1
timestamp 1623107852
transform 1 0 273 0 1 170
box 82 -113 390 189
use sky130_hilas_decoup_cap_00  CapDeco_0
timestamp 1623107852
transform 1 0 273 0 -1 548
box 82 -113 390 189
<< end >>
