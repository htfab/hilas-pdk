* Copyright 2020 The Hilas PDK Authors
* 
* This file is part of HILAS.
* 
* HILAS is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published by
* the Free Software Foundation, version 3 of the License.
* 
* HILAS is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
* 
* You should have received a copy of the GNU Lesser General Public License
* along with HILAS.  If not, see <https://www.gnu.org/licenses/>.
* 
* Licensed under the Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
* https://www.gnu.org/licenses/lgpl-3.0.en.html
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
* SPDX-License-Identifier: LGPL-3.0
* 
* 

* NGSPICE file created from sky130_hilas_WTA4stage01.ext - technology: sky130A

.subckt sky130_hilas_WTAsinglestage01 a_4_n68# sky130_hilas_li2m2_1/SUB
X0 sky130_hilas_li2m2_1/SUB a_4_n68# a_n126_n150# sky130_hilas_li2m2_1/SUB sky130_fd_pr__nfet_01v8 w=590000u l=200000u
X1 a_4_n68# a_n126_n150# a_n94_n68# sky130_hilas_li2m2_1/SUB sky130_fd_pr__nfet_01v8 w=590000u l=200000u
.ends


* Top level circuit sky130_hilas_WTA4stage01

Xsky130_hilas_WTAsinglestage01_0 a_284_2# SUB sky130_hilas_WTAsinglestage01
Xsky130_hilas_WTAsinglestage01_1 a_284_2# SUB sky130_hilas_WTAsinglestage01
Xsky130_hilas_WTAsinglestage01_2 a_284_2# SUB sky130_hilas_WTAsinglestage01
Xsky130_hilas_WTAsinglestage01_3 a_284_2# SUB sky130_hilas_WTAsinglestage01
.end

