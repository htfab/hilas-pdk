magic
tech sky130A
timestamp 1634057707
<< poly >>
rect 0 25 27 33
rect 0 8 5 25
rect 22 8 27 25
rect 0 0 27 8
<< polycont >>
rect 5 8 22 25
<< locali >>
rect 5 25 22 33
rect 5 0 22 8
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
