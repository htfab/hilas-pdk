magic
tech sky130A
timestamp 1628707275
<< poly >>
rect 0 43 33 51
rect 0 26 8 43
rect 25 26 33 43
rect 0 18 33 26
<< polycont >>
rect 8 26 25 43
<< locali >>
rect 6 43 27 51
rect 6 26 8 43
rect 25 26 27 43
rect 6 23 27 26
rect 6 8 8 23
rect 25 8 27 23
<< viali >>
rect 8 6 25 23
<< metal1 >>
rect 6 29 28 51
rect 5 23 28 29
rect 5 6 8 23
rect 25 6 28 23
rect 5 0 28 6
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
