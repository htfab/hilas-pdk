magic
tech sky130A
timestamp 1628707342
<< nwell >>
rect 0 0 223 185
<< mvvaractor >>
rect 56 59 167 123
<< mvnsubdiff >>
rect 56 123 167 151
rect 56 34 167 59
<< poly >>
rect 16 59 56 123
rect 167 59 208 123
<< metal1 >>
rect 65 0 103 186
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
