magic
tech sky130A
timestamp 1629137213
<< checkpaint >>
rect -470 -628 823 683
<< nwell >>
rect 0 12 161 133
<< pmos >>
rect 61 71 100 110
<< pdiff >>
rect 34 71 61 110
rect 100 71 127 110
<< poly >>
rect 61 110 100 123
rect 61 63 100 71
rect 61 48 150 63
rect 135 27 150 48
rect 135 12 187 27
rect 159 11 164 12
rect 172 0 187 12
use sky130_hilas_poly2m1  sky130_hilas_poly2m1_0
timestamp 1629137133
transform 1 0 160 0 1 2
box 0 0 33 51
<< end >>
