magic
tech sky130A
timestamp 1634057829
<< checkpaint >>
rect -366 -248 2918 2102
rect 368 -434 1816 -248
rect 477 -521 1816 -434
<< error_s >>
rect 432 542 438 548
rect 537 542 543 548
rect 58 532 64 538
rect 111 532 117 538
rect 52 482 58 488
rect 117 482 123 488
rect 426 478 432 484
rect 543 478 549 484
rect 58 423 64 429
rect 111 423 117 429
rect 432 425 438 431
rect 537 425 543 431
rect 52 373 58 379
rect 117 373 123 379
rect 426 361 432 367
rect 543 361 549 367
rect 3635 285 3637 313
rect 432 240 438 246
rect 537 240 543 246
rect 58 234 64 240
rect 111 234 117 240
rect 52 184 58 190
rect 117 184 123 190
rect 426 176 432 182
rect 543 176 549 182
rect 432 124 438 130
rect 537 124 543 130
rect 58 117 64 123
rect 111 117 117 123
rect 52 67 58 73
rect 117 67 123 73
rect 426 60 432 66
rect 543 60 549 66
<< nwell >>
rect 1007 604 3542 605
rect 1008 597 3542 604
rect 1 537 12 555
rect 0 351 12 369
rect 2 52 12 69
rect 1006 6 3542 597
rect 1007 1 3542 6
rect 1200 0 3542 1
<< metal1 >>
rect 36 591 76 605
rect 280 599 304 605
rect 442 597 479 605
rect 673 598 697 605
rect 912 600 931 605
rect 956 600 972 605
rect 441 592 479 597
rect 440 13 441 15
rect 36 0 75 12
rect 280 0 304 7
rect 440 1 479 13
rect 440 0 441 1
rect 673 0 697 7
rect 875 1 891 7
rect 912 1 931 7
rect 956 1 972 7
<< metal2 >>
rect 1074 602 1125 605
rect 1074 600 1167 602
rect 1074 593 1130 600
rect 888 574 1130 593
rect 1117 572 1130 574
rect 1158 572 1167 600
rect 1 537 12 555
rect 898 537 3670 555
rect 892 494 3670 512
rect 898 394 3670 412
rect 3569 369 3670 370
rect 0 351 12 369
rect 894 351 3670 369
rect 3601 313 3670 320
rect 3601 285 3608 313
rect 3637 285 3670 313
rect 3601 279 3670 285
rect 2 236 12 253
rect 877 236 3670 253
rect 887 194 3670 211
rect 885 96 3670 113
rect 2 52 12 69
rect 881 52 3670 69
<< via2 >>
rect 1130 572 1158 600
rect 3608 285 3637 313
<< metal3 >>
rect 1125 600 1163 603
rect 1125 574 1130 600
rect 1117 572 1130 574
rect 1158 574 1163 600
rect 1158 572 1171 574
rect 1117 449 1171 572
rect 3523 313 3638 384
rect 3523 285 3608 313
rect 3637 285 3638 313
rect 1037 200 1055 230
rect 3523 220 3638 285
rect 3568 219 3638 220
rect 1146 79 1164 109
<< metal4 >>
rect 1279 538 1689 568
rect 1110 477 1380 488
rect 1110 447 1401 477
rect 1350 413 1401 447
rect 1651 418 1689 538
rect 1935 421 2263 451
rect 1041 375 1177 405
rect 1147 319 1177 375
rect 1935 319 1965 421
rect 2233 319 2263 421
rect 1147 289 2263 319
rect 2503 419 3392 449
rect 1371 230 1690 233
rect 1935 230 1965 233
rect 1037 200 2257 230
rect 1371 163 1401 200
rect 1660 166 1690 200
rect 1935 166 1965 200
rect 1660 163 1965 166
rect 2227 163 2257 200
rect 1371 133 2257 163
rect 2503 167 2533 419
rect 2786 416 3097 419
rect 2786 167 2816 416
rect 3067 167 3097 416
rect 3362 167 3392 419
rect 2503 137 3398 167
rect 3067 136 3398 137
rect 1134 79 1185 109
rect 1155 55 1185 79
rect 3368 55 3398 136
rect 1155 25 3398 55
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_1
timestamp 1634057717
transform 1 0 264 0 1 382
box 0 0 2024 1090
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_0
timestamp 1634057717
transform 1 0 264 0 1 382
box 0 0 2024 1090
use sky130_hilas_m22m4  sky130_hilas_m22m4_1
timestamp 1634057755
transform 1 0 1002 0 1 405
box 0 0 79 75
use sky130_hilas_m22m4  sky130_hilas_m22m4_2
timestamp 1634057755
transform 1 0 998 0 1 196
box 0 0 79 75
use sky130_hilas_m22m4  sky130_hilas_m22m4_3
timestamp 1634057755
transform 1 0 1107 0 1 109
box 0 0 79 75
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1634057711
transform 1 0 876 0 1 581
box 0 0 32 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1634057711
transform 1 0 876 0 1 581
box 0 0 32 32
<< labels >>
rlabel metal2 3658 279 3670 320 0 CAPTERM2
port 1 nsew analog default
rlabel metal2 1074 592 1125 605 0 CAPTERM1
port 2 nsew analog default
rlabel metal1 912 600 931 605 0 GATESELECT
port 4 nsew
rlabel metal1 956 600 972 605 0 VINJ
port 3 nsew power default
rlabel metal1 442 592 479 605 0 GATE
port 6 nsew analog default
rlabel metal1 36 591 76 605 0 VTUN
port 5 nsew
rlabel metal1 36 0 75 12 0 VTUN
port 5 nsew
rlabel metal1 440 1 479 13 0 GATE
port 6 nsew
rlabel metal1 956 1 972 7 0 VINJ
rlabel metal1 875 1 891 7 0 CAPTERM1
rlabel metal1 912 1 931 7 0 GATESELECT
rlabel metal2 1 537 12 555 0 DRAIN1
port 8 nsew
rlabel metal2 0 351 12 369 0 DRAIN2
port 7 nsew
rlabel metal2 3660 52 3670 69 0 DRAIN4
port 10 nsew
rlabel metal2 3660 537 3670 555 0 DRAIN1
port 8 nsew
rlabel metal2 3659 351 3670 370 0 DRAIN2
port 7 nsew
rlabel metal2 3659 236 3670 253 0 DRAIN3
port 11 nsew
rlabel metal2 2 236 12 253 0 DRAIN3
port 11 nsew
rlabel metal2 2 52 12 69 0 DRAIN4
port 10 nsew
rlabel metal1 280 599 304 605 0 VGND
port 12 nsew
rlabel metal1 673 598 697 605 0 VGND
port 12 nsew
rlabel metal1 280 0 304 7 0 VGND
port 12 nsew
rlabel metal1 673 0 697 7 0 VGND
port 12 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
