magic
tech sky130A
timestamp 1637804567
<< error_s >>
rect 1412 612 1462 617
rect 1592 612 1642 618
rect 766 583 818 591
rect 818 578 846 583
rect 1120 579 1170 589
rect 1706 582 1707 599
rect 1089 578 1120 579
rect 1412 570 1462 575
rect 1592 570 1642 576
rect 766 541 818 549
rect 1120 537 1170 547
rect 1412 545 1462 551
rect 1732 545 1782 551
rect 692 518 745 527
rect 839 518 891 528
rect 665 512 692 518
rect 891 513 918 518
rect 1049 517 1099 528
rect 1191 517 1241 528
rect 1020 513 1049 517
rect 665 493 668 512
rect 1412 503 1462 509
rect 1732 503 1782 509
rect 692 476 745 485
rect 839 476 891 486
rect 1049 475 1099 486
rect 1191 475 1241 486
rect 1412 442 1462 448
rect 1732 442 1782 448
rect 766 432 818 440
rect 818 427 846 432
rect 1120 428 1170 438
rect 1089 427 1120 428
rect 1412 400 1462 406
rect 1732 400 1782 406
rect 766 390 818 398
rect 1120 386 1170 396
rect 692 367 745 376
rect 839 367 891 377
rect 665 361 692 367
rect 891 362 918 367
rect 1049 366 1099 377
rect 1191 366 1241 377
rect 1412 376 1462 381
rect 1592 375 1642 381
rect 1020 362 1049 366
rect 665 342 668 361
rect 1706 352 1707 369
rect 692 325 745 334
rect 839 325 891 335
rect 1049 324 1099 335
rect 1191 324 1241 335
rect 1412 334 1462 339
rect 1592 333 1642 339
rect 1412 292 1462 297
rect 1592 292 1642 298
rect 766 281 818 289
rect 818 276 846 281
rect 1120 277 1170 287
rect 1089 276 1120 277
rect 1706 262 1707 279
rect 1412 250 1462 255
rect 1592 250 1642 256
rect 766 239 818 247
rect 1120 235 1170 245
rect 692 216 745 225
rect 839 216 891 226
rect 665 210 692 216
rect 891 211 918 216
rect 1049 215 1099 226
rect 1191 215 1241 226
rect 1412 225 1462 231
rect 1732 225 1782 231
rect 1020 211 1049 215
rect 665 191 668 210
rect 692 174 745 183
rect 839 174 891 184
rect 1049 173 1099 184
rect 1191 173 1241 184
rect 1412 183 1462 189
rect 1732 183 1782 189
rect 839 171 891 172
rect 1049 171 1099 172
rect 766 131 818 139
rect 818 126 846 131
rect 1120 127 1170 137
rect 1089 126 1120 127
rect 1412 122 1462 128
rect 1732 122 1782 128
rect 766 89 818 97
rect 1120 85 1170 95
rect 1412 80 1462 86
rect 1732 80 1782 86
rect 692 66 745 75
rect 839 66 891 76
rect 665 60 692 66
rect 891 61 918 66
rect 1049 65 1099 76
rect 1191 65 1241 76
rect 1020 61 1049 65
rect 665 41 668 60
rect 1412 56 1462 61
rect 1592 55 1642 61
rect 692 24 745 33
rect 839 24 891 34
rect 1049 23 1099 34
rect 1191 23 1241 34
rect 1706 32 1707 49
rect 1412 14 1462 19
rect 1592 13 1642 19
<< psubdiff >>
rect 3042 604 3093 621
rect 3042 11 3058 604
rect 3075 11 3093 604
rect 3042 0 3093 11
<< psubdiffcont >>
rect 3058 11 3075 604
<< poly >>
rect 1921 592 1959 600
rect 1921 575 1931 592
rect 1948 575 1959 592
rect 1921 567 1959 575
rect 2978 592 3012 600
rect 2978 575 2988 592
rect 3005 575 3012 592
rect 2978 567 3012 575
rect 1921 516 1959 525
rect 1921 499 1930 516
rect 1947 499 1959 516
rect 1921 492 1959 499
rect 2978 517 3012 525
rect 2978 500 2988 517
rect 3005 500 3012 517
rect 2978 492 3012 500
rect 1921 421 1959 429
rect 1921 404 1930 421
rect 1947 404 1959 421
rect 1921 396 1959 404
rect 2978 421 3012 429
rect 2978 404 2987 421
rect 3004 404 3012 421
rect 2978 396 3012 404
rect 1921 349 1959 357
rect 1921 332 1930 349
rect 1947 332 1959 349
rect 1921 324 1959 332
rect 2978 348 3012 357
rect 2978 331 2987 348
rect 3004 331 3012 348
rect 2978 324 3012 331
rect 1921 259 1959 268
rect 1921 242 1931 259
rect 1948 242 1959 259
rect 1921 235 1959 242
rect 2978 260 3012 268
rect 2978 243 2986 260
rect 3003 243 3012 260
rect 2978 235 3012 243
rect 1921 186 1959 194
rect 1921 169 1931 186
rect 1948 169 1959 186
rect 1921 161 1959 169
rect 2978 186 3012 194
rect 2978 169 2986 186
rect 3003 169 3012 186
rect 2978 161 3012 169
rect 1921 102 1959 110
rect 1921 85 1930 102
rect 1947 85 1959 102
rect 1921 77 1959 85
rect 2978 102 3012 110
rect 2978 85 2987 102
rect 3004 85 3012 102
rect 2978 77 3012 85
rect 1921 36 1959 44
rect 1921 19 1930 36
rect 1947 19 1959 36
rect 1921 11 1959 19
rect 2978 35 3012 44
rect 2978 18 2987 35
rect 3004 18 3012 35
rect 2978 11 3012 18
<< polycont >>
rect 1931 575 1948 592
rect 2988 575 3005 592
rect 1930 499 1947 516
rect 2988 500 3005 517
rect 1930 404 1947 421
rect 2987 404 3004 421
rect 1930 332 1947 349
rect 2987 331 3004 348
rect 1931 242 1948 259
rect 2986 243 3003 260
rect 1931 169 1948 186
rect 2986 169 3003 186
rect 1930 85 1947 102
rect 2987 85 3004 102
rect 1930 19 1947 36
rect 2987 18 3004 35
<< npolyres >>
rect 1959 567 2978 600
rect 1959 492 2978 525
rect 1959 396 2978 429
rect 1959 324 2978 357
rect 1959 235 2978 268
rect 1959 161 2978 194
rect 1959 77 2978 110
rect 1959 11 2978 44
<< locali >>
rect 1927 592 1950 600
rect 1927 575 1931 592
rect 1948 575 1950 592
rect 1927 555 1950 575
rect 2988 592 3005 645
rect 2988 566 3005 575
rect 3043 605 3075 612
rect 1927 538 1930 555
rect 1947 538 1950 555
rect 1927 516 1950 538
rect 1927 499 1930 516
rect 1947 499 1950 516
rect 2988 517 3005 526
rect 1927 491 1950 499
rect 2987 500 2988 509
rect 2987 492 3005 500
rect 1926 421 1949 429
rect 1926 404 1930 421
rect 1947 404 1949 421
rect 1926 383 1949 404
rect 2987 421 3004 492
rect 2987 395 3004 404
rect 1926 366 1929 383
rect 1946 366 1949 383
rect 1926 349 1949 366
rect 1926 332 1930 349
rect 1947 332 1949 349
rect 1926 323 1949 332
rect 2987 348 3004 359
rect 2987 323 3004 331
rect 2986 268 3004 323
rect 1928 259 1951 267
rect 1928 242 1931 259
rect 1948 242 1951 259
rect 1928 220 1951 242
rect 2986 260 3003 268
rect 2986 234 3003 243
rect 1928 203 1931 220
rect 1948 203 1951 220
rect 1928 186 1951 203
rect 1928 169 1931 186
rect 1948 169 1951 186
rect 1928 161 1951 169
rect 2986 186 3003 195
rect 3003 169 3004 178
rect 2986 161 3004 169
rect 1925 102 1949 110
rect 1925 85 1930 102
rect 1947 85 1949 102
rect 1925 69 1949 85
rect 2987 102 3004 161
rect 2987 76 3004 85
rect 1925 52 1929 69
rect 1946 52 1949 69
rect 1925 36 1949 52
rect 1925 19 1930 36
rect 1947 19 1949 36
rect 1925 11 1949 19
rect 2987 35 3004 45
rect 2987 -14 3004 18
rect 3043 11 3049 605
rect 3066 604 3075 605
rect 3043 4 3075 11
rect 3058 3 3075 4
<< viali >>
rect 1930 538 1947 555
rect 1929 366 1946 383
rect 1931 203 1948 220
rect 1929 52 1946 69
rect 3049 604 3066 605
rect 3049 11 3058 604
rect 3058 11 3066 604
<< metal1 >>
rect 3042 605 3069 645
rect 1899 561 1953 570
rect 1899 535 1902 561
rect 1928 555 1953 561
rect 1928 538 1930 555
rect 1947 538 1953 555
rect 1928 535 1953 538
rect 1899 527 1953 535
rect 1901 391 1952 399
rect 1901 365 1904 391
rect 1930 383 1952 391
rect 1946 366 1952 383
rect 1930 365 1952 366
rect 1901 356 1952 365
rect 1912 235 1954 240
rect 1899 230 1954 235
rect 1899 204 1902 230
rect 1928 220 1954 230
rect 1928 204 1931 220
rect 1899 203 1931 204
rect 1948 203 1954 220
rect 1899 197 1954 203
rect 1896 69 1949 75
rect 1896 43 1899 69
rect 1925 52 1929 69
rect 1946 52 1949 69
rect 1925 43 1949 52
rect 1896 40 1949 43
rect 1907 32 1949 40
rect 3042 11 3049 605
rect 3066 604 3069 605
rect 3066 11 3075 604
rect 3042 -14 3069 11
<< via1 >>
rect 1902 535 1928 561
rect 1904 383 1930 391
rect 1904 366 1929 383
rect 1929 366 1930 383
rect 1904 365 1930 366
rect 1902 204 1928 230
rect 1899 43 1925 69
<< metal2 >>
rect 1848 585 1932 602
rect 1906 565 1923 585
rect 1900 561 1929 565
rect 1285 531 1306 554
rect 1900 535 1902 561
rect 1928 535 1929 561
rect 1900 532 1929 535
rect 1285 524 1309 531
rect 1285 516 1306 524
rect 1279 500 1306 516
rect 1285 483 1306 500
rect 1289 365 1310 420
rect 1903 391 1931 394
rect 1903 376 1904 391
rect 1279 349 1310 365
rect 1849 365 1904 376
rect 1930 365 1931 391
rect 1849 360 1931 365
rect 1849 358 1926 360
rect 1289 332 1310 349
rect 1851 264 1925 280
rect 1907 234 1923 264
rect 1901 230 1929 234
rect 1279 210 1295 212
rect 1279 198 1309 210
rect 1901 204 1902 230
rect 1928 204 1929 230
rect 1901 201 1929 204
rect 1289 64 1309 100
rect 1279 32 1309 64
rect 1897 69 1926 72
rect 1897 50 1899 69
rect 1849 43 1899 50
rect 1925 43 1926 69
rect 1849 40 1925 43
rect 1849 32 1921 40
rect 1289 31 1309 32
use sky130_hilas_VinjTgate4Single  sky130_hilas_VinjTgate4Single_0
timestamp 1637803711
transform -1 0 2917 0 -1 617
box 1050 -28 1622 631
use sky130_hilas_VinjDecode2to4  sky130_hilas_VinjDecode2to4_0
timestamp 1637801776
transform 1 0 637 0 1 -54
box -637 54 658 670
<< end >>
