magic
tech sky130A
timestamp 1607178257
<< poly >>
rect -9 11 18 19
rect -9 -6 -4 11
rect 13 -6 18 11
rect -9 -14 18 -6
<< polycont >>
rect -4 -6 13 11
<< locali >>
rect -4 11 13 19
rect -4 -14 13 -6
<< end >>
