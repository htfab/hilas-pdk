magic
tech sky130A
timestamp 1628698563
<< checkpaint >>
rect -456 -684 837 627
<< error_s >>
rect 90 368 129 371
rect 90 326 129 329
rect 89 272 128 275
rect 89 230 128 233
rect 89 176 128 179
rect 89 134 128 137
rect 89 80 128 83
rect 89 38 128 41
rect 89 -16 128 -13
rect 89 -58 128 -55
rect 90 -112 129 -109
rect 90 -154 129 -151
use sky130_hilas_pFETdevice01b  sky130_hilas_pFETdevice01b_1
timestamp 1628698535
transform 1 0 107 0 1 60
box -79 -114 108 43
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_0
timestamp 1628698561
transform 1 0 107 0 1 -36
box -79 -78 82 43
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_3
timestamp 1628698561
transform 1 0 107 0 1 156
box -79 -78 82 43
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_6
timestamp 1628698561
transform 1 0 107 0 1 252
box -79 -78 82 43
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_0
timestamp 1628698452
transform 1 0 108 0 1 348
box -80 -78 92 43
use sky130_hilas_pFETdevice01a  sky130_hilas_pFETdevice01a_0
timestamp 1628698547
transform 1 0 108 0 1 -132
box -80 -42 81 43
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
