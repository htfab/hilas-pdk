magic
tech sky130A
timestamp 1632410747
<< nwell >>
rect -173 126 244 333
<< pmos >>
rect -116 243 137 314
rect -116 144 137 214
<< pdiff >>
rect -154 308 -116 314
rect -154 249 -145 308
rect -127 249 -116 308
rect -154 243 -116 249
rect 137 306 182 314
rect 137 243 155 306
rect 146 214 155 243
rect -152 208 -116 214
rect -152 149 -145 208
rect -127 149 -116 208
rect -152 144 -116 149
rect 137 149 155 214
rect 173 149 182 306
rect 137 144 182 149
<< pdiffc >>
rect -145 249 -127 308
rect -145 149 -127 208
rect 155 149 173 306
<< nsubdiff >>
rect 182 304 224 314
rect 182 149 194 304
rect 212 149 224 304
rect 182 144 224 149
<< nsubdiffcont >>
rect 194 149 212 304
<< poly >>
rect -116 314 137 330
rect -116 214 137 243
rect -116 120 137 144
rect -116 103 -108 120
rect 129 103 137 120
rect -116 98 137 103
<< polycont >>
rect -108 103 129 120
<< locali >>
rect -145 308 -127 316
rect -145 241 -127 249
rect 146 306 216 318
rect -145 208 -127 216
rect -145 141 -127 149
rect 146 149 155 306
rect 173 304 216 306
rect 173 149 194 304
rect 212 149 216 304
rect -145 120 -128 141
rect 146 138 216 149
rect -145 103 -108 120
rect 129 103 137 120
<< end >>
