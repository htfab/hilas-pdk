magic
tech sky130A
timestamp 1632257797
<< checkpaint >>
rect -412 2223 1039 2249
rect -425 2207 1039 2223
rect -473 2181 1039 2207
rect -486 1449 1039 2181
rect -568 1407 2331 1449
rect -630 -434 2331 1407
rect -630 -454 2279 -434
rect -602 -623 2279 -454
rect -602 -628 830 -623
rect 847 -628 2279 -623
<< error_s >>
rect 361 502 1371 579
rect 1477 495 1498 567
rect 23 480 27 494
rect 37 462 41 480
<< nwell >>
rect 361 495 1371 502
<< locali >>
rect 389 502 406 503
rect 1286 502 1307 580
rect 1353 502 1370 570
rect 228 479 1371 502
rect 228 123 245 479
rect 294 0 311 446
rect 389 123 406 479
rect 457 0 474 442
rect 548 123 565 479
rect 617 0 634 450
rect 710 123 727 479
rect 779 0 796 445
rect 872 125 889 479
rect 939 0 956 450
rect 1032 126 1049 479
rect 1101 0 1118 450
rect 1193 125 1210 479
rect 1261 0 1278 448
rect 1354 122 1371 479
rect 1422 0 1439 466
<< metal1 >>
rect 665 355 1010 372
rect 820 102 838 256
rect 990 171 1010 355
rect 295 0 1639 23
<< metal2 >>
rect 27 577 696 596
rect 27 495 197 501
rect 339 495 361 541
rect 831 496 856 572
rect 831 495 859 496
rect 27 480 859 495
rect 27 456 37 480
rect 181 465 859 480
rect 1002 308 1022 564
rect 27 287 1022 308
rect 1162 210 1177 584
rect 1262 568 1378 596
rect 1337 567 1378 568
rect 27 190 1178 210
rect 27 78 845 98
use sky130_hilas_DAC6TransistorStack01a  sky130_hilas_DAC6TransistorStack01a_0
timestamp 1632256322
transform 1 0 0 0 1 176
box 0 0 172 601
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_8
timestamp 1632251409
transform 1 0 193 0 1 565
box 0 0 33 55
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_9
timestamp 1632251409
transform 1 0 34 0 1 564
box 0 0 33 55
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_10
timestamp 1632251409
transform 1 0 20 0 1 433
box 0 0 33 55
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_11
timestamp 1632251409
transform 1 0 26 0 1 338
box 0 0 33 55
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_12
timestamp 1632251409
transform 1 0 26 0 1 244
box 0 0 33 55
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1632251332
transform 1 0 302 0 1 7
box 0 0 23 29
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_7
timestamp 1632251409
transform 0 1 348 -1 0 548
box 0 0 33 55
use sky130_hilas_li2m1  sky130_hilas_li2m1_6
timestamp 1632251332
transform 1 0 464 0 1 7
box 0 0 23 29
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_6
timestamp 1632251409
transform 1 0 513 0 1 564
box 0 0 33 55
use sky130_hilas_li2m1  sky130_hilas_li2m1_7
timestamp 1632251332
transform 1 0 624 0 1 7
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1632251332
transform 1 0 786 0 1 7
box 0 0 23 29
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_5
timestamp 1632251409
transform 1 0 674 0 1 564
box 0 0 33 55
use sky130_hilas_li2m1  sky130_hilas_li2m1_5
timestamp 1632251332
transform 1 0 946 0 1 7
box 0 0 23 29
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_3
timestamp 1632251409
transform 1 0 997 0 1 565
box 0 0 33 55
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_4
timestamp 1632251409
transform 1 0 836 0 1 564
box 0 0 33 55
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1632251372
transform 1 0 826 0 1 82
box 0 0 32 32
use sky130_hilas_li2m1  sky130_hilas_li2m1_2
timestamp 1632251332
transform 1 0 1108 0 1 7
box 0 0 23 29
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_2
timestamp 1632251409
transform 1 0 1158 0 1 565
box 0 0 33 55
use sky130_hilas_li2m1  sky130_hilas_li2m1_3
timestamp 1632251332
transform 1 0 1268 0 1 7
box 0 0 23 29
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1632251356
transform 1 0 1355 0 1 565
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1632251356
transform 1 0 1288 0 1 565
box 0 0 34 33
use sky130_hilas_li2m1  sky130_hilas_li2m1_4
timestamp 1632251332
transform 1 0 1429 0 1 7
box 0 0 23 29
use sky130_hilas_DAC6TransistorStack01a  sky130_hilas_DAC6TransistorStack01a_1
timestamp 1632256322
transform 1 0 1449 0 1 176
box 0 0 172 601
use sky130_hilas_DAC6TransistorStack01  sky130_hilas_DAC6TransistorStack01_1
timestamp 1632256321
transform 1 0 157 0 1 976
box 0 0 173 601
use sky130_hilas_DAC6TransistorStack01  sky130_hilas_DAC6TransistorStack01_0
timestamp 1632256321
transform 1 0 144 0 1 950
box 0 0 173 601
<< labels >>
rlabel metal2 1262 582 1337 596 0 Vdd
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
