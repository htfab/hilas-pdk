magic
tech sky130A
magscale 1 2
timestamp 1632256325
<< error_s >>
rect 96 154 102 182
rect 164 156 166 178
rect 68 116 74 154
rect 96 146 132 154
rect 96 140 102 146
rect 128 116 132 146
rect 324 106 330 156
rect 358 126 364 178
rect 150 84 201 97
<< nwell >>
rect 0 12 406 210
<< pmos >>
rect 206 84 284 168
<< pdiff >>
rect 150 140 206 168
rect 150 106 160 140
rect 194 106 206 140
rect 150 84 206 106
rect 284 140 338 168
rect 284 106 296 140
rect 330 106 338 140
rect 284 84 338 106
<< pdiffc >>
rect 160 106 194 140
rect 296 106 330 140
<< poly >>
rect 206 168 284 194
rect 82 68 134 84
rect 206 68 284 84
rect 82 38 284 68
<< locali >>
rect 132 140 194 156
rect 132 120 160 140
rect 128 116 160 120
rect 160 90 194 106
rect 296 140 330 156
rect 296 90 330 106
<< metal2 >>
rect 0 116 74 154
rect 0 32 76 70
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1632251356
transform 1 0 356 0 1 120
box 0 0 68 66
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1632251356
transform 1 0 96 0 1 140
box 0 0 68 66
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_0
timestamp 1632251409
transform 0 1 68 -1 0 66
box 0 0 66 110
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
