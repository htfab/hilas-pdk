magic
tech sky130A
timestamp 1628616702
<< metal1 >>
rect 3 29 29 32
rect 3 0 29 3
<< via1 >>
rect 3 3 29 29
<< metal2 >>
rect 0 3 3 29
rect 29 3 32 29
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
