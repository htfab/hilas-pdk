* NGSPICE file created from /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_nFET03a.ext - technology: sky130A


* Top level circuit /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_nFET03a

X0 m2_150_6# a_n184_n58# m2_n222_4# $SUB sky130_fd_pr__nfet_01v8 w=350000u l=270000u
.end

