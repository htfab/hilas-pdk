magic
tech sky130A
timestamp 1628617012
<< error_p >>
rect 83 112 84 113
rect 111 112 112 113
rect 162 112 163 113
rect 190 112 191 113
rect 241 112 242 113
rect 269 112 270 113
rect 320 112 321 113
rect 348 112 349 113
rect 82 111 83 112
rect 112 111 113 112
rect 161 111 162 112
rect 191 111 192 112
rect 240 111 241 112
rect 270 111 271 112
rect 319 111 320 112
rect 349 111 350 112
rect 82 83 83 84
rect 112 83 113 84
rect 161 83 162 84
rect 191 83 192 84
rect 240 83 241 84
rect 270 83 271 84
rect 319 83 320 84
rect 349 83 350 84
rect 83 82 84 83
rect 111 82 112 83
rect 162 82 163 83
rect 190 82 191 83
rect 241 82 242 83
rect 269 82 270 83
rect 320 82 321 83
rect 348 82 349 83
<< nwell >>
rect 0 0 432 195
<< mvpmos >>
rect 33 112 399 162
rect 33 83 83 112
rect 112 83 162 112
rect 191 83 241 112
rect 270 83 320 112
rect 349 83 399 112
rect 33 33 399 83
<< mvpdiff >>
rect 83 106 112 112
rect 83 89 89 106
rect 106 89 112 106
rect 83 83 112 89
rect 162 106 191 112
rect 162 89 168 106
rect 185 89 191 106
rect 162 83 191 89
rect 241 106 270 112
rect 241 89 247 106
rect 264 89 270 106
rect 241 83 270 89
rect 320 106 349 112
rect 320 89 326 106
rect 343 89 349 106
rect 320 83 349 89
<< mvpdiffc >>
rect 89 89 106 106
rect 168 89 185 106
rect 247 89 264 106
rect 326 89 343 106
<< poly >>
rect 19 162 413 175
rect 19 33 33 162
rect 399 33 413 162
rect 19 19 413 33
<< locali >>
rect 25 140 405 167
rect 25 123 208 140
rect 225 123 405 140
rect 25 106 405 123
rect 25 89 89 106
rect 106 89 168 106
rect 185 105 247 106
rect 185 89 208 105
rect 25 88 208 89
rect 225 89 247 105
rect 264 89 326 106
rect 343 89 405 106
rect 225 88 405 89
rect 25 71 405 88
rect 25 54 208 71
rect 225 54 405 71
rect 25 26 405 54
<< viali >>
rect 208 123 225 140
rect 208 88 225 105
rect 208 54 225 71
<< metal1 >>
rect 204 140 228 146
rect 204 123 208 140
rect 225 123 228 140
rect 204 105 228 123
rect 204 88 208 105
rect 225 88 228 105
rect 204 82 228 88
rect 205 71 228 82
rect 205 54 208 71
rect 225 54 228 71
rect 205 17 228 54
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
