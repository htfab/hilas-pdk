magic
tech sky130A
timestamp 1634057796
<< checkpaint >>
rect -630 -603 719 929
<< error_s >>
rect 363 173 380 174
rect 387 162 388 203
rect 351 150 355 162
rect 387 150 392 162
rect 387 134 388 150
rect 387 102 388 133
rect 387 44 388 73
<< nwell >>
rect 217 304 436 477
<< nmos >>
rect 270 203 303 232
rect 355 203 388 232
rect 270 73 303 102
rect 355 73 388 102
<< pmos >>
rect 238 356 306 386
rect 342 356 410 386
<< ndiff >>
rect 270 256 303 260
rect 270 239 278 256
rect 295 239 303 256
rect 270 232 303 239
rect 355 256 388 260
rect 355 239 363 256
rect 380 239 388 256
rect 355 232 388 239
rect 270 196 303 203
rect 270 179 278 196
rect 295 179 303 196
rect 270 173 303 179
rect 270 125 303 132
rect 270 108 278 125
rect 295 108 303 125
rect 270 102 303 108
rect 355 196 388 203
rect 355 179 363 196
rect 380 179 388 196
rect 355 173 388 179
rect 355 126 388 133
rect 355 109 363 126
rect 380 109 388 126
rect 355 102 388 109
rect 270 66 303 73
rect 270 49 277 66
rect 295 49 303 66
rect 270 45 303 49
rect 355 67 388 73
rect 355 50 362 67
rect 381 50 388 67
rect 355 44 388 50
<< pdiff >>
rect 238 410 306 416
rect 238 393 246 410
rect 264 393 282 410
rect 300 393 306 410
rect 238 386 306 393
rect 342 410 410 416
rect 342 393 350 410
rect 368 393 387 410
rect 406 393 410 410
rect 342 386 410 393
rect 238 349 306 356
rect 238 332 246 349
rect 264 332 282 349
rect 300 332 306 349
rect 238 323 306 332
rect 342 349 410 356
rect 342 332 348 349
rect 366 332 384 349
rect 402 332 410 349
rect 342 328 410 332
rect 349 323 410 328
<< ndiffc >>
rect 278 239 295 256
rect 363 239 380 256
rect 278 179 295 196
rect 278 108 295 125
rect 363 179 380 196
rect 363 109 380 126
rect 277 49 295 66
rect 362 50 381 67
<< pdiffc >>
rect 246 393 264 410
rect 282 393 300 410
rect 350 393 368 410
rect 387 393 406 410
rect 246 332 264 349
rect 282 332 300 349
rect 348 332 366 349
rect 384 332 402 349
<< psubdiff >>
rect 270 161 303 173
rect 270 144 278 161
rect 295 144 303 161
rect 270 132 303 144
rect 355 162 388 173
rect 355 145 363 162
rect 380 145 388 162
rect 355 134 388 145
rect 355 133 387 134
<< nsubdiff >>
rect 238 445 306 457
rect 238 428 246 445
rect 264 428 282 445
rect 300 428 306 445
rect 238 416 306 428
rect 342 445 410 457
rect 342 428 350 445
rect 368 428 387 445
rect 406 428 410 445
rect 342 416 410 428
<< psubdiffcont >>
rect 278 144 295 161
rect 363 145 380 162
<< nsubdiffcont >>
rect 246 428 264 445
rect 282 428 300 445
rect 350 428 368 445
rect 387 428 406 445
<< poly >>
rect 225 356 238 386
rect 306 356 342 386
rect 410 356 423 386
rect 314 312 331 356
rect 308 304 335 312
rect 308 287 313 304
rect 330 287 335 304
rect 308 279 335 287
rect 0 215 27 219
rect 245 203 270 232
rect 303 203 316 232
rect 341 203 355 232
rect 388 203 411 232
rect 245 102 261 203
rect 395 102 411 203
rect 245 73 270 102
rect 303 73 316 102
rect 340 73 355 102
rect 388 73 411 102
rect 0 69 27 72
rect 245 34 261 73
rect 245 26 304 34
rect 395 33 411 73
rect 245 9 277 26
rect 295 9 304 26
rect 245 3 304 9
rect 355 25 411 33
rect 355 8 364 25
rect 381 8 411 25
rect 355 3 411 8
<< polycont >>
rect 313 287 330 304
rect 277 9 295 26
rect 364 8 381 25
<< locali >>
rect 238 428 246 445
rect 264 428 282 445
rect 300 428 350 445
rect 368 428 387 445
rect 406 428 414 445
rect 238 410 414 428
rect 238 393 246 410
rect 264 393 282 410
rect 300 393 350 410
rect 368 393 387 410
rect 406 393 414 410
rect 238 332 246 349
rect 264 332 282 349
rect 300 332 309 349
rect 340 332 348 349
rect 366 332 384 349
rect 402 332 410 349
rect 273 315 309 332
rect 273 304 338 315
rect 273 287 313 304
rect 330 287 338 304
rect 273 279 338 287
rect 273 256 300 279
rect 363 257 388 332
rect 355 256 388 257
rect 270 239 278 256
rect 295 239 303 256
rect 355 239 363 256
rect 380 239 388 256
rect 266 179 278 196
rect 295 179 307 196
rect 266 172 307 179
rect 351 179 363 196
rect 380 179 392 196
rect 351 172 392 179
rect 266 162 392 172
rect 266 161 363 162
rect 266 144 278 161
rect 295 145 363 161
rect 380 145 392 162
rect 295 144 392 145
rect 266 134 392 144
rect 266 125 307 134
rect 266 108 278 125
rect 295 108 307 125
rect 351 126 392 134
rect 351 109 363 126
rect 380 109 392 126
rect 269 49 277 66
rect 295 49 303 66
rect 354 50 362 67
rect 381 50 390 67
rect 354 49 390 50
rect 277 26 295 49
rect 277 0 295 9
rect 362 25 381 49
rect 362 8 364 25
rect 362 0 381 8
use sky130_hilas_nFET03  sky130_hilas_nFET03_3
timestamp 1634057709
transform 1 0 0 0 1 238
box 0 0 89 61
use sky130_hilas_nFET03  sky130_hilas_nFET03_2
timestamp 1634057709
transform 1 0 0 0 1 173
box 0 0 89 61
use sky130_hilas_nFET03  sky130_hilas_nFET03_1
timestamp 1634057709
transform 1 0 0 0 1 91
box 0 0 89 61
use sky130_hilas_nFET03  sky130_hilas_nFET03_0
timestamp 1634057709
transform 1 0 0 0 1 27
box 0 0 89 61
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
