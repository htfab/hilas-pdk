* NGSPICE file created from /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_TAcoreblock.ext - technology: sky130A

.subckt sky130_hilas_TACoreBlock2 VSUBS
X0 w_n122_224# a_n106_328# a_n106_328# w_n122_224# sky130_fd_pr__pfet_01v8 w=680000u l=300000u
X1 VSUBS a_n66_n378# a_n66_n378# VSUBS sky130_fd_pr__nfet_01v8 w=330000u l=290000u
X2 a_n106_328# a_n66_n378# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=330000u l=290000u
X3 a_128_272# a_124_n238# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=330000u l=290000u
X4 w_n122_224# a_n106_328# a_128_272# w_n122_224# sky130_fd_pr__pfet_01v8 w=680000u l=300000u
X5 VSUBS a_124_n238# a_124_n238# VSUBS sky130_fd_pr__nfet_01v8 w=330000u l=290000u
.ends


* Top level circuit /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_TAcoreblock

Xsky130_hilas_TACoreBlock2_0 VSUBS sky130_hilas_TACoreBlock2
.end

