magic
tech sky130A
timestamp 1627744303
<< error_p >>
rect -24 41 39 42
<< mvndiff >>
rect -24 35 39 41
rect -24 18 -18 35
rect -1 18 16 35
rect 33 18 39 35
rect -24 13 39 18
<< mvndiffc >>
rect -18 18 -1 35
rect 16 18 33 35
<< locali >>
rect -26 18 -18 35
rect 33 18 41 35
<< viali >>
rect -1 18 16 35
<< metal1 >>
rect -12 35 27 38
rect -12 18 -1 35
rect 16 18 27 35
rect -12 15 27 18
<< end >>
