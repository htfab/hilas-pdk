magic
tech sky130A
timestamp 1628707372
<< checkpaint >>
rect -699 1227 900 1249
rect -699 -581 1047 1227
rect -601 -582 1047 -581
rect -600 -603 1047 -582
rect -600 -614 708 -603
rect -600 -629 694 -614
<< nwell >>
rect 81 309 149 310
rect 81 306 157 309
rect 364 306 365 310
rect 402 18 464 588
<< nsubdiff >>
rect 420 551 446 570
rect 420 534 425 551
rect 442 534 446 551
rect 420 517 446 534
rect 420 500 425 517
rect 442 500 446 517
rect 420 488 446 500
<< nsubdiffcont >>
rect 425 534 442 551
rect 425 500 442 517
<< poly >>
rect 62 582 365 599
rect 62 310 81 582
rect 62 295 365 310
rect 62 104 82 295
rect 14 94 82 104
rect 14 77 19 94
rect 36 77 82 94
rect 14 60 82 77
rect 14 43 20 60
rect 37 43 82 60
rect 14 28 82 43
rect 14 26 364 28
rect 14 9 20 26
rect 37 11 364 26
rect 37 9 97 11
rect 14 4 97 9
rect 14 1 83 4
<< polycont >>
rect 19 77 36 94
rect 20 43 37 60
rect 20 9 37 26
<< locali >>
rect 425 532 442 534
rect 425 492 442 500
rect 96 316 112 319
rect 96 282 113 316
rect 151 315 167 319
rect 151 282 168 315
rect 206 282 223 322
rect 261 315 277 319
rect 316 315 332 319
rect 371 317 387 319
rect 261 282 278 315
rect 316 282 333 315
rect 371 282 388 317
rect 96 281 112 282
rect 151 281 167 282
rect 206 281 222 282
rect 261 281 277 282
rect 316 281 332 282
rect 371 281 387 282
rect 19 94 70 102
rect 36 77 71 94
rect 19 69 71 77
rect 20 60 71 69
rect 37 43 71 60
rect 20 26 71 43
rect 37 9 71 26
rect 20 1 71 9
<< viali >>
rect 425 551 442 568
rect 425 517 442 532
rect 425 515 442 517
<< metal1 >>
rect 414 579 440 599
rect 414 568 445 579
rect 414 551 425 568
rect 442 551 445 568
rect 414 532 445 551
rect 414 515 425 532
rect 442 515 445 532
rect 414 498 445 515
rect 414 0 440 498
<< metal2 >>
rect 33 560 339 561
rect 24 527 339 560
rect 24 282 56 527
rect 143 459 437 489
rect 362 455 437 459
rect 399 442 437 455
rect 402 355 437 442
rect 142 322 437 355
rect 24 249 340 282
rect 24 145 56 249
rect 24 113 340 145
rect 0 1 60 83
rect 402 78 437 322
rect 143 46 437 78
rect 143 45 414 46
use sky130_hilas_li2m2  sky130_hilas_li2m2_8
timestamp 1628707307
transform 1 0 43 0 1 63
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_7
timestamp 1628707307
transform 1 0 44 0 1 16
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_15
timestamp 1628707307
transform 1 0 156 0 1 59
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_17
timestamp 1628707307
transform 1 0 265 0 1 59
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_19
timestamp 1628707307
transform 1 0 375 0 1 60
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_9
timestamp 1628707307
transform 1 0 100 0 1 127
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_10
timestamp 1628707307
transform 1 0 210 0 1 127
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_6
timestamp 1628707307
transform 1 0 320 0 1 127
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628707307
transform 1 0 100 0 1 264
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628707307
transform 1 0 210 0 1 264
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1628707307
transform 1 0 320 0 1 264
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1628707307
transform 1 0 265 0 1 337
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_4
timestamp 1628707307
transform 1 0 156 0 1 337
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_5
timestamp 1628707307
transform 1 0 375 0 1 337
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_14
timestamp 1628707307
transform 1 0 210 0 1 542
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_18
timestamp 1628707307
transform 1 0 320 0 1 541
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_11
timestamp 1628707307
transform 1 0 101 0 1 542
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_16
timestamp 1628707307
transform 1 0 156 0 1 474
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_12
timestamp 1628707307
transform 1 0 265 0 1 472
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_13
timestamp 1628707307
transform 1 0 376 0 1 471
box 0 0 34 33
use sky130_hilas_pFETLargePart1  sky130_hilas_pFETLargePart1_0
timestamp 1628707368
transform 1 0 78 0 1 310
box 0 0 339 287
use sky130_hilas_pFETLargePart1  sky130_hilas_pFETLargePart1_1
timestamp 1628707368
transform 1 0 78 0 1 27
box 0 0 339 287
<< labels >>
rlabel metal2 422 415 436 489 0 DRAIN
port 3 nsew analog default
rlabel metal2 24 486 38 560 0 SOURCE
port 2 nsew analog default
rlabel metal2 0 1 10 83 0 GATE
port 1 nsew
rlabel metal1 414 591 440 599 0 WELL
port 4 nsew analog default
rlabel metal1 414 0 440 8 0 WELL
port 4 nsew analog default
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
