magic
tech sky130A
timestamp 1629137206
<< checkpaint >>
rect -574 1111 925 1204
rect -574 956 934 1111
rect -589 -352 934 956
rect -574 -507 934 -352
rect -574 -600 925 -507
<< nwell >>
rect 308 156 389 448
<< psubdiff >>
rect 315 562 359 586
rect 315 545 328 562
rect 345 545 359 562
rect 315 528 359 545
rect 315 511 328 528
rect 345 511 359 528
rect 315 494 359 511
rect 315 477 328 494
rect 345 477 359 494
rect 315 468 359 477
rect 316 104 359 130
rect 316 87 329 104
rect 346 87 359 104
rect 316 70 359 87
rect 316 53 329 70
rect 346 53 359 70
rect 316 36 359 53
rect 316 19 329 36
rect 346 19 359 36
rect 316 14 359 19
<< nsubdiff >>
rect 316 405 358 417
rect 316 387 327 405
rect 345 387 358 405
rect 316 368 358 387
rect 316 350 327 368
rect 345 350 358 368
rect 316 332 358 350
rect 316 314 327 332
rect 345 314 358 332
rect 316 296 358 314
rect 316 278 327 296
rect 345 278 358 296
rect 316 261 358 278
rect 316 243 328 261
rect 346 243 358 261
rect 316 225 358 243
rect 316 207 328 225
rect 346 207 358 225
rect 316 198 358 207
<< psubdiffcont >>
rect 328 545 345 562
rect 328 511 345 528
rect 328 477 345 494
rect 329 87 346 104
rect 329 53 346 70
rect 329 19 346 36
<< nsubdiffcont >>
rect 327 387 345 405
rect 327 350 345 368
rect 327 314 345 332
rect 327 278 345 296
rect 328 243 346 261
rect 328 207 346 225
<< locali >>
rect 291 562 353 579
rect 291 545 328 562
rect 345 545 353 562
rect 291 528 353 545
rect 291 511 328 528
rect 345 511 353 528
rect 291 494 353 511
rect 291 490 328 494
rect 317 477 328 490
rect 345 477 353 494
rect 317 475 353 477
rect 289 405 347 413
rect 289 387 327 405
rect 345 387 347 405
rect 289 374 347 387
rect 289 368 352 374
rect 289 350 327 368
rect 345 350 352 368
rect 289 332 352 350
rect 289 328 327 332
rect 289 311 292 328
rect 309 311 326 328
rect 345 314 352 332
rect 343 311 352 314
rect 289 296 352 311
rect 289 293 327 296
rect 289 276 292 293
rect 309 276 326 293
rect 345 278 352 296
rect 343 276 352 278
rect 289 261 352 276
rect 289 243 328 261
rect 346 243 352 261
rect 289 236 352 243
rect 289 225 347 236
rect 289 207 328 225
rect 346 207 347 225
rect 289 199 347 207
rect 291 104 346 114
rect 291 87 329 104
rect 291 70 346 87
rect 291 53 329 70
rect 291 36 346 53
rect 291 25 329 36
rect 329 11 346 19
<< viali >>
rect 292 311 309 328
rect 326 314 327 328
rect 327 314 343 328
rect 326 311 343 314
rect 292 276 309 293
rect 326 278 327 293
rect 327 278 343 293
rect 326 276 343 278
<< metal1 >>
rect 0 541 21 604
rect 0 525 248 541
rect 282 550 389 604
rect 282 541 301 550
rect 274 525 301 541
rect 0 524 301 525
rect 327 524 389 550
rect 0 510 389 524
rect 0 509 301 510
rect 0 483 246 509
rect 272 484 301 509
rect 327 484 389 510
rect 272 483 389 484
rect 0 473 389 483
rect 0 419 389 442
rect 0 392 37 419
rect 64 392 92 419
rect 119 392 389 419
rect 0 362 389 392
rect 0 361 92 362
rect 0 334 36 361
rect 63 335 92 361
rect 119 335 389 362
rect 63 334 389 335
rect 0 328 389 334
rect 0 311 292 328
rect 309 311 326 328
rect 343 311 389 328
rect 0 293 389 311
rect 0 278 292 293
rect 0 277 92 278
rect 0 258 37 277
rect 0 257 17 258
rect 0 250 37 257
rect 64 258 92 277
rect 64 251 92 257
rect 119 276 292 278
rect 309 276 326 293
rect 343 276 389 293
rect 119 258 389 276
rect 252 257 389 258
rect 119 251 389 257
rect 64 250 389 251
rect 0 227 389 250
rect 0 200 37 227
rect 64 225 389 227
rect 64 200 90 225
rect 0 198 90 200
rect 117 198 389 225
rect 0 163 389 198
rect 0 100 389 127
rect 0 74 262 100
rect 288 74 310 100
rect 336 74 389 100
rect 0 59 389 74
rect 0 33 260 59
rect 286 33 309 59
rect 335 33 389 59
rect 0 3 389 33
rect 0 0 17 3
rect 291 1 389 3
rect 290 0 389 1
<< via1 >>
rect 248 525 274 551
rect 301 524 327 550
rect 246 483 272 509
rect 301 484 327 510
rect 37 392 64 419
rect 92 392 119 419
rect 36 334 63 361
rect 92 335 119 362
rect 37 250 64 277
rect 92 251 119 278
rect 37 200 64 227
rect 90 198 117 225
rect 262 74 288 100
rect 310 74 336 100
rect 260 33 286 59
rect 309 33 335 59
<< metal2 >>
rect 22 419 152 604
rect 22 392 37 419
rect 64 392 92 419
rect 119 392 152 419
rect 22 362 152 392
rect 22 361 92 362
rect 22 334 36 361
rect 63 335 92 361
rect 119 335 152 362
rect 63 334 152 335
rect 22 278 152 334
rect 22 277 92 278
rect 22 250 37 277
rect 64 251 92 277
rect 119 251 152 278
rect 64 250 152 251
rect 22 227 152 250
rect 22 200 37 227
rect 64 225 152 227
rect 64 200 90 225
rect 22 198 90 200
rect 117 198 152 225
rect 22 0 152 198
rect 230 551 360 604
rect 230 525 248 551
rect 274 550 360 551
rect 274 525 301 550
rect 230 524 301 525
rect 327 524 360 550
rect 230 510 360 524
rect 230 509 301 510
rect 230 483 246 509
rect 272 484 301 509
rect 327 484 360 510
rect 272 483 360 484
rect 230 100 360 483
rect 230 74 262 100
rect 288 74 310 100
rect 336 74 360 100
rect 230 59 360 74
rect 230 33 260 59
rect 286 33 309 59
rect 335 33 360 59
rect 230 0 360 33
use sky130_hilas_decoup_cap_00  CapDeco_1
timestamp 1623107852
transform 1 0 -82 0 1 113
box 82 -113 390 194
use sky130_hilas_decoup_cap_00  CapDeco_0
timestamp 1623107852
transform 1 0 -82 0 -1 491
box 82 -113 390 194
<< labels >>
rlabel metal1 0 254 17 350 0 VPWR
port 1 nsew
rlabel metal1 372 256 389 350 0 VPWR
port 1 nsew
rlabel metal1 379 541 389 604 0 VGND
port 1 nsew
rlabel metal1 0 541 8 604 0 VGND
port 1 nsew
rlabel metal1 0 0 9 63 0 VGND
port 1 nsew
rlabel metal1 374 0 389 63 0 VGND
port 1 nsew
rlabel metal2 22 594 152 604 0 VPWR
port 1 nsew
rlabel metal2 230 596 360 604 0 VGND
port 2 nsew
rlabel metal2 22 0 152 12 0 VPWR
port 1 nsew
rlabel metal2 230 0 360 12 0 VGND
port 2 nsew
<< end >>
