VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_poly2m2
  CLASS BLOCK ;
  FOREIGN /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_poly2m2 ;
  ORIGIN 0.090 0.260 ;
  SIZE 0.330 BY 0.550 ;
  OBS
      LAYER li1 ;
        RECT -0.030 -0.200 0.180 0.250 ;
      LAYER met1 ;
        RECT -0.080 -0.260 0.240 0.290 ;
      LAYER met2 ;
        RECT -0.080 -0.030 0.240 0.290 ;
  END
END /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_poly2m2
END LIBRARY

