* SPICE3 file created from sky130_hilas_cellAttempt01.ext - technology: sky130A

.option scale=10000u

.subckt sky130_hilas_cellAttempt01 Vtun Vinj GateSel1 col1 Gate1 Drain1 Col1 Drain2
+ Col2 Drain3 Col4 Drain4
X0 FG3 Vtun Vtun xchvnwc w=59 l=50
X1 FG4 Vtun Vtun xchvnwc w=59 l=50
X2 FG2 Vtun Vtun xchvnwc w=59 l=50
X3 FG1 Vtun Vtun xchvnwc w=59 l=50
M1000 Vinj GateSel1 sky130_hilas_horizPcell01_0/a_n172_81# Vinj phv w=31 l=50
+  ad=4216 pd=520 as=682 ps=106
M1001 col1 FG2 Col2 Vinj phv w=30 l=50
+  ad=3720 pd=488 as=870 ps=118
M1002 sky130_hilas_horizPcell01_0/a_n172_81# FG2 Drain2 Vinj phv w=31 l=50
+  ad=0 pd=0 as=992 ps=126
M1003 Vinj GateSel1 sky130_hilas_horizPcell01_1/a_n172_81# Vinj phv w=31 l=50
+  ad=0 pd=0 as=682 ps=106
M1004 col1 FG4 Col4 Vinj phv w=30 l=50
+  ad=0 pd=0 as=870 ps=118
M1005 sky130_hilas_horizPcell01_1/a_n172_81# FG4 Drain4 Vinj phv w=31 l=50
+  ad=0 pd=0 as=992 ps=126
M1006 Vinj GateSel1 sky130_hilas_horizPcell01_2/a_n172_81# Vinj phv w=31 l=50
+  ad=0 pd=0 as=682 ps=106
M1007 col1 FG3 Col1 Vinj phv w=30 l=50
+  ad=0 pd=0 as=1740 ps=236
M1008 sky130_hilas_horizPcell01_2/a_n172_81# FG3 Drain3 Vinj phv w=31 l=50
+  ad=0 pd=0 as=992 ps=126
M1009 Vinj GateSel1 sky130_hilas_horizPcell01_3/a_n172_81# Vinj phv w=31 l=50
+  ad=0 pd=0 as=682 ps=106
M1010 col1 FG1 Col1 Vinj phv w=30 l=50
+  ad=0 pd=0 as=0 ps=0
M1011 sky130_hilas_horizPcell01_3/a_n172_81# FG1 Drain1 Vinj phv w=31 l=50
+  ad=0 pd=0 as=992 ps=126
X4 FG4 Gate1 Gate1 xchvnwc w=111 l=64
X5 FG2 Gate1 Gate1 xchvnwc w=111 l=64
X6 FG3 Gate1 Gate1 xchvnwc w=111 l=64
X7 FG1 Gate1 Gate1 xchvnwc w=111 l=64
C0 Col1 Drain3 2.14fF
C1 Col1 Drain1 2.14fF
C2 Drain2 Col2 2.14fF
C3 Drain4 Col4 2.17fF
C4 Gate1 SUB 2.93fF
C5 Vinj SUB 2.30fF
C6 Vtun SUB 2.73fF
.ends
