magic
tech sky130A
timestamp 1627401173
<< error_s >>
rect 1432 532 1438 538
rect 1485 532 1491 538
rect 1597 532 1603 538
rect 1650 532 1656 538
rect 1426 482 1432 488
rect 1491 482 1497 488
rect 1591 482 1597 488
rect 1656 482 1662 488
rect 957 473 963 479
rect 1062 473 1068 479
rect 2020 473 2026 479
rect 2125 473 2131 479
rect 951 423 957 429
rect 1068 423 1074 429
rect 2014 423 2020 429
rect 2131 423 2137 429
rect 1825 288 1842 289
rect 1825 271 1842 272
rect 1263 254 1264 267
rect 957 172 963 178
rect 1062 172 1068 178
rect 2020 172 2026 178
rect 2125 172 2131 178
rect 951 122 957 128
rect 1068 122 1074 128
rect 1432 118 1438 124
rect 1485 118 1491 124
rect 1597 118 1603 124
rect 1650 118 1656 124
rect 2014 122 2020 128
rect 2131 122 2137 128
rect 1426 68 1432 74
rect 1491 68 1497 74
rect 1591 68 1597 74
rect 1656 68 1662 74
<< nwell >>
rect 396 604 594 605
rect 2692 604 2839 605
rect 3077 587 3205 605
rect 396 537 403 555
rect 396 50 404 68
rect 3077 0 3205 19
<< locali >>
rect 1245 340 1265 348
rect 1245 323 1246 340
rect 1263 323 1265 340
rect 1245 271 1265 323
rect 1245 254 1247 271
rect 1264 254 1265 271
rect 1245 247 1265 254
rect 1820 340 1849 348
rect 1820 323 1825 340
rect 1842 323 1849 340
rect 1820 272 1849 323
rect 1820 255 1825 272
rect 1842 255 1849 272
rect 1820 247 1849 255
<< viali >>
rect 1246 323 1263 340
rect 1247 254 1264 271
rect 1825 323 1842 340
rect 1825 255 1842 272
<< metal1 >>
rect 420 600 448 605
rect 420 599 452 600
rect 473 599 492 605
rect 420 573 423 599
rect 449 573 452 599
rect 1121 596 1144 604
rect 1243 596 1266 604
rect 1472 589 1616 605
rect 1822 596 1845 605
rect 1944 597 1967 605
rect 2596 597 2615 605
rect 2640 600 2668 605
rect 2640 598 2672 600
rect 420 572 452 573
rect 2640 572 2643 598
rect 2669 572 2672 598
rect 3009 591 3043 605
rect 3075 590 3103 605
rect 2640 570 2672 572
rect 1244 292 1276 294
rect 1244 264 1247 292
rect 1273 266 1276 292
rect 1264 264 1276 266
rect 1814 286 1846 289
rect 1814 260 1817 286
rect 1843 260 1846 286
rect 1814 257 1825 260
rect 1842 257 1846 260
rect 2858 47 2891 49
rect 1814 34 1846 36
rect 1814 8 1817 34
rect 1843 8 1846 34
rect 2858 21 2861 47
rect 2888 21 2891 47
rect 2858 20 2891 21
rect 1814 6 1846 8
rect 2857 19 3009 20
rect 2857 6 3043 19
rect 2596 0 2615 5
rect 2640 0 2668 5
rect 3009 0 3043 6
rect 3076 0 3103 21
<< via1 >>
rect 423 573 449 599
rect 2643 572 2669 598
rect 1247 271 1273 292
rect 1247 266 1264 271
rect 1264 266 1273 271
rect 1817 272 1843 286
rect 1817 260 1825 272
rect 1825 260 1842 272
rect 1842 260 1843 272
rect 1817 8 1843 34
rect 2861 21 2888 47
<< metal2 >>
rect 420 599 452 600
rect 420 573 423 599
rect 449 588 452 599
rect 2640 598 2672 600
rect 2640 588 2643 598
rect 449 573 2643 588
rect 420 572 2643 573
rect 2669 572 2672 598
rect 2752 578 2783 602
rect 420 570 2672 572
rect 396 537 403 555
rect 2863 515 2885 517
rect 1286 477 1370 497
rect 2858 481 2885 515
rect 1331 430 2345 452
rect 2684 431 2719 453
rect 1326 333 2227 355
rect 1244 292 1276 294
rect 1244 266 1247 292
rect 1273 289 1276 292
rect 1273 286 1846 289
rect 1273 266 1817 286
rect 1244 264 1817 266
rect 1814 260 1817 264
rect 1843 260 1846 286
rect 1814 257 1846 260
rect 1331 155 1897 177
rect 1281 125 1329 126
rect 1281 101 1370 125
rect 1875 122 1897 155
rect 2205 172 2227 333
rect 2323 310 2345 430
rect 2865 424 2885 425
rect 2865 391 2887 424
rect 2867 390 2887 391
rect 2760 311 2792 335
rect 3194 334 3205 357
rect 2320 306 2345 310
rect 2320 242 2346 306
rect 3194 252 3205 274
rect 2320 221 2733 242
rect 2712 207 2733 221
rect 2712 186 2899 207
rect 2205 150 2490 172
rect 2312 122 2899 127
rect 1875 106 2899 122
rect 1875 100 2351 106
rect 396 50 404 68
rect 2858 47 2891 49
rect 1814 35 1846 36
rect 2858 35 2861 47
rect 1814 34 2861 35
rect 1814 8 1817 34
rect 1843 21 2861 34
rect 2888 21 2891 47
rect 1843 19 2891 21
rect 1843 18 1883 19
rect 1843 8 1846 18
rect 1814 6 1846 8
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1608069483
transform 1 0 3050 0 1 41
box -172 -22 155 550
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1608384750
transform 1 0 2558 0 -1 165
box 133 -440 320 165
use sky130_hilas_FGBiasWeakGate2x1cell  sky130_hilas_FGBiasWeakGate2x1cell_0
timestamp 1625491133
transform -1 0 1153 0 1 382
box -396 -382 757 223
use sky130_hilas_FGBias2x1cell  sky130_hilas_FGBias2x1cell_0
timestamp 1625491133
transform 1 0 1935 0 1 382
box -396 -382 757 223
<< labels >>
rlabel metal2 1286 477 1322 496 0 VIN11
port 2 nsew analog default
rlabel metal2 1281 101 1317 126 0 VIN12
port 1 nsew analog default
rlabel metal1 3009 599 3043 605 0 VGND
port 7 nsew analog default
rlabel metal1 3075 599 3103 605 0 VPWR
port 6 nsew analog default
rlabel metal1 3076 0 3103 6 0 VPWR
port 6 nsew power default
rlabel metal1 3009 0 3043 6 0 VGND
port 7 nsew ground default
rlabel metal2 2760 311 2792 335 0 VIN21
port 3 nsew analog default
rlabel metal2 2752 578 2783 602 1 VIN22
port 4 n analog default
rlabel metal1 2640 597 2668 605 0 VINJ
port 8 nsew power default
rlabel metal1 2640 0 2668 5 0 VINJ
port 8 nsew power default
rlabel metal2 3194 334 3205 357 0 OUTPUT1
port 9 nsew analog default
rlabel metal2 3194 252 3205 274 0 OUTPUT2
port 10 nsew analog default
rlabel metal2 396 537 403 555 0 DRAIN1
port 11 nsew
rlabel metal2 396 50 404 68 0 DRAIN2
port 12 nsew
rlabel metal1 420 598 448 605 0 VINJ
port 8 nsew
rlabel metal1 473 599 492 605 0 COLSEL2
port 13 nsew
rlabel metal1 1121 596 1144 604 0 GATE2
port 14 nsew
rlabel metal1 1243 596 1266 604 0 VGND
port 7 nsew
rlabel metal1 1944 597 1967 605 0 GATE1
port 15 nsew
rlabel metal1 1822 597 1845 605 0 VGND
port 7 nsew
rlabel metal1 2596 597 2615 605 0 COLSEL1
port 16 nsew
rlabel metal1 2596 0 2615 5 0 COLSEL1
port 16 nsew
rlabel metal1 1514 593 1574 605 0 VTUN
port 17 nsew
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
