magic
tech sky130A
timestamp 1607478930
use pFETdevice01aa  pFETdevice01aa_0
timestamp 1607478455
transform 1 0 108 0 1 348
box -80 -78 92 43
use pFETdevice01a  pFETdevice01a_0
timestamp 1607477942
transform 1 0 108 0 1 -132
box -80 -42 81 43
use pFETdevice01  pFETdevice01_0
timestamp 1607471549
transform 1 0 107 0 1 -36
box -79 -78 82 43
use pFETdevice01  pFETdevice01_3
timestamp 1607471549
transform 1 0 107 0 1 156
box -79 -78 82 43
use pFETdevice01  pFETdevice01_6
timestamp 1607471549
transform 1 0 107 0 1 252
box -79 -78 82 43
use pFETdevice01b  pFETdevice01b_1
timestamp 1607475333
transform 1 0 107 0 1 60
box -79 -114 108 43
<< end >>
