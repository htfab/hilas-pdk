magic
tech sky130A
timestamp 1632172832
<< nwell >>
rect -289 41 -33 232
<< mvpmos >>
rect -222 126 -172 180
<< mvpdiff >>
rect -251 174 -222 180
rect -251 132 -247 174
rect -229 132 -222 174
rect -251 126 -222 132
rect -172 169 -143 180
rect -172 152 -166 169
rect -147 152 -143 169
rect -172 126 -143 152
<< mvpdiffc >>
rect -247 132 -229 174
rect -166 152 -147 169
<< mvnsubdiff >>
rect -100 169 -66 183
rect -100 151 -93 169
rect -73 151 -66 169
rect -100 139 -66 151
<< mvnsubdiffcont >>
rect -93 151 -73 169
<< poly >>
rect -222 180 -172 193
rect -222 117 -172 126
rect -289 100 -172 117
<< locali >>
rect -255 174 -221 176
rect -255 132 -247 174
rect -229 132 -221 174
rect -166 169 -146 177
rect -147 152 -146 169
rect -166 138 -146 152
rect -166 121 -165 138
rect -148 121 -146 138
rect -166 117 -146 121
rect -94 169 -72 177
rect -94 151 -93 169
rect -73 151 -72 169
rect -94 135 -72 151
rect -94 118 -92 135
rect -75 118 -72 135
rect -93 115 -72 118
rect -93 111 -73 115
<< viali >>
rect -165 121 -148 138
rect -92 118 -75 135
<< metal1 >>
rect -166 146 -150 232
rect -85 181 -69 232
rect -85 172 -68 181
rect -96 167 -68 172
rect -166 141 -145 146
rect -168 138 -145 141
rect -168 121 -165 138
rect -148 121 -145 138
rect -168 117 -145 121
rect -96 135 -69 167
rect -96 118 -92 135
rect -75 118 -69 135
rect -166 115 -146 117
rect -166 42 -150 115
rect -96 112 -69 118
rect -85 42 -69 112
<< metal2 >>
rect -289 140 -280 158
rect -250 140 -33 158
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1629420194
transform 1 0 -266 0 -1 156
box -14 -15 20 18
<< end >>
