magic
tech sky130A
magscale 1 2
timestamp 1632256354
<< checkpaint >>
rect -1260 1300 10648 5924
rect 7050 618 10286 1300
<< error_s >>
rect 1498 4334 1508 4362
rect 9088 4354 9098 4362
rect 9088 4334 9216 4354
rect 9088 4323 9099 4334
rect 2282 3770 2314 3798
rect 2364 3768 2402 3796
rect 7724 3780 8386 3946
rect 9118 3820 9130 3890
rect 9146 3820 9158 3862
rect 8960 3808 9060 3820
rect 9104 3808 9204 3820
rect 9118 3796 9130 3808
rect 8194 3778 8232 3780
rect 8194 3772 8362 3778
rect 8892 3736 8960 3780
rect 9060 3736 9104 3780
rect 9146 3768 9158 3808
rect 9204 3736 9272 3780
rect 8904 3726 8928 3728
rect 8960 3726 9060 3736
rect 9104 3726 9204 3736
rect 2720 3710 2758 3716
rect 8904 3710 9274 3726
rect 1404 3606 1450 3678
rect 1482 3606 1498 3674
rect 2210 3644 2238 3680
rect 2720 3676 2722 3710
rect 2742 3676 2758 3710
rect 2720 3670 2758 3676
rect 2776 3660 2792 3694
rect 8910 3688 9274 3710
rect 8910 3674 8954 3688
rect 9052 3682 9274 3688
rect 9052 3674 9058 3682
rect 9146 3674 9192 3682
rect 8910 3634 8956 3674
rect 1324 3592 1380 3606
rect 1482 3506 1538 3606
rect 1762 3520 1768 3620
rect 1846 3520 1852 3620
rect 2034 3520 2038 3620
rect 2118 3520 2122 3620
rect 2802 3582 2814 3592
rect 8910 3544 8954 3634
rect 9052 3524 9114 3674
rect 9168 3656 9274 3674
rect 9218 3620 9274 3656
rect 9146 3572 9192 3574
rect 9138 3524 9192 3572
rect 9216 3524 9274 3574
rect 9016 3506 9114 3524
rect 1388 3446 1458 3506
rect 1482 3438 1498 3506
rect 1762 3364 1768 3462
rect 1846 3364 1852 3462
rect 1740 3240 1920 3364
rect 2034 3362 2038 3462
rect 2118 3362 2122 3462
rect 9098 3454 9114 3506
rect 9126 3496 9216 3506
rect 9138 3462 9216 3496
rect 9138 3454 9208 3462
rect 2720 3312 2758 3318
rect 2720 3278 2722 3312
rect 2746 3278 2758 3300
rect 2720 3272 2758 3278
rect 2780 3232 2814 3266
rect 2454 3216 2468 3222
rect 2452 3170 2468 3216
rect 2482 3188 2496 3196
rect 2480 3150 2496 3188
rect 2862 3158 2870 3316
rect 2890 3186 2898 3288
rect 2814 3134 2852 3140
rect 2814 3130 2830 3134
rect 2836 3130 2852 3134
rect 2814 3118 2852 3130
rect 2722 3098 2760 3104
rect 2722 3064 2724 3098
rect 2752 3064 2760 3098
rect 2786 3094 2852 3118
rect 3000 3114 3662 3172
rect 2870 3112 2904 3114
rect 2996 3112 3662 3114
rect 2870 3106 2886 3112
rect 2786 3084 2820 3094
rect 2862 3072 2886 3106
rect 2980 3084 3662 3112
rect 2722 3058 2760 3064
rect 2542 3002 2598 3028
rect 3000 3006 3662 3084
rect 3000 3004 3358 3006
rect 3040 3002 3104 3004
rect 3130 3002 3132 3004
rect 1762 2888 1768 2988
rect 1846 2888 1852 2988
rect 2034 2888 2038 2988
rect 2118 2888 2122 2988
rect 2570 2974 2626 3000
rect 3102 2942 3208 3002
rect 3528 2984 3570 3006
rect 3622 2990 3660 3006
rect 3704 2994 3746 3022
rect 3950 3006 3956 3020
rect 3130 2914 3132 2942
rect 3000 2870 3028 2906
rect 1762 2730 1768 2830
rect 1846 2730 1852 2830
rect 2034 2730 2038 2830
rect 2118 2730 2122 2830
rect 2800 2802 2812 2812
rect 2962 2802 2998 2804
rect 2996 2800 2998 2802
rect 4220 2784 4464 3400
rect 6132 3018 6376 3400
rect 8676 3240 9338 3454
rect 8126 3228 8190 3236
rect 8116 3200 8218 3208
rect 7494 3018 7558 3110
rect 6098 2990 6376 3018
rect 7402 2990 7440 3018
rect 7490 3006 7558 3018
rect 7494 3002 7558 3006
rect 7594 3006 7862 3172
rect 8364 3058 8620 3138
rect 8830 3110 8874 3200
rect 9030 3196 9042 3206
rect 8996 3154 9008 3188
rect 9030 3162 9096 3196
rect 8996 3138 9014 3154
rect 8676 3072 8874 3110
rect 8648 3066 8874 3072
rect 8986 3070 9008 3098
rect 8956 3066 9008 3070
rect 8648 3064 9008 3066
rect 8648 3058 8874 3064
rect 7594 3004 7812 3006
rect 6132 2784 6376 2990
rect 6894 2940 6940 2974
rect 7558 2942 7662 3002
rect 8332 2948 8338 3034
rect 8364 3032 8874 3058
rect 8956 3050 9008 3064
rect 8986 3044 9008 3050
rect 8892 3032 9008 3044
rect 8364 3030 9008 3032
rect 8364 3010 8874 3030
rect 8892 3010 9008 3030
rect 8364 3006 9008 3010
rect 8360 2976 8416 3006
rect 8548 2989 8599 3006
rect 8608 2990 9008 3006
rect 8620 2989 9008 2990
rect 8548 2988 9008 2989
rect 8548 2970 8608 2988
rect 8648 2980 9008 2988
rect 8648 2976 8874 2980
rect 8892 2976 9008 2980
rect 8648 2970 9008 2976
rect 8660 2962 8844 2970
rect 8676 2954 8844 2962
rect 8664 2952 8844 2954
rect 8382 2944 8414 2952
rect 8488 2944 8606 2946
rect 8660 2926 8844 2952
rect 8872 2946 9008 2970
rect 8888 2942 9008 2946
rect 8892 2930 9008 2942
rect 8354 2916 8386 2924
rect 8516 2916 8578 2918
rect 8484 2900 8516 2916
rect 8598 2914 8660 2926
rect 8518 2900 8550 2910
rect 8484 2868 8550 2900
rect 8574 2902 8582 2910
rect 8574 2868 8584 2902
rect 8598 2889 8618 2914
rect 8608 2872 8618 2889
rect 8630 2872 8648 2914
rect 8652 2911 8660 2914
rect 8664 2886 8682 2926
rect 8714 2925 8844 2926
rect 8726 2888 8766 2904
rect 8776 2888 8844 2925
rect 8872 2906 9008 2930
rect 8872 2900 8888 2906
rect 8892 2900 9008 2906
rect 8714 2886 8776 2888
rect 8676 2878 8782 2886
rect 8660 2872 8782 2878
rect 8598 2868 8782 2872
rect 8484 2858 8782 2868
rect 8484 2852 8522 2858
rect 8484 2850 8516 2852
rect 8488 2830 8494 2850
rect 8548 2846 8782 2858
rect 8536 2818 8782 2846
rect 8598 2817 8782 2818
rect 8796 2817 8822 2888
rect 8872 2848 9008 2900
rect 8892 2832 9008 2848
rect 8598 2816 8822 2817
rect 8548 2766 8702 2816
rect 8888 2800 9008 2832
rect 8598 2748 8652 2752
rect 8676 2748 8782 2766
rect 2672 2708 2724 2722
rect 2210 2670 2238 2706
rect 2704 2704 2724 2708
rect 2764 2700 2784 2710
rect 2678 2672 2680 2698
rect 2678 2670 2706 2672
rect 2282 2570 2314 2598
rect 2364 2570 2402 2598
rect 4362 2586 4446 2740
rect 8548 2726 8782 2748
rect 8536 2724 8782 2726
rect 7872 2708 7924 2722
rect 7872 2704 7892 2708
rect 8536 2698 8822 2724
rect 8598 2696 8822 2698
rect 8548 2694 8739 2696
rect 8740 2694 8822 2696
rect 8488 2664 8494 2684
rect 8548 2664 8822 2694
rect 8892 2686 9008 2800
rect 8872 2670 9008 2686
rect 9052 2676 9114 2806
rect 9127 2795 9203 2806
rect 9138 2778 9192 2795
rect 9146 2756 9192 2778
rect 9168 2730 9274 2756
rect 9218 2694 9274 2730
rect 8452 2630 8472 2664
rect 8484 2662 8516 2664
rect 8484 2656 8522 2662
rect 8548 2656 8796 2664
rect 8484 2636 8796 2656
rect 8910 2642 8954 2670
rect 9010 2642 9060 2656
rect 9146 2646 9192 2656
rect 9146 2642 9204 2646
rect 8910 2636 9060 2642
rect 8484 2630 8660 2636
rect 8714 2630 8796 2636
rect 8904 2630 9060 2636
rect 8484 2614 8550 2630
rect 8484 2598 8516 2614
rect 8518 2604 8550 2614
rect 8574 2612 8584 2630
rect 8574 2604 8582 2612
rect 8598 2610 8618 2630
rect 8630 2610 8648 2630
rect 8664 2618 8682 2628
rect 8714 2626 8822 2630
rect 8776 2618 8844 2626
rect 8910 2622 9060 2630
rect 8904 2620 9060 2622
rect 8598 2603 8652 2610
rect 8660 2603 8844 2618
rect 8910 2614 9060 2620
rect 9104 2614 9204 2642
rect 4446 2572 4530 2586
rect 8194 2570 8232 2598
rect 8598 2590 8844 2603
rect 8892 2604 9272 2614
rect 8892 2602 8948 2604
rect 8856 2596 8962 2602
rect 8856 2590 8948 2596
rect 8598 2588 8992 2590
rect 8618 2580 8652 2588
rect 8660 2564 8822 2588
rect 8842 2586 8992 2588
rect 8842 2584 8948 2586
rect 8856 2568 8948 2584
rect 8660 2563 8776 2564
rect 8660 2562 8725 2563
rect 8796 2562 8822 2564
rect 8882 2562 8948 2568
rect 8664 2560 8736 2562
rect 8676 2544 8736 2560
rect 8548 2538 8608 2544
rect 8648 2542 8736 2544
rect 8796 2556 8868 2562
rect 8882 2558 8964 2562
rect 8648 2538 8772 2542
rect 8548 2530 8772 2538
rect 8796 2530 8822 2556
rect 8882 2544 8948 2558
rect 8892 2542 8948 2544
rect 8548 2526 9338 2530
rect 8548 2522 8648 2526
rect 8536 2516 8652 2522
rect 8536 2494 8628 2516
rect 8648 2494 8652 2516
rect 8570 2492 8594 2494
rect 8598 2492 8648 2494
rect 8660 2492 9338 2526
rect 8548 2490 8628 2492
rect 8548 2476 8648 2490
rect 8676 2476 9338 2492
rect 8526 2468 8648 2476
rect 8526 2466 8652 2468
rect 8548 2464 8648 2466
rect 8548 2450 8598 2464
rect 8608 2458 8648 2464
rect 8608 2450 8648 2456
rect 8536 2448 8652 2450
rect 8526 2438 8652 2448
rect 8536 2424 8652 2438
rect 8536 2422 8628 2424
rect 8648 2422 8652 2424
rect 8574 2420 8594 2422
rect 8608 2420 8648 2422
rect 8660 2420 8694 2464
rect 8726 2458 8766 2476
rect 8726 2422 8766 2456
rect 8548 2388 8598 2420
rect 8608 2390 8628 2420
rect 8714 2394 8776 2422
rect 8660 2388 8776 2394
rect 8548 2372 8608 2388
rect 8648 2380 8764 2388
rect 8648 2372 8796 2380
rect 8548 2370 8796 2372
rect 8570 2352 8648 2370
rect 8660 2362 8796 2370
rect 8664 2352 8702 2354
rect 8704 2352 8796 2362
rect 8598 2326 8626 2344
rect 8660 2340 8694 2352
rect 8714 2350 8796 2352
rect 8660 2326 8714 2340
rect 8484 2300 8516 2316
rect 8570 2310 8578 2318
rect 8598 2314 8660 2326
rect 8518 2300 8550 2310
rect 8484 2268 8550 2300
rect 8570 2302 8582 2310
rect 8570 2272 8584 2302
rect 8598 2300 8626 2314
rect 8598 2289 8618 2300
rect 8608 2272 8618 2289
rect 8630 2272 8648 2314
rect 8652 2311 8660 2314
rect 8664 2286 8682 2326
rect 8714 2325 8776 2326
rect 8762 2304 8776 2325
rect 8726 2288 8776 2304
rect 8714 2278 8776 2288
rect 8660 2272 8776 2278
rect 8574 2268 8584 2272
rect 8598 2268 8776 2272
rect 8484 2258 8776 2268
rect 8484 2252 8522 2258
rect 8548 2256 8776 2258
rect 8484 2250 8516 2252
rect 8488 2230 8494 2250
rect 8548 2246 8764 2256
rect 8536 2238 8764 2246
rect 8536 2236 8738 2238
rect 8536 2218 8739 2236
rect 8598 2216 8714 2218
rect 8548 2166 8702 2216
rect 8598 2148 8652 2152
rect 8548 2126 8702 2148
rect 7514 2032 7532 2060
rect 7542 2038 7544 2104
rect 8536 2098 8744 2126
rect 8544 2096 8714 2098
rect 8488 2064 8494 2084
rect 8548 2072 8702 2096
rect 8714 2078 8739 2096
rect 8714 2076 8738 2078
rect 8714 2074 8764 2076
rect 8714 2072 8772 2074
rect 8484 2062 8516 2064
rect 8484 2056 8522 2062
rect 8548 2058 8772 2072
rect 8548 2056 8598 2058
rect 8484 2046 8598 2056
rect 8484 2014 8550 2046
rect 8484 1998 8516 2014
rect 8518 2004 8550 2014
rect 8574 2012 8584 2046
rect 8608 2025 8618 2056
rect 8574 2004 8582 2012
rect 8598 2010 8618 2025
rect 8630 2010 8648 2056
rect 8660 2036 8776 2058
rect 8664 2018 8682 2028
rect 8714 2026 8776 2036
rect 8598 2003 8652 2010
rect 8660 2003 8776 2018
rect 8598 1988 8776 2003
rect 8618 1980 8652 1988
rect 8660 1964 8714 1988
rect 3000 1896 3028 1932
rect 8364 1924 8620 1964
rect 8660 1963 8776 1964
rect 8660 1962 8725 1963
rect 8664 1960 8702 1962
rect 8648 1940 8702 1944
rect 8704 1942 8736 1962
rect 8704 1940 8772 1942
rect 8648 1926 8772 1940
rect 8364 1902 8628 1924
rect 8648 1902 8652 1922
rect 8660 1902 8694 1926
rect 7570 1872 7680 1894
rect 8364 1892 8694 1902
rect 8714 1892 8776 1926
rect 7542 1844 7708 1866
rect 8364 1856 8688 1892
rect 8364 1838 8620 1856
rect 8648 1842 8714 1856
rect 8362 1834 8620 1838
rect 3530 1798 3576 1826
rect 7402 1796 7440 1824
rect 7490 1796 7546 1824
rect 8362 1796 8416 1834
rect 8830 1796 8874 2088
rect 7410 1768 7474 1792
rect 8996 1754 9014 1770
rect 9024 1754 9058 1788
rect 8996 1720 9008 1754
rect 9030 1720 9046 1736
rect 9030 1702 9042 1720
rect 7594 1652 7684 1678
rect 7326 1556 7698 1652
rect 7326 1510 7762 1556
rect 7326 1498 7698 1510
rect 7530 1478 7554 1498
rect 7564 1478 7620 1498
rect 7564 1464 7588 1478
rect 7598 1472 7620 1478
rect 7538 1450 7554 1464
rect 7510 1426 7528 1448
rect 7564 1444 7572 1464
rect 7626 1444 7648 1498
rect 7626 1394 7668 1416
rect 7642 1374 7688 1388
rect 7618 1366 7688 1374
rect 7618 1358 7668 1366
rect 7642 1342 7648 1358
rect 7642 1330 7688 1342
rect 8052 610 8424 852
<< nwell >>
rect 3000 3004 3662 3006
rect 7594 3004 7862 3006
rect 3040 2942 3104 3002
rect 7494 2942 7558 3002
rect 8364 2970 8620 3006
rect 8364 1796 8620 1834
<< metal1 >>
rect 3072 3002 3104 3006
rect 3040 2998 3104 3002
rect 3040 2946 3046 2998
rect 3098 2946 3104 2998
rect 3154 2994 3192 3006
rect 3528 2984 3570 3006
rect 3622 2990 3660 3006
rect 3704 2994 3746 3006
rect 3920 2992 3956 3006
rect 5152 2976 5236 3006
rect 5358 2976 5442 3006
rect 6098 2990 6144 3006
rect 7402 2990 7440 3006
rect 7490 3002 7546 3006
rect 7490 2998 7558 3002
rect 7490 2990 7500 2998
rect 5152 2948 5442 2976
rect 3040 2942 3104 2946
rect 7494 2946 7500 2990
rect 7552 2946 7558 2998
rect 8228 2978 8296 3006
rect 8360 2976 8416 3006
rect 7494 2942 7558 2946
rect 7922 1892 7986 1896
rect 4684 1862 4748 1866
rect 3530 1798 3576 1822
rect 4684 1810 4690 1862
rect 4742 1810 4748 1862
rect 4684 1806 4748 1810
rect 5844 1862 5908 1866
rect 5844 1810 5850 1862
rect 5902 1810 5908 1862
rect 7922 1840 7928 1892
rect 7980 1840 7986 1892
rect 7922 1836 7986 1840
rect 7922 1830 8008 1836
rect 8128 1834 8230 1836
rect 8128 1830 8296 1834
rect 7922 1824 8296 1830
rect 7952 1814 8296 1824
rect 5844 1806 5908 1810
rect 7958 1808 8296 1814
rect 7402 1796 7440 1806
rect 7490 1796 7546 1806
rect 7964 1804 8296 1808
rect 7978 1802 8170 1804
rect 8228 1796 8296 1804
rect 8362 1796 8416 1838
<< via1 >>
rect 3046 2946 3098 2998
rect 7500 2946 7552 2998
rect 4690 1810 4742 1862
rect 5850 1810 5902 1862
rect 7928 1840 7980 1892
<< metal2 >>
rect 3040 2998 3104 3002
rect 3040 2946 3046 2998
rect 3098 2978 3104 2998
rect 7494 2998 7558 3002
rect 7494 2978 7500 2998
rect 3098 2946 7500 2978
rect 7552 2946 7558 2998
rect 7714 2952 7776 3000
rect 3040 2942 7558 2946
rect 3000 2870 3016 2906
rect 7936 2826 7980 2830
rect 7926 2758 7980 2826
rect 7578 2658 7648 2702
rect 7940 2644 7980 2646
rect 5302 2560 6900 2600
rect 7940 2578 7984 2644
rect 7944 2576 7984 2578
rect 6620 2424 6664 2426
rect 5304 2374 6670 2424
rect 6856 2416 6900 2560
rect 7730 2418 7794 2466
rect 8598 2464 8620 2510
rect 5304 2190 6006 2228
rect 5960 2070 6006 2190
rect 6612 2140 6670 2374
rect 6850 2408 6900 2416
rect 6850 2280 6902 2408
rect 8598 2300 8620 2344
rect 6850 2238 7676 2280
rect 7634 2210 7676 2238
rect 7634 2168 8036 2210
rect 6612 2096 7190 2140
rect 6612 2094 6670 2096
rect 5960 2040 6004 2070
rect 6834 2040 8034 2050
rect 5960 2010 8034 2040
rect 5960 2008 8008 2010
rect 5960 1996 6912 2008
rect 3000 1896 3016 1932
rect 7922 1892 7986 1896
rect 7922 1866 7928 1892
rect 4684 1862 7928 1866
rect 4684 1810 4690 1862
rect 4742 1836 5850 1862
rect 4742 1810 4748 1836
rect 4684 1806 4748 1810
rect 5844 1810 5850 1836
rect 5902 1840 7928 1862
rect 7980 1840 7986 1892
rect 5902 1836 7986 1840
rect 5902 1810 5908 1836
rect 5844 1806 5908 1810
use sky130_hilas_FGtrans2x1cell  sky130_hilas_FGtrans2x1cell_0
timestamp 1632256330
transform -1 0 4514 0 1 2560
box 0 0 4514 2104
use sky130_hilas_FGBias2x1cell  sky130_hilas_FGBias2x1cell_0
timestamp 1632256332
transform 1 0 6080 0 1 2560
box 0 0 3308 2104
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1632256331
transform 1 0 8310 0 1 1878
box 0 0 716 1504
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1632255311
transform 1 0 7326 0 -1 2126
box 0 0 1098 2126
<< labels >>
rlabel metal1 8228 2994 8296 3006 0 VGND
port 11 nsew
rlabel metal1 8360 2994 8416 3006 0 VPWR
port 10 nsew
rlabel metal1 8362 1796 8416 1808 0 VPWR
port 10 nsew
rlabel metal1 8228 1796 8296 1808 0 VGND
port 11 nsew
rlabel metal2 7730 2418 7794 2466 0 VIN21
port 9 nsew
rlabel metal2 7714 2952 7776 3000 1 VIN22
port 8 n
rlabel metal1 3530 1798 3576 1822 0 VIN12
port 18 nsew
rlabel metal1 3528 2984 3570 3006 0 VIN11
port 5 nsew
rlabel metal1 5358 2992 5442 3006 0 VTUN
port 1 nsew
rlabel metal1 5152 2992 5236 3006 0 VTUN
rlabel metal1 3704 2994 3746 3006 0 PROG
port 3 nsew
rlabel metal1 3072 2994 3104 3006 0 VINJ
port 6 nsew
rlabel metal1 7490 2990 7546 3006 0 VINJ
port 6 nsew
rlabel metal2 8598 2464 8620 2510 0 OUTPUT1
port 13 nsew
rlabel metal2 8598 2300 8620 2344 0 OUTPUT2
port 12 nsew
rlabel metal1 3154 2994 3192 3006 0 GATESEL1
port 14 nsew
rlabel metal1 7402 1796 7440 1806 0 GATESEL2
port 15 nsew
rlabel metal1 7490 1796 7546 1806 0 VINJ
port 6 nsew
rlabel metal1 7402 2990 7440 3006 0 GATESEL2
port 15 nsew
rlabel metal2 3000 2870 3016 2906 0 DRAIN1
port 16 nsew
rlabel metal2 3000 1896 3016 1932 0 DRAIN2
port 17 nsew
rlabel metal1 6098 2990 6144 3006 0 GATE1
port 4 nsew
rlabel metal1 3622 2990 3660 3006 0 GATE2
port 19 nsew
rlabel metal1 3920 2992 3956 3006 0 RUN
port 20 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
