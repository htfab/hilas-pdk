magic
tech sky130A
timestamp 1628166556
<< error_s >>
rect -937 590 -887 596
rect -865 590 -815 596
rect 819 590 869 596
rect 891 590 941 596
rect -942 579 -788 582
rect -757 579 761 582
rect 792 579 956 582
rect -743 569 725 579
rect -942 565 -788 568
rect -757 565 761 568
rect 792 565 956 568
rect -757 555 739 565
rect -937 548 -887 554
rect -865 548 -815 554
rect 819 548 869 554
rect 891 548 941 554
rect 1008 539 1013 564
rect -1004 533 -990 539
rect 999 533 1013 539
rect -1004 519 -976 525
rect -865 521 -815 527
rect 819 521 869 527
rect 985 521 1008 525
rect 985 519 1013 521
rect 1008 490 1013 519
rect -865 479 -815 485
rect 819 479 869 485
rect -865 436 -815 442
rect 819 436 869 442
rect 1008 408 1010 410
rect -865 394 -815 400
rect 819 394 869 400
rect 1009 390 1010 408
rect -937 367 -887 373
rect -865 367 -815 373
rect 819 367 869 373
rect 891 367 941 373
rect -1005 353 -1004 367
rect 1008 365 1009 367
rect -991 347 -990 353
rect -937 325 -887 331
rect -865 325 -815 331
rect 819 325 869 331
rect 891 325 941 331
rect -937 266 -887 272
rect -865 266 -815 272
rect 819 266 869 272
rect 891 266 941 272
rect -997 244 -990 250
rect 994 244 1000 246
rect 1009 244 1014 250
rect -937 224 -887 230
rect -865 224 -815 230
rect 819 224 869 230
rect 891 224 941 230
rect -997 201 -990 207
rect -865 197 -815 203
rect 819 197 869 203
rect 994 201 1000 203
rect 1009 201 1014 207
rect -865 155 -815 161
rect 819 155 869 161
rect -865 113 -815 119
rect 819 113 869 119
rect -997 91 -990 108
rect 994 91 1000 104
rect 1009 91 1014 108
rect -1004 73 -983 79
rect -865 71 -815 77
rect 819 71 869 77
rect 986 73 1008 79
rect -1004 59 -990 65
rect 1000 61 1014 65
rect -997 48 -990 59
rect 994 59 1014 61
rect -937 44 -887 50
rect -865 44 -815 50
rect 819 44 869 50
rect 891 44 941 50
rect 994 48 1000 59
rect 1009 48 1014 59
rect -937 2 -887 8
rect -865 2 -815 8
rect 819 2 869 8
rect 891 2 941 8
<< metal1 >>
rect -968 597 -952 601
rect -984 595 -952 597
rect -927 596 -908 601
rect -887 596 -871 601
rect -984 569 -981 595
rect -955 569 -952 595
rect -693 592 -669 601
rect -475 591 -437 601
rect -300 595 -276 601
rect -72 588 -32 601
rect 36 591 76 601
rect 280 596 304 601
rect 441 591 479 601
rect 673 594 697 601
rect 875 596 891 601
rect 912 596 931 601
rect 956 597 972 601
rect 956 595 988 597
rect -984 567 -952 569
rect -32 565 36 587
rect 956 569 959 595
rect 985 569 988 595
rect 956 567 988 569
rect -968 -4 -952 2
rect -927 -3 -908 3
rect -887 -3 -871 3
rect -693 -4 -669 4
rect -475 -4 -437 5
rect -300 -4 -276 3
rect -72 -4 -32 8
rect 36 -4 76 8
rect 280 -4 304 3
rect 441 -4 479 11
rect 673 -4 697 2
rect 875 -3 891 3
rect 912 -3 931 3
rect 956 -3 972 3
<< via1 >>
rect -981 569 -955 595
rect 959 569 985 595
<< metal2 >>
rect -984 595 -699 597
rect -984 569 -981 595
rect -955 587 -699 595
rect 705 595 988 597
rect 705 587 959 595
rect -955 579 959 587
rect -955 569 -942 579
rect -743 569 725 579
rect 956 569 959 579
rect 985 569 988 595
rect -984 567 -942 569
rect 956 567 988 569
rect -1004 533 -990 552
rect 999 533 1008 551
rect -1004 490 -990 509
rect 999 490 1008 508
rect -1004 390 -989 409
rect 996 390 1009 408
rect -1004 347 -991 365
rect 995 347 1009 365
rect -1004 232 -997 250
rect 1000 232 1009 250
rect -1004 189 -997 207
rect 1000 189 1009 207
rect -334 134 342 152
rect -1004 90 -997 108
rect 1000 90 1009 108
rect -1004 47 -997 65
rect 1000 47 1009 65
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_0
timestamp 1628166556
transform 1 0 264 0 1 378
box -263 -404 744 246
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_1
timestamp 1628166556
transform -1 0 -260 0 1 378
box -263 -404 744 246
<< labels >>
rlabel metal1 441 591 479 601 0 GATE2
port 1 nsew analog default
rlabel metal1 -72 -4 -32 8 0 VTUN
port 2 nsew power default
rlabel metal1 36 -4 76 8 0 VTUN
port 2 nsew power default
rlabel metal1 36 591 76 601 0 VTUN
port 2 nsew power default
rlabel metal1 -72 588 -32 601 0 VTUN
port 2 nsew power default
rlabel metal1 -475 591 -437 601 0 GATE1
port 3 nsew analog default
rlabel metal1 -475 -4 -437 5 0 GATE1
port 3 nsew analog default
rlabel metal1 956 -3 972 3 0 VINJ
port 4 nsew power default
rlabel metal1 441 -4 479 11 0 GATE2
port 1 nsew analog default
rlabel metal1 912 596 931 601 0 SelectGate2
rlabel metal1 956 596 972 601 0 VINJ
port 6 nsew power default
rlabel metal1 -968 596 -952 601 0 VINJ
port 6 nsew power default
rlabel metal1 -927 596 -908 601 0 GATESELECT1
port 10 nsew analog default
rlabel metal1 -968 -4 -952 2 0 VINJ
port 6 nsew power default
rlabel metal1 -927 -3 -908 3 0 GATESELECT1
port 10 nsew analog default
rlabel metal1 -887 596 -871 601 0 COL1
port 12 nsew analog default
rlabel metal1 -887 -3 -871 3 0 COL1
port 12 nsew analog default
rlabel metal1 912 -3 931 3 0 GATESELECT2
port 11 nsew analog default
rlabel metal1 875 -3 891 3 0 COL2
port 13 nsew analog default
rlabel metal1 875 596 891 601 0 COL2
port 13 nsew analog default
rlabel metal2 -1004 490 -997 509 0 ROW1
port 14 nsew analog default
rlabel metal2 -1004 390 -997 409 0 ROW2
port 15 nsew analog default
rlabel metal2 -1004 533 -997 552 0 DRAIN1
port 16 nsew analog default
rlabel metal2 -1004 347 -997 365 0 DRAIN2
port 17 nsew analog default
rlabel metal2 -1004 232 -997 250 0 DRAIN3
port 18 nsew analog default
rlabel metal2 -1004 189 -997 207 0 ROW3
port 19 nsew analog default
rlabel metal2 -1004 90 -997 108 0 ROW4
port 20 nsew analog default
rlabel metal2 -1004 47 -997 65 0 DRAIN4
port 21 nsew analog default
rlabel metal2 999 533 1008 551 0 DRAIN1
port 16 nsew analog default
rlabel metal2 999 490 1008 508 0 ROW1
port 14 nsew analog default
rlabel metal2 1000 390 1009 408 0 ROW2
port 15 nsew
rlabel metal2 1000 347 1009 365 0 DRAIN2
port 17 nsew analog default
rlabel metal2 1000 232 1009 250 0 DRAIN3
port 18 nsew analog default
rlabel metal2 1000 189 1009 207 0 ROW3
port 19 nsew analog default
rlabel metal2 1000 90 1009 108 0 ROW4
port 20 nsew analog default
rlabel metal2 1000 47 1009 65 0 DRAIN4
port 21 nsew
rlabel metal1 -693 595 -669 601 0 VGND
port 22 nsew
rlabel metal1 -693 -4 -669 4 0 VGND
port 22 nsew
rlabel metal1 -300 -4 -276 3 0 VGND
port 22 nsew
rlabel metal1 -300 595 -276 601 0 VGND
port 22 nsew
rlabel metal1 280 -4 304 3 0 VGND
port 22 nsew
rlabel metal1 673 -4 697 2 0 VGND
port 22 nsew
rlabel metal1 280 596 304 601 0 VGND
port 22 nsew
rlabel metal1 673 594 697 601 0 VGND
port 22 nsew
<< end >>
