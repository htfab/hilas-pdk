magic
tech sky130A
timestamp 1627400660
<< nwell >>
rect 210 63 264 309
rect 192 18 264 63
rect 7 0 264 18
<< psubdiff >>
rect 206 518 248 525
rect 206 501 219 518
rect 236 501 248 518
rect 206 494 248 501
<< nsubdiff >>
rect 205 40 246 45
rect 205 23 217 40
rect 234 23 246 40
rect 205 18 246 23
<< psubdiffcont >>
rect 219 501 236 518
<< nsubdiffcont >>
rect 217 23 234 40
<< locali >>
rect 220 526 237 531
rect 219 523 237 526
rect 219 518 262 523
rect 236 501 262 518
rect 219 498 262 501
rect 219 492 236 498
rect 205 23 217 40
rect 234 23 247 40
<< metal1 >>
rect 218 0 240 588
rect 258 0 280 588
<< metal2 >>
rect 0 548 7 565
rect 198 549 280 566
rect 0 507 7 524
rect 0 456 7 473
rect 198 457 280 474
rect 0 415 7 432
rect 0 364 7 381
rect 198 365 280 382
rect 0 323 7 340
rect 0 262 7 281
rect 200 255 280 275
rect 0 220 7 239
rect 0 166 7 185
rect 200 159 280 179
rect 0 124 7 143
rect 0 70 7 89
rect 199 63 280 83
rect 0 28 7 47
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1607179295
transform 1 0 267 0 1 504
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1607179295
transform 0 1 220 -1 0 30
box -10 -8 13 21
use sky130_hilas_pFETdevice01e  sky130_hilas_pFETdevice01e_0
timestamp 1608055794
transform 1 0 128 0 1 265
box -121 -55 82 44
use sky130_hilas_pFETdevice01e  sky130_hilas_pFETdevice01e_1
timestamp 1608055794
transform 1 0 128 0 1 169
box -121 -55 82 44
use sky130_hilas_pFETdevice01e  sky130_hilas_pFETdevice01e_2
timestamp 1608055794
transform 1 0 128 0 1 73
box -121 -55 82 44
use sky130_hilas_nFET03a  sky130_hilas_nFET03a_0
timestamp 1608056777
transform 1 0 118 0 1 362
box -111 -47 97 42
use sky130_hilas_nFET03a  sky130_hilas_nFET03a_1
timestamp 1608056777
transform 1 0 118 0 1 454
box -111 -47 97 42
use sky130_hilas_nFET03a  sky130_hilas_nFET03a_3
timestamp 1608056777
transform 1 0 118 0 1 546
box -111 -47 97 42
<< labels >>
rlabel metal1 218 0 240 9 0 WELL
port 13 nsew power default
rlabel metal1 258 0 280 9 0 VGND
port 14 nsew ground default
rlabel metal1 218 579 240 588 0 WELL
port 13 nsew ground default
rlabel metal1 258 579 280 588 0 VGND
port 14 nsew power default
rlabel metal2 0 548 7 565 0 NFET_SOURCE1
port 1 nsew analog default
rlabel metal2 0 507 7 524 0 NFET_GATE1
port 2 nsew analog default
rlabel metal2 0 456 7 473 0 NFET_SOURCE2
port 3 nsew analog default
rlabel metal2 0 415 7 432 0 NFET_GATE2
port 4 nsew analog default
rlabel metal2 0 364 7 381 0 NFET_SOURCE3
port 5 nsew analog default
rlabel metal2 0 323 7 340 0 NFET_GATE3
port 6 nsew analog default
rlabel metal2 0 220 7 239 0 PFET_GATE1
port 8 nsew analog default
rlabel metal2 0 262 7 281 0 PFET_SOURCE1
port 7 nsew analog default
rlabel metal2 0 166 7 185 0 PFET_SOURCE2
port 9 nsew analog default
rlabel metal2 0 124 7 143 0 PFET_GATE2
port 10 nsew analog default
rlabel metal2 0 70 7 89 0 PFET_SOURCE3
port 11 nsew analog default
rlabel metal2 0 28 7 47 0 PFET_GATE3
port 12 nsew analog default
rlabel metal2 274 255 280 275 0 PFET_DRAIN1
port 17 nsew analog default
rlabel metal2 274 159 280 179 0 PFET_DRAIN2
port 16 nsew analog default
rlabel metal2 274 63 280 83 0 PFET_DRAIN3
port 15 nsew analog default
rlabel metal2 275 549 280 566 0 NFET_DRAIN1
port 20 nsew analog default
rlabel metal2 275 457 280 474 0 NFET_DRAIN2
port 19 nsew analog default
rlabel metal2 275 365 280 382 0 NFET_DRAIN3
port 18 nsew analog default
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
