magic
tech sky130A
timestamp 1628704386
<< checkpaint >>
rect -544 -629 749 658
<< nwell >>
rect 0 0 128 284
<< pmos >>
rect 21 206 89 236
rect 21 75 89 105
<< pdiff >>
rect 21 260 89 265
rect 21 242 28 260
rect 46 242 64 260
rect 82 242 89 260
rect 21 236 89 242
rect 21 200 89 206
rect 21 182 29 200
rect 46 182 65 200
rect 83 182 89 200
rect 21 176 89 182
rect 21 129 89 135
rect 21 112 29 129
rect 47 112 65 129
rect 83 112 89 129
rect 21 105 89 112
rect 21 68 89 75
rect 21 51 29 68
rect 47 51 65 68
rect 83 51 89 68
rect 21 47 89 51
<< pdiffc >>
rect 28 242 46 260
rect 64 242 82 260
rect 29 182 46 200
rect 65 182 83 200
rect 29 112 47 129
rect 65 112 83 129
rect 29 51 47 68
rect 65 51 83 68
<< nsubdiff >>
rect 21 164 89 176
rect 21 147 29 164
rect 47 147 65 164
rect 83 147 89 164
rect 21 135 89 147
<< nsubdiffcont >>
rect 29 147 47 164
rect 65 147 83 164
<< poly >>
rect 8 206 21 236
rect 89 206 114 236
rect 97 105 114 206
rect 8 75 21 105
rect 89 75 114 105
rect 97 23 114 75
<< locali >>
rect 20 242 28 260
rect 46 242 64 260
rect 82 242 90 260
rect 21 182 29 200
rect 46 182 65 200
rect 83 182 91 200
rect 21 164 91 182
rect 21 147 29 164
rect 47 147 65 164
rect 83 147 91 164
rect 21 129 91 147
rect 21 112 29 129
rect 47 112 65 129
rect 83 112 91 129
rect 21 51 29 68
rect 47 51 65 68
rect 83 51 92 68
rect 56 23 92 51
rect 56 6 89 23
use sky130_hilas_poly2li  sky130_hilas_poly2li_0
timestamp 1628704338
transform 0 1 100 -1 0 19
box 0 0 27 33
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
