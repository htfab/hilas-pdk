magic
tech sky130A
timestamp 1628617048
<< checkpaint >>
rect -630 895 969 917
rect -630 -630 1116 895
rect -483 -652 1116 -630
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_3
timestamp 1628616750
transform 1 0 220 0 1 0
box 0 0 119 287
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_4
timestamp 1628616750
transform 1 0 0 0 1 0
box 0 0 119 287
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_0
timestamp 1628616750
transform 1 0 55 0 1 0
box 0 0 119 287
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_1
timestamp 1628616750
transform 1 0 110 0 1 0
box 0 0 119 287
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_2
timestamp 1628616750
transform 1 0 165 0 1 0
box 0 0 119 287
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
