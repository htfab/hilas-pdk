magic
tech sky130A
timestamp 1627744303
<< error_s >>
rect -626 12757 -597 12773
rect -547 12757 -518 12773
rect -468 12757 -439 12773
rect -389 12757 -360 12773
rect -502 12734 -485 12735
rect -626 12723 -625 12724
rect -598 12723 -597 12724
rect -547 12723 -546 12724
rect -519 12723 -518 12724
rect -468 12723 -467 12724
rect -440 12723 -439 12724
rect -389 12723 -388 12724
rect -361 12723 -360 12724
rect -676 12694 -659 12723
rect -627 12722 -596 12723
rect -548 12722 -517 12723
rect -469 12722 -438 12723
rect -390 12722 -359 12723
rect -626 12715 -597 12722
rect -547 12715 -518 12722
rect -502 12715 -485 12716
rect -468 12715 -439 12722
rect -389 12715 -360 12722
rect -626 12701 -617 12715
rect -370 12701 -360 12715
rect -626 12695 -597 12701
rect -547 12695 -518 12701
rect -502 12699 -485 12701
rect -468 12695 -439 12701
rect -389 12695 -360 12701
rect -627 12694 -596 12695
rect -548 12694 -517 12695
rect -469 12694 -438 12695
rect -390 12694 -359 12695
rect -328 12694 -310 12723
rect -626 12693 -625 12694
rect -598 12693 -597 12694
rect -547 12693 -546 12694
rect -519 12693 -518 12694
rect -468 12693 -467 12694
rect -440 12693 -439 12694
rect -389 12693 -388 12694
rect -361 12693 -360 12694
rect -502 12680 -485 12682
rect -626 12644 -597 12659
rect -547 12644 -518 12659
rect -468 12644 -439 12659
rect -389 12644 -360 12659
rect -553 12607 -514 12610
rect -553 12565 -514 12568
rect -626 12477 -597 12493
rect -547 12477 -518 12493
rect -468 12477 -439 12493
rect -389 12477 -360 12493
rect -502 12454 -485 12455
rect -626 12443 -625 12444
rect -598 12443 -597 12444
rect -547 12443 -546 12444
rect -519 12443 -518 12444
rect -468 12443 -467 12444
rect -440 12443 -439 12444
rect -389 12443 -388 12444
rect -361 12443 -360 12444
rect -676 12414 -659 12443
rect -627 12442 -596 12443
rect -548 12442 -517 12443
rect -469 12442 -438 12443
rect -390 12442 -359 12443
rect -626 12435 -597 12442
rect -547 12435 -518 12442
rect -502 12435 -485 12436
rect -468 12435 -439 12442
rect -389 12435 -360 12442
rect -626 12421 -617 12435
rect -370 12421 -360 12435
rect -626 12415 -597 12421
rect -547 12415 -518 12421
rect -502 12419 -485 12421
rect -468 12415 -439 12421
rect -389 12415 -360 12421
rect -627 12414 -596 12415
rect -548 12414 -517 12415
rect -469 12414 -438 12415
rect -390 12414 -359 12415
rect -328 12414 -310 12443
rect -626 12413 -625 12414
rect -598 12413 -597 12414
rect -547 12413 -546 12414
rect -519 12413 -518 12414
rect -468 12413 -467 12414
rect -440 12413 -439 12414
rect -389 12413 -388 12414
rect -361 12413 -360 12414
rect -502 12400 -485 12402
rect 470 12395 499 12413
rect -626 12364 -597 12379
rect -547 12364 -518 12379
rect -468 12364 -439 12379
rect -389 12364 -360 12379
rect 470 12363 471 12364
rect 498 12363 499 12364
rect -626 12322 -597 12338
rect -547 12322 -518 12338
rect -468 12322 -439 12338
rect -389 12322 -360 12338
rect 420 12334 438 12363
rect 469 12362 500 12363
rect 470 12353 499 12362
rect 470 12344 480 12353
rect 489 12344 499 12353
rect 470 12335 499 12344
rect 469 12334 500 12335
rect 531 12334 549 12363
rect 470 12333 471 12334
rect 498 12333 499 12334
rect -502 12299 -485 12300
rect -626 12288 -625 12289
rect -598 12288 -597 12289
rect -547 12288 -546 12289
rect -519 12288 -518 12289
rect -468 12288 -467 12289
rect -440 12288 -439 12289
rect -389 12288 -388 12289
rect -361 12288 -360 12289
rect -676 12259 -659 12288
rect -627 12287 -596 12288
rect -548 12287 -517 12288
rect -469 12287 -438 12288
rect -390 12287 -359 12288
rect -626 12280 -597 12287
rect -547 12280 -518 12287
rect -502 12280 -485 12281
rect -468 12280 -439 12287
rect -389 12280 -360 12287
rect -626 12266 -617 12280
rect -370 12266 -360 12280
rect -626 12260 -597 12266
rect -547 12260 -518 12266
rect -502 12264 -485 12266
rect -468 12260 -439 12266
rect -389 12260 -360 12266
rect -627 12259 -596 12260
rect -548 12259 -517 12260
rect -469 12259 -438 12260
rect -390 12259 -359 12260
rect -328 12259 -310 12288
rect 470 12284 499 12302
rect -626 12258 -625 12259
rect -598 12258 -597 12259
rect -547 12258 -546 12259
rect -519 12258 -518 12259
rect -468 12258 -467 12259
rect -440 12258 -439 12259
rect -389 12258 -388 12259
rect -361 12258 -360 12259
rect -502 12245 -485 12247
rect -626 12209 -597 12224
rect -547 12209 -518 12224
rect -468 12209 -439 12224
rect -389 12209 -360 12224
rect 1242 11570 1270 11586
rect 1384 11570 1412 11586
rect 1519 11576 1569 11585
rect 1852 11579 1902 11590
rect 1488 11570 1519 11576
rect 1818 11573 1852 11579
rect 1296 11544 1301 11549
rect 1242 11528 1270 11544
rect 1384 11528 1412 11544
rect 1519 11534 1569 11543
rect 1736 11536 1753 11541
rect 1852 11537 1902 11548
rect 1909 11528 1926 11529
rect 1193 11507 1221 11524
rect 1433 11507 1461 11524
rect 1590 11508 1641 11518
rect 1781 11517 1831 11528
rect 1909 11509 1926 11510
rect 1654 11503 1673 11508
rect 1193 11465 1221 11482
rect 1433 11465 1461 11482
rect 1559 11476 1590 11482
rect 1668 11476 1673 11503
rect 1749 11486 1781 11491
rect 1590 11466 1641 11476
rect 1781 11475 1831 11486
rect 1242 11415 1270 11431
rect 1384 11415 1412 11431
rect 1519 11421 1569 11430
rect 1852 11424 1902 11435
rect 1488 11415 1519 11421
rect 1818 11418 1852 11424
rect 1296 11389 1301 11394
rect 1242 11373 1270 11389
rect 1384 11373 1412 11389
rect 1519 11379 1569 11388
rect 1736 11381 1753 11386
rect 1852 11382 1902 11393
rect 1909 11373 1926 11374
rect 1193 11352 1221 11369
rect 1433 11352 1461 11369
rect 1590 11353 1641 11363
rect 1781 11362 1831 11373
rect 1909 11354 1926 11355
rect 1654 11348 1673 11353
rect -943 11308 -916 11315
rect 1193 11310 1221 11327
rect 1433 11310 1461 11327
rect 1559 11321 1590 11327
rect 1668 11321 1673 11348
rect 1749 11331 1781 11336
rect 1590 11311 1641 11321
rect 1781 11320 1831 11331
rect -943 11266 -916 11273
rect 1242 11260 1270 11276
rect 1384 11260 1412 11276
rect 1519 11266 1569 11275
rect 1852 11269 1902 11280
rect 2696 11271 2746 11282
rect 2768 11271 2818 11282
rect 4737 11271 4787 11282
rect 4809 11271 4859 11282
rect 5197 11277 5224 11284
rect 1488 11260 1519 11266
rect 1818 11263 1852 11269
rect 5400 11264 5417 11269
rect 2818 11240 2852 11241
rect 4703 11240 4737 11241
rect 1296 11234 1301 11239
rect -943 11216 -916 11223
rect 1242 11218 1270 11234
rect 1384 11218 1412 11234
rect 1519 11224 1569 11233
rect 1736 11226 1753 11231
rect 1852 11227 1902 11238
rect 2696 11229 2746 11240
rect 2768 11229 2818 11240
rect 4737 11229 4787 11240
rect 4809 11229 4859 11240
rect 5197 11235 5224 11242
rect 1909 11218 1926 11219
rect 1193 11197 1221 11214
rect 1433 11197 1461 11214
rect 1590 11198 1641 11208
rect 1781 11207 1831 11218
rect 5197 11211 5224 11218
rect 2760 11208 2769 11210
rect 2820 11208 2852 11210
rect 2884 11208 2923 11210
rect 3019 11208 3059 11210
rect 4496 11208 4536 11210
rect 4632 11208 4671 11210
rect 4703 11208 4735 11210
rect 4786 11208 4795 11210
rect 1909 11199 1926 11200
rect 1654 11193 1673 11198
rect -943 11174 -916 11181
rect 1193 11155 1221 11172
rect 1433 11155 1461 11172
rect 1559 11166 1590 11172
rect 1668 11166 1673 11193
rect 1749 11176 1781 11181
rect 1590 11156 1641 11166
rect 1781 11165 1831 11176
rect -943 11124 -916 11131
rect 1242 11105 1270 11121
rect 1384 11105 1412 11121
rect 1519 11111 1569 11120
rect 1852 11114 1902 11125
rect 1488 11105 1519 11111
rect 1818 11108 1852 11114
rect 2741 11104 2746 11145
rect 2881 11133 2884 11183
rect 2923 11133 2926 11183
rect 3017 11133 3019 11183
rect 3059 11133 3061 11183
rect 4494 11133 4496 11183
rect 4536 11133 4538 11183
rect 4629 11133 4632 11183
rect 4671 11133 4674 11183
rect 5197 11169 5224 11176
rect 4809 11121 4814 11145
rect 5197 11129 5224 11136
rect 4833 11104 4838 11121
rect -943 11082 -916 11089
rect 1296 11079 1301 11084
rect 1242 11063 1270 11079
rect 1384 11063 1412 11079
rect 1519 11069 1569 11078
rect 1736 11071 1753 11076
rect 1852 11072 1902 11083
rect 1909 11063 1926 11064
rect 1193 11042 1221 11059
rect 1433 11042 1461 11059
rect 1590 11043 1641 11053
rect 1781 11052 1831 11063
rect 2881 11054 2884 11104
rect 2923 11054 2926 11104
rect 3017 11054 3019 11104
rect 3059 11054 3061 11104
rect 4494 11054 4496 11104
rect 4536 11054 4538 11104
rect 4629 11054 4632 11104
rect 4671 11054 4674 11104
rect 5197 11087 5224 11094
rect 5197 11063 5224 11070
rect 1909 11044 1926 11045
rect 1654 11038 1673 11043
rect -951 11018 -912 11021
rect 1193 11000 1221 11017
rect 1433 11000 1461 11017
rect 1559 11011 1590 11017
rect 1668 11011 1673 11038
rect 1749 11021 1781 11026
rect 5197 11021 5224 11028
rect 1590 11001 1641 11011
rect 1781 11010 1831 11021
rect 7955 11011 7995 11022
rect 8105 11011 8145 11022
rect 5197 10981 5224 10988
rect -951 10976 -912 10979
rect 7955 10969 7995 10980
rect 8105 10969 8145 10980
rect 1193 10950 1221 10967
rect 1433 10950 1461 10967
rect 1590 10956 1641 10966
rect 1559 10950 1590 10956
rect 1668 10929 1673 10956
rect 1781 10946 1831 10957
rect 1749 10941 1781 10946
rect 2106 10931 2156 10942
rect 2286 10931 2336 10942
rect 2426 10931 2476 10941
rect -951 10922 -912 10925
rect 1193 10908 1221 10925
rect 1320 10907 1325 10912
rect 1433 10908 1461 10925
rect 1654 10924 1673 10929
rect 1590 10914 1641 10924
rect 1909 10922 1926 10923
rect 1749 10915 1777 10920
rect 2522 10919 2539 10921
rect 1781 10904 1831 10915
rect 1242 10888 1270 10904
rect 1384 10888 1412 10904
rect 1909 10903 1926 10904
rect 2336 10900 2366 10904
rect 1519 10889 1569 10898
rect 1852 10884 1902 10895
rect 2106 10889 2156 10900
rect 2286 10889 2336 10900
rect 2396 10899 2401 10904
rect 2522 10900 2539 10902
rect 2426 10889 2476 10899
rect 2522 10885 2539 10887
rect 2741 10884 2746 10925
rect 2881 10901 2884 10951
rect 2923 10901 2926 10951
rect 3017 10901 3019 10951
rect 3059 10901 3061 10951
rect 4494 10901 4496 10951
rect 4536 10901 4538 10951
rect 4629 10901 4632 10951
rect 4671 10901 4674 10951
rect 7879 10950 7919 10960
rect 8105 10948 8145 10960
rect 5197 10939 5224 10946
rect 4809 10901 4814 10925
rect 5197 10915 5224 10922
rect 7879 10908 7919 10918
rect 8105 10906 8145 10918
rect 4833 10884 4838 10901
rect -951 10880 -912 10883
rect 2106 10869 2156 10880
rect 2372 10869 2377 10880
rect 2426 10869 2476 10880
rect 5197 10873 5224 10880
rect 2396 10863 2401 10869
rect 2522 10866 2539 10868
rect 1242 10846 1270 10862
rect 1384 10846 1412 10862
rect 1488 10856 1519 10862
rect 1519 10847 1569 10856
rect 1818 10853 1852 10859
rect 1852 10842 1902 10853
rect 2078 10838 2106 10844
rect 2156 10838 2184 10844
rect 2396 10838 2426 10844
rect -951 10826 -912 10829
rect 2106 10827 2156 10838
rect 2426 10827 2476 10838
rect 2881 10822 2884 10872
rect 2923 10822 2926 10872
rect 3017 10822 3019 10872
rect 3059 10822 3061 10872
rect 4494 10822 4496 10872
rect 4536 10822 4538 10872
rect 4629 10822 4632 10872
rect 4671 10822 4674 10872
rect 7879 10849 7919 10859
rect 8105 10849 8145 10861
rect 5197 10833 5224 10840
rect 1193 10795 1221 10812
rect 1433 10795 1461 10812
rect 1590 10801 1641 10811
rect 7879 10807 7919 10817
rect 8105 10807 8145 10819
rect 1559 10795 1590 10801
rect -951 10784 -912 10787
rect 1668 10774 1673 10801
rect 1781 10791 1831 10802
rect 2760 10795 2769 10797
rect 2820 10795 2852 10797
rect 2884 10795 2923 10797
rect 3019 10795 3059 10797
rect 4496 10795 4536 10797
rect 4632 10795 4671 10797
rect 4703 10795 4735 10797
rect 4786 10795 4795 10797
rect 5197 10791 5224 10798
rect 1749 10786 1781 10791
rect 2106 10778 2156 10789
rect 2426 10778 2476 10789
rect 7955 10787 7995 10798
rect 8105 10787 8145 10798
rect 1193 10753 1221 10770
rect 1320 10752 1325 10757
rect 1433 10753 1461 10770
rect 1654 10769 1673 10774
rect 2078 10772 2106 10778
rect 2156 10772 2184 10778
rect 2396 10772 2426 10778
rect 1590 10759 1641 10769
rect 1909 10767 1926 10768
rect 1749 10760 1777 10765
rect 1781 10749 1831 10760
rect 1242 10733 1270 10749
rect 1384 10733 1412 10749
rect 1909 10748 1926 10749
rect 2396 10747 2401 10772
rect 2696 10765 2746 10776
rect 2768 10765 2818 10776
rect 4737 10765 4787 10776
rect 4809 10765 4859 10776
rect 5197 10767 5224 10774
rect 2818 10764 2852 10765
rect 4703 10764 4737 10765
rect 5376 10761 5400 10766
rect 2522 10748 2539 10750
rect 1519 10734 1569 10743
rect 1852 10729 1902 10740
rect 2106 10736 2156 10747
rect 2372 10740 2377 10741
rect 2360 10736 2377 10740
rect 2426 10736 2476 10747
rect 7955 10745 7995 10756
rect 8105 10745 8145 10756
rect 2522 10729 2539 10731
rect 2106 10716 2156 10727
rect 2286 10716 2336 10727
rect 2426 10717 2476 10727
rect 2696 10723 2746 10734
rect 2768 10723 2818 10734
rect 4737 10723 4787 10734
rect 4809 10723 4859 10734
rect 5197 10725 5224 10732
rect 2522 10714 2539 10716
rect 7955 10709 7995 10720
rect 8105 10709 8145 10720
rect 1242 10691 1270 10707
rect 1384 10691 1412 10707
rect 1488 10701 1519 10707
rect 1519 10692 1569 10701
rect 1818 10698 1852 10704
rect 1852 10687 1902 10698
rect 2522 10695 2539 10697
rect 2106 10674 2156 10685
rect 2286 10674 2336 10685
rect 2426 10675 2476 10685
rect 2697 10668 2747 10679
rect 2769 10668 2819 10679
rect 4737 10668 4787 10679
rect 4809 10668 4859 10679
rect 5197 10674 5224 10681
rect 7955 10667 7995 10678
rect 8105 10667 8145 10678
rect 5400 10661 5417 10666
rect 1193 10640 1221 10657
rect 1433 10640 1461 10657
rect 1590 10646 1641 10656
rect 1559 10640 1590 10646
rect 1668 10619 1673 10646
rect 1781 10636 1831 10647
rect 2106 10638 2156 10649
rect 2286 10638 2336 10649
rect 7879 10648 7919 10658
rect 2426 10638 2476 10648
rect 8105 10646 8145 10658
rect 2819 10637 2853 10638
rect 4703 10637 4737 10638
rect 1749 10631 1781 10636
rect 2522 10626 2539 10628
rect 2697 10626 2747 10637
rect 2769 10626 2819 10637
rect 4737 10626 4787 10637
rect 4809 10626 4859 10637
rect 5197 10632 5224 10639
rect 1193 10598 1221 10615
rect 1320 10597 1325 10602
rect 1433 10598 1461 10615
rect 1654 10614 1673 10619
rect 1590 10604 1641 10614
rect 1909 10612 1926 10613
rect 1749 10605 1777 10610
rect 2336 10607 2366 10611
rect 1781 10594 1831 10605
rect 2106 10596 2156 10607
rect 2286 10596 2336 10607
rect 2396 10606 2401 10611
rect 2522 10607 2539 10609
rect 5197 10608 5224 10615
rect 2426 10596 2476 10606
rect 2761 10605 2770 10607
rect 2821 10605 2853 10607
rect 2885 10605 2924 10607
rect 3020 10605 3060 10607
rect 4496 10605 4536 10607
rect 4632 10605 4671 10607
rect 4703 10605 4735 10607
rect 4786 10605 4795 10607
rect 7879 10606 7919 10616
rect 3058 10597 3060 10605
rect 8105 10604 8145 10616
rect 1242 10578 1270 10594
rect 1384 10578 1412 10594
rect 1909 10593 1926 10594
rect 2522 10592 2539 10594
rect 1519 10579 1569 10588
rect 1852 10574 1902 10585
rect 2106 10576 2156 10587
rect 2372 10576 2377 10587
rect 2426 10576 2476 10587
rect 2396 10570 2401 10576
rect 2522 10573 2539 10575
rect 1242 10536 1270 10552
rect 1384 10536 1412 10552
rect 1488 10546 1519 10552
rect 1519 10537 1569 10546
rect 1818 10543 1852 10549
rect 2078 10545 2106 10551
rect 2156 10545 2184 10551
rect 2396 10545 2426 10551
rect 1852 10532 1902 10543
rect 2106 10534 2156 10545
rect 2426 10534 2476 10545
rect 1193 10485 1221 10502
rect 1433 10485 1461 10502
rect 2742 10501 2747 10542
rect 2882 10530 2885 10580
rect 2924 10530 2927 10580
rect 3018 10530 3020 10580
rect 3060 10530 3062 10580
rect 4494 10530 4496 10580
rect 4536 10530 4538 10580
rect 4629 10530 4632 10580
rect 4671 10530 4674 10580
rect 5197 10566 5224 10573
rect 7879 10547 7919 10557
rect 8105 10547 8145 10559
rect 4809 10518 4814 10542
rect 5197 10526 5224 10533
rect 4833 10501 4838 10518
rect 7879 10505 7919 10515
rect 8105 10505 8145 10517
rect 1590 10491 1641 10501
rect 1559 10485 1590 10491
rect 1668 10464 1673 10491
rect 1781 10481 1831 10492
rect 2106 10485 2156 10496
rect 2426 10485 2476 10496
rect 1749 10476 1781 10481
rect 2078 10479 2106 10485
rect 2156 10479 2184 10485
rect 2396 10479 2426 10485
rect 1193 10443 1221 10460
rect 1320 10442 1325 10447
rect 1433 10443 1461 10460
rect 1654 10459 1673 10464
rect 1590 10449 1641 10459
rect 1909 10457 1926 10458
rect 1749 10450 1777 10455
rect 2396 10454 2401 10479
rect 2522 10455 2539 10457
rect 1781 10439 1831 10450
rect 2106 10443 2156 10454
rect 2372 10447 2377 10448
rect 2360 10443 2377 10447
rect 2426 10443 2476 10454
rect 2882 10451 2885 10501
rect 2924 10451 2927 10501
rect 3018 10451 3020 10501
rect 3060 10451 3062 10501
rect 4494 10451 4496 10501
rect 4536 10451 4538 10501
rect 4629 10451 4632 10501
rect 4671 10451 4674 10501
rect 5197 10484 5224 10491
rect 7955 10485 7995 10496
rect 8105 10485 8145 10496
rect 5197 10460 5224 10467
rect 7955 10443 7995 10454
rect 8105 10443 8145 10454
rect 1242 10423 1270 10439
rect 1384 10423 1412 10439
rect 1909 10438 1926 10439
rect 2522 10436 2539 10438
rect 1519 10424 1569 10433
rect 1852 10419 1902 10430
rect 2106 10423 2156 10434
rect 2286 10423 2336 10434
rect 2426 10424 2476 10434
rect 2522 10421 2539 10423
rect 3480 10420 3497 10421
rect 4059 10420 4076 10421
rect 5197 10418 5224 10425
rect 2522 10402 2539 10404
rect 3480 10401 3497 10402
rect 4059 10401 4076 10402
rect 1242 10381 1270 10397
rect 1384 10381 1412 10397
rect 1488 10391 1519 10397
rect 1519 10382 1569 10391
rect 1818 10388 1852 10394
rect 1852 10377 1902 10388
rect 2106 10381 2156 10392
rect 2286 10381 2336 10392
rect 2426 10382 2476 10392
rect 3480 10385 3497 10387
rect 4059 10385 4076 10387
rect 5197 10378 5224 10385
rect 3481 10366 3498 10368
rect 4059 10366 4076 10368
rect 2742 10281 2747 10322
rect 2882 10298 2885 10348
rect 2924 10298 2927 10348
rect 3018 10298 3020 10348
rect 3060 10298 3062 10348
rect 4494 10298 4496 10348
rect 4536 10298 4538 10348
rect 4629 10298 4632 10348
rect 4671 10298 4674 10348
rect 5197 10336 5224 10343
rect 4809 10298 4814 10322
rect 5197 10312 5224 10319
rect 4833 10281 4838 10298
rect 5197 10270 5224 10277
rect 2882 10219 2885 10269
rect 2924 10219 2927 10269
rect 3018 10219 3020 10269
rect 3060 10219 3062 10269
rect 4494 10219 4496 10269
rect 4536 10219 4538 10269
rect 4629 10219 4632 10269
rect 4671 10219 4674 10269
rect 5197 10230 5224 10237
rect 2761 10192 2770 10194
rect 2821 10192 2853 10194
rect 2885 10192 2924 10194
rect 3020 10192 3060 10194
rect 4496 10192 4536 10194
rect 4632 10192 4671 10194
rect 4703 10192 4735 10194
rect 4786 10192 4795 10194
rect 5197 10188 5224 10195
rect 2697 10162 2747 10173
rect 2769 10162 2819 10173
rect 4737 10162 4787 10173
rect 4809 10162 4859 10173
rect 5197 10164 5224 10171
rect 2819 10161 2853 10162
rect 4703 10161 4737 10162
rect 5376 10158 5400 10163
rect 2697 10120 2747 10131
rect 2769 10120 2819 10131
rect 4737 10120 4787 10131
rect 4809 10120 4859 10131
rect 5197 10122 5224 10129
rect 1193 9937 1221 9954
rect 1433 9937 1461 9954
rect 1590 9943 1641 9953
rect 1559 9937 1590 9943
rect 1668 9916 1673 9943
rect 1781 9933 1831 9944
rect 1749 9928 1781 9933
rect 2106 9924 2156 9935
rect 2286 9924 2336 9935
rect 2426 9924 2476 9934
rect 2841 9933 2891 9944
rect 2913 9933 2963 9944
rect 4597 9933 4647 9944
rect 4669 9933 4719 9944
rect 1193 9895 1221 9912
rect 1320 9894 1325 9899
rect 1433 9895 1461 9912
rect 1654 9911 1673 9916
rect 2522 9912 2539 9914
rect 1590 9901 1641 9911
rect 1909 9909 1926 9910
rect 1749 9902 1777 9907
rect 2963 9902 2995 9903
rect 4565 9902 4597 9903
rect 1781 9891 1831 9902
rect 2336 9893 2366 9897
rect 1242 9875 1270 9891
rect 1384 9875 1412 9891
rect 1909 9890 1926 9891
rect 1519 9876 1569 9885
rect 2106 9882 2156 9893
rect 2286 9882 2336 9893
rect 2396 9892 2401 9897
rect 2522 9893 2539 9895
rect 2426 9882 2476 9892
rect 2841 9891 2891 9902
rect 2913 9891 2963 9902
rect 4597 9891 4647 9902
rect 4669 9891 4719 9902
rect 1852 9871 1902 9882
rect 2522 9878 2539 9880
rect 2106 9862 2156 9873
rect 2372 9862 2377 9873
rect 2426 9862 2476 9873
rect 2913 9871 2963 9883
rect 4597 9871 4647 9883
rect 2396 9856 2401 9862
rect 2522 9859 2539 9861
rect 1242 9833 1270 9849
rect 1384 9833 1412 9849
rect 1488 9843 1519 9849
rect 1519 9834 1569 9843
rect 1818 9840 1852 9846
rect 2882 9841 2886 9871
rect 2963 9870 2992 9871
rect 4568 9870 4597 9871
rect 4674 9841 4678 9871
rect 1852 9829 1902 9840
rect 2078 9831 2106 9837
rect 2156 9831 2184 9837
rect 2396 9831 2426 9837
rect 2106 9820 2156 9831
rect 2426 9820 2476 9831
rect 2913 9829 2963 9841
rect 4597 9829 4647 9841
rect 3088 9825 3105 9827
rect 3482 9826 3499 9828
rect 4061 9826 4078 9828
rect 4455 9825 4472 9827
rect 3088 9806 3105 9808
rect 3482 9807 3499 9809
rect 4061 9807 4078 9809
rect 4455 9806 4472 9808
rect 1193 9782 1221 9799
rect 1433 9782 1461 9799
rect 1590 9788 1641 9798
rect 2913 9789 2963 9801
rect 4597 9789 4647 9801
rect 1559 9782 1590 9788
rect 1668 9761 1673 9788
rect 1781 9778 1831 9789
rect 1749 9773 1781 9778
rect 2106 9771 2156 9782
rect 2426 9771 2476 9782
rect 2078 9765 2106 9771
rect 2156 9765 2184 9771
rect 2396 9765 2426 9771
rect 1193 9740 1221 9757
rect 1320 9739 1325 9744
rect 1433 9740 1461 9757
rect 1654 9756 1673 9761
rect 1590 9746 1641 9756
rect 1909 9754 1926 9755
rect 1749 9747 1777 9752
rect 1781 9736 1831 9747
rect 2396 9740 2401 9765
rect 2882 9759 2886 9789
rect 2963 9759 2992 9760
rect 4568 9759 4597 9760
rect 4674 9759 4678 9789
rect 2913 9747 2963 9759
rect 4597 9747 4647 9759
rect 2522 9741 2539 9743
rect 1242 9720 1270 9736
rect 1384 9720 1412 9736
rect 1909 9735 1926 9736
rect 1519 9721 1569 9730
rect 2106 9729 2156 9740
rect 2372 9733 2377 9734
rect 2360 9729 2377 9733
rect 2426 9729 2476 9740
rect 2841 9728 2891 9739
rect 2913 9728 2963 9739
rect 4597 9728 4647 9739
rect 4669 9728 4719 9739
rect 2963 9727 2995 9728
rect 4565 9727 4597 9728
rect 1852 9716 1902 9727
rect 2522 9722 2539 9724
rect 2106 9709 2156 9720
rect 2286 9709 2336 9720
rect 2426 9710 2476 9720
rect 2522 9707 2539 9709
rect 1242 9678 1270 9694
rect 1384 9678 1412 9694
rect 1488 9688 1519 9694
rect 1519 9679 1569 9688
rect 1818 9685 1852 9691
rect 2522 9688 2539 9690
rect 2841 9686 2891 9697
rect 2913 9686 2963 9697
rect 4597 9686 4647 9697
rect 4669 9686 4719 9697
rect 1852 9674 1902 9685
rect 3481 9680 3498 9682
rect 4062 9680 4079 9682
rect 2106 9667 2156 9678
rect 2286 9667 2336 9678
rect 2426 9668 2476 9678
rect 3088 9666 3105 9668
rect 4455 9666 4472 9668
rect 3481 9661 3498 9663
rect 4062 9661 4079 9663
rect 3088 9647 3105 9649
rect 4455 9647 4472 9649
rect 1193 9627 1221 9644
rect 1433 9627 1461 9644
rect 1590 9633 1641 9643
rect 1559 9627 1590 9633
rect 1668 9606 1673 9633
rect 1781 9623 1831 9634
rect 2106 9631 2156 9642
rect 2286 9631 2336 9642
rect 2426 9631 2476 9641
rect 2841 9632 2891 9643
rect 2913 9632 2963 9643
rect 4597 9632 4647 9643
rect 4669 9632 4719 9643
rect 1749 9618 1781 9623
rect 2522 9619 2539 9621
rect 1193 9585 1221 9602
rect 1320 9584 1325 9589
rect 1433 9585 1461 9602
rect 1654 9601 1673 9606
rect 1590 9591 1641 9601
rect 2336 9600 2366 9604
rect 1909 9599 1926 9600
rect 1749 9592 1777 9597
rect 1781 9581 1831 9592
rect 2106 9589 2156 9600
rect 2286 9589 2336 9600
rect 2396 9599 2401 9604
rect 2522 9600 2539 9602
rect 2963 9601 2995 9602
rect 4565 9601 4597 9602
rect 2426 9589 2476 9599
rect 2841 9590 2891 9601
rect 2913 9590 2963 9601
rect 4597 9590 4647 9601
rect 4669 9590 4719 9601
rect 2522 9585 2539 9587
rect 1242 9565 1270 9581
rect 1384 9565 1412 9581
rect 1909 9580 1926 9581
rect 1519 9566 1569 9575
rect 1852 9561 1902 9572
rect 2106 9569 2156 9580
rect 2372 9569 2377 9580
rect 2426 9569 2476 9580
rect 2913 9570 2963 9582
rect 4597 9570 4647 9582
rect 2396 9563 2401 9569
rect 2522 9566 2539 9568
rect 1242 9523 1270 9539
rect 1384 9523 1412 9539
rect 1488 9533 1519 9539
rect 2078 9538 2106 9544
rect 2156 9538 2184 9544
rect 2396 9538 2426 9544
rect 2882 9540 2886 9570
rect 2963 9569 2992 9570
rect 4568 9569 4597 9570
rect 4674 9540 4678 9570
rect 1519 9524 1569 9533
rect 1818 9530 1852 9536
rect 1852 9519 1902 9530
rect 2106 9527 2156 9538
rect 2426 9527 2476 9538
rect 2913 9528 2963 9540
rect 4597 9528 4647 9540
rect 2913 9489 2963 9501
rect 4597 9489 4647 9501
rect 1193 9472 1221 9489
rect 1433 9472 1461 9489
rect 1590 9478 1641 9488
rect 1559 9472 1590 9478
rect 1668 9451 1673 9478
rect 1781 9468 1831 9479
rect 2106 9478 2156 9489
rect 2426 9478 2476 9489
rect 2078 9472 2106 9478
rect 2156 9472 2184 9478
rect 2396 9472 2426 9478
rect 1749 9463 1781 9468
rect 1193 9430 1221 9447
rect 1320 9429 1325 9434
rect 1433 9430 1461 9447
rect 1654 9446 1673 9451
rect 2396 9447 2401 9472
rect 2882 9459 2886 9489
rect 2963 9459 2992 9460
rect 4568 9459 4597 9460
rect 4674 9459 4678 9489
rect 2522 9448 2539 9450
rect 2913 9447 2963 9459
rect 4597 9447 4647 9459
rect 1590 9436 1641 9446
rect 1909 9444 1926 9445
rect 1749 9437 1777 9442
rect 1781 9426 1831 9437
rect 2106 9436 2156 9447
rect 2372 9440 2377 9441
rect 2360 9436 2377 9440
rect 2426 9436 2476 9447
rect 2522 9429 2539 9431
rect 2841 9428 2891 9439
rect 2913 9428 2963 9439
rect 4597 9428 4647 9439
rect 4669 9428 4719 9439
rect 2963 9427 2995 9428
rect 4565 9427 4597 9428
rect 1242 9410 1270 9426
rect 1384 9410 1412 9426
rect 1909 9425 1926 9426
rect 1519 9411 1569 9420
rect 1852 9406 1902 9417
rect 2106 9416 2156 9427
rect 2286 9416 2336 9427
rect 2426 9417 2476 9427
rect 2522 9414 2539 9416
rect 2522 9395 2539 9397
rect 2841 9386 2891 9397
rect 2913 9386 2963 9397
rect 4597 9386 4647 9397
rect 4669 9386 4719 9397
rect 1242 9368 1270 9384
rect 1384 9368 1412 9384
rect 1488 9378 1519 9384
rect 1519 9369 1569 9378
rect 1818 9375 1852 9381
rect 1852 9364 1902 9375
rect 2106 9374 2156 9385
rect 2286 9374 2336 9385
rect 2426 9375 2476 9385
rect 1193 8960 1221 8977
rect 1433 8960 1461 8977
rect 1590 8966 1641 8976
rect 1559 8960 1590 8966
rect 1668 8939 1673 8966
rect 1781 8956 1831 8967
rect 1749 8951 1781 8956
rect 2106 8948 2156 8959
rect 2286 8948 2336 8959
rect 2426 8948 2476 8958
rect 2841 8955 2891 8966
rect 2913 8955 2963 8966
rect 1193 8918 1221 8935
rect 1320 8917 1325 8922
rect 1433 8918 1461 8935
rect 1654 8934 1673 8939
rect 2522 8936 2539 8938
rect 1590 8924 1641 8934
rect 1909 8932 1926 8933
rect 1749 8925 1777 8930
rect 1781 8914 1831 8925
rect 2963 8924 2995 8925
rect 2336 8917 2366 8921
rect 1242 8898 1270 8914
rect 1384 8898 1412 8914
rect 1909 8913 1926 8914
rect 1519 8899 1569 8908
rect 2106 8906 2156 8917
rect 2286 8906 2336 8917
rect 2396 8916 2401 8921
rect 2522 8917 2539 8919
rect 2426 8906 2476 8916
rect 2841 8913 2891 8924
rect 2913 8913 2963 8924
rect 1852 8894 1902 8905
rect 2522 8902 2539 8904
rect 2106 8886 2156 8897
rect 2372 8886 2377 8897
rect 2426 8886 2476 8897
rect 2913 8893 2963 8905
rect 2396 8880 2401 8886
rect 2522 8883 2539 8885
rect 1242 8856 1270 8872
rect 1384 8856 1412 8872
rect 1488 8866 1519 8872
rect 1519 8857 1569 8866
rect 1818 8863 1852 8869
rect 2882 8863 2886 8893
rect 2963 8892 2992 8893
rect 1852 8852 1902 8863
rect 2078 8855 2106 8861
rect 2156 8855 2184 8861
rect 2396 8855 2426 8861
rect 2106 8844 2156 8855
rect 2426 8844 2476 8855
rect 2913 8851 2963 8863
rect 3503 8848 3520 8850
rect 3101 8845 3118 8847
rect 3503 8829 3520 8831
rect 3101 8826 3118 8828
rect 1193 8805 1221 8822
rect 1433 8805 1461 8822
rect 1590 8811 1641 8821
rect 1559 8805 1590 8811
rect 1668 8784 1673 8811
rect 1781 8801 1831 8812
rect 2913 8811 2963 8823
rect 1749 8796 1781 8801
rect 2106 8795 2156 8806
rect 2426 8795 2476 8806
rect 2078 8789 2106 8795
rect 2156 8789 2184 8795
rect 2396 8789 2426 8795
rect 1193 8763 1221 8780
rect 1320 8762 1325 8767
rect 1433 8763 1461 8780
rect 1654 8779 1673 8784
rect 1590 8769 1641 8779
rect 1909 8777 1926 8778
rect 1749 8770 1777 8775
rect 1781 8759 1831 8770
rect 2396 8764 2401 8789
rect 2882 8781 2886 8811
rect 2963 8781 2992 8782
rect 2913 8769 2963 8781
rect 2522 8765 2539 8767
rect 1242 8743 1270 8759
rect 1384 8743 1412 8759
rect 1909 8758 1926 8759
rect 2106 8753 2156 8764
rect 2372 8757 2377 8758
rect 2360 8753 2377 8757
rect 2426 8753 2476 8764
rect 1519 8744 1569 8753
rect 2841 8750 2891 8761
rect 2913 8750 2963 8761
rect 1852 8739 1902 8750
rect 2963 8749 2995 8750
rect 2522 8746 2539 8748
rect 2106 8733 2156 8744
rect 2286 8733 2336 8744
rect 2426 8734 2476 8744
rect 2522 8731 2539 8733
rect 3100 8727 3117 8729
rect 3502 8721 3519 8723
rect 1242 8701 1270 8717
rect 1384 8701 1412 8717
rect 1488 8711 1519 8717
rect 1519 8702 1569 8711
rect 1818 8708 1852 8714
rect 2522 8712 2539 8714
rect 2841 8708 2891 8719
rect 2913 8708 2963 8719
rect 3100 8708 3117 8710
rect 1852 8697 1902 8708
rect 3502 8702 3519 8704
rect 2106 8691 2156 8702
rect 2286 8691 2336 8702
rect 2426 8692 2476 8702
rect 3100 8693 3117 8695
rect 3502 8687 3519 8689
rect 3100 8674 3117 8676
rect 3502 8668 3519 8670
rect 1193 8650 1221 8667
rect 1433 8650 1461 8667
rect 1590 8656 1641 8666
rect 1559 8650 1590 8656
rect 1668 8629 1673 8656
rect 1781 8646 1831 8657
rect 2106 8655 2156 8666
rect 2286 8655 2336 8666
rect 2426 8655 2476 8665
rect 2841 8654 2891 8665
rect 2913 8654 2963 8665
rect 3100 8659 3117 8661
rect 3502 8653 3519 8655
rect 1749 8641 1781 8646
rect 2522 8643 2539 8645
rect 3100 8640 3117 8642
rect 3502 8634 3519 8636
rect 1193 8608 1221 8625
rect 1320 8607 1325 8612
rect 1433 8608 1461 8625
rect 1654 8624 1673 8629
rect 2336 8624 2366 8628
rect 1590 8614 1641 8624
rect 1909 8622 1926 8623
rect 1749 8615 1777 8620
rect 1781 8604 1831 8615
rect 2106 8613 2156 8624
rect 2286 8613 2336 8624
rect 2396 8623 2401 8628
rect 2522 8624 2539 8626
rect 2963 8623 2995 8624
rect 2426 8613 2476 8623
rect 2841 8612 2891 8623
rect 2913 8612 2963 8623
rect 3502 8619 3519 8621
rect 2522 8609 2539 8611
rect 1242 8588 1270 8604
rect 1384 8588 1412 8604
rect 1909 8603 1926 8604
rect 1519 8589 1569 8598
rect 1852 8584 1902 8595
rect 2106 8593 2156 8604
rect 2372 8593 2377 8604
rect 2426 8593 2476 8604
rect 2396 8587 2401 8593
rect 2913 8592 2963 8604
rect 2522 8590 2539 8592
rect 2078 8562 2106 8568
rect 2156 8562 2184 8568
rect 2396 8562 2426 8568
rect 2882 8562 2886 8592
rect 2963 8591 2992 8592
rect 1242 8546 1270 8562
rect 1384 8546 1412 8562
rect 1488 8556 1519 8562
rect 1519 8547 1569 8556
rect 1818 8553 1852 8559
rect 1852 8542 1902 8553
rect 2106 8551 2156 8562
rect 2426 8551 2476 8562
rect 2913 8550 2963 8562
rect 1193 8495 1221 8512
rect 1433 8495 1461 8512
rect 1590 8501 1641 8511
rect 2106 8502 2156 8513
rect 2426 8502 2476 8513
rect 2913 8511 2963 8523
rect 1559 8495 1590 8501
rect 1668 8474 1673 8501
rect 1781 8491 1831 8502
rect 2078 8496 2106 8502
rect 2156 8496 2184 8502
rect 2396 8496 2426 8502
rect 1749 8486 1781 8491
rect 1193 8453 1221 8470
rect 1320 8452 1325 8457
rect 1433 8453 1461 8470
rect 1654 8469 1673 8474
rect 2396 8471 2401 8496
rect 2882 8481 2886 8511
rect 2963 8481 2992 8482
rect 2522 8472 2539 8474
rect 1590 8459 1641 8469
rect 1909 8467 1926 8468
rect 1749 8460 1777 8465
rect 2106 8460 2156 8471
rect 2372 8464 2377 8465
rect 2360 8460 2377 8464
rect 2426 8460 2476 8471
rect 2913 8469 2963 8481
rect 1781 8449 1831 8460
rect 2522 8453 2539 8455
rect 1242 8433 1270 8449
rect 1384 8433 1412 8449
rect 1909 8448 1926 8449
rect 1519 8434 1569 8443
rect 2106 8440 2156 8451
rect 2286 8440 2336 8451
rect 2426 8441 2476 8451
rect 2841 8450 2891 8461
rect 2913 8450 2963 8461
rect 2963 8449 2995 8450
rect 1852 8429 1902 8440
rect 2522 8438 2539 8440
rect 2522 8419 2539 8421
rect 1242 8391 1270 8407
rect 1384 8391 1412 8407
rect 1488 8401 1519 8407
rect 1519 8392 1569 8401
rect 1818 8398 1852 8404
rect 2106 8398 2156 8409
rect 2286 8398 2336 8409
rect 2426 8399 2476 8409
rect 2841 8408 2891 8419
rect 2913 8408 2963 8419
rect 1852 8387 1902 8398
rect 7469 7523 7472 7562
rect 7511 7523 7514 7562
rect 7565 7523 7568 7562
rect 7607 7523 7610 7562
rect 7661 7523 7664 7562
rect 7703 7523 7706 7562
rect 7757 7523 7760 7562
rect 7799 7523 7802 7562
rect 7853 7523 7856 7562
rect 7895 7523 7898 7562
rect 7949 7523 7952 7562
rect 7991 7523 7994 7562
rect 7469 7362 7472 7401
rect 7511 7362 7514 7401
rect 7565 7361 7568 7400
rect 7607 7361 7610 7400
rect 7661 7361 7664 7400
rect 7703 7361 7706 7400
rect 7757 7361 7760 7400
rect 7799 7361 7802 7400
rect 7853 7361 7856 7400
rect 7895 7361 7898 7400
rect 7949 7362 7952 7401
rect 7991 7362 7994 7401
rect 7469 7201 7472 7240
rect 7511 7201 7514 7240
rect 7565 7200 7568 7239
rect 7607 7200 7610 7239
rect 7661 7200 7664 7239
rect 7703 7200 7706 7239
rect 7757 7200 7760 7239
rect 7799 7200 7802 7239
rect 7853 7200 7856 7239
rect 7895 7200 7898 7239
rect 7949 7201 7952 7240
rect 7991 7201 7994 7240
rect 8041 7134 8045 7166
rect 8055 7120 8059 7180
rect 7469 7040 7472 7079
rect 7511 7040 7514 7079
rect 7565 7039 7568 7078
rect 7607 7039 7610 7078
rect 7661 7039 7664 7078
rect 7703 7039 7706 7078
rect 7757 7039 7760 7078
rect 7799 7039 7802 7078
rect 7853 7039 7856 7078
rect 7895 7039 7898 7078
rect 7949 7040 7952 7079
rect 7991 7040 7994 7079
rect 7571 7012 7607 7017
rect 8041 6973 8045 7005
rect 8055 6959 8059 7019
rect 7469 6879 7472 6918
rect 7511 6879 7514 6918
rect 7565 6878 7568 6917
rect 7607 6878 7610 6917
rect 7661 6878 7664 6917
rect 7703 6878 7706 6917
rect 7757 6878 7760 6917
rect 7799 6878 7802 6917
rect 7853 6878 7856 6917
rect 7895 6878 7898 6917
rect 7949 6879 7952 6918
rect 7991 6879 7994 6918
rect 7737 6828 7741 6829
rect 8040 6812 8044 6844
rect 8054 6798 8058 6858
rect 7469 6718 7472 6757
rect 7511 6718 7514 6757
rect 7565 6717 7568 6756
rect 7607 6717 7610 6756
rect 7661 6717 7664 6756
rect 7703 6717 7706 6756
rect 7757 6717 7760 6756
rect 7799 6717 7802 6756
rect 7853 6717 7856 6756
rect 7895 6717 7898 6756
rect 7949 6718 7952 6757
rect 7991 6718 7994 6757
rect 8040 6650 8045 6682
rect 8054 6636 8059 6696
rect 7469 6557 7472 6596
rect 7511 6557 7514 6596
rect 7565 6556 7568 6595
rect 7607 6556 7610 6595
rect 7661 6556 7664 6595
rect 7703 6556 7706 6595
rect 7757 6556 7760 6595
rect 7799 6556 7802 6595
rect 7853 6556 7856 6595
rect 7895 6556 7898 6595
rect 7949 6557 7952 6596
rect 7991 6557 7994 6596
rect 8040 6489 8044 6521
rect 8054 6475 8058 6535
rect 7469 6396 7472 6435
rect 7511 6396 7514 6435
rect 7565 6395 7568 6434
rect 7607 6395 7610 6434
rect 7661 6395 7664 6434
rect 7703 6395 7706 6434
rect 7757 6395 7760 6434
rect 7799 6395 7802 6434
rect 7853 6395 7856 6434
rect 7895 6395 7898 6434
rect 7949 6396 7952 6435
rect 7991 6396 7994 6435
rect 7469 6235 7472 6274
rect 7511 6235 7514 6274
rect 7565 6234 7568 6273
rect 7607 6234 7610 6273
rect 7661 6234 7664 6273
rect 7703 6234 7706 6273
rect 7757 6234 7760 6273
rect 7799 6234 7802 6273
rect 7853 6234 7856 6273
rect 7895 6234 7898 6273
rect 7949 6235 7952 6274
rect 7991 6235 7994 6274
rect 8041 6169 8044 6201
rect 8055 6155 8058 6215
rect 7469 6074 7472 6113
rect 7511 6074 7514 6113
rect 7565 6074 7568 6113
rect 7607 6074 7610 6113
rect 7661 6074 7664 6113
rect 7703 6074 7706 6113
rect 7757 6074 7760 6113
rect 7799 6074 7802 6113
rect 7853 6074 7856 6113
rect 7895 6074 7898 6113
rect 7949 6074 7952 6113
rect 7991 6074 7994 6113
<< metal1 >>
rect -13106 14454 -12717 14571
rect -10247 14453 -9858 14570
rect -7388 14453 -6999 14570
rect -3198 14456 -2809 14573
rect 1014 14454 1403 14571
rect 3873 14454 4262 14571
rect 6733 14454 7122 14571
rect 9592 14454 9981 14571
rect 12451 14454 12840 14571
rect 15310 14453 15699 14570
rect 18169 14453 18558 14570
rect -12554 12222 -12231 13533
rect -9695 12563 -9372 13533
rect -6836 12992 -6513 13533
rect -5582 13312 -5565 13324
rect -6879 12961 -6496 12992
rect -6879 12736 -6836 12961
rect -6513 12736 -6496 12961
rect -6879 12718 -6496 12736
rect -5617 12656 -5565 13312
rect -5623 12645 -5558 12656
rect -5623 12608 -5617 12645
rect -5565 12608 -5558 12645
rect -5623 12605 -5558 12608
rect -9711 12512 -9361 12563
rect -9711 12287 -9695 12512
rect -9372 12287 -9361 12512
rect -9711 12274 -9361 12287
rect -12771 12183 -12231 12222
rect -12771 11860 -12737 12183
rect -12512 11860 -12231 12183
rect -14015 11852 -13676 11859
rect -14112 11843 -13676 11852
rect -14435 11520 -13890 11843
rect -13704 11520 -13676 11843
rect -12771 11842 -12477 11860
rect -5617 11837 -5565 12605
rect -5277 12214 -5236 13335
rect -2566 13135 -2450 13326
rect -2566 13022 170 13135
rect -2566 13002 189 13022
rect 37 12862 170 13002
rect 1566 12911 1889 13534
rect 2730 13326 2791 13340
rect 2728 13130 2846 13326
rect 2648 13039 2846 13130
rect 2648 13021 2829 13039
rect 3172 13023 3244 13409
rect 2648 12952 2721 13021
rect 4425 12911 4748 13533
rect 7284 12911 7607 13533
rect 8177 13272 8196 13273
rect 8890 13272 8962 13409
rect 8177 13237 8962 13272
rect 8177 13024 8196 13237
rect 10143 13218 10466 13533
rect 10067 13190 10466 13218
rect 10065 13170 10466 13190
rect 10047 13073 10482 13170
rect 10047 12867 10143 13073
rect 10466 12867 10482 13073
rect 10047 12800 10482 12867
rect 13002 12752 13325 13533
rect 12972 12708 13327 12752
rect 12972 12378 13002 12708
rect 13208 12378 13327 12708
rect 12972 12347 13327 12378
rect -5289 12211 -5236 12214
rect -5289 12170 -5283 12211
rect -5242 12170 -5236 12211
rect 15861 12189 16184 13533
rect -5289 12167 -5236 12170
rect -5637 11828 -5565 11837
rect -5637 11776 -5631 11828
rect -5579 11776 -5565 11828
rect -5637 11764 -5565 11776
rect -14112 11452 -13676 11520
rect -15468 10968 -15343 11357
rect -13098 8984 -12872 8988
rect -14435 8661 -13085 8984
rect -12877 8661 -12872 8984
rect -13098 8657 -12872 8661
rect -15467 8110 -15342 8499
rect -5617 8229 -5565 11764
rect -5277 11742 -5236 12167
rect 15841 12159 16200 12189
rect 15841 11953 15861 12159
rect 16184 11953 16200 12159
rect 15841 11936 16200 11953
rect 18720 11840 19043 13533
rect -5291 11732 -5229 11742
rect -5291 11691 -5278 11732
rect -5237 11691 -5229 11732
rect -5291 11683 -5229 11691
rect 18689 11717 19065 11840
rect -5625 8226 -5562 8229
rect -5625 8174 -5621 8226
rect -5569 8174 -5562 8226
rect -5625 8169 -5562 8174
rect -5277 8127 -5236 11683
rect 18689 11512 18720 11717
rect 19043 11512 19065 11717
rect 18689 11478 19065 11512
rect 20124 11771 20465 11803
rect 20124 11448 20154 11771
rect 20353 11448 20788 11771
rect 10956 11382 11398 11443
rect 20124 11399 20465 11448
rect 10956 11350 10980 11382
rect 11202 11350 11398 11382
rect 10956 8432 11398 11350
rect 21692 10898 21817 11287
rect 19283 8912 19515 8920
rect 19283 8589 19299 8912
rect 19508 8589 20787 8912
rect 19283 8583 19515 8589
rect 10953 8420 11400 8432
rect 10953 8311 10964 8420
rect 11392 8311 11400 8420
rect 10953 8300 11400 8311
rect -5282 8124 -5234 8127
rect -5282 8080 -5278 8124
rect -5237 8080 -5234 8124
rect -5282 8077 -5234 8080
rect -12707 6125 -12484 6133
rect -14434 5802 -12695 6125
rect -12487 5802 -12484 6125
rect -12707 5787 -12484 5802
rect -15468 5250 -15343 5639
rect -12256 3266 -12015 3276
rect -14435 2943 -12232 3266
rect -12024 2943 -12015 3266
rect -12256 2933 -12015 2943
rect -15466 2391 -15341 2780
rect -11800 407 -11573 414
rect -14434 84 -11791 407
rect -11583 84 -11573 407
rect -11800 74 -11573 84
rect -15467 -467 -15342 -78
rect -11364 -2452 -11139 -2446
rect -14435 -2775 -11357 -2452
rect -11149 -2775 -11139 -2452
rect -11364 -2783 -11139 -2775
rect -15468 -3327 -15343 -2938
rect -10932 -5311 -10707 -5300
rect -14435 -5634 -10692 -5311
rect -10932 -5645 -10707 -5634
rect -15467 -6185 -15342 -5796
rect 10956 -7830 11398 8300
rect 21691 8038 21816 8427
rect 18866 6053 19102 6066
rect 18866 5730 18874 6053
rect 19083 5730 20789 6053
rect 18866 5720 19102 5730
rect 21691 5178 21816 5567
rect 18465 3194 18693 3210
rect 18465 2871 18476 3194
rect 18685 2871 20787 3194
rect 18465 2860 18693 2871
rect 21692 2322 21817 2711
rect 18035 335 18277 347
rect 18035 12 18051 335
rect 18260 12 20787 335
rect 18035 -4 18277 12
rect 21690 -539 21815 -150
rect 17646 -2524 17873 -2513
rect 17646 -2847 17657 -2524
rect 17866 -2847 20788 -2524
rect 17646 -2860 17873 -2847
rect 21692 -3397 21817 -3008
rect 17206 -5383 17436 -5375
rect 17206 -5706 20788 -5383
rect 17206 -5716 17436 -5706
rect 21692 -6258 21817 -5869
rect 10864 -7841 11398 -7830
rect -10526 -8170 -10285 -8160
rect -14435 -8493 -10503 -8170
rect -10295 -8493 -10285 -8170
rect 10864 -8283 10882 -7841
rect 11324 -8204 11398 -7841
rect 11324 -8283 11340 -8204
rect 10864 -8300 11340 -8283
rect -10526 -8511 -10285 -8493
rect -15464 -9043 -15339 -8654
rect -10098 -11029 -9852 -11022
rect -14435 -11352 -9852 -11029
rect -10098 -11357 -9852 -11352
rect -15466 -11904 -15341 -11515
rect -9661 -13888 -9421 -13874
rect -14436 -14211 -9641 -13888
rect -9433 -14211 -9421 -13888
rect -9661 -14221 -9421 -14211
rect -15467 -14763 -15342 -14374
rect -9267 -16747 -9018 -16739
rect -14436 -17070 -9244 -16747
rect -9036 -17070 -9018 -16747
rect -9267 -17089 -9018 -17070
rect -15467 -17622 -15342 -17233
rect -8820 -19606 -8585 -19596
rect -14434 -19929 -8800 -19606
rect -8592 -19929 -8585 -19606
rect -8820 -19942 -8585 -19929
rect -15466 -20481 -15341 -20092
rect -8420 -22465 -8149 -22459
rect -14434 -22788 -8370 -22465
rect -8162 -22788 -8149 -22465
rect -8420 -22800 -8149 -22788
rect -15466 -23339 -15341 -22950
<< via1 >>
rect -6836 12736 -6513 12961
rect -5617 12608 -5565 12645
rect -9695 12287 -9372 12512
rect -12737 11860 -12512 12183
rect -13890 11520 -13704 11843
rect 10143 12867 10466 13073
rect 13002 12378 13208 12708
rect -5283 12170 -5242 12211
rect -5631 11776 -5579 11828
rect -13085 8661 -12877 8984
rect 15861 11953 16184 12159
rect -5278 11691 -5237 11732
rect -5621 8174 -5569 8226
rect 18720 11512 19043 11717
rect 20154 11448 20353 11771
rect 10980 11350 11202 11382
rect 19299 8589 19508 8912
rect 10964 8311 11392 8420
rect -5278 8080 -5237 8124
rect -12695 5802 -12487 6125
rect -12232 2943 -12024 3266
rect -11791 84 -11583 407
rect -11357 -2775 -11149 -2452
rect 18874 5730 19083 6053
rect 18476 2871 18685 3194
rect 18051 12 18260 335
rect 17657 -2847 17866 -2524
rect -10503 -8493 -10295 -8170
rect 10882 -8283 11324 -7841
rect -9641 -14211 -9433 -13888
rect -9244 -17070 -9036 -16747
rect -8800 -19929 -8592 -19606
rect -8370 -22788 -8162 -22465
<< metal2 >>
rect 21381 14165 21500 14166
rect -15126 14164 -13833 14165
rect -15139 14025 -13833 14164
rect 20201 14113 21500 14165
rect 20180 14037 21500 14113
rect -15139 13873 -14910 14025
rect -15094 13869 -14910 13873
rect -15050 13017 -14910 13869
rect 21284 13905 21500 14037
rect -14423 13388 -13848 13528
rect 20116 13395 20783 13535
rect -14423 12916 -14283 13388
rect 10028 13073 10508 13153
rect -6892 12987 -6483 13012
rect -6892 12961 -2695 12987
rect -6892 12736 -6836 12961
rect -6513 12762 -2695 12961
rect 10028 12944 10143 13073
rect 8858 12867 10143 12944
rect 10466 12944 10508 13073
rect 10466 12867 10513 12944
rect -6513 12736 -6483 12762
rect 8858 12738 10513 12867
rect 20642 12844 20782 13395
rect 21284 12982 21412 13905
rect 21336 12908 21412 12982
rect -6892 12702 -6483 12736
rect 12987 12708 13318 12737
rect -5622 12651 -5560 12653
rect -5622 12645 -2707 12651
rect -5622 12608 -5617 12645
rect -5565 12614 -2707 12645
rect -5565 12608 -5560 12614
rect -5622 12607 -5560 12608
rect -9704 12538 -9366 12549
rect -9745 12512 -2695 12538
rect 12987 12531 13002 12708
rect -9745 12313 -9695 12512
rect -9704 12287 -9695 12313
rect -9372 12313 -2695 12512
rect 8858 12378 13002 12531
rect 13208 12531 13318 12708
rect 13208 12378 13350 12531
rect 8858 12325 13350 12378
rect -9372 12287 -9366 12313
rect -9704 12281 -9366 12287
rect -5287 12211 -5239 12212
rect -12758 12183 -12494 12207
rect -12758 12089 -12737 12183
rect -12766 11864 -12737 12089
rect -12758 11860 -12737 11864
rect -12512 12089 -12494 12183
rect -5287 12170 -5283 12211
rect -5242 12209 -5239 12211
rect -5242 12171 -2708 12209
rect -5242 12170 -5239 12171
rect -5287 12169 -5239 12170
rect 15826 12159 16219 12168
rect 15826 12123 15861 12159
rect -12512 11864 -2735 12089
rect 8858 11953 15861 12123
rect 16184 11953 16219 12159
rect 8858 11917 16219 11953
rect 15826 11916 16219 11917
rect -12512 11860 -12494 11864
rect -13981 11843 -13692 11851
rect -12758 11847 -12494 11860
rect -13981 11655 -13890 11843
rect -13984 11520 -13890 11655
rect -13704 11655 -13692 11843
rect -5634 11828 -5572 11831
rect -5634 11776 -5631 11828
rect -5579 11822 -5572 11828
rect -5579 11781 -2740 11822
rect -5579 11776 -5572 11781
rect -5634 11772 -5572 11776
rect 19876 11771 20447 11846
rect -5287 11732 -5233 11735
rect -5287 11691 -5278 11732
rect -5237 11691 -2744 11732
rect 18706 11717 19056 11743
rect -5287 11687 -5233 11691
rect 18706 11689 18720 11717
rect -13704 11520 -2772 11655
rect -13984 11469 -2772 11520
rect 8858 11512 18720 11689
rect 19043 11689 19056 11717
rect 19043 11512 19065 11689
rect 8858 11484 19065 11512
rect 19876 11448 20154 11771
rect 20353 11448 20447 11771
rect 8876 11382 11209 11387
rect 8876 11350 10980 11382
rect 11202 11350 11209 11382
rect 8876 11344 11209 11350
rect 19876 11282 20447 11448
rect 19832 11278 20447 11282
rect 8858 11232 20447 11278
rect -13095 11003 -2743 11211
rect 8858 11042 20431 11232
rect -13095 8992 -12887 11003
rect 19298 10804 19507 10822
rect -12679 10515 -2695 10723
rect 8858 10595 19507 10804
rect -13102 8984 -12868 8992
rect -13102 8661 -13085 8984
rect -12877 8661 -12868 8984
rect -13102 8655 -12868 8661
rect -13095 8568 -12887 8655
rect -12679 6132 -12471 10515
rect -12701 6125 -12471 6132
rect -12701 5802 -12695 6125
rect -12487 5802 -12471 6125
rect -12701 5791 -12471 5802
rect -12679 5758 -12471 5791
rect -12245 10033 -2695 10241
rect 8858 10055 19093 10264
rect -12245 3284 -12037 10033
rect -11791 9563 -2695 9771
rect 8858 9567 18685 9776
rect -12266 3266 -12009 3284
rect -12266 2943 -12232 3266
rect -12024 2943 -12009 3266
rect -12266 2924 -12009 2943
rect -12245 2920 -12037 2924
rect -11791 422 -11583 9563
rect -11356 9137 -2695 9345
rect -11807 407 -11568 422
rect -11807 84 -11791 407
rect -11583 84 -11568 407
rect -11807 65 -11568 84
rect -11791 12 -11583 65
rect -11356 -2439 -11148 9137
rect 8858 9047 18276 9256
rect -10922 8730 -2695 8938
rect -11374 -2452 -11129 -2439
rect -11374 -2775 -11357 -2452
rect -11149 -2775 -11129 -2452
rect -11374 -2791 -11129 -2775
rect -11356 -2803 -11148 -2791
rect -10922 -5290 -10714 8730
rect 8858 8543 17863 8752
rect -10506 8315 -2695 8523
rect 10955 8421 11408 8429
rect 8886 8420 11415 8421
rect -10947 -5663 -10687 -5290
rect -10922 -5696 -10714 -5663
rect -10506 -8153 -10298 8315
rect 8886 8311 10964 8420
rect 11392 8311 11415 8420
rect 8886 8306 11415 8311
rect 10955 8304 11408 8306
rect -5624 8226 -5564 8227
rect -5624 8174 -5621 8226
rect -5569 8222 -5564 8226
rect -5569 8178 -2690 8222
rect -5569 8174 -5564 8178
rect -5624 8171 -5564 8174
rect -5281 8124 -5235 8125
rect -5281 8080 -5278 8124
rect -5237 8080 -2694 8124
rect -5281 8078 -5235 8080
rect -10081 7800 -2695 8008
rect 8890 7992 17439 8201
rect -10548 -8170 -10277 -8153
rect -10548 -8493 -10503 -8170
rect -10295 -8493 -10277 -8170
rect -10548 -8520 -10277 -8493
rect -10506 -8592 -10298 -8520
rect -10081 -11015 -9873 7800
rect -9655 7374 -2695 7582
rect -10114 -11363 -9840 -11015
rect -10081 -11444 -9873 -11363
rect -9655 -13844 -9447 7374
rect -9240 6870 -2695 7078
rect -9677 -13888 -9398 -13844
rect -9677 -14211 -9641 -13888
rect -9433 -14211 -9398 -13888
rect -9677 -14249 -9398 -14211
rect -9655 -14277 -9447 -14249
rect -9240 -16722 -9032 6870
rect -8805 6309 -2695 6517
rect -9289 -16747 -9006 -16722
rect -9289 -17070 -9244 -16747
rect -9036 -17070 -9006 -16747
rect -9289 -17100 -9006 -17070
rect -9240 -17156 -9032 -17100
rect -8805 -19580 -8597 6309
rect -8389 5839 -2695 6047
rect -8840 -19606 -8575 -19580
rect -8840 -19929 -8800 -19606
rect -8592 -19929 -8575 -19606
rect -8840 -19952 -8575 -19929
rect -8805 -19953 -8597 -19952
rect -8389 -22450 -8181 5839
rect -8408 -22465 -8141 -22450
rect -8408 -22788 -8370 -22465
rect -8162 -22788 -8141 -22465
rect -8408 -22803 -8141 -22788
rect -2235 -23386 -1901 5853
rect -1269 -23816 -1067 5843
rect -863 -23659 -661 5843
rect -863 -23815 -660 -23659
rect -466 -23660 -264 5843
rect -66 -23660 136 5843
rect -863 -23816 -661 -23815
rect -467 -23816 -264 -23660
rect -67 -23816 136 -23660
rect 339 -23816 541 5843
rect 740 -23659 942 5843
rect 739 -23815 942 -23659
rect 740 -23816 942 -23815
rect 1140 -23816 1342 5843
rect 1549 -23816 1751 5843
rect 1962 -23660 2164 5843
rect 2362 -23660 2564 5843
rect 2758 -23660 2960 5843
rect 1961 -23816 2164 -23660
rect 2361 -23816 2564 -23660
rect 2757 -23816 2960 -23660
rect 3163 -23659 3365 5843
rect 3163 -23815 3366 -23659
rect 3163 -23816 3365 -23815
rect 3572 -23816 3774 5843
rect 3973 -23661 4175 5843
rect 4377 -23660 4579 5843
rect 3973 -23816 4176 -23661
rect 4377 -23816 4580 -23660
rect 4786 -23662 4988 5843
rect 4786 -23816 4989 -23662
rect 5191 -23816 5393 5843
rect 5588 -23816 5790 5843
rect 6000 -23816 6202 5843
rect 3974 -23817 4176 -23816
rect 4787 -23818 4989 -23816
rect 6413 -23817 6615 5843
rect 6814 -23816 7016 5843
rect 7215 -23648 7417 5843
rect 7215 -23814 7419 -23648
rect 7624 -23650 7826 5843
rect 7624 -23816 7827 -23650
rect 8041 -23816 8243 5843
rect 8441 -23650 8643 5843
rect 8842 -23650 9044 5843
rect 9238 -23650 9440 5843
rect 8441 -23816 8644 -23650
rect 8839 -23816 9044 -23650
rect 9237 -23816 9440 -23650
rect 9643 -23650 9845 5843
rect 10049 -23650 10251 5843
rect 17230 -5151 17439 7992
rect 17654 -2504 17863 8543
rect 18067 344 18276 9047
rect 18476 3221 18685 9567
rect 18884 6071 19093 10055
rect 19298 8927 19507 10595
rect 19278 8912 19521 8927
rect 19278 8589 19299 8912
rect 19508 8589 19521 8912
rect 19278 8573 19521 8589
rect 19298 8506 19507 8573
rect 18860 6053 19111 6071
rect 18860 5730 18874 6053
rect 19083 5730 19111 6053
rect 18860 5714 19111 5730
rect 18456 3194 18708 3221
rect 18456 2871 18476 3194
rect 18685 2871 18708 3194
rect 18456 2850 18708 2871
rect 18476 2847 18685 2850
rect 18040 335 18276 344
rect 18040 12 18051 335
rect 18260 12 18276 335
rect 18040 2 18276 12
rect 18067 -69 18276 2
rect 17637 -2524 17880 -2504
rect 17637 -2847 17657 -2524
rect 17866 -2847 17880 -2524
rect 17637 -2875 17880 -2847
rect 17231 -5341 17439 -5151
rect 17231 -5353 17440 -5341
rect 17220 -5359 17440 -5353
rect 17194 -5727 17447 -5359
rect 17220 -5729 17429 -5727
rect 21338 -6998 21412 -6964
rect 20640 -7101 20780 -7023
rect 21272 -7038 21413 -6998
rect 20639 -7113 20780 -7101
rect 21274 -7107 21412 -7038
rect 20638 -7128 20780 -7113
rect 20638 -7218 20779 -7128
rect 21273 -7224 21413 -7107
rect 10871 -7841 11331 -7836
rect 10871 -8283 10882 -7841
rect 11324 -7914 11331 -7841
rect 11324 -8082 20786 -7914
rect 11324 -8211 20799 -8082
rect 11324 -8283 11331 -8211
rect 10871 -8293 11331 -8283
rect 9643 -23816 9847 -23650
rect 10049 -23816 10253 -23650
rect -15053 -24304 -14913 -24107
rect -14423 -24337 -14283 -23971
use sky130_hilas_TopProtection  sky130_hilas_TopProtection_0
timestamp 1627737364
transform 1 0 -13875 0 1 13286
box -2 -76 34131 1170
use sky130_hilas_LeftProtection  sky130_hilas_LeftProtection_0
timestamp 1627737364
transform 1 0 -13278 0 1 -15672
box -2065 -8439 -833 28728
use sky130_hilas_RightProtection  sky130_hilas_RightProtection_0
timestamp 1627737364
transform 1 0 22518 0 1 -15744
box -2054 8715 -826 28728
use sky130_hilas_TopLevelTextStructure  sky130_hilas_TopLevelTextStructure_0
timestamp 1627744303
transform 1 0 -2990 0 1 6624
box 218 -793 13243 6785
<< labels >>
rlabel metal1 21692 -6258 21817 -5869 0 IO07
port 1 nsew
rlabel metal1 21692 -3397 21817 -3008 0 IO08
port 2 nsew
rlabel metal1 21690 -539 21815 -150 0 IO09
port 3 nsew
rlabel metal1 21692 2322 21817 2711 0 IO10
port 4 nsew
rlabel metal1 21691 5178 21816 5567 0 IO11
port 5 nsew
rlabel metal1 21691 8038 21816 8427 0 IO12
port 6 nsew
rlabel metal1 21692 10898 21817 11287 0 IO13
port 7 nsew
rlabel metal1 -15468 10968 -15343 11357 0 IO25
port 8 nsew
rlabel metal1 -15467 8110 -15342 8499 0 IO26
port 9 nsew
rlabel metal1 -15468 5250 -15343 5639 0 IO27
port 10 nsew
rlabel metal1 -15466 2391 -15341 2780 0 IO28
port 11 nsew
rlabel metal1 -15467 -467 -15342 -78 0 IO29
port 12 nsew
rlabel metal1 -15468 -3327 -15343 -2938 0 IO30
port 13 nsew
rlabel metal1 -15467 -6185 -15342 -5796 0 IO31
port 14 nsew
rlabel metal1 -15464 -9043 -15339 -8654 0 IO32
port 15 nsew
rlabel metal1 -15466 -11904 -15341 -11515 0 IO33
port 16 nsew
rlabel metal1 -15467 -14763 -15342 -14374 0 IO34
port 17 nsew
rlabel metal1 -15467 -17622 -15342 -17233 0 IO35
port 18 nsew
rlabel metal1 -15466 -20481 -15341 -20092 0 IO36
port 19 nsew
rlabel metal1 -15466 -23339 -15341 -22950 0 IO37
port 20 nsew
rlabel metal2 -15139 13873 -14971 14164 0 VSSA1
port 21 nsew
rlabel metal1 -13106 14454 -12717 14571 0 ANALOG10
port 22 nsew
rlabel metal1 -10247 14453 -9858 14570 0 ANALOG09
port 23 nsew
rlabel metal1 -7388 14453 -6999 14570 0 ANALOG08
port 24 nsew
rlabel metal1 -3198 14456 -2809 14573 0 ANALOG07
port 25 nsew
rlabel metal1 1014 14454 1403 14571 0 ANALOG06
port 26 nsew
rlabel metal1 3873 14454 4262 14571 0 ANALOG05
port 27 nsew
rlabel metal1 6733 14454 7122 14571 0 ANALOG04
port 28 nsew
rlabel metal1 9592 14454 9981 14571 0 ANALOG03
port 29 nsew
rlabel metal1 12451 14454 12840 14571 0 ANALOG02
port 30 nsew
rlabel metal1 15310 14453 15699 14570 0 ANALOG01
port 31 nsew
rlabel metal1 18169 14453 18558 14570 0 ANALOG00
port 32 nsew
rlabel metal2 21381 13908 21500 14166 0 VSSA1
port 33 nsew
rlabel metal2 -14423 -24337 -14283 -24197 0 VDDA1
port 34 nsew
rlabel metal2 -15053 -24304 -14913 -24164 0 VSSA1
port 33 nsew
rlabel metal2 20639 -7218 20779 -7101 0 VDDA1
port 34 nsew
rlabel metal2 21273 -7224 21413 -7107 0 VSSA1
port 33 nsew
rlabel metal2 -1269 -23816 -1067 -23660 0 LADATAOUT00
port 36 nsew
rlabel metal2 -862 -23815 -660 -23659 0 LADATAOUT01
port 35 nsew
rlabel metal2 -467 -23816 -265 -23660 0 LADATAOUT02
port 37 nsew
rlabel metal2 -67 -23816 135 -23660 0 LADATAOUT03
port 38 nsew
rlabel metal2 339 -23816 541 -23660 0 LADATAOUT04
port 39 nsew
rlabel metal2 739 -23815 941 -23659 0 LADATAOUT05
port 40 nsew
rlabel metal2 1140 -23816 1342 -23660 0 LADATAOUT06
port 41 nsew
rlabel metal2 1549 -23816 1751 -23660 0 LADATAOUT07
port 42 nsew
rlabel metal2 1961 -23816 2163 -23660 0 LADATAOUT08
port 43 nsew
rlabel metal2 2361 -23816 2563 -23660 0 LADATAOUT09
port 44 nsew
rlabel metal2 2757 -23816 2959 -23660 0 LADATAOUT10
port 45 nsew
rlabel metal2 3164 -23815 3366 -23659 0 LADATAOUT11
port 46 nsew
rlabel metal2 3572 -23816 3774 -23660 0 LADATAOUT12
port 47 nsew
rlabel metal2 3974 -23817 4176 -23661 0 LADATAOUT13
port 48 nsew
rlabel metal2 4378 -23816 4580 -23660 0 LADATAOUT14
port 49 nsew
rlabel metal2 4787 -23818 4989 -23662 0 LADATAOUT15
port 50 nsew
rlabel metal2 5191 -23816 5393 -23660 0 LADATA16
port 51 nsew
rlabel metal2 5588 -23816 5790 -23660 0 LADATAOUT17
port 52 nsew
rlabel metal2 6000 -23815 6202 -23659 0 LADATAOUT18
port 53 nsew
rlabel metal2 6413 -23817 6615 -23661 0 LADATAOUT19
port 54 nsew
rlabel metal2 6814 -23816 7016 -23660 0 LADATAOUT20
port 55 nsew
rlabel metal2 7215 -23814 7419 -23648 0 LADATAOUT21
port 56 nsew
rlabel metal2 7624 -23816 7827 -23650 0 LADATAOUT22
port 57 nsew
rlabel metal2 8039 -23816 8242 -23650 0 LADATAOUT23
port 58 nsew
rlabel metal2 8441 -23816 8644 -23650 0 LADATAOUT24
port 59 nsew
rlabel metal2 8839 -23816 9042 -23650 0 LADATAIN00
port 60 nsew
rlabel metal2 9237 -23816 9440 -23650 0 LADATAIN01
port 61 nsew
rlabel metal2 9644 -23816 9847 -23650 0 LADATAIN02
port 62 nsew
rlabel metal2 10050 -23816 10253 -23650 0 LADATAIN03
port 63 nsew
rlabel metal2 20683 -8211 20799 -8085 0 VCCA
port 64 nsew
<< end >>
