VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_ta2cell_1fg
  CLASS BLOCK ;
  FOREIGN sky130_hilas_ta2cell_1fg ;
  ORIGIN 26.160 -1.400 ;
  SIZE 28.090 BY 6.050 ;
  OBS
      LAYER nwell ;
        RECT 0.650 7.270 1.930 7.450 ;
        RECT 0.650 1.400 1.930 1.590 ;
      LAYER met1 ;
        RECT -4.160 7.370 -3.970 7.450 ;
        RECT -3.720 7.370 -3.440 7.450 ;
        RECT -0.030 7.310 0.310 7.450 ;
        RECT 0.630 7.300 0.910 7.450 ;
        RECT -0.030 1.400 0.310 1.590 ;
        RECT 0.640 1.400 0.910 1.610 ;
      LAYER met2 ;
        RECT -2.600 7.180 -2.290 7.420 ;
        RECT -1.490 6.550 -1.270 6.570 ;
        RECT -17.260 6.170 -16.420 6.370 ;
        RECT -1.540 6.210 -1.270 6.550 ;
        RECT -16.810 5.700 -6.670 5.920 ;
        RECT -3.280 5.710 -2.930 5.930 ;
        RECT -16.860 4.730 -7.850 4.950 ;
        RECT -16.810 2.950 -11.150 3.170 ;
        RECT -17.310 2.410 -16.420 2.650 ;
        RECT -11.370 2.620 -11.150 2.950 ;
        RECT -8.070 3.120 -7.850 4.730 ;
        RECT -6.890 4.500 -6.670 5.700 ;
        RECT -1.470 5.640 -1.270 5.650 ;
        RECT -1.470 5.310 -1.250 5.640 ;
        RECT -1.450 5.300 -1.250 5.310 ;
        RECT -2.520 4.510 -2.200 4.750 ;
        RECT -6.920 4.460 -6.670 4.500 ;
        RECT -6.920 3.820 -6.660 4.460 ;
        RECT -6.920 3.610 -2.790 3.820 ;
        RECT -3.000 3.470 -2.790 3.610 ;
        RECT -3.000 3.260 -1.130 3.470 ;
        RECT -8.070 2.900 -5.220 3.120 ;
        RECT -7.000 2.620 -1.130 2.670 ;
        RECT -11.370 2.460 -1.130 2.620 ;
        RECT -11.370 2.400 -6.610 2.460 ;
  END
END sky130_hilas_ta2cell_1fg
END LIBRARY

