magic
tech sky130A
timestamp 1628285143
<< nmos >>
rect 16 -31 42 215
<< ndiff >>
rect -12 206 16 215
rect -12 189 -7 206
rect 10 189 16 206
rect -12 172 16 189
rect -12 155 -7 172
rect 10 155 16 172
rect -12 138 16 155
rect -12 121 -7 138
rect 10 121 16 138
rect -12 104 16 121
rect -12 87 -7 104
rect 10 87 16 104
rect -12 70 16 87
rect -12 53 -7 70
rect 10 53 16 70
rect -12 36 16 53
rect -12 19 -7 36
rect 10 19 16 36
rect -12 2 16 19
rect -12 -15 -7 2
rect 10 -15 16 2
rect -12 -31 16 -15
rect 42 206 70 215
rect 42 189 48 206
rect 65 189 70 206
rect 42 172 70 189
rect 42 155 48 172
rect 65 155 70 172
rect 42 138 70 155
rect 42 121 48 138
rect 65 121 70 138
rect 42 104 70 121
rect 42 87 48 104
rect 65 87 70 104
rect 42 70 70 87
rect 42 53 48 70
rect 65 53 70 70
rect 42 36 70 53
rect 42 19 48 36
rect 65 19 70 36
rect 42 2 70 19
rect 42 -15 48 2
rect 65 -15 70 2
rect 42 -31 70 -15
<< ndiffc >>
rect -7 189 10 206
rect -7 155 10 172
rect -7 121 10 138
rect -7 87 10 104
rect -7 53 10 70
rect -7 19 10 36
rect -7 -15 10 2
rect 48 189 65 206
rect 48 155 65 172
rect 48 121 65 138
rect 48 87 65 104
rect 48 53 65 70
rect 48 19 65 36
rect 48 -15 65 2
<< poly >>
rect 16 215 42 228
rect 16 -44 42 -31
<< locali >>
rect -7 206 10 214
rect -7 172 10 189
rect -7 138 10 155
rect -7 104 10 121
rect -7 70 10 87
rect -7 36 10 53
rect -7 2 10 19
rect -7 -26 10 -15
rect 48 206 65 214
rect 48 172 65 189
rect 48 138 65 155
rect 48 104 65 121
rect 48 70 65 87
rect 48 36 65 53
rect 48 2 65 19
rect 48 -26 65 -15
<< end >>
