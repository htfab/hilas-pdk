magic
tech sky130A
timestamp 1634057841
<< checkpaint >>
rect 359 2962 2168 3031
rect -234 650 2680 2962
rect 515 309 2625 650
rect 515 -630 2324 309
<< error_s >>
rect 58 1430 64 1436
rect 111 1430 117 1436
rect 52 1380 58 1386
rect 117 1380 123 1386
rect 481 1371 487 1377
rect 586 1371 592 1377
rect 475 1321 481 1327
rect 592 1321 598 1327
rect 481 1070 487 1076
rect 586 1070 592 1076
rect 58 1016 64 1022
rect 111 1016 117 1022
rect 475 1020 481 1026
rect 592 1020 598 1026
rect 52 966 58 972
rect 117 966 123 972
<< nwell >>
rect 1665 1485 1792 1503
rect 1145 1329 1311 1351
rect 1191 1168 1219 1192
rect 1664 898 1792 917
<< locali >>
rect 283 1237 329 1246
rect 283 1220 286 1237
rect 303 1220 329 1237
rect 283 1168 329 1220
rect 283 1151 286 1168
rect 303 1151 329 1168
rect 283 1145 329 1151
<< viali >>
rect 286 1220 303 1237
rect 286 1151 303 1168
<< metal1 >>
rect 35 1496 77 1503
rect 405 1495 428 1503
rect 1057 1495 1076 1503
rect 1101 1495 1129 1503
rect 1596 1489 1630 1503
rect 1663 1488 1690 1503
rect 279 1242 317 1246
rect 279 1149 283 1242
rect 312 1149 317 1242
rect 279 1145 317 1149
rect 1596 898 1630 917
rect 1663 898 1690 919
<< via1 >>
rect 1600 1337 1626 1363
rect 283 1237 312 1242
rect 283 1220 286 1237
rect 286 1220 303 1237
rect 303 1220 312 1237
rect 283 1168 312 1220
rect 283 1151 286 1168
rect 286 1151 303 1168
rect 303 1151 312 1168
rect 283 1149 312 1151
<< metal2 >>
rect 1343 1476 1368 1502
rect 0 1435 7 1453
rect 1449 1378 1474 1415
rect 1596 1363 1630 1367
rect 1596 1358 1600 1363
rect 1145 1329 1311 1351
rect 1361 1339 1600 1358
rect 1361 1282 1380 1339
rect 1596 1337 1600 1339
rect 1626 1337 1630 1363
rect 1596 1334 1630 1337
rect 1452 1293 1473 1322
rect 282 1263 1380 1282
rect 282 1245 301 1263
rect 280 1242 315 1245
rect 280 1149 283 1242
rect 312 1149 315 1242
rect 1777 1232 1792 1254
rect 1347 1209 1372 1232
rect 1191 1168 1219 1192
rect 1777 1150 1792 1172
rect 280 1146 315 1149
rect 1296 1085 1473 1105
rect 1139 1036 1155 1076
rect 1267 1004 1473 1025
rect 0 950 8 965
rect 1187 900 1213 925
use sky130_hilas_FGBias2x1cell  sky130_hilas_FGBias2x1cell_0
timestamp 1634057765
transform 1 0 396 0 1 1280
box 0 0 1654 1052
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_0
timestamp 1634057767
transform 1 0 989 0 1 1338
box 0 0 549 1063
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1634057767
transform 1 0 1145 0 -1 1063
box 0 0 549 1063
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1634057763
transform 1 0 1637 0 1 939
box 0 0 358 746
<< labels >>
rlabel metal1 1596 898 1630 904 0 VGND
port 7 nsew ground default
rlabel metal1 1663 898 1690 904 0 VPWR
port 8 nsew power default
rlabel metal1 1596 1498 1630 1503 0 VGND
port 7 nsew ground default
rlabel metal1 1663 1498 1690 1503 0 VPWR
port 8 nsew power default
rlabel metal2 1347 1209 1372 1232 0 VIN21
port 3 nsew
rlabel metal2 1187 900 1210 925 0 VIN12
port 2 nsew analog default
rlabel metal2 1343 1476 1368 1502 0 VIN22
port 4 nsew
rlabel metal2 1777 1150 1792 1172 0 OUTPUT1
port 5 nsew
rlabel metal2 1777 1232 1792 1254 0 OUTPUT2
port 6 nsew
rlabel metal1 1057 1495 1076 1503 0 COLSEL1
port 1 nsew
rlabel metal2 0 1435 7 1453 0 DRAIN1
port 9 nsew
rlabel metal2 0 950 8 965 0 DRAIN2
port 10 nsew
rlabel metal1 35 1496 77 1503 0 VTUN
port 11 nsew
rlabel metal1 405 1495 428 1503 0 GATE1
port 12 nsew
rlabel metal1 1101 1495 1129 1503 0 VINJ
port 13 nsew
rlabel metal2 1191 1168 1214 1192 0 VIN11
port 14 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
