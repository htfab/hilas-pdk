magic
tech sky130A
timestamp 1628698514
<< error_p >>
rect -454 43 -453 44
rect -426 43 -425 44
rect -375 43 -374 44
rect -347 43 -346 44
rect -296 43 -295 44
rect -268 43 -267 44
rect -217 43 -216 44
rect -189 43 -188 44
rect -455 42 -454 43
rect -425 42 -424 43
rect -376 42 -375 43
rect -346 42 -345 43
rect -297 42 -296 43
rect -267 42 -266 43
rect -218 42 -217 43
rect -188 42 -187 43
rect -455 14 -454 15
rect -425 14 -424 15
rect -376 14 -375 15
rect -346 14 -345 15
rect -297 14 -296 15
rect -267 14 -266 15
rect -218 14 -217 15
rect -188 14 -187 15
rect -454 13 -453 14
rect -426 13 -425 14
rect -375 13 -374 14
rect -347 13 -346 14
rect -296 13 -295 14
rect -268 13 -267 14
rect -217 13 -216 14
rect -189 13 -188 14
<< nwell >>
rect -537 -69 -105 126
<< mvpmos >>
rect -504 43 -138 93
rect -504 14 -454 43
rect -425 14 -375 43
rect -346 14 -296 43
rect -267 14 -217 43
rect -188 14 -138 43
rect -504 -36 -138 14
<< mvpdiff >>
rect -454 37 -425 43
rect -454 20 -448 37
rect -431 20 -425 37
rect -454 14 -425 20
rect -375 37 -346 43
rect -375 20 -369 37
rect -352 20 -346 37
rect -375 14 -346 20
rect -296 37 -267 43
rect -296 20 -290 37
rect -273 20 -267 37
rect -296 14 -267 20
rect -217 37 -188 43
rect -217 20 -211 37
rect -194 20 -188 37
rect -217 14 -188 20
<< mvpdiffc >>
rect -448 20 -431 37
rect -369 20 -352 37
rect -290 20 -273 37
rect -211 20 -194 37
<< poly >>
rect -518 93 -124 106
rect -518 -36 -504 93
rect -138 -36 -124 93
rect -518 -50 -124 -36
<< locali >>
rect -512 71 -132 98
rect -512 54 -329 71
rect -312 54 -132 71
rect -512 37 -132 54
rect -512 20 -448 37
rect -431 20 -369 37
rect -352 36 -290 37
rect -352 20 -329 36
rect -512 19 -329 20
rect -312 20 -290 36
rect -273 20 -211 37
rect -194 20 -132 37
rect -312 19 -132 20
rect -512 2 -132 19
rect -512 -15 -329 2
rect -312 -15 -132 2
rect -512 -43 -132 -15
<< viali >>
rect -329 54 -312 71
rect -329 19 -312 36
rect -329 -15 -312 2
<< metal1 >>
rect -333 71 -309 77
rect -333 54 -329 71
rect -312 54 -309 71
rect -333 36 -309 54
rect -333 19 -329 36
rect -312 19 -309 36
rect -333 13 -309 19
rect -332 2 -309 13
rect -332 -15 -329 2
rect -312 -15 -309 2
rect -332 -52 -309 -15
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
