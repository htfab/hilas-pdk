magic
tech sky130A
timestamp 1627063084
<< nwell >>
rect 0 -80 251 79
<< mvpmos >>
rect 65 15 115 46
rect 136 -47 186 -16
<< mvpdiff >>
rect 34 39 65 46
rect 34 22 42 39
rect 59 22 65 39
rect 34 15 65 22
rect 115 40 149 46
rect 115 23 121 40
rect 138 23 149 40
rect 115 15 149 23
rect 105 -24 136 -16
rect 105 -41 111 -24
rect 129 -41 136 -24
rect 105 -47 136 -41
rect 186 -22 218 -16
rect 186 -39 192 -22
rect 210 -39 218 -22
rect 186 -47 218 -39
<< mvpdiffc >>
rect 42 22 59 39
rect 121 23 138 40
rect 111 -41 129 -24
rect 192 -39 210 -22
<< mvnsubdiff >>
rect 35 -24 105 -16
rect 35 -41 61 -24
rect 78 -41 105 -24
rect 35 -47 105 -41
<< mvnsubdiffcont >>
rect 61 -41 78 -24
<< poly >>
rect 65 48 236 64
rect 65 46 115 48
rect 209 20 236 48
rect 65 0 115 15
rect 209 3 214 20
rect 231 3 236 20
rect 136 -16 186 -1
rect 209 -5 236 3
rect 136 -50 186 -47
rect 136 -65 266 -50
<< polycont >>
rect 214 3 231 20
<< locali >>
rect 128 47 351 55
rect 128 40 145 47
rect 34 22 42 39
rect 59 22 67 39
rect 113 23 121 40
rect 138 30 145 40
rect 162 38 351 47
rect 162 30 173 38
rect 138 23 173 30
rect 41 12 59 22
rect 58 -5 59 12
rect 41 -23 59 -5
rect 206 3 214 20
rect 231 3 239 20
rect 206 -22 231 3
rect 58 -24 59 -23
rect 58 -40 61 -24
rect 41 -41 61 -40
rect 78 -41 111 -24
rect 129 -41 137 -24
rect 184 -39 192 -22
rect 210 -32 231 -22
rect 210 -33 248 -32
rect 210 -39 266 -33
rect 192 -50 266 -39
<< viali >>
rect 145 30 162 47
rect 41 -5 58 12
rect 41 -40 58 -23
<< metal1 >>
rect 34 12 63 79
rect 138 52 170 55
rect 138 26 141 52
rect 167 26 170 52
rect 138 25 170 26
rect 34 -5 41 12
rect 58 -5 63 12
rect 34 -23 63 -5
rect 34 -40 41 -23
rect 58 -40 63 -23
rect 34 -80 63 -40
<< via1 >>
rect 141 47 167 52
rect 141 30 145 47
rect 145 30 162 47
rect 162 30 167 47
rect 141 26 167 30
<< metal2 >>
rect 138 47 141 52
rect 7 27 141 47
rect 138 26 141 27
rect 167 26 170 52
use sky130_hilas_StepUpDigitalPart1  StepUpDigitalPart1_0
timestamp 1624113415
transform 1 0 -12 0 1 -40
box 278 -40 892 119
<< labels >>
rlabel metal2 7 27 14 47 0 Output
rlabel metal1 34 71 63 79 0 Vinj
rlabel metal1 34 -80 63 -72 0 Vinj
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
