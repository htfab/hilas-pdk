magic
tech sky130A
timestamp 1634057735
<< nwell >>
rect 0 28 417 235
<< pmos >>
rect 57 145 310 216
rect 57 46 310 116
<< pdiff >>
rect 19 210 57 216
rect 19 151 28 210
rect 46 151 57 210
rect 19 145 57 151
rect 310 208 355 216
rect 310 145 328 208
rect 319 116 328 145
rect 21 110 57 116
rect 21 51 28 110
rect 46 51 57 110
rect 21 46 57 51
rect 310 51 328 116
rect 346 51 355 208
rect 310 46 355 51
<< pdiffc >>
rect 28 151 46 210
rect 28 51 46 110
rect 328 51 346 208
<< nsubdiff >>
rect 355 206 397 216
rect 355 51 367 206
rect 385 51 397 206
rect 355 46 397 51
<< nsubdiffcont >>
rect 367 51 385 206
<< poly >>
rect 57 216 310 232
rect 57 116 310 145
rect 57 22 310 46
rect 57 5 65 22
rect 302 5 310 22
rect 57 0 310 5
<< polycont >>
rect 65 5 302 22
<< locali >>
rect 28 210 46 218
rect 28 143 46 151
rect 319 208 389 220
rect 28 110 46 118
rect 28 43 46 51
rect 319 51 328 208
rect 346 206 389 208
rect 346 189 348 206
rect 365 189 367 206
rect 346 169 367 189
rect 346 152 348 169
rect 365 152 367 169
rect 346 133 367 152
rect 346 116 348 133
rect 365 116 367 133
rect 346 97 367 116
rect 346 80 348 97
rect 365 80 367 97
rect 346 61 367 80
rect 346 51 348 61
rect 319 44 348 51
rect 365 51 367 61
rect 385 51 389 206
rect 365 44 389 51
rect 28 22 45 43
rect 319 40 389 44
rect 28 5 65 22
rect 302 5 310 22
<< viali >>
rect 348 189 365 206
rect 348 152 365 169
rect 348 116 365 133
rect 348 80 365 97
rect 348 44 365 61
<< metal1 >>
rect 334 206 377 223
rect 334 189 348 206
rect 365 189 377 206
rect 334 169 377 189
rect 334 152 348 169
rect 365 152 377 169
rect 334 133 377 152
rect 334 116 348 133
rect 365 116 377 133
rect 334 97 377 116
rect 334 80 348 97
rect 365 80 377 97
rect 334 61 377 80
rect 334 44 348 61
rect 365 44 377 61
rect 334 34 377 44
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
