magic
tech sky130A
timestamp 1627744303
<< error_s >>
rect -994 528 -944 539
rect -922 528 -872 539
rect -872 497 -840 498
rect -994 486 -944 497
rect -922 486 -872 497
rect -922 466 -872 478
rect -953 436 -949 466
rect -872 465 -843 466
rect -922 424 -872 436
rect -332 421 -315 423
rect -734 418 -717 420
rect -332 402 -315 404
rect -734 399 -717 401
rect -922 384 -872 396
rect -953 354 -949 384
rect -872 354 -843 355
rect -922 342 -872 354
rect -994 323 -944 334
rect -922 323 -872 334
rect -872 322 -840 323
rect -735 300 -718 302
rect -333 294 -316 296
rect -994 281 -944 292
rect -922 281 -872 292
rect -735 281 -718 283
rect -333 275 -316 277
rect -735 266 -718 268
rect -333 260 -316 262
rect -735 247 -718 249
rect -333 241 -316 243
rect -994 227 -944 238
rect -922 227 -872 238
rect -735 232 -718 234
rect -333 226 -316 228
rect -735 213 -718 215
rect -333 207 -316 209
rect -872 196 -840 197
rect -994 185 -944 196
rect -922 185 -872 196
rect -333 192 -316 194
rect -922 165 -872 177
rect -953 135 -949 165
rect -872 164 -843 165
rect -922 123 -872 135
rect -922 84 -872 96
rect -953 54 -949 84
rect -872 54 -843 55
rect -922 42 -872 54
rect -994 23 -944 34
rect -922 23 -872 34
rect -872 22 -840 23
rect -994 -19 -944 -8
rect -922 -19 -872 -8
<< nwell >>
rect -1101 561 -805 562
rect -1101 546 -1060 561
rect -532 552 -494 562
rect -129 548 -89 562
rect -1101 545 -1042 546
rect -1101 369 -1060 545
rect -1112 254 -1060 369
rect -1101 -42 -1060 254
<< poly >>
rect 209 516 229 562
rect 209 -43 229 -18
<< locali >>
rect -1115 -22 -1097 67
<< metal1 >>
rect -1025 555 -1009 562
rect -984 555 -965 562
rect -944 555 -928 562
rect -532 552 -494 562
rect -129 534 -89 562
rect 131 516 154 562
rect 257 516 280 562
rect -782 430 -761 504
rect -1112 254 -1091 369
rect -784 93 -768 243
rect 257 127 280 132
rect 253 126 281 127
rect 253 124 283 126
rect 253 97 254 124
rect 281 97 283 124
rect 253 94 283 97
rect -532 -43 -494 -33
rect 131 -43 154 -18
rect 257 -43 280 -18
<< via1 >>
rect 254 97 281 124
<< metal2 >>
rect -758 512 7 531
rect -1116 494 -1061 512
rect -758 510 24 512
rect -14 491 24 510
rect -1112 418 -1097 469
rect -65 457 -50 469
rect -65 437 56 457
rect 170 426 296 442
rect -1112 402 -769 418
rect -1112 352 -1086 378
rect -1107 351 -1090 352
rect -55 351 66 371
rect 170 333 296 349
rect -1118 308 -1061 326
rect -791 304 -768 305
rect -791 301 -34 304
rect -791 284 -28 301
rect -791 274 -767 284
rect -1112 256 -767 274
rect -47 264 24 284
rect -1112 254 -775 256
rect -777 234 -32 236
rect -777 214 24 234
rect -777 213 -745 214
rect -1116 193 -1061 211
rect -1116 192 -1100 193
rect -1118 118 -1098 168
rect -56 152 44 168
rect 170 149 296 165
rect 251 124 284 125
rect -1118 98 -763 118
rect 251 116 254 124
rect -384 99 254 116
rect 251 97 254 99
rect 281 97 284 124
rect 251 96 284 97
rect -1119 47 -1091 74
rect -55 54 45 71
rect 172 56 296 72
rect -55 53 39 54
rect -1114 26 -1098 27
rect -1114 8 -1061 26
rect -32 8 23 9
rect -790 -14 23 8
rect -790 -15 -31 -14
rect -790 -16 -713 -15
rect -790 -20 -766 -16
rect -1114 -40 -766 -20
rect -1114 -41 -847 -40
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1627744303
transform 1 0 -1107 0 1 59
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1627744303
transform 1 0 -1102 0 1 -26
box -14 -15 20 18
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1627744303
transform 1 0 -1107 0 1 258
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_3
timestamp 1627744303
transform 1 0 -1105 0 1 359
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1627744303
transform 1 0 -776 0 1 514
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_2
timestamp 1627744303
transform 1 0 -778 0 1 409
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_5
timestamp 1627744303
transform 1 0 -794 0 1 103
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_4
timestamp 1627744303
transform 1 0 -778 0 1 221
box -9 -10 23 22
use sky130_hilas_WTA4stage01  sky130_hilas_WTA4stage01_0
timestamp 1627744303
transform 1 0 67 0 1 -19
box -54 1 229 535
use sky130_hilas_swc4x1BiasCell  sky130_hilas_swc4x1BiasCell_0
timestamp 1627744303
transform -1 0 -317 0 1 339
box -266 -382 745 223
<< labels >>
rlabel metal2 289 426 296 442 0 OUTPUT1
port 4 nsew analog default
rlabel metal2 291 333 296 349 0 OUTPUT2
port 5 nsew analog default
rlabel metal2 291 149 296 165 0 OUTPUT3
port 6 nsew analog default
rlabel metal2 291 56 296 72 0 OUTPUT4
port 7 nsew analog default
rlabel metal1 257 556 280 562 0 VGND
port 1 nsew ground default
rlabel metal1 257 -43 280 -37 0 VGND
port 1 nsew ground default
rlabel metal2 -1112 449 -1097 469 0 INPUT1
port 8 nsew analog default
rlabel metal2 -1112 352 -1086 378 0 INPUT2
port 9 nsew analog default
rlabel metal2 -1118 151 -1098 168 0 INPUT3
port 10 nsew analog default
rlabel metal2 -1119 47 -1091 74 0 INPUT4
port 11 nsew analog default
rlabel metal2 -1100 494 -1088 512 0 DRAIN1
port 12 nsew
rlabel metal2 -1100 308 -1088 326 0 DRAIN2
port 13 nsew
rlabel metal2 -1100 193 -1088 211 0 DRAIN3
port 14 nsew
rlabel metal2 -1100 8 -1088 26 0 DRAIN4
port 15 nsew
rlabel metal1 -531 552 -495 562 0 GATE1
port 16 nsew
rlabel metal1 -129 548 -89 562 0 VTUN
port 17 nsew
rlabel metal1 131 -43 154 -37 0 WTAMIDDLENODE
port 18 nsew
rlabel metal1 131 556 154 562 0 WTAMIDDLENODE
port 18 nsew
rlabel metal1 -984 555 -965 562 0 COLSEL1
port 19 nsew
rlabel metal1 -1025 555 -1009 562 0 VINJ
port 21 nsew
rlabel metal1 -944 555 -928 562 0 VPWR
port 20 nsew
<< end >>
