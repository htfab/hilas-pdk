magic
tech sky130A
timestamp 1634057750
<< checkpaint >>
rect 822 1716 2255 1721
rect 703 1543 2255 1716
rect 703 1362 2655 1543
rect 411 97 2655 1362
rect 411 -189 2255 97
rect 411 -194 2186 -189
rect 411 -630 1927 -194
<< error_s >>
rect 912 657 931 671
rect 956 657 972 671
rect 752 615 773 632
rect 999 617 1013 635
rect 731 444 752 461
rect 752 410 766 424
rect 999 422 1013 440
rect 898 381 944 384
rect 891 376 944 381
rect 888 371 944 376
rect 888 368 901 371
rect 891 367 901 368
rect 896 364 901 367
rect 908 370 944 371
rect 908 369 929 370
rect 931 369 944 370
rect 908 367 944 369
rect 908 366 913 367
rect 941 366 944 367
rect 956 366 972 380
rect 908 364 918 366
rect 896 359 918 364
rect 929 359 944 366
rect 896 358 904 359
rect 905 354 918 359
rect 905 351 913 354
rect 931 346 934 356
rect 749 308 764 312
rect 749 295 773 308
rect 752 291 773 295
rect 997 293 1011 311
rect 731 119 752 136
rect 997 97 1011 115
rect 912 60 931 74
rect 956 60 972 74
<< nwell >>
rect 58 518 117 534
rect 432 512 543 539
rect 752 420 761 428
rect 896 370 913 376
rect 896 369 931 370
rect 896 359 913 369
rect 930 359 931 369
rect 58 194 117 209
rect 432 192 543 211
<< psubdiff >>
rect 258 523 283 546
rect 258 506 262 523
rect 279 506 283 523
rect 660 520 685 548
rect 258 478 283 506
rect 660 503 664 520
rect 681 503 685 520
rect 660 477 685 503
rect 258 396 284 438
rect 258 379 263 396
rect 280 379 284 396
rect 258 362 284 379
rect 258 345 263 362
rect 280 345 284 362
rect 258 328 284 345
rect 258 311 263 328
rect 280 311 284 328
rect 258 300 284 311
rect 660 402 687 423
rect 660 385 665 402
rect 682 385 687 402
rect 660 368 687 385
rect 660 351 665 368
rect 682 351 687 368
rect 660 334 687 351
rect 660 317 665 334
rect 682 317 687 334
rect 263 296 280 300
rect 660 299 687 317
<< mvnsubdiff >>
rect 58 518 117 534
rect 432 512 543 539
rect 58 194 117 209
rect 432 192 543 211
<< psubdiffcont >>
rect 262 506 279 523
rect 664 503 681 520
rect 263 379 280 396
rect 263 345 280 362
rect 263 311 280 328
rect 665 385 682 402
rect 665 351 682 368
rect 665 317 682 334
<< poly >>
rect 584 596 752 613
rect 159 568 392 592
rect 157 446 392 470
rect 584 444 752 461
rect 891 366 896 367
rect 913 369 931 370
rect 929 367 931 369
rect 913 366 941 367
rect 929 359 931 366
rect 157 266 394 290
rect 584 272 752 289
rect 159 134 396 158
rect 584 119 752 136
<< polycont >>
rect 896 359 913 376
<< locali >>
rect 262 523 279 525
rect 664 520 681 522
rect 263 362 280 379
rect 263 328 280 332
rect 665 368 682 385
rect 887 359 896 376
rect 665 334 682 336
<< viali >>
rect 262 525 279 542
rect 262 489 279 506
rect 664 522 681 539
rect 664 486 681 503
rect 263 396 280 413
rect 263 345 280 349
rect 263 332 280 345
rect 263 311 280 313
rect 263 296 280 311
rect 665 402 682 419
rect 913 359 931 376
rect 665 351 682 353
rect 665 336 682 351
rect 665 300 682 317
<< metal1 >>
rect 36 41 76 691
rect 257 542 284 691
rect 441 654 479 691
rect 257 525 262 542
rect 279 525 284 542
rect 257 506 284 525
rect 257 489 262 506
rect 279 489 284 506
rect 257 413 284 489
rect 257 396 263 413
rect 280 396 284 413
rect 257 349 284 396
rect 257 332 263 349
rect 280 332 284 349
rect 257 313 284 332
rect 257 296 263 313
rect 280 296 284 313
rect 257 217 284 296
rect 660 539 685 691
rect 875 657 891 664
rect 912 657 931 664
rect 956 657 972 664
rect 660 522 664 539
rect 681 522 685 539
rect 660 503 685 522
rect 660 486 664 503
rect 681 486 685 503
rect 660 419 685 486
rect 660 402 665 419
rect 682 402 685 419
rect 660 353 685 402
rect 910 376 934 379
rect 891 367 913 376
rect 875 366 913 367
rect 891 359 913 366
rect 931 359 934 376
rect 956 366 972 367
rect 910 356 934 359
rect 660 336 665 353
rect 682 336 685 353
rect 920 346 931 356
rect 660 317 685 336
rect 660 300 665 317
rect 682 300 685 317
rect 660 220 685 300
rect 659 217 687 220
rect 255 214 286 217
rect 255 188 257 214
rect 284 188 286 214
rect 658 216 688 217
rect 658 190 660 216
rect 686 190 688 216
rect 658 189 688 190
rect 255 186 286 188
rect 659 187 687 189
rect 257 41 284 186
rect 441 41 479 69
rect 660 41 685 187
rect 875 60 891 67
rect 912 60 931 67
rect 956 60 972 67
<< via1 >>
rect 257 188 284 214
rect 660 190 686 216
<< metal2 >>
rect 999 617 1008 635
rect 1 573 762 592
rect 999 574 1008 592
rect 1 465 764 483
rect 999 465 1008 483
rect 752 421 761 424
rect 999 422 1008 440
rect 752 410 764 421
rect 749 295 764 312
rect 997 293 1008 311
rect 1 254 48 270
rect 2 253 48 254
rect 78 251 764 268
rect 997 250 1008 268
rect 657 216 689 217
rect 254 188 257 214
rect 284 211 287 214
rect 657 211 660 216
rect 284 194 660 211
rect 284 188 287 194
rect 657 190 660 194
rect 686 190 689 216
rect 657 189 689 190
rect 1 155 764 172
rect 997 140 1008 158
rect 997 97 1008 115
use sky130_hilas_horizPcell01d3  sky130_hilas_horizPcell01d3_2
timestamp 1634057722
transform 1 0 1041 0 -1 408
box 0 0 256 191
use sky130_hilas_horizPcell01d3  sky130_hilas_horizPcell01d3_1
timestamp 1634057722
transform 1 0 1041 0 1 0
box 0 0 256 191
use sky130_hilas_horizPcell01d3  sky130_hilas_horizPcell01d3_3
timestamp 1634057722
transform 1 0 1041 0 -1 732
box 0 0 256 191
use sky130_hilas_horizPcell01d3  sky130_hilas_horizPcell01d3_0
timestamp 1634057722
transform 1 0 1041 0 1 325
box 0 0 256 191
use sky130_hilas_wellContact  sky130_hilas_wellContact_1
timestamp 1634057703
transform 1 0 1449 0 1 734
box 0 0 173 186
use sky130_hilas_wellContact  sky130_hilas_wellContact_0
timestamp 1634057703
transform 1 0 1852 0 1 727
box 0 0 173 186
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_0
timestamp 1634057705
transform 1 0 1333 0 1 436
box 0 0 223 186
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_2
timestamp 1634057705
transform 1 0 1333 0 1 756
box 0 0 223 186
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_1
timestamp 1634057705
transform 1 0 1333 0 1 571
box 0 0 223 186
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_3
timestamp 1634057705
transform 1 0 1333 0 1 900
box 0 0 223 186
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_1
timestamp 1634057702
transform 1 0 1452 0 1 441
box 0 0 173 190
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_2
timestamp 1634057702
transform 1 0 1452 0 1 765
box 0 0 173 190
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_0
timestamp 1634057702
transform 1 0 1452 0 1 576
box 0 0 173 190
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_3
timestamp 1634057702
transform 1 0 1452 0 1 901
box 0 0 173 190
<< labels >>
rlabel metal2 1 254 13 270 0 ROW3
port 3 nsew analog default
rlabel metal2 1 156 15 171 0 ROW4
port 4 nsew analog default
rlabel metal1 36 650 76 664 0 VTUN
port 5 nsew analog default
rlabel metal1 36 59 76 69 0 VTUN
port 5 nsew analog default
rlabel metal1 441 59 479 69 0 GATE1
port 6 nsew analog default
rlabel metal1 441 654 479 664 0 GATE1
port 6 nsew analog default
rlabel metal1 956 657 972 664 0 VINJ
port 7 nsew power default
rlabel metal1 875 657 891 664 0 VPWR
port 8 nsew power default
rlabel metal1 912 657 931 664 0 COLSEL1
rlabel metal1 956 60 972 67 0 VINJ
port 7 nsew power default
rlabel metal1 875 60 891 67 0 VPWR
port 8 nsew power default
rlabel metal1 912 60 931 67 0 COLSEL1
port 9 nsew analog default
rlabel metal1 257 656 284 664 0 VGND
port 18 nsew
rlabel metal1 660 659 685 664 0 VGND
port 18 nsew
rlabel metal1 257 59 284 66 0 VGND
port 18 nsew
rlabel metal1 660 59 685 66 0 VGND
port 18 nsew
rlabel metal2 997 250 1008 268 0 ROW3
port 3 nsew
rlabel metal2 997 293 1008 311 0 DRAIN3
port 19 nsew
rlabel metal2 997 97 1008 115 0 DRAIN4
port 20 nsew
rlabel metal2 997 140 1008 158 0 ROW4
port 4 nsew
rlabel metal2 999 617 1008 635 0 DRAIN1
port 21 nsew
rlabel metal2 999 574 1008 592 0 ROW1
port 1 nsew
rlabel metal2 999 465 1008 483 0 ROW2
port 2 nsew
rlabel metal2 999 422 1008 440 0 DRAIN2
port 22 nsew
rlabel space 0 573 12 592 0 ROW1
port 1 nsew
rlabel metal2 1 465 7 483 0 ROW2
port 2 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
