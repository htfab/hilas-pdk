* NGSPICE file created from /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_Tgate4Double01.ext - technology: sky130A

.subckt sky130_hilas_TgateDouble01 VSUBS a_n40_n314# a_n468_n112# output w_n502_n362#
+ a_290_n314#
X0 a_n196_n192# a_n468_n112# w_n502_n362# w_n502_n362# sky130_fd_pr__pfet_01v8 w=320000u l=400000u
X1 VSUBS a_n468_n112# a_n196_n192# VSUBS sky130_fd_pr__nfet_01v8 w=300000u l=400000u
X2 output a_n468_n112# a_n40_n314# VSUBS sky130_fd_pr__nfet_01v8 w=310000u l=400000u
X3 output a_n468_n112# a_290_n314# w_n502_n362# sky130_fd_pr__pfet_01v8 w=310000u l=400000u
X4 output a_n196_n192# a_n40_n314# w_n502_n362# sky130_fd_pr__pfet_01v8 w=310000u l=400000u
X5 output a_n196_n192# a_290_n314# VSUBS sky130_fd_pr__nfet_01v8 w=310000u l=400000u
.ends

.subckt home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_Tgate4Double01
+ Vdd Input1_1 Input2_1 Select1 Select2 Input2_2 Input1_2 Select3 Input2_3 Select4
+ Input2_4 Input1_4 Output4 Output3 Output2 Output1
Xsky130_hilas_TgateDouble01_0 Vdd Input1_1 Select1 Output1 Vdd Input2_1 sky130_hilas_TgateDouble01
Xsky130_hilas_TgateDouble01_1 Vdd Input1_4 Select4 Output4 Vdd Input2_4 sky130_hilas_TgateDouble01
Xsky130_hilas_TgateDouble01_2 Vdd Input1_3 Select3 Output3 Vdd Input2_3 sky130_hilas_TgateDouble01
Xsky130_hilas_TgateDouble01_3 Vdd Input1_2 Select2 Output2 Vdd Input2_2 sky130_hilas_TgateDouble01
.ends

