magic
tech sky130A
timestamp 1628698551
<< psubdiff >>
rect -131 148 491 156
rect -131 131 -116 148
rect -99 131 491 148
rect -131 124 491 131
<< psubdiffcont >>
rect -116 131 -99 148
<< poly >>
rect -119 193 -75 206
rect -119 176 -106 193
rect -89 176 -75 193
rect -119 164 -75 176
rect 438 195 484 206
rect 438 178 453 195
rect 470 178 487 195
rect 438 164 484 178
<< polycont >>
rect -106 176 -89 193
rect 453 178 470 195
<< npolyres >>
rect -75 164 438 206
<< locali >>
rect -89 176 -81 193
rect 445 178 453 195
rect 445 176 487 178
rect -127 131 -116 148
<< viali >>
rect -123 176 -106 193
rect 470 178 487 195
rect -99 131 -82 148
<< metal1 >>
rect -143 193 -86 198
rect -143 176 -123 193
rect -106 176 -86 193
rect -143 171 -86 176
rect 453 195 506 201
rect 453 178 470 195
rect 487 178 506 195
rect 453 171 506 178
rect -102 148 -76 151
rect -128 144 -99 148
rect -143 131 -99 144
rect -82 131 -76 148
rect -143 128 -76 131
<< labels >>
rlabel metal1 -142 171 -133 198 0 TERM1
port 1 nsew
rlabel metal1 494 171 506 201 0 TERM2
port 2 nsew
rlabel metal1 -143 128 -134 144 0 VGND
port 3 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
