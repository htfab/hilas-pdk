VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_hilas_TA2Cell_1FG_Strong
  CLASS CORE ;
  FOREIGN sky130_hilas_TA2Cell_1FG_Strong ;
  ORIGIN 0.000 0.000 ;
  SIZE 32.050 BY 9.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 14.710 5.900 15.130 6.050 ;
        RECT 15.740 5.900 16.160 6.050 ;
        RECT 14.710 5.760 16.160 5.900 ;
    END
  END VTUN
  PIN PROG
    PORT
      LAYER met1 ;
        RECT 7.470 5.990 7.680 6.050 ;
    END
  END PROG
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT 19.440 5.970 19.670 6.050 ;
    END
  END GATE1
  PIN VIN11
    PORT
      LAYER met1 ;
        RECT 6.590 5.940 6.800 6.050 ;
    END
  END VIN11
  PIN VINJ
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 1.770 5.970 2.080 6.160 ;
        RECT 4.150 5.970 4.470 6.030 ;
        RECT 1.770 5.910 11.520 5.970 ;
        RECT 26.420 5.910 26.740 6.030 ;
        RECT 1.770 5.830 26.740 5.910 ;
        RECT 1.800 5.780 26.740 5.830 ;
        RECT 4.150 5.730 26.740 5.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 26.400 6.030 26.680 6.050 ;
        RECT 26.400 5.970 26.740 6.030 ;
        RECT 26.420 5.730 26.740 5.970 ;
      LAYER via ;
        RECT 26.450 5.750 26.710 6.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 26.400 0.000 26.680 0.050 ;
    END
  END VINJ
  PIN VIN22
    ANTENNAGATEAREA 4.153100 ;
    ANTENNADIFFAREA 8.050300 ;
    PORT
      LAYER nwell ;
        RECT 27.570 6.050 30.880 9.870 ;
        RECT 26.920 6.040 32.050 6.050 ;
        RECT 26.910 3.830 32.050 6.040 ;
        RECT 26.910 0.000 28.770 3.830 ;
        RECT 30.770 0.000 32.050 3.830 ;
      LAYER met2 ;
        RECT 29.490 7.010 29.810 7.270 ;
        RECT 29.530 6.990 30.710 7.010 ;
        RECT 29.530 6.730 30.750 6.990 ;
        RECT 29.530 6.670 30.710 6.730 ;
        RECT 29.490 6.660 30.710 6.670 ;
        RECT 29.490 6.410 29.810 6.660 ;
        RECT 28.160 6.030 28.470 6.040 ;
        RECT 27.590 6.020 28.470 6.030 ;
        RECT 27.520 5.780 28.470 6.020 ;
        RECT 28.160 5.710 28.470 5.780 ;
        RECT 29.130 5.710 29.440 5.760 ;
        RECT 31.380 5.710 31.690 5.810 ;
        RECT 28.550 5.590 28.860 5.660 ;
        RECT 29.130 5.590 31.690 5.710 ;
        RECT 28.550 5.480 31.690 5.590 ;
        RECT 28.550 5.380 30.880 5.480 ;
        RECT 28.550 5.330 28.860 5.380 ;
        RECT 28.310 5.170 28.620 5.210 ;
        RECT 28.130 5.030 28.850 5.170 ;
        RECT 29.080 5.030 29.390 5.110 ;
        RECT 28.130 4.920 29.390 5.030 ;
        RECT 28.310 4.880 29.390 4.920 ;
        RECT 28.580 4.820 29.390 4.880 ;
        RECT 28.580 4.810 28.850 4.820 ;
        RECT 29.080 4.780 29.390 4.820 ;
        RECT 27.190 4.530 27.500 4.670 ;
        RECT 26.840 4.490 27.500 4.530 ;
        RECT 28.400 4.500 28.710 4.640 ;
        RECT 28.400 4.490 30.880 4.500 ;
        RECT 19.350 4.340 30.880 4.490 ;
        RECT 26.840 4.310 27.190 4.340 ;
        RECT 28.400 4.320 30.880 4.340 ;
        RECT 28.400 4.310 28.710 4.320 ;
        RECT 28.650 4.240 28.850 4.250 ;
        RECT 28.650 4.230 28.870 4.240 ;
        RECT 29.080 4.230 29.390 4.270 ;
        RECT 28.650 4.160 29.390 4.230 ;
        RECT 28.360 4.140 29.390 4.160 ;
        RECT 28.310 4.020 29.390 4.140 ;
        RECT 28.310 3.900 28.870 4.020 ;
        RECT 29.080 3.940 29.390 4.020 ;
        RECT 28.310 3.890 28.780 3.900 ;
        RECT 28.560 0.350 28.880 0.500 ;
        RECT 12.370 0.200 28.880 0.350 ;
        RECT 12.370 0.050 12.690 0.200 ;
        RECT 18.170 0.050 18.490 0.200 ;
    END
  END VIN22
  PIN VIN21
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT 27.920 3.350 28.230 3.390 ;
        RECT 27.600 3.340 28.260 3.350 ;
        RECT 27.600 3.110 28.700 3.340 ;
        RECT 27.920 3.060 28.230 3.110 ;
    END
  END VIN21
  PIN VPWR
    ANTENNADIFFAREA 1.373600 ;
    PORT
      LAYER met1 ;
        RECT 30.750 5.900 31.030 6.050 ;
        RECT 30.760 4.470 31.030 5.900 ;
        RECT 30.760 4.180 31.040 4.470 ;
        RECT 30.760 1.880 31.030 4.180 ;
        RECT 30.760 1.590 31.040 1.880 ;
        RECT 30.760 0.000 31.030 1.590 ;
    END
  END VPWR
  PIN VGND
    ANTENNAGATEAREA 3.745100 ;
    ANTENNADIFFAREA 3.678400 ;
    PORT
      LAYER met1 ;
        RECT 29.920 8.410 30.110 9.870 ;
        RECT 30.360 9.220 30.640 9.870 ;
        RECT 30.250 8.620 30.640 9.220 ;
        RECT 29.920 8.380 30.140 8.410 ;
        RECT 29.900 8.110 30.150 8.380 ;
        RECT 29.910 8.100 30.150 8.110 ;
        RECT 29.910 7.860 30.140 8.100 ;
        RECT 29.520 6.380 29.780 6.700 ;
        RECT 29.520 6.260 29.760 6.380 ;
        RECT 29.950 6.050 30.110 7.860 ;
        RECT 30.360 7.020 30.640 8.620 ;
        RECT 30.360 6.700 30.720 7.020 ;
        RECT 30.360 6.050 30.640 6.700 ;
        RECT 28.150 5.710 28.470 6.030 ;
        RECT 29.950 5.830 30.640 6.050 ;
        RECT 29.130 5.430 29.450 5.750 ;
        RECT 29.910 5.580 30.640 5.830 ;
        RECT 29.900 5.310 30.640 5.580 ;
        RECT 29.080 4.780 29.400 5.100 ;
        RECT 28.400 4.200 28.710 4.640 ;
        RECT 28.410 4.190 28.620 4.200 ;
        RECT 28.390 3.870 28.650 4.190 ;
        RECT 29.080 3.950 29.400 4.270 ;
        RECT 28.410 2.580 28.620 3.870 ;
        RECT 29.920 3.820 30.640 5.310 ;
        RECT 28.390 2.290 28.620 2.580 ;
        RECT 28.560 0.200 28.880 0.500 ;
        RECT 30.090 0.200 30.430 3.820 ;
        RECT 28.560 0.140 30.430 0.200 ;
        RECT 28.610 0.060 30.430 0.140 ;
        RECT 30.090 0.000 30.430 0.060 ;
      LAYER via ;
        RECT 29.520 6.410 29.780 6.670 ;
        RECT 30.460 6.730 30.720 6.990 ;
        RECT 28.180 5.740 28.440 6.000 ;
        RECT 29.160 5.460 29.420 5.720 ;
        RECT 29.110 4.810 29.370 5.070 ;
        RECT 28.430 4.350 28.690 4.610 ;
        RECT 28.390 3.900 28.650 4.160 ;
        RECT 29.110 3.980 29.370 4.240 ;
        RECT 28.590 0.220 28.850 0.480 ;
    END
  END VGND
  PIN OUTPUT2
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER met2 ;
        RECT 29.130 2.740 29.440 2.800 ;
        RECT 31.420 2.740 31.730 2.870 ;
        RECT 29.130 2.520 32.050 2.740 ;
        RECT 29.130 2.470 29.440 2.520 ;
    END
  END OUTPUT2
  PIN OUTPUT1
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER met2 ;
        RECT 29.130 3.570 29.440 3.620 ;
        RECT 31.430 3.570 31.740 3.590 ;
        RECT 29.130 3.340 32.050 3.570 ;
        RECT 29.130 3.290 29.440 3.340 ;
        RECT 31.430 3.260 31.740 3.340 ;
    END
  END OUTPUT1
  PIN GATESEL1
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER met1 ;
        RECT 4.600 6.050 4.780 9.870 ;
        RECT 4.600 5.990 4.910 6.050 ;
        RECT 4.600 5.340 4.780 5.990 ;
        RECT 4.540 5.000 4.830 5.340 ;
        RECT 4.600 3.820 4.780 5.000 ;
    END
  END GATESEL1
  PIN GATESEL2
    PORT
      LAYER met1 ;
        RECT 25.960 0.000 26.150 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.960 5.970 26.150 6.050 ;
    END
  END GATESEL2
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 3.950 5.370 4.030 5.550 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 3.950 0.500 4.030 0.680 ;
    END
  END DRAIN2
  PIN VIN12
    PORT
      LAYER met1 ;
        RECT 6.600 0.010 6.830 0.130 ;
    END
  END VIN12
  PIN GATE2
    PORT
      LAYER met1 ;
        RECT 7.060 5.970 7.250 6.050 ;
    END
  END GATE2
  PIN RUN
    ANTENNADIFFAREA 1.850000 ;
    PORT
      LAYER met1 ;
        RECT 8.470 6.050 8.700 9.870 ;
        RECT 8.470 5.980 8.730 6.050 ;
        RECT 8.470 3.820 8.700 5.980 ;
    END
  END RUN
  OBS
      LAYER nwell ;
        RECT 0.000 3.830 3.310 9.860 ;
        RECT 5.040 7.480 7.760 9.130 ;
        RECT 9.790 9.120 11.520 9.870 ;
        RECT 5.040 7.440 7.750 7.480 ;
        RECT 5.040 6.110 7.750 6.150 ;
        RECT 5.040 6.050 7.760 6.110 ;
        RECT 3.950 6.040 7.760 6.050 ;
        RECT 4.150 5.730 4.470 6.030 ;
        RECT 5.040 4.460 7.760 6.040 ;
        RECT 9.780 5.550 11.520 9.120 ;
        RECT 9.790 3.830 11.520 5.550 ;
        RECT 19.360 9.120 21.090 9.870 ;
        RECT 19.360 5.550 21.100 9.120 ;
        RECT 23.120 7.480 25.840 9.130 ;
        RECT 23.120 7.440 25.830 7.480 ;
        RECT 23.120 6.110 25.830 6.150 ;
        RECT 19.360 3.830 21.090 5.550 ;
        RECT 23.120 4.460 25.840 6.110 ;
        RECT 26.420 5.730 26.740 6.030 ;
      LAYER li1 ;
        RECT 0.400 9.190 0.600 9.540 ;
        RECT 1.880 9.290 2.410 9.460 ;
        RECT 2.650 9.440 2.840 9.470 ;
        RECT 2.650 9.270 3.710 9.440 ;
        RECT 28.470 9.290 29.000 9.460 ;
        RECT 2.650 9.240 2.840 9.270 ;
        RECT 0.390 9.160 0.600 9.190 ;
        RECT 0.390 8.580 0.610 9.160 ;
        RECT 0.390 8.570 0.600 8.580 ;
        RECT 0.770 8.400 0.960 8.410 ;
        RECT 0.760 8.110 0.960 8.400 ;
        RECT 0.730 7.780 0.970 8.110 ;
        RECT 1.160 7.300 1.330 8.910 ;
        RECT 1.990 7.810 2.160 8.900 ;
        RECT 3.120 8.880 3.310 8.910 ;
        RECT 2.580 8.710 3.310 8.880 ;
        RECT 3.540 8.880 3.710 9.270 ;
        RECT 30.280 9.190 30.480 9.540 ;
        RECT 30.280 9.160 30.490 9.190 ;
        RECT 3.540 8.710 4.280 8.880 ;
        RECT 26.600 8.710 26.950 8.880 ;
        RECT 27.970 8.710 28.300 8.880 ;
        RECT 3.120 8.680 3.310 8.710 ;
        RECT 5.340 8.090 5.570 8.610 ;
        RECT 2.580 7.920 5.570 8.090 ;
        RECT 1.760 7.770 2.160 7.810 ;
        RECT 1.750 7.580 2.160 7.770 ;
        RECT 10.540 7.730 11.090 8.160 ;
        RECT 19.790 7.730 20.340 8.160 ;
        RECT 23.420 7.920 23.650 8.610 ;
        RECT 28.720 8.380 28.890 8.900 ;
        RECT 28.560 8.120 28.890 8.380 ;
        RECT 26.600 7.920 26.950 8.090 ;
        RECT 27.970 7.920 28.300 8.090 ;
        RECT 1.760 7.550 2.160 7.580 ;
        RECT 1.150 7.110 1.330 7.300 ;
        RECT 1.990 7.210 2.160 7.550 ;
        RECT 2.650 7.300 2.840 7.480 ;
        RECT 2.580 7.130 2.930 7.300 ;
        RECT 3.500 6.720 3.710 7.150 ;
        RECT 3.930 7.130 4.270 7.300 ;
        RECT 3.520 6.700 3.690 6.720 ;
        RECT 1.150 6.390 1.330 6.580 ;
        RECT 0.730 5.580 0.970 5.910 ;
        RECT 0.760 5.290 0.960 5.580 ;
        RECT 0.770 5.280 0.960 5.290 ;
        RECT 0.390 5.110 0.600 5.120 ;
        RECT 0.390 4.530 0.610 5.110 ;
        RECT 1.160 4.780 1.330 6.390 ;
        RECT 1.990 6.120 2.160 6.480 ;
        RECT 2.580 6.390 2.930 6.560 ;
        RECT 3.120 6.540 3.310 6.590 ;
        RECT 4.020 6.560 4.190 7.130 ;
        RECT 8.300 6.900 8.490 7.300 ;
        RECT 22.390 6.900 22.580 7.300 ;
        RECT 26.610 7.130 26.950 7.300 ;
        RECT 27.970 7.130 28.300 7.300 ;
        RECT 28.720 7.210 28.890 8.120 ;
        RECT 29.550 7.300 29.720 8.910 ;
        RECT 30.270 8.580 30.490 9.160 ;
        RECT 30.280 8.570 30.490 8.580 ;
        RECT 29.920 8.400 30.110 8.410 ;
        RECT 29.920 8.110 30.120 8.400 ;
        RECT 29.910 7.780 30.150 8.110 ;
        RECT 8.300 6.890 8.680 6.900 ;
        RECT 4.940 6.710 8.680 6.890 ;
        RECT 8.300 6.670 8.680 6.710 ;
        RECT 22.200 6.890 22.580 6.900 ;
        RECT 22.200 6.710 25.940 6.890 ;
        RECT 22.200 6.670 22.580 6.710 ;
        RECT 3.120 6.530 3.350 6.540 ;
        RECT 3.930 6.530 4.270 6.560 ;
        RECT 3.120 6.390 4.270 6.530 ;
        RECT 2.660 6.180 2.850 6.390 ;
        RECT 3.120 6.360 4.100 6.390 ;
        RECT 3.260 6.330 4.100 6.360 ;
        RECT 8.300 6.290 8.490 6.670 ;
        RECT 1.750 6.080 2.160 6.120 ;
        RECT 1.740 5.890 2.160 6.080 ;
        RECT 10.540 6.000 11.090 6.430 ;
        RECT 19.790 6.000 20.340 6.430 ;
        RECT 22.390 6.290 22.580 6.670 ;
        RECT 28.050 6.560 28.220 7.130 ;
        RECT 29.550 7.110 29.730 7.300 ;
        RECT 26.610 6.390 26.950 6.560 ;
        RECT 27.970 6.390 28.300 6.560 ;
        RECT 27.900 6.000 28.070 6.050 ;
        RECT 1.750 5.860 2.160 5.890 ;
        RECT 1.990 4.790 2.160 5.860 ;
        RECT 2.580 5.670 5.510 5.770 ;
        RECT 2.580 5.600 5.570 5.670 ;
        RECT 4.600 5.280 4.770 5.340 ;
        RECT 4.580 5.070 4.790 5.280 ;
        RECT 3.110 4.980 3.300 5.010 ;
        RECT 4.600 5.000 4.770 5.070 ;
        RECT 5.340 4.980 5.570 5.600 ;
        RECT 23.420 4.980 23.650 5.710 ;
        RECT 26.600 5.600 26.950 5.770 ;
        RECT 27.900 5.740 28.460 6.000 ;
        RECT 27.900 5.720 28.300 5.740 ;
        RECT 27.970 5.600 28.300 5.720 ;
        RECT 28.720 5.620 28.890 6.480 ;
        RECT 29.550 6.390 29.730 6.580 ;
        RECT 29.550 5.760 29.720 6.390 ;
        RECT 29.370 5.720 29.720 5.760 ;
        RECT 2.580 4.810 3.300 4.980 ;
        RECT 3.110 4.780 3.300 4.810 ;
        RECT 3.470 4.810 4.280 4.980 ;
        RECT 26.600 4.810 26.950 4.980 ;
        RECT 0.390 4.500 0.600 4.530 ;
        RECT 0.400 4.150 0.600 4.500 ;
        RECT 2.680 4.470 2.870 4.500 ;
        RECT 3.470 4.470 3.660 4.810 ;
        RECT 27.320 4.640 27.500 5.570 ;
        RECT 28.050 5.310 28.380 5.480 ;
        RECT 28.560 5.360 28.890 5.620 ;
        RECT 29.140 5.460 29.720 5.720 ;
        RECT 29.910 5.760 30.150 5.910 ;
        RECT 29.910 5.580 30.510 5.760 ;
        RECT 29.370 5.430 29.720 5.460 ;
        RECT 28.130 5.170 28.380 5.310 ;
        RECT 28.130 4.980 28.610 5.170 ;
        RECT 27.970 4.910 28.610 4.980 ;
        RECT 27.970 4.810 28.300 4.910 ;
        RECT 1.880 4.230 2.410 4.400 ;
        RECT 2.680 4.290 3.660 4.470 ;
        RECT 27.200 4.610 27.520 4.640 ;
        RECT 27.200 4.420 27.530 4.610 ;
        RECT 27.200 4.380 27.520 4.420 ;
        RECT 2.680 4.270 2.870 4.290 ;
        RECT 27.320 0.470 27.500 4.380 ;
        RECT 28.130 3.530 28.300 4.810 ;
        RECT 28.720 4.790 28.890 5.360 ;
        RECT 28.960 5.070 29.130 5.110 ;
        RECT 29.550 5.100 29.720 5.430 ;
        RECT 29.920 5.280 30.510 5.580 ;
        RECT 31.330 5.640 31.910 5.810 ;
        RECT 31.330 5.540 31.720 5.640 ;
        RECT 31.330 5.510 31.710 5.540 ;
        RECT 31.330 5.360 31.690 5.510 ;
        RECT 29.370 5.070 29.720 5.100 ;
        RECT 28.960 4.810 29.720 5.070 ;
        RECT 28.960 4.780 29.130 4.810 ;
        RECT 29.370 4.780 29.720 4.810 ;
        RECT 29.370 4.770 29.570 4.780 ;
        RECT 29.960 4.770 30.510 5.280 ;
        RECT 30.980 5.190 31.690 5.360 ;
        RECT 30.270 4.530 30.490 4.770 ;
        RECT 30.280 4.500 30.490 4.530 ;
        RECT 28.470 4.270 29.000 4.400 ;
        RECT 30.280 4.280 30.480 4.500 ;
        RECT 30.980 4.440 31.680 4.750 ;
        RECT 28.470 4.240 29.130 4.270 ;
        RECT 29.370 4.240 29.570 4.280 ;
        RECT 28.470 4.230 29.570 4.240 ;
        RECT 28.960 3.980 29.570 4.230 ;
        RECT 28.960 3.940 29.130 3.980 ;
        RECT 29.370 3.950 29.570 3.980 ;
        RECT 29.370 3.590 29.570 3.620 ;
        RECT 27.930 3.330 28.250 3.360 ;
        RECT 29.140 3.330 29.570 3.590 ;
        RECT 27.930 3.140 28.260 3.330 ;
        RECT 29.370 3.290 29.570 3.330 ;
        RECT 29.960 3.290 30.510 4.280 ;
        RECT 30.830 4.210 31.680 4.440 ;
        RECT 30.980 3.870 31.680 4.210 ;
        RECT 31.440 3.510 31.760 3.550 ;
        RECT 31.440 3.450 31.770 3.510 ;
        RECT 30.970 3.320 31.770 3.450 ;
        RECT 30.970 3.290 31.760 3.320 ;
        RECT 30.970 3.270 31.670 3.290 ;
        RECT 27.930 3.100 28.250 3.140 ;
        RECT 27.930 3.020 28.100 3.100 ;
        RECT 27.880 2.850 28.100 3.020 ;
        RECT 27.880 2.690 28.050 2.850 ;
        RECT 29.370 2.760 29.570 2.800 ;
        RECT 28.410 2.430 28.600 2.550 ;
        RECT 29.140 2.500 29.570 2.760 ;
        RECT 29.370 2.470 29.570 2.500 ;
        RECT 28.050 2.320 28.600 2.430 ;
        RECT 28.050 2.260 28.590 2.320 ;
        RECT 28.130 0.480 28.300 2.260 ;
        RECT 28.960 2.110 29.130 2.150 ;
        RECT 29.370 2.110 29.570 2.140 ;
        RECT 28.960 1.850 29.570 2.110 ;
        RECT 28.960 1.820 29.130 1.850 ;
        RECT 29.370 1.810 29.570 1.850 ;
        RECT 29.960 1.810 30.510 2.800 ;
        RECT 31.430 2.790 31.750 2.830 ;
        RECT 30.970 2.610 31.760 2.790 ;
        RECT 31.430 2.600 31.760 2.610 ;
        RECT 31.430 2.570 31.750 2.600 ;
        RECT 30.980 1.850 31.680 2.190 ;
        RECT 30.830 1.620 31.680 1.850 ;
        RECT 28.960 1.280 29.130 1.310 ;
        RECT 29.370 1.280 29.570 1.320 ;
        RECT 28.960 1.020 29.570 1.280 ;
        RECT 28.960 0.980 29.130 1.020 ;
        RECT 29.370 0.990 29.570 1.020 ;
        RECT 29.370 0.630 29.570 0.660 ;
        RECT 29.140 0.370 29.570 0.630 ;
        RECT 29.370 0.330 29.570 0.370 ;
        RECT 29.960 0.330 30.510 1.320 ;
        RECT 30.980 1.310 31.680 1.620 ;
        RECT 30.980 0.700 31.690 0.870 ;
        RECT 31.330 0.420 31.690 0.700 ;
        RECT 31.330 0.250 31.910 0.420 ;
      LAYER mcon ;
        RECT 2.230 9.290 2.410 9.460 ;
        RECT 2.660 9.270 2.830 9.440 ;
        RECT 0.420 8.990 0.590 9.160 ;
        RECT 0.770 8.150 0.950 8.340 ;
        RECT 3.130 8.710 3.300 8.880 ;
        RECT 30.290 8.990 30.460 9.160 ;
        RECT 5.370 8.410 5.540 8.580 ;
        RECT 23.450 8.410 23.620 8.580 ;
        RECT 5.370 7.960 5.540 8.130 ;
        RECT 1.850 7.590 2.020 7.760 ;
        RECT 10.820 7.810 11.090 8.080 ;
        RECT 19.790 7.810 20.060 8.080 ;
        RECT 23.450 7.960 23.620 8.130 ;
        RECT 28.620 8.160 28.790 8.330 ;
        RECT 2.660 7.280 2.830 7.450 ;
        RECT 29.930 8.150 30.110 8.340 ;
        RECT 8.500 6.700 8.670 6.870 ;
        RECT 22.210 6.700 22.380 6.870 ;
        RECT 0.770 5.350 0.950 5.540 ;
        RECT 3.130 6.390 3.300 6.560 ;
        RECT 2.670 6.210 2.840 6.380 ;
        RECT 1.840 5.900 2.010 6.070 ;
        RECT 10.820 6.080 11.090 6.350 ;
        RECT 19.790 6.080 20.060 6.350 ;
        RECT 28.230 5.780 28.400 5.950 ;
        RECT 5.370 5.460 5.540 5.630 ;
        RECT 5.370 5.010 5.540 5.180 ;
        RECT 23.450 5.460 23.620 5.630 ;
        RECT 23.450 5.010 23.620 5.180 ;
        RECT 3.120 4.810 3.290 4.980 ;
        RECT 0.420 4.530 0.590 4.700 ;
        RECT 28.620 5.400 28.790 5.570 ;
        RECT 29.200 5.500 29.370 5.670 ;
        RECT 28.380 4.950 28.550 5.120 ;
        RECT 2.230 4.230 2.410 4.400 ;
        RECT 2.690 4.300 2.860 4.470 ;
        RECT 27.260 4.430 27.430 4.600 ;
        RECT 29.930 5.350 30.110 5.540 ;
        RECT 31.450 5.550 31.620 5.720 ;
        RECT 29.150 4.850 29.320 5.020 ;
        RECT 30.180 5.180 30.350 5.350 ;
        RECT 30.290 4.530 30.460 4.700 ;
        RECT 29.150 4.030 29.320 4.200 ;
        RECT 30.840 4.240 31.010 4.410 ;
        RECT 30.180 3.700 30.350 3.870 ;
        RECT 29.200 3.380 29.370 3.550 ;
        RECT 27.990 3.150 28.160 3.320 ;
        RECT 31.500 3.330 31.670 3.500 ;
        RECT 28.420 2.350 28.590 2.520 ;
        RECT 29.200 2.540 29.370 2.710 ;
        RECT 31.490 2.610 31.660 2.780 ;
        RECT 30.180 2.220 30.350 2.390 ;
        RECT 29.150 1.890 29.320 2.060 ;
        RECT 30.840 1.650 31.010 1.820 ;
        RECT 29.150 1.070 29.320 1.240 ;
        RECT 30.180 0.740 30.350 0.910 ;
        RECT 29.200 0.420 29.370 0.590 ;
        RECT 31.410 0.360 31.580 0.530 ;
      LAYER met1 ;
        RECT 0.360 9.220 0.520 9.870 ;
        RECT 0.360 8.670 0.630 9.220 ;
        RECT 0.350 8.620 0.630 8.670 ;
        RECT 0.350 8.530 0.520 8.620 ;
        RECT 0.360 5.160 0.520 8.530 ;
        RECT 0.770 8.410 0.960 9.870 ;
        RECT 2.640 9.500 2.850 9.870 ;
        RECT 2.170 9.050 2.480 9.490 ;
        RECT 2.630 9.210 2.860 9.500 ;
        RECT 0.740 8.380 0.960 8.410 ;
        RECT 0.730 8.110 0.980 8.380 ;
        RECT 0.730 8.100 0.970 8.110 ;
        RECT 0.740 7.860 0.970 8.100 ;
        RECT 0.770 5.830 0.930 7.860 ;
        RECT 1.770 7.520 2.090 7.840 ;
        RECT 2.640 7.510 2.850 9.210 ;
        RECT 3.110 8.940 3.300 9.870 ;
        RECT 3.100 8.650 3.330 8.940 ;
        RECT 1.120 7.010 1.360 7.430 ;
        RECT 2.630 7.220 2.860 7.510 ;
        RECT 2.640 7.080 2.850 7.220 ;
        RECT 1.090 6.690 1.360 7.010 ;
        RECT 1.120 6.260 1.360 6.690 ;
        RECT 3.110 6.620 3.300 8.650 ;
        RECT 3.520 7.150 3.730 9.870 ;
        RECT 5.320 7.870 5.580 8.660 ;
        RECT 3.490 6.640 3.730 7.150 ;
        RECT 2.660 6.440 2.850 6.570 ;
        RECT 2.640 6.150 2.870 6.440 ;
        RECT 3.100 6.330 3.330 6.620 ;
        RECT 1.760 5.830 2.080 6.150 ;
        RECT 0.740 5.590 0.970 5.830 ;
        RECT 0.730 5.580 0.970 5.590 ;
        RECT 0.730 5.310 0.980 5.580 ;
        RECT 0.740 5.280 0.960 5.310 ;
        RECT 0.350 5.070 0.520 5.160 ;
        RECT 0.350 5.020 0.630 5.070 ;
        RECT 0.360 4.470 0.630 5.020 ;
        RECT 0.360 3.820 0.520 4.470 ;
        RECT 0.770 3.820 0.960 5.280 ;
        RECT 2.170 4.200 2.480 4.640 ;
        RECT 2.660 4.530 2.850 6.150 ;
        RECT 3.110 5.040 3.300 6.330 ;
        RECT 3.090 4.750 3.320 5.040 ;
        RECT 2.660 4.320 2.890 4.530 ;
        RECT 2.650 4.240 2.890 4.320 ;
        RECT 2.650 3.820 2.880 4.240 ;
        RECT 3.110 3.820 3.300 4.750 ;
        RECT 3.520 3.820 3.730 6.640 ;
        RECT 4.310 6.030 4.470 6.050 ;
        RECT 4.150 5.730 4.470 6.030 ;
        RECT 5.320 4.930 5.580 5.720 ;
        RECT 10.760 3.820 11.180 9.870 ;
        RECT 19.700 3.820 20.120 9.870 ;
        RECT 22.180 3.820 22.410 9.870 ;
        RECT 23.400 8.660 23.630 9.870 ;
        RECT 28.400 9.050 28.710 9.490 ;
        RECT 23.400 7.870 23.660 8.660 ;
        RECT 28.550 8.090 28.870 8.410 ;
        RECT 23.400 5.720 23.630 7.870 ;
        RECT 29.520 7.300 29.760 7.430 ;
        RECT 29.520 6.980 29.780 7.300 ;
        RECT 23.400 4.930 23.660 5.720 ;
        RECT 28.550 5.330 28.870 5.650 ;
        RECT 31.380 5.480 31.700 5.800 ;
        RECT 23.400 3.820 23.630 4.930 ;
        RECT 28.300 4.880 28.620 5.200 ;
        RECT 27.190 4.350 27.510 4.670 ;
        RECT 27.920 3.070 28.240 3.390 ;
        RECT 29.130 3.300 29.450 3.620 ;
        RECT 31.430 3.260 31.750 3.580 ;
        RECT 29.130 2.470 29.450 2.790 ;
        RECT 31.420 2.540 31.740 2.860 ;
        RECT 29.080 1.820 29.400 2.140 ;
        RECT 29.080 0.990 29.400 1.310 ;
        RECT 12.370 0.050 12.690 0.350 ;
        RECT 18.170 0.050 18.490 0.350 ;
        RECT 29.130 0.340 29.450 0.660 ;
        RECT 31.340 0.290 31.660 0.610 ;
      LAYER via ;
        RECT 2.190 9.080 2.450 9.340 ;
        RECT 1.800 7.550 2.060 7.810 ;
        RECT 1.090 6.720 1.350 6.980 ;
        RECT 1.790 5.860 2.050 6.120 ;
        RECT 2.190 4.350 2.450 4.610 ;
        RECT 4.180 5.750 4.440 6.010 ;
        RECT 28.430 9.080 28.690 9.340 ;
        RECT 28.580 8.120 28.840 8.380 ;
        RECT 29.520 7.010 29.780 7.270 ;
        RECT 28.580 5.360 28.840 5.620 ;
        RECT 31.410 5.510 31.670 5.770 ;
        RECT 28.330 4.910 28.590 5.170 ;
        RECT 27.220 4.380 27.480 4.640 ;
        RECT 27.950 3.100 28.210 3.360 ;
        RECT 29.160 3.330 29.420 3.590 ;
        RECT 31.460 3.290 31.720 3.550 ;
        RECT 29.160 2.500 29.420 2.760 ;
        RECT 31.450 2.570 31.710 2.830 ;
        RECT 29.110 1.850 29.370 2.110 ;
        RECT 29.110 1.020 29.370 1.280 ;
        RECT 29.160 0.370 29.420 0.630 ;
        RECT 12.400 0.070 12.660 0.330 ;
        RECT 18.200 0.070 18.460 0.330 ;
        RECT 31.370 0.320 31.630 0.580 ;
      LAYER met2 ;
        RECT 2.410 9.380 2.730 9.390 ;
        RECT 2.170 9.370 2.730 9.380 ;
        RECT 28.400 9.370 28.710 9.380 ;
        RECT 0.000 9.190 11.520 9.370 ;
        RECT 19.350 9.190 30.880 9.370 ;
        RECT 2.170 9.050 2.480 9.190 ;
        RECT 28.400 9.050 28.710 9.190 ;
        RECT 28.550 8.350 28.860 8.420 ;
        RECT 28.550 8.130 30.880 8.350 ;
        RECT 28.550 8.090 28.860 8.130 ;
        RECT 1.780 7.830 2.090 7.850 ;
        RECT 1.780 7.640 11.520 7.830 ;
        RECT 1.780 7.520 2.090 7.640 ;
        RECT 1.060 6.950 1.380 6.980 ;
        RECT 1.060 6.720 11.520 6.950 ;
        RECT 2.170 4.500 2.480 4.640 ;
        RECT 0.000 4.490 2.480 4.500 ;
        RECT 0.000 4.340 11.520 4.490 ;
        RECT 0.000 4.320 2.480 4.340 ;
        RECT 2.170 4.310 2.480 4.320 ;
        RECT 15.460 3.820 23.450 4.020 ;
        RECT 22.050 3.140 22.270 3.150 ;
        RECT 15.470 2.890 22.300 3.140 ;
        RECT 23.230 3.100 23.450 3.820 ;
        RECT 15.470 1.970 18.980 2.160 ;
        RECT 18.750 1.370 18.980 1.970 ;
        RECT 22.010 1.720 22.300 2.890 ;
        RECT 23.200 3.060 23.450 3.100 ;
        RECT 23.200 2.420 23.460 3.060 ;
        RECT 23.200 2.210 27.330 2.420 ;
        RECT 27.120 2.070 27.330 2.210 ;
        RECT 29.080 2.070 29.390 2.150 ;
        RECT 27.120 1.860 29.390 2.070 ;
        RECT 29.080 1.820 29.390 1.860 ;
        RECT 22.010 1.500 24.900 1.720 ;
        RECT 22.010 1.490 22.300 1.500 ;
        RECT 18.750 1.220 18.970 1.370 ;
        RECT 29.080 1.270 29.390 1.310 ;
        RECT 23.120 1.220 29.390 1.270 ;
        RECT 18.750 1.060 29.390 1.220 ;
        RECT 18.750 1.000 23.510 1.060 ;
        RECT 29.080 0.980 29.390 1.060 ;
        RECT 29.130 0.580 29.440 0.660 ;
        RECT 31.340 0.580 31.650 0.620 ;
        RECT 29.130 0.350 31.840 0.580 ;
        RECT 29.130 0.330 29.440 0.350 ;
        RECT 31.340 0.290 31.650 0.350 ;
  END
END sky130_hilas_TA2Cell_1FG_Strong

MACRO sky130_hilas_TA2Cell_NoFG
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TA2Cell_NoFG ;
  ORIGIN 14.730 -1.400 ;
  SIZE 17.920 BY 9.870 ;
  PIN COLSEL1
    PORT
      LAYER met1 ;
        RECT -4.160 7.370 -3.970 7.450 ;
    END
  END COLSEL1
  PIN VIN12
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -2.260 1.670 -1.950 1.740 ;
        RECT -2.860 1.420 -1.950 1.670 ;
        RECT -2.260 1.410 -1.950 1.420 ;
    END
  END VIN12
  PIN VIN21
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -0.940 4.750 -0.630 4.790 ;
        RECT -1.030 4.740 -0.600 4.750 ;
        RECT -1.260 4.510 -0.160 4.740 ;
        RECT -0.940 4.460 -0.630 4.510 ;
    END
  END VIN21
  PIN VIN22
    ANTENNAGATEAREA 4.299400 ;
    ANTENNADIFFAREA 6.715500 ;
    PORT
      LAYER nwell ;
        RECT -2.550 7.450 0.760 11.270 ;
        RECT -3.510 5.230 0.760 7.450 ;
        RECT -3.510 1.410 -0.090 5.230 ;
        RECT -1.950 1.400 -0.090 1.410 ;
      LAYER met2 ;
        RECT -0.630 8.410 -0.310 8.670 ;
        RECT -0.590 8.390 0.590 8.410 ;
        RECT -0.590 8.130 0.630 8.390 ;
        RECT -0.590 8.070 0.590 8.130 ;
        RECT -0.630 8.060 0.590 8.070 ;
        RECT -0.630 7.810 -0.310 8.060 ;
        RECT -1.300 7.430 -1.050 7.440 ;
        RECT -0.700 7.430 -0.390 7.440 ;
        RECT -1.300 7.180 -0.390 7.430 ;
        RECT -0.700 7.110 -0.390 7.180 ;
        RECT 0.270 7.110 0.580 7.160 ;
        RECT 2.520 7.110 2.830 7.210 ;
        RECT -1.570 6.990 -1.260 7.060 ;
        RECT 0.270 6.990 2.830 7.110 ;
        RECT -1.570 6.880 2.830 6.990 ;
        RECT -1.570 6.780 0.760 6.880 ;
        RECT -1.570 6.730 -1.260 6.780 ;
        RECT -0.550 6.570 -0.240 6.610 ;
        RECT -0.730 6.430 0.010 6.570 ;
        RECT 0.220 6.430 0.530 6.510 ;
        RECT -0.730 6.320 0.530 6.430 ;
        RECT -0.550 6.280 0.530 6.320 ;
        RECT -0.240 6.220 0.530 6.280 ;
        RECT -0.240 6.200 0.010 6.220 ;
        RECT 0.220 6.180 0.530 6.220 ;
        RECT -1.670 6.040 -1.360 6.070 ;
        RECT -1.720 5.930 -1.360 6.040 ;
        RECT 1.230 6.000 1.570 6.090 ;
        RECT -3.280 5.900 -1.360 5.930 ;
        RECT -1.120 5.900 1.570 6.000 ;
        RECT -3.280 5.890 1.570 5.900 ;
        RECT -10.770 5.810 1.570 5.890 ;
        RECT -10.770 5.740 0.760 5.810 ;
        RECT 1.230 5.760 1.570 5.810 ;
        RECT -3.280 5.720 0.760 5.740 ;
        RECT -3.280 5.710 -1.410 5.720 ;
        RECT -1.120 5.240 -0.930 5.720 ;
        RECT -0.210 5.630 0.000 5.640 ;
        RECT 0.220 5.630 0.530 5.670 ;
        RECT -0.210 5.560 0.530 5.630 ;
        RECT -0.500 5.540 0.530 5.560 ;
        RECT -0.550 5.420 0.530 5.540 ;
        RECT -0.550 5.350 0.000 5.420 ;
        RECT -0.550 5.290 -0.080 5.350 ;
        RECT 0.220 5.340 0.530 5.420 ;
        RECT -11.910 5.050 -0.930 5.240 ;
        RECT -11.910 4.870 -11.720 5.050 ;
        RECT -11.930 3.880 -11.580 4.870 ;
        RECT -2.500 4.340 -2.190 4.390 ;
        RECT -2.820 4.110 -1.720 4.340 ;
        RECT -2.820 4.100 -2.160 4.110 ;
        RECT -2.500 4.060 -2.190 4.100 ;
    END
  END VIN22
  PIN OUTPUT1
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER met2 ;
        RECT 0.270 4.140 0.580 4.200 ;
        RECT 2.560 4.140 2.870 4.270 ;
        RECT 0.270 3.920 3.190 4.140 ;
        RECT 0.270 3.870 0.580 3.920 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER met2 ;
        RECT 0.270 4.970 0.580 5.020 ;
        RECT 2.570 4.970 2.880 4.990 ;
        RECT 0.270 4.740 3.190 4.970 ;
        RECT 0.270 4.690 0.580 4.740 ;
        RECT 2.570 4.660 2.880 4.740 ;
    END
  END OUTPUT2
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 1.230 1.400 1.570 7.450 ;
      LAYER via ;
        RECT 1.270 5.790 1.530 6.050 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 1.920 7.270 3.190 7.450 ;
        RECT 1.910 1.400 3.190 7.270 ;
      LAYER met1 ;
        RECT 1.900 5.870 2.170 7.450 ;
        RECT 1.900 5.580 2.180 5.870 ;
        RECT 1.900 3.280 2.170 5.580 ;
        RECT 1.900 2.990 2.180 3.280 ;
        RECT 1.900 1.400 2.170 2.990 ;
    END
  END VPWR
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT -14.730 6.770 -14.660 6.950 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT -14.730 1.920 -14.650 2.070 ;
    END
  END DRAIN2
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT -14.380 7.380 -13.960 7.450 ;
    END
  END VTUN
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT -10.680 7.370 -10.450 7.450 ;
    END
  END GATE1
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT -3.720 7.370 -3.440 7.450 ;
    END
  END VINJ
  OBS
      LAYER nwell ;
        RECT -10.760 10.520 -9.030 11.270 ;
        RECT -10.760 6.950 -9.020 10.520 ;
        RECT -7.000 8.880 -4.280 10.530 ;
        RECT -7.000 8.840 -4.290 8.880 ;
        RECT -7.000 7.510 -4.290 7.550 ;
        RECT -10.760 5.230 -9.030 6.950 ;
        RECT -7.000 5.860 -4.280 7.510 ;
      LAYER li1 ;
        RECT -1.650 10.690 -1.120 10.860 ;
        RECT 0.160 10.590 0.360 10.940 ;
        RECT 0.160 10.560 0.370 10.590 ;
        RECT -3.520 10.110 -3.170 10.280 ;
        RECT -2.150 10.110 -1.820 10.280 ;
        RECT -10.330 9.130 -9.780 9.560 ;
        RECT -6.700 9.320 -6.470 10.010 ;
        RECT -1.400 9.780 -1.230 10.300 ;
        RECT -1.560 9.520 -1.230 9.780 ;
        RECT -3.520 9.320 -3.170 9.490 ;
        RECT -2.150 9.320 -1.820 9.490 ;
        RECT -7.730 8.300 -7.540 8.700 ;
        RECT -3.510 8.530 -3.170 8.700 ;
        RECT -2.150 8.530 -1.820 8.700 ;
        RECT -1.400 8.610 -1.230 9.520 ;
        RECT -0.570 8.700 -0.400 10.310 ;
        RECT 0.150 9.980 0.370 10.560 ;
        RECT 0.160 9.970 0.370 9.980 ;
        RECT -0.200 9.800 -0.010 9.810 ;
        RECT -0.200 9.510 0.000 9.800 ;
        RECT -0.210 9.180 0.030 9.510 ;
        RECT -7.920 8.290 -7.540 8.300 ;
        RECT -7.920 8.110 -4.180 8.290 ;
        RECT -7.920 8.070 -7.540 8.110 ;
        RECT -10.330 7.400 -9.780 7.830 ;
        RECT -7.730 7.690 -7.540 8.070 ;
        RECT -2.070 7.960 -1.900 8.530 ;
        RECT -0.570 8.510 -0.390 8.700 ;
        RECT -3.510 7.790 -3.170 7.960 ;
        RECT -2.150 7.790 -1.820 7.960 ;
        RECT -6.700 6.380 -6.470 7.110 ;
        RECT -3.520 7.000 -3.170 7.170 ;
        RECT -2.150 7.000 -1.820 7.170 ;
        RECT -1.400 7.020 -1.230 7.880 ;
        RECT -0.570 7.790 -0.390 7.980 ;
        RECT -0.960 7.400 -0.790 7.450 ;
        RECT -0.570 7.400 -0.400 7.790 ;
        RECT -0.960 7.140 -0.400 7.400 ;
        RECT -0.960 7.120 -0.790 7.140 ;
        RECT -3.520 6.210 -3.170 6.380 ;
        RECT -11.900 3.870 -11.440 4.880 ;
        RECT -3.100 3.070 -2.920 6.980 ;
        RECT -2.290 6.380 -2.120 6.970 ;
        RECT -1.560 6.760 -1.230 7.020 ;
        RECT -0.570 6.880 -0.400 7.140 ;
        RECT -0.210 6.980 0.030 7.310 ;
        RECT 0.510 7.120 0.710 7.160 ;
        RECT -2.290 6.210 -1.820 6.380 ;
        RECT -2.290 5.190 -2.120 6.210 ;
        RECT -1.540 6.190 -1.230 6.760 ;
        RECT -0.810 6.710 -0.400 6.880 ;
        RECT -0.730 6.570 -0.400 6.710 ;
        RECT -0.200 6.690 0.000 6.980 ;
        RECT 0.280 6.860 0.710 7.120 ;
        RECT 0.510 6.830 0.710 6.860 ;
        RECT -0.200 6.680 -0.010 6.690 ;
        RECT -0.730 6.310 -0.250 6.570 ;
        RECT 0.160 6.510 0.370 6.520 ;
        RECT 0.100 6.470 0.370 6.510 ;
        RECT 0.510 6.470 0.710 6.500 ;
        RECT -1.540 6.040 -1.360 6.190 ;
        RECT -0.730 6.180 -0.400 6.310 ;
        RECT 0.100 6.210 0.710 6.470 ;
        RECT 0.100 6.180 0.370 6.210 ;
        RECT -1.660 6.010 -1.340 6.040 ;
        RECT -1.660 5.820 -1.330 6.010 ;
        RECT -1.660 5.800 -1.340 5.820 ;
        RECT -1.660 5.780 -1.120 5.800 ;
        RECT -1.650 5.630 -1.120 5.780 ;
        RECT -2.370 5.130 -1.830 5.190 ;
        RECT -2.370 5.020 -1.820 5.130 ;
        RECT -2.010 4.900 -1.820 5.020 ;
        RECT -2.540 4.600 -2.370 4.760 ;
        RECT -2.540 4.430 -2.320 4.600 ;
        RECT -2.490 4.350 -2.320 4.430 ;
        RECT -2.490 4.310 -2.170 4.350 ;
        RECT -2.490 4.120 -2.160 4.310 ;
        RECT -2.490 4.090 -2.170 4.120 ;
        RECT -3.220 3.030 -2.900 3.070 ;
        RECT -3.220 2.840 -2.890 3.030 ;
        RECT -3.220 2.810 -2.900 2.840 ;
        RECT -3.100 1.880 -2.920 2.810 ;
        RECT -2.290 2.540 -2.120 3.920 ;
        RECT -2.290 2.280 -1.810 2.540 ;
        RECT -2.290 2.140 -2.040 2.280 ;
        RECT -2.370 1.970 -2.040 2.140 ;
        RECT -1.540 1.870 -1.360 5.630 ;
        RECT -0.730 4.930 -0.560 6.180 ;
        RECT 0.150 5.930 0.370 6.180 ;
        RECT 0.510 6.170 0.710 6.210 ;
        RECT 1.100 6.170 1.650 7.160 ;
        RECT 2.470 7.040 3.050 7.210 ;
        RECT 2.470 6.940 2.860 7.040 ;
        RECT 2.470 6.910 2.850 6.940 ;
        RECT 2.470 6.760 2.830 6.910 ;
        RECT 2.120 6.590 2.830 6.760 ;
        RECT 0.160 5.900 0.370 5.930 ;
        RECT 0.160 5.670 0.360 5.900 ;
        RECT 2.120 5.840 2.820 6.150 ;
        RECT 0.100 5.640 0.360 5.670 ;
        RECT 0.510 5.640 0.710 5.680 ;
        RECT 0.100 5.380 0.710 5.640 ;
        RECT 0.100 5.340 0.270 5.380 ;
        RECT 0.510 5.350 0.710 5.380 ;
        RECT 0.510 4.990 0.710 5.020 ;
        RECT -0.930 4.730 -0.610 4.760 ;
        RECT 0.280 4.730 0.710 4.990 ;
        RECT -0.930 4.540 -0.600 4.730 ;
        RECT 0.510 4.690 0.710 4.730 ;
        RECT 1.100 4.690 1.650 5.680 ;
        RECT 1.970 5.610 2.820 5.840 ;
        RECT 2.120 5.270 2.820 5.610 ;
        RECT 2.580 4.910 2.900 4.950 ;
        RECT 2.580 4.850 2.910 4.910 ;
        RECT 2.110 4.720 2.910 4.850 ;
        RECT 2.110 4.690 2.900 4.720 ;
        RECT 2.110 4.670 2.810 4.690 ;
        RECT -0.930 4.500 -0.610 4.540 ;
        RECT -0.930 4.420 -0.760 4.500 ;
        RECT -0.980 4.250 -0.760 4.420 ;
        RECT -0.980 4.090 -0.810 4.250 ;
        RECT 0.510 4.160 0.710 4.200 ;
        RECT -0.450 3.830 -0.260 3.950 ;
        RECT 0.280 3.900 0.710 4.160 ;
        RECT 0.510 3.870 0.710 3.900 ;
        RECT -0.810 3.720 -0.260 3.830 ;
        RECT -0.810 3.660 -0.270 3.720 ;
        RECT -0.730 1.880 -0.560 3.660 ;
        RECT 0.100 3.510 0.270 3.550 ;
        RECT 0.510 3.510 0.710 3.540 ;
        RECT 0.100 3.250 0.710 3.510 ;
        RECT 0.100 3.220 0.270 3.250 ;
        RECT 0.510 3.210 0.710 3.250 ;
        RECT 1.100 3.210 1.650 4.200 ;
        RECT 2.570 4.190 2.890 4.230 ;
        RECT 2.110 4.010 2.900 4.190 ;
        RECT 2.570 4.000 2.900 4.010 ;
        RECT 2.570 3.970 2.890 4.000 ;
        RECT 2.120 3.250 2.820 3.590 ;
        RECT 1.970 3.020 2.820 3.250 ;
        RECT 0.100 2.680 0.270 2.710 ;
        RECT 0.510 2.680 0.710 2.720 ;
        RECT 0.100 2.420 0.710 2.680 ;
        RECT 0.100 2.380 0.270 2.420 ;
        RECT 0.510 2.390 0.710 2.420 ;
        RECT 0.510 2.030 0.710 2.060 ;
        RECT 0.280 1.770 0.710 2.030 ;
        RECT 0.510 1.730 0.710 1.770 ;
        RECT 1.100 1.730 1.650 2.720 ;
        RECT 2.120 2.710 2.820 3.020 ;
        RECT 2.120 2.100 2.830 2.270 ;
        RECT 2.470 1.820 2.830 2.100 ;
        RECT -2.520 1.710 -2.350 1.730 ;
        RECT -2.520 1.450 -1.960 1.710 ;
        RECT 2.470 1.650 3.050 1.820 ;
        RECT -2.520 1.400 -2.350 1.450 ;
      LAYER mcon ;
        RECT 0.170 10.390 0.340 10.560 ;
        RECT -6.670 9.810 -6.500 9.980 ;
        RECT -10.330 9.210 -10.060 9.480 ;
        RECT -6.670 9.360 -6.500 9.530 ;
        RECT -1.500 9.560 -1.330 9.730 ;
        RECT -0.190 9.550 -0.010 9.740 ;
        RECT -7.910 8.100 -7.740 8.270 ;
        RECT -10.330 7.480 -10.060 7.750 ;
        RECT -6.670 6.860 -6.500 7.030 ;
        RECT -0.630 7.180 -0.460 7.350 ;
        RECT -6.670 6.410 -6.500 6.580 ;
        RECT -11.870 4.620 -11.700 4.790 ;
        RECT -11.870 3.930 -11.700 4.100 ;
        RECT -1.500 6.800 -1.330 6.970 ;
        RECT -0.190 6.750 -0.010 6.940 ;
        RECT 0.340 6.900 0.510 7.070 ;
        RECT 2.590 6.950 2.760 7.120 ;
        RECT 1.320 6.580 1.490 6.750 ;
        RECT -0.480 6.350 -0.310 6.520 ;
        RECT 0.290 6.250 0.460 6.420 ;
        RECT -1.600 5.830 -1.430 6.000 ;
        RECT -2.000 4.930 -1.830 5.100 ;
        RECT -2.430 4.130 -2.260 4.300 ;
        RECT -3.160 2.850 -2.990 3.020 ;
        RECT -2.040 2.330 -1.870 2.500 ;
        RECT 0.170 5.930 0.340 6.100 ;
        RECT 0.290 5.430 0.460 5.600 ;
        RECT 1.980 5.640 2.150 5.810 ;
        RECT 1.320 5.100 1.490 5.270 ;
        RECT 0.340 4.780 0.510 4.950 ;
        RECT -0.870 4.550 -0.700 4.720 ;
        RECT 2.640 4.730 2.810 4.900 ;
        RECT -0.440 3.750 -0.270 3.920 ;
        RECT 0.340 3.940 0.510 4.110 ;
        RECT 2.630 4.010 2.800 4.180 ;
        RECT 1.320 3.620 1.490 3.790 ;
        RECT 0.290 3.290 0.460 3.460 ;
        RECT 1.980 3.050 2.150 3.220 ;
        RECT 0.290 2.470 0.460 2.640 ;
        RECT 1.320 2.140 1.490 2.310 ;
        RECT 0.340 1.820 0.510 1.990 ;
        RECT 2.550 1.760 2.720 1.930 ;
        RECT -2.190 1.500 -2.020 1.670 ;
      LAYER met1 ;
        RECT -10.420 5.220 -10.000 11.270 ;
        RECT -7.940 5.220 -7.710 11.270 ;
        RECT -6.720 10.060 -6.490 11.270 ;
        RECT -1.720 10.450 -1.410 10.890 ;
        RECT -6.720 9.270 -6.460 10.060 ;
        RECT -0.200 9.810 -0.010 11.270 ;
        RECT 0.240 10.620 0.520 11.270 ;
        RECT 0.130 10.020 0.520 10.620 ;
        RECT -1.570 9.490 -1.250 9.810 ;
        RECT -0.200 9.780 0.020 9.810 ;
        RECT -0.220 9.510 0.030 9.780 ;
        RECT -0.210 9.500 0.030 9.510 ;
        RECT -6.720 7.120 -6.490 9.270 ;
        RECT -0.210 9.260 0.020 9.500 ;
        RECT -0.600 8.700 -0.360 8.830 ;
        RECT -0.600 8.380 -0.340 8.700 ;
        RECT -0.600 7.780 -0.340 8.100 ;
        RECT -0.600 7.660 -0.360 7.780 ;
        RECT -6.720 6.330 -6.460 7.120 ;
        RECT -0.710 7.110 -0.390 7.430 ;
        RECT -0.170 7.230 -0.010 9.260 ;
        RECT 0.240 8.420 0.520 10.020 ;
        RECT 0.240 8.100 0.600 8.420 ;
        RECT -1.570 6.730 -1.250 7.050 ;
        RECT -0.210 6.990 0.020 7.230 ;
        RECT 0.240 7.150 0.520 8.100 ;
        RECT -0.210 6.980 0.030 6.990 ;
        RECT -0.220 6.710 0.030 6.980 ;
        RECT 0.240 6.830 0.590 7.150 ;
        RECT 2.520 6.880 2.840 7.200 ;
        RECT -0.200 6.680 0.020 6.710 ;
        RECT -6.720 5.220 -6.490 6.330 ;
        RECT -0.560 6.280 -0.240 6.600 ;
        RECT -1.670 6.040 -1.350 6.070 ;
        RECT -1.720 5.750 -1.350 6.040 ;
        RECT -1.720 5.600 -1.410 5.750 ;
        RECT -0.450 5.590 -0.240 5.700 ;
        RECT -0.470 5.270 -0.210 5.590 ;
        RECT -11.940 3.870 -11.560 4.880 ;
        RECT -2.030 4.870 -1.800 5.160 ;
        RECT -2.500 4.060 -2.180 4.380 ;
        RECT -2.010 3.580 -1.800 4.870 ;
        RECT -0.940 4.470 -0.620 4.790 ;
        RECT -0.450 3.980 -0.240 5.270 ;
        RECT -0.200 5.220 -0.010 6.680 ;
        RECT 0.240 6.500 0.520 6.830 ;
        RECT 0.220 6.470 0.540 6.500 ;
        RECT 0.130 6.180 0.540 6.470 ;
        RECT 0.130 5.870 0.520 6.180 ;
        RECT 0.240 5.670 0.520 5.870 ;
        RECT 0.220 5.350 0.540 5.670 ;
        RECT 0.240 5.220 0.520 5.350 ;
        RECT 0.270 4.700 0.590 5.020 ;
        RECT 2.570 4.660 2.890 4.980 ;
        RECT -0.470 3.690 -0.240 3.980 ;
        RECT 0.270 3.870 0.590 4.190 ;
        RECT 2.560 3.940 2.880 4.260 ;
        RECT -2.030 3.260 -1.770 3.580 ;
        RECT -2.010 3.150 -1.800 3.260 ;
        RECT 0.220 3.220 0.540 3.540 ;
        RECT -3.230 2.780 -2.910 3.100 ;
        RECT -2.120 2.250 -1.800 2.570 ;
        RECT 0.220 2.390 0.540 2.710 ;
        RECT 0.270 1.740 0.590 2.060 ;
        RECT -2.270 1.420 -1.950 1.740 ;
        RECT 2.480 1.690 2.800 2.010 ;
      LAYER via ;
        RECT -1.690 10.480 -1.430 10.740 ;
        RECT -1.540 9.520 -1.280 9.780 ;
        RECT -0.600 8.410 -0.340 8.670 ;
        RECT -0.600 7.810 -0.340 8.070 ;
        RECT -0.680 7.140 -0.420 7.400 ;
        RECT 0.340 8.130 0.600 8.390 ;
        RECT -1.540 6.760 -1.280 7.020 ;
        RECT 0.300 6.860 0.560 7.120 ;
        RECT 2.550 6.910 2.810 7.170 ;
        RECT -0.530 6.310 -0.270 6.570 ;
        RECT -1.640 6.010 -1.380 6.040 ;
        RECT -1.690 5.780 -1.380 6.010 ;
        RECT -1.690 5.750 -1.430 5.780 ;
        RECT -0.470 5.300 -0.210 5.560 ;
        RECT -11.900 3.910 -11.610 4.840 ;
        RECT -2.470 4.090 -2.210 4.350 ;
        RECT -0.910 4.500 -0.650 4.760 ;
        RECT 0.250 6.210 0.510 6.470 ;
        RECT 0.250 5.380 0.510 5.640 ;
        RECT 0.300 4.730 0.560 4.990 ;
        RECT 2.600 4.690 2.860 4.950 ;
        RECT 0.300 3.900 0.560 4.160 ;
        RECT 2.590 3.970 2.850 4.230 ;
        RECT -2.030 3.290 -1.770 3.550 ;
        RECT 0.250 3.250 0.510 3.510 ;
        RECT -3.200 2.810 -2.940 3.070 ;
        RECT -2.090 2.280 -1.830 2.540 ;
        RECT 0.250 2.420 0.510 2.680 ;
        RECT 0.300 1.770 0.560 2.030 ;
        RECT -2.240 1.450 -1.980 1.710 ;
        RECT 2.510 1.720 2.770 1.980 ;
      LAYER met2 ;
        RECT -1.720 10.770 -1.410 10.780 ;
        RECT -10.770 10.590 0.760 10.770 ;
        RECT -1.720 10.450 -1.410 10.590 ;
        RECT -1.570 9.750 -1.260 9.820 ;
        RECT -1.570 9.530 0.760 9.750 ;
        RECT -1.570 9.490 -1.260 9.530 ;
        RECT -2.110 3.470 -1.640 3.560 ;
        RECT 0.220 3.470 0.530 3.550 ;
        RECT -2.110 3.310 0.530 3.470 ;
        RECT -2.060 3.290 0.530 3.310 ;
        RECT -1.770 3.270 0.530 3.290 ;
        RECT -0.080 3.260 0.530 3.270 ;
        RECT 0.220 3.220 0.530 3.260 ;
        RECT -3.340 3.110 -3.180 3.180 ;
        RECT -3.340 2.780 -2.920 3.110 ;
        RECT 0.220 2.670 0.530 2.710 ;
        RECT -2.060 2.570 0.530 2.670 ;
        RECT -2.110 2.530 0.530 2.570 ;
        RECT -2.290 2.460 0.530 2.530 ;
        RECT -2.290 2.280 -1.740 2.460 ;
        RECT 0.220 2.380 0.530 2.460 ;
        RECT -2.110 2.240 -1.800 2.280 ;
        RECT 0.270 1.980 0.580 2.060 ;
        RECT 2.480 1.980 2.790 2.020 ;
        RECT 0.270 1.750 2.980 1.980 ;
        RECT 0.270 1.730 0.580 1.750 ;
        RECT 2.480 1.690 2.790 1.750 ;
  END
END sky130_hilas_TA2Cell_NoFG

MACRO sky130_hilas_TopLevelTextStructure
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TopLevelTextStructure ;
  ORIGIN -2.180 10.310 ;
  SIZE 130.250 BY 78.160 ;
  PIN DIG24 
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 67.710 22.600 67.750 22.690 ;
        RECT 67.600 22.510 68.810 22.600 ;
        RECT 67.600 22.450 68.940 22.510 ;
        RECT 75.910 22.450 76.230 22.500 ;
        RECT 67.600 22.400 76.230 22.450 ;
        RECT 68.630 22.290 76.230 22.400 ;
        RECT 68.630 22.180 68.940 22.290 ;
        RECT 75.910 22.240 76.230 22.290 ;
        RECT 75.890 13.290 131.720 13.330 ;
        RECT 75.890 12.830 132.430 13.290 ;
        RECT 130.420 -7.170 132.430 12.830 ;
        RECT 130.390 -7.750 132.430 -7.170 ;
        RECT 130.390 -7.820 132.420 -7.750 ;
    END
  END DIG24 
  PIN DIG23
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 67.700 21.630 68.910 21.740 ;
        RECT 67.700 21.540 68.940 21.630 ;
        RECT 68.630 21.520 68.940 21.540 ;
        RECT 75.390 21.520 75.710 21.570 ;
        RECT 68.630 21.360 75.710 21.520 ;
        RECT 68.630 21.300 68.940 21.360 ;
        RECT 75.390 21.310 75.710 21.360 ;
        RECT 126.330 12.430 128.340 12.450 ;
        RECT 75.350 11.930 128.340 12.430 ;
        RECT 126.330 -7.190 128.340 11.930 ;
        RECT 126.330 -7.840 128.370 -7.190 ;
        RECT 126.330 -7.920 128.340 -7.840 ;
    END
  END DIG23
  PIN DIG22
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 68.630 19.710 68.940 19.740 ;
        RECT 67.690 19.680 68.940 19.710 ;
        RECT 74.920 19.680 75.240 19.730 ;
        RECT 67.690 19.550 75.240 19.680 ;
        RECT 68.630 19.520 75.240 19.550 ;
        RECT 68.630 19.410 68.940 19.520 ;
        RECT 74.920 19.470 75.240 19.520 ;
        RECT 74.880 11.510 124.150 11.530 ;
        RECT 74.880 11.030 124.260 11.510 ;
        RECT 122.250 -7.170 124.260 11.030 ;
        RECT 122.250 -7.820 124.320 -7.170 ;
        RECT 122.250 -7.860 124.260 -7.820 ;
    END
  END DIG22
  PIN DIG21
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 68.630 18.750 68.940 18.860 ;
        RECT 74.420 18.750 74.740 18.800 ;
        RECT 68.630 18.740 74.740 18.750 ;
        RECT 67.700 18.590 74.740 18.740 ;
        RECT 67.700 18.560 68.940 18.590 ;
        RECT 68.630 18.530 68.940 18.560 ;
        RECT 74.420 18.540 74.740 18.590 ;
        RECT 74.400 10.620 120.190 10.630 ;
        RECT 74.400 10.130 120.400 10.620 ;
        RECT 118.390 -7.170 120.400 10.130 ;
        RECT 118.330 -7.690 120.400 -7.170 ;
        RECT 118.330 -7.820 120.360 -7.690 ;
    END
  END DIG21
  PIN DIG29
    PORT
      LAYER met2 ;
        RECT 110.140 -6.470 110.330 -6.300 ;
        RECT 110.140 -6.660 115.140 -6.470 ;
        RECT 114.950 -7.190 115.140 -6.660 ;
        RECT 115.790 -7.190 115.980 -7.120 ;
        RECT 114.280 -7.840 116.310 -7.190 ;
    END
  END DIG29
  PIN DIG28
    PORT
      LAYER met2 ;
        RECT 109.170 -7.260 109.380 -6.280 ;
        RECT 110.300 -7.260 112.330 -7.170 ;
        RECT 109.170 -7.470 112.330 -7.260 ;
        RECT 110.300 -7.820 112.330 -7.470 ;
    END
  END DIG28
  PIN DIG27
    PORT
      LAYER met2 ;
        RECT 107.240 -7.170 107.450 -6.280 ;
        RECT 106.120 -7.820 108.150 -7.170 ;
    END
  END DIG27
  PIN DIG26
    ANTENNAGATEAREA 49.910000 ;
    ANTENNADIFFAREA 293.818481 ;
    PORT
      LAYER nwell ;
        RECT 28.530 61.660 31.240 61.700 ;
        RECT 28.520 60.010 31.240 61.660 ;
        RECT 28.530 58.670 31.240 58.710 ;
        RECT 28.520 56.010 31.240 58.670 ;
        RECT 41.220 44.250 42.990 50.490 ;
        RECT 82.360 44.600 85.670 49.220 ;
        RECT 92.150 48.480 93.880 49.230 ;
        RECT 92.140 44.910 93.880 48.480 ;
        RECT 105.480 46.840 108.200 48.490 ;
        RECT 105.480 46.800 108.190 46.840 ;
        RECT 19.360 41.090 21.930 44.180 ;
        RECT 62.020 43.850 63.750 44.600 ;
        RECT 62.010 43.450 63.750 43.850 ;
        RECT 62.010 40.280 66.010 43.450 ;
        RECT 79.810 43.190 85.670 44.600 ;
        RECT 92.150 43.190 93.880 44.910 ;
        RECT 105.480 45.470 108.190 45.510 ;
        RECT 105.480 44.110 108.200 45.470 ;
        RECT 109.930 45.410 113.240 49.230 ;
        RECT 109.280 45.400 114.410 45.410 ;
        RECT 109.270 44.110 114.410 45.400 ;
        RECT 105.480 43.820 114.410 44.110 ;
        RECT 107.560 43.190 114.410 43.820 ;
        RECT 79.810 40.780 83.120 43.190 ;
        RECT 79.160 40.770 84.290 40.780 ;
        RECT 62.020 38.560 66.010 40.280 ;
        RECT 62.590 37.400 66.010 38.560 ;
        RECT 79.150 38.560 84.290 40.770 ;
        RECT 79.150 34.730 81.010 38.560 ;
        RECT 83.010 37.290 84.290 38.560 ;
        RECT 107.560 39.360 111.130 43.190 ;
        RECT 113.130 39.360 114.410 43.190 ;
        RECT 107.560 38.060 110.320 39.360 ;
        RECT 83.010 35.430 84.740 37.290 ;
        RECT 83.000 33.590 84.740 35.430 ;
        RECT 54.990 27.460 57.540 27.470 ;
        RECT 54.980 23.650 57.540 27.460 ;
        RECT 59.070 23.650 61.300 27.470 ;
        RECT 62.590 27.330 66.010 33.380 ;
        RECT 83.010 31.240 84.740 33.590 ;
        RECT 90.520 37.280 93.070 37.290 ;
        RECT 90.520 31.260 93.080 37.280 ;
        RECT 90.520 31.250 93.070 31.260 ;
        RECT 63.320 26.840 65.050 27.330 ;
        RECT 63.320 23.770 65.060 26.840 ;
        RECT 54.980 23.640 61.300 23.650 ;
        RECT 54.980 23.490 57.650 23.640 ;
        RECT 54.980 23.480 57.830 23.490 ;
        RECT 19.900 19.290 20.460 21.260 ;
        RECT 41.220 16.790 42.990 23.030 ;
        RECT 46.950 16.790 49.460 23.030 ;
        RECT 54.980 21.440 57.650 23.480 ;
        RECT 54.990 21.430 57.650 21.440 ;
        RECT 55.500 17.610 57.650 21.430 ;
        RECT 59.070 21.420 61.300 23.640 ;
        RECT 62.930 23.620 63.310 23.650 ;
        RECT 63.320 23.620 65.050 23.770 ;
        RECT 55.500 17.590 57.250 17.610 ;
        RECT 62.590 17.570 66.010 23.620 ;
        RECT 110.040 -5.660 111.390 9.810 ;
        RECT 110.030 -6.130 111.390 -5.660 ;
      LAYER met3 ;
        RECT 79.410 46.940 79.860 47.690 ;
        RECT 79.410 40.780 79.780 46.940 ;
        RECT 80.450 46.930 80.900 47.680 ;
        RECT 80.530 44.290 80.900 46.930 ;
        RECT 80.530 43.690 80.970 44.290 ;
        RECT 79.410 40.450 79.900 40.780 ;
        RECT 79.460 40.290 79.900 40.450 ;
        RECT 80.530 38.580 80.900 43.690 ;
        RECT 80.520 37.710 80.990 38.580 ;
    END
  END DIG26
  PIN DIG25
    ANTENNAGATEAREA 43.185299 ;
    ANTENNADIFFAREA 248.747787 ;
    PORT
      LAYER met2 ;
        RECT 2.950 62.460 3.630 63.680 ;
        RECT 4.180 62.460 4.630 62.560 ;
        RECT 2.950 62.230 4.630 62.460 ;
        RECT 2.950 61.360 3.630 62.230 ;
        RECT 4.180 62.130 4.630 62.230 ;
        RECT 9.150 59.710 9.470 60.030 ;
        RECT 4.280 58.660 4.710 59.130 ;
        RECT 9.170 58.670 9.440 59.710 ;
        RECT 6.650 58.660 9.440 58.670 ;
        RECT 4.280 58.650 9.440 58.660 ;
        RECT 4.370 58.440 9.440 58.650 ;
        RECT 4.370 58.430 8.920 58.440 ;
        RECT 34.590 52.740 34.900 52.760 ;
        RECT 24.800 52.660 25.120 52.670 ;
        RECT 34.590 52.660 34.910 52.740 ;
        RECT 58.770 52.670 59.090 52.690 ;
        RECT 58.770 52.660 59.100 52.670 ;
        RECT 65.540 52.660 65.860 52.690 ;
        RECT 80.310 52.660 80.630 52.680 ;
        RECT 94.970 52.660 95.530 52.800 ;
        RECT 24.800 52.430 95.530 52.660 ;
        RECT 24.800 52.350 25.120 52.430 ;
        RECT 34.590 52.420 34.900 52.430 ;
        RECT 58.770 52.410 59.100 52.430 ;
        RECT 65.540 52.410 65.860 52.430 ;
        RECT 80.310 52.420 80.630 52.430 ;
        RECT 94.970 52.290 95.530 52.430 ;
        RECT 30.590 52.210 30.960 52.270 ;
        RECT 93.790 52.210 94.330 52.230 ;
        RECT 30.590 51.980 94.330 52.210 ;
        RECT 30.590 51.920 30.960 51.980 ;
        RECT 62.390 51.760 62.670 51.770 ;
        RECT 33.420 51.750 33.730 51.760 ;
        RECT 62.370 51.750 62.690 51.760 ;
        RECT 65.100 51.750 65.420 51.780 ;
        RECT 79.420 51.750 79.740 51.810 ;
        RECT 92.710 51.750 93.250 51.760 ;
        RECT 33.420 51.520 93.250 51.750 ;
        RECT 93.790 51.670 94.330 51.980 ;
        RECT 33.420 51.490 33.750 51.520 ;
        RECT 62.370 51.500 62.690 51.520 ;
        RECT 65.100 51.500 65.420 51.520 ;
        RECT 62.390 51.490 62.670 51.500 ;
        RECT 33.420 51.470 33.730 51.490 ;
        RECT 27.340 51.290 27.660 51.300 ;
        RECT 91.770 51.290 92.300 51.320 ;
        RECT 2.460 51.060 2.970 51.080 ;
        RECT 22.100 51.060 22.500 51.070 ;
        RECT 2.460 50.710 22.500 51.060 ;
        RECT 27.340 51.060 92.300 51.290 ;
        RECT 92.710 51.200 93.250 51.520 ;
        RECT 27.340 51.000 27.660 51.060 ;
        RECT 91.770 50.710 92.300 51.060 ;
        RECT 2.460 50.670 2.970 50.710 ;
        RECT 22.100 50.680 22.500 50.710 ;
        RECT 71.660 50.130 71.940 50.150 ;
        RECT 71.640 50.100 71.960 50.130 ;
        RECT 103.780 50.100 105.120 50.640 ;
        RECT 71.640 49.890 105.120 50.100 ;
        RECT 71.640 49.870 71.960 49.890 ;
        RECT 71.660 49.850 71.940 49.870 ;
        RECT 103.780 49.360 105.120 49.890 ;
        RECT 22.480 48.050 22.770 48.070 ;
        RECT 10.030 47.650 22.790 48.050 ;
        RECT 2.470 44.960 3.740 45.830 ;
        RECT 10.030 44.960 10.430 47.650 ;
        RECT 22.480 47.640 22.770 47.650 ;
        RECT 79.360 47.340 79.940 47.780 ;
        RECT 79.360 47.150 80.000 47.340 ;
        RECT 20.980 46.750 21.290 46.840 ;
        RECT 22.490 46.750 22.810 46.800 ;
        RECT 20.980 46.580 22.870 46.750 ;
        RECT 20.980 46.510 21.290 46.580 ;
        RECT 22.490 46.540 22.810 46.580 ;
        RECT 79.760 46.540 80.000 47.150 ;
        RECT 80.380 47.140 80.960 47.770 ;
        RECT 18.720 46.330 19.040 46.380 ;
        RECT 19.420 46.330 19.740 46.410 ;
        RECT 111.850 46.370 112.170 46.630 ;
        RECT 118.130 46.520 118.490 46.530 ;
        RECT 104.280 46.340 104.580 46.360 ;
        RECT 111.890 46.350 113.070 46.370 ;
        RECT 111.890 46.340 113.110 46.350 ;
        RECT 117.570 46.340 118.490 46.520 ;
        RECT 18.720 46.160 19.740 46.330 ;
        RECT 18.720 46.120 19.040 46.160 ;
        RECT 19.420 46.090 19.740 46.160 ;
        RECT 104.270 46.240 118.490 46.340 ;
        RECT 104.270 45.920 118.530 46.240 ;
        RECT 20.980 45.830 21.290 45.920 ;
        RECT 104.280 45.900 104.580 45.920 ;
        RECT 22.490 45.830 22.810 45.880 ;
        RECT 20.980 45.660 22.870 45.830 ;
        RECT 111.850 45.770 112.170 45.920 ;
        RECT 20.980 45.590 21.290 45.660 ;
        RECT 22.490 45.620 22.810 45.660 ;
        RECT 117.570 45.580 118.530 45.920 ;
        RECT 18.690 45.410 19.010 45.460 ;
        RECT 19.420 45.410 19.740 45.490 ;
        RECT 18.690 45.240 19.740 45.410 ;
        RECT 110.520 45.390 110.830 45.400 ;
        RECT 109.950 45.380 110.830 45.390 ;
        RECT 18.690 45.200 19.010 45.240 ;
        RECT 19.420 45.170 19.740 45.240 ;
        RECT 109.880 45.140 110.830 45.380 ;
        RECT 110.520 45.070 110.830 45.140 ;
        RECT 111.490 45.070 111.800 45.120 ;
        RECT 113.740 45.070 114.050 45.170 ;
        RECT 2.470 44.560 10.430 44.960 ;
        RECT 20.980 44.910 21.290 45.000 ;
        RECT 22.460 44.910 22.780 44.960 ;
        RECT 110.910 44.950 111.220 45.020 ;
        RECT 111.490 44.950 114.050 45.070 ;
        RECT 20.980 44.740 22.870 44.910 ;
        RECT 110.910 44.840 114.050 44.950 ;
        RECT 110.910 44.740 113.240 44.840 ;
        RECT 20.980 44.670 21.290 44.740 ;
        RECT 22.460 44.700 22.780 44.740 ;
        RECT 110.910 44.690 111.220 44.740 ;
        RECT 2.470 43.950 3.740 44.560 ;
        RECT 18.700 44.490 19.020 44.540 ;
        RECT 19.420 44.490 19.740 44.570 ;
        RECT 110.670 44.530 110.980 44.570 ;
        RECT 18.700 44.320 19.740 44.490 ;
        RECT 110.490 44.390 111.210 44.530 ;
        RECT 111.440 44.390 111.750 44.470 ;
        RECT 18.700 44.280 19.020 44.320 ;
        RECT 19.420 44.250 19.740 44.320 ;
        RECT 89.660 44.100 98.810 44.330 ;
        RECT 110.490 44.280 111.750 44.390 ;
        RECT 110.670 44.240 111.750 44.280 ;
        RECT 110.940 44.180 111.750 44.240 ;
        RECT 110.940 44.170 111.210 44.180 ;
        RECT 111.440 44.140 111.750 44.180 ;
        RECT 117.630 44.150 118.530 45.580 ;
        RECT 98.520 44.000 98.810 44.100 ;
        RECT 108.310 44.000 109.430 44.010 ;
        RECT 109.550 44.000 109.860 44.030 ;
        RECT 98.520 43.860 111.070 44.000 ;
        RECT 98.520 43.800 113.240 43.860 ;
        RECT 98.520 43.790 98.810 43.800 ;
        RECT 101.710 43.700 113.240 43.800 ;
        RECT 109.080 43.670 109.550 43.700 ;
        RECT 110.650 43.680 113.240 43.700 ;
        RECT 110.650 43.670 111.070 43.680 ;
        RECT 111.010 43.600 111.210 43.610 ;
        RECT 111.010 43.590 111.230 43.600 ;
        RECT 111.440 43.590 111.750 43.630 ;
        RECT 18.050 43.480 18.370 43.520 ;
        RECT 19.700 43.480 20.020 43.540 ;
        RECT 111.010 43.520 111.750 43.590 ;
        RECT 110.720 43.500 111.750 43.520 ;
        RECT 18.050 43.290 20.020 43.480 ;
        RECT 18.050 43.260 18.370 43.290 ;
        RECT 19.700 43.220 20.020 43.290 ;
        RECT 89.660 43.380 97.870 43.500 ;
        RECT 110.670 43.380 111.750 43.500 ;
        RECT 89.660 43.280 105.810 43.380 ;
        RECT 97.650 43.180 105.810 43.280 ;
        RECT 110.670 43.260 111.230 43.380 ;
        RECT 111.440 43.300 111.750 43.380 ;
        RECT 110.670 43.250 111.140 43.260 ;
        RECT 18.010 42.520 18.330 42.560 ;
        RECT 19.700 42.520 20.020 42.580 ;
        RECT 18.010 42.330 20.020 42.520 ;
        RECT 18.010 42.300 18.330 42.330 ;
        RECT 19.700 42.260 20.020 42.330 ;
        RECT 97.650 42.500 97.870 43.180 ;
        RECT 100.270 43.020 100.730 43.150 ;
        RECT 105.590 43.020 105.810 43.180 ;
        RECT 110.000 43.020 110.320 43.060 ;
        RECT 111.010 43.020 111.330 43.050 ;
        RECT 100.270 42.820 108.050 43.020 ;
        RECT 109.950 42.930 113.710 43.020 ;
        RECT 113.790 42.930 114.100 42.950 ;
        RECT 109.950 42.820 114.410 42.930 ;
        RECT 100.270 42.700 100.730 42.820 ;
        RECT 104.410 42.500 104.630 42.510 ;
        RECT 97.650 42.370 104.660 42.500 ;
        RECT 105.590 42.460 105.810 42.820 ;
        RECT 107.730 42.730 108.050 42.820 ;
        RECT 110.000 42.800 110.320 42.820 ;
        RECT 111.010 42.790 111.330 42.820 ;
        RECT 110.280 42.710 110.590 42.750 ;
        RECT 109.960 42.700 110.620 42.710 ;
        RECT 111.490 42.700 114.410 42.820 ;
        RECT 109.960 42.470 111.060 42.700 ;
        RECT 111.490 42.650 111.800 42.700 ;
        RECT 105.560 42.420 105.810 42.460 ;
        RECT 105.560 42.370 105.820 42.420 ;
        RECT 107.730 42.370 108.050 42.460 ;
        RECT 110.280 42.420 110.590 42.470 ;
        RECT 110.000 42.370 110.320 42.390 ;
        RECT 111.010 42.370 111.330 42.400 ;
        RECT 113.510 42.370 113.710 42.700 ;
        RECT 113.790 42.620 114.100 42.700 ;
        RECT 97.650 42.250 108.050 42.370 ;
        RECT 18.050 41.560 18.370 41.600 ;
        RECT 19.700 41.560 20.020 41.620 ;
        RECT 18.050 41.370 20.020 41.560 ;
        RECT 18.050 41.340 18.370 41.370 ;
        RECT 19.700 41.300 20.020 41.370 ;
        RECT 97.650 41.520 97.870 42.250 ;
        RECT 101.280 42.170 108.050 42.250 ;
        RECT 109.950 42.170 113.710 42.370 ;
        RECT 101.280 42.050 101.640 42.170 ;
        RECT 97.650 41.390 101.340 41.520 ;
        RECT 104.370 41.390 104.660 42.170 ;
        RECT 105.560 41.780 105.820 42.170 ;
        RECT 110.000 42.130 110.320 42.170 ;
        RECT 111.010 42.140 111.330 42.170 ;
        RECT 111.490 42.100 111.800 42.160 ;
        RECT 113.510 42.100 113.710 42.170 ;
        RECT 113.780 42.100 114.090 42.230 ;
        RECT 111.490 41.880 114.410 42.100 ;
        RECT 111.490 41.830 111.800 41.880 ;
        RECT 105.560 41.570 109.690 41.780 ;
        RECT 109.080 41.400 109.390 41.520 ;
        RECT 109.480 41.430 109.690 41.570 ;
        RECT 110.650 41.430 110.960 41.520 ;
        RECT 111.440 41.430 111.750 41.510 ;
        RECT 108.310 41.390 109.430 41.400 ;
        RECT 109.480 41.390 111.750 41.430 ;
        RECT 97.650 41.220 111.750 41.390 ;
        RECT 97.650 41.190 110.960 41.220 ;
        RECT 97.650 41.180 99.250 41.190 ;
        RECT 62.370 41.090 62.680 41.100 ;
        RECT 62.360 41.030 62.690 41.090 ;
        RECT 62.010 40.980 62.690 41.030 ;
        RECT 58.780 40.900 62.690 40.980 ;
        RECT 64.010 40.950 65.960 41.090 ;
        RECT 101.110 40.980 101.340 41.190 ;
        RECT 104.370 41.080 104.660 41.190 ;
        RECT 108.310 41.180 109.430 41.190 ;
        RECT 111.440 41.180 111.750 41.220 ;
        RECT 113.510 41.120 113.710 41.880 ;
        RECT 117.600 41.120 118.500 41.790 ;
        RECT 104.370 40.980 107.260 41.080 ;
        RECT 108.310 40.980 109.430 40.990 ;
        RECT 63.940 40.930 65.960 40.950 ;
        RECT 63.940 40.900 64.260 40.930 ;
        RECT 64.740 40.920 65.960 40.930 ;
        RECT 65.440 40.910 65.960 40.920 ;
        RECT 58.780 40.760 64.260 40.900 ;
        RECT 89.660 40.780 110.960 40.980 ;
        RECT 61.530 40.710 64.260 40.760 ;
        RECT 61.530 40.660 61.850 40.710 ;
        RECT 63.940 40.690 64.260 40.710 ;
        RECT 101.110 40.730 101.340 40.780 ;
        RECT 108.310 40.770 109.430 40.780 ;
        RECT 101.110 40.580 101.330 40.730 ;
        RECT 109.080 40.650 109.390 40.770 ;
        RECT 110.650 40.650 110.960 40.780 ;
        RECT 113.510 40.690 118.500 41.120 ;
        RECT 111.440 40.630 111.750 40.670 ;
        RECT 105.480 40.580 111.750 40.630 ;
        RECT 101.110 40.420 111.750 40.580 ;
        RECT 101.110 40.360 105.870 40.420 ;
        RECT 111.440 40.340 111.750 40.420 ;
        RECT 102.200 40.110 102.590 40.130 ;
        RECT 102.190 40.000 102.600 40.110 ;
        RECT 110.000 40.000 110.320 40.040 ;
        RECT 111.010 40.000 111.330 40.030 ;
        RECT 111.490 40.000 111.800 40.020 ;
        RECT 113.510 40.000 113.710 40.690 ;
        RECT 102.190 39.800 108.050 40.000 ;
        RECT 109.950 39.980 113.710 40.000 ;
        RECT 109.950 39.940 114.010 39.980 ;
        RECT 109.950 39.800 114.200 39.940 ;
        RECT 102.190 39.710 102.600 39.800 ;
        RECT 107.730 39.710 108.050 39.800 ;
        RECT 110.000 39.780 110.320 39.800 ;
        RECT 110.920 39.770 111.330 39.800 ;
        RECT 110.920 39.710 111.240 39.770 ;
        RECT 94.730 39.560 111.240 39.710 ;
        RECT 111.490 39.710 114.200 39.800 ;
        RECT 111.490 39.690 111.800 39.710 ;
        RECT 113.510 39.650 114.010 39.710 ;
        RECT 117.600 39.700 118.500 40.690 ;
        RECT 94.730 39.410 95.050 39.560 ;
        RECT 100.530 39.410 100.850 39.560 ;
        RECT 103.020 39.410 103.420 39.420 ;
        RECT 103.000 39.350 103.440 39.410 ;
        RECT 107.730 39.350 108.050 39.440 ;
        RECT 110.000 39.350 110.320 39.370 ;
        RECT 111.010 39.350 111.330 39.380 ;
        RECT 113.510 39.350 113.710 39.650 ;
        RECT 103.000 39.150 108.050 39.350 ;
        RECT 109.950 39.230 113.710 39.350 ;
        RECT 109.950 39.150 113.680 39.230 ;
        RECT 103.020 39.140 103.420 39.150 ;
        RECT 110.000 39.110 110.320 39.150 ;
        RECT 111.010 39.120 111.330 39.150 ;
        RECT 94.880 30.500 95.480 30.560 ;
        RECT 117.600 30.500 118.500 31.530 ;
        RECT 94.880 30.030 118.500 30.500 ;
        RECT 94.880 29.980 95.480 30.030 ;
        RECT 117.600 29.440 118.500 30.030 ;
        RECT 18.010 26.530 18.320 26.550 ;
        RECT 18.670 26.530 18.980 26.550 ;
        RECT 18.010 26.060 25.330 26.530 ;
        RECT 18.010 26.040 18.320 26.060 ;
        RECT 18.670 26.040 18.980 26.060 ;
        RECT 24.860 25.380 25.330 26.060 ;
        RECT 57.140 25.540 57.450 25.670 ;
        RECT 64.940 25.540 65.080 25.560 ;
        RECT 54.970 25.380 65.080 25.540 ;
        RECT 117.630 25.380 118.530 26.350 ;
        RECT 16.680 25.250 16.940 25.320 ;
        RECT 18.730 25.250 19.050 25.270 ;
        RECT 20.490 25.250 20.820 25.290 ;
        RECT 16.680 25.060 20.820 25.250 ;
        RECT 16.680 25.000 16.940 25.060 ;
        RECT 18.730 25.010 19.050 25.060 ;
        RECT 20.490 25.020 20.820 25.060 ;
        RECT 24.860 24.910 118.530 25.380 ;
        RECT 16.130 24.850 16.450 24.890 ;
        RECT 18.070 24.850 18.390 24.910 ;
        RECT 20.990 24.850 21.310 24.890 ;
        RECT 16.130 24.660 21.310 24.850 ;
        RECT 57.140 24.790 57.450 24.910 ;
        RECT 93.790 24.790 94.360 24.910 ;
        RECT 16.130 24.630 16.450 24.660 ;
        RECT 18.070 24.650 18.390 24.660 ;
        RECT 20.990 24.630 21.310 24.660 ;
        RECT 19.470 24.270 19.780 24.340 ;
        RECT 22.470 24.290 22.770 24.310 ;
        RECT 22.460 24.270 22.780 24.290 ;
        RECT 19.470 24.060 22.780 24.270 ;
        RECT 117.630 24.260 118.530 24.910 ;
        RECT 19.470 24.010 19.780 24.060 ;
        RECT 20.240 24.050 22.780 24.060 ;
        RECT 18.300 23.830 18.610 23.900 ;
        RECT 20.240 23.830 20.460 24.050 ;
        RECT 22.460 24.030 22.780 24.050 ;
        RECT 22.470 24.010 22.770 24.030 ;
        RECT 18.300 23.610 20.460 23.830 ;
        RECT 18.300 23.570 18.610 23.610 ;
        RECT 57.140 23.530 57.450 23.550 ;
        RECT 54.980 23.370 65.050 23.530 ;
        RECT 54.980 23.360 65.040 23.370 ;
        RECT 54.980 23.350 57.540 23.360 ;
        RECT 57.140 23.220 57.450 23.350 ;
        RECT 60.400 23.340 60.720 23.360 ;
        RECT 19.980 23.110 20.300 23.170 ;
        RECT 21.850 23.140 22.140 23.160 ;
        RECT 60.400 23.150 68.320 23.340 ;
        RECT 68.480 23.150 68.790 23.190 ;
        RECT 19.980 23.100 20.460 23.110 ;
        RECT 21.840 23.100 22.160 23.140 ;
        RECT 60.400 23.130 68.790 23.150 ;
        RECT 60.400 23.100 60.720 23.130 ;
        RECT 61.530 23.100 64.260 23.130 ;
        RECT 19.980 22.910 22.160 23.100 ;
        RECT 61.530 23.050 65.960 23.100 ;
        RECT 61.530 22.970 61.850 23.050 ;
        RECT 63.940 23.000 65.960 23.050 ;
        RECT 63.980 22.930 65.960 23.000 ;
        RECT 68.110 22.940 68.790 23.130 ;
        RECT 65.440 22.920 65.960 22.930 ;
        RECT 19.980 22.900 20.460 22.910 ;
        RECT 19.980 22.850 20.300 22.900 ;
        RECT 21.840 22.880 22.160 22.910 ;
        RECT 21.850 22.860 22.140 22.880 ;
        RECT 68.480 22.860 68.790 22.940 ;
        RECT 57.130 22.710 57.280 22.720 ;
        RECT 56.110 22.670 57.280 22.710 ;
        RECT 56.110 22.560 57.450 22.670 ;
        RECT 56.050 22.540 56.330 22.560 ;
        RECT 57.130 22.550 57.450 22.560 ;
        RECT 60.290 22.550 60.770 22.760 ;
        RECT 57.130 22.540 65.050 22.550 ;
        RECT 17.150 22.500 17.470 22.520 ;
        RECT 16.930 22.280 17.470 22.500 ;
        RECT 54.980 22.380 65.050 22.540 ;
        RECT 54.980 22.360 57.540 22.380 ;
        RECT 17.150 22.260 17.470 22.280 ;
        RECT 56.050 22.230 56.330 22.360 ;
        RECT 57.130 22.340 57.450 22.360 ;
        RECT 57.130 22.210 57.280 22.340 ;
        RECT 60.380 22.210 60.700 22.310 ;
        RECT 62.720 22.290 64.260 22.380 ;
        RECT 57.130 22.110 60.700 22.210 ;
        RECT 54.980 22.050 60.700 22.110 ;
        RECT 19.900 21.920 20.220 22.040 ;
        RECT 54.980 21.940 57.550 22.050 ;
        RECT 54.980 21.930 57.450 21.940 ;
        RECT 16.930 21.720 20.220 21.920 ;
        RECT 57.140 21.810 57.450 21.930 ;
        RECT 57.110 21.790 57.450 21.810 ;
        RECT 16.930 21.710 19.910 21.720 ;
        RECT 57.110 21.550 57.430 21.790 ;
        RECT 60.430 21.590 60.770 21.660 ;
        RECT 57.180 21.540 57.350 21.550 ;
        RECT 16.930 21.500 19.910 21.520 ;
        RECT 16.930 21.310 20.230 21.500 ;
        RECT 60.290 21.360 60.770 21.590 ;
        RECT 19.910 21.180 20.230 21.310 ;
        RECT 60.340 21.070 60.570 21.080 ;
        RECT 61.530 21.070 61.850 21.150 ;
        RECT 64.010 21.120 65.960 21.260 ;
        RECT 63.940 21.100 65.960 21.120 ;
        RECT 63.940 21.070 64.260 21.100 ;
        RECT 64.740 21.090 65.960 21.100 ;
        RECT 65.440 21.080 65.960 21.090 ;
        RECT 60.340 21.040 67.910 21.070 ;
        RECT 16.160 20.980 16.450 20.990 ;
        RECT 16.150 20.960 16.470 20.980 ;
        RECT 17.150 20.960 17.470 20.970 ;
        RECT 16.150 20.740 17.470 20.960 ;
        RECT 60.340 20.870 67.970 21.040 ;
        RECT 68.480 20.870 68.790 20.950 ;
        RECT 16.150 20.720 16.470 20.740 ;
        RECT 16.160 20.700 16.450 20.720 ;
        RECT 17.150 20.710 17.470 20.740 ;
        RECT 57.090 20.770 57.410 20.800 ;
        RECT 60.340 20.770 60.580 20.870 ;
        RECT 61.530 20.830 61.850 20.870 ;
        RECT 63.940 20.860 64.260 20.870 ;
        RECT 57.090 20.590 60.580 20.770 ;
        RECT 67.780 20.670 68.790 20.870 ;
        RECT 68.380 20.660 68.790 20.670 ;
        RECT 68.480 20.620 68.790 20.660 ;
        RECT 57.090 20.570 60.500 20.590 ;
        RECT 19.960 20.500 20.280 20.550 ;
        RECT 21.420 20.500 21.740 20.550 ;
        RECT 57.090 20.540 57.410 20.570 ;
        RECT 19.960 20.290 21.740 20.500 ;
        RECT 19.960 20.230 20.280 20.290 ;
        RECT 21.420 20.250 21.740 20.290 ;
        RECT 60.380 20.390 60.700 20.430 ;
        RECT 60.380 20.370 67.930 20.390 ;
        RECT 68.480 20.380 68.790 20.420 ;
        RECT 68.380 20.370 68.790 20.380 ;
        RECT 60.380 20.170 68.790 20.370 ;
        RECT 60.480 20.160 60.800 20.170 ;
        RECT 61.530 20.120 64.260 20.170 ;
        RECT 61.530 20.040 61.850 20.120 ;
        RECT 63.940 20.110 64.260 20.120 ;
        RECT 63.940 20.070 65.960 20.110 ;
        RECT 68.480 20.090 68.790 20.170 ;
        RECT 92.670 20.140 93.220 20.150 ;
        RECT 92.670 20.120 93.230 20.140 ;
        RECT 117.600 20.120 118.500 21.270 ;
        RECT 64.050 19.950 65.960 20.070 ;
        RECT 64.770 19.930 65.960 19.950 ;
        RECT 56.660 19.710 56.980 19.760 ;
        RECT 56.660 19.440 57.270 19.710 ;
        RECT 60.290 19.600 60.770 19.830 ;
        RECT 92.670 19.650 118.500 20.120 ;
        RECT 92.670 19.640 93.230 19.650 ;
        RECT 92.670 19.620 93.220 19.640 ;
        RECT 60.430 19.530 60.770 19.600 ;
        RECT 57.070 19.210 57.270 19.440 ;
        RECT 60.220 19.210 60.540 19.250 ;
        RECT 57.070 19.010 60.620 19.210 ;
        RECT 117.600 19.180 118.500 19.650 ;
        RECT 60.220 18.990 60.540 19.010 ;
        RECT 17.260 17.920 17.570 17.930 ;
        RECT 18.350 17.920 18.660 17.930 ;
        RECT 15.940 17.910 18.660 17.920 ;
        RECT 15.710 17.600 18.660 17.910 ;
        RECT 15.710 17.590 18.650 17.600 ;
        RECT 15.710 15.970 16.060 17.590 ;
        RECT 49.450 17.340 49.770 17.390 ;
        RECT 56.060 17.340 56.380 17.440 ;
        RECT 16.710 17.240 17.020 17.250 ;
        RECT 17.810 17.240 18.120 17.250 ;
        RECT 18.910 17.240 19.220 17.250 ;
        RECT 16.680 16.920 19.840 17.240 ;
        RECT 49.450 17.180 56.380 17.340 ;
        RECT 49.450 17.130 49.770 17.180 ;
        RECT 56.060 17.160 56.380 17.180 ;
        RECT 97.860 17.310 98.420 17.380 ;
        RECT 110.580 17.310 111.260 17.370 ;
        RECT 118.110 17.310 118.770 17.950 ;
        RECT 56.650 17.100 56.930 17.110 ;
        RECT 48.920 17.050 49.250 17.070 ;
        RECT 19.520 15.970 19.840 16.920 ;
        RECT 48.910 16.970 49.260 17.050 ;
        RECT 54.660 16.970 54.980 17.030 ;
        RECT 56.630 17.010 56.950 17.100 ;
        RECT 58.870 17.010 59.190 17.040 ;
        RECT 48.910 16.810 54.980 16.970 ;
        RECT 56.600 16.850 59.190 17.010 ;
        RECT 97.860 16.900 118.770 17.310 ;
        RECT 97.860 16.850 98.420 16.900 ;
        RECT 56.630 16.840 56.950 16.850 ;
        RECT 56.650 16.830 56.930 16.840 ;
        RECT 48.910 16.740 49.270 16.810 ;
        RECT 54.660 16.760 54.980 16.810 ;
        RECT 58.870 16.780 59.190 16.850 ;
        RECT 110.580 16.840 111.260 16.900 ;
        RECT 118.110 16.800 118.770 16.900 ;
        RECT 58.890 16.770 59.170 16.780 ;
        RECT 49.160 16.710 49.270 16.740 ;
        RECT 44.490 16.350 44.820 16.590 ;
        RECT 50.350 16.480 50.650 16.490 ;
        RECT 50.340 16.350 50.660 16.480 ;
        RECT 60.880 16.350 61.160 16.650 ;
        RECT 64.910 16.350 65.210 16.630 ;
        RECT 44.490 16.330 65.210 16.350 ;
        RECT 44.490 16.300 65.200 16.330 ;
        RECT 44.490 16.190 65.140 16.300 ;
        RECT 48.300 15.970 48.740 15.980 ;
        RECT 2.980 15.960 48.740 15.970 ;
        RECT 2.980 15.550 48.760 15.960 ;
        RECT 15.710 15.150 16.060 15.550 ;
        RECT 15.710 15.000 18.660 15.150 ;
        RECT 19.520 15.000 19.840 15.550 ;
        RECT 41.450 15.540 41.930 15.550 ;
        RECT 48.280 15.540 48.760 15.550 ;
        RECT 48.300 15.530 48.740 15.540 ;
        RECT 57.670 15.500 58.050 15.890 ;
        RECT 58.820 15.460 59.220 15.800 ;
        RECT 2.960 14.580 44.940 15.000 ;
        RECT 15.710 13.950 16.060 14.580 ;
        RECT 15.710 13.820 16.090 13.950 ;
        RECT 15.710 13.780 16.460 13.820 ;
        RECT 17.260 13.780 17.570 13.800 ;
        RECT 15.710 13.480 18.660 13.780 ;
        RECT 17.260 13.470 17.570 13.480 ;
        RECT 18.350 13.450 18.660 13.480 ;
        RECT 16.710 13.100 17.020 13.110 ;
        RECT 19.520 13.100 19.840 14.580 ;
        RECT 26.010 14.080 26.840 14.580 ;
        RECT 48.970 14.460 49.350 14.840 ;
        RECT 91.620 14.820 92.220 14.870 ;
        RECT 118.030 14.820 120.130 15.760 ;
        RECT 91.620 14.350 120.130 14.820 ;
        RECT 91.620 14.310 92.220 14.350 ;
        RECT 118.030 13.680 120.130 14.350 ;
        RECT 118.050 13.670 118.820 13.680 ;
        RECT 16.690 12.770 19.840 13.100 ;
        RECT 16.690 12.760 19.750 12.770 ;
        RECT 19.600 12.560 19.890 12.580 ;
        RECT 21.830 12.560 22.140 12.580 ;
        RECT 19.590 12.200 22.140 12.560 ;
        RECT 19.600 12.180 19.890 12.200 ;
        RECT 21.830 12.180 22.140 12.200 ;
        RECT 58.380 11.690 61.440 11.700 ;
        RECT 58.290 11.670 61.440 11.690 ;
        RECT 48.570 11.660 51.630 11.670 ;
        RECT 48.480 11.330 51.630 11.660 ;
        RECT 55.410 11.360 61.440 11.670 ;
        RECT 65.220 11.690 68.280 11.700 ;
        RECT 65.220 11.360 68.370 11.690 ;
        RECT 55.410 11.330 58.610 11.360 ;
        RECT 61.110 11.350 61.420 11.360 ;
        RECT 65.240 11.350 65.550 11.360 ;
        RECT 17.300 10.360 17.610 10.370 ;
        RECT 18.390 10.360 18.700 10.370 ;
        RECT 15.980 10.350 18.700 10.360 ;
        RECT 15.750 10.040 18.700 10.350 ;
        RECT 15.750 10.030 18.690 10.040 ;
        RECT 15.750 7.590 16.100 10.030 ;
        RECT 16.750 9.680 17.060 9.690 ;
        RECT 17.850 9.680 18.160 9.690 ;
        RECT 18.950 9.680 19.260 9.690 ;
        RECT 16.720 9.360 19.880 9.680 ;
        RECT 19.560 8.900 19.880 9.360 ;
        RECT 22.460 8.900 22.740 8.910 ;
        RECT 18.870 8.570 22.760 8.900 ;
        RECT 48.480 8.880 48.800 11.330 ;
        RECT 51.300 11.320 51.610 11.330 ;
        RECT 55.430 11.320 55.740 11.330 ;
        RECT 49.660 10.950 49.970 10.980 ;
        RECT 50.750 10.950 51.060 10.960 ;
        RECT 55.980 10.950 56.290 10.960 ;
        RECT 57.070 10.950 57.380 10.980 ;
        RECT 49.660 10.650 52.610 10.950 ;
        RECT 50.750 10.630 51.060 10.650 ;
        RECT 51.860 10.610 52.610 10.650 ;
        RECT 52.230 10.480 52.610 10.610 ;
        RECT 52.260 9.610 52.610 10.480 ;
        RECT 54.430 10.650 57.380 10.950 ;
        RECT 54.430 10.610 55.180 10.650 ;
        RECT 55.980 10.630 56.290 10.650 ;
        RECT 54.430 10.480 54.810 10.610 ;
        RECT 54.430 10.050 54.780 10.480 ;
        RECT 58.240 10.050 58.610 11.330 ;
        RECT 59.470 10.980 59.780 11.010 ;
        RECT 60.560 10.980 60.870 10.990 ;
        RECT 65.790 10.980 66.100 10.990 ;
        RECT 66.880 10.980 67.190 11.010 ;
        RECT 59.470 10.680 62.420 10.980 ;
        RECT 60.560 10.660 60.870 10.680 ;
        RECT 61.670 10.640 62.420 10.680 ;
        RECT 62.040 10.510 62.420 10.640 ;
        RECT 62.070 10.050 62.420 10.510 ;
        RECT 64.240 10.680 67.190 10.980 ;
        RECT 64.240 10.640 64.990 10.680 ;
        RECT 65.790 10.660 66.100 10.680 ;
        RECT 64.240 10.510 64.620 10.640 ;
        RECT 52.990 10.020 63.890 10.050 ;
        RECT 52.980 9.770 63.890 10.020 ;
        RECT 52.980 9.740 53.320 9.770 ;
        RECT 53.720 9.760 54.060 9.770 ;
        RECT 49.660 9.280 52.610 9.610 ;
        RECT 49.060 9.230 49.560 9.240 ;
        RECT 52.260 9.230 52.610 9.280 ;
        RECT 54.430 9.610 54.780 9.770 ;
        RECT 54.430 9.280 57.380 9.610 ;
        RECT 54.430 9.230 54.780 9.280 ;
        RECT 58.240 9.230 58.610 9.770 ;
        RECT 62.070 9.640 62.420 9.770 ;
        RECT 62.790 9.740 63.130 9.770 ;
        RECT 59.470 9.310 62.420 9.640 ;
        RECT 62.070 9.230 62.420 9.310 ;
        RECT 64.240 9.640 64.590 10.510 ;
        RECT 64.240 9.310 67.190 9.640 ;
        RECT 64.240 9.230 64.590 9.310 ;
        RECT 68.050 9.230 68.370 11.360 ;
        RECT 70.960 11.670 74.020 11.680 ;
        RECT 70.960 11.340 74.110 11.670 ;
        RECT 70.980 11.330 71.290 11.340 ;
        RECT 71.530 10.960 71.840 10.970 ;
        RECT 72.620 10.960 72.930 10.990 ;
        RECT 69.980 10.660 72.930 10.960 ;
        RECT 69.980 10.620 70.730 10.660 ;
        RECT 71.530 10.640 71.840 10.660 ;
        RECT 69.980 10.490 70.360 10.620 ;
        RECT 69.980 9.620 70.330 10.490 ;
        RECT 69.980 9.290 72.930 9.620 ;
        RECT 69.980 9.230 70.330 9.290 ;
        RECT 73.790 9.230 74.110 11.340 ;
        RECT 94.990 9.230 95.550 9.250 ;
        RECT 49.060 8.880 95.550 9.230 ;
        RECT 48.480 8.770 95.550 8.880 ;
        RECT 19.560 8.320 19.880 8.570 ;
        RECT 22.460 8.550 22.740 8.570 ;
        RECT 48.480 8.550 51.640 8.770 ;
        RECT 16.720 7.990 19.880 8.320 ;
        RECT 15.750 7.260 18.700 7.590 ;
        RECT 15.040 7.220 15.390 7.250 ;
        RECT 15.750 7.220 16.100 7.260 ;
        RECT 19.560 7.220 19.880 7.990 ;
        RECT 48.480 7.510 48.800 8.550 ;
        RECT 21.420 7.240 21.750 7.280 ;
        RECT 21.410 7.220 21.760 7.240 ;
        RECT 15.040 6.960 25.070 7.220 ;
        RECT 48.480 7.190 51.640 7.510 ;
        RECT 49.100 7.180 49.410 7.190 ;
        RECT 50.200 7.180 50.510 7.190 ;
        RECT 51.300 7.180 51.610 7.190 ;
        RECT 15.080 6.930 25.070 6.960 ;
        RECT 15.750 6.390 16.100 6.930 ;
        RECT 19.560 6.590 19.880 6.930 ;
        RECT 21.420 6.910 21.750 6.930 ;
        RECT 15.750 6.260 16.130 6.390 ;
        RECT 15.750 6.220 16.500 6.260 ;
        RECT 18.880 6.250 21.220 6.590 ;
        RECT 17.300 6.220 17.610 6.240 ;
        RECT 15.750 5.920 18.700 6.220 ;
        RECT 18.880 6.010 21.260 6.250 ;
        RECT 18.880 5.990 21.220 6.010 ;
        RECT 17.300 5.910 17.610 5.920 ;
        RECT 18.390 5.890 18.700 5.920 ;
        RECT 16.750 5.540 17.060 5.550 ;
        RECT 19.560 5.540 19.880 5.990 ;
        RECT 20.250 5.920 20.910 5.990 ;
        RECT 20.280 5.910 20.880 5.920 ;
        RECT 16.730 5.210 19.880 5.540 ;
        RECT 16.730 5.200 19.790 5.210 ;
        RECT 24.770 4.850 25.060 6.930 ;
        RECT 52.260 6.840 52.610 8.770 ;
        RECT 49.670 6.830 52.610 6.840 ;
        RECT 49.660 6.520 52.610 6.830 ;
        RECT 54.430 6.840 54.780 8.770 ;
        RECT 55.400 8.580 61.450 8.770 ;
        RECT 55.400 8.550 58.610 8.580 ;
        RECT 58.240 8.320 58.610 8.550 ;
        RECT 62.070 8.320 62.420 8.770 ;
        RECT 64.240 8.320 64.590 8.770 ;
        RECT 65.210 8.580 68.370 8.770 ;
        RECT 68.050 8.320 68.370 8.580 ;
        RECT 69.980 8.320 70.330 8.770 ;
        RECT 70.950 8.560 74.110 8.770 ;
        RECT 94.990 8.750 95.550 8.770 ;
        RECT 73.790 8.320 74.110 8.560 ;
        RECT 57.370 7.860 94.450 8.320 ;
        RECT 57.440 7.760 57.960 7.860 ;
        RECT 58.240 7.540 58.610 7.860 ;
        RECT 58.240 7.510 61.450 7.540 ;
        RECT 55.400 7.410 61.450 7.510 ;
        RECT 62.070 7.410 62.420 7.860 ;
        RECT 64.240 7.410 64.590 7.860 ;
        RECT 68.050 7.540 68.370 7.860 ;
        RECT 65.210 7.410 68.370 7.540 ;
        RECT 69.980 7.410 70.330 7.860 ;
        RECT 73.790 7.520 74.110 7.860 ;
        RECT 93.800 7.800 94.360 7.860 ;
        RECT 70.950 7.410 74.110 7.520 ;
        RECT 55.400 7.220 93.360 7.410 ;
        RECT 55.400 7.190 58.560 7.220 ;
        RECT 55.430 7.180 55.740 7.190 ;
        RECT 56.530 7.180 56.840 7.190 ;
        RECT 57.630 7.180 57.940 7.190 ;
        RECT 58.800 6.950 93.360 7.220 ;
        RECT 58.050 6.890 58.650 6.920 ;
        RECT 58.800 6.890 59.450 6.950 ;
        RECT 54.430 6.830 57.370 6.840 ;
        RECT 54.430 6.520 57.380 6.830 ;
        RECT 49.660 6.510 52.380 6.520 ;
        RECT 54.660 6.510 57.380 6.520 ;
        RECT 49.660 6.500 49.970 6.510 ;
        RECT 50.750 6.500 51.060 6.510 ;
        RECT 55.980 6.500 56.290 6.510 ;
        RECT 57.070 6.500 57.380 6.510 ;
        RECT 58.050 6.820 59.450 6.890 ;
        RECT 62.070 6.870 62.420 6.950 ;
        RECT 59.480 6.860 62.420 6.870 ;
        RECT 58.050 6.100 58.800 6.820 ;
        RECT 59.470 6.550 62.420 6.860 ;
        RECT 64.240 6.870 64.590 6.950 ;
        RECT 64.240 6.860 67.180 6.870 ;
        RECT 64.240 6.550 67.190 6.860 ;
        RECT 59.470 6.540 62.190 6.550 ;
        RECT 64.470 6.540 67.190 6.550 ;
        RECT 59.470 6.530 59.780 6.540 ;
        RECT 60.560 6.530 60.870 6.540 ;
        RECT 65.790 6.530 66.100 6.540 ;
        RECT 66.880 6.530 67.190 6.540 ;
        RECT 58.190 6.070 58.800 6.100 ;
        RECT 67.250 6.470 67.770 6.490 ;
        RECT 68.010 6.470 68.610 6.920 ;
        RECT 69.980 6.850 70.330 6.950 ;
        RECT 92.670 6.930 93.230 6.950 ;
        RECT 69.980 6.840 72.920 6.850 ;
        RECT 69.980 6.530 72.930 6.840 ;
        RECT 70.210 6.520 72.930 6.530 ;
        RECT 71.530 6.510 71.840 6.520 ;
        RECT 72.620 6.510 72.930 6.520 ;
        RECT 73.750 6.470 74.350 6.900 ;
        RECT 91.740 6.470 92.300 6.480 ;
        RECT 67.250 6.010 92.390 6.470 ;
        RECT 67.250 5.960 67.780 6.010 ;
        RECT 67.250 5.910 67.770 5.960 ;
        RECT 41.190 4.850 41.510 4.870 ;
        RECT 97.190 4.850 98.350 4.880 ;
        RECT 24.580 3.730 98.350 4.850 ;
        RECT 41.190 3.710 41.510 3.730 ;
        RECT 52.560 3.650 54.480 3.730 ;
        RECT 62.370 3.620 64.300 3.730 ;
        RECT 97.190 3.700 98.350 3.730 ;
        RECT 101.030 1.550 101.230 1.560 ;
        RECT 104.750 1.550 105.070 1.600 ;
        RECT 101.030 1.400 105.070 1.550 ;
        RECT 4.110 0.400 4.610 0.510 ;
        RECT 73.080 0.430 73.470 0.440 ;
        RECT 73.070 0.400 73.470 0.430 ;
        RECT 4.110 0.120 73.470 0.400 ;
        RECT 4.110 0.040 4.610 0.120 ;
        RECT 73.070 0.100 73.470 0.120 ;
        RECT 73.080 0.090 73.470 0.100 ;
        RECT 100.350 -0.690 100.780 -0.670 ;
        RECT 81.850 -0.720 83.810 -0.690 ;
        RECT 100.330 -0.720 100.790 -0.690 ;
        RECT 81.850 -1.070 100.790 -0.720 ;
        RECT 81.850 -7.170 83.810 -1.070 ;
        RECT 100.330 -1.090 100.790 -1.070 ;
        RECT 100.350 -1.100 100.780 -1.090 ;
        RECT 101.030 -1.510 101.230 1.400 ;
        RECT 104.750 1.280 105.070 1.400 ;
        RECT 102.000 -0.010 104.770 0.000 ;
        RECT 102.000 -0.200 105.070 -0.010 ;
        RECT 101.250 -1.500 101.680 -1.480 ;
        RECT 101.240 -1.510 101.690 -1.500 ;
        RECT 85.780 -1.890 101.690 -1.510 ;
        RECT 81.820 -7.820 83.850 -7.170 ;
        RECT 85.780 -7.190 87.740 -1.890 ;
        RECT 99.880 -2.050 100.140 -1.890 ;
        RECT 99.910 -2.330 100.110 -2.050 ;
        RECT 101.030 -2.330 101.230 -1.890 ;
        RECT 101.250 -1.910 101.680 -1.890 ;
        RECT 102.000 -2.320 102.210 -0.200 ;
        RECT 104.750 -0.330 105.070 -0.200 ;
        RECT 103.780 -1.660 104.090 -1.630 ;
        RECT 104.740 -1.660 105.060 -1.620 ;
        RECT 103.780 -1.910 105.060 -1.660 ;
        RECT 102.000 -2.330 102.620 -2.320 ;
        RECT 89.930 -2.710 102.620 -2.330 ;
        RECT 89.930 -7.170 91.910 -2.710 ;
        RECT 99.910 -3.120 100.110 -2.710 ;
        RECT 101.030 -3.120 101.230 -2.710 ;
        RECT 102.000 -3.120 102.210 -2.710 ;
        RECT 103.010 -3.120 103.430 -3.090 ;
        RECT 94.040 -3.500 103.430 -3.120 ;
        RECT 85.770 -7.840 87.800 -7.190 ;
        RECT 89.890 -7.820 91.920 -7.170 ;
        RECT 94.040 -7.200 96.020 -3.500 ;
        RECT 99.910 -6.290 100.110 -3.500 ;
        RECT 101.030 -6.290 101.230 -3.500 ;
        RECT 102.000 -6.290 102.210 -3.500 ;
        RECT 103.010 -3.530 103.430 -3.500 ;
        RECT 103.780 -6.290 104.080 -1.910 ;
        RECT 104.740 -1.940 105.060 -1.910 ;
        RECT 104.740 -3.260 105.060 -3.240 ;
        RECT 104.740 -3.560 105.090 -3.260 ;
        RECT 104.900 -4.850 105.090 -3.560 ;
        RECT 104.740 -5.170 105.090 -4.850 ;
        RECT 104.900 -6.290 105.090 -5.170 ;
        RECT 99.110 -6.490 105.350 -6.290 ;
        RECT 99.110 -7.170 99.310 -6.490 ;
        RECT 99.910 -7.170 100.110 -6.490 ;
        RECT 94.030 -7.850 96.060 -7.200 ;
        RECT 98.020 -7.820 100.110 -7.170 ;
        RECT 99.910 -10.310 100.110 -7.820 ;
        RECT 101.030 -10.170 101.230 -6.490 ;
        RECT 101.020 -10.310 101.230 -10.170 ;
        RECT 102.000 -7.170 102.210 -6.490 ;
        RECT 103.780 -6.610 104.080 -6.490 ;
        RECT 104.370 -6.610 104.690 -6.490 ;
        RECT 103.780 -6.700 104.690 -6.610 ;
        RECT 104.900 -6.700 105.090 -6.490 ;
        RECT 106.270 -6.700 106.470 -6.290 ;
        RECT 103.780 -6.900 106.470 -6.700 ;
        RECT 103.780 -7.170 104.240 -6.900 ;
        RECT 102.000 -7.470 104.240 -7.170 ;
        RECT 102.000 -7.820 104.080 -7.470 ;
        RECT 102.000 -10.310 102.210 -7.820 ;
        RECT 103.780 -8.250 104.080 -7.820 ;
        RECT 104.900 -8.050 105.090 -6.900 ;
        RECT 103.780 -8.410 104.140 -8.250 ;
        RECT 104.750 -8.370 105.090 -8.050 ;
        RECT 103.430 -9.850 103.750 -9.780 ;
        RECT 103.930 -9.850 104.140 -8.410 ;
        RECT 104.900 -9.640 105.090 -8.370 ;
        RECT 103.430 -10.050 104.140 -9.850 ;
        RECT 104.740 -9.960 105.090 -9.640 ;
        RECT 103.430 -10.100 103.750 -10.050 ;
        RECT 103.930 -10.310 104.140 -10.050 ;
        RECT 104.900 -10.160 105.090 -9.960 ;
        RECT 104.880 -10.310 105.090 -10.160 ;
      LAYER via2 ;
        RECT 79.480 47.310 79.800 47.630 ;
        RECT 80.510 47.300 80.830 47.620 ;
    END
  END DIG25
  PIN DIG16
    PORT
      LAYER met2 ;
        RECT 39.510 48.650 39.900 48.740 ;
        RECT 39.510 48.480 41.240 48.650 ;
        RECT 39.490 -0.230 39.910 -0.220 ;
        RECT 39.490 -0.480 79.760 -0.230 ;
        RECT 39.490 -0.560 79.770 -0.480 ;
        RECT 39.490 -0.570 39.910 -0.560 ;
        RECT 73.730 -0.580 79.770 -0.560 ;
        RECT 77.830 -1.080 79.770 -0.580 ;
        RECT 77.830 -7.150 79.760 -1.080 ;
        RECT 77.740 -7.930 79.770 -7.150 ;
    END
  END DIG16
  PIN DIG15
    PORT
      LAYER met2 ;
        RECT 38.910 47.110 39.240 47.120 ;
        RECT 38.890 47.010 39.260 47.110 ;
        RECT 38.890 46.840 41.240 47.010 ;
        RECT 38.890 46.730 39.260 46.840 ;
        RECT 38.890 -0.850 39.270 -0.840 ;
        RECT 38.890 -1.180 75.690 -0.850 ;
        RECT 38.890 -1.190 39.270 -1.180 ;
        RECT 69.620 -1.190 75.690 -1.180 ;
        RECT 73.730 -1.510 75.690 -1.190 ;
        RECT 73.730 -7.170 75.680 -1.510 ;
        RECT 73.670 -7.820 75.700 -7.170 ;
    END
  END DIG15
  PIN DIG14
    PORT
      LAYER met2 ;
        RECT 38.310 45.530 38.700 45.630 ;
        RECT 38.310 45.360 41.240 45.530 ;
        RECT 38.310 45.260 38.700 45.360 ;
        RECT 38.250 -1.480 38.670 -1.470 ;
        RECT 38.250 -1.810 71.610 -1.480 ;
        RECT 38.250 -1.820 38.670 -1.810 ;
        RECT 69.620 -7.170 71.610 -1.810 ;
        RECT 69.620 -7.820 71.650 -7.170 ;
    END
  END DIG14
  PIN DIG13
    PORT
      LAYER met2 ;
        RECT 37.670 43.930 38.060 44.020 ;
        RECT 37.670 43.760 41.240 43.930 ;
        RECT 37.670 43.670 38.060 43.760 ;
        RECT 37.660 -2.120 38.060 -2.100 ;
        RECT 37.660 -2.450 67.600 -2.120 ;
        RECT 37.660 -2.460 38.060 -2.450 ;
        RECT 65.640 -7.170 67.590 -2.450 ;
        RECT 65.590 -7.820 67.620 -7.170 ;
    END
  END DIG13
  PIN DIG12
    PORT
      LAYER met2 ;
        RECT 37.030 43.360 37.420 43.470 ;
        RECT 37.030 43.190 41.240 43.360 ;
        RECT 37.030 43.090 37.420 43.190 ;
        RECT 37.000 -2.790 37.410 -2.780 ;
        RECT 36.990 -3.120 63.510 -2.790 ;
        RECT 37.000 -3.140 37.410 -3.120 ;
        RECT 61.600 -7.190 63.510 -3.120 ;
        RECT 61.520 -7.840 63.550 -7.190 ;
    END
  END DIG12
  PIN DIG11
    PORT
      LAYER met2 ;
        RECT 36.420 41.790 36.810 41.890 ;
        RECT 36.420 41.620 41.240 41.790 ;
        RECT 36.420 41.520 36.810 41.620 ;
        RECT 36.420 -3.410 36.830 -3.400 ;
        RECT 36.420 -3.430 59.490 -3.410 ;
        RECT 36.420 -3.740 59.500 -3.430 ;
        RECT 36.420 -3.750 36.830 -3.740 ;
        RECT 57.500 -7.120 59.500 -3.740 ;
        RECT 57.470 -7.820 59.500 -7.120 ;
    END
  END DIG11
  PIN DIG10
    PORT
      LAYER met2 ;
        RECT 35.790 40.260 36.210 40.350 ;
        RECT 35.790 40.090 41.240 40.260 ;
        RECT 35.790 40.000 36.210 40.090 ;
        RECT 35.820 -4.060 36.210 -4.050 ;
        RECT 35.820 -4.380 55.510 -4.060 ;
        RECT 35.920 -4.390 55.510 -4.380 ;
        RECT 53.520 -7.100 55.510 -4.390 ;
        RECT 53.510 -7.850 55.540 -7.100 ;
    END
  END DIG10
  PIN DIG09
    PORT
      LAYER met2 ;
        RECT 35.230 38.690 35.620 38.780 ;
        RECT 35.230 38.520 41.240 38.690 ;
        RECT 35.230 38.430 35.620 38.520 ;
        RECT 35.240 -4.670 35.630 -4.620 ;
        RECT 35.240 -4.950 51.600 -4.670 ;
        RECT 35.500 -5.000 51.600 -4.950 ;
        RECT 49.530 -7.820 51.560 -5.000 ;
    END
  END DIG09
  PIN DIG08
    PORT
      LAYER met2 ;
        RECT 34.620 33.220 34.990 33.340 ;
        RECT 34.620 33.050 40.940 33.220 ;
        RECT 34.620 32.940 34.990 33.050 ;
        RECT 34.660 -5.640 47.400 -5.310 ;
        RECT 45.350 -7.170 47.380 -5.640 ;
        RECT 45.350 -7.180 47.370 -7.170 ;
        RECT 45.350 -7.230 47.390 -7.180 ;
        RECT 45.360 -7.840 47.390 -7.230 ;
    END
  END DIG08
  PIN DIG07
    PORT
      LAYER met2 ;
        RECT 33.980 31.630 34.370 31.720 ;
        RECT 33.980 31.460 40.940 31.630 ;
        RECT 33.980 31.370 34.370 31.460 ;
        RECT 41.270 -5.940 43.290 -5.920 ;
        RECT 34.110 -5.950 43.290 -5.940 ;
        RECT 34.010 -6.270 43.290 -5.950 ;
        RECT 34.010 -6.280 34.400 -6.270 ;
        RECT 41.250 -7.150 43.290 -6.270 ;
        RECT 41.250 -7.160 43.270 -7.150 ;
        RECT 41.250 -7.230 43.300 -7.160 ;
        RECT 41.270 -7.820 43.300 -7.230 ;
    END
  END DIG07
  PIN DIG06
    PORT
      LAYER met2 ;
        RECT 33.360 30.080 33.750 30.160 ;
        RECT 33.360 29.910 40.940 30.080 ;
        RECT 33.360 29.830 33.750 29.910 ;
        RECT 33.370 -6.930 39.350 -6.590 ;
        RECT 37.340 -7.180 39.350 -6.930 ;
        RECT 39.010 -7.190 39.350 -7.180 ;
        RECT 37.310 -7.370 39.350 -7.190 ;
        RECT 37.310 -7.850 39.340 -7.370 ;
    END
  END DIG06
  PIN DIG05
    PORT
      LAYER met2 ;
        RECT 32.750 28.600 33.170 28.690 ;
        RECT 32.750 28.430 40.940 28.600 ;
        RECT 32.750 28.330 33.170 28.430 ;
        RECT 32.760 -7.180 33.310 -7.160 ;
        RECT 32.760 -7.610 35.310 -7.180 ;
        RECT 33.280 -7.840 35.310 -7.610 ;
    END
  END DIG05
  PIN DIG04
    PORT
      LAYER met2 ;
        RECT 32.110 23.430 32.520 23.530 ;
        RECT 32.110 23.260 40.940 23.430 ;
        RECT 32.110 23.170 32.520 23.260 ;
        RECT 31.260 -7.160 31.910 -7.150 ;
        RECT 29.230 -7.790 31.910 -7.160 ;
        RECT 29.230 -7.820 31.260 -7.790 ;
    END
  END DIG04
  PIN DIG03
    PORT
      LAYER met2 ;
        RECT 31.450 21.860 31.840 21.970 ;
        RECT 31.450 21.690 40.940 21.860 ;
        RECT 31.450 21.590 31.840 21.690 ;
        RECT 31.430 -6.530 31.920 -6.330 ;
        RECT 25.820 -6.550 31.920 -6.530 ;
        RECT 25.250 -6.830 31.920 -6.550 ;
        RECT 25.250 -6.930 31.830 -6.830 ;
        RECT 25.250 -7.160 27.230 -6.930 ;
        RECT 25.230 -7.820 27.260 -7.160 ;
    END
  END DIG03
  PIN DIG02
    PORT
      LAYER met2 ;
        RECT 30.840 20.320 31.210 20.330 ;
        RECT 30.840 20.150 40.940 20.320 ;
        RECT 30.840 19.940 31.210 20.150 ;
        RECT 30.750 -5.720 31.290 -5.650 ;
        RECT 21.320 -6.150 31.290 -5.720 ;
        RECT 21.320 -7.160 23.300 -6.150 ;
        RECT 21.270 -7.820 23.300 -7.160 ;
    END
  END DIG02
  PIN DIG01
    PORT
      LAYER met2 ;
        RECT 30.150 18.780 30.540 18.880 ;
        RECT 30.150 18.610 40.940 18.780 ;
        RECT 30.150 18.510 30.540 18.610 ;
        RECT 30.100 -4.880 30.640 -4.840 ;
        RECT 17.270 -4.920 30.640 -4.880 ;
        RECT 17.220 -5.310 30.640 -4.920 ;
        RECT 17.220 -7.190 19.230 -5.310 ;
        RECT 30.100 -5.340 30.640 -5.310 ;
        RECT 17.200 -7.850 19.230 -7.190 ;
    END
  END DIG01
  PIN OUTPUTTA1    
    ANTENNAGATEAREA 0.477400 ;
    PORT
      LAYER met2 ;
        RECT 8.730 57.790 9.040 58.020 ;
        RECT 5.640 57.690 9.040 57.790 ;
        RECT 5.640 57.560 9.020 57.690 ;
        RECT 5.640 57.530 5.960 57.560 ;
        RECT 115.050 55.250 115.820 55.400 ;
        RECT 5.560 54.830 115.820 55.250 ;
        RECT 115.050 54.690 115.820 54.830 ;
        RECT 114.860 35.490 115.640 35.640 ;
        RECT 117.600 35.490 118.500 36.410 ;
        RECT 114.860 35.020 118.500 35.490 ;
        RECT 114.860 34.870 115.640 35.020 ;
        RECT 117.600 34.320 118.500 35.020 ;
    END
  END OUTPUTTA1    
  PIN DRAINOUT
    ANTENNAGATEAREA 4.652100 ;
    ANTENNADIFFAREA 30.025099 ;
    PORT
      LAYER met2 ;
        RECT 44.420 56.610 44.920 56.630 ;
        RECT 50.160 56.610 50.600 56.660 ;
        RECT 64.530 56.610 65.030 56.630 ;
        RECT 44.420 56.190 70.930 56.610 ;
        RECT 44.570 56.170 70.930 56.190 ;
        RECT 50.160 56.160 50.600 56.170 ;
        RECT 70.330 56.150 70.830 56.170 ;
        RECT 41.670 53.400 41.970 53.460 ;
        RECT 82.990 53.400 83.290 53.430 ;
        RECT 41.670 53.170 83.360 53.400 ;
        RECT 41.670 53.140 41.970 53.170 ;
        RECT 82.990 53.090 83.290 53.170 ;
        RECT 84.770 48.740 85.090 48.750 ;
        RECT 84.530 48.730 85.090 48.740 ;
        RECT 110.760 48.730 111.070 48.740 ;
        RECT 82.360 48.650 93.880 48.730 ;
        RECT 101.710 48.650 113.240 48.730 ;
        RECT 117.640 48.650 118.500 50.630 ;
        RECT 82.360 48.550 118.500 48.650 ;
        RECT 84.530 48.410 84.840 48.550 ;
        RECT 89.290 48.530 118.500 48.550 ;
        RECT 89.290 48.280 118.390 48.530 ;
        RECT 89.290 48.250 89.700 48.280 ;
        RECT 110.910 47.710 111.220 47.780 ;
        RECT 83.200 47.630 83.670 47.690 ;
        RECT 108.100 47.640 108.390 47.650 ;
        RECT 108.100 47.630 108.400 47.640 ;
        RECT 110.910 47.630 113.240 47.710 ;
        RECT 118.630 47.630 119.080 47.650 ;
        RECT 83.200 47.200 119.090 47.630 ;
        RECT 84.140 47.190 84.450 47.200 ;
        RECT 108.100 47.190 108.400 47.200 ;
        RECT 84.140 47.000 93.880 47.190 ;
        RECT 108.100 47.170 108.390 47.190 ;
        RECT 84.140 46.880 84.450 47.000 ;
        RECT 83.420 46.310 83.740 46.340 ;
        RECT 83.420 46.080 93.880 46.310 ;
        RECT 81.730 41.740 82.050 42.000 ;
        RECT 81.770 41.720 82.950 41.740 ;
        RECT 81.770 41.460 82.990 41.720 ;
        RECT 81.770 41.400 82.950 41.460 ;
        RECT 81.730 41.390 82.950 41.400 ;
        RECT 81.730 41.140 82.050 41.390 ;
        RECT 79.400 40.760 79.960 40.780 ;
        RECT 80.400 40.760 80.710 40.770 ;
        RECT 79.400 40.510 80.710 40.760 ;
        RECT 79.400 40.240 79.960 40.510 ;
        RECT 80.400 40.440 80.710 40.510 ;
        RECT 81.370 40.440 81.680 40.490 ;
        RECT 83.620 40.440 83.930 40.540 ;
        RECT 80.790 40.320 81.100 40.390 ;
        RECT 81.370 40.320 83.930 40.440 ;
        RECT 80.790 40.210 83.930 40.320 ;
        RECT 80.790 40.110 83.120 40.210 ;
        RECT 80.790 40.060 81.100 40.110 ;
        RECT 80.550 39.900 80.860 39.940 ;
        RECT 80.370 39.760 81.090 39.900 ;
        RECT 81.320 39.760 81.630 39.840 ;
        RECT 80.370 39.650 81.630 39.760 ;
        RECT 80.550 39.610 81.630 39.650 ;
        RECT 80.820 39.550 81.630 39.610 ;
        RECT 80.820 39.540 81.090 39.550 ;
        RECT 81.320 39.510 81.630 39.550 ;
        RECT 79.430 39.260 79.740 39.400 ;
        RECT 65.550 39.220 75.690 39.250 ;
        RECT 79.080 39.220 79.740 39.260 ;
        RECT 80.640 39.230 80.950 39.370 ;
        RECT 80.640 39.220 83.120 39.230 ;
        RECT 65.550 39.070 83.120 39.220 ;
        RECT 65.550 39.030 75.690 39.070 ;
        RECT 79.080 39.040 79.430 39.070 ;
        RECT 80.640 39.050 83.120 39.070 ;
        RECT 80.640 39.040 80.950 39.050 ;
        RECT 75.470 37.830 75.690 39.030 ;
        RECT 80.890 38.970 81.090 38.980 ;
        RECT 80.890 38.960 81.110 38.970 ;
        RECT 81.320 38.960 81.630 39.000 ;
        RECT 80.890 38.890 81.630 38.960 ;
        RECT 80.600 38.870 81.630 38.890 ;
        RECT 80.550 38.750 81.630 38.870 ;
        RECT 80.550 38.630 81.110 38.750 ;
        RECT 81.320 38.670 81.630 38.750 ;
        RECT 80.550 38.620 81.020 38.630 ;
        RECT 75.440 37.790 75.690 37.830 ;
        RECT 75.440 37.150 75.700 37.790 ;
        RECT 75.440 36.940 79.570 37.150 ;
        RECT 79.360 36.800 79.570 36.940 ;
        RECT 81.320 36.800 81.630 36.880 ;
        RECT 79.360 36.590 81.630 36.800 ;
        RECT 81.320 36.550 81.630 36.590 ;
        RECT 70.380 35.080 70.700 35.090 ;
        RECT 80.820 35.080 81.150 35.220 ;
        RECT 69.840 34.930 70.150 34.940 ;
        RECT 70.380 34.930 81.150 35.080 ;
        RECT 67.680 34.920 81.150 34.930 ;
        RECT 67.680 34.750 77.760 34.920 ;
        RECT 69.840 34.610 70.150 34.750 ;
        RECT 69.840 33.350 70.150 33.370 ;
        RECT 70.520 33.350 73.370 33.430 ;
        RECT 87.410 33.350 90.240 33.430 ;
        RECT 90.610 33.350 90.920 33.370 ;
        RECT 67.680 33.330 77.740 33.350 ;
        RECT 83.020 33.330 93.080 33.350 ;
        RECT 67.680 33.180 93.080 33.330 ;
        RECT 67.680 33.170 70.240 33.180 ;
        RECT 69.840 33.040 70.150 33.170 ;
        RECT 70.520 33.130 70.940 33.180 ;
        RECT 72.930 33.150 87.610 33.180 ;
        RECT 89.920 33.130 90.240 33.180 ;
        RECT 90.520 33.170 93.080 33.180 ;
        RECT 90.610 33.040 90.920 33.170 ;
        RECT 70.750 32.800 71.070 32.880 ;
        RECT 74.680 32.800 75.000 32.810 ;
        RECT 70.750 32.620 75.000 32.800 ;
        RECT 70.750 32.560 71.070 32.620 ;
        RECT 74.680 32.550 75.000 32.620 ;
        RECT 85.760 32.800 86.080 32.810 ;
        RECT 89.690 32.800 90.010 32.880 ;
        RECT 85.760 32.620 90.010 32.800 ;
        RECT 85.760 32.550 86.080 32.620 ;
        RECT 89.690 32.560 90.010 32.620 ;
        RECT 57.140 26.540 57.450 26.560 ;
        RECT 51.630 26.390 51.940 26.410 ;
        RECT 54.980 26.390 65.060 26.540 ;
        RECT 89.270 26.390 89.720 26.420 ;
        RECT 51.630 25.980 89.720 26.390 ;
        RECT 51.630 25.960 51.940 25.980 ;
        RECT 89.270 25.960 89.720 25.980 ;
      LAYER via2 ;
        RECT 79.520 40.340 79.850 40.690 ;
    END
  END DRAINOUT
  PIN ROWTERM2
    PORT
      LAYER met2 ;
        RECT 88.410 53.720 88.830 53.740 ;
        RECT 117.640 53.720 118.500 55.020 ;
        RECT 88.410 53.350 118.500 53.720 ;
        RECT 88.410 53.330 88.830 53.350 ;
        RECT 117.640 52.920 118.500 53.350 ;
        RECT 88.350 31.500 88.790 31.620 ;
        RECT 77.590 31.320 88.790 31.500 ;
        RECT 88.350 31.220 88.790 31.320 ;
    END
  END ROWTERM2
  PIN COLUMN2
    ANTENNADIFFAREA 5.542100 ;
    PORT
      LAYER nwell ;
        RECT 87.400 46.840 90.120 48.490 ;
        RECT 87.400 46.800 90.110 46.840 ;
        RECT 87.400 45.470 90.110 45.510 ;
        RECT 87.400 45.410 90.120 45.470 ;
        RECT 86.310 45.400 90.120 45.410 ;
        RECT 87.400 43.820 90.120 45.400 ;
        RECT 86.760 31.240 88.990 37.290 ;
      LAYER met2 ;
        RECT 87.630 58.430 88.070 58.450 ;
        RECT 117.670 58.430 118.530 59.110 ;
        RECT 87.630 58.060 118.530 58.430 ;
        RECT 87.630 58.040 88.070 58.060 ;
        RECT 117.670 57.010 118.530 58.060 ;
        RECT 69.840 33.780 70.150 33.920 ;
        RECT 87.610 33.870 88.040 33.950 ;
        RECT 67.680 33.770 70.150 33.780 ;
        RECT 76.350 33.770 88.040 33.870 ;
        RECT 90.610 33.780 90.920 33.920 ;
        RECT 90.610 33.770 93.080 33.780 ;
        RECT 67.680 33.610 93.080 33.770 ;
        RECT 67.680 33.600 77.740 33.610 ;
        RECT 83.020 33.600 93.080 33.610 ;
        RECT 69.840 33.590 70.150 33.600 ;
        RECT 87.610 33.540 88.040 33.600 ;
        RECT 90.610 33.590 90.920 33.600 ;
    END
  END COLUMN2
  PIN COLUMN1
    ANTENNAGATEAREA 0.790000 ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 86.800 61.890 87.260 61.910 ;
        RECT 117.670 61.890 118.530 63.240 ;
        RECT 86.800 61.520 118.530 61.890 ;
        RECT 86.800 61.500 87.260 61.520 ;
        RECT 117.670 61.140 118.530 61.520 ;
        RECT 84.130 45.330 84.440 45.520 ;
        RECT 86.510 45.330 86.830 45.390 ;
        RECT 84.130 45.270 93.880 45.330 ;
        RECT 108.780 45.270 109.100 45.390 ;
        RECT 84.130 45.190 109.100 45.270 ;
        RECT 84.160 45.140 109.100 45.190 ;
        RECT 86.510 45.090 109.100 45.140 ;
        RECT 59.010 34.470 59.330 34.480 ;
        RECT 86.820 34.470 87.280 34.540 ;
        RECT 59.010 34.190 87.280 34.470 ;
        RECT 59.010 34.140 59.330 34.190 ;
        RECT 86.820 34.130 87.280 34.190 ;
    END
  END COLUMN1
  PIN GATE2
    ANTENNADIFFAREA 1.847500 ;
    PORT
      LAYER met1 ;
        RECT 102.730 62.870 105.920 63.990 ;
        RECT 103.820 50.670 105.100 62.870 ;
        RECT 103.810 49.330 105.100 50.670 ;
        RECT 103.820 48.840 105.100 49.330 ;
        RECT 104.540 46.370 104.770 48.840 ;
        RECT 104.270 45.890 104.770 46.370 ;
        RECT 104.370 43.180 104.770 45.890 ;
        RECT 104.370 15.900 104.600 43.180 ;
        RECT 104.370 15.670 104.610 15.900 ;
        RECT 104.370 9.860 104.600 15.670 ;
      LAYER via ;
        RECT 103.810 49.360 105.090 50.640 ;
        RECT 104.300 45.920 104.560 46.340 ;
    END
  END GATE2
  PIN DRAININJECT
    ANTENNADIFFAREA 0.105300 ;
    PORT
      LAYER met2 ;
        RECT 47.180 60.000 47.630 60.020 ;
        RECT 47.170 59.940 47.650 60.000 ;
        RECT 24.780 59.800 47.650 59.940 ;
        RECT 24.760 59.640 47.650 59.800 ;
        RECT 24.760 59.480 25.080 59.640 ;
        RECT 47.170 59.580 47.650 59.640 ;
        RECT 47.180 59.560 47.630 59.580 ;
        RECT 24.760 59.470 25.070 59.480 ;
    END
  END DRAININJECT
  PIN VTUN
    ANTENNADIFFAREA 0.604400 ;
    PORT
      LAYER nwell ;
        RECT 33.720 59.960 35.940 61.650 ;
      LAYER met2 ;
        RECT 43.330 59.240 43.780 59.260 ;
        RECT 43.320 59.230 43.800 59.240 ;
        RECT 66.940 59.230 68.360 59.270 ;
        RECT 43.320 58.830 68.410 59.230 ;
        RECT 43.320 58.820 43.800 58.830 ;
        RECT 43.330 58.800 43.780 58.820 ;
        RECT 66.940 58.790 68.360 58.830 ;
    END
  END VTUN
  PIN CHAROUTPUT
    ANTENNADIFFAREA 0.359600 ;
    PORT
      LAYER met2 ;
        RECT 2.950 58.270 3.630 59.150 ;
        RECT 2.950 58.240 6.610 58.270 ;
        RECT 2.950 57.980 6.910 58.240 ;
        RECT 2.950 57.950 6.610 57.980 ;
        RECT 2.950 56.830 3.630 57.950 ;
    END
  END CHAROUTPUT
  PIN LARGECAPACITOR
    ANTENNADIFFAREA 6.082200 ;
    PORT
      LAYER nwell ;
        RECT 11.700 57.080 21.390 61.680 ;
        RECT 11.100 55.690 21.390 57.080 ;
      LAYER met2 ;
        RECT 2.500 54.010 3.180 54.680 ;
        RECT 11.420 54.010 11.890 54.030 ;
        RECT 2.500 53.430 11.890 54.010 ;
        RECT 2.500 53.190 3.220 53.430 ;
        RECT 11.420 53.410 11.890 53.430 ;
        RECT 2.500 52.360 3.180 53.190 ;
    END
  END LARGECAPACITOR
  PIN DRAIN6N
    PORT
      LAYER met2 ;
        RECT 13.790 9.600 14.160 9.610 ;
        RECT 2.900 8.780 4.170 9.480 ;
        RECT 12.470 9.220 15.000 9.600 ;
        RECT 12.470 8.780 12.850 9.220 ;
        RECT 13.790 9.200 14.160 9.220 ;
        RECT 2.900 8.400 12.850 8.780 ;
        RECT 2.900 7.600 4.170 8.400 ;
    END
  END DRAIN6N
  PIN DRAIN6P
    PORT
      LAYER met2 ;
        RECT 2.900 3.550 4.170 4.460 ;
        RECT 2.900 3.170 12.870 3.550 ;
        RECT 2.900 2.580 4.170 3.170 ;
        RECT 12.490 2.320 12.870 3.170 ;
        RECT 13.790 2.320 14.160 2.330 ;
        RECT 12.490 1.940 15.210 2.320 ;
        RECT 13.790 1.920 14.160 1.940 ;
    END
  END DRAIN6P
  PIN DRAIN5P
    PORT
      LAYER met2 ;
        RECT 12.060 19.230 12.470 19.250 ;
        RECT 13.830 19.230 15.820 19.250 ;
        RECT 12.060 19.190 15.820 19.230 ;
        RECT 18.800 19.190 19.110 19.240 ;
        RECT 12.060 18.970 19.110 19.190 ;
        RECT 12.060 18.860 14.210 18.970 ;
        RECT 18.800 18.910 19.110 18.970 ;
        RECT 12.060 18.840 12.470 18.860 ;
        RECT 13.830 18.840 14.200 18.860 ;
        RECT 2.840 12.990 4.110 13.770 ;
        RECT 12.070 12.990 12.480 13.010 ;
        RECT 2.840 12.620 12.480 12.990 ;
        RECT 2.840 11.890 4.110 12.620 ;
        RECT 12.070 12.600 12.480 12.620 ;
    END
  END DRAIN5P
  PIN DARIN4P
    ANTENNADIFFAREA 0.727900 ;
    PORT
      LAYER met2 ;
        RECT 2.900 22.240 4.170 23.010 ;
        RECT 2.900 21.870 8.890 22.240 ;
        RECT 2.900 21.130 4.170 21.870 ;
        RECT 8.520 20.210 8.890 21.870 ;
        RECT 8.520 20.030 14.470 20.210 ;
        RECT 8.520 19.960 14.540 20.030 ;
        RECT 15.930 19.960 17.200 19.970 ;
        RECT 17.630 19.960 17.940 20.020 ;
        RECT 8.520 19.840 17.940 19.960 ;
        RECT 13.830 19.800 17.940 19.840 ;
        RECT 14.190 19.750 17.940 19.800 ;
        RECT 17.630 19.690 17.940 19.750 ;
    END
  END DARIN4P
  PIN DRAIN5N
    ANTENNADIFFAREA 0.688800 ;
    PORT
      LAYER met2 ;
        RECT 6.830 23.890 7.600 24.080 ;
        RECT 13.830 23.890 14.220 23.910 ;
        RECT 6.830 23.850 14.220 23.890 ;
        RECT 17.600 23.850 17.910 23.900 ;
        RECT 6.830 23.640 17.910 23.850 ;
        RECT 6.830 23.520 14.210 23.640 ;
        RECT 17.600 23.570 17.910 23.640 ;
        RECT 6.830 23.340 7.600 23.520 ;
        RECT 13.830 23.500 14.200 23.520 ;
        RECT 2.900 18.100 4.170 18.920 ;
        RECT 6.830 18.100 7.630 18.240 ;
        RECT 2.900 17.600 7.630 18.100 ;
        RECT 2.900 17.040 4.170 17.600 ;
        RECT 6.830 17.470 7.630 17.600 ;
    END
  END DRAIN5N
  PIN DRAIN4N
    ANTENNADIFFAREA 0.688800 ;
    PORT
      LAYER met2 ;
        RECT 2.840 26.270 4.110 27.110 ;
        RECT 2.840 25.900 12.540 26.270 ;
        RECT 2.840 25.230 4.110 25.900 ;
        RECT 12.170 24.550 12.540 25.900 ;
        RECT 12.170 24.540 14.200 24.550 ;
        RECT 12.170 24.360 14.420 24.540 ;
        RECT 12.170 24.300 15.820 24.360 ;
        RECT 18.820 24.300 19.130 24.340 ;
        RECT 12.170 24.180 19.130 24.300 ;
        RECT 13.830 24.140 19.130 24.180 ;
        RECT 14.200 24.080 19.130 24.140 ;
        RECT 18.820 24.010 19.130 24.080 ;
    END
  END DRAIN4N
  PIN DRAIN3P
    ANTENNADIFFAREA 0.109200 ;
    PORT
      LAYER met2 ;
        RECT 19.700 41.980 20.010 42.090 ;
        RECT 13.830 41.790 20.010 41.980 ;
        RECT 2.900 30.420 4.170 31.330 ;
        RECT 13.830 30.420 14.200 41.790 ;
        RECT 19.700 41.760 20.010 41.790 ;
        RECT 2.900 30.050 14.200 30.420 ;
        RECT 2.900 29.450 4.170 30.050 ;
    END
  END DRAIN3P
  PIN DRAIN2P
    ANTENNADIFFAREA 0.218400 ;
    PORT
      LAYER met2 ;
        RECT 19.700 43.900 20.010 44.010 ;
        RECT 12.990 43.880 20.010 43.900 ;
        RECT 12.700 43.710 20.010 43.880 ;
        RECT 12.700 43.530 14.200 43.710 ;
        RECT 19.700 43.680 20.010 43.710 ;
        RECT 12.700 42.940 13.360 43.530 ;
        RECT 13.830 43.490 14.200 43.530 ;
        RECT 19.700 42.940 20.010 43.050 ;
        RECT 12.700 42.750 20.010 42.940 ;
        RECT 12.700 42.570 14.200 42.750 ;
        RECT 19.700 42.720 20.010 42.750 ;
        RECT 12.700 42.560 13.370 42.570 ;
        RECT 12.700 42.520 13.360 42.560 ;
        RECT 13.830 42.530 14.200 42.570 ;
        RECT 2.840 35.260 4.110 36.150 ;
        RECT 12.700 35.260 13.070 42.520 ;
        RECT 2.840 34.890 13.070 35.260 ;
        RECT 2.840 34.270 4.110 34.890 ;
    END
  END DRAIN2P
  PIN DRAIN3N
    ANTENNADIFFAREA 0.325500 ;
    PORT
      LAYER met2 ;
        RECT 13.830 46.970 14.200 46.980 ;
        RECT 12.040 46.740 14.200 46.970 ;
        RECT 19.890 46.740 20.200 46.830 ;
        RECT 12.040 46.610 20.200 46.740 ;
        RECT 12.040 45.910 12.660 46.610 ;
        RECT 13.830 46.570 20.200 46.610 ;
        RECT 19.890 46.500 20.200 46.570 ;
        RECT 13.830 45.910 14.200 45.950 ;
        RECT 11.510 45.820 14.200 45.910 ;
        RECT 19.890 45.820 20.200 45.910 ;
        RECT 11.510 45.650 20.200 45.820 ;
        RECT 11.510 45.540 14.200 45.650 ;
        RECT 19.890 45.580 20.200 45.650 ;
        RECT 11.510 45.430 12.660 45.540 ;
        RECT 11.510 44.980 12.620 45.430 ;
        RECT 13.830 44.980 14.200 45.020 ;
        RECT 11.510 44.900 14.200 44.980 ;
        RECT 19.890 44.900 20.200 44.990 ;
        RECT 11.510 44.730 20.200 44.900 ;
        RECT 11.510 44.610 14.200 44.730 ;
        RECT 19.890 44.660 20.200 44.730 ;
        RECT 11.510 44.570 12.410 44.610 ;
        RECT 2.900 40.020 4.170 40.900 ;
        RECT 11.510 40.020 11.880 44.570 ;
        RECT 2.900 39.650 11.880 40.020 ;
        RECT 2.900 39.020 4.170 39.650 ;
    END
  END DRAIN3N
  PIN SOURCEP
    ANTENNADIFFAREA 0.315900 ;
    PORT
      LAYER met2 ;
        RECT 2.180 48.860 3.450 50.320 ;
        RECT 13.530 48.860 13.830 48.870 ;
        RECT 23.120 48.860 23.410 48.880 ;
        RECT 2.180 48.470 23.440 48.860 ;
        RECT 2.180 48.440 3.450 48.470 ;
        RECT 23.120 48.450 23.410 48.470 ;
        RECT 21.000 43.840 21.310 43.910 ;
        RECT 23.100 43.840 23.420 43.870 ;
        RECT 21.000 43.640 23.520 43.840 ;
        RECT 21.000 43.580 21.310 43.640 ;
        RECT 23.100 43.610 23.420 43.640 ;
        RECT 21.000 42.880 21.310 42.950 ;
        RECT 23.110 42.880 23.430 42.910 ;
        RECT 21.000 42.680 23.520 42.880 ;
        RECT 21.000 42.620 21.310 42.680 ;
        RECT 23.110 42.650 23.430 42.680 ;
        RECT 21.000 41.920 21.310 41.990 ;
        RECT 23.100 41.920 23.420 41.950 ;
        RECT 21.000 41.720 23.520 41.920 ;
        RECT 21.000 41.660 21.310 41.720 ;
        RECT 23.100 41.690 23.420 41.720 ;
        RECT 18.320 19.940 18.630 20.010 ;
        RECT 23.110 19.960 23.400 19.980 ;
        RECT 18.320 19.930 20.460 19.940 ;
        RECT 23.100 19.930 23.420 19.960 ;
        RECT 18.320 19.730 23.420 19.930 ;
        RECT 18.320 19.680 18.630 19.730 ;
        RECT 20.250 19.720 23.420 19.730 ;
        RECT 19.510 19.110 19.820 19.180 ;
        RECT 20.250 19.110 20.460 19.720 ;
        RECT 23.100 19.700 23.420 19.720 ;
        RECT 23.110 19.680 23.400 19.700 ;
        RECT 19.510 18.900 20.460 19.110 ;
        RECT 19.510 18.850 19.820 18.900 ;
        RECT 23.040 1.350 23.350 1.370 ;
        RECT 18.810 1.010 23.350 1.350 ;
        RECT 23.040 0.990 23.350 1.010 ;
    END
  END SOURCEP
  PIN GATE1
    PORT
      LAYER met2 ;
        RECT 59.240 50.710 59.560 50.750 ;
        RECT 74.890 50.710 76.170 50.810 ;
        RECT 59.240 50.500 76.170 50.710 ;
        RECT 59.240 50.470 59.560 50.500 ;
    END
  END GATE1
  PIN VINJ
    ANTENNADIFFAREA 1.921700 ;
    PORT
      LAYER nwell ;
        RECT 6.090 58.170 8.830 61.670 ;
        RECT 22.970 55.670 26.970 61.660 ;
      LAYER met2 ;
        RECT 2.800 60.260 5.280 60.270 ;
        RECT 6.590 60.260 6.910 60.460 ;
        RECT 7.320 60.260 7.630 60.470 ;
        RECT 8.000 60.260 8.320 60.470 ;
        RECT 8.660 60.260 23.310 60.390 ;
        RECT 2.800 60.180 23.310 60.260 ;
        RECT 2.800 60.010 8.800 60.180 ;
        RECT 22.730 60.170 23.480 60.180 ;
        RECT 2.800 59.870 8.660 60.010 ;
        RECT 5.070 59.500 8.660 59.870 ;
        RECT 22.730 59.870 24.350 60.170 ;
        RECT 22.730 59.730 22.970 59.870 ;
        RECT 24.050 59.810 24.350 59.870 ;
        RECT 6.590 59.330 6.910 59.500 ;
        RECT 7.320 59.300 7.630 59.500 ;
        RECT 8.020 59.350 8.340 59.500 ;
        RECT 22.710 59.400 23.020 59.730 ;
        RECT 24.050 59.490 24.380 59.810 ;
        RECT 24.070 59.480 24.380 59.490 ;
    END
    PORT
      LAYER met2 ;
        RECT 2.500 51.860 3.010 51.980 ;
        RECT 2.500 51.570 5.600 51.860 ;
        RECT 3.010 51.560 5.600 51.570 ;
    END
    PORT
      LAYER nwell ;
        RECT 46.950 44.250 49.460 50.490 ;
      LAYER met2 ;
        RECT 48.840 57.620 49.340 57.650 ;
        RECT 54.560 57.620 55.060 57.650 ;
        RECT 48.840 57.210 79.000 57.620 ;
        RECT 48.990 57.180 79.000 57.210 ;
        RECT 56.110 46.140 56.400 46.320 ;
        RECT 54.400 44.100 54.710 44.110 ;
        RECT 56.110 44.100 56.290 46.140 ;
        RECT 52.230 43.920 63.760 44.100 ;
        RECT 54.400 43.780 54.710 43.920 ;
        RECT 54.250 43.080 54.560 43.150 ;
        RECT 52.230 43.070 54.560 43.080 ;
        RECT 56.110 43.070 56.290 43.920 ;
        RECT 61.530 43.070 61.850 43.120 ;
        RECT 63.940 43.070 64.260 43.090 ;
        RECT 52.230 42.930 64.260 43.070 ;
        RECT 52.230 42.880 65.960 42.930 ;
        RECT 52.230 42.860 63.760 42.880 ;
        RECT 53.540 42.850 63.760 42.860 ;
        RECT 54.250 42.820 54.560 42.850 ;
        RECT 55.280 42.700 56.290 42.850 ;
        RECT 61.530 42.800 61.850 42.850 ;
        RECT 63.940 42.830 65.960 42.880 ;
        RECT 63.980 42.760 65.960 42.830 ;
        RECT 65.440 42.750 65.960 42.760 ;
    END
  END VINJ
  PIN VGND
    ANTENNADIFFAREA 5.176000 ;
    PORT
      LAYER met2 ;
        RECT 7.300 56.620 7.610 56.830 ;
        RECT 8.730 56.620 9.040 56.850 ;
        RECT 4.950 56.460 9.870 56.620 ;
        RECT 3.140 56.290 9.870 56.460 ;
        RECT 3.140 56.240 9.880 56.290 ;
        RECT 3.140 56.130 9.900 56.240 ;
        RECT 3.140 56.060 5.410 56.130 ;
        RECT 3.140 55.860 3.540 56.060 ;
        RECT 6.510 55.920 6.820 56.130 ;
        RECT 7.440 55.920 7.750 56.130 ;
        RECT 8.140 55.920 8.450 56.130 ;
        RECT 8.880 55.950 9.900 56.130 ;
        RECT 21.990 55.950 22.300 56.070 ;
        RECT 31.850 55.950 32.160 56.090 ;
        RECT 8.880 55.920 32.160 55.950 ;
        RECT 2.790 55.460 3.540 55.860 ;
        RECT 8.900 55.760 32.160 55.920 ;
        RECT 8.900 55.740 32.130 55.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.530 63.860 62.510 64.010 ;
        RECT 61.540 56.610 62.510 63.860 ;
        RECT 61.520 56.140 62.530 56.610 ;
      LAYER via ;
        RECT 61.550 56.180 62.500 56.590 ;
    END
  END VGND
  PIN VPWR
    PORT
      LAYER met1 ;
        RECT 53.020 10.050 53.280 10.510 ;
        RECT 53.760 10.070 54.020 10.510 ;
        RECT 53.010 9.710 53.290 10.050 ;
        RECT 53.750 9.730 54.030 10.070 ;
        RECT 53.020 8.300 53.280 9.710 ;
        RECT 53.760 8.300 54.020 9.730 ;
        RECT 53.020 4.870 54.020 8.300 ;
        RECT 52.540 4.830 54.470 4.870 ;
        RECT 52.000 3.640 54.470 4.830 ;
        RECT 52.000 -7.850 52.940 3.640 ;
      LAYER via ;
        RECT 53.010 9.740 53.290 10.020 ;
        RECT 53.750 9.760 54.030 10.040 ;
        RECT 53.330 4.790 54.450 4.810 ;
        RECT 52.590 3.690 54.450 4.790 ;
        RECT 52.590 3.670 53.710 3.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 62.830 10.050 63.090 10.540 ;
        RECT 62.820 9.710 63.100 10.050 ;
        RECT 62.830 8.530 63.090 9.710 ;
        RECT 63.570 8.530 63.830 10.540 ;
        RECT 62.830 4.890 63.830 8.530 ;
        RECT 63.960 4.890 64.850 4.930 ;
        RECT 62.350 3.610 64.850 4.890 ;
        RECT 63.960 -6.390 64.850 3.610 ;
        RECT 63.960 -7.120 64.880 -6.390 ;
        RECT 63.930 -7.850 64.850 -7.120 ;
      LAYER via ;
        RECT 62.820 9.740 63.100 10.020 ;
        RECT 62.400 3.640 64.260 4.830 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 101.720 48.480 103.450 49.230 ;
        RECT 86.510 45.090 86.830 45.390 ;
        RECT 101.720 44.910 103.460 48.480 ;
        RECT 108.780 45.090 109.100 45.390 ;
        RECT 41.870 43.640 42.110 43.690 ;
        RECT 41.630 43.630 43.100 43.640 ;
        RECT 41.330 43.550 43.100 43.630 ;
        RECT 47.360 43.550 49.570 43.640 ;
        RECT 52.230 43.400 55.540 44.590 ;
        RECT 52.230 43.390 56.190 43.400 ;
        RECT 41.220 36.690 42.990 42.930 ;
        RECT 46.950 36.690 49.460 42.930 ;
        RECT 52.230 40.780 56.200 43.390 ;
        RECT 57.270 42.210 59.990 43.860 ;
        RECT 57.280 42.170 59.990 42.210 ;
        RECT 71.600 43.850 73.330 44.600 ;
        RECT 57.280 40.840 59.990 40.880 ;
        RECT 57.270 40.780 59.990 40.840 ;
        RECT 52.230 40.770 59.990 40.780 ;
        RECT 52.230 40.280 56.200 40.770 ;
        RECT 52.230 40.100 56.270 40.280 ;
        RECT 52.230 38.560 56.200 40.100 ;
        RECT 57.270 39.190 59.990 40.770 ;
        RECT 71.600 40.280 73.340 43.850 ;
        RECT 75.360 42.210 78.080 43.860 ;
        RECT 101.720 43.190 103.450 44.910 ;
        RECT 75.360 42.170 78.070 42.210 ;
        RECT 75.360 40.840 78.070 40.880 ;
        RECT 71.600 38.560 73.330 40.280 ;
        RECT 75.360 39.190 78.080 40.840 ;
        RECT 55.500 37.340 56.200 38.560 ;
        RECT 67.690 37.280 70.240 37.290 ;
        RECT 56.200 35.230 56.280 35.410 ;
        RECT 41.220 26.560 42.990 32.800 ;
        RECT 46.950 26.560 49.460 32.800 ;
        RECT 67.680 31.260 70.240 37.280 ;
        RECT 67.690 31.250 70.240 31.260 ;
        RECT 71.770 31.240 74.000 37.290 ;
        RECT 76.020 35.430 77.750 37.290 ;
        RECT 76.020 33.590 77.760 35.430 ;
        RECT 76.020 31.240 77.750 33.590 ;
        RECT 66.960 23.510 67.360 23.650 ;
        RECT 16.060 18.370 18.430 21.240 ;
        RECT 57.400 12.190 59.420 16.150 ;
        RECT 57.300 12.160 60.690 12.190 ;
        RECT 15.480 4.930 16.100 10.630 ;
        RECT 16.470 7.710 16.480 7.750 ;
        RECT 17.480 4.710 20.870 10.410 ;
        RECT 47.490 6.460 50.880 12.160 ;
        RECT 51.880 9.120 51.890 9.160 ;
        RECT 52.260 6.240 52.880 11.940 ;
        RECT 54.160 6.240 54.780 11.940 ;
        RECT 55.150 9.120 55.160 9.160 ;
        RECT 56.160 6.490 60.690 12.160 ;
        RECT 61.690 9.150 61.700 9.190 ;
        RECT 56.160 6.460 59.550 6.490 ;
        RECT 62.070 6.270 62.690 11.970 ;
        RECT 63.970 6.270 64.590 11.970 ;
        RECT 64.960 9.150 64.970 9.190 ;
        RECT 65.970 6.490 69.360 12.190 ;
        RECT 99.150 -9.940 104.800 6.160 ;
      LAYER li1 ;
        RECT 6.090 61.250 6.260 61.550 ;
        RECT 6.090 61.070 7.090 61.250 ;
        RECT 7.490 61.240 7.660 61.550 ;
        RECT 9.290 61.280 9.960 61.450 ;
        RECT 7.490 61.070 8.500 61.240 ;
        RECT 9.290 60.490 9.960 60.660 ;
        RECT 7.300 60.390 7.620 60.430 ;
        RECT 6.420 60.220 8.500 60.390 ;
        RECT 23.310 60.350 26.620 61.330 ;
        RECT 30.710 60.530 30.940 61.220 ;
        RECT 35.410 60.480 35.640 61.170 ;
        RECT 7.290 60.200 7.620 60.220 ;
        RECT 7.300 60.170 7.620 60.200 ;
        RECT 6.600 59.810 8.420 59.980 ;
        RECT 7.300 59.570 7.620 59.590 ;
        RECT 6.420 59.400 8.500 59.570 ;
        RECT 9.210 59.560 9.420 59.990 ;
        RECT 23.420 59.690 23.590 60.040 ;
        RECT 24.140 59.770 24.310 59.800 ;
        RECT 24.050 59.730 24.370 59.770 ;
        RECT 24.820 59.760 24.990 59.800 ;
        RECT 22.690 59.650 23.590 59.690 ;
        RECT 9.230 59.540 9.400 59.560 ;
        RECT 22.680 59.460 23.590 59.650 ;
        RECT 24.040 59.540 24.370 59.730 ;
        RECT 24.740 59.720 25.060 59.760 ;
        RECT 24.050 59.510 24.370 59.540 ;
        RECT 24.730 59.530 25.060 59.720 ;
        RECT 24.140 59.470 24.310 59.510 ;
        RECT 24.740 59.500 25.060 59.530 ;
        RECT 24.820 59.470 24.990 59.500 ;
        RECT 22.690 59.430 23.590 59.460 ;
        RECT 31.920 59.450 32.090 59.470 ;
        RECT 7.290 59.360 7.620 59.400 ;
        RECT 7.300 59.330 7.620 59.360 ;
        RECT 9.290 59.060 9.960 59.230 ;
        RECT 6.420 58.560 7.090 58.730 ;
        RECT 7.820 58.560 8.500 58.730 ;
        RECT 8.800 58.440 8.990 58.500 ;
        RECT 8.800 58.270 9.970 58.440 ;
        RECT 8.730 57.990 8.900 58.020 ;
        RECT 8.730 57.960 9.060 57.990 ;
        RECT 8.730 57.770 9.070 57.960 ;
        RECT 8.730 57.730 9.060 57.770 ;
        RECT 8.730 57.690 8.900 57.730 ;
        RECT 7.480 57.610 7.650 57.670 ;
        RECT 9.300 57.660 9.970 57.830 ;
        RECT 6.420 57.440 7.090 57.610 ;
        RECT 7.480 57.440 8.500 57.610 ;
        RECT 7.480 57.340 7.650 57.440 ;
        RECT 7.280 56.770 7.600 56.790 ;
        RECT 8.710 56.770 9.030 56.810 ;
        RECT 6.410 56.600 9.990 56.770 ;
        RECT 7.270 56.560 7.600 56.600 ;
        RECT 8.700 56.580 9.030 56.600 ;
        RECT 7.280 56.530 7.600 56.560 ;
        RECT 8.710 56.550 9.030 56.580 ;
        RECT 6.490 56.170 6.810 56.210 ;
        RECT 7.420 56.170 7.740 56.210 ;
        RECT 8.120 56.170 8.440 56.210 ;
        RECT 8.860 56.170 9.180 56.210 ;
        RECT 6.480 56.100 6.810 56.170 ;
        RECT 7.410 56.100 7.740 56.170 ;
        RECT 8.110 56.100 8.440 56.170 ;
        RECT 8.850 56.150 9.180 56.170 ;
        RECT 9.570 56.160 9.890 56.200 ;
        RECT 9.560 56.150 9.890 56.160 ;
        RECT 8.850 56.100 9.890 56.150 ;
        RECT 6.460 55.930 9.890 56.100 ;
        RECT 11.560 55.990 11.730 56.660 ;
        RECT 22.050 56.570 22.220 59.220 ;
        RECT 23.420 59.030 23.590 59.430 ;
        RECT 29.030 59.280 32.090 59.450 ;
        RECT 31.920 58.630 32.090 59.280 ;
        RECT 23.310 57.550 26.620 58.530 ;
        RECT 31.920 58.460 33.190 58.630 ;
        RECT 30.710 57.540 30.940 58.230 ;
        RECT 22.050 56.030 22.230 56.570 ;
        RECT 21.970 55.990 22.290 56.030 ;
        RECT 23.310 56.000 26.620 56.980 ;
        RECT 30.710 56.530 30.940 57.220 ;
        RECT 31.920 56.050 32.090 58.460 ;
        RECT 34.660 56.810 34.830 57.700 ;
        RECT 31.830 56.010 32.150 56.050 ;
        RECT 9.040 55.920 9.890 55.930 ;
        RECT 21.960 55.800 22.290 55.990 ;
        RECT 31.820 55.820 32.150 56.010 ;
        RECT 21.970 55.770 22.290 55.800 ;
        RECT 31.830 55.790 32.150 55.820 ;
        RECT 22.000 52.210 23.520 52.220 ;
        RECT 22.000 51.420 23.550 52.210 ;
        RECT 42.880 50.020 43.230 50.120 ;
        RECT 45.950 50.100 48.180 50.250 ;
        RECT 45.950 50.080 48.330 50.100 ;
        RECT 45.950 50.070 46.130 50.080 ;
        RECT 45.490 50.050 46.130 50.070 ;
        RECT 44.540 50.020 45.000 50.050 ;
        RECT 41.470 49.850 42.230 50.020 ;
        RECT 42.480 49.850 43.650 50.020 ;
        RECT 43.890 49.880 45.000 50.020 ;
        RECT 45.450 49.880 46.130 50.050 ;
        RECT 47.730 49.930 48.330 50.080 ;
        RECT 48.790 49.920 49.120 50.090 ;
        RECT 43.890 49.850 44.710 49.880 ;
        RECT 41.470 49.840 41.700 49.850 ;
        RECT 41.430 49.400 41.700 49.840 ;
        RECT 44.450 49.710 44.710 49.850 ;
        RECT 45.950 49.820 46.130 49.880 ;
        RECT 47.070 49.730 47.400 49.900 ;
        RECT 42.910 49.400 43.240 49.660 ;
        RECT 44.450 49.540 45.630 49.710 ;
        RECT 44.450 49.400 44.710 49.540 ;
        RECT 40.880 49.260 41.050 49.320 ;
        RECT 40.850 49.040 41.070 49.260 ;
        RECT 41.400 49.220 41.730 49.400 ;
        RECT 41.980 49.230 44.140 49.400 ;
        RECT 44.380 49.230 44.710 49.400 ;
        RECT 44.540 49.180 44.710 49.230 ;
        RECT 45.000 49.040 45.210 49.370 ;
        RECT 45.450 49.100 45.630 49.540 ;
        RECT 47.150 49.480 47.400 49.730 ;
        RECT 47.150 49.380 47.620 49.480 ;
        RECT 48.870 49.460 49.050 49.920 ;
        RECT 46.980 49.370 47.620 49.380 ;
        RECT 46.180 49.310 47.620 49.370 ;
        RECT 46.180 49.200 47.540 49.310 ;
        RECT 48.090 49.290 49.050 49.460 ;
        RECT 40.880 48.990 41.050 49.040 ;
        RECT 42.880 48.470 43.230 48.570 ;
        RECT 45.950 48.550 48.180 48.700 ;
        RECT 45.950 48.530 48.330 48.550 ;
        RECT 45.950 48.520 46.130 48.530 ;
        RECT 45.490 48.500 46.130 48.520 ;
        RECT 44.540 48.470 45.000 48.500 ;
        RECT 41.470 48.300 42.230 48.470 ;
        RECT 42.480 48.300 43.650 48.470 ;
        RECT 43.890 48.330 45.000 48.470 ;
        RECT 45.450 48.330 46.130 48.500 ;
        RECT 47.730 48.380 48.330 48.530 ;
        RECT 48.790 48.370 49.120 48.540 ;
        RECT 43.890 48.300 44.710 48.330 ;
        RECT 41.470 48.290 41.700 48.300 ;
        RECT 41.430 47.850 41.700 48.290 ;
        RECT 44.450 48.160 44.710 48.300 ;
        RECT 45.950 48.270 46.130 48.330 ;
        RECT 47.070 48.180 47.400 48.350 ;
        RECT 42.910 47.850 43.240 48.110 ;
        RECT 44.450 47.990 45.630 48.160 ;
        RECT 44.450 47.850 44.710 47.990 ;
        RECT 40.880 47.710 41.050 47.770 ;
        RECT 40.850 47.490 41.070 47.710 ;
        RECT 41.400 47.670 41.730 47.850 ;
        RECT 41.980 47.680 44.140 47.850 ;
        RECT 44.380 47.680 44.710 47.850 ;
        RECT 44.540 47.630 44.710 47.680 ;
        RECT 45.000 47.490 45.210 47.820 ;
        RECT 45.450 47.550 45.630 47.990 ;
        RECT 47.150 47.930 47.400 48.180 ;
        RECT 47.150 47.830 47.620 47.930 ;
        RECT 48.870 47.910 49.050 48.370 ;
        RECT 69.970 48.260 70.640 49.130 ;
        RECT 82.250 48.820 84.350 49.130 ;
        RECT 82.250 48.650 84.770 48.820 ;
        RECT 85.010 48.800 85.200 48.830 ;
        RECT 82.250 48.280 84.350 48.650 ;
        RECT 85.010 48.630 86.070 48.800 ;
        RECT 110.830 48.650 111.360 48.820 ;
        RECT 85.010 48.600 85.200 48.630 ;
        RECT 82.750 47.940 82.970 48.280 ;
        RECT 82.750 47.930 82.960 47.940 ;
        RECT 46.980 47.820 47.620 47.830 ;
        RECT 46.180 47.760 47.620 47.820 ;
        RECT 46.180 47.650 47.540 47.760 ;
        RECT 48.090 47.740 49.050 47.910 ;
        RECT 83.130 47.760 83.320 47.770 ;
        RECT 40.880 47.440 41.050 47.490 ;
        RECT 83.120 47.470 83.320 47.760 ;
        RECT 42.880 46.920 43.230 47.020 ;
        RECT 45.950 47.000 48.180 47.150 ;
        RECT 83.090 47.140 83.330 47.470 ;
        RECT 45.950 46.980 48.330 47.000 ;
        RECT 45.950 46.970 46.130 46.980 ;
        RECT 45.490 46.950 46.130 46.970 ;
        RECT 44.540 46.920 45.000 46.950 ;
        RECT 20.210 46.790 20.410 46.830 ;
        RECT 19.900 46.530 20.410 46.790 ;
        RECT 20.210 46.500 20.410 46.530 ;
        RECT 20.800 46.800 21.000 46.830 ;
        RECT 20.800 46.760 21.310 46.800 ;
        RECT 20.800 46.570 21.320 46.760 ;
        RECT 41.470 46.750 42.230 46.920 ;
        RECT 42.480 46.750 43.650 46.920 ;
        RECT 43.890 46.780 45.000 46.920 ;
        RECT 45.450 46.780 46.130 46.950 ;
        RECT 47.730 46.830 48.330 46.980 ;
        RECT 48.790 46.820 49.120 46.990 ;
        RECT 43.890 46.750 44.710 46.780 ;
        RECT 41.470 46.740 41.700 46.750 ;
        RECT 20.800 46.540 21.310 46.570 ;
        RECT 20.800 46.500 21.000 46.540 ;
        RECT 21.490 46.350 21.660 46.400 ;
        RECT 19.460 46.330 19.890 46.350 ;
        RECT 19.460 46.160 19.910 46.330 ;
        RECT 21.480 46.320 21.660 46.350 ;
        RECT 21.480 46.310 21.910 46.320 ;
        RECT 19.460 46.140 19.890 46.160 ;
        RECT 21.480 46.080 22.070 46.310 ;
        RECT 41.430 46.300 41.700 46.740 ;
        RECT 44.450 46.610 44.710 46.750 ;
        RECT 45.950 46.720 46.130 46.780 ;
        RECT 47.070 46.630 47.400 46.800 ;
        RECT 42.910 46.300 43.240 46.560 ;
        RECT 44.450 46.440 45.630 46.610 ;
        RECT 44.450 46.300 44.710 46.440 ;
        RECT 40.880 46.160 41.050 46.220 ;
        RECT 21.480 46.070 21.910 46.080 ;
        RECT 21.480 46.010 21.650 46.070 ;
        RECT 40.850 45.940 41.070 46.160 ;
        RECT 41.400 46.120 41.730 46.300 ;
        RECT 41.980 46.130 44.140 46.300 ;
        RECT 44.380 46.130 44.710 46.300 ;
        RECT 44.540 46.080 44.710 46.130 ;
        RECT 45.000 45.940 45.210 46.270 ;
        RECT 45.450 46.000 45.630 46.440 ;
        RECT 47.150 46.380 47.400 46.630 ;
        RECT 47.150 46.280 47.620 46.380 ;
        RECT 48.870 46.360 49.050 46.820 ;
        RECT 83.520 46.660 83.690 48.270 ;
        RECT 84.350 47.170 84.520 48.260 ;
        RECT 85.480 48.240 85.670 48.270 ;
        RECT 84.940 48.070 85.670 48.240 ;
        RECT 85.900 48.240 86.070 48.630 ;
        RECT 112.640 48.550 112.840 48.900 ;
        RECT 112.640 48.520 112.850 48.550 ;
        RECT 85.900 48.070 86.640 48.240 ;
        RECT 108.960 48.070 109.310 48.240 ;
        RECT 110.330 48.070 110.660 48.240 ;
        RECT 85.480 48.040 85.670 48.070 ;
        RECT 87.700 47.450 87.930 47.970 ;
        RECT 84.940 47.280 87.930 47.450 ;
        RECT 84.120 47.130 84.520 47.170 ;
        RECT 84.110 46.940 84.520 47.130 ;
        RECT 92.900 47.090 93.450 47.520 ;
        RECT 102.150 47.090 102.700 47.520 ;
        RECT 105.780 47.280 106.010 47.970 ;
        RECT 111.080 47.740 111.250 48.260 ;
        RECT 110.920 47.480 111.250 47.740 ;
        RECT 108.960 47.280 109.310 47.450 ;
        RECT 110.330 47.280 110.660 47.450 ;
        RECT 84.120 46.910 84.520 46.940 ;
        RECT 83.510 46.470 83.690 46.660 ;
        RECT 84.350 46.570 84.520 46.910 ;
        RECT 85.010 46.660 85.200 46.840 ;
        RECT 84.940 46.490 85.290 46.660 ;
        RECT 46.980 46.270 47.620 46.280 ;
        RECT 46.180 46.210 47.620 46.270 ;
        RECT 46.180 46.100 47.540 46.210 ;
        RECT 48.090 46.190 49.050 46.360 ;
        RECT 85.860 46.080 86.070 46.510 ;
        RECT 86.290 46.490 86.630 46.660 ;
        RECT 85.880 46.060 86.050 46.080 ;
        RECT 20.210 45.870 20.410 45.910 ;
        RECT 19.900 45.610 20.410 45.870 ;
        RECT 20.210 45.580 20.410 45.610 ;
        RECT 20.800 45.880 21.000 45.910 ;
        RECT 40.880 45.890 41.050 45.940 ;
        RECT 20.800 45.840 21.310 45.880 ;
        RECT 20.800 45.650 21.320 45.840 ;
        RECT 83.510 45.750 83.690 45.940 ;
        RECT 20.800 45.620 21.310 45.650 ;
        RECT 20.800 45.580 21.000 45.620 ;
        RECT 19.460 45.410 19.890 45.430 ;
        RECT 19.460 45.240 19.910 45.410 ;
        RECT 42.880 45.370 43.230 45.470 ;
        RECT 45.950 45.450 48.180 45.600 ;
        RECT 45.950 45.430 48.330 45.450 ;
        RECT 45.950 45.420 46.130 45.430 ;
        RECT 45.490 45.400 46.130 45.420 ;
        RECT 44.540 45.370 45.000 45.400 ;
        RECT 19.460 45.220 19.890 45.240 ;
        RECT 41.470 45.200 42.230 45.370 ;
        RECT 42.480 45.200 43.650 45.370 ;
        RECT 43.890 45.230 45.000 45.370 ;
        RECT 45.450 45.230 46.130 45.400 ;
        RECT 47.730 45.280 48.330 45.430 ;
        RECT 48.790 45.270 49.120 45.440 ;
        RECT 43.890 45.200 44.710 45.230 ;
        RECT 41.470 45.190 41.700 45.200 ;
        RECT 20.210 44.950 20.410 44.990 ;
        RECT 19.900 44.690 20.410 44.950 ;
        RECT 20.210 44.660 20.410 44.690 ;
        RECT 20.800 44.960 21.000 44.990 ;
        RECT 20.800 44.920 21.310 44.960 ;
        RECT 20.800 44.730 21.320 44.920 ;
        RECT 41.430 44.750 41.700 45.190 ;
        RECT 44.450 45.060 44.710 45.200 ;
        RECT 45.950 45.170 46.130 45.230 ;
        RECT 47.070 45.080 47.400 45.250 ;
        RECT 42.910 44.750 43.240 45.010 ;
        RECT 44.450 44.890 45.630 45.060 ;
        RECT 44.450 44.750 44.710 44.890 ;
        RECT 20.800 44.700 21.310 44.730 ;
        RECT 20.800 44.660 21.000 44.700 ;
        RECT 40.880 44.610 41.050 44.670 ;
        RECT 19.460 44.490 19.890 44.510 ;
        RECT 19.460 44.320 19.910 44.490 ;
        RECT 40.850 44.390 41.070 44.610 ;
        RECT 41.400 44.570 41.730 44.750 ;
        RECT 41.980 44.580 44.140 44.750 ;
        RECT 44.380 44.580 44.710 44.750 ;
        RECT 44.540 44.530 44.710 44.580 ;
        RECT 45.000 44.390 45.210 44.720 ;
        RECT 45.450 44.450 45.630 44.890 ;
        RECT 47.150 44.830 47.400 45.080 ;
        RECT 47.150 44.730 47.620 44.830 ;
        RECT 48.870 44.810 49.050 45.270 ;
        RECT 83.090 44.940 83.330 45.270 ;
        RECT 46.980 44.720 47.620 44.730 ;
        RECT 46.180 44.660 47.620 44.720 ;
        RECT 46.180 44.550 47.540 44.660 ;
        RECT 48.090 44.640 49.050 44.810 ;
        RECT 83.120 44.650 83.320 44.940 ;
        RECT 83.130 44.640 83.320 44.650 ;
        RECT 82.750 44.470 82.960 44.480 ;
        RECT 40.880 44.340 41.050 44.390 ;
        RECT 19.460 44.300 19.890 44.320 ;
        RECT 19.710 43.930 20.030 43.970 ;
        RECT 19.710 43.910 20.040 43.930 ;
        RECT 52.630 43.920 52.830 44.270 ;
        RECT 54.110 44.020 54.640 44.190 ;
        RECT 19.710 43.710 20.330 43.910 ;
        RECT 20.160 43.580 20.330 43.710 ;
        RECT 20.840 43.870 21.010 43.910 ;
        RECT 52.620 43.890 52.830 43.920 ;
        RECT 20.840 43.830 21.330 43.870 ;
        RECT 20.840 43.640 21.340 43.830 ;
        RECT 20.840 43.610 21.330 43.640 ;
        RECT 20.840 43.580 21.010 43.610 ;
        RECT 19.550 43.470 19.980 43.490 ;
        RECT 19.530 43.300 19.980 43.470 ;
        RECT 52.620 43.310 52.840 43.890 ;
        RECT 52.620 43.300 52.830 43.310 ;
        RECT 19.550 43.280 19.980 43.300 ;
        RECT 53.000 43.130 53.190 43.140 ;
        RECT 19.710 42.970 20.030 43.010 ;
        RECT 19.710 42.950 20.040 42.970 ;
        RECT 19.710 42.750 20.330 42.950 ;
        RECT 20.160 42.620 20.330 42.750 ;
        RECT 20.840 42.910 21.010 42.950 ;
        RECT 20.840 42.870 21.330 42.910 ;
        RECT 20.840 42.680 21.340 42.870 ;
        RECT 52.990 42.840 53.190 43.130 ;
        RECT 40.880 42.790 41.050 42.840 ;
        RECT 20.840 42.650 21.330 42.680 ;
        RECT 20.840 42.620 21.010 42.650 ;
        RECT 40.850 42.570 41.070 42.790 ;
        RECT 19.550 42.510 19.980 42.530 ;
        RECT 40.880 42.510 41.050 42.570 ;
        RECT 19.530 42.340 19.980 42.510 ;
        RECT 41.400 42.430 41.730 42.610 ;
        RECT 44.540 42.600 44.710 42.650 ;
        RECT 41.980 42.430 44.140 42.600 ;
        RECT 44.380 42.430 44.710 42.600 ;
        RECT 45.000 42.460 45.210 42.790 ;
        RECT 19.550 42.320 19.980 42.340 ;
        RECT 19.710 42.010 20.030 42.050 ;
        RECT 19.710 41.990 20.040 42.010 ;
        RECT 41.430 41.990 41.700 42.430 ;
        RECT 42.910 42.170 43.240 42.430 ;
        RECT 44.450 42.290 44.710 42.430 ;
        RECT 45.450 42.290 45.630 42.730 ;
        RECT 46.180 42.520 47.540 42.630 ;
        RECT 46.180 42.460 47.620 42.520 ;
        RECT 46.980 42.450 47.620 42.460 ;
        RECT 19.710 41.790 20.330 41.990 ;
        RECT 20.160 41.660 20.330 41.790 ;
        RECT 20.840 41.950 21.010 41.990 ;
        RECT 41.470 41.980 41.700 41.990 ;
        RECT 44.450 42.120 45.630 42.290 ;
        RECT 47.150 42.350 47.620 42.450 ;
        RECT 48.090 42.370 49.050 42.540 ;
        RECT 52.960 42.510 53.200 42.840 ;
        RECT 44.450 41.980 44.710 42.120 ;
        RECT 47.150 42.100 47.400 42.350 ;
        RECT 20.840 41.910 21.330 41.950 ;
        RECT 20.840 41.720 21.340 41.910 ;
        RECT 41.470 41.810 42.230 41.980 ;
        RECT 42.480 41.810 43.650 41.980 ;
        RECT 43.890 41.950 44.710 41.980 ;
        RECT 45.950 41.950 46.130 42.010 ;
        RECT 43.890 41.810 45.000 41.950 ;
        RECT 20.840 41.690 21.330 41.720 ;
        RECT 42.880 41.710 43.230 41.810 ;
        RECT 44.540 41.780 45.000 41.810 ;
        RECT 45.450 41.780 46.130 41.950 ;
        RECT 47.070 41.930 47.400 42.100 ;
        RECT 48.870 41.910 49.050 42.370 ;
        RECT 53.390 42.030 53.560 43.640 ;
        RECT 45.490 41.760 46.130 41.780 ;
        RECT 45.950 41.750 46.130 41.760 ;
        RECT 47.730 41.750 48.330 41.900 ;
        RECT 45.950 41.730 48.330 41.750 ;
        RECT 48.790 41.740 49.120 41.910 ;
        RECT 53.380 41.840 53.560 42.030 ;
        RECT 54.220 43.110 54.390 43.630 ;
        RECT 54.810 43.440 55.140 43.610 ;
        RECT 56.160 43.440 56.510 43.610 ;
        RECT 56.830 43.590 61.890 44.420 ;
        RECT 80.710 44.020 81.240 44.190 ;
        RECT 82.520 43.920 82.720 44.270 ;
        RECT 82.520 43.890 82.730 43.920 ;
        RECT 61.340 43.510 61.820 43.590 ;
        RECT 54.220 42.850 54.550 43.110 ;
        RECT 54.220 41.940 54.390 42.850 ;
        RECT 54.810 42.650 55.140 42.820 ;
        RECT 56.160 42.650 56.510 42.820 ;
        RECT 59.460 42.650 59.690 43.340 ;
        RECT 61.340 43.260 61.810 43.510 ;
        RECT 78.840 43.440 79.190 43.610 ;
        RECT 80.210 43.440 80.540 43.610 ;
        RECT 60.650 42.750 60.820 43.170 ;
        RECT 61.460 43.050 61.700 43.080 ;
        RECT 61.130 42.880 61.700 43.050 ;
        RECT 61.940 42.890 63.280 43.050 ;
        RECT 61.940 42.880 63.320 42.890 ;
        RECT 63.730 42.880 64.690 43.050 ;
        RECT 61.460 42.840 61.700 42.880 ;
        RECT 60.580 42.530 60.750 42.570 ;
        RECT 60.520 42.360 60.750 42.530 ;
        RECT 62.770 42.460 63.320 42.880 ;
        RECT 64.240 42.870 64.410 42.880 ;
        RECT 60.580 42.030 60.750 42.360 ;
        RECT 60.920 42.430 61.110 42.450 ;
        RECT 63.920 42.430 64.250 42.610 ;
        RECT 60.920 42.260 61.480 42.430 ;
        RECT 61.940 42.260 64.690 42.430 ;
        RECT 60.920 42.220 61.110 42.260 ;
        RECT 65.220 42.190 65.390 43.120 ;
        RECT 65.620 42.320 65.790 43.170 ;
        RECT 72.030 42.460 72.580 42.890 ;
        RECT 75.660 42.650 75.890 43.340 ;
        RECT 80.960 43.110 81.130 43.630 ;
        RECT 80.800 42.850 81.130 43.110 ;
        RECT 78.840 42.650 79.190 42.820 ;
        RECT 80.210 42.650 80.540 42.820 ;
        RECT 54.810 41.860 55.140 42.030 ;
        RECT 56.160 41.860 56.500 42.030 ;
        RECT 60.530 42.010 60.750 42.030 ;
        RECT 20.840 41.660 21.010 41.690 ;
        RECT 45.950 41.580 48.180 41.730 ;
        RECT 19.550 41.550 19.980 41.570 ;
        RECT 19.530 41.380 19.980 41.550 ;
        RECT 19.550 41.360 19.980 41.380 ;
        RECT 21.340 41.320 21.760 41.490 ;
        RECT 21.440 41.280 21.670 41.320 ;
        RECT 40.880 41.240 41.050 41.290 ;
        RECT 40.850 41.020 41.070 41.240 ;
        RECT 40.880 40.960 41.050 41.020 ;
        RECT 41.400 40.880 41.730 41.060 ;
        RECT 44.540 41.050 44.710 41.100 ;
        RECT 41.980 40.880 44.140 41.050 ;
        RECT 44.380 40.880 44.710 41.050 ;
        RECT 45.000 40.910 45.210 41.240 ;
        RECT 41.430 40.440 41.700 40.880 ;
        RECT 42.910 40.620 43.240 40.880 ;
        RECT 44.450 40.740 44.710 40.880 ;
        RECT 45.450 40.740 45.630 41.180 ;
        RECT 53.380 41.120 53.560 41.310 ;
        RECT 54.890 41.290 55.060 41.860 ;
        RECT 60.530 41.770 60.720 42.010 ;
        RECT 60.530 41.630 60.750 41.770 ;
        RECT 74.630 41.630 74.820 42.030 ;
        RECT 78.850 41.860 79.190 42.030 ;
        RECT 80.210 41.860 80.540 42.030 ;
        RECT 80.960 41.940 81.130 42.850 ;
        RECT 81.790 42.030 81.960 43.640 ;
        RECT 82.510 43.310 82.730 43.890 ;
        RECT 82.750 43.890 82.970 44.470 ;
        RECT 83.520 44.140 83.690 45.750 ;
        RECT 84.350 45.480 84.520 45.840 ;
        RECT 84.940 45.750 85.290 45.920 ;
        RECT 85.480 45.900 85.670 45.950 ;
        RECT 86.380 45.920 86.550 46.490 ;
        RECT 90.660 46.260 90.850 46.660 ;
        RECT 104.750 46.260 104.940 46.660 ;
        RECT 108.970 46.490 109.310 46.660 ;
        RECT 110.330 46.490 110.660 46.660 ;
        RECT 111.080 46.570 111.250 47.480 ;
        RECT 111.910 46.660 112.080 48.270 ;
        RECT 112.630 47.940 112.850 48.520 ;
        RECT 112.640 47.930 112.850 47.940 ;
        RECT 112.280 47.760 112.470 47.770 ;
        RECT 112.280 47.470 112.480 47.760 ;
        RECT 112.270 47.140 112.510 47.470 ;
        RECT 90.660 46.250 91.040 46.260 ;
        RECT 87.300 46.070 91.040 46.250 ;
        RECT 90.660 46.030 91.040 46.070 ;
        RECT 104.560 46.250 104.940 46.260 ;
        RECT 104.560 46.070 108.300 46.250 ;
        RECT 104.560 46.030 104.940 46.070 ;
        RECT 85.480 45.890 85.710 45.900 ;
        RECT 86.290 45.890 86.630 45.920 ;
        RECT 85.480 45.750 86.630 45.890 ;
        RECT 85.020 45.540 85.210 45.750 ;
        RECT 85.480 45.720 86.460 45.750 ;
        RECT 85.620 45.690 86.460 45.720 ;
        RECT 90.660 45.650 90.850 46.030 ;
        RECT 84.110 45.440 84.520 45.480 ;
        RECT 84.100 45.250 84.520 45.440 ;
        RECT 92.900 45.360 93.450 45.790 ;
        RECT 102.150 45.360 102.700 45.790 ;
        RECT 104.750 45.650 104.940 46.030 ;
        RECT 110.410 45.920 110.580 46.490 ;
        RECT 111.910 46.470 112.090 46.660 ;
        RECT 108.970 45.750 109.310 45.920 ;
        RECT 110.330 45.750 110.660 45.920 ;
        RECT 110.260 45.360 110.430 45.410 ;
        RECT 84.110 45.220 84.520 45.250 ;
        RECT 84.350 44.150 84.520 45.220 ;
        RECT 84.940 45.030 87.870 45.130 ;
        RECT 84.940 44.960 87.930 45.030 ;
        RECT 86.960 44.640 87.130 44.700 ;
        RECT 86.940 44.430 87.150 44.640 ;
        RECT 85.470 44.340 85.660 44.370 ;
        RECT 86.960 44.360 87.130 44.430 ;
        RECT 87.700 44.340 87.930 44.960 ;
        RECT 105.780 44.340 106.010 45.070 ;
        RECT 108.960 44.960 109.310 45.130 ;
        RECT 110.260 45.100 110.820 45.360 ;
        RECT 110.260 45.080 110.660 45.100 ;
        RECT 110.330 44.960 110.660 45.080 ;
        RECT 111.080 44.980 111.250 45.840 ;
        RECT 111.910 45.750 112.090 45.940 ;
        RECT 111.910 45.120 112.080 45.750 ;
        RECT 111.730 45.080 112.080 45.120 ;
        RECT 84.940 44.170 85.660 44.340 ;
        RECT 85.470 44.140 85.660 44.170 ;
        RECT 85.830 44.170 86.640 44.340 ;
        RECT 108.960 44.170 109.310 44.340 ;
        RECT 82.750 43.860 82.960 43.890 ;
        RECT 82.760 43.510 82.960 43.860 ;
        RECT 85.040 43.830 85.230 43.860 ;
        RECT 85.830 43.830 86.020 44.170 ;
        RECT 109.680 44.000 109.860 44.930 ;
        RECT 110.410 44.670 110.740 44.840 ;
        RECT 110.920 44.720 111.250 44.980 ;
        RECT 111.500 44.820 112.080 45.080 ;
        RECT 112.270 45.120 112.510 45.270 ;
        RECT 112.270 44.940 112.870 45.120 ;
        RECT 111.730 44.790 112.080 44.820 ;
        RECT 110.490 44.530 110.740 44.670 ;
        RECT 110.490 44.340 110.970 44.530 ;
        RECT 110.330 44.270 110.970 44.340 ;
        RECT 110.330 44.170 110.660 44.270 ;
        RECT 109.560 43.970 109.880 44.000 ;
        RECT 110.490 43.970 110.660 44.170 ;
        RECT 111.080 44.150 111.250 44.720 ;
        RECT 111.320 44.430 111.490 44.470 ;
        RECT 111.910 44.460 112.080 44.790 ;
        RECT 112.280 44.640 112.870 44.940 ;
        RECT 113.690 45.000 114.270 45.170 ;
        RECT 113.690 44.900 114.080 45.000 ;
        RECT 113.690 44.870 114.070 44.900 ;
        RECT 113.690 44.720 114.050 44.870 ;
        RECT 111.730 44.430 112.080 44.460 ;
        RECT 111.320 44.170 112.080 44.430 ;
        RECT 111.320 44.140 111.490 44.170 ;
        RECT 111.730 44.140 112.080 44.170 ;
        RECT 111.730 44.130 111.930 44.140 ;
        RECT 112.320 44.130 112.870 44.640 ;
        RECT 113.340 44.550 114.050 44.720 ;
        RECT 109.090 43.940 109.410 43.970 ;
        RECT 84.240 43.590 84.770 43.760 ;
        RECT 85.040 43.650 86.020 43.830 ;
        RECT 85.040 43.630 85.230 43.650 ;
        RECT 107.870 43.600 108.040 43.880 ;
        RECT 109.090 43.750 109.420 43.940 ;
        RECT 109.560 43.800 109.890 43.970 ;
        RECT 110.490 43.940 110.980 43.970 ;
        RECT 110.100 43.800 110.290 43.820 ;
        RECT 109.090 43.710 109.410 43.750 ;
        RECT 109.560 43.740 110.290 43.800 ;
        RECT 107.870 43.560 108.080 43.600 ;
        RECT 107.870 43.540 108.100 43.560 ;
        RECT 109.220 43.550 109.390 43.710 ;
        RECT 109.680 43.630 110.290 43.740 ;
        RECT 107.870 43.520 108.130 43.540 ;
        RECT 107.870 43.470 108.210 43.520 ;
        RECT 107.870 43.410 108.360 43.470 ;
        RECT 107.870 43.380 108.380 43.410 ;
        RECT 107.910 43.350 108.380 43.380 ;
        RECT 82.520 43.300 82.730 43.310 ;
        RECT 108.040 43.300 108.380 43.350 ;
        RECT 109.680 43.300 109.860 43.630 ;
        RECT 110.080 43.620 110.290 43.630 ;
        RECT 110.100 43.590 110.290 43.620 ;
        RECT 110.490 43.760 110.990 43.940 ;
        RECT 112.630 43.890 112.850 44.130 ;
        RECT 111.230 43.800 111.420 43.830 ;
        RECT 111.230 43.760 111.670 43.800 ;
        RECT 110.490 43.710 111.670 43.760 ;
        RECT 108.160 43.290 108.380 43.300 ;
        RECT 108.170 43.260 108.380 43.290 ;
        RECT 108.190 43.180 108.380 43.260 ;
        RECT 109.550 43.180 109.880 43.300 ;
        RECT 110.490 43.180 110.660 43.710 ;
        RECT 110.720 43.630 111.670 43.710 ;
        RECT 110.720 43.600 111.490 43.630 ;
        RECT 111.730 43.600 111.930 43.640 ;
        RECT 110.720 43.590 111.930 43.600 ;
        RECT 110.720 43.550 110.890 43.590 ;
        RECT 111.320 43.340 111.930 43.590 ;
        RECT 111.320 43.300 111.490 43.340 ;
        RECT 111.730 43.310 111.930 43.340 ;
        RECT 111.950 43.210 112.120 43.890 ;
        RECT 112.640 43.860 112.850 43.890 ;
        RECT 112.640 43.640 112.840 43.860 ;
        RECT 113.340 43.800 114.040 44.110 ;
        RECT 82.160 43.130 82.350 43.140 ;
        RECT 107.700 43.130 107.870 43.150 ;
        RECT 82.160 42.840 82.360 43.130 ;
        RECT 82.150 42.510 82.390 42.840 ;
        RECT 107.680 42.700 107.890 43.130 ;
        RECT 108.190 43.010 108.710 43.180 ;
        RECT 108.190 42.980 108.380 43.010 ;
        RECT 109.060 43.000 110.960 43.180 ;
        RECT 111.690 43.170 112.120 43.210 ;
        RECT 111.340 43.010 112.120 43.170 ;
        RECT 111.340 43.000 111.880 43.010 ;
        RECT 107.680 42.060 107.890 42.490 ;
        RECT 108.190 42.180 108.380 42.210 ;
        RECT 109.680 42.190 109.860 43.000 ;
        RECT 110.490 42.890 110.660 43.000 ;
        RECT 111.690 42.980 111.880 43.000 ;
        RECT 111.730 42.950 111.930 42.980 ;
        RECT 110.290 42.690 110.610 42.720 ;
        RECT 111.500 42.690 111.930 42.950 ;
        RECT 110.290 42.500 110.620 42.690 ;
        RECT 111.730 42.650 111.930 42.690 ;
        RECT 112.320 42.650 112.870 43.640 ;
        RECT 113.190 43.570 114.040 43.800 ;
        RECT 113.340 43.230 114.040 43.570 ;
        RECT 113.800 42.870 114.120 42.910 ;
        RECT 113.800 42.810 114.130 42.870 ;
        RECT 113.330 42.680 114.130 42.810 ;
        RECT 113.330 42.650 114.120 42.680 ;
        RECT 113.330 42.630 114.030 42.650 ;
        RECT 110.290 42.460 110.610 42.500 ;
        RECT 110.290 42.380 110.460 42.460 ;
        RECT 110.240 42.210 110.460 42.380 ;
        RECT 110.240 42.190 110.410 42.210 ;
        RECT 111.690 42.190 111.880 42.210 ;
        RECT 107.700 42.040 107.870 42.060 ;
        RECT 60.530 41.620 60.910 41.630 ;
        RECT 57.170 41.440 60.910 41.620 ;
        RECT 74.440 41.620 74.820 41.630 ;
        RECT 60.530 41.420 60.910 41.440 ;
        RECT 60.520 41.400 60.910 41.420 ;
        RECT 60.920 41.520 61.110 41.560 ;
        RECT 46.180 40.970 47.540 41.080 ;
        RECT 46.180 40.910 47.620 40.970 ;
        RECT 46.980 40.900 47.620 40.910 ;
        RECT 41.470 40.430 41.700 40.440 ;
        RECT 44.450 40.570 45.630 40.740 ;
        RECT 47.150 40.800 47.620 40.900 ;
        RECT 48.090 40.820 49.050 40.990 ;
        RECT 44.450 40.430 44.710 40.570 ;
        RECT 47.150 40.550 47.400 40.800 ;
        RECT 41.470 40.260 42.230 40.430 ;
        RECT 42.480 40.260 43.650 40.430 ;
        RECT 43.890 40.400 44.710 40.430 ;
        RECT 45.950 40.400 46.130 40.460 ;
        RECT 43.890 40.260 45.000 40.400 ;
        RECT 42.880 40.160 43.230 40.260 ;
        RECT 44.540 40.230 45.000 40.260 ;
        RECT 45.450 40.230 46.130 40.400 ;
        RECT 47.070 40.380 47.400 40.550 ;
        RECT 48.870 40.360 49.050 40.820 ;
        RECT 45.490 40.210 46.130 40.230 ;
        RECT 45.950 40.200 46.130 40.210 ;
        RECT 47.730 40.200 48.330 40.350 ;
        RECT 45.950 40.180 48.330 40.200 ;
        RECT 48.790 40.190 49.120 40.360 ;
        RECT 52.960 40.310 53.200 40.640 ;
        RECT 45.950 40.030 48.180 40.180 ;
        RECT 52.990 40.020 53.190 40.310 ;
        RECT 53.000 40.010 53.190 40.020 ;
        RECT 52.620 39.840 52.830 39.850 ;
        RECT 40.880 39.690 41.050 39.740 ;
        RECT 40.850 39.470 41.070 39.690 ;
        RECT 40.880 39.410 41.050 39.470 ;
        RECT 41.400 39.330 41.730 39.510 ;
        RECT 44.540 39.500 44.710 39.550 ;
        RECT 41.980 39.330 44.140 39.500 ;
        RECT 44.380 39.330 44.710 39.500 ;
        RECT 45.000 39.360 45.210 39.690 ;
        RECT 41.430 38.890 41.700 39.330 ;
        RECT 42.910 39.070 43.240 39.330 ;
        RECT 44.450 39.190 44.710 39.330 ;
        RECT 45.450 39.190 45.630 39.630 ;
        RECT 46.180 39.420 47.540 39.530 ;
        RECT 46.180 39.360 47.620 39.420 ;
        RECT 46.980 39.350 47.620 39.360 ;
        RECT 41.470 38.880 41.700 38.890 ;
        RECT 44.450 39.020 45.630 39.190 ;
        RECT 47.150 39.250 47.620 39.350 ;
        RECT 48.090 39.270 49.050 39.440 ;
        RECT 44.450 38.880 44.710 39.020 ;
        RECT 47.150 39.000 47.400 39.250 ;
        RECT 41.470 38.710 42.230 38.880 ;
        RECT 42.480 38.710 43.650 38.880 ;
        RECT 43.890 38.850 44.710 38.880 ;
        RECT 45.950 38.850 46.130 38.910 ;
        RECT 43.890 38.710 45.000 38.850 ;
        RECT 42.880 38.610 43.230 38.710 ;
        RECT 44.540 38.680 45.000 38.710 ;
        RECT 45.450 38.680 46.130 38.850 ;
        RECT 47.070 38.830 47.400 39.000 ;
        RECT 48.870 38.810 49.050 39.270 ;
        RECT 52.620 39.260 52.840 39.840 ;
        RECT 53.390 39.510 53.560 41.120 ;
        RECT 54.220 40.350 54.390 41.210 ;
        RECT 54.810 41.120 55.140 41.290 ;
        RECT 56.160 41.120 56.500 41.290 ;
        RECT 60.520 41.250 60.750 41.400 ;
        RECT 60.920 41.350 61.480 41.520 ;
        RECT 61.940 41.350 64.690 41.520 ;
        RECT 60.920 41.330 61.110 41.350 ;
        RECT 60.530 41.210 60.750 41.250 ;
        RECT 60.530 41.030 60.720 41.210 ;
        RECT 63.920 41.170 64.250 41.350 ;
        RECT 60.530 41.020 60.820 41.030 ;
        RECT 60.650 40.610 60.820 41.020 ;
        RECT 61.460 40.900 61.700 40.940 ;
        RECT 62.770 40.900 63.320 41.160 ;
        RECT 64.240 40.900 64.410 40.910 ;
        RECT 61.130 40.730 61.700 40.900 ;
        RECT 61.940 40.730 63.320 40.900 ;
        RECT 63.730 40.730 64.690 40.900 ;
        RECT 61.460 40.700 61.700 40.730 ;
        RECT 65.220 40.660 65.390 41.590 ;
        RECT 65.620 40.610 65.790 41.460 ;
        RECT 74.440 41.440 78.180 41.620 ;
        RECT 74.440 41.400 74.820 41.440 ;
        RECT 72.030 40.730 72.580 41.160 ;
        RECT 74.630 41.020 74.820 41.400 ;
        RECT 80.290 41.290 80.460 41.860 ;
        RECT 81.790 41.840 81.970 42.030 ;
        RECT 108.190 42.010 108.710 42.180 ;
        RECT 109.060 42.010 110.960 42.190 ;
        RECT 111.340 42.180 111.880 42.190 ;
        RECT 111.340 42.020 112.120 42.180 ;
        RECT 108.190 41.930 108.380 42.010 ;
        RECT 108.170 41.900 108.380 41.930 ;
        RECT 108.160 41.890 108.380 41.900 ;
        RECT 109.550 41.890 109.880 42.010 ;
        RECT 111.500 41.980 112.120 42.020 ;
        RECT 108.040 41.840 108.380 41.890 ;
        RECT 107.910 41.810 108.380 41.840 ;
        RECT 107.870 41.780 108.380 41.810 ;
        RECT 107.870 41.720 108.360 41.780 ;
        RECT 107.870 41.670 108.210 41.720 ;
        RECT 107.870 41.650 108.130 41.670 ;
        RECT 107.870 41.630 108.100 41.650 ;
        RECT 107.870 41.590 108.080 41.630 ;
        RECT 107.870 41.310 108.040 41.590 ;
        RECT 109.220 41.480 109.390 41.640 ;
        RECT 109.680 41.560 109.860 41.890 ;
        RECT 110.770 41.790 110.960 41.910 ;
        RECT 111.500 41.860 111.930 41.980 ;
        RECT 111.730 41.830 111.930 41.860 ;
        RECT 110.410 41.680 110.960 41.790 ;
        RECT 110.410 41.620 110.950 41.680 ;
        RECT 110.100 41.570 110.290 41.600 ;
        RECT 110.080 41.560 110.290 41.570 ;
        RECT 109.090 41.440 109.410 41.480 ;
        RECT 78.850 41.120 79.190 41.290 ;
        RECT 80.210 41.120 80.540 41.290 ;
        RECT 80.140 40.730 80.310 40.780 ;
        RECT 54.220 40.090 54.550 40.350 ;
        RECT 54.810 40.330 55.140 40.500 ;
        RECT 56.160 40.330 56.510 40.500 ;
        RECT 54.220 39.520 54.390 40.090 ;
        RECT 59.460 39.710 59.690 40.440 ;
        RECT 60.650 39.820 60.820 40.240 ;
        RECT 61.460 40.120 61.700 40.150 ;
        RECT 61.130 39.950 61.700 40.120 ;
        RECT 61.940 39.950 63.280 40.120 ;
        RECT 63.730 39.950 64.690 40.120 ;
        RECT 61.460 39.910 61.700 39.950 ;
        RECT 64.240 39.940 64.410 39.950 ;
        RECT 54.810 39.540 55.140 39.710 ;
        RECT 56.160 39.540 56.510 39.710 ;
        RECT 60.580 39.600 60.750 39.640 ;
        RECT 60.520 39.500 60.750 39.600 ;
        RECT 61.500 39.580 61.840 39.830 ;
        RECT 60.920 39.500 61.110 39.520 ;
        RECT 61.500 39.500 61.850 39.580 ;
        RECT 63.920 39.500 64.250 39.680 ;
        RECT 52.620 39.230 52.830 39.260 ;
        RECT 52.630 38.880 52.830 39.230 ;
        RECT 54.110 38.960 54.640 39.130 ;
        RECT 45.490 38.660 46.130 38.680 ;
        RECT 45.950 38.650 46.130 38.660 ;
        RECT 47.730 38.650 48.330 38.800 ;
        RECT 45.950 38.630 48.330 38.650 ;
        RECT 48.790 38.640 49.120 38.810 ;
        RECT 56.800 38.650 61.850 39.500 ;
        RECT 61.940 39.330 64.690 39.500 ;
        RECT 65.220 39.260 65.390 40.190 ;
        RECT 65.620 39.390 65.790 40.240 ;
        RECT 75.660 39.710 75.890 40.440 ;
        RECT 78.840 40.330 79.190 40.500 ;
        RECT 80.140 40.470 80.700 40.730 ;
        RECT 80.140 40.450 80.540 40.470 ;
        RECT 80.210 40.330 80.540 40.450 ;
        RECT 80.960 40.350 81.130 41.210 ;
        RECT 81.790 41.120 81.970 41.310 ;
        RECT 109.090 41.250 109.420 41.440 ;
        RECT 109.680 41.390 110.290 41.560 ;
        RECT 109.090 41.220 109.410 41.250 ;
        RECT 81.790 40.490 81.960 41.120 ;
        RECT 109.090 40.920 109.410 40.950 ;
        RECT 81.610 40.450 81.960 40.490 ;
        RECT 78.840 39.540 79.190 39.710 ;
        RECT 79.560 39.370 79.740 40.300 ;
        RECT 80.290 40.040 80.620 40.210 ;
        RECT 80.800 40.090 81.130 40.350 ;
        RECT 81.380 40.190 81.960 40.450 ;
        RECT 82.150 40.490 82.390 40.640 ;
        RECT 107.870 40.580 108.040 40.860 ;
        RECT 109.090 40.730 109.420 40.920 ;
        RECT 109.680 40.780 109.860 41.390 ;
        RECT 110.100 41.370 110.290 41.390 ;
        RECT 110.490 41.480 110.660 41.620 ;
        RECT 110.720 41.480 110.890 41.620 ;
        RECT 111.230 41.560 111.420 41.590 ;
        RECT 110.490 41.440 110.980 41.480 ;
        RECT 111.230 41.470 111.670 41.560 ;
        RECT 111.730 41.470 111.930 41.500 ;
        RECT 110.490 41.250 110.990 41.440 ;
        RECT 111.230 41.360 111.930 41.470 ;
        RECT 110.490 41.220 110.980 41.250 ;
        RECT 110.490 40.950 110.660 41.220 ;
        RECT 111.320 41.210 111.930 41.360 ;
        RECT 111.950 41.300 112.120 41.980 ;
        RECT 111.320 41.180 111.490 41.210 ;
        RECT 111.730 41.170 111.930 41.210 ;
        RECT 112.320 41.170 112.870 42.160 ;
        RECT 113.790 42.150 114.110 42.190 ;
        RECT 113.330 41.970 114.120 42.150 ;
        RECT 113.790 41.960 114.120 41.970 ;
        RECT 113.790 41.930 114.110 41.960 ;
        RECT 113.340 41.210 114.040 41.550 ;
        RECT 113.190 40.980 114.040 41.210 ;
        RECT 110.490 40.920 110.980 40.950 ;
        RECT 110.100 40.780 110.290 40.800 ;
        RECT 109.090 40.690 109.410 40.730 ;
        RECT 107.870 40.540 108.080 40.580 ;
        RECT 82.150 40.310 82.750 40.490 ;
        RECT 81.610 40.160 81.960 40.190 ;
        RECT 80.370 39.900 80.620 40.040 ;
        RECT 80.370 39.710 80.850 39.900 ;
        RECT 80.210 39.640 80.850 39.710 ;
        RECT 80.210 39.540 80.540 39.640 ;
        RECT 79.440 39.340 79.760 39.370 ;
        RECT 79.440 39.150 79.770 39.340 ;
        RECT 79.440 39.110 79.760 39.150 ;
        RECT 45.950 38.480 48.180 38.630 ;
        RECT 60.580 38.490 60.750 38.650 ;
        RECT 60.520 38.320 60.750 38.490 ;
        RECT 60.920 38.590 61.110 38.630 ;
        RECT 60.920 38.420 61.480 38.590 ;
        RECT 61.940 38.420 64.690 38.590 ;
        RECT 60.920 38.400 61.110 38.420 ;
        RECT 60.580 38.280 60.750 38.320 ;
        RECT 63.920 38.240 64.250 38.420 ;
        RECT 40.880 38.140 41.050 38.190 ;
        RECT 40.850 37.920 41.070 38.140 ;
        RECT 40.880 37.860 41.050 37.920 ;
        RECT 41.400 37.780 41.730 37.960 ;
        RECT 44.540 37.950 44.710 38.000 ;
        RECT 41.980 37.780 44.140 37.950 ;
        RECT 44.380 37.780 44.710 37.950 ;
        RECT 45.000 37.810 45.210 38.140 ;
        RECT 41.430 37.340 41.700 37.780 ;
        RECT 42.910 37.520 43.240 37.780 ;
        RECT 44.450 37.640 44.710 37.780 ;
        RECT 45.450 37.640 45.630 38.080 ;
        RECT 46.180 37.870 47.540 37.980 ;
        RECT 46.180 37.810 47.620 37.870 ;
        RECT 46.980 37.800 47.620 37.810 ;
        RECT 41.470 37.330 41.700 37.340 ;
        RECT 44.450 37.470 45.630 37.640 ;
        RECT 47.150 37.700 47.620 37.800 ;
        RECT 48.090 37.720 49.050 37.890 ;
        RECT 44.450 37.330 44.710 37.470 ;
        RECT 47.150 37.450 47.400 37.700 ;
        RECT 41.470 37.160 42.230 37.330 ;
        RECT 42.480 37.160 43.650 37.330 ;
        RECT 43.890 37.300 44.710 37.330 ;
        RECT 45.950 37.300 46.130 37.360 ;
        RECT 43.890 37.160 45.000 37.300 ;
        RECT 42.880 37.060 43.230 37.160 ;
        RECT 44.540 37.130 45.000 37.160 ;
        RECT 45.450 37.130 46.130 37.300 ;
        RECT 47.070 37.280 47.400 37.450 ;
        RECT 48.870 37.260 49.050 37.720 ;
        RECT 60.650 37.680 60.820 38.100 ;
        RECT 61.460 37.970 61.700 38.010 ;
        RECT 64.240 37.970 64.410 37.980 ;
        RECT 64.690 37.970 64.890 38.210 ;
        RECT 61.130 37.800 61.700 37.970 ;
        RECT 61.940 37.800 63.280 37.970 ;
        RECT 63.730 37.800 64.890 37.970 ;
        RECT 61.460 37.770 61.700 37.800 ;
        RECT 45.490 37.110 46.130 37.130 ;
        RECT 45.950 37.100 46.130 37.110 ;
        RECT 47.730 37.100 48.330 37.250 ;
        RECT 45.950 37.080 48.330 37.100 ;
        RECT 48.790 37.090 49.120 37.260 ;
        RECT 64.690 37.200 64.890 37.800 ;
        RECT 65.220 37.730 65.390 38.660 ;
        RECT 65.620 37.680 65.790 38.530 ;
        RECT 70.440 37.200 70.730 38.210 ;
        RECT 45.950 36.930 48.180 37.080 ;
        RECT 68.080 36.610 68.280 36.960 ;
        RECT 69.820 36.880 70.140 36.890 ;
        RECT 69.560 36.710 70.140 36.880 ;
        RECT 69.810 36.660 70.140 36.710 ;
        RECT 69.820 36.630 70.140 36.660 ;
        RECT 68.070 36.580 68.280 36.610 ;
        RECT 68.070 35.990 68.290 36.580 ;
        RECT 68.810 36.020 69.010 36.590 ;
        RECT 69.820 36.300 70.140 36.340 ;
        RECT 69.810 36.260 70.140 36.300 ;
        RECT 69.560 36.090 70.140 36.260 ;
        RECT 69.820 36.080 70.140 36.090 ;
        RECT 68.070 34.960 68.290 35.550 ;
        RECT 70.820 35.530 70.990 36.040 ;
        RECT 74.760 35.540 74.930 36.050 ;
        RECT 68.070 34.930 68.280 34.960 ;
        RECT 68.810 34.950 69.010 35.520 ;
        RECT 69.820 35.450 70.140 35.460 ;
        RECT 69.560 35.280 70.140 35.450 ;
        RECT 69.810 35.240 70.140 35.280 ;
        RECT 69.820 35.200 70.140 35.240 ;
        RECT 79.560 35.200 79.740 39.110 ;
        RECT 80.370 38.260 80.540 39.540 ;
        RECT 80.960 39.520 81.130 40.090 ;
        RECT 81.200 39.800 81.370 39.840 ;
        RECT 81.790 39.830 81.960 40.160 ;
        RECT 82.160 40.010 82.750 40.310 ;
        RECT 83.570 40.370 84.150 40.540 ;
        RECT 107.870 40.520 108.100 40.540 ;
        RECT 109.220 40.530 109.390 40.690 ;
        RECT 109.680 40.610 110.290 40.780 ;
        RECT 107.870 40.500 108.130 40.520 ;
        RECT 107.870 40.450 108.210 40.500 ;
        RECT 107.870 40.390 108.360 40.450 ;
        RECT 83.570 40.270 83.960 40.370 ;
        RECT 107.870 40.360 108.380 40.390 ;
        RECT 107.910 40.330 108.380 40.360 ;
        RECT 108.040 40.280 108.380 40.330 ;
        RECT 109.680 40.280 109.860 40.610 ;
        RECT 110.080 40.600 110.290 40.610 ;
        RECT 110.100 40.570 110.290 40.600 ;
        RECT 110.490 40.730 110.990 40.920 ;
        RECT 111.230 40.780 111.420 40.810 ;
        RECT 110.490 40.690 110.980 40.730 ;
        RECT 108.160 40.270 108.380 40.280 ;
        RECT 83.570 40.240 83.950 40.270 ;
        RECT 108.170 40.240 108.380 40.270 ;
        RECT 83.570 40.090 83.930 40.240 ;
        RECT 108.190 40.160 108.380 40.240 ;
        RECT 109.550 40.160 109.880 40.280 ;
        RECT 110.490 40.160 110.660 40.690 ;
        RECT 110.720 40.530 110.890 40.690 ;
        RECT 111.230 40.640 111.670 40.780 ;
        RECT 111.730 40.640 111.930 40.680 ;
        RECT 111.230 40.580 111.930 40.640 ;
        RECT 111.320 40.380 111.930 40.580 ;
        RECT 111.320 40.340 111.490 40.380 ;
        RECT 111.730 40.350 111.930 40.380 ;
        RECT 111.950 40.190 112.120 40.870 ;
        RECT 107.700 40.110 107.870 40.130 ;
        RECT 81.610 39.800 81.960 39.830 ;
        RECT 81.200 39.540 81.960 39.800 ;
        RECT 81.200 39.510 81.370 39.540 ;
        RECT 81.610 39.510 81.960 39.540 ;
        RECT 81.610 39.500 81.810 39.510 ;
        RECT 82.200 39.500 82.750 40.010 ;
        RECT 83.220 39.920 83.930 40.090 ;
        RECT 107.680 39.680 107.890 40.110 ;
        RECT 108.190 39.990 108.710 40.160 ;
        RECT 108.190 39.960 108.380 39.990 ;
        RECT 109.060 39.980 110.960 40.160 ;
        RECT 111.690 40.150 112.120 40.190 ;
        RECT 111.340 39.990 112.120 40.150 ;
        RECT 111.340 39.980 111.930 39.990 ;
        RECT 109.680 39.830 109.860 39.980 ;
        RECT 110.490 39.840 110.660 39.980 ;
        RECT 111.500 39.730 111.930 39.980 ;
        RECT 111.730 39.690 111.930 39.730 ;
        RECT 112.320 39.690 112.870 40.680 ;
        RECT 113.340 40.670 114.040 40.980 ;
        RECT 113.340 40.060 114.050 40.230 ;
        RECT 113.690 39.780 114.050 40.060 ;
        RECT 113.690 39.610 114.270 39.780 ;
        RECT 82.510 39.260 82.730 39.500 ;
        RECT 82.520 39.230 82.730 39.260 ;
        RECT 80.710 39.000 81.240 39.130 ;
        RECT 82.520 39.010 82.720 39.230 ;
        RECT 83.220 39.170 83.920 39.480 ;
        RECT 80.710 38.970 81.370 39.000 ;
        RECT 81.610 38.970 81.810 39.010 ;
        RECT 80.710 38.960 81.810 38.970 ;
        RECT 81.200 38.710 81.810 38.960 ;
        RECT 81.200 38.670 81.370 38.710 ;
        RECT 81.610 38.680 81.810 38.710 ;
        RECT 81.610 38.320 81.810 38.350 ;
        RECT 80.170 38.060 80.490 38.090 ;
        RECT 81.380 38.060 81.810 38.320 ;
        RECT 80.170 37.870 80.500 38.060 ;
        RECT 81.610 38.020 81.810 38.060 ;
        RECT 82.200 38.020 82.750 39.010 ;
        RECT 83.070 38.940 83.920 39.170 ;
        RECT 107.680 39.040 107.890 39.470 ;
        RECT 108.190 39.160 108.380 39.190 ;
        RECT 111.690 39.170 111.880 39.190 ;
        RECT 107.700 39.020 107.870 39.040 ;
        RECT 83.220 38.600 83.920 38.940 ;
        RECT 108.190 38.990 108.710 39.160 ;
        RECT 109.060 38.990 110.960 39.170 ;
        RECT 111.340 39.160 111.880 39.170 ;
        RECT 111.340 39.000 112.120 39.160 ;
        RECT 108.190 38.910 108.380 38.990 ;
        RECT 108.170 38.880 108.380 38.910 ;
        RECT 108.160 38.870 108.380 38.880 ;
        RECT 109.550 38.870 109.880 38.990 ;
        RECT 111.690 38.960 112.120 39.000 ;
        RECT 108.040 38.820 108.380 38.870 ;
        RECT 107.910 38.790 108.380 38.820 ;
        RECT 107.870 38.760 108.380 38.790 ;
        RECT 107.870 38.700 108.360 38.760 ;
        RECT 107.870 38.650 108.210 38.700 ;
        RECT 107.870 38.630 108.130 38.650 ;
        RECT 107.870 38.610 108.100 38.630 ;
        RECT 107.870 38.570 108.080 38.610 ;
        RECT 107.870 38.290 108.040 38.570 ;
        RECT 109.220 38.460 109.390 38.620 ;
        RECT 110.100 38.550 110.290 38.580 ;
        RECT 110.080 38.540 110.290 38.550 ;
        RECT 109.090 38.420 109.410 38.460 ;
        RECT 83.680 38.240 84.000 38.280 ;
        RECT 83.680 38.180 84.010 38.240 ;
        RECT 109.090 38.230 109.420 38.420 ;
        RECT 109.830 38.370 110.290 38.540 ;
        RECT 110.720 38.460 110.890 38.620 ;
        RECT 111.230 38.540 111.420 38.570 ;
        RECT 110.100 38.350 110.290 38.370 ;
        RECT 110.660 38.420 110.980 38.460 ;
        RECT 110.660 38.230 110.990 38.420 ;
        RECT 111.230 38.370 111.670 38.540 ;
        RECT 111.230 38.340 111.420 38.370 ;
        RECT 111.950 38.280 112.120 38.960 ;
        RECT 109.090 38.200 109.410 38.230 ;
        RECT 110.660 38.200 110.980 38.230 ;
        RECT 83.210 38.050 84.010 38.180 ;
        RECT 83.210 38.020 84.000 38.050 ;
        RECT 83.210 38.000 83.910 38.020 ;
        RECT 80.170 37.830 80.490 37.870 ;
        RECT 80.170 37.750 80.340 37.830 ;
        RECT 80.120 37.580 80.340 37.750 ;
        RECT 80.120 37.420 80.290 37.580 ;
        RECT 81.610 37.490 81.810 37.530 ;
        RECT 80.650 37.160 80.840 37.280 ;
        RECT 81.380 37.230 81.810 37.490 ;
        RECT 81.610 37.200 81.810 37.230 ;
        RECT 80.290 37.050 80.840 37.160 ;
        RECT 80.290 36.990 80.830 37.050 ;
        RECT 80.370 35.210 80.540 36.990 ;
        RECT 81.200 36.840 81.370 36.880 ;
        RECT 81.610 36.840 81.810 36.870 ;
        RECT 81.200 36.580 81.810 36.840 ;
        RECT 81.200 36.550 81.370 36.580 ;
        RECT 81.610 36.540 81.810 36.580 ;
        RECT 82.200 36.540 82.750 37.530 ;
        RECT 83.670 37.520 83.990 37.560 ;
        RECT 83.210 37.340 84.000 37.520 ;
        RECT 83.670 37.330 84.000 37.340 ;
        RECT 83.670 37.300 83.990 37.330 ;
        RECT 83.220 36.580 83.920 36.920 ;
        RECT 90.620 36.880 90.940 36.890 ;
        RECT 90.620 36.710 91.200 36.880 ;
        RECT 90.620 36.660 90.950 36.710 ;
        RECT 90.620 36.630 90.940 36.660 ;
        RECT 92.480 36.610 92.680 36.960 ;
        RECT 83.070 36.350 83.920 36.580 ;
        RECT 81.200 36.010 81.370 36.040 ;
        RECT 81.610 36.010 81.810 36.050 ;
        RECT 81.200 35.750 81.810 36.010 ;
        RECT 81.200 35.710 81.370 35.750 ;
        RECT 81.610 35.720 81.810 35.750 ;
        RECT 81.610 35.360 81.810 35.390 ;
        RECT 81.380 35.100 81.810 35.360 ;
        RECT 81.610 35.060 81.810 35.100 ;
        RECT 82.200 35.060 82.750 36.050 ;
        RECT 83.220 36.040 83.920 36.350 ;
        RECT 90.620 36.300 90.940 36.340 ;
        RECT 90.620 36.260 90.950 36.300 ;
        RECT 90.620 36.090 91.200 36.260 ;
        RECT 90.620 36.080 90.940 36.090 ;
        RECT 83.220 35.430 83.930 35.600 ;
        RECT 85.830 35.540 86.000 36.050 ;
        RECT 89.770 35.530 89.940 36.040 ;
        RECT 91.750 36.020 91.950 36.590 ;
        RECT 92.480 36.580 92.690 36.610 ;
        RECT 92.470 35.990 92.690 36.580 ;
        RECT 83.570 35.150 83.930 35.430 ;
        RECT 90.620 35.450 90.940 35.460 ;
        RECT 90.620 35.280 91.200 35.450 ;
        RECT 90.620 35.240 90.950 35.280 ;
        RECT 90.620 35.200 90.940 35.240 ;
        RECT 83.570 34.980 84.150 35.150 ;
        RECT 91.750 34.950 91.950 35.520 ;
        RECT 92.470 34.960 92.690 35.550 ;
        RECT 68.080 34.580 68.280 34.930 ;
        RECT 92.480 34.930 92.690 34.960 ;
        RECT 69.820 34.880 70.140 34.910 ;
        RECT 69.810 34.830 70.140 34.880 ;
        RECT 90.620 34.880 90.940 34.910 ;
        RECT 69.560 34.660 70.140 34.830 ;
        RECT 69.820 34.650 70.140 34.660 ;
        RECT 68.450 34.180 68.890 34.350 ;
        RECT 68.080 33.600 68.280 33.950 ;
        RECT 69.820 33.870 70.140 33.880 ;
        RECT 69.560 33.700 70.140 33.870 ;
        RECT 69.810 33.650 70.140 33.700 ;
        RECT 70.820 33.690 70.990 34.700 ;
        RECT 72.750 33.970 73.300 34.400 ;
        RECT 74.750 33.830 74.920 34.840 ;
        RECT 76.780 34.040 77.330 34.470 ;
        RECT 83.430 34.040 83.980 34.470 ;
        RECT 85.840 33.830 86.010 34.840 ;
        RECT 90.620 34.830 90.950 34.880 ;
        RECT 87.460 33.970 88.010 34.400 ;
        RECT 89.770 33.690 89.940 34.700 ;
        RECT 90.620 34.660 91.200 34.830 ;
        RECT 90.620 34.650 90.940 34.660 ;
        RECT 92.480 34.580 92.680 34.930 ;
        RECT 91.870 34.180 92.310 34.350 ;
        RECT 90.620 33.870 90.940 33.880 ;
        RECT 90.620 33.700 91.200 33.870 ;
        RECT 69.820 33.620 70.140 33.650 ;
        RECT 90.620 33.650 90.950 33.700 ;
        RECT 90.620 33.620 90.940 33.650 ;
        RECT 68.070 33.570 68.280 33.600 ;
        RECT 92.480 33.600 92.680 33.950 ;
        RECT 40.880 32.660 41.050 32.710 ;
        RECT 60.650 32.680 60.820 33.100 ;
        RECT 61.460 32.980 61.700 33.010 ;
        RECT 61.130 32.810 61.700 32.980 ;
        RECT 61.940 32.810 63.280 32.980 ;
        RECT 63.730 32.810 64.690 32.980 ;
        RECT 61.460 32.770 61.700 32.810 ;
        RECT 64.240 32.800 64.410 32.810 ;
        RECT 40.850 32.440 41.070 32.660 ;
        RECT 40.880 32.380 41.050 32.440 ;
        RECT 41.400 32.300 41.730 32.480 ;
        RECT 44.540 32.470 44.710 32.520 ;
        RECT 41.980 32.300 44.140 32.470 ;
        RECT 44.380 32.300 44.710 32.470 ;
        RECT 45.000 32.330 45.210 32.660 ;
        RECT 41.430 31.860 41.700 32.300 ;
        RECT 42.910 32.040 43.240 32.300 ;
        RECT 44.450 32.160 44.710 32.300 ;
        RECT 45.450 32.160 45.630 32.600 ;
        RECT 46.180 32.390 47.540 32.500 ;
        RECT 60.580 32.460 60.750 32.500 ;
        RECT 46.180 32.330 47.620 32.390 ;
        RECT 46.980 32.320 47.620 32.330 ;
        RECT 41.470 31.850 41.700 31.860 ;
        RECT 44.450 31.990 45.630 32.160 ;
        RECT 47.150 32.220 47.620 32.320 ;
        RECT 48.090 32.240 49.050 32.410 ;
        RECT 60.520 32.290 60.750 32.460 ;
        RECT 44.450 31.850 44.710 31.990 ;
        RECT 47.150 31.970 47.400 32.220 ;
        RECT 41.470 31.680 42.230 31.850 ;
        RECT 42.480 31.680 43.650 31.850 ;
        RECT 43.890 31.820 44.710 31.850 ;
        RECT 45.950 31.820 46.130 31.880 ;
        RECT 43.890 31.680 45.000 31.820 ;
        RECT 42.880 31.580 43.230 31.680 ;
        RECT 44.540 31.650 45.000 31.680 ;
        RECT 45.450 31.650 46.130 31.820 ;
        RECT 47.070 31.800 47.400 31.970 ;
        RECT 48.870 31.780 49.050 32.240 ;
        RECT 60.580 31.940 60.750 32.290 ;
        RECT 60.920 32.360 61.110 32.380 ;
        RECT 63.920 32.360 64.250 32.540 ;
        RECT 60.920 32.190 61.480 32.360 ;
        RECT 61.940 32.190 64.690 32.360 ;
        RECT 60.920 32.150 61.110 32.190 ;
        RECT 65.220 32.120 65.390 33.050 ;
        RECT 65.620 32.250 65.790 33.100 ;
        RECT 68.070 32.980 68.290 33.570 ;
        RECT 68.810 33.010 69.010 33.580 ;
        RECT 69.820 33.290 70.140 33.330 ;
        RECT 69.810 33.250 70.140 33.290 ;
        RECT 69.560 33.080 70.140 33.250 ;
        RECT 69.820 33.070 70.140 33.080 ;
        RECT 90.620 33.290 90.940 33.330 ;
        RECT 90.620 33.250 90.950 33.290 ;
        RECT 90.620 33.080 91.200 33.250 ;
        RECT 90.620 33.070 90.940 33.080 ;
        RECT 91.750 33.010 91.950 33.580 ;
        RECT 92.480 33.570 92.690 33.600 ;
        RECT 92.470 32.980 92.690 33.570 ;
        RECT 68.070 31.960 68.290 32.550 ;
        RECT 68.070 31.930 68.280 31.960 ;
        RECT 68.810 31.950 69.010 32.520 ;
        RECT 69.820 32.450 70.140 32.460 ;
        RECT 69.560 32.280 70.140 32.450 ;
        RECT 69.810 32.240 70.140 32.280 ;
        RECT 69.820 32.200 70.140 32.240 ;
        RECT 90.620 32.450 90.940 32.460 ;
        RECT 90.620 32.280 91.200 32.450 ;
        RECT 90.620 32.240 90.950 32.280 ;
        RECT 90.620 32.200 90.940 32.240 ;
        RECT 91.750 31.950 91.950 32.520 ;
        RECT 92.470 31.960 92.690 32.550 ;
        RECT 45.490 31.630 46.130 31.650 ;
        RECT 45.950 31.620 46.130 31.630 ;
        RECT 47.730 31.620 48.330 31.770 ;
        RECT 45.950 31.600 48.330 31.620 ;
        RECT 48.790 31.610 49.120 31.780 ;
        RECT 45.950 31.450 48.180 31.600 ;
        RECT 60.580 31.350 60.750 31.700 ;
        RECT 68.080 31.580 68.280 31.930 ;
        RECT 92.480 31.930 92.690 31.960 ;
        RECT 69.820 31.880 70.140 31.910 ;
        RECT 69.810 31.830 70.140 31.880 ;
        RECT 69.560 31.660 70.140 31.830 ;
        RECT 69.820 31.650 70.140 31.660 ;
        RECT 90.620 31.880 90.940 31.910 ;
        RECT 90.620 31.830 90.950 31.880 ;
        RECT 90.620 31.660 91.200 31.830 ;
        RECT 90.620 31.650 90.940 31.660 ;
        RECT 92.480 31.580 92.680 31.930 ;
        RECT 60.520 31.180 60.750 31.350 ;
        RECT 60.920 31.450 61.110 31.490 ;
        RECT 60.920 31.280 61.480 31.450 ;
        RECT 61.940 31.280 64.690 31.450 ;
        RECT 60.920 31.260 61.110 31.280 ;
        RECT 40.880 31.110 41.050 31.160 ;
        RECT 60.580 31.140 60.750 31.180 ;
        RECT 40.850 30.890 41.070 31.110 ;
        RECT 40.880 30.830 41.050 30.890 ;
        RECT 41.400 30.750 41.730 30.930 ;
        RECT 44.540 30.920 44.710 30.970 ;
        RECT 41.980 30.750 44.140 30.920 ;
        RECT 44.380 30.750 44.710 30.920 ;
        RECT 45.000 30.780 45.210 31.110 ;
        RECT 63.920 31.100 64.250 31.280 ;
        RECT 41.430 30.310 41.700 30.750 ;
        RECT 42.910 30.490 43.240 30.750 ;
        RECT 44.450 30.610 44.710 30.750 ;
        RECT 45.450 30.610 45.630 31.050 ;
        RECT 46.180 30.840 47.540 30.950 ;
        RECT 46.180 30.780 47.620 30.840 ;
        RECT 46.980 30.770 47.620 30.780 ;
        RECT 41.470 30.300 41.700 30.310 ;
        RECT 44.450 30.440 45.630 30.610 ;
        RECT 47.150 30.670 47.620 30.770 ;
        RECT 48.090 30.690 49.050 30.860 ;
        RECT 44.450 30.300 44.710 30.440 ;
        RECT 47.150 30.420 47.400 30.670 ;
        RECT 41.470 30.130 42.230 30.300 ;
        RECT 42.480 30.130 43.650 30.300 ;
        RECT 43.890 30.270 44.710 30.300 ;
        RECT 45.950 30.270 46.130 30.330 ;
        RECT 43.890 30.130 45.000 30.270 ;
        RECT 42.880 30.030 43.230 30.130 ;
        RECT 44.540 30.100 45.000 30.130 ;
        RECT 45.450 30.100 46.130 30.270 ;
        RECT 47.070 30.250 47.400 30.420 ;
        RECT 48.870 30.230 49.050 30.690 ;
        RECT 60.650 30.540 60.820 30.960 ;
        RECT 61.460 30.830 61.700 30.870 ;
        RECT 64.240 30.830 64.410 30.840 ;
        RECT 61.130 30.660 61.700 30.830 ;
        RECT 61.940 30.660 63.280 30.830 ;
        RECT 63.730 30.660 64.690 30.830 ;
        RECT 61.460 30.630 61.700 30.660 ;
        RECT 65.220 30.590 65.390 31.520 ;
        RECT 65.620 30.540 65.790 31.390 ;
        RECT 45.490 30.080 46.130 30.100 ;
        RECT 45.950 30.070 46.130 30.080 ;
        RECT 47.730 30.070 48.330 30.220 ;
        RECT 45.950 30.050 48.330 30.070 ;
        RECT 48.790 30.060 49.120 30.230 ;
        RECT 45.950 29.900 48.180 30.050 ;
        RECT 60.650 29.750 60.820 30.170 ;
        RECT 61.460 30.050 61.700 30.080 ;
        RECT 61.130 29.880 61.700 30.050 ;
        RECT 61.940 29.880 63.280 30.050 ;
        RECT 63.730 29.880 64.690 30.050 ;
        RECT 61.460 29.840 61.700 29.880 ;
        RECT 64.240 29.870 64.410 29.880 ;
        RECT 40.880 29.560 41.050 29.610 ;
        RECT 40.850 29.340 41.070 29.560 ;
        RECT 40.880 29.280 41.050 29.340 ;
        RECT 41.400 29.200 41.730 29.380 ;
        RECT 44.540 29.370 44.710 29.420 ;
        RECT 41.980 29.200 44.140 29.370 ;
        RECT 44.380 29.200 44.710 29.370 ;
        RECT 45.000 29.230 45.210 29.560 ;
        RECT 60.580 29.530 60.750 29.570 ;
        RECT 41.430 28.760 41.700 29.200 ;
        RECT 42.910 28.940 43.240 29.200 ;
        RECT 44.450 29.060 44.710 29.200 ;
        RECT 45.450 29.060 45.630 29.500 ;
        RECT 46.180 29.290 47.540 29.400 ;
        RECT 60.520 29.360 60.750 29.530 ;
        RECT 46.180 29.230 47.620 29.290 ;
        RECT 46.980 29.220 47.620 29.230 ;
        RECT 41.470 28.750 41.700 28.760 ;
        RECT 44.450 28.890 45.630 29.060 ;
        RECT 47.150 29.120 47.620 29.220 ;
        RECT 48.090 29.140 49.050 29.310 ;
        RECT 44.450 28.750 44.710 28.890 ;
        RECT 47.150 28.870 47.400 29.120 ;
        RECT 41.470 28.580 42.230 28.750 ;
        RECT 42.480 28.580 43.650 28.750 ;
        RECT 43.890 28.720 44.710 28.750 ;
        RECT 45.950 28.720 46.130 28.780 ;
        RECT 43.890 28.580 45.000 28.720 ;
        RECT 42.880 28.480 43.230 28.580 ;
        RECT 44.540 28.550 45.000 28.580 ;
        RECT 45.450 28.550 46.130 28.720 ;
        RECT 47.070 28.700 47.400 28.870 ;
        RECT 48.870 28.680 49.050 29.140 ;
        RECT 60.580 29.010 60.750 29.360 ;
        RECT 60.920 29.430 61.110 29.450 ;
        RECT 63.920 29.430 64.250 29.610 ;
        RECT 60.920 29.260 61.480 29.430 ;
        RECT 61.940 29.260 64.690 29.430 ;
        RECT 60.920 29.220 61.110 29.260 ;
        RECT 65.220 29.190 65.390 30.120 ;
        RECT 65.620 29.320 65.790 30.170 ;
        RECT 45.490 28.530 46.130 28.550 ;
        RECT 45.950 28.520 46.130 28.530 ;
        RECT 47.730 28.520 48.330 28.670 ;
        RECT 45.950 28.500 48.330 28.520 ;
        RECT 48.790 28.510 49.120 28.680 ;
        RECT 45.950 28.350 48.180 28.500 ;
        RECT 60.580 28.420 60.750 28.770 ;
        RECT 60.520 28.250 60.750 28.420 ;
        RECT 60.920 28.520 61.110 28.560 ;
        RECT 60.920 28.350 61.480 28.520 ;
        RECT 61.940 28.350 64.690 28.520 ;
        RECT 60.920 28.330 61.110 28.350 ;
        RECT 60.580 28.210 60.750 28.250 ;
        RECT 63.920 28.170 64.250 28.350 ;
        RECT 40.880 28.010 41.050 28.060 ;
        RECT 40.850 27.790 41.070 28.010 ;
        RECT 40.880 27.730 41.050 27.790 ;
        RECT 41.400 27.650 41.730 27.830 ;
        RECT 44.540 27.820 44.710 27.870 ;
        RECT 41.980 27.650 44.140 27.820 ;
        RECT 44.380 27.650 44.710 27.820 ;
        RECT 45.000 27.680 45.210 28.010 ;
        RECT 41.430 27.210 41.700 27.650 ;
        RECT 42.910 27.390 43.240 27.650 ;
        RECT 44.450 27.510 44.710 27.650 ;
        RECT 45.450 27.510 45.630 27.950 ;
        RECT 46.180 27.740 47.540 27.850 ;
        RECT 46.180 27.680 47.620 27.740 ;
        RECT 46.980 27.670 47.620 27.680 ;
        RECT 41.470 27.200 41.700 27.210 ;
        RECT 44.450 27.340 45.630 27.510 ;
        RECT 47.150 27.570 47.620 27.670 ;
        RECT 48.090 27.590 49.050 27.760 ;
        RECT 60.650 27.610 60.820 28.030 ;
        RECT 61.460 27.900 61.700 27.940 ;
        RECT 64.240 27.900 64.410 27.910 ;
        RECT 61.130 27.730 61.700 27.900 ;
        RECT 61.940 27.730 63.280 27.900 ;
        RECT 63.730 27.730 64.690 27.900 ;
        RECT 61.460 27.700 61.700 27.730 ;
        RECT 65.220 27.660 65.390 28.590 ;
        RECT 65.620 27.610 65.790 28.460 ;
        RECT 44.450 27.200 44.710 27.340 ;
        RECT 47.150 27.320 47.400 27.570 ;
        RECT 41.470 27.030 42.230 27.200 ;
        RECT 42.480 27.030 43.650 27.200 ;
        RECT 43.890 27.170 44.710 27.200 ;
        RECT 45.950 27.170 46.130 27.230 ;
        RECT 43.890 27.030 45.000 27.170 ;
        RECT 42.880 26.930 43.230 27.030 ;
        RECT 44.540 27.000 45.000 27.030 ;
        RECT 45.450 27.000 46.130 27.170 ;
        RECT 47.070 27.150 47.400 27.320 ;
        RECT 48.870 27.130 49.050 27.590 ;
        RECT 45.490 26.980 46.130 27.000 ;
        RECT 45.950 26.970 46.130 26.980 ;
        RECT 47.730 26.970 48.330 27.120 ;
        RECT 45.950 26.950 48.330 26.970 ;
        RECT 48.790 26.960 49.120 27.130 ;
        RECT 45.950 26.800 48.180 26.950 ;
        RECT 55.380 26.790 55.580 27.140 ;
        RECT 57.120 27.060 57.440 27.070 ;
        RECT 56.860 26.890 57.440 27.060 ;
        RECT 57.110 26.840 57.440 26.890 ;
        RECT 57.120 26.810 57.440 26.840 ;
        RECT 55.370 26.760 55.580 26.790 ;
        RECT 55.370 26.170 55.590 26.760 ;
        RECT 56.110 26.200 56.310 26.770 ;
        RECT 57.120 26.480 57.440 26.520 ;
        RECT 57.110 26.440 57.440 26.480 ;
        RECT 56.860 26.270 57.440 26.440 ;
        RECT 57.120 26.260 57.440 26.270 ;
        RECT 55.370 25.140 55.590 25.730 ;
        RECT 55.370 25.110 55.580 25.140 ;
        RECT 56.110 25.130 56.310 25.700 ;
        RECT 58.250 25.690 58.420 26.200 ;
        RECT 62.270 25.720 62.440 26.230 ;
        RECT 57.120 25.630 57.440 25.640 ;
        RECT 56.860 25.460 57.440 25.630 ;
        RECT 57.110 25.420 57.440 25.460 ;
        RECT 57.120 25.380 57.440 25.420 ;
        RECT 55.380 24.760 55.580 25.110 ;
        RECT 57.120 25.060 57.440 25.090 ;
        RECT 57.110 25.010 57.440 25.060 ;
        RECT 56.860 24.840 57.440 25.010 ;
        RECT 57.120 24.830 57.440 24.840 ;
        RECT 55.750 24.360 56.190 24.530 ;
        RECT 17.760 23.870 17.930 24.360 ;
        RECT 17.610 23.840 17.930 23.870 ;
        RECT 18.310 23.870 18.480 24.360 ;
        RECT 18.950 24.310 19.120 24.360 ;
        RECT 19.500 24.310 19.670 24.360 ;
        RECT 18.830 24.280 19.150 24.310 ;
        RECT 19.480 24.280 19.800 24.310 ;
        RECT 18.830 24.090 19.160 24.280 ;
        RECT 19.480 24.090 19.810 24.280 ;
        RECT 18.830 24.050 19.150 24.090 ;
        RECT 19.480 24.050 19.800 24.090 ;
        RECT 18.310 23.840 18.630 23.870 ;
        RECT 17.610 23.650 17.940 23.840 ;
        RECT 18.310 23.650 18.640 23.840 ;
        RECT 17.610 23.610 17.930 23.650 ;
        RECT 17.220 22.150 17.390 22.170 ;
        RECT 17.200 21.720 17.410 22.150 ;
        RECT 17.760 21.960 17.930 23.610 ;
        RECT 18.310 23.610 18.630 23.650 ;
        RECT 18.310 21.960 18.480 23.610 ;
        RECT 18.950 21.960 19.120 24.050 ;
        RECT 19.500 21.960 19.670 24.050 ;
        RECT 55.380 23.780 55.580 24.130 ;
        RECT 57.120 24.050 57.440 24.060 ;
        RECT 56.860 23.880 57.440 24.050 ;
        RECT 57.110 23.830 57.440 23.880 ;
        RECT 58.240 23.830 58.410 25.020 ;
        RECT 60.050 24.150 60.600 24.580 ;
        RECT 57.120 23.800 57.440 23.830 ;
        RECT 55.370 23.750 55.580 23.780 ;
        RECT 62.260 23.770 62.430 24.960 ;
        RECT 64.080 24.220 64.630 24.650 ;
        RECT 20.050 22.600 20.220 23.450 ;
        RECT 55.370 23.160 55.590 23.750 ;
        RECT 56.110 23.190 56.310 23.760 ;
        RECT 57.120 23.470 57.440 23.510 ;
        RECT 57.110 23.430 57.440 23.470 ;
        RECT 56.860 23.260 57.440 23.430 ;
        RECT 57.120 23.250 57.440 23.260 ;
        RECT 40.880 22.890 41.050 22.940 ;
        RECT 60.650 22.920 60.820 23.340 ;
        RECT 61.460 23.220 61.700 23.250 ;
        RECT 61.130 23.050 61.700 23.220 ;
        RECT 61.940 23.050 63.280 23.220 ;
        RECT 63.730 23.050 64.690 23.220 ;
        RECT 61.460 23.010 61.700 23.050 ;
        RECT 64.240 23.040 64.410 23.050 ;
        RECT 40.850 22.670 41.070 22.890 ;
        RECT 40.880 22.610 41.050 22.670 ;
        RECT 41.400 22.530 41.730 22.710 ;
        RECT 44.540 22.700 44.710 22.750 ;
        RECT 41.980 22.530 44.140 22.700 ;
        RECT 44.380 22.530 44.710 22.700 ;
        RECT 45.000 22.560 45.210 22.890 ;
        RECT 41.430 22.090 41.700 22.530 ;
        RECT 42.910 22.270 43.240 22.530 ;
        RECT 44.450 22.390 44.710 22.530 ;
        RECT 45.450 22.390 45.630 22.830 ;
        RECT 46.180 22.620 47.540 22.730 ;
        RECT 46.180 22.560 47.620 22.620 ;
        RECT 46.980 22.550 47.620 22.560 ;
        RECT 41.470 22.080 41.700 22.090 ;
        RECT 44.450 22.220 45.630 22.390 ;
        RECT 47.150 22.450 47.620 22.550 ;
        RECT 48.090 22.470 49.050 22.640 ;
        RECT 44.450 22.080 44.710 22.220 ;
        RECT 47.150 22.200 47.400 22.450 ;
        RECT 19.940 21.970 20.370 21.990 ;
        RECT 19.940 21.800 20.390 21.970 ;
        RECT 41.470 21.910 42.230 22.080 ;
        RECT 42.480 21.910 43.650 22.080 ;
        RECT 43.890 22.050 44.710 22.080 ;
        RECT 45.950 22.050 46.130 22.110 ;
        RECT 43.890 21.910 45.000 22.050 ;
        RECT 42.880 21.810 43.230 21.910 ;
        RECT 44.540 21.880 45.000 21.910 ;
        RECT 45.450 21.880 46.130 22.050 ;
        RECT 47.070 22.030 47.400 22.200 ;
        RECT 48.870 22.010 49.050 22.470 ;
        RECT 55.370 22.140 55.590 22.730 ;
        RECT 60.580 22.700 60.750 22.740 ;
        RECT 55.370 22.110 55.580 22.140 ;
        RECT 56.110 22.130 56.310 22.700 ;
        RECT 57.120 22.630 57.440 22.640 ;
        RECT 56.860 22.460 57.440 22.630 ;
        RECT 60.520 22.530 60.750 22.700 ;
        RECT 57.110 22.420 57.440 22.460 ;
        RECT 57.120 22.380 57.440 22.420 ;
        RECT 60.580 22.180 60.750 22.530 ;
        RECT 60.920 22.600 61.110 22.620 ;
        RECT 63.920 22.600 64.250 22.780 ;
        RECT 60.920 22.430 61.480 22.600 ;
        RECT 61.940 22.430 64.690 22.600 ;
        RECT 60.920 22.390 61.110 22.430 ;
        RECT 65.220 22.360 65.390 23.290 ;
        RECT 65.620 22.490 65.790 23.340 ;
        RECT 68.490 23.130 68.810 23.160 ;
        RECT 68.490 22.960 70.280 23.130 ;
        RECT 68.490 22.940 68.820 22.960 ;
        RECT 68.490 22.900 68.810 22.940 ;
        RECT 70.110 22.730 70.280 22.960 ;
        RECT 68.960 22.480 69.300 22.730 ;
        RECT 69.470 22.560 69.800 22.730 ;
        RECT 70.020 22.560 70.360 22.730 ;
        RECT 68.640 22.220 69.300 22.480 ;
        RECT 69.550 22.390 69.720 22.560 ;
        RECT 70.110 22.390 70.280 22.560 ;
        RECT 69.470 22.220 69.800 22.390 ;
        RECT 70.020 22.220 70.360 22.390 ;
        RECT 45.490 21.860 46.130 21.880 ;
        RECT 45.950 21.850 46.130 21.860 ;
        RECT 47.730 21.850 48.330 22.000 ;
        RECT 45.950 21.830 48.330 21.850 ;
        RECT 48.790 21.840 49.120 22.010 ;
        RECT 19.940 21.780 20.370 21.800 ;
        RECT 45.950 21.680 48.180 21.830 ;
        RECT 55.380 21.760 55.580 22.110 ;
        RECT 57.120 22.060 57.440 22.090 ;
        RECT 57.110 22.010 57.440 22.060 ;
        RECT 56.860 21.840 57.440 22.010 ;
        RECT 69.550 21.990 69.800 22.220 ;
        RECT 70.680 22.140 71.190 22.810 ;
        RECT 57.120 21.830 57.440 21.840 ;
        RECT 60.580 21.590 60.750 21.940 ;
        RECT 69.550 21.820 70.220 21.990 ;
        RECT 16.300 18.600 16.470 21.090 ;
        RECT 16.850 18.600 17.020 21.100 ;
        RECT 17.210 21.080 17.420 21.510 ;
        RECT 19.950 21.430 20.380 21.450 ;
        RECT 19.950 21.260 20.400 21.430 ;
        RECT 60.520 21.420 60.750 21.590 ;
        RECT 60.920 21.690 61.110 21.730 ;
        RECT 60.920 21.520 61.480 21.690 ;
        RECT 61.940 21.520 64.690 21.690 ;
        RECT 60.920 21.500 61.110 21.520 ;
        RECT 40.880 21.340 41.050 21.390 ;
        RECT 60.580 21.380 60.750 21.420 ;
        RECT 63.920 21.340 64.250 21.520 ;
        RECT 19.950 21.240 20.380 21.260 ;
        RECT 40.850 21.120 41.070 21.340 ;
        RECT 17.230 21.060 17.400 21.080 ;
        RECT 17.480 19.990 17.650 21.090 ;
        RECT 17.480 19.960 17.960 19.990 ;
        RECT 17.480 19.770 17.970 19.960 ;
        RECT 17.480 19.730 17.960 19.770 ;
        RECT 17.480 18.600 17.650 19.730 ;
        RECT 18.030 18.600 18.200 21.100 ;
        RECT 40.880 21.060 41.050 21.120 ;
        RECT 41.400 20.980 41.730 21.160 ;
        RECT 44.540 21.150 44.710 21.200 ;
        RECT 41.980 20.980 44.140 21.150 ;
        RECT 44.380 20.980 44.710 21.150 ;
        RECT 45.000 21.010 45.210 21.340 ;
        RECT 20.040 20.050 20.210 20.720 ;
        RECT 41.430 20.540 41.700 20.980 ;
        RECT 42.910 20.720 43.240 20.980 ;
        RECT 44.450 20.840 44.710 20.980 ;
        RECT 45.450 20.840 45.630 21.280 ;
        RECT 46.180 21.070 47.540 21.180 ;
        RECT 46.180 21.010 47.620 21.070 ;
        RECT 46.980 21.000 47.620 21.010 ;
        RECT 41.470 20.530 41.700 20.540 ;
        RECT 44.450 20.670 45.630 20.840 ;
        RECT 47.150 20.900 47.620 21.000 ;
        RECT 48.090 20.920 49.050 21.090 ;
        RECT 44.450 20.530 44.710 20.670 ;
        RECT 47.150 20.650 47.400 20.900 ;
        RECT 41.470 20.360 42.230 20.530 ;
        RECT 42.480 20.360 43.650 20.530 ;
        RECT 43.890 20.500 44.710 20.530 ;
        RECT 45.950 20.500 46.130 20.560 ;
        RECT 43.890 20.360 45.000 20.500 ;
        RECT 42.880 20.260 43.230 20.360 ;
        RECT 44.540 20.330 45.000 20.360 ;
        RECT 45.450 20.330 46.130 20.500 ;
        RECT 47.070 20.480 47.400 20.650 ;
        RECT 48.870 20.460 49.050 20.920 ;
        RECT 60.650 20.780 60.820 21.200 ;
        RECT 61.460 21.070 61.700 21.110 ;
        RECT 64.240 21.070 64.410 21.080 ;
        RECT 61.130 20.900 61.700 21.070 ;
        RECT 61.940 20.900 63.280 21.070 ;
        RECT 63.730 20.900 64.690 21.070 ;
        RECT 61.460 20.870 61.700 20.900 ;
        RECT 65.220 20.830 65.390 21.760 ;
        RECT 65.620 20.780 65.790 21.630 ;
        RECT 69.550 21.590 69.800 21.820 ;
        RECT 68.640 21.330 69.300 21.590 ;
        RECT 69.470 21.420 69.800 21.590 ;
        RECT 70.020 21.420 70.360 21.590 ;
        RECT 68.960 21.080 69.300 21.330 ;
        RECT 69.550 21.250 69.720 21.420 ;
        RECT 70.110 21.250 70.280 21.420 ;
        RECT 69.470 21.080 69.800 21.250 ;
        RECT 70.020 21.080 70.360 21.250 ;
        RECT 68.490 20.870 68.810 20.910 ;
        RECT 68.490 20.850 68.820 20.870 ;
        RECT 70.110 20.850 70.280 21.080 ;
        RECT 70.680 21.000 71.190 21.670 ;
        RECT 68.490 20.680 70.280 20.850 ;
        RECT 68.490 20.650 68.810 20.680 ;
        RECT 45.490 20.310 46.130 20.330 ;
        RECT 45.950 20.300 46.130 20.310 ;
        RECT 47.730 20.300 48.330 20.450 ;
        RECT 45.950 20.280 48.330 20.300 ;
        RECT 48.790 20.290 49.120 20.460 ;
        RECT 45.950 20.130 48.180 20.280 ;
        RECT 60.650 19.990 60.820 20.410 ;
        RECT 61.460 20.290 61.700 20.320 ;
        RECT 61.130 20.120 61.700 20.290 ;
        RECT 61.940 20.120 63.280 20.290 ;
        RECT 63.730 20.120 64.690 20.290 ;
        RECT 61.460 20.080 61.700 20.120 ;
        RECT 64.240 20.110 64.410 20.120 ;
        RECT 18.330 19.950 18.650 19.980 ;
        RECT 18.330 19.760 18.660 19.950 ;
        RECT 40.880 19.790 41.050 19.840 ;
        RECT 18.330 19.720 18.650 19.760 ;
        RECT 40.850 19.570 41.070 19.790 ;
        RECT 40.880 19.510 41.050 19.570 ;
        RECT 41.400 19.430 41.730 19.610 ;
        RECT 44.540 19.600 44.710 19.650 ;
        RECT 41.980 19.430 44.140 19.600 ;
        RECT 44.380 19.430 44.710 19.600 ;
        RECT 45.000 19.460 45.210 19.790 ;
        RECT 60.580 19.770 60.750 19.810 ;
        RECT 18.810 19.180 19.130 19.210 ;
        RECT 18.810 18.990 19.140 19.180 ;
        RECT 19.520 19.120 19.840 19.150 ;
        RECT 18.810 18.950 19.130 18.990 ;
        RECT 19.520 18.930 19.850 19.120 ;
        RECT 41.430 18.990 41.700 19.430 ;
        RECT 42.910 19.170 43.240 19.430 ;
        RECT 44.450 19.290 44.710 19.430 ;
        RECT 45.450 19.290 45.630 19.730 ;
        RECT 46.180 19.520 47.540 19.630 ;
        RECT 60.520 19.600 60.750 19.770 ;
        RECT 46.180 19.460 47.620 19.520 ;
        RECT 46.980 19.450 47.620 19.460 ;
        RECT 41.470 18.980 41.700 18.990 ;
        RECT 44.450 19.120 45.630 19.290 ;
        RECT 47.150 19.350 47.620 19.450 ;
        RECT 48.090 19.370 49.050 19.540 ;
        RECT 44.450 18.980 44.710 19.120 ;
        RECT 47.150 19.100 47.400 19.350 ;
        RECT 19.520 18.890 19.840 18.930 ;
        RECT 41.470 18.810 42.230 18.980 ;
        RECT 42.480 18.810 43.650 18.980 ;
        RECT 43.890 18.950 44.710 18.980 ;
        RECT 45.950 18.950 46.130 19.010 ;
        RECT 43.890 18.810 45.000 18.950 ;
        RECT 42.880 18.710 43.230 18.810 ;
        RECT 44.540 18.780 45.000 18.810 ;
        RECT 45.450 18.780 46.130 18.950 ;
        RECT 47.070 18.930 47.400 19.100 ;
        RECT 48.870 18.910 49.050 19.370 ;
        RECT 60.580 19.250 60.750 19.600 ;
        RECT 60.920 19.670 61.110 19.690 ;
        RECT 63.920 19.670 64.250 19.850 ;
        RECT 60.920 19.500 61.480 19.670 ;
        RECT 61.940 19.500 64.690 19.670 ;
        RECT 60.920 19.460 61.110 19.500 ;
        RECT 65.220 19.430 65.390 20.360 ;
        RECT 65.620 19.560 65.790 20.410 ;
        RECT 68.490 20.360 68.810 20.390 ;
        RECT 68.490 20.190 70.280 20.360 ;
        RECT 68.490 20.170 68.820 20.190 ;
        RECT 68.490 20.130 68.810 20.170 ;
        RECT 70.110 19.960 70.280 20.190 ;
        RECT 68.960 19.710 69.300 19.960 ;
        RECT 69.470 19.790 69.800 19.960 ;
        RECT 70.020 19.790 70.360 19.960 ;
        RECT 68.640 19.450 69.300 19.710 ;
        RECT 69.550 19.620 69.720 19.790 ;
        RECT 70.110 19.620 70.280 19.790 ;
        RECT 69.470 19.450 69.800 19.620 ;
        RECT 70.020 19.450 70.360 19.620 ;
        RECT 69.550 19.220 69.800 19.450 ;
        RECT 70.680 19.370 71.190 20.040 ;
        RECT 69.550 19.050 70.220 19.220 ;
        RECT 45.490 18.760 46.130 18.780 ;
        RECT 45.950 18.750 46.130 18.760 ;
        RECT 47.730 18.750 48.330 18.900 ;
        RECT 45.950 18.730 48.330 18.750 ;
        RECT 48.790 18.740 49.120 18.910 ;
        RECT 45.950 18.580 48.180 18.730 ;
        RECT 57.050 18.720 57.370 18.760 ;
        RECT 57.050 18.530 57.380 18.720 ;
        RECT 60.580 18.660 60.750 19.010 ;
        RECT 57.050 18.500 57.370 18.530 ;
        RECT 16.210 17.890 16.380 17.960 ;
        RECT 16.140 17.860 16.460 17.890 ;
        RECT 16.130 17.670 16.460 17.860 ;
        RECT 16.140 17.630 16.460 17.670 ;
        RECT 16.210 15.120 16.380 17.630 ;
        RECT 16.760 17.220 16.930 17.960 ;
        RECT 17.310 17.900 17.480 17.960 ;
        RECT 17.240 17.870 17.560 17.900 ;
        RECT 17.230 17.680 17.560 17.870 ;
        RECT 17.240 17.640 17.560 17.680 ;
        RECT 16.690 17.190 17.010 17.220 ;
        RECT 16.680 17.000 17.010 17.190 ;
        RECT 16.690 16.960 17.010 17.000 ;
        RECT 16.760 15.850 16.930 16.960 ;
        RECT 16.690 15.820 17.010 15.850 ;
        RECT 16.680 15.630 17.010 15.820 ;
        RECT 16.690 15.590 17.010 15.630 ;
        RECT 16.140 15.090 16.460 15.120 ;
        RECT 16.130 14.900 16.460 15.090 ;
        RECT 16.140 14.860 16.460 14.900 ;
        RECT 16.210 13.780 16.380 14.860 ;
        RECT 16.130 13.750 16.450 13.780 ;
        RECT 16.120 13.560 16.450 13.750 ;
        RECT 16.130 13.520 16.450 13.560 ;
        RECT 16.210 12.780 16.380 13.520 ;
        RECT 16.760 13.080 16.930 15.590 ;
        RECT 17.310 15.120 17.480 17.640 ;
        RECT 17.860 17.220 18.030 17.960 ;
        RECT 18.410 17.900 18.580 17.960 ;
        RECT 18.330 17.870 18.650 17.900 ;
        RECT 18.320 17.680 18.650 17.870 ;
        RECT 18.330 17.640 18.650 17.680 ;
        RECT 17.790 17.190 18.110 17.220 ;
        RECT 17.780 17.000 18.110 17.190 ;
        RECT 17.790 16.960 18.110 17.000 ;
        RECT 17.860 15.850 18.030 16.960 ;
        RECT 17.790 15.820 18.110 15.850 ;
        RECT 17.780 15.630 18.110 15.820 ;
        RECT 17.790 15.590 18.110 15.630 ;
        RECT 17.240 15.090 17.560 15.120 ;
        RECT 17.230 14.900 17.560 15.090 ;
        RECT 17.240 14.860 17.560 14.900 ;
        RECT 17.310 13.770 17.480 14.860 ;
        RECT 17.240 13.740 17.560 13.770 ;
        RECT 17.230 13.550 17.560 13.740 ;
        RECT 17.240 13.510 17.560 13.550 ;
        RECT 16.690 13.050 17.010 13.080 ;
        RECT 16.680 12.860 17.010 13.050 ;
        RECT 16.690 12.820 17.010 12.860 ;
        RECT 16.760 12.780 16.930 12.820 ;
        RECT 17.310 12.780 17.480 13.510 ;
        RECT 17.860 13.070 18.030 15.590 ;
        RECT 18.410 15.120 18.580 17.640 ;
        RECT 18.960 17.220 19.130 17.960 ;
        RECT 19.370 17.680 19.880 18.360 ;
        RECT 40.880 18.240 41.050 18.290 ;
        RECT 40.850 18.020 41.070 18.240 ;
        RECT 40.880 17.960 41.050 18.020 ;
        RECT 41.400 17.880 41.730 18.060 ;
        RECT 44.540 18.050 44.710 18.100 ;
        RECT 41.980 17.880 44.140 18.050 ;
        RECT 44.380 17.880 44.710 18.050 ;
        RECT 45.000 17.910 45.210 18.240 ;
        RECT 19.370 17.610 19.890 17.680 ;
        RECT 19.380 17.350 19.890 17.610 ;
        RECT 41.430 17.440 41.700 17.880 ;
        RECT 42.910 17.620 43.240 17.880 ;
        RECT 44.450 17.740 44.710 17.880 ;
        RECT 45.450 17.740 45.630 18.180 ;
        RECT 46.180 17.970 47.540 18.080 ;
        RECT 46.180 17.910 47.620 17.970 ;
        RECT 46.980 17.900 47.620 17.910 ;
        RECT 41.470 17.430 41.700 17.440 ;
        RECT 44.450 17.570 45.630 17.740 ;
        RECT 47.150 17.800 47.620 17.900 ;
        RECT 48.090 17.820 49.050 17.990 ;
        RECT 44.450 17.430 44.710 17.570 ;
        RECT 47.150 17.550 47.400 17.800 ;
        RECT 41.470 17.260 42.230 17.430 ;
        RECT 42.480 17.260 43.650 17.430 ;
        RECT 43.890 17.400 44.710 17.430 ;
        RECT 45.950 17.400 46.130 17.460 ;
        RECT 43.890 17.260 45.000 17.400 ;
        RECT 18.890 17.190 19.210 17.220 ;
        RECT 18.880 17.000 19.210 17.190 ;
        RECT 42.880 17.160 43.230 17.260 ;
        RECT 44.540 17.230 45.000 17.260 ;
        RECT 45.450 17.230 46.130 17.400 ;
        RECT 47.070 17.380 47.400 17.550 ;
        RECT 48.870 17.360 49.050 17.820 ;
        RECT 57.100 17.910 57.280 18.500 ;
        RECT 60.520 18.490 60.750 18.660 ;
        RECT 60.920 18.760 61.110 18.800 ;
        RECT 60.920 18.590 61.480 18.760 ;
        RECT 61.940 18.590 64.690 18.760 ;
        RECT 60.920 18.570 61.110 18.590 ;
        RECT 60.580 18.450 60.750 18.490 ;
        RECT 63.920 18.410 64.250 18.590 ;
        RECT 57.100 17.870 57.420 17.910 ;
        RECT 57.100 17.680 57.430 17.870 ;
        RECT 60.650 17.850 60.820 18.270 ;
        RECT 61.460 18.140 61.700 18.180 ;
        RECT 64.240 18.140 64.410 18.150 ;
        RECT 61.130 17.970 61.700 18.140 ;
        RECT 61.940 17.970 63.280 18.140 ;
        RECT 63.730 17.970 64.690 18.140 ;
        RECT 61.460 17.940 61.700 17.970 ;
        RECT 65.220 17.900 65.390 18.830 ;
        RECT 69.550 18.820 69.800 19.050 ;
        RECT 65.620 17.850 65.790 18.700 ;
        RECT 68.640 18.560 69.300 18.820 ;
        RECT 69.470 18.650 69.800 18.820 ;
        RECT 70.020 18.650 70.360 18.820 ;
        RECT 68.960 18.310 69.300 18.560 ;
        RECT 69.550 18.480 69.720 18.650 ;
        RECT 70.110 18.480 70.280 18.650 ;
        RECT 69.470 18.310 69.800 18.480 ;
        RECT 70.020 18.310 70.360 18.480 ;
        RECT 68.490 18.100 68.810 18.140 ;
        RECT 68.490 18.080 68.820 18.100 ;
        RECT 70.110 18.080 70.280 18.310 ;
        RECT 70.680 18.230 71.190 18.900 ;
        RECT 68.490 17.910 70.280 18.080 ;
        RECT 68.490 17.880 68.810 17.910 ;
        RECT 57.100 17.650 57.420 17.680 ;
        RECT 45.490 17.210 46.130 17.230 ;
        RECT 45.950 17.200 46.130 17.210 ;
        RECT 47.730 17.200 48.330 17.350 ;
        RECT 45.950 17.180 48.330 17.200 ;
        RECT 48.790 17.190 49.120 17.360 ;
        RECT 18.890 16.960 19.210 17.000 ;
        RECT 18.960 15.850 19.130 16.960 ;
        RECT 19.670 15.970 19.840 17.160 ;
        RECT 45.950 17.030 48.180 17.180 ;
        RECT 18.890 15.820 19.210 15.850 ;
        RECT 18.880 15.630 19.210 15.820 ;
        RECT 18.890 15.590 19.210 15.630 ;
        RECT 18.330 15.090 18.650 15.120 ;
        RECT 18.320 14.900 18.650 15.090 ;
        RECT 18.330 14.860 18.650 14.900 ;
        RECT 18.410 13.750 18.580 14.860 ;
        RECT 18.330 13.720 18.650 13.750 ;
        RECT 18.320 13.530 18.650 13.720 ;
        RECT 18.330 13.490 18.650 13.530 ;
        RECT 17.790 13.040 18.110 13.070 ;
        RECT 17.780 12.850 18.110 13.040 ;
        RECT 17.790 12.810 18.110 12.850 ;
        RECT 17.860 12.780 18.030 12.810 ;
        RECT 18.410 12.780 18.580 13.490 ;
        RECT 18.960 13.070 19.130 15.590 ;
        RECT 26.000 13.660 26.760 14.080 ;
        RECT 18.880 13.040 19.200 13.070 ;
        RECT 18.870 12.850 19.200 13.040 ;
        RECT 26.020 12.870 26.760 13.660 ;
        RECT 18.880 12.810 19.200 12.850 ;
        RECT 18.960 12.780 19.130 12.810 ;
        RECT 57.540 11.930 57.710 11.960 ;
        RECT 58.090 11.930 58.260 11.960 ;
        RECT 58.640 11.930 58.810 11.960 ;
        RECT 59.190 11.930 59.360 11.960 ;
        RECT 16.180 10.300 16.500 10.330 ;
        RECT 17.280 10.310 17.600 10.340 ;
        RECT 18.370 10.310 18.690 10.340 ;
        RECT 16.170 10.110 16.500 10.300 ;
        RECT 17.270 10.120 17.600 10.310 ;
        RECT 18.360 10.270 18.690 10.310 ;
        RECT 19.410 10.270 19.920 10.800 ;
        RECT 16.180 10.070 16.500 10.110 ;
        RECT 17.280 10.080 17.600 10.120 ;
        RECT 17.710 9.660 17.880 10.270 ;
        RECT 18.260 10.080 18.690 10.270 ;
        RECT 16.730 9.630 17.050 9.660 ;
        RECT 16.720 9.440 17.050 9.630 ;
        RECT 16.730 9.400 17.050 9.440 ;
        RECT 17.710 9.400 18.150 9.660 ;
        RECT 17.710 8.290 17.880 9.400 ;
        RECT 16.730 8.260 17.050 8.290 ;
        RECT 16.720 8.070 17.050 8.260 ;
        RECT 16.730 8.030 17.050 8.070 ;
        RECT 17.710 8.030 18.150 8.290 ;
        RECT 16.250 7.990 16.410 8.000 ;
        RECT 16.800 7.990 16.960 8.000 ;
        RECT 17.350 7.990 17.510 8.000 ;
        RECT 16.240 7.640 16.410 7.990 ;
        RECT 16.790 7.660 16.960 7.990 ;
        RECT 17.340 7.660 17.510 7.990 ;
        RECT 17.710 7.770 17.880 8.030 ;
        RECT 17.900 7.990 18.060 8.000 ;
        RECT 16.250 7.620 16.410 7.640 ;
        RECT 16.800 7.620 16.960 7.660 ;
        RECT 17.350 7.620 17.510 7.660 ;
        RECT 17.890 7.590 18.060 7.990 ;
        RECT 18.260 7.770 18.430 10.080 ;
        RECT 18.810 9.660 18.980 10.270 ;
        RECT 19.360 9.790 20.080 10.270 ;
        RECT 18.810 9.400 19.250 9.660 ;
        RECT 18.810 8.290 18.980 9.400 ;
        RECT 18.810 8.030 19.250 8.290 ;
        RECT 18.450 7.990 18.610 8.000 ;
        RECT 18.440 7.660 18.610 7.990 ;
        RECT 18.810 7.770 18.980 8.030 ;
        RECT 19.000 7.990 19.160 8.000 ;
        RECT 18.450 7.620 18.610 7.660 ;
        RECT 18.990 7.650 19.160 7.990 ;
        RECT 19.360 7.770 19.530 9.790 ;
        RECT 19.910 7.770 20.080 9.790 ;
        RECT 20.460 7.770 20.630 10.260 ;
        RECT 47.730 9.440 47.900 11.930 ;
        RECT 48.280 9.430 48.450 11.930 ;
        RECT 48.830 9.430 49.000 11.930 ;
        RECT 49.380 11.620 49.550 11.930 ;
        RECT 49.120 11.360 49.550 11.620 ;
        RECT 49.380 9.430 49.550 11.360 ;
        RECT 49.930 10.940 50.100 11.930 ;
        RECT 50.480 11.620 50.650 11.930 ;
        RECT 50.210 11.360 50.650 11.620 ;
        RECT 49.670 10.680 50.100 10.940 ;
        RECT 49.930 9.570 50.100 10.680 ;
        RECT 49.670 9.430 50.100 9.570 ;
        RECT 50.480 9.430 50.650 11.360 ;
        RECT 51.310 11.570 51.630 11.610 ;
        RECT 51.310 11.380 51.640 11.570 ;
        RECT 51.310 11.350 51.630 11.380 ;
        RECT 52.490 10.980 52.660 11.740 ;
        RECT 54.380 10.980 54.550 11.740 ;
        RECT 56.390 11.620 56.560 11.930 ;
        RECT 55.410 11.570 55.730 11.610 ;
        RECT 55.400 11.380 55.730 11.570 ;
        RECT 55.410 11.350 55.730 11.380 ;
        RECT 56.390 11.360 56.830 11.620 ;
        RECT 50.760 10.880 51.080 10.920 ;
        RECT 50.760 10.690 51.090 10.880 ;
        RECT 51.870 10.870 52.190 10.910 ;
        RECT 54.850 10.870 55.170 10.910 ;
        RECT 55.960 10.880 56.280 10.920 ;
        RECT 50.760 10.660 51.080 10.690 ;
        RECT 51.870 10.680 52.200 10.870 ;
        RECT 54.840 10.680 55.170 10.870 ;
        RECT 55.950 10.690 56.280 10.880 ;
        RECT 51.870 10.650 52.190 10.680 ;
        RECT 54.850 10.650 55.170 10.680 ;
        RECT 55.960 10.660 56.280 10.690 ;
        RECT 50.760 9.530 51.080 9.570 ;
        RECT 51.860 9.530 52.180 9.570 ;
        RECT 54.860 9.530 55.180 9.570 ;
        RECT 55.960 9.530 56.280 9.570 ;
        RECT 49.670 9.340 50.000 9.430 ;
        RECT 50.760 9.340 51.090 9.530 ;
        RECT 51.860 9.340 52.190 9.530 ;
        RECT 54.850 9.340 55.180 9.530 ;
        RECT 55.950 9.340 56.280 9.530 ;
        RECT 56.390 9.430 56.560 11.360 ;
        RECT 56.940 10.940 57.110 11.930 ;
        RECT 57.490 11.620 57.710 11.930 ;
        RECT 57.490 11.360 57.920 11.620 ;
        RECT 56.940 10.680 57.370 10.940 ;
        RECT 56.940 9.570 57.110 10.680 ;
        RECT 56.940 9.430 57.370 9.570 ;
        RECT 57.490 9.470 57.710 11.360 ;
        RECT 57.490 9.430 57.660 9.470 ;
        RECT 58.040 9.460 58.260 11.930 ;
        RECT 58.590 9.460 58.810 11.930 ;
        RECT 59.140 11.650 59.360 11.930 ;
        RECT 58.930 11.390 59.360 11.650 ;
        RECT 59.140 9.460 59.360 11.390 ;
        RECT 59.740 10.970 59.910 11.960 ;
        RECT 60.290 11.650 60.460 11.960 ;
        RECT 60.020 11.390 60.460 11.650 ;
        RECT 59.480 10.710 59.910 10.970 ;
        RECT 59.740 9.600 59.910 10.710 ;
        RECT 59.480 9.460 59.910 9.600 ;
        RECT 60.290 9.460 60.460 11.390 ;
        RECT 61.120 11.600 61.440 11.640 ;
        RECT 61.120 11.410 61.450 11.600 ;
        RECT 61.120 11.380 61.440 11.410 ;
        RECT 62.300 11.010 62.470 11.770 ;
        RECT 64.190 11.010 64.360 11.770 ;
        RECT 66.200 11.650 66.370 11.960 ;
        RECT 65.220 11.600 65.540 11.640 ;
        RECT 65.210 11.410 65.540 11.600 ;
        RECT 65.220 11.380 65.540 11.410 ;
        RECT 66.200 11.390 66.640 11.650 ;
        RECT 60.570 10.910 60.890 10.950 ;
        RECT 60.570 10.720 60.900 10.910 ;
        RECT 61.680 10.900 62.000 10.940 ;
        RECT 64.660 10.900 64.980 10.940 ;
        RECT 65.770 10.910 66.090 10.950 ;
        RECT 60.570 10.690 60.890 10.720 ;
        RECT 61.680 10.710 62.010 10.900 ;
        RECT 64.650 10.710 64.980 10.900 ;
        RECT 65.760 10.720 66.090 10.910 ;
        RECT 61.680 10.680 62.000 10.710 ;
        RECT 64.660 10.680 64.980 10.710 ;
        RECT 65.770 10.690 66.090 10.720 ;
        RECT 60.570 9.560 60.890 9.600 ;
        RECT 61.670 9.560 61.990 9.600 ;
        RECT 64.670 9.560 64.990 9.600 ;
        RECT 65.770 9.560 66.090 9.600 ;
        RECT 58.040 9.430 58.210 9.460 ;
        RECT 58.590 9.430 58.760 9.460 ;
        RECT 59.140 9.440 59.310 9.460 ;
        RECT 57.040 9.340 57.370 9.430 ;
        RECT 59.480 9.370 59.810 9.460 ;
        RECT 60.570 9.370 60.900 9.560 ;
        RECT 61.670 9.370 62.000 9.560 ;
        RECT 64.660 9.370 64.990 9.560 ;
        RECT 65.760 9.370 66.090 9.560 ;
        RECT 66.200 9.460 66.370 11.390 ;
        RECT 66.750 10.970 66.920 11.960 ;
        RECT 67.300 11.650 67.470 11.960 ;
        RECT 67.300 11.390 67.730 11.650 ;
        RECT 66.750 10.710 67.180 10.970 ;
        RECT 66.750 9.600 66.920 10.710 ;
        RECT 66.750 9.460 67.180 9.600 ;
        RECT 67.300 9.460 67.470 11.390 ;
        RECT 67.850 9.460 68.020 11.960 ;
        RECT 68.400 9.460 68.570 11.960 ;
        RECT 68.950 9.470 69.120 11.960 ;
        RECT 70.480 10.920 70.650 11.660 ;
        RECT 71.030 11.620 71.200 11.660 ;
        RECT 70.960 11.580 71.280 11.620 ;
        RECT 70.950 11.390 71.280 11.580 ;
        RECT 70.960 11.360 71.280 11.390 ;
        RECT 70.400 10.880 70.720 10.920 ;
        RECT 70.390 10.690 70.720 10.880 ;
        RECT 70.400 10.660 70.720 10.690 ;
        RECT 70.480 9.580 70.650 10.660 ;
        RECT 70.410 9.540 70.730 9.580 ;
        RECT 66.850 9.370 67.180 9.460 ;
        RECT 59.480 9.340 59.800 9.370 ;
        RECT 60.570 9.340 60.890 9.370 ;
        RECT 61.670 9.340 61.990 9.370 ;
        RECT 64.670 9.340 64.990 9.370 ;
        RECT 65.770 9.340 66.090 9.370 ;
        RECT 66.860 9.340 67.180 9.370 ;
        RECT 70.400 9.350 70.730 9.540 ;
        RECT 49.670 9.310 49.990 9.340 ;
        RECT 50.760 9.310 51.080 9.340 ;
        RECT 51.860 9.310 52.180 9.340 ;
        RECT 54.860 9.310 55.180 9.340 ;
        RECT 55.960 9.310 56.280 9.340 ;
        RECT 57.050 9.310 57.370 9.340 ;
        RECT 70.410 9.320 70.730 9.350 ;
        RECT 49.200 9.220 49.360 9.250 ;
        RECT 19.000 7.620 19.160 7.650 ;
        RECT 16.180 7.530 16.500 7.560 ;
        RECT 17.280 7.530 17.600 7.560 ;
        RECT 18.370 7.530 18.690 7.560 ;
        RECT 16.170 7.340 16.500 7.530 ;
        RECT 17.270 7.340 17.600 7.530 ;
        RECT 18.360 7.440 18.690 7.530 ;
        RECT 16.180 7.300 16.500 7.340 ;
        RECT 17.280 7.300 17.600 7.340 ;
        RECT 16.170 6.190 16.490 6.220 ;
        RECT 16.160 6.000 16.490 6.190 ;
        RECT 17.280 6.180 17.600 6.210 ;
        RECT 16.170 5.960 16.490 6.000 ;
        RECT 17.270 5.990 17.600 6.180 ;
        RECT 17.280 5.950 17.600 5.990 ;
        RECT 15.700 5.130 15.870 5.890 ;
        RECT 16.730 5.490 17.050 5.520 ;
        RECT 16.720 5.300 17.050 5.490 ;
        RECT 16.730 5.260 17.050 5.300 ;
        RECT 17.710 5.510 17.880 7.440 ;
        RECT 18.260 7.300 18.690 7.440 ;
        RECT 18.260 6.190 18.430 7.300 ;
        RECT 18.260 5.930 18.690 6.190 ;
        RECT 17.710 5.250 18.150 5.510 ;
        RECT 17.710 4.940 17.880 5.250 ;
        RECT 18.260 4.940 18.430 5.930 ;
        RECT 18.810 5.510 18.980 7.440 ;
        RECT 18.810 5.250 19.240 5.510 ;
        RECT 18.810 4.940 18.980 5.250 ;
        RECT 19.360 4.940 19.530 7.440 ;
        RECT 19.910 4.940 20.080 7.440 ;
        RECT 20.460 5.340 20.630 7.430 ;
        RECT 47.730 6.610 47.900 9.100 ;
        RECT 48.280 7.080 48.450 9.100 ;
        RECT 48.830 7.080 49.000 9.100 ;
        RECT 49.200 8.880 49.370 9.220 ;
        RECT 49.750 9.210 49.910 9.250 ;
        RECT 49.200 8.870 49.360 8.880 ;
        RECT 49.380 8.840 49.550 9.100 ;
        RECT 49.750 8.880 49.920 9.210 ;
        RECT 49.750 8.870 49.910 8.880 ;
        RECT 49.110 8.580 49.550 8.840 ;
        RECT 49.380 7.470 49.550 8.580 ;
        RECT 49.110 7.210 49.550 7.470 ;
        RECT 48.280 6.600 49.000 7.080 ;
        RECT 49.380 6.600 49.550 7.210 ;
        RECT 49.930 6.790 50.100 9.100 ;
        RECT 50.300 8.880 50.470 9.280 ;
        RECT 50.850 9.210 51.010 9.250 ;
        RECT 51.400 9.210 51.560 9.250 ;
        RECT 51.950 9.230 52.110 9.250 ;
        RECT 54.930 9.230 55.090 9.250 ;
        RECT 50.300 8.870 50.460 8.880 ;
        RECT 50.480 8.840 50.650 9.100 ;
        RECT 50.850 8.880 51.020 9.210 ;
        RECT 51.400 8.880 51.570 9.210 ;
        RECT 51.950 8.880 52.120 9.230 ;
        RECT 54.920 8.880 55.090 9.230 ;
        RECT 55.480 9.210 55.640 9.250 ;
        RECT 56.030 9.210 56.190 9.250 ;
        RECT 55.470 8.880 55.640 9.210 ;
        RECT 56.020 8.880 56.190 9.210 ;
        RECT 50.850 8.870 51.010 8.880 ;
        RECT 51.400 8.870 51.560 8.880 ;
        RECT 51.950 8.870 52.110 8.880 ;
        RECT 54.930 8.870 55.090 8.880 ;
        RECT 55.480 8.870 55.640 8.880 ;
        RECT 56.030 8.870 56.190 8.880 ;
        RECT 56.390 8.840 56.560 9.100 ;
        RECT 56.570 8.880 56.740 9.280 ;
        RECT 59.010 9.250 59.170 9.280 ;
        RECT 57.130 9.210 57.290 9.250 ;
        RECT 57.680 9.220 57.840 9.250 ;
        RECT 56.580 8.870 56.740 8.880 ;
        RECT 50.210 8.580 50.650 8.840 ;
        RECT 51.310 8.800 51.630 8.840 ;
        RECT 55.410 8.800 55.730 8.840 ;
        RECT 51.310 8.610 51.640 8.800 ;
        RECT 55.400 8.610 55.730 8.800 ;
        RECT 51.310 8.580 51.630 8.610 ;
        RECT 55.410 8.580 55.730 8.610 ;
        RECT 56.390 8.580 56.830 8.840 ;
        RECT 50.480 7.470 50.650 8.580 ;
        RECT 56.390 7.470 56.560 8.580 ;
        RECT 50.210 7.210 50.650 7.470 ;
        RECT 51.310 7.430 51.630 7.470 ;
        RECT 55.410 7.430 55.730 7.470 ;
        RECT 51.310 7.240 51.640 7.430 ;
        RECT 55.400 7.240 55.730 7.430 ;
        RECT 51.310 7.210 51.630 7.240 ;
        RECT 55.410 7.210 55.730 7.240 ;
        RECT 56.390 7.210 56.830 7.470 ;
        RECT 49.670 6.600 50.100 6.790 ;
        RECT 50.480 6.600 50.650 7.210 ;
        RECT 50.760 6.750 51.080 6.790 ;
        RECT 51.860 6.760 52.180 6.800 ;
        RECT 54.860 6.760 55.180 6.800 ;
        RECT 48.440 6.070 48.950 6.600 ;
        RECT 49.670 6.560 50.000 6.600 ;
        RECT 50.760 6.560 51.090 6.750 ;
        RECT 51.860 6.570 52.190 6.760 ;
        RECT 54.850 6.570 55.180 6.760 ;
        RECT 55.960 6.750 56.280 6.790 ;
        RECT 49.670 6.530 49.990 6.560 ;
        RECT 50.760 6.530 51.080 6.560 ;
        RECT 51.860 6.540 52.180 6.570 ;
        RECT 54.860 6.540 55.180 6.570 ;
        RECT 55.950 6.560 56.280 6.750 ;
        RECT 56.390 6.600 56.560 7.210 ;
        RECT 56.940 6.790 57.110 9.100 ;
        RECT 57.120 8.880 57.290 9.210 ;
        RECT 57.670 9.130 57.840 9.220 ;
        RECT 57.540 9.100 57.840 9.130 ;
        RECT 58.090 9.100 58.260 9.130 ;
        RECT 58.640 9.100 58.810 9.130 ;
        RECT 57.130 8.870 57.290 8.880 ;
        RECT 57.490 8.870 57.840 9.100 ;
        RECT 57.490 8.840 57.710 8.870 ;
        RECT 57.490 8.580 57.930 8.840 ;
        RECT 57.490 7.470 57.710 8.580 ;
        RECT 57.490 7.210 57.930 7.470 ;
        RECT 56.940 6.600 57.370 6.790 ;
        RECT 57.490 6.640 57.710 7.210 ;
        RECT 58.040 7.110 58.260 9.100 ;
        RECT 58.590 7.110 58.810 9.100 ;
        RECT 59.010 9.100 59.180 9.250 ;
        RECT 59.560 9.240 59.720 9.280 ;
        RECT 59.190 9.100 59.360 9.130 ;
        RECT 59.010 8.900 59.360 9.100 ;
        RECT 59.560 8.910 59.730 9.240 ;
        RECT 59.560 8.900 59.720 8.910 ;
        RECT 59.140 8.870 59.360 8.900 ;
        RECT 58.920 8.610 59.360 8.870 ;
        RECT 59.140 7.500 59.360 8.610 ;
        RECT 58.920 7.240 59.360 7.500 ;
        RECT 57.490 6.600 57.660 6.640 ;
        RECT 58.040 6.630 58.810 7.110 ;
        RECT 59.140 6.630 59.360 7.240 ;
        RECT 59.740 6.820 59.910 9.130 ;
        RECT 60.110 8.910 60.280 9.310 ;
        RECT 60.660 9.240 60.820 9.280 ;
        RECT 61.210 9.240 61.370 9.280 ;
        RECT 61.760 9.260 61.920 9.280 ;
        RECT 64.740 9.260 64.900 9.280 ;
        RECT 60.110 8.900 60.270 8.910 ;
        RECT 60.290 8.870 60.460 9.130 ;
        RECT 60.660 8.910 60.830 9.240 ;
        RECT 61.210 8.910 61.380 9.240 ;
        RECT 61.760 8.910 61.930 9.260 ;
        RECT 64.730 8.910 64.900 9.260 ;
        RECT 65.290 9.240 65.450 9.280 ;
        RECT 65.840 9.240 66.000 9.280 ;
        RECT 65.280 8.910 65.450 9.240 ;
        RECT 65.830 8.910 66.000 9.240 ;
        RECT 60.660 8.900 60.820 8.910 ;
        RECT 61.210 8.900 61.370 8.910 ;
        RECT 61.760 8.900 61.920 8.910 ;
        RECT 64.740 8.900 64.900 8.910 ;
        RECT 65.290 8.900 65.450 8.910 ;
        RECT 65.840 8.900 66.000 8.910 ;
        RECT 66.200 8.870 66.370 9.130 ;
        RECT 66.380 8.910 66.550 9.310 ;
        RECT 66.940 9.240 67.100 9.280 ;
        RECT 67.490 9.250 67.650 9.280 ;
        RECT 66.390 8.900 66.550 8.910 ;
        RECT 60.020 8.610 60.460 8.870 ;
        RECT 61.120 8.830 61.440 8.870 ;
        RECT 65.220 8.830 65.540 8.870 ;
        RECT 61.120 8.640 61.450 8.830 ;
        RECT 65.210 8.640 65.540 8.830 ;
        RECT 61.120 8.610 61.440 8.640 ;
        RECT 65.220 8.610 65.540 8.640 ;
        RECT 66.200 8.610 66.640 8.870 ;
        RECT 60.290 7.500 60.460 8.610 ;
        RECT 66.200 7.500 66.370 8.610 ;
        RECT 60.020 7.240 60.460 7.500 ;
        RECT 61.120 7.460 61.440 7.500 ;
        RECT 65.220 7.460 65.540 7.500 ;
        RECT 61.120 7.270 61.450 7.460 ;
        RECT 65.210 7.270 65.540 7.460 ;
        RECT 61.120 7.240 61.440 7.270 ;
        RECT 65.220 7.240 65.540 7.270 ;
        RECT 66.200 7.240 66.640 7.500 ;
        RECT 59.480 6.630 59.910 6.820 ;
        RECT 60.290 6.630 60.460 7.240 ;
        RECT 60.570 6.780 60.890 6.820 ;
        RECT 61.670 6.790 61.990 6.830 ;
        RECT 64.670 6.790 64.990 6.830 ;
        RECT 58.040 6.600 58.760 6.630 ;
        RECT 59.140 6.610 59.310 6.630 ;
        RECT 57.040 6.560 57.370 6.600 ;
        RECT 55.960 6.530 56.280 6.560 ;
        RECT 57.050 6.530 57.370 6.560 ;
        RECT 58.090 6.100 58.760 6.600 ;
        RECT 59.480 6.590 59.810 6.630 ;
        RECT 60.570 6.590 60.900 6.780 ;
        RECT 61.670 6.600 62.000 6.790 ;
        RECT 64.660 6.600 64.990 6.790 ;
        RECT 65.770 6.780 66.090 6.820 ;
        RECT 59.480 6.560 59.800 6.590 ;
        RECT 60.570 6.560 60.890 6.590 ;
        RECT 61.670 6.570 61.990 6.600 ;
        RECT 64.670 6.570 64.990 6.600 ;
        RECT 65.760 6.590 66.090 6.780 ;
        RECT 66.200 6.630 66.370 7.240 ;
        RECT 66.750 6.820 66.920 9.130 ;
        RECT 66.930 8.910 67.100 9.240 ;
        RECT 66.940 8.900 67.100 8.910 ;
        RECT 67.300 8.870 67.470 9.130 ;
        RECT 67.480 8.910 67.650 9.250 ;
        RECT 67.490 8.900 67.650 8.910 ;
        RECT 67.300 8.610 67.740 8.870 ;
        RECT 67.300 7.500 67.470 8.610 ;
        RECT 67.300 7.240 67.740 7.500 ;
        RECT 66.750 6.630 67.180 6.820 ;
        RECT 67.300 6.630 67.470 7.240 ;
        RECT 67.850 7.110 68.020 9.130 ;
        RECT 68.400 7.110 68.570 9.130 ;
        RECT 67.850 6.630 68.570 7.110 ;
        RECT 68.950 6.640 69.120 9.130 ;
        RECT 70.480 6.810 70.650 9.320 ;
        RECT 71.030 8.850 71.200 11.360 ;
        RECT 71.580 10.930 71.750 11.660 ;
        RECT 72.130 11.630 72.300 11.660 ;
        RECT 72.060 11.590 72.380 11.630 ;
        RECT 72.050 11.400 72.380 11.590 ;
        RECT 72.060 11.370 72.380 11.400 ;
        RECT 71.510 10.890 71.830 10.930 ;
        RECT 71.500 10.700 71.830 10.890 ;
        RECT 71.510 10.670 71.830 10.700 ;
        RECT 71.580 9.580 71.750 10.670 ;
        RECT 71.510 9.540 71.830 9.580 ;
        RECT 71.500 9.350 71.830 9.540 ;
        RECT 71.510 9.320 71.830 9.350 ;
        RECT 70.960 8.810 71.280 8.850 ;
        RECT 70.950 8.620 71.280 8.810 ;
        RECT 70.960 8.590 71.280 8.620 ;
        RECT 71.030 7.480 71.200 8.590 ;
        RECT 70.960 7.440 71.280 7.480 ;
        RECT 70.950 7.250 71.280 7.440 ;
        RECT 70.960 7.220 71.280 7.250 ;
        RECT 70.410 6.770 70.730 6.810 ;
        RECT 66.850 6.590 67.180 6.630 ;
        RECT 65.770 6.560 66.090 6.590 ;
        RECT 66.860 6.560 67.180 6.590 ;
        RECT 67.900 6.100 68.410 6.630 ;
        RECT 70.400 6.580 70.730 6.770 ;
        RECT 70.410 6.550 70.730 6.580 ;
        RECT 70.480 6.480 70.650 6.550 ;
        RECT 71.030 6.480 71.200 7.220 ;
        RECT 71.580 6.800 71.750 9.320 ;
        RECT 72.130 8.850 72.300 11.370 ;
        RECT 72.680 10.950 72.850 11.660 ;
        RECT 73.230 11.630 73.400 11.660 ;
        RECT 73.150 11.590 73.470 11.630 ;
        RECT 73.140 11.400 73.470 11.590 ;
        RECT 73.150 11.370 73.470 11.400 ;
        RECT 72.600 10.910 72.920 10.950 ;
        RECT 72.590 10.720 72.920 10.910 ;
        RECT 72.600 10.690 72.920 10.720 ;
        RECT 72.680 9.580 72.850 10.690 ;
        RECT 72.600 9.540 72.920 9.580 ;
        RECT 72.590 9.350 72.920 9.540 ;
        RECT 72.600 9.320 72.920 9.350 ;
        RECT 72.060 8.810 72.380 8.850 ;
        RECT 72.050 8.620 72.380 8.810 ;
        RECT 72.060 8.590 72.380 8.620 ;
        RECT 72.130 7.480 72.300 8.590 ;
        RECT 72.060 7.440 72.380 7.480 ;
        RECT 72.050 7.250 72.380 7.440 ;
        RECT 72.060 7.220 72.380 7.250 ;
        RECT 71.510 6.760 71.830 6.800 ;
        RECT 71.500 6.570 71.830 6.760 ;
        RECT 71.510 6.540 71.830 6.570 ;
        RECT 71.580 6.480 71.750 6.540 ;
        RECT 72.130 6.480 72.300 7.220 ;
        RECT 72.680 6.800 72.850 9.320 ;
        RECT 73.230 8.850 73.400 11.370 ;
        RECT 73.160 8.810 73.480 8.850 ;
        RECT 73.150 8.620 73.480 8.810 ;
        RECT 73.160 8.590 73.480 8.620 ;
        RECT 73.230 7.480 73.400 8.590 ;
        RECT 73.160 7.440 73.480 7.480 ;
        RECT 73.150 7.250 73.480 7.440 ;
        RECT 73.940 7.280 74.110 8.470 ;
        RECT 73.160 7.220 73.480 7.250 ;
        RECT 72.600 6.760 72.920 6.800 ;
        RECT 72.590 6.570 72.920 6.760 ;
        RECT 72.600 6.540 72.920 6.570 ;
        RECT 72.680 6.480 72.850 6.540 ;
        RECT 73.230 6.480 73.400 7.220 ;
        RECT 73.650 6.830 74.160 7.090 ;
        RECT 73.640 6.760 74.160 6.830 ;
        RECT 58.090 6.070 58.600 6.100 ;
        RECT 73.640 6.080 74.150 6.760 ;
        RECT 20.350 4.970 22.740 5.340 ;
        RECT 20.400 1.710 22.740 4.970 ;
        RECT 99.150 4.170 99.380 4.180 ;
        RECT 99.130 4.000 103.790 4.170 ;
        RECT 99.150 3.990 99.380 4.000 ;
        RECT 104.690 3.520 104.880 3.530 ;
        RECT 100.350 3.480 104.150 3.490 ;
        RECT 104.660 3.480 104.920 3.520 ;
        RECT 100.350 3.320 104.920 3.480 ;
        RECT 103.920 3.310 104.920 3.320 ;
        RECT 103.920 2.850 104.150 3.310 ;
        RECT 104.660 3.200 104.920 3.310 ;
        RECT 104.690 2.850 104.880 2.860 ;
        RECT 103.920 2.640 104.930 2.850 ;
        RECT 99.150 2.560 99.380 2.570 ;
        RECT 99.130 2.390 103.610 2.560 ;
        RECT 99.150 2.380 99.380 2.390 ;
        RECT 103.920 1.880 104.150 2.640 ;
        RECT 104.660 2.530 104.920 2.640 ;
        RECT 100.370 1.710 104.150 1.880 ;
        RECT 20.400 1.700 22.730 1.710 ;
        RECT 99.150 0.960 99.380 0.970 ;
        RECT 99.130 0.790 103.630 0.960 ;
        RECT 99.150 0.780 99.380 0.790 ;
        RECT 100.370 0.780 100.700 0.790 ;
        RECT 101.330 0.780 101.660 0.790 ;
        RECT 102.290 0.780 102.620 0.790 ;
        RECT 103.250 0.780 103.580 0.790 ;
        RECT 103.920 0.270 104.150 1.710 ;
        RECT 104.600 1.520 105.030 1.540 ;
        RECT 104.580 1.350 105.030 1.520 ;
        RECT 104.600 1.330 105.030 1.350 ;
        RECT 100.370 0.100 104.150 0.270 ;
        RECT 100.430 -0.130 100.860 -0.110 ;
        RECT 100.410 -0.300 100.860 -0.130 ;
        RECT 100.430 -0.320 100.860 -0.300 ;
        RECT 99.150 -0.660 99.380 -0.650 ;
        RECT 99.130 -0.830 103.630 -0.660 ;
        RECT 99.150 -0.840 99.380 -0.830 ;
        RECT 103.920 -1.330 104.150 0.100 ;
        RECT 104.600 -0.090 105.030 -0.070 ;
        RECT 104.580 -0.260 105.030 -0.090 ;
        RECT 104.600 -0.280 105.030 -0.260 ;
        RECT 100.380 -1.340 104.150 -1.330 ;
        RECT 100.370 -1.500 104.150 -1.340 ;
        RECT 100.370 -1.510 100.700 -1.500 ;
        RECT 102.290 -1.510 102.620 -1.500 ;
        RECT 103.250 -1.510 103.580 -1.500 ;
        RECT 101.430 -1.870 101.860 -1.850 ;
        RECT 101.430 -2.040 101.880 -1.870 ;
        RECT 101.430 -2.060 101.860 -2.040 ;
        RECT 99.150 -2.260 99.380 -2.250 ;
        RECT 99.130 -2.430 103.580 -2.260 ;
        RECT 99.150 -2.440 99.380 -2.430 ;
        RECT 100.370 -2.440 100.700 -2.430 ;
        RECT 101.330 -2.440 101.660 -2.430 ;
        RECT 102.290 -2.440 102.620 -2.430 ;
        RECT 103.250 -2.440 103.580 -2.430 ;
        RECT 103.920 -2.950 104.150 -1.500 ;
        RECT 104.590 -1.700 105.020 -1.680 ;
        RECT 104.570 -1.870 105.020 -1.700 ;
        RECT 104.590 -1.890 105.020 -1.870 ;
        RECT 100.360 -3.120 104.150 -2.950 ;
        RECT 102.340 -3.380 102.770 -3.360 ;
        RECT 102.320 -3.550 102.770 -3.380 ;
        RECT 102.340 -3.570 102.770 -3.550 ;
        RECT 99.150 -3.880 99.380 -3.870 ;
        RECT 99.130 -4.050 103.630 -3.880 ;
        RECT 99.150 -4.060 99.380 -4.050 ;
        RECT 100.370 -4.570 100.700 -4.560 ;
        RECT 101.330 -4.570 101.660 -4.560 ;
        RECT 102.290 -4.570 102.620 -4.560 ;
        RECT 103.250 -4.570 103.580 -4.560 ;
        RECT 103.920 -4.570 104.150 -3.120 ;
        RECT 104.590 -3.320 105.020 -3.300 ;
        RECT 104.570 -3.490 105.020 -3.320 ;
        RECT 104.590 -3.510 105.020 -3.490 ;
        RECT 100.360 -4.740 104.150 -4.570 ;
        RECT 99.150 -5.480 99.380 -5.470 ;
        RECT 99.130 -5.490 103.550 -5.480 ;
        RECT 99.130 -5.650 103.580 -5.490 ;
        RECT 99.150 -5.660 99.380 -5.650 ;
        RECT 100.370 -5.660 100.700 -5.650 ;
        RECT 101.330 -5.660 101.660 -5.650 ;
        RECT 102.290 -5.660 102.620 -5.650 ;
        RECT 103.250 -5.660 103.580 -5.650 ;
        RECT 103.920 -6.160 104.150 -4.740 ;
        RECT 104.590 -4.930 105.020 -4.910 ;
        RECT 104.570 -5.100 105.020 -4.930 ;
        RECT 104.590 -5.120 105.020 -5.100 ;
        RECT 110.580 -5.290 110.950 9.580 ;
        RECT 110.580 -5.540 110.960 -5.290 ;
        RECT 100.360 -6.330 104.160 -6.160 ;
        RECT 100.370 -6.340 100.700 -6.330 ;
        RECT 101.330 -6.340 101.660 -6.330 ;
        RECT 102.290 -6.340 102.620 -6.330 ;
        RECT 103.250 -6.340 103.580 -6.330 ;
        RECT 99.150 -7.110 99.380 -7.090 ;
        RECT 100.370 -7.110 100.700 -7.100 ;
        RECT 101.330 -7.110 101.660 -7.100 ;
        RECT 102.290 -7.110 102.620 -7.100 ;
        RECT 103.250 -7.110 103.580 -7.100 ;
        RECT 99.130 -7.280 103.590 -7.110 ;
        RECT 103.920 -7.770 104.150 -6.330 ;
        RECT 104.430 -6.920 104.640 -6.490 ;
        RECT 104.450 -6.940 104.620 -6.920 ;
        RECT 100.360 -7.940 104.150 -7.770 ;
        RECT 100.370 -7.950 100.700 -7.940 ;
        RECT 101.330 -7.950 101.660 -7.940 ;
        RECT 102.290 -7.950 102.620 -7.940 ;
        RECT 103.250 -7.950 103.580 -7.940 ;
        RECT 104.600 -8.130 105.030 -8.110 ;
        RECT 104.580 -8.300 105.030 -8.130 ;
        RECT 104.600 -8.320 105.030 -8.300 ;
        RECT 104.590 -9.720 105.020 -9.700 ;
        RECT 101.390 -9.800 101.820 -9.780 ;
        RECT 102.330 -9.800 102.760 -9.780 ;
        RECT 101.370 -9.970 101.820 -9.800 ;
        RECT 102.310 -9.970 102.760 -9.800 ;
        RECT 103.280 -9.860 103.710 -9.840 ;
        RECT 101.390 -9.990 101.820 -9.970 ;
        RECT 102.330 -9.990 102.760 -9.970 ;
        RECT 103.260 -10.030 103.710 -9.860 ;
        RECT 104.570 -9.890 105.020 -9.720 ;
        RECT 104.590 -9.910 105.020 -9.890 ;
        RECT 103.280 -10.050 103.710 -10.030 ;
      LAYER mcon ;
        RECT 6.670 61.070 6.840 61.240 ;
        RECT 9.540 61.280 9.710 61.450 ;
        RECT 8.080 61.070 8.250 61.240 ;
        RECT 24.880 61.100 25.050 61.270 ;
        RECT 24.880 60.750 25.050 60.920 ;
        RECT 9.540 60.490 9.710 60.660 ;
        RECT 24.880 60.410 25.050 60.580 ;
        RECT 30.740 61.010 30.910 61.180 ;
        RECT 30.740 60.560 30.910 60.730 ;
        RECT 35.440 60.960 35.610 61.130 ;
        RECT 35.440 60.510 35.610 60.680 ;
        RECT 6.670 60.220 6.840 60.390 ;
        RECT 7.390 60.210 7.560 60.380 ;
        RECT 8.080 60.220 8.250 60.390 ;
        RECT 6.850 59.810 7.020 59.980 ;
        RECT 7.910 59.810 8.080 59.980 ;
        RECT 6.670 59.400 6.840 59.570 ;
        RECT 7.390 59.370 7.560 59.540 ;
        RECT 8.080 59.400 8.250 59.570 ;
        RECT 22.780 59.470 22.950 59.640 ;
        RECT 24.140 59.550 24.310 59.720 ;
        RECT 24.830 59.540 25.000 59.710 ;
        RECT 9.540 59.060 9.710 59.230 ;
        RECT 6.670 58.560 6.840 58.730 ;
        RECT 8.080 58.560 8.250 58.730 ;
        RECT 8.810 58.300 8.980 58.470 ;
        RECT 8.800 57.780 8.970 57.950 ;
        RECT 9.550 57.660 9.720 57.830 ;
        RECT 6.670 57.440 6.840 57.610 ;
        RECT 8.080 57.440 8.250 57.610 ;
        RECT 7.370 56.570 7.540 56.740 ;
        RECT 8.800 56.590 8.970 56.760 ;
        RECT 11.560 56.240 11.730 56.410 ;
        RECT 6.580 55.990 6.750 56.160 ;
        RECT 7.510 55.990 7.680 56.160 ;
        RECT 8.210 55.990 8.380 56.160 ;
        RECT 8.950 55.990 9.120 56.160 ;
        RECT 9.660 55.980 9.830 56.150 ;
        RECT 24.880 58.300 25.050 58.470 ;
        RECT 24.880 57.950 25.050 58.120 ;
        RECT 24.880 57.610 25.050 57.780 ;
        RECT 30.740 58.020 30.910 58.190 ;
        RECT 30.740 57.570 30.910 57.740 ;
        RECT 30.740 57.010 30.910 57.180 ;
        RECT 24.880 56.750 25.050 56.920 ;
        RECT 24.880 56.400 25.050 56.570 ;
        RECT 30.740 56.560 30.910 56.730 ;
        RECT 24.880 56.060 25.050 56.230 ;
        RECT 34.660 57.500 34.830 57.670 ;
        RECT 22.060 55.810 22.230 55.980 ;
        RECT 31.920 55.830 32.090 56.000 ;
        RECT 22.070 51.450 22.500 52.190 ;
        RECT 42.960 49.890 43.170 50.100 ;
        RECT 47.840 50.000 48.010 50.170 ;
        RECT 41.490 49.520 41.660 49.690 ;
        RECT 48.880 49.650 49.050 49.820 ;
        RECT 48.880 49.300 49.050 49.470 ;
        RECT 42.960 48.340 43.170 48.550 ;
        RECT 47.840 48.450 48.010 48.620 ;
        RECT 41.490 47.970 41.660 48.140 ;
        RECT 48.880 48.100 49.050 48.270 ;
        RECT 70.360 48.290 70.620 49.110 ;
        RECT 82.310 48.320 82.630 49.110 ;
        RECT 84.590 48.650 84.770 48.820 ;
        RECT 85.020 48.630 85.190 48.800 ;
        RECT 82.780 48.350 82.950 48.520 ;
        RECT 48.880 47.750 49.050 47.920 ;
        RECT 83.130 47.510 83.310 47.700 ;
        RECT 19.960 46.570 20.130 46.740 ;
        RECT 21.050 46.580 21.220 46.750 ;
        RECT 42.960 46.790 43.170 47.000 ;
        RECT 47.840 46.900 48.010 47.070 ;
        RECT 41.490 46.420 41.660 46.590 ;
        RECT 19.740 46.160 19.910 46.330 ;
        RECT 21.890 46.110 22.060 46.280 ;
        RECT 48.880 46.550 49.050 46.720 ;
        RECT 85.490 48.070 85.660 48.240 ;
        RECT 112.650 48.350 112.820 48.520 ;
        RECT 87.730 47.770 87.900 47.940 ;
        RECT 105.810 47.770 105.980 47.940 ;
        RECT 87.730 47.320 87.900 47.490 ;
        RECT 84.210 46.950 84.380 47.120 ;
        RECT 93.180 47.170 93.450 47.440 ;
        RECT 102.150 47.170 102.420 47.440 ;
        RECT 105.810 47.320 105.980 47.490 ;
        RECT 110.980 47.520 111.150 47.690 ;
        RECT 85.020 46.640 85.190 46.810 ;
        RECT 48.880 46.200 49.050 46.370 ;
        RECT 19.960 45.650 20.130 45.820 ;
        RECT 21.050 45.660 21.220 45.830 ;
        RECT 112.290 47.510 112.470 47.700 ;
        RECT 90.860 46.060 91.030 46.230 ;
        RECT 104.570 46.060 104.740 46.230 ;
        RECT 19.740 45.240 19.910 45.410 ;
        RECT 42.960 45.240 43.170 45.450 ;
        RECT 47.840 45.350 48.010 45.520 ;
        RECT 19.960 44.730 20.130 44.900 ;
        RECT 21.050 44.740 21.220 44.910 ;
        RECT 41.490 44.870 41.660 45.040 ;
        RECT 19.740 44.320 19.910 44.490 ;
        RECT 48.880 45.000 49.050 45.170 ;
        RECT 48.880 44.650 49.050 44.820 ;
        RECT 83.130 44.710 83.310 44.900 ;
        RECT 54.460 44.020 54.640 44.190 ;
        RECT 19.770 43.750 19.940 43.920 ;
        RECT 21.070 43.650 21.240 43.820 ;
        RECT 52.650 43.720 52.820 43.890 ;
        RECT 19.770 42.790 19.940 42.960 ;
        RECT 53.000 42.880 53.180 43.070 ;
        RECT 21.070 42.690 21.240 42.860 ;
        RECT 41.490 42.140 41.660 42.310 ;
        RECT 19.770 41.830 19.940 42.000 ;
        RECT 48.880 42.360 49.050 42.530 ;
        RECT 21.070 41.730 21.240 41.900 ;
        RECT 42.960 41.730 43.170 41.940 ;
        RECT 48.880 42.010 49.050 42.180 ;
        RECT 47.840 41.660 48.010 41.830 ;
        RECT 85.490 45.750 85.660 45.920 ;
        RECT 85.030 45.570 85.200 45.740 ;
        RECT 84.200 45.260 84.370 45.430 ;
        RECT 93.180 45.440 93.450 45.710 ;
        RECT 102.150 45.440 102.420 45.710 ;
        RECT 110.590 45.140 110.760 45.310 ;
        RECT 87.730 44.820 87.900 44.990 ;
        RECT 87.730 44.370 87.900 44.540 ;
        RECT 105.810 44.820 105.980 44.990 ;
        RECT 105.810 44.370 105.980 44.540 ;
        RECT 85.480 44.170 85.650 44.340 ;
        RECT 82.530 43.720 82.700 43.890 ;
        RECT 82.780 43.890 82.950 44.060 ;
        RECT 59.490 43.140 59.660 43.310 ;
        RECT 61.580 43.300 61.750 43.470 ;
        RECT 54.320 42.890 54.490 43.060 ;
        RECT 59.490 42.690 59.660 42.860 ;
        RECT 60.650 43.000 60.820 43.170 ;
        RECT 61.490 42.880 61.660 43.050 ;
        RECT 62.240 42.880 62.410 43.050 ;
        RECT 63.050 42.540 63.320 42.810 ;
        RECT 65.220 42.550 65.390 42.720 ;
        RECT 60.930 42.250 61.100 42.420 ;
        RECT 65.620 43.000 65.790 43.170 ;
        RECT 75.690 43.140 75.860 43.310 ;
        RECT 65.620 42.660 65.790 42.830 ;
        RECT 72.030 42.540 72.300 42.810 ;
        RECT 75.690 42.690 75.860 42.860 ;
        RECT 80.860 42.890 81.030 43.060 ;
        RECT 21.470 41.290 21.640 41.460 ;
        RECT 41.490 40.590 41.660 40.760 ;
        RECT 110.980 44.760 111.150 44.930 ;
        RECT 111.560 44.860 111.730 45.030 ;
        RECT 110.740 44.310 110.910 44.480 ;
        RECT 112.290 44.710 112.470 44.900 ;
        RECT 113.810 44.910 113.980 45.080 ;
        RECT 111.510 44.210 111.680 44.380 ;
        RECT 112.540 44.540 112.710 44.710 ;
        RECT 84.590 43.590 84.770 43.760 ;
        RECT 85.050 43.660 85.220 43.830 ;
        RECT 109.150 43.760 109.320 43.930 ;
        RECT 109.620 43.790 109.790 43.960 ;
        RECT 110.110 43.620 110.280 43.790 ;
        RECT 110.720 43.760 110.890 43.930 ;
        RECT 112.650 43.890 112.820 44.060 ;
        RECT 110.830 43.590 111.010 43.760 ;
        RECT 111.240 43.630 111.410 43.800 ;
        RECT 111.510 43.390 111.680 43.560 ;
        RECT 82.170 42.880 82.350 43.070 ;
        RECT 107.700 42.980 107.870 43.150 ;
        RECT 108.200 43.010 108.370 43.180 ;
        RECT 111.700 43.010 111.870 43.180 ;
        RECT 113.200 43.600 113.370 43.770 ;
        RECT 112.540 43.060 112.710 43.230 ;
        RECT 111.560 42.740 111.730 42.910 ;
        RECT 110.350 42.510 110.520 42.680 ;
        RECT 113.860 42.690 114.030 42.860 ;
        RECT 60.730 41.430 60.900 41.600 ;
        RECT 48.880 40.810 49.050 40.980 ;
        RECT 42.960 40.180 43.170 40.390 ;
        RECT 48.880 40.460 49.050 40.630 ;
        RECT 47.840 40.110 48.010 40.280 ;
        RECT 53.000 40.080 53.180 40.270 ;
        RECT 41.490 39.040 41.660 39.210 ;
        RECT 48.880 39.260 49.050 39.430 ;
        RECT 42.960 38.630 43.170 38.840 ;
        RECT 60.520 41.250 60.690 41.420 ;
        RECT 60.930 41.360 61.100 41.530 ;
        RECT 61.490 40.730 61.660 40.900 ;
        RECT 62.240 40.730 62.410 40.900 ;
        RECT 63.050 40.810 63.320 41.080 ;
        RECT 65.220 41.060 65.390 41.230 ;
        RECT 64.240 40.740 64.410 40.910 ;
        RECT 65.620 41.290 65.790 41.460 ;
        RECT 74.450 41.430 74.620 41.600 ;
        RECT 65.620 40.950 65.790 41.120 ;
        RECT 72.030 40.810 72.300 41.080 ;
        RECT 108.200 42.010 108.370 42.180 ;
        RECT 111.700 42.070 111.870 42.180 ;
        RECT 110.780 41.710 110.950 41.880 ;
        RECT 111.560 42.010 111.870 42.070 ;
        RECT 111.560 41.900 111.730 42.010 ;
        RECT 80.470 40.510 80.640 40.680 ;
        RECT 54.320 40.130 54.490 40.300 ;
        RECT 59.490 40.190 59.660 40.360 ;
        RECT 59.490 39.740 59.660 39.910 ;
        RECT 60.650 40.070 60.820 40.240 ;
        RECT 61.490 39.950 61.660 40.120 ;
        RECT 62.240 39.950 62.410 40.120 ;
        RECT 52.650 39.260 52.820 39.430 ;
        RECT 60.520 39.430 60.690 39.600 ;
        RECT 61.610 39.610 61.780 39.780 ;
        RECT 65.220 39.620 65.390 39.790 ;
        RECT 60.930 39.320 61.100 39.490 ;
        RECT 48.880 38.910 49.050 39.080 ;
        RECT 54.460 38.960 54.640 39.130 ;
        RECT 47.840 38.560 48.010 38.730 ;
        RECT 65.620 40.070 65.790 40.240 ;
        RECT 65.620 39.730 65.790 39.900 ;
        RECT 75.690 40.190 75.860 40.360 ;
        RECT 109.150 41.260 109.320 41.430 ;
        RECT 110.110 41.400 110.280 41.570 ;
        RECT 75.690 39.740 75.860 39.910 ;
        RECT 80.860 40.130 81.030 40.300 ;
        RECT 81.440 40.230 81.610 40.400 ;
        RECT 109.150 40.740 109.320 40.910 ;
        RECT 110.720 41.260 110.890 41.430 ;
        RECT 111.240 41.390 111.410 41.560 ;
        RECT 111.510 41.250 111.680 41.420 ;
        RECT 113.850 41.970 114.020 42.140 ;
        RECT 112.540 41.580 112.710 41.750 ;
        RECT 113.200 41.010 113.370 41.180 ;
        RECT 80.620 39.680 80.790 39.850 ;
        RECT 79.500 39.160 79.670 39.330 ;
        RECT 60.930 38.430 61.100 38.600 ;
        RECT 41.490 37.490 41.660 37.660 ;
        RECT 48.880 37.710 49.050 37.880 ;
        RECT 42.960 37.080 43.170 37.290 ;
        RECT 61.490 37.800 61.660 37.970 ;
        RECT 62.240 37.800 62.410 37.970 ;
        RECT 64.240 37.810 64.410 37.980 ;
        RECT 64.700 37.960 64.870 38.130 ;
        RECT 48.880 37.360 49.050 37.530 ;
        RECT 65.220 38.130 65.390 38.300 ;
        RECT 65.620 38.360 65.790 38.530 ;
        RECT 65.620 38.020 65.790 38.190 ;
        RECT 70.490 37.960 70.660 38.130 ;
        RECT 64.710 37.270 64.880 37.440 ;
        RECT 47.840 37.010 48.010 37.180 ;
        RECT 70.490 37.280 70.660 37.450 ;
        RECT 69.910 36.670 70.080 36.840 ;
        RECT 68.100 36.410 68.270 36.580 ;
        RECT 68.830 36.380 69.000 36.550 ;
        RECT 69.910 36.120 70.080 36.290 ;
        RECT 70.820 35.870 70.990 36.040 ;
        RECT 74.760 35.880 74.930 36.050 ;
        RECT 68.100 34.960 68.270 35.130 ;
        RECT 69.910 35.250 70.080 35.420 ;
        RECT 82.170 40.080 82.350 40.270 ;
        RECT 83.690 40.280 83.860 40.450 ;
        RECT 110.110 40.600 110.280 40.770 ;
        RECT 110.720 40.740 110.890 40.910 ;
        RECT 111.240 40.610 111.410 40.780 ;
        RECT 111.510 40.430 111.680 40.600 ;
        RECT 81.390 39.580 81.560 39.750 ;
        RECT 82.420 39.910 82.590 40.080 ;
        RECT 107.700 39.960 107.870 40.130 ;
        RECT 108.200 39.990 108.370 40.160 ;
        RECT 111.700 39.990 111.870 40.160 ;
        RECT 112.540 40.100 112.710 40.270 ;
        RECT 111.560 39.780 111.730 39.950 ;
        RECT 113.770 39.720 113.940 39.890 ;
        RECT 82.530 39.260 82.700 39.430 ;
        RECT 81.390 38.760 81.560 38.930 ;
        RECT 83.080 38.970 83.250 39.140 ;
        RECT 108.200 38.990 108.370 39.160 ;
        RECT 111.700 38.990 111.870 39.160 ;
        RECT 82.420 38.430 82.590 38.600 ;
        RECT 81.440 38.110 81.610 38.280 ;
        RECT 80.230 37.880 80.400 38.050 ;
        RECT 109.150 38.240 109.320 38.410 ;
        RECT 110.110 38.380 110.280 38.550 ;
        RECT 83.740 38.060 83.910 38.230 ;
        RECT 110.720 38.240 110.890 38.410 ;
        RECT 111.240 38.370 111.410 38.540 ;
        RECT 80.660 37.080 80.830 37.250 ;
        RECT 81.440 37.270 81.610 37.440 ;
        RECT 83.730 37.340 83.900 37.510 ;
        RECT 82.420 36.950 82.590 37.120 ;
        RECT 81.390 36.620 81.560 36.790 ;
        RECT 90.680 36.670 90.850 36.840 ;
        RECT 83.080 36.380 83.250 36.550 ;
        RECT 81.390 35.800 81.560 35.970 ;
        RECT 91.760 36.380 91.930 36.550 ;
        RECT 90.680 36.120 90.850 36.290 ;
        RECT 82.420 35.470 82.590 35.640 ;
        RECT 85.830 35.880 86.000 36.050 ;
        RECT 68.830 34.990 69.000 35.160 ;
        RECT 81.440 35.150 81.610 35.320 ;
        RECT 89.770 35.870 89.940 36.040 ;
        RECT 92.490 36.410 92.660 36.580 ;
        RECT 83.650 35.090 83.820 35.260 ;
        RECT 90.680 35.250 90.850 35.420 ;
        RECT 91.760 34.990 91.930 35.160 ;
        RECT 92.490 34.960 92.660 35.130 ;
        RECT 69.910 34.700 70.080 34.870 ;
        RECT 70.820 34.280 70.990 34.450 ;
        RECT 74.750 34.420 74.920 34.590 ;
        RECT 90.680 34.700 90.850 34.870 ;
        RECT 70.820 33.940 70.990 34.110 ;
        RECT 73.030 34.050 73.300 34.320 ;
        RECT 74.750 34.080 74.920 34.250 ;
        RECT 69.910 33.660 70.080 33.830 ;
        RECT 77.060 34.120 77.330 34.390 ;
        RECT 83.430 34.120 83.700 34.390 ;
        RECT 85.840 34.420 86.010 34.590 ;
        RECT 85.840 34.080 86.010 34.250 ;
        RECT 87.460 34.050 87.730 34.320 ;
        RECT 89.770 34.280 89.940 34.450 ;
        RECT 92.130 34.180 92.310 34.350 ;
        RECT 89.770 33.940 89.940 34.110 ;
        RECT 90.680 33.660 90.850 33.830 ;
        RECT 68.100 33.400 68.270 33.570 ;
        RECT 60.650 32.930 60.820 33.100 ;
        RECT 61.490 32.810 61.660 32.980 ;
        RECT 62.240 32.810 62.410 32.980 ;
        RECT 41.490 32.010 41.660 32.180 ;
        RECT 48.880 32.230 49.050 32.400 ;
        RECT 42.960 31.600 43.170 31.810 ;
        RECT 48.880 31.880 49.050 32.050 ;
        RECT 65.220 32.480 65.390 32.650 ;
        RECT 60.930 32.180 61.100 32.350 ;
        RECT 65.620 32.930 65.790 33.100 ;
        RECT 68.830 33.370 69.000 33.540 ;
        RECT 91.760 33.370 91.930 33.540 ;
        RECT 69.910 33.110 70.080 33.280 ;
        RECT 90.680 33.110 90.850 33.280 ;
        RECT 92.490 33.400 92.660 33.570 ;
        RECT 65.620 32.590 65.790 32.760 ;
        RECT 68.100 31.960 68.270 32.130 ;
        RECT 69.910 32.250 70.080 32.420 ;
        RECT 90.680 32.250 90.850 32.420 ;
        RECT 68.830 31.990 69.000 32.160 ;
        RECT 91.760 31.990 91.930 32.160 ;
        RECT 92.490 31.960 92.660 32.130 ;
        RECT 47.840 31.530 48.010 31.700 ;
        RECT 69.910 31.700 70.080 31.870 ;
        RECT 90.680 31.700 90.850 31.870 ;
        RECT 60.930 31.290 61.100 31.460 ;
        RECT 41.490 30.460 41.660 30.630 ;
        RECT 65.220 30.990 65.390 31.160 ;
        RECT 48.880 30.680 49.050 30.850 ;
        RECT 42.960 30.050 43.170 30.260 ;
        RECT 61.490 30.660 61.660 30.830 ;
        RECT 62.240 30.660 62.410 30.830 ;
        RECT 64.240 30.670 64.410 30.840 ;
        RECT 65.620 31.220 65.790 31.390 ;
        RECT 65.620 30.880 65.790 31.050 ;
        RECT 48.880 30.330 49.050 30.500 ;
        RECT 47.840 29.980 48.010 30.150 ;
        RECT 60.650 30.000 60.820 30.170 ;
        RECT 61.490 29.880 61.660 30.050 ;
        RECT 62.240 29.880 62.410 30.050 ;
        RECT 41.490 28.910 41.660 29.080 ;
        RECT 48.880 29.130 49.050 29.300 ;
        RECT 42.960 28.500 43.170 28.710 ;
        RECT 65.220 29.550 65.390 29.720 ;
        RECT 60.930 29.250 61.100 29.420 ;
        RECT 65.620 30.000 65.790 30.170 ;
        RECT 65.620 29.660 65.790 29.830 ;
        RECT 48.880 28.780 49.050 28.950 ;
        RECT 47.840 28.430 48.010 28.600 ;
        RECT 60.930 28.360 61.100 28.530 ;
        RECT 65.220 28.060 65.390 28.230 ;
        RECT 41.490 27.360 41.660 27.530 ;
        RECT 48.880 27.580 49.050 27.750 ;
        RECT 61.490 27.730 61.660 27.900 ;
        RECT 62.240 27.730 62.410 27.900 ;
        RECT 64.240 27.740 64.410 27.910 ;
        RECT 65.620 28.290 65.790 28.460 ;
        RECT 65.620 27.950 65.790 28.120 ;
        RECT 42.960 26.950 43.170 27.160 ;
        RECT 48.880 27.230 49.050 27.400 ;
        RECT 47.840 26.880 48.010 27.050 ;
        RECT 57.210 26.850 57.380 27.020 ;
        RECT 55.400 26.590 55.570 26.760 ;
        RECT 56.130 26.560 56.300 26.730 ;
        RECT 57.210 26.300 57.380 26.470 ;
        RECT 58.250 26.030 58.420 26.200 ;
        RECT 55.400 25.140 55.570 25.310 ;
        RECT 62.270 26.060 62.440 26.230 ;
        RECT 57.210 25.430 57.380 25.600 ;
        RECT 56.130 25.170 56.300 25.340 ;
        RECT 57.210 24.880 57.380 25.050 ;
        RECT 58.240 24.850 58.410 25.020 ;
        RECT 58.240 24.510 58.410 24.680 ;
        RECT 62.260 24.790 62.430 24.960 ;
        RECT 18.890 24.100 19.060 24.270 ;
        RECT 19.540 24.100 19.710 24.270 ;
        RECT 58.240 24.170 58.410 24.340 ;
        RECT 17.670 23.660 17.840 23.830 ;
        RECT 18.370 23.660 18.540 23.830 ;
        RECT 17.220 22.000 17.390 22.170 ;
        RECT 57.210 23.840 57.380 24.010 ;
        RECT 60.330 24.230 60.600 24.500 ;
        RECT 62.260 24.450 62.430 24.620 ;
        RECT 62.260 24.110 62.430 24.280 ;
        RECT 64.360 24.300 64.630 24.570 ;
        RECT 55.400 23.580 55.570 23.750 ;
        RECT 20.050 23.280 20.220 23.450 ;
        RECT 56.130 23.550 56.300 23.720 ;
        RECT 57.210 23.290 57.380 23.460 ;
        RECT 60.650 23.170 60.820 23.340 ;
        RECT 20.050 22.940 20.220 23.110 ;
        RECT 61.490 23.050 61.660 23.220 ;
        RECT 62.240 23.050 62.410 23.220 ;
        RECT 41.490 22.240 41.660 22.410 ;
        RECT 48.880 22.460 49.050 22.630 ;
        RECT 20.220 21.800 20.390 21.970 ;
        RECT 42.960 21.830 43.170 22.040 ;
        RECT 48.880 22.110 49.050 22.280 ;
        RECT 55.400 22.140 55.570 22.310 ;
        RECT 57.210 22.430 57.380 22.600 ;
        RECT 56.130 22.170 56.300 22.340 ;
        RECT 65.220 22.720 65.390 22.890 ;
        RECT 60.930 22.420 61.100 22.590 ;
        RECT 65.620 23.170 65.790 23.340 ;
        RECT 65.620 22.830 65.790 23.000 ;
        RECT 68.550 22.950 68.720 23.120 ;
        RECT 68.700 22.270 68.870 22.440 ;
        RECT 70.850 22.390 71.020 22.560 ;
        RECT 47.840 21.760 48.010 21.930 ;
        RECT 57.210 21.880 57.380 22.050 ;
        RECT 69.590 21.820 69.760 21.990 ;
        RECT 20.230 21.260 20.400 21.430 ;
        RECT 60.930 21.530 61.100 21.700 ;
        RECT 17.700 19.780 17.870 19.950 ;
        RECT 41.490 20.690 41.660 20.860 ;
        RECT 65.220 21.230 65.390 21.400 ;
        RECT 20.040 20.300 20.210 20.470 ;
        RECT 48.880 20.910 49.050 21.080 ;
        RECT 42.960 20.280 43.170 20.490 ;
        RECT 61.490 20.900 61.660 21.070 ;
        RECT 62.240 20.900 62.410 21.070 ;
        RECT 64.240 20.910 64.410 21.080 ;
        RECT 65.620 21.460 65.790 21.630 ;
        RECT 68.700 21.370 68.870 21.540 ;
        RECT 65.620 21.120 65.790 21.290 ;
        RECT 70.850 21.250 71.020 21.420 ;
        RECT 48.880 20.560 49.050 20.730 ;
        RECT 68.550 20.690 68.720 20.860 ;
        RECT 47.840 20.210 48.010 20.380 ;
        RECT 60.650 20.240 60.820 20.410 ;
        RECT 61.490 20.120 61.660 20.290 ;
        RECT 62.240 20.120 62.410 20.290 ;
        RECT 18.390 19.770 18.560 19.940 ;
        RECT 18.870 19.000 19.040 19.170 ;
        RECT 41.490 19.140 41.660 19.310 ;
        RECT 19.580 18.940 19.750 19.110 ;
        RECT 48.880 19.360 49.050 19.530 ;
        RECT 42.960 18.730 43.170 18.940 ;
        RECT 65.220 19.790 65.390 19.960 ;
        RECT 60.930 19.490 61.100 19.660 ;
        RECT 65.620 20.240 65.790 20.410 ;
        RECT 68.550 20.180 68.720 20.350 ;
        RECT 65.620 19.900 65.790 20.070 ;
        RECT 68.700 19.500 68.870 19.670 ;
        RECT 70.850 19.620 71.020 19.790 ;
        RECT 48.880 19.010 49.050 19.180 ;
        RECT 69.590 19.050 69.760 19.220 ;
        RECT 47.840 18.660 48.010 18.830 ;
        RECT 57.110 18.540 57.280 18.710 ;
        RECT 19.540 18.120 19.710 18.290 ;
        RECT 16.230 17.680 16.400 17.850 ;
        RECT 17.330 17.690 17.500 17.860 ;
        RECT 16.780 17.010 16.950 17.180 ;
        RECT 16.780 15.640 16.950 15.810 ;
        RECT 16.230 14.910 16.400 15.080 ;
        RECT 16.220 13.570 16.390 13.740 ;
        RECT 18.420 17.690 18.590 17.860 ;
        RECT 17.880 17.010 18.050 17.180 ;
        RECT 17.880 15.640 18.050 15.810 ;
        RECT 17.330 14.910 17.500 15.080 ;
        RECT 17.330 13.560 17.500 13.730 ;
        RECT 16.780 12.870 16.950 13.040 ;
        RECT 19.550 17.650 19.720 17.820 ;
        RECT 41.490 17.590 41.660 17.760 ;
        RECT 48.880 17.810 49.050 17.980 ;
        RECT 18.980 17.010 19.150 17.180 ;
        RECT 42.960 17.180 43.170 17.390 ;
        RECT 60.930 18.600 61.100 18.770 ;
        RECT 65.220 18.300 65.390 18.470 ;
        RECT 57.160 17.690 57.330 17.860 ;
        RECT 61.490 17.970 61.660 18.140 ;
        RECT 62.240 17.970 62.410 18.140 ;
        RECT 64.240 17.980 64.410 18.150 ;
        RECT 65.620 18.530 65.790 18.700 ;
        RECT 68.700 18.600 68.870 18.770 ;
        RECT 65.620 18.190 65.790 18.360 ;
        RECT 70.850 18.480 71.020 18.650 ;
        RECT 68.550 17.920 68.720 18.090 ;
        RECT 48.880 17.460 49.050 17.630 ;
        RECT 19.670 16.990 19.840 17.160 ;
        RECT 47.840 17.110 48.010 17.280 ;
        RECT 19.670 16.650 19.840 16.820 ;
        RECT 19.670 16.310 19.840 16.480 ;
        RECT 18.980 15.640 19.150 15.810 ;
        RECT 18.420 14.910 18.590 15.080 ;
        RECT 18.420 13.540 18.590 13.710 ;
        RECT 17.880 12.860 18.050 13.030 ;
        RECT 26.250 13.740 26.420 14.080 ;
        RECT 26.590 13.740 26.760 14.080 ;
        RECT 18.970 12.860 19.140 13.030 ;
        RECT 19.580 10.560 19.750 10.730 ;
        RECT 16.270 10.120 16.440 10.290 ;
        RECT 17.370 10.130 17.540 10.300 ;
        RECT 18.460 10.130 18.630 10.300 ;
        RECT 16.820 9.450 16.990 9.620 ;
        RECT 17.920 9.450 18.090 9.620 ;
        RECT 16.820 8.080 16.990 8.250 ;
        RECT 17.920 8.080 18.090 8.250 ;
        RECT 19.590 10.090 19.760 10.260 ;
        RECT 19.020 9.450 19.190 9.620 ;
        RECT 19.020 8.080 19.190 8.250 ;
        RECT 49.180 11.400 49.350 11.570 ;
        RECT 50.270 11.400 50.440 11.570 ;
        RECT 49.730 10.720 49.900 10.890 ;
        RECT 49.730 9.350 49.900 9.520 ;
        RECT 52.490 11.570 52.660 11.740 ;
        RECT 51.370 11.390 51.540 11.560 ;
        RECT 52.490 11.230 52.660 11.400 ;
        RECT 54.380 11.570 54.550 11.740 ;
        RECT 54.380 11.230 54.550 11.400 ;
        RECT 55.500 11.390 55.670 11.560 ;
        RECT 56.600 11.400 56.770 11.570 ;
        RECT 50.820 10.700 50.990 10.870 ;
        RECT 51.930 10.690 52.100 10.860 ;
        RECT 54.940 10.690 55.110 10.860 ;
        RECT 56.050 10.700 56.220 10.870 ;
        RECT 50.820 9.350 50.990 9.520 ;
        RECT 51.920 9.350 52.090 9.520 ;
        RECT 54.950 9.350 55.120 9.520 ;
        RECT 56.050 9.350 56.220 9.520 ;
        RECT 57.690 11.400 57.860 11.570 ;
        RECT 57.140 10.720 57.310 10.890 ;
        RECT 57.140 9.350 57.310 9.520 ;
        RECT 58.990 11.430 59.160 11.600 ;
        RECT 60.080 11.430 60.250 11.600 ;
        RECT 59.540 10.750 59.710 10.920 ;
        RECT 59.540 9.380 59.710 9.550 ;
        RECT 62.300 11.600 62.470 11.770 ;
        RECT 61.180 11.420 61.350 11.590 ;
        RECT 62.300 11.260 62.470 11.430 ;
        RECT 64.190 11.600 64.360 11.770 ;
        RECT 64.190 11.260 64.360 11.430 ;
        RECT 65.310 11.420 65.480 11.590 ;
        RECT 66.410 11.430 66.580 11.600 ;
        RECT 60.630 10.730 60.800 10.900 ;
        RECT 61.740 10.720 61.910 10.890 ;
        RECT 64.750 10.720 64.920 10.890 ;
        RECT 65.860 10.730 66.030 10.900 ;
        RECT 60.630 9.380 60.800 9.550 ;
        RECT 61.730 9.380 61.900 9.550 ;
        RECT 64.760 9.380 64.930 9.550 ;
        RECT 65.860 9.380 66.030 9.550 ;
        RECT 67.500 11.430 67.670 11.600 ;
        RECT 66.950 10.750 67.120 10.920 ;
        RECT 66.950 9.380 67.120 9.550 ;
        RECT 71.050 11.400 71.220 11.570 ;
        RECT 70.490 10.700 70.660 10.870 ;
        RECT 70.500 9.360 70.670 9.530 ;
        RECT 16.270 7.350 16.440 7.520 ;
        RECT 17.370 7.350 17.540 7.520 ;
        RECT 16.260 6.010 16.430 6.180 ;
        RECT 17.370 6.000 17.540 6.170 ;
        RECT 15.700 5.470 15.870 5.640 ;
        RECT 16.820 5.310 16.990 5.480 ;
        RECT 18.460 7.350 18.630 7.520 ;
        RECT 18.460 5.980 18.630 6.150 ;
        RECT 17.920 5.300 18.090 5.470 ;
        RECT 19.010 5.300 19.180 5.470 ;
        RECT 49.170 8.620 49.340 8.790 ;
        RECT 49.170 7.250 49.340 7.420 ;
        RECT 48.600 6.610 48.770 6.780 ;
        RECT 50.270 8.620 50.440 8.790 ;
        RECT 51.370 8.620 51.540 8.790 ;
        RECT 55.500 8.620 55.670 8.790 ;
        RECT 56.600 8.620 56.770 8.790 ;
        RECT 50.270 7.250 50.440 7.420 ;
        RECT 51.370 7.250 51.540 7.420 ;
        RECT 55.500 7.250 55.670 7.420 ;
        RECT 56.600 7.250 56.770 7.420 ;
        RECT 49.730 6.570 49.900 6.740 ;
        RECT 50.820 6.570 50.990 6.740 ;
        RECT 51.920 6.580 52.090 6.750 ;
        RECT 54.950 6.580 55.120 6.750 ;
        RECT 56.050 6.570 56.220 6.740 ;
        RECT 57.700 8.620 57.870 8.790 ;
        RECT 57.700 7.250 57.870 7.420 ;
        RECT 57.140 6.570 57.310 6.740 ;
        RECT 58.980 8.650 59.150 8.820 ;
        RECT 58.980 7.280 59.150 7.450 ;
        RECT 58.410 6.780 58.580 6.810 ;
        RECT 58.270 6.640 58.580 6.780 ;
        RECT 58.270 6.610 58.440 6.640 ;
        RECT 60.080 8.650 60.250 8.820 ;
        RECT 61.180 8.650 61.350 8.820 ;
        RECT 65.310 8.650 65.480 8.820 ;
        RECT 66.410 8.650 66.580 8.820 ;
        RECT 60.080 7.280 60.250 7.450 ;
        RECT 61.180 7.280 61.350 7.450 ;
        RECT 65.310 7.280 65.480 7.450 ;
        RECT 66.410 7.280 66.580 7.450 ;
        RECT 48.610 6.140 48.780 6.310 ;
        RECT 59.540 6.600 59.710 6.770 ;
        RECT 60.630 6.600 60.800 6.770 ;
        RECT 61.730 6.610 61.900 6.780 ;
        RECT 64.760 6.610 64.930 6.780 ;
        RECT 65.860 6.600 66.030 6.770 ;
        RECT 67.510 8.650 67.680 8.820 ;
        RECT 67.510 7.280 67.680 7.450 ;
        RECT 66.950 6.600 67.120 6.770 ;
        RECT 68.080 6.640 68.250 6.810 ;
        RECT 72.150 11.410 72.320 11.580 ;
        RECT 71.600 10.710 71.770 10.880 ;
        RECT 71.600 9.360 71.770 9.530 ;
        RECT 71.050 8.630 71.220 8.800 ;
        RECT 71.050 7.260 71.220 7.430 ;
        RECT 58.420 6.310 58.590 6.340 ;
        RECT 58.260 6.170 58.590 6.310 ;
        RECT 58.260 6.140 58.430 6.170 ;
        RECT 70.500 6.590 70.670 6.760 ;
        RECT 73.240 11.410 73.410 11.580 ;
        RECT 72.690 10.730 72.860 10.900 ;
        RECT 72.690 9.360 72.860 9.530 ;
        RECT 72.150 8.630 72.320 8.800 ;
        RECT 72.150 7.260 72.320 7.430 ;
        RECT 71.600 6.580 71.770 6.750 ;
        RECT 73.250 8.630 73.420 8.800 ;
        RECT 73.940 8.300 74.110 8.470 ;
        RECT 73.940 7.960 74.110 8.130 ;
        RECT 73.940 7.620 74.110 7.790 ;
        RECT 73.250 7.260 73.420 7.430 ;
        RECT 72.690 6.580 72.860 6.750 ;
        RECT 73.820 6.620 73.990 6.790 ;
        RECT 68.070 6.170 68.240 6.340 ;
        RECT 73.810 6.150 73.980 6.320 ;
        RECT 20.410 1.770 20.580 5.290 ;
        RECT 20.780 1.770 20.950 5.290 ;
        RECT 21.130 1.770 21.300 5.290 ;
        RECT 21.470 1.770 21.640 5.290 ;
        RECT 21.820 1.770 21.990 5.290 ;
        RECT 22.180 1.770 22.350 5.290 ;
        RECT 22.540 1.770 22.710 5.290 ;
        RECT 99.180 4.000 99.350 4.170 ;
        RECT 104.700 3.260 104.870 3.430 ;
        RECT 99.180 2.390 99.350 2.560 ;
        RECT 104.700 2.590 104.870 2.760 ;
        RECT 99.180 0.790 99.350 0.960 ;
        RECT 99.180 -0.830 99.350 -0.660 ;
        RECT 101.710 -2.040 101.880 -1.870 ;
        RECT 99.180 -2.430 99.350 -2.260 ;
        RECT 99.180 -4.050 99.350 -3.880 ;
        RECT 99.180 -5.650 99.350 -5.480 ;
        RECT 110.780 -5.440 110.950 9.510 ;
        RECT 99.180 -7.270 99.350 -7.100 ;
      LAYER met1 ;
        RECT 82.330 66.110 82.670 66.250 ;
        RECT 90.210 66.110 90.930 67.850 ;
        RECT 82.330 65.390 90.930 66.110 ;
        RECT 30.260 62.940 31.600 63.390 ;
        RECT 4.160 62.100 4.660 62.580 ;
        RECT 30.260 62.520 43.780 62.940 ;
        RECT 45.570 62.850 48.760 63.970 ;
        RECT 30.260 62.380 31.600 62.520 ;
        RECT 4.260 59.140 4.650 62.100 ;
        RECT 24.850 61.780 27.620 62.020 ;
        RECT 6.630 61.320 6.890 61.520 ;
        RECT 9.490 61.480 9.750 61.570 ;
        RECT 6.570 61.010 6.950 61.320 ;
        RECT 7.980 61.010 9.010 61.320 ;
        RECT 9.480 61.250 9.770 61.480 ;
        RECT 6.620 60.220 6.880 60.490 ;
        RECT 7.310 60.220 7.630 60.460 ;
        RECT 8.030 60.220 8.290 60.500 ;
        RECT 6.580 59.560 8.330 60.220 ;
        RECT 6.620 59.300 6.880 59.560 ;
        RECT 7.310 59.300 7.630 59.560 ;
        RECT 8.050 59.320 8.310 59.560 ;
        RECT 4.260 58.650 4.730 59.140 ;
        RECT 4.260 58.640 4.710 58.650 ;
        RECT 4.260 0.530 4.650 58.640 ;
        RECT 6.640 58.270 6.870 58.790 ;
        RECT 6.620 57.950 6.880 58.270 ;
        RECT 5.670 57.500 5.930 57.820 ;
        RECT 5.680 55.280 5.920 57.500 ;
        RECT 6.640 57.380 6.870 57.950 ;
        RECT 8.050 57.380 8.280 58.790 ;
        RECT 8.770 58.240 9.010 61.010 ;
        RECT 24.850 60.690 25.090 61.780 ;
        RECT 9.430 60.560 9.820 60.690 ;
        RECT 9.430 60.270 9.850 60.560 ;
        RECT 24.850 60.430 25.080 60.690 ;
        RECT 9.150 59.710 9.470 60.030 ;
        RECT 9.200 59.480 9.430 59.710 ;
        RECT 9.620 59.330 9.850 60.270 ;
        RECT 24.840 60.210 25.080 60.430 ;
        RECT 22.700 59.400 23.020 59.720 ;
        RECT 24.060 59.480 24.380 59.800 ;
        RECT 24.750 59.470 25.070 59.790 ;
        RECT 9.490 59.260 9.850 59.330 ;
        RECT 9.430 59.150 9.850 59.260 ;
        RECT 9.430 59.030 9.820 59.150 ;
        RECT 8.730 57.700 9.050 58.020 ;
        RECT 9.490 57.860 9.760 59.030 ;
        RECT 24.850 57.890 25.090 58.530 ;
        RECT 9.490 57.630 9.820 57.860 ;
        RECT 24.850 57.630 25.080 57.890 ;
        RECT 24.840 56.980 25.080 57.630 ;
        RECT 7.290 56.500 7.610 56.820 ;
        RECT 8.720 56.520 9.040 56.840 ;
        RECT 6.500 55.920 6.820 56.240 ;
        RECT 7.430 55.920 7.750 56.240 ;
        RECT 8.130 55.920 8.450 56.240 ;
        RECT 8.870 55.920 9.190 56.240 ;
        RECT 9.580 55.910 9.900 56.230 ;
        RECT 5.590 54.800 6.010 55.280 ;
        RECT 11.480 54.040 11.770 56.730 ;
        RECT 24.840 56.340 25.090 56.980 ;
        RECT 21.980 55.740 22.300 56.060 ;
        RECT 11.460 53.370 11.870 54.040 ;
        RECT 24.840 52.680 25.080 56.340 ;
        RECT 24.790 52.340 25.130 52.680 ;
        RECT 22.040 52.240 22.530 52.250 ;
        RECT 18.110 43.550 18.340 47.030 ;
        RECT 18.780 46.410 19.000 47.030 ;
        RECT 19.890 46.500 20.210 46.820 ;
        RECT 20.980 46.510 21.300 46.830 ;
        RECT 18.750 46.090 19.010 46.410 ;
        RECT 19.420 46.360 19.740 46.410 ;
        RECT 19.420 46.130 19.970 46.360 ;
        RECT 19.420 46.090 19.740 46.130 ;
        RECT 18.780 45.490 19.000 46.090 ;
        RECT 19.890 45.580 20.210 45.900 ;
        RECT 20.980 45.590 21.300 45.910 ;
        RECT 18.720 45.170 19.000 45.490 ;
        RECT 19.420 45.440 19.740 45.490 ;
        RECT 19.420 45.210 19.970 45.440 ;
        RECT 19.420 45.170 19.740 45.210 ;
        RECT 18.780 44.570 19.000 45.170 ;
        RECT 19.890 44.660 20.210 44.980 ;
        RECT 20.980 44.670 21.300 44.990 ;
        RECT 18.730 44.250 19.000 44.570 ;
        RECT 19.420 44.520 19.740 44.570 ;
        RECT 19.420 44.290 19.970 44.520 ;
        RECT 19.420 44.250 19.740 44.290 ;
        RECT 18.080 43.230 18.340 43.550 ;
        RECT 18.110 42.590 18.340 43.230 ;
        RECT 18.040 42.270 18.340 42.590 ;
        RECT 18.110 41.630 18.340 42.270 ;
        RECT 18.080 41.310 18.340 41.630 ;
        RECT 18.110 26.560 18.340 41.310 ;
        RECT 18.780 26.560 19.000 44.250 ;
        RECT 19.700 43.680 20.020 44.000 ;
        RECT 21.000 43.580 21.320 43.900 ;
        RECT 19.700 43.500 20.020 43.540 ;
        RECT 19.470 43.270 20.020 43.500 ;
        RECT 19.700 43.220 20.020 43.270 ;
        RECT 19.700 42.720 20.020 43.040 ;
        RECT 21.000 42.620 21.320 42.940 ;
        RECT 19.700 42.540 20.020 42.580 ;
        RECT 19.470 42.310 20.020 42.540 ;
        RECT 19.700 42.260 20.020 42.310 ;
        RECT 19.700 41.760 20.020 42.080 ;
        RECT 21.000 41.660 21.320 41.980 ;
        RECT 19.700 41.580 20.020 41.620 ;
        RECT 19.470 41.350 20.020 41.580 ;
        RECT 21.470 41.490 21.690 51.300 ;
        RECT 22.030 51.090 22.540 52.240 ;
        RECT 27.380 51.310 27.620 61.780 ;
        RECT 30.690 61.450 33.720 61.720 ;
        RECT 30.690 60.470 30.960 61.450 ;
        RECT 30.700 58.260 30.960 58.280 ;
        RECT 30.660 52.280 30.970 58.260 ;
        RECT 31.840 55.760 32.160 56.080 ;
        RECT 30.580 51.910 30.970 52.280 ;
        RECT 33.450 51.770 33.720 61.450 ;
        RECT 35.400 60.430 35.660 62.520 ;
        RECT 43.360 59.270 43.780 62.520 ;
        RECT 47.170 60.030 47.590 62.850 ;
        RECT 47.170 59.550 47.640 60.030 ;
        RECT 43.320 58.790 43.800 59.270 ;
        RECT 34.630 57.720 34.860 57.890 ;
        RECT 34.620 55.850 34.870 57.720 ;
        RECT 48.870 57.180 49.310 57.680 ;
        RECT 54.590 57.180 55.030 57.680 ;
        RECT 44.450 56.160 44.890 56.660 ;
        RECT 34.620 55.670 34.880 55.850 ;
        RECT 34.620 52.770 34.870 55.670 ;
        RECT 41.660 53.420 41.980 53.470 ;
        RECT 41.570 53.130 41.980 53.420 ;
        RECT 34.580 52.410 34.910 52.770 ;
        RECT 33.410 51.460 33.750 51.770 ;
        RECT 21.980 50.990 22.540 51.090 ;
        RECT 27.330 50.990 27.670 51.310 ;
        RECT 21.870 50.590 22.540 50.990 ;
        RECT 41.270 50.840 41.510 50.890 ;
        RECT 21.870 50.560 22.530 50.590 ;
        RECT 21.870 46.340 22.090 50.560 ;
        RECT 41.570 50.490 41.810 53.130 ;
        RECT 44.510 50.890 44.820 56.160 ;
        RECT 44.210 50.820 44.820 50.890 ;
        RECT 48.640 50.840 48.930 50.890 ;
        RECT 44.510 50.490 44.820 50.820 ;
        RECT 48.940 50.490 49.230 57.180 ;
        RECT 50.130 56.190 50.630 56.630 ;
        RECT 41.460 49.630 41.810 50.490 ;
        RECT 42.880 49.850 43.230 50.140 ;
        RECT 42.880 49.830 43.080 49.850 ;
        RECT 40.720 48.990 41.130 49.320 ;
        RECT 23.090 48.440 23.440 48.900 ;
        RECT 39.520 48.460 39.890 48.770 ;
        RECT 22.490 48.080 22.740 48.200 ;
        RECT 22.460 47.620 22.780 48.080 ;
        RECT 21.860 46.050 22.090 46.340 ;
        RECT 19.700 41.300 20.020 41.350 ;
        RECT 21.410 41.260 21.700 41.490 ;
        RECT 18.000 26.030 18.340 26.560 ;
        RECT 18.660 26.030 19.000 26.560 ;
        RECT 16.690 25.290 16.920 25.360 ;
        RECT 16.650 25.030 16.970 25.290 ;
        RECT 16.200 24.920 16.430 24.960 ;
        RECT 16.160 24.600 16.430 24.920 ;
        RECT 6.850 23.360 7.570 24.060 ;
        RECT 6.860 18.210 7.520 23.360 ;
        RECT 16.200 21.080 16.430 24.600 ;
        RECT 16.690 22.560 16.920 25.030 ;
        RECT 18.110 24.940 18.340 26.030 ;
        RECT 18.780 25.300 19.000 26.030 ;
        RECT 20.540 25.320 20.810 25.360 ;
        RECT 18.760 24.980 19.020 25.300 ;
        RECT 20.520 24.990 20.810 25.320 ;
        RECT 18.100 24.620 18.360 24.940 ;
        RECT 18.820 24.020 19.140 24.340 ;
        RECT 19.470 24.020 19.790 24.340 ;
        RECT 17.600 23.580 17.920 23.900 ;
        RECT 18.300 23.580 18.620 23.900 ;
        RECT 19.990 22.570 20.280 23.480 ;
        RECT 16.690 22.550 17.420 22.560 ;
        RECT 16.690 22.230 17.440 22.550 ;
        RECT 16.690 22.190 17.420 22.230 ;
        RECT 16.200 21.010 16.460 21.080 ;
        RECT 16.180 21.000 16.460 21.010 ;
        RECT 16.150 20.690 16.470 21.000 ;
        RECT 12.050 18.830 12.480 19.260 ;
        RECT 6.860 17.490 7.600 18.210 ;
        RECT 12.100 13.020 12.470 18.830 ;
        RECT 16.150 17.600 16.470 17.920 ;
        RECT 16.690 17.250 16.920 22.190 ;
        RECT 17.190 21.940 17.420 22.190 ;
        RECT 19.900 22.000 20.220 22.040 ;
        RECT 20.540 22.020 20.810 24.990 ;
        RECT 20.420 22.000 20.810 22.020 ;
        RECT 17.190 21.720 17.410 21.940 ;
        RECT 19.900 21.770 20.810 22.000 ;
        RECT 21.020 24.920 21.260 24.960 ;
        RECT 21.020 24.600 21.280 24.920 ;
        RECT 19.900 21.720 20.220 21.770 ;
        RECT 17.210 21.290 17.430 21.510 ;
        RECT 17.200 21.000 17.430 21.290 ;
        RECT 19.910 21.460 20.230 21.500 ;
        RECT 21.020 21.460 21.260 24.600 ;
        RECT 19.910 21.230 21.260 21.460 ;
        RECT 19.910 21.180 20.230 21.230 ;
        RECT 17.180 20.680 17.440 21.000 ;
        RECT 19.980 20.550 20.250 20.730 ;
        RECT 19.960 20.230 20.280 20.550 ;
        RECT 19.980 20.060 20.250 20.230 ;
        RECT 17.630 19.700 17.950 20.020 ;
        RECT 18.320 19.690 18.640 20.010 ;
        RECT 18.800 18.920 19.120 19.240 ;
        RECT 19.510 18.860 19.830 19.180 ;
        RECT 19.460 18.040 19.780 18.360 ;
        RECT 17.250 17.610 17.570 17.930 ;
        RECT 18.340 17.610 18.660 17.930 ;
        RECT 19.470 17.570 19.790 17.890 ;
        RECT 16.690 16.930 17.020 17.250 ;
        RECT 17.800 16.930 18.120 17.250 ;
        RECT 18.900 16.930 19.220 17.250 ;
        RECT 16.690 15.880 16.920 16.930 ;
        RECT 19.610 16.760 19.900 17.190 ;
        RECT 19.610 16.740 20.080 16.760 ;
        RECT 19.620 16.440 20.080 16.740 ;
        RECT 19.620 15.910 19.900 16.440 ;
        RECT 16.690 15.560 17.020 15.880 ;
        RECT 17.800 15.560 18.120 15.880 ;
        RECT 18.900 15.560 19.220 15.880 ;
        RECT 16.150 14.830 16.470 15.150 ;
        RECT 16.690 14.690 16.920 15.560 ;
        RECT 17.250 14.830 17.570 15.150 ;
        RECT 18.340 14.830 18.660 15.150 ;
        RECT 16.690 14.460 19.140 14.690 ;
        RECT 18.820 14.130 19.140 14.460 ;
        RECT 16.140 13.490 16.460 13.810 ;
        RECT 17.250 13.480 17.570 13.800 ;
        RECT 18.340 13.460 18.660 13.780 ;
        RECT 12.060 12.590 12.490 13.020 ;
        RECT 16.700 12.790 17.020 13.110 ;
        RECT 17.800 12.780 18.120 13.100 ;
        RECT 18.890 12.780 19.210 13.100 ;
        RECT 19.580 12.560 19.910 12.590 ;
        RECT 19.440 12.480 19.910 12.560 ;
        RECT 19.200 12.240 19.910 12.480 ;
        RECT 19.580 12.170 19.910 12.240 ;
        RECT 15.070 6.930 15.360 7.280 ;
        RECT 15.080 6.360 15.340 6.930 ;
        RECT 15.720 5.830 15.980 10.810 ;
        RECT 19.500 10.480 19.820 10.800 ;
        RECT 16.190 10.040 16.510 10.360 ;
        RECT 17.290 10.050 17.610 10.370 ;
        RECT 18.380 10.050 18.700 10.370 ;
        RECT 19.510 10.010 19.830 10.330 ;
        RECT 16.740 9.370 17.060 9.690 ;
        RECT 17.840 9.370 18.160 9.690 ;
        RECT 18.940 9.370 19.260 9.690 ;
        RECT 16.740 8.000 17.060 8.320 ;
        RECT 17.840 8.000 18.160 8.320 ;
        RECT 18.940 8.000 19.260 8.320 ;
        RECT 16.190 7.270 16.510 7.590 ;
        RECT 17.290 7.270 17.610 7.590 ;
        RECT 18.380 7.270 18.700 7.590 ;
        RECT 21.020 6.570 21.260 21.230 ;
        RECT 21.470 20.560 21.690 41.260 ;
        RECT 21.870 23.170 22.090 46.050 ;
        RECT 22.490 46.830 22.740 47.620 ;
        RECT 22.490 46.510 22.780 46.830 ;
        RECT 22.490 45.910 22.740 46.510 ;
        RECT 22.490 45.590 22.780 45.910 ;
        RECT 22.490 44.990 22.740 45.590 ;
        RECT 22.490 44.670 22.750 44.990 ;
        RECT 22.490 24.320 22.740 44.670 ;
        RECT 23.110 43.900 23.370 48.440 ;
        RECT 38.880 46.740 39.270 47.110 ;
        RECT 38.300 45.250 38.690 45.640 ;
        RECT 23.110 43.580 23.390 43.900 ;
        RECT 37.660 43.660 38.050 44.040 ;
        RECT 37.690 43.650 38.030 43.660 ;
        RECT 23.110 42.940 23.370 43.580 ;
        RECT 37.050 43.460 37.390 43.470 ;
        RECT 37.040 43.070 37.400 43.460 ;
        RECT 23.110 42.620 23.400 42.940 ;
        RECT 23.110 41.980 23.370 42.620 ;
        RECT 23.110 41.660 23.390 41.980 ;
        RECT 22.490 24.300 22.750 24.320 ;
        RECT 22.480 24.020 22.760 24.300 ;
        RECT 22.490 24.000 22.750 24.020 ;
        RECT 21.830 22.850 22.150 23.170 ;
        RECT 21.430 20.240 21.710 20.560 ;
        RECT 21.470 7.270 21.690 20.240 ;
        RECT 21.870 15.030 22.090 22.850 ;
        RECT 21.870 14.550 22.160 15.030 ;
        RECT 21.870 12.590 22.090 14.550 ;
        RECT 21.850 12.170 22.110 12.590 ;
        RECT 21.870 7.550 22.090 12.170 ;
        RECT 22.490 8.930 22.740 24.000 ;
        RECT 23.110 19.990 23.370 41.660 ;
        RECT 36.430 41.510 36.790 41.900 ;
        RECT 35.780 39.970 36.190 40.370 ;
        RECT 35.250 38.410 35.610 38.800 ;
        RECT 34.670 33.350 35.000 33.370 ;
        RECT 34.610 32.930 35.000 33.350 ;
        RECT 34.040 31.740 34.370 31.760 ;
        RECT 33.990 31.350 34.380 31.740 ;
        RECT 33.420 30.190 33.750 30.200 ;
        RECT 33.390 29.800 33.750 30.190 ;
        RECT 32.770 28.320 33.160 28.720 ;
        RECT 32.100 23.150 32.530 23.550 ;
        RECT 31.440 21.580 31.850 21.980 ;
        RECT 23.100 19.670 23.410 19.990 ;
        RECT 30.830 19.940 31.220 20.340 ;
        RECT 22.450 8.530 22.750 8.930 ;
        RECT 21.870 7.410 22.110 7.550 ;
        RECT 21.430 6.920 21.740 7.270 ;
        RECT 21.880 6.780 22.110 7.410 ;
        RECT 16.180 5.930 16.500 6.250 ;
        RECT 17.290 5.920 17.610 6.240 ;
        RECT 18.380 5.900 18.700 6.220 ;
        RECT 20.230 6.010 21.260 6.570 ;
        RECT 21.870 6.750 22.110 6.780 ;
        RECT 20.230 5.900 21.020 6.010 ;
        RECT 15.670 5.020 15.980 5.830 ;
        RECT 16.740 5.230 17.060 5.550 ;
        RECT 17.840 5.220 18.160 5.540 ;
        RECT 18.930 5.220 19.250 5.540 ;
        RECT 21.870 5.360 22.090 6.750 ;
        RECT 15.720 4.820 15.980 5.020 ;
        RECT 20.340 1.680 22.760 5.360 ;
        RECT 23.110 1.390 23.370 19.670 ;
        RECT 30.140 18.500 30.550 18.890 ;
        RECT 25.930 13.350 26.860 15.000 ;
        RECT 26.020 12.870 26.760 13.350 ;
        RECT 23.020 0.980 23.370 1.390 ;
        RECT 4.090 0.010 4.650 0.530 ;
        RECT 30.200 -4.840 30.530 18.500 ;
        RECT 30.150 -4.850 30.580 -4.840 ;
        RECT 30.120 -5.310 30.610 -4.850 ;
        RECT 30.150 -5.330 30.580 -5.310 ;
        RECT 30.850 -5.630 31.180 19.940 ;
        RECT 30.760 -6.120 31.250 -5.630 ;
        RECT 31.500 -6.340 31.830 21.580 ;
        RECT 31.470 -6.800 31.870 -6.340 ;
        RECT 31.260 -7.290 31.840 -7.180 ;
        RECT 32.170 -7.290 32.500 23.150 ;
        RECT 32.810 -2.710 33.140 28.320 ;
        RECT 32.810 -7.170 33.130 -2.710 ;
        RECT 33.420 -6.560 33.750 29.800 ;
        RECT 34.040 -6.310 34.370 31.350 ;
        RECT 34.670 -5.280 35.000 32.930 ;
        RECT 35.270 -4.980 35.600 38.410 ;
        RECT 35.850 -4.410 36.180 39.970 ;
        RECT 36.460 -3.380 36.790 41.510 ;
        RECT 37.050 -2.770 37.380 43.070 ;
        RECT 37.690 -2.100 38.020 43.650 ;
        RECT 38.310 -1.450 38.640 45.250 ;
        RECT 38.910 -0.820 39.240 46.740 ;
        RECT 39.540 -0.210 39.870 48.460 ;
        RECT 40.720 47.440 41.130 47.770 ;
        RECT 40.720 45.890 41.130 46.220 ;
        RECT 41.460 44.700 41.700 49.630 ;
        RECT 44.400 49.560 44.820 50.490 ;
        RECT 47.760 49.950 48.080 50.250 ;
        RECT 48.830 49.580 49.230 50.490 ;
        RECT 42.880 48.300 43.230 48.590 ;
        RECT 42.880 48.280 43.080 48.300 ;
        RECT 42.880 46.750 43.230 47.040 ;
        RECT 42.880 46.730 43.080 46.750 ;
        RECT 42.880 45.200 43.230 45.490 ;
        RECT 42.880 45.180 43.080 45.200 ;
        RECT 44.400 44.710 44.710 49.560 ;
        RECT 44.960 49.100 45.240 49.430 ;
        RECT 47.760 48.400 48.080 48.700 ;
        RECT 44.960 47.550 45.240 47.880 ;
        RECT 47.760 46.850 48.080 47.150 ;
        RECT 44.960 46.000 45.240 46.330 ;
        RECT 47.760 45.300 48.080 45.600 ;
        RECT 40.720 44.340 41.130 44.670 ;
        RECT 41.270 44.650 41.700 44.700 ;
        RECT 44.210 44.650 44.710 44.710 ;
        RECT 41.460 44.250 41.700 44.650 ;
        RECT 44.400 44.250 44.710 44.650 ;
        RECT 44.960 44.450 45.240 44.780 ;
        RECT 48.830 44.700 49.120 49.580 ;
        RECT 48.640 44.650 49.120 44.700 ;
        RECT 48.830 44.250 49.120 44.650 ;
        RECT 44.810 43.630 44.820 43.640 ;
        RECT 41.570 43.550 41.810 43.630 ;
        RECT 44.510 43.550 44.820 43.630 ;
        RECT 48.940 43.550 49.230 43.630 ;
        RECT 50.400 43.190 50.590 56.190 ;
        RECT 52.470 43.950 52.750 44.600 ;
        RECT 52.470 43.350 52.860 43.950 ;
        RECT 40.720 42.510 41.130 42.840 ;
        RECT 41.460 42.530 41.700 42.930 ;
        RECT 44.400 42.530 44.710 42.930 ;
        RECT 41.270 42.480 41.700 42.530 ;
        RECT 40.720 40.960 41.130 41.290 ;
        RECT 40.720 39.410 41.130 39.740 ;
        RECT 40.720 37.860 41.130 38.190 ;
        RECT 41.460 37.550 41.700 42.480 ;
        RECT 44.210 42.470 44.710 42.530 ;
        RECT 42.880 41.980 43.080 42.000 ;
        RECT 42.880 41.690 43.230 41.980 ;
        RECT 42.880 40.430 43.080 40.450 ;
        RECT 42.880 40.140 43.230 40.430 ;
        RECT 42.880 38.880 43.080 38.900 ;
        RECT 42.880 38.590 43.230 38.880 ;
        RECT 44.400 37.620 44.710 42.470 ;
        RECT 44.960 42.400 45.240 42.730 ;
        RECT 48.830 42.530 49.120 42.930 ;
        RECT 48.640 42.480 49.120 42.530 ;
        RECT 47.760 41.580 48.080 41.880 ;
        RECT 44.960 40.850 45.240 41.180 ;
        RECT 47.760 40.030 48.080 40.330 ;
        RECT 44.960 39.300 45.240 39.630 ;
        RECT 47.760 38.480 48.080 38.780 ;
        RECT 44.960 37.750 45.240 38.080 ;
        RECT 41.460 36.690 41.810 37.550 ;
        RECT 42.880 37.330 43.080 37.350 ;
        RECT 42.880 37.040 43.230 37.330 ;
        RECT 44.400 36.690 44.820 37.620 ;
        RECT 48.830 37.600 49.120 42.480 ;
        RECT 52.470 39.800 52.750 43.350 ;
        RECT 53.000 43.140 53.190 44.600 ;
        RECT 54.680 44.220 54.930 57.180 ;
        RECT 56.380 57.140 57.110 64.010 ;
        RECT 74.160 62.840 77.350 63.960 ;
        RECT 66.930 58.770 68.400 59.300 ;
        RECT 56.540 46.750 56.710 57.140 ;
        RECT 64.560 56.160 65.000 56.660 ;
        RECT 58.760 52.410 59.100 52.700 ;
        RECT 58.810 52.380 59.070 52.410 ;
        RECT 56.930 48.850 57.190 49.170 ;
        RECT 56.960 46.620 57.150 48.850 ;
        RECT 58.830 46.600 59.040 52.380 ;
        RECT 62.400 51.780 62.660 51.790 ;
        RECT 62.380 51.480 62.680 51.780 ;
        RECT 62.400 51.470 62.660 51.480 ;
        RECT 59.230 50.450 59.570 50.770 ;
        RECT 59.300 46.620 59.490 50.450 ;
        RECT 59.670 48.360 59.960 48.680 ;
        RECT 59.710 46.600 59.920 48.360 ;
        RECT 60.710 47.880 61.050 48.200 ;
        RECT 60.790 46.630 60.970 47.880 ;
        RECT 54.400 43.780 54.930 44.220 ;
        RECT 54.680 43.150 54.930 43.780 ;
        RECT 59.480 43.390 59.710 44.600 ;
        RECT 60.700 43.630 60.930 44.600 ;
        RECT 52.970 43.110 53.190 43.140 ;
        RECT 52.960 42.840 53.210 43.110 ;
        RECT 52.960 42.830 53.200 42.840 ;
        RECT 52.970 42.590 53.200 42.830 ;
        RECT 54.240 42.820 54.560 43.140 ;
        RECT 59.450 42.600 59.710 43.390 ;
        RECT 60.690 43.450 60.930 43.630 ;
        RECT 60.690 43.380 61.090 43.450 ;
        RECT 60.700 43.230 61.090 43.380 ;
        RECT 61.500 43.230 61.820 43.550 ;
        RECT 62.430 43.450 62.630 51.470 ;
        RECT 64.660 46.580 64.890 56.160 ;
        RECT 65.560 52.390 65.840 52.710 ;
        RECT 65.120 51.480 65.400 51.800 ;
        RECT 60.620 42.740 61.090 43.230 ;
        RECT 61.480 43.090 61.850 43.110 ;
        RECT 61.430 42.830 61.850 43.090 ;
        RECT 61.480 42.820 61.850 42.830 ;
        RECT 53.000 40.560 53.160 42.590 ;
        RECT 53.350 42.030 53.590 42.160 ;
        RECT 53.330 41.710 53.590 42.030 ;
        RECT 53.330 41.110 53.590 41.430 ;
        RECT 53.350 40.990 53.590 41.110 ;
        RECT 56.440 40.730 56.720 40.780 ;
        RECT 52.970 40.320 53.200 40.560 ;
        RECT 56.440 40.450 56.760 40.730 ;
        RECT 56.970 40.720 57.160 40.780 ;
        RECT 59.480 40.450 59.710 42.600 ;
        RECT 60.700 42.580 61.090 42.740 ;
        RECT 60.440 42.480 61.090 42.580 ;
        RECT 60.440 42.300 61.130 42.480 ;
        RECT 60.700 42.190 61.130 42.300 ;
        RECT 60.700 41.590 61.090 42.190 ;
        RECT 60.700 41.480 61.130 41.590 ;
        RECT 60.440 41.300 61.130 41.480 ;
        RECT 60.440 41.200 61.090 41.300 ;
        RECT 60.700 41.040 61.090 41.200 ;
        RECT 60.620 40.550 61.090 41.040 ;
        RECT 62.210 41.110 62.630 43.450 ;
        RECT 61.480 40.950 61.850 40.960 ;
        RECT 61.430 40.690 61.850 40.950 ;
        RECT 61.480 40.670 61.850 40.690 ;
        RECT 62.210 40.780 62.690 41.110 ;
        RECT 52.960 40.310 53.200 40.320 ;
        RECT 52.960 40.040 53.210 40.310 ;
        RECT 54.240 40.060 54.560 40.380 ;
        RECT 52.970 40.010 53.190 40.040 ;
        RECT 52.470 39.200 52.860 39.800 ;
        RECT 52.470 38.550 52.750 39.200 ;
        RECT 53.000 38.550 53.190 40.010 ;
        RECT 59.450 39.660 59.710 40.450 ;
        RECT 60.700 40.300 61.090 40.550 ;
        RECT 60.620 39.810 61.090 40.300 ;
        RECT 61.480 40.160 61.850 40.180 ;
        RECT 61.430 39.900 61.850 40.160 ;
        RECT 61.480 39.890 61.850 39.900 ;
        RECT 54.400 38.930 54.710 39.370 ;
        RECT 59.480 38.550 59.710 39.660 ;
        RECT 60.700 39.650 61.090 39.810 ;
        RECT 60.440 39.550 61.090 39.650 ;
        RECT 60.440 39.370 61.130 39.550 ;
        RECT 61.530 39.540 61.850 39.860 ;
        RECT 60.700 39.260 61.130 39.370 ;
        RECT 60.700 38.660 61.090 39.260 ;
        RECT 60.700 38.550 61.130 38.660 ;
        RECT 60.440 38.270 60.760 38.550 ;
        RECT 60.900 38.370 61.130 38.550 ;
        RECT 60.900 38.110 61.090 38.370 ;
        RECT 60.620 37.620 61.090 38.110 ;
        RECT 61.480 38.020 61.850 38.030 ;
        RECT 61.430 37.760 61.850 38.020 ;
        RECT 61.480 37.740 61.850 37.760 ;
        RECT 47.760 36.930 48.080 37.230 ;
        RECT 48.830 36.690 49.230 37.600 ;
        RECT 41.270 36.290 41.510 36.340 ;
        RECT 41.570 33.180 41.810 36.690 ;
        RECT 44.510 36.360 44.820 36.690 ;
        RECT 44.210 36.290 44.820 36.360 ;
        RECT 48.640 36.290 48.930 36.340 ;
        RECT 44.510 33.110 44.820 36.290 ;
        RECT 48.940 33.130 49.230 36.690 ;
        RECT 50.400 33.140 50.590 37.540 ;
        RECT 51.710 33.330 51.940 37.580 ;
        RECT 54.680 33.330 54.930 37.600 ;
        RECT 60.900 37.400 61.090 37.620 ;
        RECT 62.210 37.400 62.440 40.780 ;
        RECT 62.990 38.560 63.410 44.600 ;
        RECT 65.150 43.450 65.370 51.480 ;
        RECT 65.150 43.230 65.430 43.450 ;
        RECT 65.580 43.230 65.810 52.390 ;
        RECT 66.950 46.390 67.370 58.770 ;
        RECT 67.980 46.390 68.400 58.770 ;
        RECT 70.360 56.120 70.800 56.620 ;
        RECT 70.460 49.140 70.690 56.120 ;
        RECT 74.880 50.870 76.160 62.840 ;
        RECT 78.640 57.650 78.920 57.770 ;
        RECT 78.640 57.150 78.970 57.650 ;
        RECT 74.880 50.790 76.180 50.870 ;
        RECT 74.870 50.490 76.180 50.790 ;
        RECT 71.650 49.840 71.950 50.160 ;
        RECT 70.330 49.130 70.690 49.140 ;
        RECT 70.300 48.280 70.690 49.130 ;
        RECT 70.330 48.270 70.690 48.280 ;
        RECT 70.460 46.580 70.690 48.270 ;
        RECT 71.680 46.580 71.910 49.840 ;
        RECT 77.960 49.290 78.390 49.630 ;
        RECT 78.200 46.620 78.390 49.290 ;
        RECT 78.640 46.530 78.920 57.150 ;
        RECT 80.340 52.390 80.600 52.710 ;
        RECT 79.450 51.520 79.710 51.840 ;
        RECT 79.480 47.800 79.670 51.520 ;
        RECT 80.360 47.800 80.580 52.390 ;
        RECT 82.330 49.170 82.670 65.390 ;
        RECT 86.830 61.930 87.200 61.940 ;
        RECT 86.780 61.480 87.280 61.930 ;
        RECT 82.980 53.070 83.300 53.440 ;
        RECT 83.000 49.230 83.270 53.070 ;
        RECT 82.280 49.090 82.670 49.170 ;
        RECT 82.270 48.320 82.670 49.090 ;
        RECT 82.280 48.250 82.670 48.320 ;
        RECT 79.310 47.110 79.990 47.800 ;
        RECT 80.350 47.110 81.030 47.800 ;
        RECT 82.330 46.470 82.670 48.250 ;
        RECT 82.720 48.580 82.880 49.230 ;
        RECT 82.720 48.030 82.990 48.580 ;
        RECT 82.710 47.980 82.990 48.030 ;
        RECT 82.710 47.890 82.880 47.980 ;
        RECT 82.720 44.600 82.880 47.890 ;
        RECT 83.000 47.740 83.320 49.230 ;
        RECT 85.000 48.860 85.210 49.230 ;
        RECT 84.530 48.410 84.840 48.850 ;
        RECT 84.990 48.570 85.220 48.860 ;
        RECT 83.000 47.690 83.340 47.740 ;
        RECT 83.000 47.190 83.680 47.690 ;
        RECT 83.000 46.540 83.290 47.190 ;
        RECT 84.130 46.880 84.450 47.200 ;
        RECT 85.000 46.870 85.210 48.570 ;
        RECT 85.470 48.300 85.660 49.230 ;
        RECT 85.460 48.010 85.690 48.300 ;
        RECT 83.130 45.190 83.290 46.540 ;
        RECT 83.480 46.370 83.720 46.790 ;
        RECT 84.990 46.580 85.220 46.870 ;
        RECT 85.000 46.440 85.210 46.580 ;
        RECT 83.450 46.050 83.720 46.370 ;
        RECT 83.480 45.620 83.720 46.050 ;
        RECT 85.470 45.980 85.660 48.010 ;
        RECT 85.880 46.510 86.090 49.230 ;
        RECT 85.850 46.000 86.090 46.510 ;
        RECT 85.020 45.800 85.210 45.930 ;
        RECT 85.000 45.510 85.230 45.800 ;
        RECT 85.460 45.690 85.690 45.980 ;
        RECT 84.120 45.190 84.440 45.510 ;
        RECT 83.100 44.950 83.330 45.190 ;
        RECT 83.090 44.940 83.330 44.950 ;
        RECT 83.090 44.670 83.340 44.940 ;
        RECT 83.100 44.640 83.320 44.670 ;
        RECT 63.940 43.070 64.280 43.120 ;
        RECT 63.940 43.050 64.500 43.070 ;
        RECT 63.820 42.880 64.500 43.050 ;
        RECT 63.940 42.840 64.500 42.880 ;
        RECT 63.940 42.800 64.280 42.840 ;
        RECT 65.150 42.160 65.820 43.230 ;
        RECT 65.150 41.620 65.430 42.160 ;
        RECT 65.580 41.620 65.810 42.160 ;
        RECT 63.940 40.940 64.280 40.980 ;
        RECT 63.940 40.900 64.500 40.940 ;
        RECT 63.450 40.690 63.680 40.770 ;
        RECT 63.820 40.730 64.500 40.900 ;
        RECT 63.940 40.710 64.500 40.730 ;
        RECT 63.940 40.660 64.280 40.710 ;
        RECT 64.670 40.690 64.900 40.770 ;
        RECT 65.150 40.550 65.820 41.620 ;
        RECT 66.960 40.620 68.400 40.780 ;
        RECT 70.460 40.690 70.690 40.780 ;
        RECT 71.680 40.700 71.910 40.780 ;
        RECT 65.150 40.300 65.430 40.550 ;
        RECT 65.580 40.300 65.810 40.550 ;
        RECT 63.940 40.140 64.280 40.190 ;
        RECT 63.940 40.120 64.500 40.140 ;
        RECT 63.820 39.950 64.500 40.120 ;
        RECT 63.940 39.910 64.500 39.950 ;
        RECT 65.150 39.940 65.820 40.300 ;
        RECT 63.940 39.870 64.280 39.910 ;
        RECT 65.140 39.870 65.820 39.940 ;
        RECT 65.130 39.270 65.820 39.870 ;
        RECT 65.140 39.240 65.820 39.270 ;
        RECT 65.150 39.230 65.820 39.240 ;
        RECT 65.150 38.690 65.430 39.230 ;
        RECT 63.940 38.010 64.280 38.050 ;
        RECT 63.940 37.970 64.500 38.010 ;
        RECT 63.820 37.800 64.500 37.970 ;
        RECT 64.700 37.960 64.870 38.130 ;
        RECT 63.940 37.780 64.500 37.800 ;
        RECT 63.940 37.730 64.280 37.780 ;
        RECT 64.680 37.370 65.000 37.670 ;
        RECT 65.150 37.620 65.820 38.690 ;
        RECT 71.940 38.550 72.360 44.600 ;
        RECT 74.420 38.550 74.650 44.600 ;
        RECT 75.640 43.390 75.870 44.600 ;
        RECT 80.640 43.780 80.950 44.220 ;
        RECT 75.640 42.600 75.900 43.390 ;
        RECT 82.160 43.140 82.350 44.600 ;
        RECT 82.600 44.430 82.880 44.600 ;
        RECT 82.600 43.950 82.990 44.430 ;
        RECT 82.490 43.830 82.990 43.950 ;
        RECT 82.490 43.350 82.880 43.830 ;
        RECT 80.790 42.820 81.110 43.140 ;
        RECT 82.160 43.110 82.380 43.140 ;
        RECT 82.140 42.840 82.390 43.110 ;
        RECT 82.150 42.830 82.390 42.840 ;
        RECT 75.640 40.450 75.870 42.600 ;
        RECT 82.150 42.590 82.380 42.830 ;
        RECT 81.760 42.030 82.000 42.160 ;
        RECT 81.760 41.710 82.020 42.030 ;
        RECT 81.760 41.110 82.020 41.430 ;
        RECT 81.760 40.990 82.000 41.110 ;
        RECT 82.190 40.780 82.350 42.590 ;
        RECT 82.600 41.750 82.880 43.350 ;
        RECT 83.130 43.180 83.320 44.640 ;
        RECT 84.530 43.560 84.840 44.000 ;
        RECT 85.020 43.890 85.210 45.510 ;
        RECT 85.470 44.400 85.660 45.690 ;
        RECT 85.450 44.110 85.680 44.400 ;
        RECT 85.020 43.680 85.250 43.890 ;
        RECT 85.010 43.600 85.250 43.680 ;
        RECT 85.010 43.180 85.240 43.600 ;
        RECT 85.470 43.180 85.660 44.110 ;
        RECT 85.880 43.180 86.090 46.000 ;
        RECT 86.830 45.410 87.200 61.480 ;
        RECT 87.620 58.030 88.080 58.460 ;
        RECT 86.670 45.390 87.270 45.410 ;
        RECT 86.510 45.350 87.270 45.390 ;
        RECT 86.510 45.090 87.200 45.350 ;
        RECT 82.600 41.430 82.960 41.750 ;
        RECT 82.600 40.780 82.880 41.430 ;
        RECT 78.200 40.700 78.390 40.780 ;
        RECT 78.640 40.730 78.920 40.780 ;
        RECT 75.640 39.660 75.900 40.450 ;
        RECT 78.640 40.430 78.960 40.730 ;
        RECT 80.390 40.440 80.710 40.760 ;
        RECT 82.190 40.560 82.880 40.780 ;
        RECT 82.990 40.630 83.270 40.780 ;
        RECT 80.790 40.060 81.110 40.380 ;
        RECT 81.370 40.160 81.690 40.480 ;
        RECT 82.150 40.310 82.880 40.560 ;
        RECT 82.140 40.040 82.880 40.310 ;
        RECT 75.640 38.550 75.870 39.660 ;
        RECT 80.540 39.610 80.860 39.930 ;
        RECT 81.320 39.510 81.640 39.830 ;
        RECT 79.430 39.080 79.750 39.400 ;
        RECT 80.640 38.930 80.950 39.370 ;
        RECT 80.650 38.920 80.860 38.930 ;
        RECT 80.630 38.600 80.890 38.920 ;
        RECT 81.320 38.680 81.640 39.000 ;
        RECT 70.490 37.960 70.660 38.130 ;
        RECT 80.160 37.800 80.480 38.120 ;
        RECT 65.150 37.400 65.430 37.620 ;
        RECT 64.710 37.270 64.880 37.370 ;
        RECT 65.150 36.040 65.370 37.400 ;
        RECT 70.380 37.300 70.700 37.620 ;
        RECT 80.650 37.310 80.860 38.600 ;
        RECT 82.160 38.550 82.880 40.040 ;
        RECT 83.000 39.200 83.270 40.630 ;
        RECT 83.620 40.210 83.940 40.530 ;
        RECT 83.000 38.910 83.280 39.200 ;
        RECT 81.370 38.030 81.690 38.350 ;
        RECT 68.040 36.640 68.200 37.290 ;
        RECT 68.040 36.090 68.310 36.640 ;
        RECT 68.030 36.040 68.310 36.090 ;
        RECT 68.450 36.300 68.640 37.290 ;
        RECT 68.850 36.610 69.010 37.290 ;
        RECT 70.490 37.280 70.660 37.300 ;
        RECT 68.810 36.590 69.010 36.610 ;
        RECT 69.830 36.600 70.150 36.920 ;
        RECT 68.800 36.350 69.030 36.590 ;
        RECT 68.450 36.180 68.620 36.300 ;
        RECT 65.150 35.950 65.500 36.040 ;
        RECT 68.030 35.950 68.200 36.040 ;
        RECT 65.150 35.730 65.660 35.950 ;
        RECT 68.040 35.590 68.200 35.950 ;
        RECT 68.030 35.500 68.200 35.590 ;
        RECT 68.030 35.450 68.310 35.500 ;
        RECT 68.040 35.150 68.310 35.450 ;
        RECT 68.450 35.360 68.610 36.180 ;
        RECT 68.810 36.130 69.010 36.350 ;
        RECT 68.850 35.410 69.010 36.130 ;
        RECT 69.830 36.050 70.150 36.370 ;
        RECT 70.790 36.130 71.030 37.290 ;
        RECT 68.450 35.240 68.620 35.360 ;
        RECT 56.440 33.900 56.720 35.010 ;
        RECT 56.970 34.320 57.160 34.920 ;
        RECT 58.970 34.480 59.360 34.500 ;
        RECT 58.960 34.390 59.360 34.480 ;
        RECT 56.970 34.130 58.600 34.320 ;
        RECT 56.440 33.620 58.160 33.900 ;
        RECT 57.880 33.390 58.160 33.620 ;
        RECT 58.410 33.350 58.600 34.130 ;
        RECT 58.810 34.140 59.360 34.390 ;
        RECT 58.810 34.120 59.350 34.140 ;
        RECT 58.810 33.270 58.970 34.120 ;
        RECT 62.930 34.050 63.310 34.070 ;
        RECT 63.450 34.050 63.680 34.960 ;
        RECT 62.930 33.820 63.680 34.050 ;
        RECT 64.670 33.960 64.900 34.960 ;
        RECT 67.980 33.970 68.400 35.150 ;
        RECT 68.450 34.380 68.640 35.240 ;
        RECT 68.810 35.190 69.010 35.410 ;
        RECT 68.800 34.950 69.030 35.190 ;
        RECT 69.830 35.170 70.150 35.490 ;
        RECT 70.780 35.470 71.050 36.130 ;
        RECT 68.810 34.930 69.010 34.950 ;
        RECT 68.420 34.150 68.660 34.380 ;
        RECT 60.900 33.160 61.090 33.380 ;
        RECT 40.720 32.380 41.130 32.710 ;
        RECT 41.460 32.400 41.700 32.800 ;
        RECT 44.400 32.400 44.710 32.800 ;
        RECT 41.270 32.350 41.700 32.400 ;
        RECT 40.720 30.830 41.130 31.160 ;
        RECT 40.720 29.280 41.130 29.610 ;
        RECT 40.720 27.730 41.130 28.060 ;
        RECT 41.460 27.420 41.700 32.350 ;
        RECT 44.210 32.340 44.710 32.400 ;
        RECT 42.880 31.850 43.080 31.870 ;
        RECT 42.880 31.560 43.230 31.850 ;
        RECT 42.880 30.300 43.080 30.320 ;
        RECT 42.880 30.010 43.230 30.300 ;
        RECT 42.880 28.750 43.080 28.770 ;
        RECT 42.880 28.460 43.230 28.750 ;
        RECT 44.400 27.490 44.710 32.340 ;
        RECT 44.960 32.270 45.240 32.600 ;
        RECT 48.830 32.400 49.120 32.800 ;
        RECT 60.620 32.670 61.090 33.160 ;
        RECT 61.480 33.020 61.850 33.040 ;
        RECT 61.430 32.760 61.850 33.020 ;
        RECT 61.480 32.750 61.850 32.760 ;
        RECT 48.640 32.350 49.120 32.400 ;
        RECT 47.760 31.450 48.080 31.750 ;
        RECT 44.960 30.720 45.240 31.050 ;
        RECT 47.760 29.900 48.080 30.200 ;
        RECT 44.960 29.170 45.240 29.500 ;
        RECT 47.760 28.350 48.080 28.650 ;
        RECT 44.960 27.620 45.240 27.950 ;
        RECT 41.460 26.560 41.810 27.420 ;
        RECT 42.880 27.200 43.080 27.220 ;
        RECT 42.880 26.910 43.230 27.200 ;
        RECT 44.400 26.560 44.820 27.490 ;
        RECT 48.830 27.470 49.120 32.350 ;
        RECT 60.440 32.230 60.760 32.510 ;
        RECT 60.900 32.410 61.090 32.670 ;
        RECT 60.900 32.120 61.130 32.410 ;
        RECT 60.900 31.520 61.090 32.120 ;
        RECT 60.440 31.130 60.760 31.410 ;
        RECT 60.900 31.230 61.130 31.520 ;
        RECT 60.900 30.970 61.090 31.230 ;
        RECT 60.620 30.480 61.090 30.970 ;
        RECT 61.480 30.880 61.850 30.890 ;
        RECT 61.430 30.620 61.850 30.880 ;
        RECT 61.480 30.600 61.850 30.620 ;
        RECT 60.900 30.230 61.090 30.480 ;
        RECT 60.620 29.740 61.090 30.230 ;
        RECT 61.480 30.090 61.850 30.110 ;
        RECT 61.430 29.830 61.850 30.090 ;
        RECT 61.480 29.820 61.850 29.830 ;
        RECT 60.440 29.300 60.760 29.580 ;
        RECT 60.900 29.480 61.090 29.740 ;
        RECT 60.900 29.190 61.130 29.480 ;
        RECT 60.900 28.590 61.090 29.190 ;
        RECT 60.440 28.200 60.760 28.480 ;
        RECT 60.900 28.300 61.130 28.590 ;
        RECT 60.900 28.040 61.090 28.300 ;
        RECT 60.620 27.550 61.090 28.040 ;
        RECT 61.480 27.950 61.850 27.960 ;
        RECT 61.430 27.690 61.850 27.950 ;
        RECT 61.480 27.670 61.850 27.690 ;
        RECT 47.760 26.800 48.080 27.100 ;
        RECT 48.830 26.560 49.230 27.470 ;
        RECT 41.270 26.160 41.510 26.210 ;
        RECT 41.570 23.650 41.810 26.560 ;
        RECT 44.510 26.230 44.820 26.560 ;
        RECT 44.210 26.160 44.820 26.230 ;
        RECT 48.640 26.160 48.930 26.210 ;
        RECT 44.510 23.650 44.820 26.160 ;
        RECT 48.940 23.650 49.230 26.560 ;
        RECT 50.400 23.380 50.590 27.470 ;
        RECT 51.710 26.430 51.940 27.510 ;
        RECT 51.620 25.950 51.950 26.430 ;
        RECT 51.710 23.340 51.940 25.950 ;
        RECT 54.680 23.550 54.930 27.530 ;
        RECT 55.340 26.820 55.500 27.470 ;
        RECT 55.340 26.270 55.610 26.820 ;
        RECT 55.330 26.220 55.610 26.270 ;
        RECT 55.750 26.480 55.940 27.470 ;
        RECT 56.150 26.790 56.310 27.470 ;
        RECT 56.110 26.770 56.310 26.790 ;
        RECT 57.130 26.780 57.450 27.100 ;
        RECT 56.100 26.530 56.330 26.770 ;
        RECT 55.750 26.360 55.920 26.480 ;
        RECT 55.330 26.130 55.500 26.220 ;
        RECT 55.340 25.770 55.500 26.130 ;
        RECT 55.330 25.680 55.500 25.770 ;
        RECT 55.330 25.630 55.610 25.680 ;
        RECT 55.340 25.080 55.610 25.630 ;
        RECT 55.750 25.540 55.910 26.360 ;
        RECT 56.110 26.310 56.310 26.530 ;
        RECT 56.150 25.590 56.310 26.310 ;
        RECT 57.130 26.230 57.450 26.550 ;
        RECT 55.750 25.420 55.920 25.540 ;
        RECT 55.340 23.810 55.500 25.080 ;
        RECT 55.750 24.560 55.940 25.420 ;
        RECT 56.110 25.370 56.310 25.590 ;
        RECT 56.100 25.130 56.330 25.370 ;
        RECT 57.130 25.350 57.450 25.670 ;
        RECT 56.110 25.110 56.310 25.130 ;
        RECT 55.720 24.330 55.960 24.560 ;
        RECT 55.340 23.260 55.610 23.810 ;
        RECT 55.330 23.210 55.610 23.260 ;
        RECT 55.750 23.470 55.940 24.330 ;
        RECT 56.150 23.780 56.310 25.110 ;
        RECT 57.130 24.800 57.450 25.120 ;
        RECT 56.110 23.760 56.310 23.780 ;
        RECT 57.130 23.770 57.450 24.090 ;
        RECT 56.100 23.520 56.330 23.760 ;
        RECT 55.750 23.350 55.920 23.470 ;
        RECT 55.330 23.120 55.500 23.210 ;
        RECT 40.720 22.610 41.130 22.940 ;
        RECT 41.460 22.630 41.700 23.030 ;
        RECT 44.400 22.630 44.710 23.030 ;
        RECT 41.270 22.580 41.700 22.630 ;
        RECT 40.720 21.060 41.130 21.390 ;
        RECT 40.720 19.510 41.130 19.840 ;
        RECT 40.720 17.960 41.130 18.290 ;
        RECT 41.460 17.650 41.700 22.580 ;
        RECT 44.210 22.570 44.710 22.630 ;
        RECT 42.880 22.080 43.080 22.100 ;
        RECT 42.880 21.790 43.230 22.080 ;
        RECT 42.880 20.530 43.080 20.550 ;
        RECT 42.880 20.240 43.230 20.530 ;
        RECT 42.880 18.980 43.080 19.000 ;
        RECT 42.880 18.690 43.230 18.980 ;
        RECT 44.400 17.720 44.710 22.570 ;
        RECT 44.960 22.500 45.240 22.830 ;
        RECT 48.830 22.630 49.120 23.030 ;
        RECT 55.340 22.770 55.500 23.120 ;
        RECT 55.330 22.680 55.500 22.770 ;
        RECT 55.330 22.630 55.610 22.680 ;
        RECT 48.640 22.580 49.120 22.630 ;
        RECT 47.760 21.680 48.080 21.980 ;
        RECT 44.960 20.950 45.240 21.280 ;
        RECT 47.760 20.130 48.080 20.430 ;
        RECT 44.960 19.400 45.240 19.730 ;
        RECT 47.760 18.580 48.080 18.880 ;
        RECT 44.960 17.850 45.240 18.180 ;
        RECT 41.460 16.790 41.810 17.650 ;
        RECT 42.880 17.430 43.080 17.450 ;
        RECT 42.880 17.140 43.230 17.430 ;
        RECT 44.400 16.790 44.820 17.720 ;
        RECT 48.830 17.700 49.120 22.580 ;
        RECT 55.340 22.080 55.610 22.630 ;
        RECT 55.750 22.540 55.910 23.350 ;
        RECT 56.110 23.300 56.310 23.520 ;
        RECT 56.150 22.590 56.310 23.300 ;
        RECT 57.130 23.220 57.450 23.540 ;
        RECT 58.000 23.490 58.160 27.540 ;
        RECT 58.210 23.650 58.460 27.470 ;
        RECT 60.270 25.550 60.650 27.470 ;
        RECT 60.750 27.330 61.090 27.550 ;
        RECT 62.210 27.470 62.440 33.380 ;
        RECT 62.930 33.050 63.310 33.820 ;
        RECT 64.670 33.660 64.920 33.960 ;
        RECT 64.680 33.190 64.920 33.660 ;
        RECT 67.980 33.580 68.440 33.970 ;
        RECT 65.180 33.160 65.430 33.380 ;
        RECT 63.940 33.000 64.280 33.050 ;
        RECT 63.940 32.980 64.500 33.000 ;
        RECT 63.820 32.810 64.500 32.980 ;
        RECT 63.940 32.770 64.500 32.810 ;
        RECT 63.940 32.730 64.280 32.770 ;
        RECT 65.180 32.090 65.820 33.160 ;
        RECT 68.040 33.080 68.440 33.580 ;
        RECT 68.030 33.030 68.440 33.080 ;
        RECT 68.450 33.290 68.640 34.150 ;
        RECT 68.850 33.600 69.010 34.930 ;
        RECT 69.830 34.620 70.150 34.940 ;
        RECT 70.380 34.790 70.700 35.090 ;
        RECT 70.460 33.980 70.690 34.790 ;
        RECT 68.810 33.580 69.010 33.600 ;
        RECT 69.830 33.590 70.150 33.910 ;
        RECT 70.460 33.630 70.720 33.980 ;
        RECT 68.800 33.340 69.030 33.580 ;
        RECT 70.480 33.470 70.720 33.630 ;
        RECT 70.790 33.470 71.030 35.470 ;
        RECT 72.970 35.370 73.350 37.290 ;
        RECT 74.720 36.110 74.960 37.290 ;
        RECT 74.710 35.450 74.970 36.110 ;
        RECT 71.680 34.070 71.910 34.960 ;
        RECT 71.660 33.690 72.470 34.070 ;
        RECT 68.450 33.170 68.620 33.290 ;
        RECT 68.030 32.940 68.200 33.030 ;
        RECT 68.040 32.590 68.200 32.940 ;
        RECT 68.030 32.500 68.200 32.590 ;
        RECT 68.030 32.450 68.310 32.500 ;
        RECT 65.180 31.550 65.430 32.090 ;
        RECT 68.040 31.900 68.310 32.450 ;
        RECT 68.450 32.360 68.610 33.170 ;
        RECT 68.810 33.120 69.010 33.340 ;
        RECT 68.850 32.410 69.010 33.120 ;
        RECT 69.830 33.040 70.150 33.360 ;
        RECT 70.480 33.190 71.030 33.470 ;
        RECT 71.090 33.420 71.280 33.470 ;
        RECT 71.490 33.420 71.650 33.470 ;
        RECT 70.520 33.130 71.030 33.190 ;
        RECT 70.790 32.880 71.030 33.130 ;
        RECT 72.090 33.050 72.470 33.690 ;
        RECT 72.970 33.510 73.360 35.370 ;
        RECT 70.780 32.560 71.040 32.880 ;
        RECT 68.450 32.240 68.620 32.360 ;
        RECT 63.940 30.870 64.280 30.910 ;
        RECT 63.940 30.830 64.500 30.870 ;
        RECT 63.820 30.660 64.500 30.830 ;
        RECT 63.940 30.640 64.500 30.660 ;
        RECT 63.940 30.590 64.280 30.640 ;
        RECT 65.180 30.480 65.820 31.550 ;
        RECT 68.040 31.250 68.200 31.900 ;
        RECT 68.450 31.250 68.640 32.240 ;
        RECT 68.810 32.190 69.010 32.410 ;
        RECT 68.800 31.950 69.030 32.190 ;
        RECT 69.830 32.170 70.150 32.490 ;
        RECT 68.810 31.930 69.010 31.950 ;
        RECT 68.850 31.250 69.010 31.930 ;
        RECT 69.830 31.620 70.150 31.940 ;
        RECT 70.790 31.240 71.030 32.560 ;
        RECT 72.970 31.240 73.350 33.510 ;
        RECT 73.430 33.380 73.670 33.470 ;
        RECT 74.720 32.840 74.960 35.450 ;
        RECT 77.000 33.940 77.400 37.290 ;
        RECT 80.630 37.020 80.860 37.310 ;
        RECT 81.370 37.200 81.690 37.520 ;
        RECT 81.320 36.550 81.640 36.870 ;
        RECT 81.320 35.720 81.640 36.040 ;
        RECT 78.200 33.940 78.390 34.920 ;
        RECT 76.370 33.570 76.650 33.890 ;
        RECT 76.800 33.750 78.390 33.940 ;
        RECT 75.610 33.370 75.990 33.470 ;
        RECT 76.430 33.270 76.590 33.570 ;
        RECT 76.800 33.400 76.990 33.750 ;
        RECT 77.000 33.560 77.400 33.750 ;
        RECT 78.640 33.560 78.920 35.010 ;
        RECT 80.820 34.930 81.150 35.220 ;
        RECT 81.370 35.070 81.690 35.390 ;
        RECT 82.330 34.930 82.670 38.550 ;
        RECT 80.810 34.790 82.670 34.930 ;
        RECT 82.330 34.730 82.670 34.790 ;
        RECT 83.000 36.610 83.270 38.910 ;
        RECT 83.670 37.990 83.990 38.310 ;
        RECT 83.660 37.290 83.980 37.590 ;
        RECT 83.360 37.270 83.980 37.290 ;
        RECT 83.000 36.320 83.280 36.610 ;
        RECT 83.000 34.730 83.270 36.320 ;
        RECT 83.360 35.340 83.760 37.270 ;
        RECT 85.800 36.110 86.040 37.290 ;
        RECT 85.790 35.450 86.050 36.110 ;
        RECT 83.360 35.020 83.900 35.340 ;
        RECT 77.000 33.280 78.920 33.560 ;
        RECT 83.360 33.470 83.760 35.020 ;
        RECT 79.640 33.340 80.040 33.470 ;
        RECT 80.720 33.370 81.120 33.470 ;
        RECT 83.160 33.420 83.760 33.470 ;
        RECT 74.710 32.520 74.970 32.840 ;
        RECT 74.720 31.240 74.960 32.520 ;
        RECT 77.000 31.240 77.400 33.280 ;
        RECT 80.040 33.110 80.720 33.330 ;
        RECT 83.360 31.240 83.760 33.420 ;
        RECT 84.770 33.370 85.150 33.470 ;
        RECT 85.800 32.840 86.040 35.450 ;
        RECT 86.830 34.570 87.200 45.090 ;
        RECT 87.640 37.290 88.010 58.030 ;
        RECT 88.390 53.320 88.840 53.750 ;
        RECT 87.410 35.370 88.010 37.290 ;
        RECT 86.800 34.110 87.250 34.570 ;
        RECT 86.830 34.070 87.200 34.110 ;
        RECT 87.400 33.980 88.010 35.370 ;
        RECT 87.400 33.520 88.050 33.980 ;
        RECT 87.400 33.510 88.010 33.520 ;
        RECT 87.410 33.470 88.010 33.510 ;
        RECT 87.090 33.400 87.330 33.470 ;
        RECT 85.790 32.520 86.050 32.840 ;
        RECT 85.800 31.240 86.040 32.520 ;
        RECT 87.410 31.240 87.790 33.470 ;
        RECT 88.410 31.630 88.780 53.320 ;
        RECT 94.960 52.270 95.540 52.830 ;
        RECT 91.750 50.700 92.310 51.350 ;
        RECT 92.700 51.190 93.260 51.770 ;
        RECT 93.780 51.650 94.340 52.240 ;
        RECT 89.280 48.240 89.710 48.680 ;
        RECT 88.950 45.300 89.160 45.410 ;
        RECT 88.960 39.370 89.190 39.490 ;
        RECT 89.290 33.470 89.660 48.240 ;
        RECT 90.830 45.410 91.060 49.230 ;
        RECT 89.830 45.350 90.040 45.410 ;
        RECT 90.830 45.340 91.090 45.410 ;
        RECT 90.830 43.180 91.060 45.340 ;
        RECT 91.770 37.290 92.270 50.700 ;
        RECT 92.700 49.230 93.200 51.190 ;
        RECT 92.700 43.180 93.540 49.230 ;
        RECT 92.700 37.290 93.200 43.180 ;
        RECT 89.730 36.130 89.970 37.290 ;
        RECT 90.610 36.600 90.930 36.920 ;
        RECT 91.750 36.590 92.310 37.290 ;
        RECT 92.560 36.640 93.200 37.290 ;
        RECT 89.710 35.470 89.980 36.130 ;
        RECT 90.610 36.050 90.930 36.370 ;
        RECT 91.730 36.350 92.310 36.590 ;
        RECT 89.730 33.470 89.970 35.470 ;
        RECT 90.610 35.170 90.930 35.490 ;
        RECT 91.750 35.190 92.310 36.350 ;
        RECT 92.450 36.040 93.200 36.640 ;
        RECT 92.560 35.500 93.200 36.040 ;
        RECT 91.730 34.950 92.310 35.190 ;
        RECT 90.610 34.620 90.930 34.940 ;
        RECT 91.750 34.380 92.310 34.950 ;
        RECT 92.450 34.900 93.200 35.500 ;
        RECT 91.750 34.150 92.340 34.380 ;
        RECT 90.610 33.590 90.930 33.910 ;
        RECT 91.750 33.580 92.310 34.150 ;
        RECT 92.560 33.630 93.200 34.900 ;
        RECT 89.110 33.420 89.270 33.470 ;
        RECT 89.290 33.420 89.670 33.470 ;
        RECT 89.730 33.430 90.080 33.470 ;
        RECT 88.380 31.620 88.780 31.630 ;
        RECT 88.370 31.200 88.790 31.620 ;
        RECT 88.410 31.190 88.780 31.200 ;
        RECT 65.180 30.230 65.430 30.480 ;
        RECT 63.940 30.070 64.280 30.120 ;
        RECT 63.940 30.050 64.500 30.070 ;
        RECT 63.820 29.880 64.500 30.050 ;
        RECT 63.940 29.840 64.500 29.880 ;
        RECT 63.940 29.800 64.280 29.840 ;
        RECT 65.180 29.160 65.820 30.230 ;
        RECT 65.180 28.620 65.430 29.160 ;
        RECT 63.940 27.940 64.280 27.980 ;
        RECT 63.940 27.900 64.500 27.940 ;
        RECT 62.210 27.330 62.490 27.470 ;
        RECT 60.270 23.690 60.660 25.550 ;
        RECT 60.750 23.900 60.990 27.330 ;
        RECT 58.210 23.580 58.600 23.650 ;
        RECT 58.810 23.580 58.970 23.650 ;
        RECT 58.210 23.030 58.460 23.580 ;
        RECT 60.270 23.400 60.650 23.690 ;
        RECT 60.730 23.650 61.120 23.900 ;
        RECT 60.870 23.400 61.120 23.650 ;
        RECT 62.220 23.620 62.490 27.330 ;
        RECT 58.190 23.000 58.470 23.030 ;
        RECT 58.180 22.720 58.480 23.000 ;
        RECT 60.270 22.910 61.090 23.400 ;
        RECT 61.480 23.260 61.850 23.280 ;
        RECT 61.430 23.000 61.850 23.260 ;
        RECT 62.210 23.000 62.490 23.620 ;
        RECT 62.930 23.270 63.310 27.760 ;
        RECT 63.820 27.730 64.500 27.900 ;
        RECT 63.940 27.710 64.500 27.730 ;
        RECT 63.940 27.660 64.280 27.710 ;
        RECT 64.680 27.470 64.920 27.620 ;
        RECT 64.300 23.880 64.920 27.470 ;
        RECT 65.180 27.550 65.820 28.620 ;
        RECT 65.180 27.330 65.430 27.550 ;
        RECT 64.300 23.610 65.150 23.880 ;
        RECT 63.940 23.240 64.280 23.290 ;
        RECT 64.300 23.240 64.700 23.610 ;
        RECT 64.880 23.380 65.150 23.610 ;
        RECT 65.180 23.400 65.430 23.620 ;
        RECT 63.940 23.220 64.700 23.240 ;
        RECT 63.820 23.050 64.700 23.220 ;
        RECT 63.940 23.010 64.700 23.050 ;
        RECT 61.480 22.990 61.850 23.000 ;
        RECT 60.270 22.750 60.650 22.910 ;
        RECT 58.190 22.700 58.470 22.720 ;
        RECT 56.110 22.560 56.310 22.590 ;
        RECT 55.750 22.420 55.920 22.540 ;
        RECT 55.340 21.430 55.500 22.080 ;
        RECT 55.750 21.430 55.940 22.420 ;
        RECT 56.030 22.220 56.350 22.560 ;
        RECT 57.130 22.350 57.450 22.670 ;
        RECT 56.100 22.130 56.330 22.220 ;
        RECT 47.760 17.030 48.080 17.330 ;
        RECT 48.830 17.080 49.230 17.700 ;
        RECT 49.440 17.100 49.780 17.420 ;
        RECT 48.830 16.790 49.260 17.080 ;
        RECT 41.270 16.390 41.510 16.440 ;
        RECT 41.570 5.020 41.810 16.790 ;
        RECT 44.510 16.570 44.820 16.790 ;
        RECT 48.910 16.730 49.260 16.790 ;
        RECT 44.470 16.460 44.840 16.570 ;
        RECT 44.210 16.390 44.840 16.460 ;
        RECT 48.640 16.390 48.930 16.440 ;
        RECT 44.470 16.240 44.840 16.390 ;
        RECT 48.940 16.270 49.230 16.730 ;
        RECT 49.440 16.490 49.690 17.100 ;
        RECT 50.400 16.510 50.590 17.710 ;
        RECT 54.680 17.040 54.930 17.770 ;
        RECT 56.110 17.460 56.320 22.130 ;
        RECT 57.130 21.800 57.450 22.120 ;
        RECT 57.140 21.720 57.400 21.800 ;
        RECT 57.130 21.520 57.400 21.720 ;
        RECT 57.130 20.830 57.340 21.520 ;
        RECT 58.210 21.420 58.460 22.700 ;
        RECT 60.270 22.470 60.760 22.750 ;
        RECT 60.900 22.650 61.090 22.910 ;
        RECT 62.200 22.690 62.510 23.000 ;
        RECT 63.940 22.970 64.280 23.010 ;
        RECT 60.270 22.340 60.650 22.470 ;
        RECT 60.900 22.360 61.130 22.650 ;
        RECT 60.270 22.020 60.670 22.340 ;
        RECT 60.270 21.650 60.650 22.020 ;
        RECT 60.900 21.760 61.090 22.360 ;
        RECT 60.270 21.420 60.760 21.650 ;
        RECT 60.440 21.370 60.760 21.420 ;
        RECT 60.900 21.470 61.130 21.760 ;
        RECT 60.900 21.210 61.090 21.470 ;
        RECT 57.120 20.780 57.380 20.830 ;
        RECT 57.120 20.530 57.760 20.780 ;
        RECT 60.620 20.720 61.090 21.210 ;
        RECT 62.210 21.420 62.490 22.690 ;
        RECT 64.300 21.420 64.700 23.010 ;
        RECT 65.180 22.330 65.820 23.400 ;
        RECT 66.960 23.250 67.360 27.780 ;
        RECT 70.480 27.480 70.720 27.620 ;
        RECT 70.480 27.420 70.840 27.480 ;
        RECT 71.090 27.430 71.280 27.490 ;
        RECT 71.490 27.430 71.650 27.490 ;
        RECT 73.430 27.420 73.670 27.500 ;
        RECT 75.610 27.420 75.990 27.510 ;
        RECT 77.360 27.420 77.600 27.490 ;
        RECT 79.640 27.420 80.040 27.540 ;
        RECT 80.720 27.420 81.120 27.540 ;
        RECT 83.160 27.420 83.400 27.490 ;
        RECT 84.770 27.420 85.150 27.570 ;
        RECT 89.290 27.490 89.660 33.420 ;
        RECT 89.730 33.130 90.240 33.430 ;
        RECT 89.730 32.880 89.970 33.130 ;
        RECT 90.610 33.040 90.930 33.360 ;
        RECT 91.730 33.340 92.310 33.580 ;
        RECT 89.720 32.560 89.980 32.880 ;
        RECT 89.730 31.240 89.970 32.560 ;
        RECT 90.610 32.170 90.930 32.490 ;
        RECT 91.750 32.190 92.310 33.340 ;
        RECT 92.450 33.030 93.200 33.630 ;
        RECT 92.560 32.500 93.200 33.030 ;
        RECT 91.730 31.950 92.310 32.190 ;
        RECT 90.610 31.620 90.930 31.940 ;
        RECT 91.750 31.250 92.310 31.950 ;
        RECT 92.450 31.900 93.200 32.500 ;
        RECT 92.560 31.250 93.200 31.900 ;
        RECT 87.090 27.420 87.330 27.480 ;
        RECT 89.110 27.430 89.270 27.490 ;
        RECT 89.290 27.430 89.670 27.490 ;
        RECT 89.920 27.430 90.080 27.490 ;
        RECT 70.480 25.110 70.720 27.420 ;
        RECT 89.290 26.450 89.660 27.430 ;
        RECT 89.250 25.940 89.740 26.450 ;
        RECT 89.290 25.910 89.660 25.940 ;
        RECT 70.480 24.870 71.060 25.110 ;
        RECT 68.480 22.870 68.800 23.190 ;
        RECT 65.180 21.790 65.430 22.330 ;
        RECT 68.630 22.190 68.950 22.510 ;
        RECT 61.480 21.120 61.850 21.130 ;
        RECT 61.430 20.860 61.850 21.120 ;
        RECT 61.480 20.840 61.850 20.860 ;
        RECT 57.120 20.510 57.380 20.530 ;
        RECT 56.650 19.430 56.990 19.770 ;
        RECT 56.690 19.410 56.910 19.430 ;
        RECT 56.080 17.140 56.360 17.460 ;
        RECT 56.690 17.130 56.890 19.410 ;
        RECT 57.040 18.470 57.360 18.790 ;
        RECT 57.150 17.940 57.340 17.950 ;
        RECT 57.090 17.620 57.410 17.940 ;
        RECT 57.150 17.450 57.340 17.620 ;
        RECT 54.650 16.750 54.990 17.040 ;
        RECT 56.650 16.810 56.930 17.130 ;
        RECT 57.110 17.120 57.390 17.450 ;
        RECT 44.510 15.030 44.820 16.240 ;
        RECT 48.370 15.990 49.230 16.270 ;
        RECT 48.290 15.980 49.230 15.990 ;
        RECT 49.390 16.380 49.690 16.490 ;
        RECT 48.290 15.510 48.750 15.980 ;
        RECT 44.460 14.550 44.880 15.030 ;
        RECT 49.390 14.870 49.580 16.380 ;
        RECT 50.340 16.190 50.660 16.510 ;
        RECT 53.020 15.980 53.770 16.170 ;
        RECT 53.270 15.140 53.770 15.980 ;
        RECT 57.580 15.900 57.760 20.530 ;
        RECT 60.900 20.470 61.090 20.720 ;
        RECT 60.620 20.460 61.090 20.470 ;
        RECT 60.410 20.140 61.090 20.460 ;
        RECT 61.480 20.330 61.850 20.350 ;
        RECT 60.410 19.820 60.570 20.140 ;
        RECT 60.620 19.980 61.090 20.140 ;
        RECT 61.430 20.070 61.850 20.330 ;
        RECT 61.480 20.060 61.850 20.070 ;
        RECT 60.410 19.540 60.760 19.820 ;
        RECT 60.900 19.720 61.090 19.980 ;
        RECT 60.410 19.280 60.570 19.540 ;
        RECT 60.250 18.960 60.570 19.280 ;
        RECT 60.900 19.430 61.130 19.720 ;
        RECT 60.900 18.830 61.090 19.430 ;
        RECT 60.440 18.440 60.760 18.720 ;
        RECT 60.900 18.540 61.130 18.830 ;
        RECT 60.900 18.280 61.090 18.540 ;
        RECT 60.620 17.850 61.090 18.280 ;
        RECT 61.480 18.190 61.850 18.200 ;
        RECT 61.430 17.930 61.850 18.190 ;
        RECT 61.480 17.910 61.850 17.930 ;
        RECT 60.620 17.790 61.120 17.850 ;
        RECT 58.900 17.060 59.160 17.090 ;
        RECT 58.880 16.760 59.180 17.060 ;
        RECT 58.900 16.750 59.160 16.760 ;
        RECT 57.580 15.600 58.060 15.900 ;
        RECT 58.910 15.830 59.130 16.750 ;
        RECT 60.870 16.620 61.120 17.790 ;
        RECT 62.210 17.570 62.440 21.420 ;
        RECT 63.940 21.110 64.280 21.150 ;
        RECT 63.940 21.070 64.500 21.110 ;
        RECT 63.820 20.900 64.500 21.070 ;
        RECT 63.940 20.880 64.500 20.900 ;
        RECT 63.940 20.830 64.280 20.880 ;
        RECT 65.180 20.720 65.820 21.790 ;
        RECT 68.630 21.300 68.950 21.620 ;
        RECT 65.180 20.470 65.430 20.720 ;
        RECT 68.480 20.620 68.800 20.940 ;
        RECT 63.940 20.310 64.280 20.360 ;
        RECT 63.940 20.290 64.500 20.310 ;
        RECT 63.820 20.120 64.500 20.290 ;
        RECT 63.940 20.080 64.500 20.120 ;
        RECT 63.940 20.040 64.280 20.080 ;
        RECT 65.180 19.400 65.820 20.470 ;
        RECT 68.480 20.100 68.800 20.420 ;
        RECT 68.630 19.420 68.950 19.740 ;
        RECT 65.180 18.860 65.430 19.400 ;
        RECT 63.940 18.180 64.280 18.220 ;
        RECT 63.940 18.140 64.500 18.180 ;
        RECT 63.820 17.970 64.500 18.140 ;
        RECT 63.940 17.950 64.500 17.970 ;
        RECT 63.940 17.900 64.280 17.950 ;
        RECT 62.930 17.600 63.310 17.700 ;
        RECT 64.880 16.640 65.150 17.870 ;
        RECT 65.180 17.790 65.820 18.860 ;
        RECT 68.630 18.530 68.950 18.850 ;
        RECT 68.480 17.850 68.800 18.170 ;
        RECT 65.180 17.570 65.430 17.790 ;
        RECT 69.560 17.600 69.790 23.650 ;
        RECT 70.820 23.530 71.060 24.870 ;
        RECT 70.820 19.300 71.050 23.530 ;
        RECT 75.940 22.470 76.200 22.530 ;
        RECT 75.930 22.210 76.200 22.470 ;
        RECT 75.420 21.280 75.680 21.600 ;
        RECT 74.950 19.440 75.210 19.760 ;
        RECT 70.780 19.290 71.060 19.300 ;
        RECT 70.780 18.970 71.080 19.290 ;
        RECT 67.700 17.070 68.130 17.470 ;
        RECT 60.860 16.360 61.180 16.620 ;
        RECT 64.880 16.330 65.230 16.640 ;
        RECT 57.660 15.490 58.060 15.600 ;
        RECT 58.850 15.430 59.190 15.830 ;
        RECT 58.910 15.350 59.130 15.430 ;
        RECT 62.860 15.160 63.800 16.090 ;
        RECT 67.740 15.280 68.090 17.070 ;
        RECT 69.560 16.510 69.780 17.600 ;
        RECT 70.820 17.110 71.050 18.970 ;
        RECT 74.450 18.510 74.710 18.830 ;
        RECT 70.820 16.880 74.030 17.110 ;
        RECT 70.820 16.870 71.050 16.880 ;
        RECT 69.270 16.270 69.780 16.510 ;
        RECT 48.950 14.550 49.580 14.870 ;
        RECT 52.780 14.820 53.020 15.140 ;
        RECT 54.020 14.820 54.260 15.140 ;
        RECT 62.590 14.840 62.830 15.160 ;
        RECT 63.830 14.840 64.070 15.160 ;
        RECT 69.270 15.020 69.500 16.270 ;
        RECT 73.800 15.910 74.030 16.880 ;
        RECT 73.750 15.510 74.060 15.910 ;
        RECT 69.160 14.580 69.620 15.020 ;
        RECT 48.950 14.450 49.390 14.550 ;
        RECT 52.780 13.480 53.020 13.800 ;
        RECT 54.020 13.470 54.260 13.790 ;
        RECT 62.590 13.500 62.830 13.820 ;
        RECT 63.830 13.490 64.070 13.810 ;
        RECT 73.800 12.340 74.030 15.510 ;
        RECT 73.670 12.120 74.030 12.340 ;
        RECT 52.380 11.850 52.640 12.050 ;
        RECT 54.400 11.850 54.660 12.050 ;
        RECT 49.110 11.330 49.430 11.650 ;
        RECT 50.200 11.330 50.520 11.650 ;
        RECT 51.300 11.320 51.620 11.640 ;
        RECT 52.380 11.040 52.690 11.850 ;
        RECT 54.350 11.040 54.660 11.850 ;
        RECT 62.190 11.880 62.450 12.080 ;
        RECT 64.210 11.880 64.470 12.080 ;
        RECT 73.470 11.890 74.030 12.120 ;
        RECT 73.470 11.880 74.010 11.890 ;
        RECT 55.420 11.320 55.740 11.640 ;
        RECT 56.520 11.330 56.840 11.650 ;
        RECT 57.610 11.330 57.930 11.650 ;
        RECT 58.920 11.360 59.240 11.680 ;
        RECT 60.010 11.360 60.330 11.680 ;
        RECT 61.110 11.350 61.430 11.670 ;
        RECT 62.190 11.070 62.500 11.880 ;
        RECT 64.160 11.070 64.470 11.880 ;
        RECT 65.230 11.350 65.550 11.670 ;
        RECT 66.330 11.360 66.650 11.680 ;
        RECT 67.420 11.360 67.740 11.680 ;
        RECT 70.970 11.330 71.290 11.650 ;
        RECT 72.070 11.340 72.390 11.660 ;
        RECT 73.160 11.340 73.480 11.660 ;
        RECT 49.160 9.270 49.480 11.020 ;
        RECT 49.660 10.650 49.980 10.970 ;
        RECT 50.750 10.630 51.070 10.950 ;
        RECT 51.860 10.620 52.180 10.940 ;
        RECT 49.660 9.280 49.980 9.600 ;
        RECT 50.750 9.280 51.070 9.600 ;
        RECT 51.850 9.280 52.170 9.600 ;
        RECT 49.040 8.670 49.580 9.270 ;
        RECT 49.100 8.550 49.420 8.670 ;
        RECT 50.200 8.550 50.520 8.870 ;
        RECT 51.300 8.550 51.620 8.870 ;
        RECT 49.100 7.180 49.420 7.500 ;
        RECT 50.200 7.180 50.520 7.500 ;
        RECT 51.300 7.180 51.620 7.500 ;
        RECT 48.530 6.540 48.850 6.860 ;
        RECT 49.660 6.500 49.980 6.820 ;
        RECT 50.750 6.500 51.070 6.820 ;
        RECT 51.850 6.510 52.170 6.830 ;
        RECT 48.540 6.070 48.860 6.390 ;
        RECT 52.380 6.060 52.640 11.040 ;
        RECT 52.780 10.710 53.020 11.030 ;
        RECT 54.020 10.700 54.260 11.020 ;
        RECT 54.400 6.060 54.660 11.040 ;
        RECT 54.860 10.620 55.180 10.940 ;
        RECT 55.970 10.630 56.290 10.950 ;
        RECT 57.060 10.650 57.380 10.970 ;
        RECT 54.870 9.280 55.190 9.600 ;
        RECT 55.970 9.280 56.290 9.600 ;
        RECT 57.060 9.280 57.380 9.600 ;
        RECT 57.530 8.870 57.870 11.040 ;
        RECT 58.960 8.900 59.300 11.030 ;
        RECT 59.470 10.680 59.790 11.000 ;
        RECT 60.560 10.660 60.880 10.980 ;
        RECT 61.670 10.650 61.990 10.970 ;
        RECT 59.470 9.310 59.790 9.630 ;
        RECT 60.560 9.310 60.880 9.630 ;
        RECT 61.660 9.310 61.980 9.630 ;
        RECT 55.420 8.550 55.740 8.870 ;
        RECT 56.520 8.550 56.840 8.870 ;
        RECT 57.530 8.550 57.940 8.870 ;
        RECT 58.910 8.580 59.300 8.900 ;
        RECT 60.010 8.580 60.330 8.900 ;
        RECT 61.110 8.580 61.430 8.900 ;
        RECT 57.530 8.250 57.870 8.550 ;
        RECT 57.470 7.730 57.930 8.250 ;
        RECT 58.960 7.530 59.300 8.580 ;
        RECT 55.420 7.180 55.740 7.500 ;
        RECT 56.520 7.180 56.840 7.500 ;
        RECT 57.620 7.180 57.940 7.500 ;
        RECT 58.910 7.360 59.300 7.530 ;
        RECT 58.340 6.860 58.660 6.890 ;
        RECT 54.870 6.510 55.190 6.830 ;
        RECT 55.970 6.500 56.290 6.820 ;
        RECT 57.060 6.500 57.380 6.820 ;
        RECT 58.190 6.570 58.660 6.860 ;
        RECT 58.870 6.840 59.390 7.360 ;
        RECT 60.010 7.210 60.330 7.530 ;
        RECT 61.110 7.210 61.430 7.530 ;
        RECT 58.190 6.540 58.510 6.570 ;
        RECT 59.470 6.530 59.790 6.850 ;
        RECT 60.560 6.530 60.880 6.850 ;
        RECT 61.660 6.540 61.980 6.860 ;
        RECT 58.350 6.390 58.670 6.420 ;
        RECT 58.180 6.100 58.670 6.390 ;
        RECT 58.180 6.070 58.500 6.100 ;
        RECT 62.190 6.090 62.450 11.070 ;
        RECT 62.590 10.730 62.830 11.050 ;
        RECT 63.830 10.730 64.070 11.050 ;
        RECT 64.210 6.090 64.470 11.070 ;
        RECT 64.670 10.650 64.990 10.970 ;
        RECT 65.780 10.660 66.100 10.980 ;
        RECT 66.870 10.680 67.190 11.000 ;
        RECT 64.680 9.310 65.000 9.630 ;
        RECT 65.780 9.310 66.100 9.630 ;
        RECT 66.870 9.310 67.190 9.630 ;
        RECT 67.380 8.900 67.650 11.070 ;
        RECT 70.410 10.630 70.730 10.950 ;
        RECT 71.520 10.640 71.840 10.960 ;
        RECT 72.610 10.660 72.930 10.980 ;
        RECT 74.450 10.670 74.700 18.510 ;
        RECT 74.950 11.570 75.200 19.440 ;
        RECT 75.430 12.480 75.680 21.280 ;
        RECT 75.930 13.370 76.180 22.210 ;
        RECT 91.770 14.870 92.270 31.250 ;
        RECT 92.700 20.150 93.200 31.250 ;
        RECT 93.830 25.380 94.330 51.650 ;
        RECT 94.960 39.710 95.460 52.270 ;
        RECT 97.070 45.260 97.490 45.410 ;
        RECT 98.100 45.260 98.520 45.410 ;
        RECT 101.800 45.330 102.030 45.410 ;
        RECT 97.070 45.120 98.520 45.260 ;
        RECT 102.060 43.180 102.480 49.230 ;
        RECT 105.760 48.020 105.990 49.230 ;
        RECT 110.760 48.410 111.070 48.850 ;
        RECT 105.760 47.230 106.020 48.020 ;
        RECT 108.180 47.660 108.380 47.690 ;
        RECT 105.760 45.080 105.990 47.230 ;
        RECT 108.090 47.160 108.400 47.660 ;
        RECT 110.910 47.450 111.230 47.770 ;
        RECT 108.180 45.410 108.380 47.160 ;
        RECT 111.690 46.790 111.880 64.190 ;
        RECT 115.030 55.340 115.850 55.430 ;
        RECT 114.970 54.650 115.850 55.340 ;
        RECT 112.280 47.770 112.470 49.230 ;
        RECT 112.720 48.580 113.000 49.230 ;
        RECT 112.610 47.980 113.000 48.580 ;
        RECT 112.280 47.740 112.500 47.770 ;
        RECT 112.260 47.470 112.510 47.740 ;
        RECT 112.270 47.460 112.510 47.470 ;
        RECT 112.270 47.220 112.500 47.460 ;
        RECT 111.690 46.660 112.120 46.790 ;
        RECT 111.690 46.340 112.140 46.660 ;
        RECT 111.690 46.060 111.880 46.340 ;
        RECT 111.690 45.740 112.140 46.060 ;
        RECT 111.690 45.620 112.120 45.740 ;
        RECT 108.180 45.330 108.510 45.410 ;
        RECT 108.760 45.390 109.040 45.410 ;
        RECT 108.760 45.330 109.100 45.390 ;
        RECT 105.760 44.290 106.020 45.080 ;
        RECT 105.760 43.180 105.990 44.290 ;
        RECT 108.180 43.240 108.380 45.330 ;
        RECT 108.780 45.090 109.100 45.330 ;
        RECT 110.510 45.070 110.830 45.390 ;
        RECT 111.690 45.110 111.880 45.620 ;
        RECT 112.310 45.410 112.470 47.220 ;
        RECT 112.720 46.380 113.000 47.980 ;
        RECT 112.720 46.060 113.080 46.380 ;
        RECT 112.720 45.410 113.000 46.060 ;
        RECT 112.310 45.190 113.000 45.410 ;
        RECT 113.110 45.260 113.390 45.410 ;
        RECT 110.910 44.690 111.230 45.010 ;
        RECT 111.490 44.790 111.880 45.110 ;
        RECT 112.270 44.940 113.000 45.190 ;
        RECT 110.660 44.240 110.980 44.560 ;
        RECT 111.690 44.460 111.880 44.790 ;
        RECT 112.260 44.670 113.000 44.940 ;
        RECT 111.440 44.140 111.880 44.460 ;
        RECT 109.080 43.680 109.400 44.000 ;
        RECT 109.550 43.710 109.870 44.030 ;
        RECT 110.080 43.560 110.310 43.850 ;
        RECT 110.650 43.680 111.070 44.000 ;
        RECT 110.760 43.560 111.070 43.680 ;
        RECT 111.210 43.630 111.440 43.860 ;
        RECT 111.690 43.630 111.880 44.140 ;
        RECT 111.210 43.570 111.880 43.630 ;
        RECT 100.280 42.690 100.750 43.180 ;
        RECT 107.670 43.020 107.900 43.210 ;
        RECT 107.670 42.920 108.020 43.020 ;
        RECT 108.170 42.950 108.400 43.240 ;
        RECT 110.100 43.090 110.290 43.560 ;
        RECT 110.770 43.550 110.980 43.560 ;
        RECT 110.750 43.230 111.010 43.550 ;
        RECT 107.680 42.700 108.020 42.920 ;
        RECT 94.730 39.410 95.460 39.710 ;
        RECT 94.960 30.550 95.460 39.410 ;
        RECT 94.910 29.990 95.460 30.550 ;
        RECT 93.820 24.820 94.340 25.380 ;
        RECT 92.690 19.630 93.210 20.150 ;
        RECT 91.610 14.300 92.270 14.870 ;
        RECT 75.880 12.790 76.250 13.370 ;
        RECT 75.350 11.900 75.720 12.480 ;
        RECT 74.860 10.990 75.230 11.570 ;
        RECT 70.420 9.290 70.740 9.610 ;
        RECT 71.520 9.290 71.840 9.610 ;
        RECT 72.610 9.290 72.930 9.610 ;
        RECT 65.230 8.580 65.550 8.900 ;
        RECT 66.330 8.580 66.650 8.900 ;
        RECT 67.380 8.580 67.750 8.900 ;
        RECT 73.120 8.880 73.450 10.450 ;
        RECT 74.390 10.100 74.740 10.670 ;
        RECT 67.380 7.530 67.650 8.580 ;
        RECT 70.970 8.560 71.290 8.880 ;
        RECT 72.070 8.560 72.390 8.880 ;
        RECT 73.120 8.560 73.490 8.880 ;
        RECT 65.230 7.210 65.550 7.530 ;
        RECT 66.330 7.210 66.650 7.530 ;
        RECT 67.380 7.210 67.750 7.530 ;
        RECT 73.120 7.510 73.450 8.560 ;
        RECT 73.890 8.000 74.170 8.530 ;
        RECT 73.890 7.700 74.350 8.000 ;
        RECT 73.880 7.680 74.350 7.700 ;
        RECT 64.680 6.540 65.000 6.860 ;
        RECT 65.780 6.530 66.100 6.850 ;
        RECT 66.870 6.530 67.190 6.850 ;
        RECT 67.380 6.480 67.650 7.210 ;
        RECT 70.970 7.190 71.290 7.510 ;
        RECT 72.070 7.190 72.390 7.510 ;
        RECT 73.120 7.190 73.490 7.510 ;
        RECT 73.880 7.250 74.170 7.680 ;
        RECT 68.000 6.570 68.320 6.890 ;
        RECT 70.420 6.520 70.740 6.840 ;
        RECT 71.520 6.510 71.840 6.830 ;
        RECT 72.610 6.510 72.930 6.830 ;
        RECT 67.270 5.920 67.760 6.480 ;
        RECT 67.990 6.100 68.310 6.420 ;
        RECT 41.170 3.700 41.820 5.020 ;
        RECT 73.120 0.460 73.450 7.190 ;
        RECT 73.740 6.550 74.060 6.870 ;
        RECT 73.730 6.080 74.050 6.400 ;
        RECT 91.770 5.990 92.270 14.300 ;
        RECT 92.700 6.900 93.200 19.630 ;
        RECT 93.830 7.770 94.330 24.820 ;
        RECT 94.960 9.280 95.460 29.990 ;
        RECT 100.330 39.710 100.730 42.690 ;
        RECT 101.250 42.080 101.670 42.440 ;
        RECT 107.680 42.270 108.020 42.490 ;
        RECT 107.670 42.170 108.020 42.270 ;
        RECT 108.180 42.240 108.380 42.950 ;
        RECT 110.030 42.770 110.290 43.090 ;
        RECT 110.280 42.430 110.600 42.750 ;
        RECT 100.330 39.410 100.850 39.710 ;
        RECT 97.850 16.840 98.430 17.400 ;
        RECT 97.880 16.830 98.390 16.840 ;
        RECT 94.960 8.720 95.520 9.280 ;
        RECT 94.960 8.590 95.460 8.720 ;
        RECT 97.880 4.960 98.380 16.830 ;
        RECT 97.250 3.680 98.380 4.960 ;
        RECT 99.130 4.200 99.360 6.270 ;
        RECT 99.120 3.970 99.410 4.200 ;
        RECT 99.130 2.590 99.360 3.970 ;
        RECT 99.120 2.360 99.410 2.590 ;
        RECT 99.130 0.990 99.360 2.360 ;
        RECT 99.120 0.760 99.410 0.990 ;
        RECT 73.060 0.070 73.490 0.460 ;
        RECT 39.520 -0.590 39.890 -0.210 ;
        RECT 99.130 -0.630 99.360 0.760 ;
        RECT 100.330 -0.100 100.730 39.410 ;
        RECT 100.330 -0.120 100.860 -0.100 ;
        RECT 101.260 -0.120 101.650 42.080 ;
        RECT 107.670 41.980 107.900 42.170 ;
        RECT 108.170 41.950 108.400 42.240 ;
        RECT 110.030 42.100 110.290 42.420 ;
        RECT 108.180 40.220 108.380 41.950 ;
        RECT 110.100 41.630 110.290 42.100 ;
        RECT 110.770 41.940 110.980 43.230 ;
        RECT 111.210 43.080 111.400 43.570 ;
        RECT 111.440 43.310 111.880 43.570 ;
        RECT 111.690 43.240 111.880 43.310 ;
        RECT 111.040 42.830 111.400 43.080 ;
        RECT 111.670 42.980 111.900 43.240 ;
        RECT 112.280 43.180 113.000 44.670 ;
        RECT 113.120 43.830 113.390 45.260 ;
        RECT 113.740 44.840 114.060 45.160 ;
        RECT 113.120 43.540 113.400 43.830 ;
        RECT 111.490 42.950 111.900 42.980 ;
        RECT 111.040 42.760 111.300 42.830 ;
        RECT 111.490 42.660 111.880 42.950 ;
        RECT 111.040 42.360 111.300 42.430 ;
        RECT 111.040 42.110 111.400 42.360 ;
        RECT 111.690 42.240 111.880 42.660 ;
        RECT 111.670 42.150 111.900 42.240 ;
        RECT 110.750 41.650 110.980 41.940 ;
        RECT 109.080 41.190 109.400 41.510 ;
        RECT 110.080 41.340 110.310 41.630 ;
        RECT 111.210 41.620 111.400 42.110 ;
        RECT 111.490 41.950 111.900 42.150 ;
        RECT 111.490 41.830 111.880 41.950 ;
        RECT 110.650 41.190 110.970 41.510 ;
        RECT 111.210 41.500 111.440 41.620 ;
        RECT 111.690 41.500 111.880 41.830 ;
        RECT 111.210 41.330 111.880 41.500 ;
        RECT 111.440 41.180 111.880 41.330 ;
        RECT 109.080 40.660 109.400 40.980 ;
        RECT 110.080 40.540 110.310 40.830 ;
        RECT 110.650 40.660 110.970 40.980 ;
        RECT 111.210 40.670 111.440 40.840 ;
        RECT 111.690 40.670 111.880 41.180 ;
        RECT 111.210 40.550 111.880 40.670 ;
        RECT 102.170 39.690 102.620 40.120 ;
        RECT 107.670 40.000 107.900 40.190 ;
        RECT 107.670 39.900 108.020 40.000 ;
        RECT 108.170 39.930 108.400 40.220 ;
        RECT 110.100 40.070 110.290 40.540 ;
        RECT 102.190 -0.120 102.580 39.690 ;
        RECT 107.680 39.680 108.020 39.900 ;
        RECT 103.030 39.430 103.410 39.440 ;
        RECT 103.010 39.130 103.430 39.430 ;
        RECT 107.680 39.250 108.020 39.470 ;
        RECT 107.670 39.150 108.020 39.250 ;
        RECT 108.180 39.410 108.380 39.930 ;
        RECT 110.030 39.750 110.290 40.070 ;
        RECT 111.210 40.060 111.400 40.550 ;
        RECT 111.440 40.350 111.880 40.550 ;
        RECT 111.690 40.220 111.880 40.350 ;
        RECT 111.040 39.860 111.400 40.060 ;
        RECT 111.670 40.020 111.900 40.220 ;
        RECT 110.920 39.810 111.400 39.860 ;
        RECT 111.490 39.930 111.900 40.020 ;
        RECT 110.920 39.740 111.300 39.810 ;
        RECT 110.920 39.560 111.240 39.740 ;
        RECT 111.490 39.700 111.880 39.930 ;
        RECT 111.690 39.560 111.880 39.700 ;
        RECT 112.450 39.560 112.790 43.180 ;
        RECT 110.920 39.500 112.790 39.560 ;
        RECT 110.970 39.420 112.790 39.500 ;
        RECT 108.180 39.360 108.510 39.410 ;
        RECT 108.760 39.360 109.040 39.410 ;
        RECT 108.180 39.220 108.380 39.360 ;
        RECT 100.330 -0.320 102.850 -0.120 ;
        RECT 38.870 -1.210 39.260 -0.820 ;
        RECT 99.120 -0.860 99.410 -0.630 ;
        RECT 100.330 -0.660 100.730 -0.320 ;
        RECT 38.270 -1.840 38.650 -1.450 ;
        RECT 37.680 -2.470 38.030 -2.100 ;
        RECT 99.130 -2.230 99.360 -0.860 ;
        RECT 100.320 -1.120 100.790 -0.660 ;
        RECT 101.260 -1.460 101.650 -0.320 ;
        RECT 99.850 -1.840 100.170 -1.760 ;
        RECT 101.230 -1.840 101.690 -1.460 ;
        RECT 99.850 -2.020 101.940 -1.840 ;
        RECT 101.430 -2.060 101.940 -2.020 ;
        RECT 101.650 -2.070 101.940 -2.060 ;
        RECT 99.120 -2.460 99.410 -2.230 ;
        RECT 102.190 -2.280 102.580 -0.320 ;
        RECT 37.040 -3.150 37.400 -2.770 ;
        RECT 36.450 -3.390 36.790 -3.380 ;
        RECT 36.430 -3.760 36.810 -3.390 ;
        RECT 36.450 -3.770 36.780 -3.760 ;
        RECT 99.130 -3.850 99.360 -2.460 ;
        RECT 102.170 -2.740 102.640 -2.280 ;
        RECT 102.680 -3.350 102.850 -0.320 ;
        RECT 103.030 -3.080 103.410 39.130 ;
        RECT 107.670 38.960 107.900 39.150 ;
        RECT 108.170 38.930 108.400 39.220 ;
        RECT 110.030 39.080 110.290 39.400 ;
        RECT 111.040 39.340 111.300 39.410 ;
        RECT 111.040 39.090 111.400 39.340 ;
        RECT 111.690 39.220 111.880 39.420 ;
        RECT 112.450 39.360 112.790 39.420 ;
        RECT 113.120 41.240 113.390 43.540 ;
        RECT 113.790 42.620 114.110 42.940 ;
        RECT 113.780 41.900 114.100 42.220 ;
        RECT 113.120 40.950 113.400 41.240 ;
        RECT 113.120 39.360 113.390 40.950 ;
        RECT 113.700 39.650 114.020 39.970 ;
        RECT 108.180 38.060 108.380 38.930 ;
        RECT 110.100 38.610 110.290 39.080 ;
        RECT 109.080 38.170 109.400 38.490 ;
        RECT 110.080 38.320 110.310 38.610 ;
        RECT 111.210 38.600 111.400 39.090 ;
        RECT 111.670 38.930 111.900 39.220 ;
        RECT 110.650 38.170 110.970 38.490 ;
        RECT 111.210 38.310 111.440 38.600 ;
        RECT 111.690 38.060 111.880 38.930 ;
        RECT 114.970 35.650 115.680 54.650 ;
        RECT 114.840 34.860 115.680 35.650 ;
        RECT 110.560 16.820 111.280 17.390 ;
        RECT 110.620 9.810 111.130 16.820 ;
        RECT 110.480 9.760 111.130 9.810 ;
        RECT 110.470 9.580 111.130 9.760 ;
        RECT 110.440 9.570 111.130 9.580 ;
        RECT 110.440 9.200 111.040 9.570 ;
        RECT 110.440 7.330 111.020 9.200 ;
        RECT 110.090 6.340 111.020 7.330 ;
        RECT 110.440 5.560 111.020 6.340 ;
        RECT 110.450 4.950 111.020 5.560 ;
        RECT 110.440 3.950 111.020 4.950 ;
        RECT 104.630 3.190 104.950 3.510 ;
        RECT 110.450 3.350 111.020 3.950 ;
        RECT 104.630 2.520 104.950 2.840 ;
        RECT 104.750 1.550 105.070 1.600 ;
        RECT 104.520 1.320 105.070 1.550 ;
        RECT 104.750 1.280 105.070 1.320 ;
        RECT 104.750 -0.060 105.070 -0.010 ;
        RECT 104.520 -0.290 105.070 -0.060 ;
        RECT 104.750 -0.330 105.070 -0.290 ;
        RECT 104.740 -1.670 105.060 -1.620 ;
        RECT 104.510 -1.900 105.060 -1.670 ;
        RECT 104.740 -1.940 105.060 -1.900 ;
        RECT 102.260 -3.570 102.850 -3.350 ;
        RECT 103.000 -3.540 103.440 -3.080 ;
        RECT 104.740 -3.290 105.060 -3.240 ;
        RECT 104.510 -3.520 105.060 -3.290 ;
        RECT 104.740 -3.560 105.060 -3.520 ;
        RECT 102.260 -3.580 102.550 -3.570 ;
        RECT 99.120 -4.080 99.410 -3.850 ;
        RECT 34.670 -5.610 35.020 -5.280 ;
        RECT 99.130 -5.450 99.360 -4.080 ;
        RECT 110.440 -4.090 111.020 3.350 ;
        RECT 110.450 -4.690 111.020 -4.090 ;
        RECT 104.740 -4.900 105.060 -4.850 ;
        RECT 104.510 -5.130 105.060 -4.900 ;
        RECT 104.740 -5.170 105.060 -5.130 ;
        RECT 34.690 -5.670 35.020 -5.610 ;
        RECT 99.120 -5.680 99.410 -5.450 ;
        RECT 110.440 -5.510 111.020 -4.690 ;
        RECT 110.440 -5.520 110.980 -5.510 ;
        RECT 33.400 -6.890 33.750 -6.560 ;
        RECT 33.400 -6.960 33.730 -6.890 ;
        RECT 99.130 -7.070 99.360 -5.680 ;
        RECT 104.370 -6.770 104.690 -6.450 ;
        RECT 104.420 -7.000 104.650 -6.770 ;
        RECT 31.260 -7.620 32.500 -7.290 ;
        RECT 32.790 -7.590 33.230 -7.170 ;
        RECT 99.120 -7.300 99.410 -7.070 ;
        RECT 31.260 -7.730 31.840 -7.620 ;
        RECT 104.750 -8.100 105.070 -8.050 ;
        RECT 104.520 -8.330 105.070 -8.100 ;
        RECT 104.750 -8.370 105.070 -8.330 ;
        RECT 104.740 -9.690 105.060 -9.640 ;
        RECT 101.540 -9.770 101.860 -9.720 ;
        RECT 102.480 -9.770 102.800 -9.720 ;
        RECT 101.310 -10.000 101.860 -9.770 ;
        RECT 102.250 -10.000 102.800 -9.770 ;
        RECT 103.430 -9.830 103.750 -9.780 ;
        RECT 101.540 -10.040 101.860 -10.000 ;
        RECT 102.480 -10.040 102.800 -10.000 ;
        RECT 103.200 -10.060 103.750 -9.830 ;
        RECT 104.510 -9.920 105.060 -9.690 ;
        RECT 104.740 -9.960 105.060 -9.920 ;
        RECT 103.430 -10.100 103.750 -10.060 ;
      LAYER via ;
        RECT 4.210 62.150 4.600 62.540 ;
        RECT 6.630 61.230 6.890 61.490 ;
        RECT 9.490 61.280 9.750 61.540 ;
        RECT 6.620 60.200 6.880 60.460 ;
        RECT 7.340 60.170 7.600 60.430 ;
        RECT 8.030 60.210 8.290 60.470 ;
        RECT 6.620 59.750 6.880 60.010 ;
        RECT 8.030 59.770 8.290 60.030 ;
        RECT 6.620 59.330 6.880 59.590 ;
        RECT 7.340 59.330 7.600 59.590 ;
        RECT 8.050 59.350 8.310 59.610 ;
        RECT 4.290 58.700 4.680 59.090 ;
        RECT 6.620 57.980 6.880 58.240 ;
        RECT 5.670 57.530 5.930 57.790 ;
        RECT 9.180 59.740 9.440 60.000 ;
        RECT 22.730 59.430 22.990 59.690 ;
        RECT 24.090 59.510 24.350 59.770 ;
        RECT 24.780 59.500 25.040 59.760 ;
        RECT 8.760 57.730 9.020 57.990 ;
        RECT 7.320 56.530 7.580 56.790 ;
        RECT 8.750 56.550 9.010 56.810 ;
        RECT 6.530 55.950 6.790 56.210 ;
        RECT 7.460 55.950 7.720 56.210 ;
        RECT 8.160 55.950 8.420 56.210 ;
        RECT 8.900 55.950 9.160 56.210 ;
        RECT 9.610 55.940 9.870 56.200 ;
        RECT 5.590 54.830 6.010 55.250 ;
        RECT 22.010 55.770 22.270 56.030 ;
        RECT 11.540 53.430 11.830 54.010 ;
        RECT 24.830 52.370 25.090 52.630 ;
        RECT 19.920 46.530 20.180 46.790 ;
        RECT 21.010 46.540 21.270 46.800 ;
        RECT 18.750 46.120 19.010 46.380 ;
        RECT 19.450 46.120 19.710 46.380 ;
        RECT 19.920 45.610 20.180 45.870 ;
        RECT 21.010 45.620 21.270 45.880 ;
        RECT 18.720 45.200 18.980 45.460 ;
        RECT 19.450 45.200 19.710 45.460 ;
        RECT 19.920 44.690 20.180 44.950 ;
        RECT 21.010 44.700 21.270 44.960 ;
        RECT 18.730 44.280 18.990 44.540 ;
        RECT 19.450 44.280 19.710 44.540 ;
        RECT 18.080 43.260 18.340 43.520 ;
        RECT 18.040 42.300 18.300 42.560 ;
        RECT 18.080 41.340 18.340 41.600 ;
        RECT 19.730 43.710 19.990 43.970 ;
        RECT 21.030 43.610 21.290 43.870 ;
        RECT 19.730 43.250 19.990 43.510 ;
        RECT 19.730 42.750 19.990 43.010 ;
        RECT 21.030 42.650 21.290 42.910 ;
        RECT 19.730 42.290 19.990 42.550 ;
        RECT 19.730 41.790 19.990 42.050 ;
        RECT 21.030 41.690 21.290 41.950 ;
        RECT 19.730 41.330 19.990 41.590 ;
        RECT 31.870 55.790 32.130 56.050 ;
        RECT 30.620 51.940 30.930 52.250 ;
        RECT 47.200 59.580 47.620 60.000 ;
        RECT 43.350 58.820 43.770 59.240 ;
        RECT 48.870 57.210 49.310 57.650 ;
        RECT 54.590 57.210 55.030 57.650 ;
        RECT 66.970 58.820 68.320 59.240 ;
        RECT 56.410 57.180 56.850 57.620 ;
        RECT 44.450 56.190 44.890 56.630 ;
        RECT 41.690 53.170 41.950 53.430 ;
        RECT 34.620 52.480 34.880 52.740 ;
        RECT 33.450 51.490 33.720 51.750 ;
        RECT 22.120 50.710 22.470 51.060 ;
        RECT 27.370 51.020 27.630 51.280 ;
        RECT 50.160 56.190 50.600 56.630 ;
        RECT 42.930 49.860 43.190 50.120 ;
        RECT 40.830 49.020 41.090 49.280 ;
        RECT 23.140 48.470 23.400 48.860 ;
        RECT 39.540 48.480 39.870 48.740 ;
        RECT 22.500 47.650 22.760 48.050 ;
        RECT 18.040 26.060 18.300 26.530 ;
        RECT 18.680 26.060 18.940 26.530 ;
        RECT 16.680 25.030 16.940 25.290 ;
        RECT 16.160 24.630 16.420 24.890 ;
        RECT 6.880 23.380 7.540 24.040 ;
        RECT 18.760 25.010 19.020 25.270 ;
        RECT 20.520 25.020 20.790 25.290 ;
        RECT 18.100 24.650 18.360 24.910 ;
        RECT 18.850 24.050 19.110 24.310 ;
        RECT 19.500 24.050 19.760 24.310 ;
        RECT 17.630 23.610 17.890 23.870 ;
        RECT 18.330 23.610 18.590 23.870 ;
        RECT 20.010 22.880 20.270 23.140 ;
        RECT 17.180 22.260 17.440 22.520 ;
        RECT 16.180 20.720 16.440 20.980 ;
        RECT 12.090 18.860 12.460 19.230 ;
        RECT 6.920 17.520 7.580 18.180 ;
        RECT 16.180 17.630 16.440 17.890 ;
        RECT 19.930 21.750 20.190 22.010 ;
        RECT 21.020 24.630 21.280 24.890 ;
        RECT 19.940 21.210 20.200 21.470 ;
        RECT 17.180 20.710 17.440 20.970 ;
        RECT 19.990 20.260 20.250 20.520 ;
        RECT 17.660 19.730 17.920 19.990 ;
        RECT 18.350 19.720 18.610 19.980 ;
        RECT 18.830 18.950 19.090 19.210 ;
        RECT 19.540 18.890 19.800 19.150 ;
        RECT 19.490 18.070 19.750 18.330 ;
        RECT 17.280 17.640 17.540 17.900 ;
        RECT 18.370 17.640 18.630 17.900 ;
        RECT 19.500 17.600 19.760 17.860 ;
        RECT 16.730 16.960 16.990 17.220 ;
        RECT 17.830 16.960 18.090 17.220 ;
        RECT 18.930 16.960 19.190 17.220 ;
        RECT 16.730 15.590 16.990 15.850 ;
        RECT 17.830 15.590 18.090 15.850 ;
        RECT 18.930 15.590 19.190 15.850 ;
        RECT 16.180 14.860 16.440 15.120 ;
        RECT 17.280 14.860 17.540 15.120 ;
        RECT 18.370 14.860 18.630 15.120 ;
        RECT 16.170 13.520 16.430 13.780 ;
        RECT 17.280 13.510 17.540 13.770 ;
        RECT 18.370 13.490 18.630 13.750 ;
        RECT 12.080 12.620 12.450 12.990 ;
        RECT 16.730 12.820 16.990 13.080 ;
        RECT 17.830 12.810 18.090 13.070 ;
        RECT 18.920 12.810 19.180 13.070 ;
        RECT 19.620 12.200 19.880 12.560 ;
        RECT 15.070 6.960 15.360 7.250 ;
        RECT 19.530 10.510 19.790 10.770 ;
        RECT 16.220 10.070 16.480 10.330 ;
        RECT 17.320 10.080 17.580 10.340 ;
        RECT 18.410 10.080 18.670 10.340 ;
        RECT 19.540 10.040 19.800 10.300 ;
        RECT 16.770 9.400 17.030 9.660 ;
        RECT 17.870 9.400 18.130 9.660 ;
        RECT 18.970 9.400 19.230 9.660 ;
        RECT 16.770 8.030 17.030 8.290 ;
        RECT 17.870 8.030 18.130 8.290 ;
        RECT 18.970 8.030 19.230 8.290 ;
        RECT 16.220 7.300 16.480 7.560 ;
        RECT 17.320 7.300 17.580 7.560 ;
        RECT 18.410 7.300 18.670 7.560 ;
        RECT 22.520 46.540 22.780 46.800 ;
        RECT 22.520 45.620 22.780 45.880 ;
        RECT 22.490 44.700 22.750 44.960 ;
        RECT 38.910 46.760 39.240 47.090 ;
        RECT 38.340 45.280 38.670 45.610 ;
        RECT 23.130 43.610 23.390 43.870 ;
        RECT 37.700 43.680 38.030 44.010 ;
        RECT 37.060 43.110 37.390 43.440 ;
        RECT 23.140 42.650 23.400 42.910 ;
        RECT 23.130 41.690 23.390 41.950 ;
        RECT 22.490 24.030 22.750 24.290 ;
        RECT 21.870 22.880 22.130 23.140 ;
        RECT 21.450 20.270 21.710 20.530 ;
        RECT 21.890 14.580 22.150 15.000 ;
        RECT 21.850 12.200 22.110 12.560 ;
        RECT 36.450 41.540 36.780 41.870 ;
        RECT 35.820 40.010 36.150 40.340 ;
        RECT 35.260 38.440 35.590 38.770 ;
        RECT 34.640 32.970 34.970 33.300 ;
        RECT 34.010 31.380 34.340 31.710 ;
        RECT 33.390 29.830 33.720 30.160 ;
        RECT 32.790 28.350 33.120 28.680 ;
        RECT 32.150 23.180 32.480 23.510 ;
        RECT 31.480 21.610 31.810 21.940 ;
        RECT 23.130 19.700 23.390 19.960 ;
        RECT 30.860 19.970 31.190 20.300 ;
        RECT 22.470 8.570 22.730 8.900 ;
        RECT 21.440 6.950 21.730 7.240 ;
        RECT 16.210 5.960 16.470 6.220 ;
        RECT 17.320 5.950 17.580 6.210 ;
        RECT 18.410 5.930 18.670 6.190 ;
        RECT 20.280 5.940 20.880 6.540 ;
        RECT 16.770 5.260 17.030 5.520 ;
        RECT 17.870 5.250 18.130 5.510 ;
        RECT 18.960 5.250 19.220 5.510 ;
        RECT 30.180 18.530 30.510 18.860 ;
        RECT 26.140 14.170 26.720 14.880 ;
        RECT 23.060 1.010 23.320 1.350 ;
        RECT 4.150 0.070 4.540 0.460 ;
        RECT 30.150 -5.300 30.580 -4.870 ;
        RECT 30.800 -6.090 31.230 -5.660 ;
        RECT 31.470 -6.770 31.870 -6.370 ;
        RECT 31.300 -7.710 31.810 -7.200 ;
        RECT 40.830 47.470 41.090 47.730 ;
        RECT 40.830 45.920 41.090 46.180 ;
        RECT 47.790 49.960 48.050 50.220 ;
        RECT 42.930 48.310 43.190 48.570 ;
        RECT 42.930 46.760 43.190 47.020 ;
        RECT 42.930 45.210 43.190 45.470 ;
        RECT 44.970 49.140 45.230 49.400 ;
        RECT 47.790 48.410 48.050 48.670 ;
        RECT 44.970 47.590 45.230 47.850 ;
        RECT 47.790 46.860 48.050 47.120 ;
        RECT 44.970 46.040 45.230 46.300 ;
        RECT 47.790 45.310 48.050 45.570 ;
        RECT 40.830 44.370 41.090 44.630 ;
        RECT 44.970 44.490 45.230 44.750 ;
        RECT 40.830 42.550 41.090 42.810 ;
        RECT 40.830 41.000 41.090 41.260 ;
        RECT 40.830 39.450 41.090 39.710 ;
        RECT 40.830 37.900 41.090 38.160 ;
        RECT 42.930 41.710 43.190 41.970 ;
        RECT 42.930 40.160 43.190 40.420 ;
        RECT 42.930 38.610 43.190 38.870 ;
        RECT 44.970 42.430 45.230 42.690 ;
        RECT 47.790 41.610 48.050 41.870 ;
        RECT 44.970 40.880 45.230 41.140 ;
        RECT 47.790 40.060 48.050 40.320 ;
        RECT 44.970 39.330 45.230 39.590 ;
        RECT 47.790 38.510 48.050 38.770 ;
        RECT 44.970 37.780 45.230 38.040 ;
        RECT 42.930 37.060 43.190 37.320 ;
        RECT 64.560 56.190 65.000 56.630 ;
        RECT 58.810 52.410 59.070 52.670 ;
        RECT 56.930 48.880 57.190 49.140 ;
        RECT 62.400 51.500 62.660 51.760 ;
        RECT 59.270 50.480 59.530 50.740 ;
        RECT 59.690 48.390 59.950 48.650 ;
        RECT 60.750 47.910 61.010 48.170 ;
        RECT 54.420 43.810 54.680 44.070 ;
        RECT 54.270 42.850 54.530 43.110 ;
        RECT 61.530 43.260 61.790 43.520 ;
        RECT 65.570 52.420 65.830 52.680 ;
        RECT 65.130 51.510 65.390 51.770 ;
        RECT 61.560 42.830 61.820 43.090 ;
        RECT 53.330 41.740 53.590 42.000 ;
        RECT 53.330 41.140 53.590 41.400 ;
        RECT 56.470 40.460 56.730 40.720 ;
        RECT 60.470 42.310 60.730 42.570 ;
        RECT 60.470 41.210 60.730 41.470 ;
        RECT 61.560 40.690 61.820 40.950 ;
        RECT 62.390 40.810 62.660 41.080 ;
        RECT 54.270 40.090 54.530 40.350 ;
        RECT 61.560 39.900 61.820 40.160 ;
        RECT 54.420 39.080 54.680 39.340 ;
        RECT 60.470 39.380 60.730 39.640 ;
        RECT 61.560 39.570 61.820 39.830 ;
        RECT 60.470 38.280 60.730 38.540 ;
        RECT 61.560 37.760 61.820 38.020 ;
        RECT 47.790 36.960 48.050 37.220 ;
        RECT 70.360 56.150 70.800 56.590 ;
        RECT 78.690 57.180 78.970 57.620 ;
        RECT 74.910 50.520 76.130 50.780 ;
        RECT 71.670 49.870 71.930 50.130 ;
        RECT 78.000 49.330 78.260 49.590 ;
        RECT 80.340 52.420 80.600 52.680 ;
        RECT 79.450 51.550 79.710 51.810 ;
        RECT 86.860 61.520 87.230 61.890 ;
        RECT 83.010 53.130 83.270 53.400 ;
        RECT 79.450 47.340 79.710 47.600 ;
        RECT 80.470 47.350 80.730 47.610 ;
        RECT 84.550 48.440 84.810 48.700 ;
        RECT 83.220 47.230 83.650 47.660 ;
        RECT 84.160 46.910 84.420 47.170 ;
        RECT 83.450 46.080 83.710 46.340 ;
        RECT 84.150 45.220 84.410 45.480 ;
        RECT 63.970 42.830 64.230 43.090 ;
        RECT 63.970 40.690 64.230 40.950 ;
        RECT 63.970 39.900 64.230 40.160 ;
        RECT 63.970 37.760 64.230 38.020 ;
        RECT 64.710 37.390 64.970 37.650 ;
        RECT 80.670 43.810 80.930 44.070 ;
        RECT 80.820 42.850 81.080 43.110 ;
        RECT 81.760 41.740 82.020 42.000 ;
        RECT 81.760 41.140 82.020 41.400 ;
        RECT 84.550 43.710 84.810 43.970 ;
        RECT 87.680 58.060 88.050 58.430 ;
        RECT 86.540 45.110 86.800 45.370 ;
        RECT 82.700 41.460 82.960 41.720 ;
        RECT 78.670 40.450 78.930 40.710 ;
        RECT 80.420 40.470 80.680 40.730 ;
        RECT 80.820 40.090 81.080 40.350 ;
        RECT 81.400 40.190 81.660 40.450 ;
        RECT 80.570 39.640 80.830 39.900 ;
        RECT 81.350 39.540 81.610 39.800 ;
        RECT 79.460 39.110 79.720 39.370 ;
        RECT 80.670 39.080 80.930 39.340 ;
        RECT 80.630 38.630 80.890 38.890 ;
        RECT 81.350 38.710 81.610 38.970 ;
        RECT 80.190 37.830 80.450 38.090 ;
        RECT 70.410 37.330 70.670 37.590 ;
        RECT 83.650 40.240 83.910 40.500 ;
        RECT 81.400 38.060 81.660 38.320 ;
        RECT 69.860 36.630 70.120 36.890 ;
        RECT 69.860 36.080 70.120 36.340 ;
        RECT 59.030 34.170 59.310 34.450 ;
        RECT 69.860 35.200 70.120 35.460 ;
        RECT 40.830 32.420 41.090 32.680 ;
        RECT 40.830 30.870 41.090 31.130 ;
        RECT 40.830 29.320 41.090 29.580 ;
        RECT 40.830 27.770 41.090 28.030 ;
        RECT 42.930 31.580 43.190 31.840 ;
        RECT 42.930 30.030 43.190 30.290 ;
        RECT 42.930 28.480 43.190 28.740 ;
        RECT 44.970 32.300 45.230 32.560 ;
        RECT 61.560 32.760 61.820 33.020 ;
        RECT 47.790 31.480 48.050 31.740 ;
        RECT 44.970 30.750 45.230 31.010 ;
        RECT 47.790 29.930 48.050 30.190 ;
        RECT 44.970 29.200 45.230 29.460 ;
        RECT 47.790 28.380 48.050 28.640 ;
        RECT 44.970 27.650 45.230 27.910 ;
        RECT 42.930 26.930 43.190 27.190 ;
        RECT 60.470 32.240 60.730 32.500 ;
        RECT 60.470 31.140 60.730 31.400 ;
        RECT 61.560 30.620 61.820 30.880 ;
        RECT 61.560 29.830 61.820 30.090 ;
        RECT 60.470 29.310 60.730 29.570 ;
        RECT 60.470 28.210 60.730 28.470 ;
        RECT 61.560 27.690 61.820 27.950 ;
        RECT 47.790 26.830 48.050 27.090 ;
        RECT 51.660 25.980 51.920 26.390 ;
        RECT 57.160 26.810 57.420 27.070 ;
        RECT 57.160 26.260 57.420 26.520 ;
        RECT 57.160 25.380 57.420 25.640 ;
        RECT 57.160 24.830 57.420 25.090 ;
        RECT 57.160 23.800 57.420 24.060 ;
        RECT 40.830 22.650 41.090 22.910 ;
        RECT 40.830 21.100 41.090 21.360 ;
        RECT 40.830 19.550 41.090 19.810 ;
        RECT 40.830 18.000 41.090 18.260 ;
        RECT 42.930 21.810 43.190 22.070 ;
        RECT 42.930 20.260 43.190 20.520 ;
        RECT 42.930 18.710 43.190 18.970 ;
        RECT 44.970 22.530 45.230 22.790 ;
        RECT 47.790 21.710 48.050 21.970 ;
        RECT 44.970 20.980 45.230 21.240 ;
        RECT 47.790 20.160 48.050 20.420 ;
        RECT 44.970 19.430 45.230 19.690 ;
        RECT 47.790 18.610 48.050 18.870 ;
        RECT 44.970 17.880 45.230 18.140 ;
        RECT 42.930 17.160 43.190 17.420 ;
        RECT 57.160 23.250 57.420 23.510 ;
        RECT 63.970 32.760 64.230 33.020 ;
        RECT 69.860 34.650 70.120 34.910 ;
        RECT 70.410 34.810 70.670 35.070 ;
        RECT 69.860 33.620 70.120 33.880 ;
        RECT 69.860 33.070 70.120 33.330 ;
        RECT 70.550 33.150 70.810 33.410 ;
        RECT 70.780 32.590 71.040 32.850 ;
        RECT 63.970 30.620 64.230 30.880 ;
        RECT 69.860 32.200 70.120 32.460 ;
        RECT 69.860 31.650 70.120 31.910 ;
        RECT 81.400 37.230 81.660 37.490 ;
        RECT 81.350 36.580 81.610 36.840 ;
        RECT 81.350 35.750 81.610 36.010 ;
        RECT 76.380 33.600 76.640 33.860 ;
        RECT 80.850 34.940 81.120 35.200 ;
        RECT 81.400 35.100 81.660 35.360 ;
        RECT 83.700 38.020 83.960 38.280 ;
        RECT 83.690 37.300 83.950 37.560 ;
        RECT 83.610 35.050 83.870 35.310 ;
        RECT 74.710 32.550 74.970 32.810 ;
        RECT 88.450 53.350 88.820 53.720 ;
        RECT 86.870 34.150 87.240 34.520 ;
        RECT 87.640 33.560 88.010 33.930 ;
        RECT 85.790 32.550 86.050 32.810 ;
        RECT 95.000 52.300 95.500 52.800 ;
        RECT 91.780 50.740 92.280 51.240 ;
        RECT 92.730 51.230 93.230 51.730 ;
        RECT 93.810 51.700 94.310 52.200 ;
        RECT 89.330 48.280 89.700 48.650 ;
        RECT 90.640 36.630 90.900 36.890 ;
        RECT 90.640 36.080 90.900 36.340 ;
        RECT 90.640 35.200 90.900 35.460 ;
        RECT 90.640 34.650 90.900 34.910 ;
        RECT 90.640 33.620 90.900 33.880 ;
        RECT 88.380 31.230 88.750 31.600 ;
        RECT 63.970 29.830 64.230 30.090 ;
        RECT 60.430 23.100 60.690 23.360 ;
        RECT 58.200 22.730 58.460 22.990 ;
        RECT 61.560 23.000 61.820 23.260 ;
        RECT 63.970 27.690 64.230 27.950 ;
        RECT 63.970 23.000 64.230 23.260 ;
        RECT 56.060 22.260 56.320 22.520 ;
        RECT 57.160 22.380 57.420 22.640 ;
        RECT 47.790 17.060 48.050 17.320 ;
        RECT 49.480 17.130 49.740 17.390 ;
        RECT 48.940 16.760 49.230 17.050 ;
        RECT 44.500 16.250 44.810 16.560 ;
        RECT 57.160 21.830 57.420 22.090 ;
        RECT 57.140 21.550 57.400 21.810 ;
        RECT 60.470 22.480 60.730 22.740 ;
        RECT 62.220 22.710 62.490 22.970 ;
        RECT 60.410 22.050 60.670 22.310 ;
        RECT 60.470 21.380 60.730 21.640 ;
        RECT 57.120 20.540 57.380 20.800 ;
        RECT 89.950 33.150 90.210 33.410 ;
        RECT 90.640 33.070 90.900 33.330 ;
        RECT 89.720 32.590 89.980 32.850 ;
        RECT 90.640 32.200 90.900 32.460 ;
        RECT 90.640 31.650 90.900 31.910 ;
        RECT 89.310 25.980 89.680 26.390 ;
        RECT 68.510 22.900 68.770 23.160 ;
        RECT 68.660 22.220 68.920 22.480 ;
        RECT 61.560 20.860 61.820 21.120 ;
        RECT 56.690 19.480 56.950 19.740 ;
        RECT 56.090 17.170 56.350 17.430 ;
        RECT 57.070 18.500 57.330 18.760 ;
        RECT 57.120 17.650 57.380 17.910 ;
        RECT 57.120 17.160 57.380 17.420 ;
        RECT 54.690 16.760 54.950 17.020 ;
        RECT 56.660 16.840 56.920 17.100 ;
        RECT 48.310 15.540 48.730 15.960 ;
        RECT 44.460 14.580 44.880 15.000 ;
        RECT 50.370 16.220 50.630 16.480 ;
        RECT 60.410 20.170 60.670 20.430 ;
        RECT 61.560 20.070 61.820 20.330 ;
        RECT 60.470 19.550 60.730 19.810 ;
        RECT 60.250 18.990 60.510 19.250 ;
        RECT 60.470 18.450 60.730 18.710 ;
        RECT 61.560 17.930 61.820 18.190 ;
        RECT 58.900 16.780 59.160 17.040 ;
        RECT 57.700 15.530 58.030 15.860 ;
        RECT 63.970 20.860 64.230 21.120 ;
        RECT 68.660 21.330 68.920 21.590 ;
        RECT 68.510 20.650 68.770 20.910 ;
        RECT 63.970 20.070 64.230 20.330 ;
        RECT 68.510 20.130 68.770 20.390 ;
        RECT 68.660 19.450 68.920 19.710 ;
        RECT 63.970 17.930 64.230 18.190 ;
        RECT 68.660 18.560 68.920 18.820 ;
        RECT 68.510 17.880 68.770 18.140 ;
        RECT 75.940 22.240 76.200 22.500 ;
        RECT 75.420 21.310 75.680 21.570 ;
        RECT 74.950 19.470 75.210 19.730 ;
        RECT 70.790 19.000 71.060 19.270 ;
        RECT 67.740 17.090 68.090 17.440 ;
        RECT 60.890 16.360 61.150 16.620 ;
        RECT 64.930 16.330 65.200 16.600 ;
        RECT 58.850 15.460 59.190 15.800 ;
        RECT 74.450 18.540 74.710 18.800 ;
        RECT 67.780 15.320 68.040 15.640 ;
        RECT 73.770 15.540 74.030 15.880 ;
        RECT 48.990 14.490 49.310 14.810 ;
        RECT 69.200 14.610 69.580 14.990 ;
        RECT 49.140 11.360 49.400 11.620 ;
        RECT 50.230 11.360 50.490 11.620 ;
        RECT 51.330 11.350 51.590 11.610 ;
        RECT 55.450 11.350 55.710 11.610 ;
        RECT 56.550 11.360 56.810 11.620 ;
        RECT 57.640 11.360 57.900 11.620 ;
        RECT 58.950 11.390 59.210 11.650 ;
        RECT 60.040 11.390 60.300 11.650 ;
        RECT 61.140 11.380 61.400 11.640 ;
        RECT 65.260 11.380 65.520 11.640 ;
        RECT 66.360 11.390 66.620 11.650 ;
        RECT 67.450 11.390 67.710 11.650 ;
        RECT 71.000 11.360 71.260 11.620 ;
        RECT 72.100 11.370 72.360 11.630 ;
        RECT 73.190 11.370 73.450 11.630 ;
        RECT 49.690 10.680 49.950 10.940 ;
        RECT 50.780 10.660 51.040 10.920 ;
        RECT 51.890 10.650 52.150 10.910 ;
        RECT 49.690 9.310 49.950 9.570 ;
        RECT 50.780 9.310 51.040 9.570 ;
        RECT 51.880 9.310 52.140 9.570 ;
        RECT 49.090 8.710 49.550 9.170 ;
        RECT 49.130 8.580 49.390 8.710 ;
        RECT 50.230 8.580 50.490 8.840 ;
        RECT 51.330 8.580 51.590 8.840 ;
        RECT 49.130 7.210 49.390 7.470 ;
        RECT 50.230 7.210 50.490 7.470 ;
        RECT 51.330 7.210 51.590 7.470 ;
        RECT 48.560 6.570 48.820 6.830 ;
        RECT 49.690 6.530 49.950 6.790 ;
        RECT 50.780 6.530 51.040 6.790 ;
        RECT 51.880 6.540 52.140 6.800 ;
        RECT 48.570 6.100 48.830 6.360 ;
        RECT 54.890 10.650 55.150 10.910 ;
        RECT 56.000 10.660 56.260 10.920 ;
        RECT 57.090 10.680 57.350 10.940 ;
        RECT 54.900 9.310 55.160 9.570 ;
        RECT 56.000 9.310 56.260 9.570 ;
        RECT 57.090 9.310 57.350 9.570 ;
        RECT 59.500 10.710 59.760 10.970 ;
        RECT 60.590 10.690 60.850 10.950 ;
        RECT 61.700 10.680 61.960 10.940 ;
        RECT 59.500 9.340 59.760 9.600 ;
        RECT 60.590 9.340 60.850 9.600 ;
        RECT 61.690 9.340 61.950 9.600 ;
        RECT 55.450 8.580 55.710 8.840 ;
        RECT 56.550 8.580 56.810 8.840 ;
        RECT 57.650 8.580 57.910 8.840 ;
        RECT 58.940 8.610 59.200 8.870 ;
        RECT 60.040 8.610 60.300 8.870 ;
        RECT 61.140 8.610 61.400 8.870 ;
        RECT 57.470 7.760 57.930 8.220 ;
        RECT 55.450 7.210 55.710 7.470 ;
        RECT 56.550 7.210 56.810 7.470 ;
        RECT 57.650 7.210 57.910 7.470 ;
        RECT 58.940 7.330 59.200 7.500 ;
        RECT 58.370 6.830 58.630 6.860 ;
        RECT 54.900 6.540 55.160 6.800 ;
        RECT 56.000 6.530 56.260 6.790 ;
        RECT 57.090 6.530 57.350 6.790 ;
        RECT 58.220 6.600 58.630 6.830 ;
        RECT 58.900 6.870 59.360 7.330 ;
        RECT 60.040 7.240 60.300 7.500 ;
        RECT 61.140 7.240 61.400 7.500 ;
        RECT 58.220 6.570 58.480 6.600 ;
        RECT 59.500 6.560 59.760 6.820 ;
        RECT 60.590 6.560 60.850 6.820 ;
        RECT 61.690 6.570 61.950 6.830 ;
        RECT 58.380 6.360 58.640 6.390 ;
        RECT 58.210 6.130 58.640 6.360 ;
        RECT 58.210 6.100 58.470 6.130 ;
        RECT 64.700 10.680 64.960 10.940 ;
        RECT 65.810 10.690 66.070 10.950 ;
        RECT 66.900 10.710 67.160 10.970 ;
        RECT 64.710 9.340 64.970 9.600 ;
        RECT 65.810 9.340 66.070 9.600 ;
        RECT 66.900 9.340 67.160 9.600 ;
        RECT 70.440 10.660 70.700 10.920 ;
        RECT 71.550 10.670 71.810 10.930 ;
        RECT 72.640 10.690 72.900 10.950 ;
        RECT 110.790 48.440 111.050 48.700 ;
        RECT 108.130 47.200 108.390 47.630 ;
        RECT 110.940 47.480 111.200 47.740 ;
        RECT 115.080 54.690 115.790 55.400 ;
        RECT 111.880 46.370 112.140 46.630 ;
        RECT 111.880 45.770 112.140 46.030 ;
        RECT 108.810 45.110 109.070 45.370 ;
        RECT 110.540 45.100 110.800 45.360 ;
        RECT 112.820 46.090 113.080 46.350 ;
        RECT 110.940 44.720 111.200 44.980 ;
        RECT 111.520 44.820 111.780 45.080 ;
        RECT 110.690 44.270 110.950 44.530 ;
        RECT 111.470 44.170 111.730 44.430 ;
        RECT 109.110 43.710 109.370 43.970 ;
        RECT 109.580 43.740 109.840 44.000 ;
        RECT 110.680 43.710 111.050 43.970 ;
        RECT 100.300 42.720 100.700 43.120 ;
        RECT 107.760 42.730 108.020 42.990 ;
        RECT 110.750 43.260 111.010 43.520 ;
        RECT 94.760 39.430 95.020 39.690 ;
        RECT 94.910 30.020 95.410 30.520 ;
        RECT 93.830 24.830 94.330 25.300 ;
        RECT 92.700 19.640 93.200 20.140 ;
        RECT 91.650 14.340 92.150 14.840 ;
        RECT 75.920 12.830 76.180 13.330 ;
        RECT 75.380 11.930 75.640 12.430 ;
        RECT 74.910 11.030 75.170 11.530 ;
        RECT 70.450 9.320 70.710 9.580 ;
        RECT 71.550 9.320 71.810 9.580 ;
        RECT 72.640 9.320 72.900 9.580 ;
        RECT 65.260 8.610 65.520 8.870 ;
        RECT 66.360 8.610 66.620 8.870 ;
        RECT 74.430 10.130 74.690 10.630 ;
        RECT 67.460 8.610 67.720 8.870 ;
        RECT 71.000 8.590 71.260 8.850 ;
        RECT 72.100 8.590 72.360 8.850 ;
        RECT 73.200 8.590 73.460 8.850 ;
        RECT 65.260 7.240 65.520 7.500 ;
        RECT 66.360 7.240 66.620 7.500 ;
        RECT 67.460 7.240 67.720 7.500 ;
        RECT 71.000 7.220 71.260 7.480 ;
        RECT 64.710 6.570 64.970 6.830 ;
        RECT 65.810 6.560 66.070 6.820 ;
        RECT 66.900 6.560 67.160 6.820 ;
        RECT 72.100 7.220 72.360 7.480 ;
        RECT 73.200 7.220 73.460 7.480 ;
        RECT 68.030 6.600 68.290 6.860 ;
        RECT 70.450 6.550 70.710 6.810 ;
        RECT 71.550 6.540 71.810 6.800 ;
        RECT 72.640 6.540 72.900 6.800 ;
        RECT 67.290 5.960 67.750 6.420 ;
        RECT 68.020 6.130 68.280 6.390 ;
        RECT 41.220 3.730 41.480 4.850 ;
        RECT 73.770 6.580 74.030 6.840 ;
        RECT 101.280 42.080 101.640 42.440 ;
        RECT 107.760 42.200 108.020 42.460 ;
        RECT 110.030 42.800 110.290 43.060 ;
        RECT 110.310 42.460 110.570 42.720 ;
        RECT 100.560 39.430 100.820 39.690 ;
        RECT 97.890 16.860 98.390 17.360 ;
        RECT 95.020 8.750 95.520 9.250 ;
        RECT 93.830 7.800 94.330 8.260 ;
        RECT 92.700 6.930 93.200 7.390 ;
        RECT 73.760 6.110 74.020 6.370 ;
        RECT 91.770 6.020 92.270 6.480 ;
        RECT 97.310 3.730 98.250 4.850 ;
        RECT 73.100 0.100 73.430 0.430 ;
        RECT 39.540 -0.560 39.870 -0.230 ;
        RECT 110.030 42.130 110.290 42.390 ;
        RECT 111.470 43.340 111.730 43.600 ;
        RECT 111.040 42.790 111.300 43.050 ;
        RECT 113.770 44.870 114.030 45.130 ;
        RECT 111.520 42.690 111.780 42.950 ;
        RECT 111.040 42.140 111.300 42.400 ;
        RECT 109.110 41.220 109.370 41.480 ;
        RECT 111.520 41.860 111.780 42.120 ;
        RECT 110.680 41.220 110.940 41.480 ;
        RECT 111.470 41.210 111.730 41.470 ;
        RECT 109.110 40.690 109.370 40.950 ;
        RECT 110.680 40.690 110.940 40.950 ;
        RECT 102.200 39.710 102.590 40.100 ;
        RECT 107.760 39.710 108.020 39.970 ;
        RECT 111.470 40.380 111.730 40.640 ;
        RECT 103.030 39.150 103.410 39.410 ;
        RECT 107.760 39.180 108.020 39.440 ;
        RECT 110.030 39.780 110.290 40.040 ;
        RECT 111.040 39.840 111.300 40.030 ;
        RECT 110.950 39.770 111.300 39.840 ;
        RECT 110.950 39.580 111.210 39.770 ;
        RECT 111.520 39.730 111.780 39.990 ;
        RECT 38.920 -1.180 39.250 -0.850 ;
        RECT 38.290 -1.810 38.620 -1.480 ;
        RECT 37.690 -2.440 38.020 -2.110 ;
        RECT 100.360 -1.090 100.760 -0.690 ;
        RECT 99.880 -2.020 100.140 -1.760 ;
        RECT 101.270 -1.890 101.660 -1.500 ;
        RECT 37.050 -3.120 37.380 -2.790 ;
        RECT 36.450 -3.740 36.780 -3.410 ;
        RECT 102.200 -2.710 102.590 -2.320 ;
        RECT 110.030 39.110 110.290 39.370 ;
        RECT 111.040 39.120 111.300 39.380 ;
        RECT 113.820 42.650 114.080 42.910 ;
        RECT 113.810 41.930 114.070 42.190 ;
        RECT 113.730 39.680 113.990 39.940 ;
        RECT 109.110 38.200 109.370 38.460 ;
        RECT 110.680 38.200 110.940 38.460 ;
        RECT 114.890 34.900 115.600 35.610 ;
        RECT 110.690 16.850 111.200 17.360 ;
        RECT 104.660 3.220 104.920 3.480 ;
        RECT 104.660 2.550 104.920 2.810 ;
        RECT 104.780 1.310 105.040 1.570 ;
        RECT 104.780 -0.300 105.040 -0.040 ;
        RECT 104.770 -1.910 105.030 -1.650 ;
        RECT 103.020 -3.500 103.400 -3.120 ;
        RECT 104.770 -3.530 105.030 -3.270 ;
        RECT 35.850 -4.380 36.180 -4.050 ;
        RECT 35.270 -4.950 35.600 -4.620 ;
        RECT 34.690 -5.640 35.020 -5.310 ;
        RECT 104.770 -5.140 105.030 -4.880 ;
        RECT 34.040 -6.280 34.370 -5.950 ;
        RECT 33.400 -6.930 33.730 -6.590 ;
        RECT 104.400 -6.740 104.660 -6.480 ;
        RECT 32.820 -7.570 33.190 -7.200 ;
        RECT 104.780 -8.340 105.040 -8.080 ;
        RECT 101.570 -10.010 101.830 -9.750 ;
        RECT 102.510 -10.010 102.770 -9.750 ;
        RECT 103.460 -10.070 103.720 -9.810 ;
        RECT 104.770 -9.930 105.030 -9.670 ;
      LAYER met2 ;
        RECT 9.460 61.490 9.780 61.540 ;
        RECT 6.600 61.250 9.780 61.490 ;
        RECT 6.600 61.230 6.920 61.250 ;
        RECT 49.160 50.370 49.270 50.570 ;
        RECT 47.760 50.170 48.080 50.220 ;
        RECT 40.470 49.390 40.560 49.710 ;
        RECT 42.930 49.350 43.190 50.150 ;
        RECT 47.760 49.970 49.390 50.170 ;
        RECT 47.760 49.960 48.080 49.970 ;
        RECT 77.970 49.560 78.280 49.620 ;
        RECT 49.670 49.550 78.280 49.560 ;
        RECT 44.930 49.350 45.270 49.410 ;
        RECT 49.340 49.360 78.280 49.550 ;
        RECT 49.340 49.350 49.920 49.360 ;
        RECT 40.660 48.990 41.120 49.310 ;
        RECT 42.830 49.130 45.270 49.350 ;
        RECT 77.970 49.300 78.280 49.360 ;
        RECT 56.900 49.090 57.220 49.140 ;
        RECT 49.160 48.820 49.270 49.020 ;
        RECT 51.900 48.890 57.270 49.090 ;
        RECT 47.760 48.620 48.080 48.670 ;
        RECT 40.470 47.840 40.560 48.160 ;
        RECT 42.930 47.800 43.190 48.600 ;
        RECT 47.760 48.420 49.390 48.620 ;
        RECT 47.760 48.410 48.080 48.420 ;
        RECT 51.900 48.010 52.100 48.890 ;
        RECT 56.900 48.880 57.220 48.890 ;
        RECT 59.660 48.650 59.970 48.660 ;
        RECT 59.660 48.620 59.980 48.650 ;
        RECT 49.660 48.000 52.100 48.010 ;
        RECT 44.930 47.800 45.270 47.860 ;
        RECT 49.370 47.810 52.100 48.000 ;
        RECT 52.410 48.420 59.980 48.620 ;
        RECT 49.370 47.800 49.860 47.810 ;
        RECT 40.660 47.440 41.120 47.760 ;
        RECT 42.830 47.580 45.270 47.800 ;
        RECT 49.160 47.270 49.270 47.470 ;
        RECT 47.760 47.070 48.080 47.120 ;
        RECT 40.470 46.290 40.560 46.610 ;
        RECT 42.930 46.250 43.190 47.050 ;
        RECT 47.760 46.870 49.390 47.070 ;
        RECT 47.760 46.860 48.080 46.870 ;
        RECT 52.410 46.460 52.610 48.420 ;
        RECT 59.660 48.390 59.980 48.420 ;
        RECT 59.660 48.380 59.970 48.390 ;
        RECT 60.720 48.140 61.040 48.180 ;
        RECT 49.660 46.450 52.610 46.460 ;
        RECT 44.930 46.250 45.270 46.310 ;
        RECT 49.370 46.260 52.610 46.450 ;
        RECT 52.960 47.940 61.120 48.140 ;
        RECT 49.370 46.250 49.870 46.260 ;
        RECT 40.660 45.890 41.120 46.210 ;
        RECT 42.830 46.030 45.270 46.250 ;
        RECT 49.160 45.720 49.270 45.920 ;
        RECT 47.760 45.520 48.080 45.570 ;
        RECT 40.470 44.740 40.560 45.060 ;
        RECT 42.930 44.700 43.190 45.500 ;
        RECT 47.760 45.320 49.390 45.520 ;
        RECT 47.760 45.310 48.080 45.320 ;
        RECT 52.960 44.910 53.160 47.940 ;
        RECT 60.720 47.900 61.040 47.940 ;
        RECT 49.670 44.900 53.160 44.910 ;
        RECT 44.930 44.700 45.270 44.760 ;
        RECT 49.370 44.710 53.160 44.900 ;
        RECT 86.310 44.730 86.390 44.910 ;
        RECT 49.370 44.700 49.830 44.710 ;
        RECT 40.660 44.340 41.120 44.660 ;
        RECT 42.830 44.480 45.270 44.700 ;
        RECT 80.460 44.100 81.060 44.270 ;
        RECT 84.060 44.100 89.290 44.330 ;
        RECT 71.590 43.920 83.120 44.100 ;
        RECT 80.460 43.710 81.060 43.920 ;
        RECT 84.530 43.860 84.840 44.000 ;
        RECT 82.360 43.850 84.840 43.860 ;
        RECT 82.360 43.700 93.880 43.850 ;
        RECT 82.360 43.680 84.840 43.700 ;
        RECT 84.530 43.670 84.840 43.680 ;
        RECT 61.510 43.510 61.820 43.560 ;
        RECT 61.510 43.500 61.970 43.510 ;
        RECT 61.510 43.320 63.760 43.500 ;
        RECT 61.510 43.230 61.820 43.320 ;
        RECT 84.070 43.280 89.290 43.500 ;
        RECT 80.790 43.080 81.100 43.150 ;
        RECT 80.790 42.860 83.120 43.080 ;
        RECT 40.660 42.520 41.120 42.840 ;
        RECT 80.790 42.820 81.100 42.860 ;
        RECT 42.830 42.480 45.270 42.700 ;
        RECT 49.670 42.490 49.970 42.520 ;
        RECT 49.670 42.480 50.060 42.490 ;
        RECT 40.470 42.120 40.560 42.440 ;
        RECT 42.930 41.680 43.190 42.480 ;
        RECT 44.930 42.420 45.270 42.480 ;
        RECT 49.370 42.280 50.060 42.480 ;
        RECT 60.290 42.360 60.770 42.590 ;
        RECT 60.430 42.290 60.770 42.360 ;
        RECT 53.300 41.880 63.760 42.100 ;
        RECT 47.760 41.860 48.080 41.870 ;
        RECT 47.760 41.660 49.390 41.860 ;
        RECT 53.300 41.740 53.620 41.880 ;
        RECT 47.760 41.610 48.080 41.660 ;
        RECT 40.660 40.970 41.120 41.290 ;
        RECT 49.160 41.260 49.270 41.460 ;
        RECT 53.320 41.400 53.580 41.740 ;
        RECT 49.640 41.170 49.970 41.370 ;
        RECT 42.830 40.930 45.270 41.150 ;
        RECT 49.640 40.950 49.820 41.170 ;
        RECT 53.300 41.140 53.620 41.400 ;
        RECT 55.670 41.250 56.400 41.430 ;
        RECT 60.430 41.420 60.770 41.490 ;
        RECT 55.670 41.040 55.850 41.250 ;
        RECT 60.290 41.190 60.770 41.420 ;
        RECT 49.620 40.930 49.820 40.950 ;
        RECT 40.470 40.570 40.560 40.890 ;
        RECT 42.930 40.130 43.190 40.930 ;
        RECT 44.930 40.870 45.270 40.930 ;
        RECT 49.370 40.730 49.820 40.930 ;
        RECT 55.280 40.860 55.850 41.040 ;
        RECT 84.840 40.820 89.290 40.980 ;
        RECT 84.810 40.780 89.290 40.820 ;
        RECT 56.440 40.610 56.760 40.730 ;
        RECT 78.640 40.610 78.960 40.730 ;
        RECT 56.440 40.430 78.960 40.610 ;
        RECT 54.250 40.320 54.560 40.390 ;
        RECT 47.760 40.310 48.080 40.320 ;
        RECT 47.760 40.110 49.390 40.310 ;
        RECT 52.230 40.140 63.760 40.320 ;
        RECT 63.940 40.140 64.260 40.160 ;
        RECT 52.230 40.110 64.260 40.140 ;
        RECT 47.760 40.060 48.080 40.110 ;
        RECT 53.540 40.100 64.260 40.110 ;
        RECT 54.250 40.060 54.560 40.100 ;
        RECT 40.660 39.420 41.120 39.740 ;
        RECT 49.160 39.710 49.270 39.910 ;
        RECT 55.770 39.890 55.950 40.100 ;
        RECT 55.280 39.710 55.950 39.890 ;
        RECT 61.530 39.950 64.260 40.100 ;
        RECT 61.530 39.870 61.850 39.950 ;
        RECT 63.940 39.940 64.260 39.950 ;
        RECT 63.940 39.900 65.960 39.940 ;
        RECT 61.540 39.790 61.850 39.870 ;
        RECT 42.830 39.380 45.270 39.600 ;
        RECT 49.620 39.540 49.970 39.610 ;
        RECT 49.620 39.380 50.010 39.540 ;
        RECT 60.290 39.430 60.770 39.660 ;
        RECT 61.540 39.580 63.760 39.790 ;
        RECT 64.050 39.780 65.960 39.900 ;
        RECT 64.770 39.760 65.960 39.780 ;
        RECT 61.540 39.540 61.850 39.580 ;
        RECT 65.100 39.500 65.940 39.700 ;
        RECT 40.470 39.020 40.560 39.340 ;
        RECT 42.930 38.580 43.190 39.380 ;
        RECT 44.930 39.320 45.270 39.380 ;
        RECT 49.430 39.310 50.010 39.380 ;
        RECT 49.430 39.180 49.820 39.310 ;
        RECT 54.400 39.230 54.710 39.370 ;
        RECT 60.430 39.360 60.770 39.430 ;
        RECT 52.230 39.220 54.710 39.230 ;
        RECT 52.230 39.070 63.760 39.220 ;
        RECT 52.230 39.050 54.710 39.070 ;
        RECT 54.400 39.040 54.710 39.050 ;
        RECT 47.760 38.760 48.080 38.770 ;
        RECT 47.760 38.560 49.390 38.760 ;
        RECT 47.760 38.510 48.080 38.560 ;
        RECT 60.430 38.490 60.770 38.560 ;
        RECT 40.660 37.870 41.120 38.190 ;
        RECT 49.160 38.160 49.270 38.360 ;
        RECT 49.710 38.230 49.970 38.440 ;
        RECT 60.290 38.260 60.770 38.490 ;
        RECT 81.370 38.300 81.680 38.350 ;
        RECT 83.670 38.300 83.980 38.320 ;
        RECT 84.810 38.300 85.040 40.780 ;
        RECT 86.310 39.860 86.390 40.040 ;
        RECT 109.080 38.380 109.390 38.500 ;
        RECT 108.310 38.370 109.430 38.380 ;
        RECT 110.650 38.370 110.960 38.500 ;
        RECT 42.830 37.830 45.270 38.050 ;
        RECT 49.710 37.830 49.910 38.230 ;
        RECT 65.500 38.080 74.510 38.280 ;
        RECT 80.440 38.120 81.060 38.220 ;
        RECT 80.160 38.080 81.060 38.120 ;
        RECT 64.710 38.070 74.510 38.080 ;
        RECT 64.020 38.060 74.510 38.070 ;
        RECT 55.280 37.850 56.050 38.030 ;
        RECT 40.470 37.470 40.560 37.790 ;
        RECT 42.930 37.030 43.190 37.830 ;
        RECT 44.930 37.770 45.270 37.830 ;
        RECT 49.570 37.630 49.910 37.830 ;
        RECT 49.710 37.620 49.910 37.630 ;
        RECT 47.760 37.210 48.080 37.220 ;
        RECT 47.760 37.010 49.390 37.210 ;
        RECT 47.760 36.960 48.080 37.010 ;
        RECT 49.160 36.610 49.270 36.810 ;
        RECT 55.870 35.410 56.050 37.850 ;
        RECT 61.530 37.970 61.850 38.050 ;
        RECT 64.020 38.020 65.960 38.060 ;
        RECT 63.940 37.970 65.960 38.020 ;
        RECT 61.530 37.910 65.960 37.970 ;
        RECT 61.530 37.780 64.260 37.910 ;
        RECT 64.710 37.900 65.960 37.910 ;
        RECT 61.530 37.730 61.850 37.780 ;
        RECT 63.940 37.760 64.260 37.780 ;
        RECT 64.680 37.620 65.000 37.670 ;
        RECT 64.680 37.370 70.700 37.620 ;
        RECT 70.380 37.300 70.700 37.370 ;
        RECT 69.840 36.790 70.150 36.930 ;
        RECT 74.290 36.790 74.510 38.060 ;
        RECT 79.840 37.840 81.060 38.080 ;
        RECT 81.370 38.070 85.040 38.300 ;
        RECT 85.650 38.170 89.290 38.370 ;
        RECT 89.660 38.170 110.960 38.370 ;
        RECT 81.370 38.020 81.680 38.070 ;
        RECT 83.670 37.990 83.980 38.070 ;
        RECT 80.160 37.790 81.060 37.840 ;
        RECT 80.440 37.690 81.060 37.790 ;
        RECT 81.370 37.470 81.680 37.530 ;
        RECT 83.660 37.470 83.970 37.600 ;
        RECT 85.650 37.470 85.850 38.170 ;
        RECT 108.310 38.160 109.430 38.170 ;
        RECT 81.370 37.320 85.850 37.470 ;
        RECT 81.370 37.250 85.820 37.320 ;
        RECT 81.370 37.200 81.680 37.250 ;
        RECT 90.610 36.790 90.920 36.930 ;
        RECT 67.680 36.610 77.750 36.790 ;
        RECT 83.010 36.610 93.080 36.790 ;
        RECT 69.840 36.600 70.150 36.610 ;
        RECT 65.550 36.360 71.210 36.500 ;
        RECT 74.290 36.450 74.510 36.610 ;
        RECT 90.610 36.600 90.920 36.610 ;
        RECT 74.290 36.360 77.140 36.450 ;
        RECT 90.610 36.360 90.920 36.380 ;
        RECT 65.550 36.280 77.750 36.360 ;
        RECT 67.680 36.180 77.750 36.280 ;
        RECT 83.010 36.180 93.080 36.360 ;
        RECT 69.840 36.050 70.150 36.180 ;
        RECT 65.050 35.980 65.530 35.990 ;
        RECT 65.050 35.740 65.940 35.980 ;
        RECT 70.990 35.950 71.210 36.180 ;
        RECT 90.610 36.050 90.920 36.180 ;
        RECT 81.320 36.000 81.630 36.040 ;
        RECT 75.360 35.950 81.630 36.000 ;
        RECT 70.990 35.790 81.630 35.950 ;
        RECT 70.990 35.730 75.750 35.790 ;
        RECT 81.320 35.710 81.630 35.790 ;
        RECT 55.870 35.230 56.410 35.410 ;
        RECT 69.840 35.360 70.150 35.490 ;
        RECT 67.680 35.180 77.760 35.360 ;
        RECT 81.370 35.310 81.680 35.390 ;
        RECT 90.610 35.360 90.920 35.490 ;
        RECT 83.000 35.310 93.080 35.360 ;
        RECT 81.370 35.180 93.080 35.310 ;
        RECT 69.840 35.160 70.150 35.180 ;
        RECT 81.370 35.080 84.080 35.180 ;
        RECT 90.610 35.160 90.920 35.180 ;
        RECT 81.370 35.060 81.680 35.080 ;
        RECT 83.580 35.020 83.890 35.080 ;
        RECT 90.610 34.930 90.920 34.940 ;
        RECT 83.000 34.750 93.080 34.930 ;
        RECT 90.610 34.610 90.920 34.750 ;
        RECT 61.530 33.000 61.850 33.050 ;
        RECT 63.940 33.000 64.260 33.020 ;
        RECT 56.040 32.810 57.820 32.930 ;
        RECT 55.450 32.750 57.820 32.810 ;
        RECT 61.530 32.860 64.260 33.000 ;
        RECT 61.530 32.810 65.960 32.860 ;
        RECT 40.660 32.390 41.120 32.710 ;
        RECT 55.450 32.630 56.290 32.750 ;
        RECT 61.530 32.730 61.850 32.810 ;
        RECT 63.940 32.760 65.960 32.810 ;
        RECT 70.320 32.790 70.460 32.980 ;
        RECT 90.350 32.790 90.440 32.970 ;
        RECT 63.980 32.690 65.960 32.760 ;
        RECT 65.440 32.680 65.960 32.690 ;
        RECT 42.830 32.350 45.270 32.570 ;
        RECT 49.710 32.450 49.960 32.470 ;
        RECT 49.710 32.350 49.970 32.450 ;
        RECT 40.470 31.990 40.560 32.310 ;
        RECT 42.930 31.550 43.190 32.350 ;
        RECT 44.930 32.290 45.270 32.350 ;
        RECT 49.370 32.150 49.970 32.350 ;
        RECT 60.290 32.290 60.770 32.520 ;
        RECT 69.840 32.370 70.150 32.490 ;
        RECT 70.320 32.370 70.460 32.550 ;
        RECT 77.580 32.370 78.140 32.500 ;
        RECT 90.350 32.370 90.440 32.540 ;
        RECT 90.610 32.370 90.920 32.490 ;
        RECT 69.840 32.360 78.140 32.370 ;
        RECT 60.430 32.220 60.770 32.290 ;
        RECT 67.680 32.320 78.140 32.360 ;
        RECT 83.020 32.360 90.920 32.370 ;
        RECT 67.680 32.200 77.740 32.320 ;
        RECT 83.020 32.200 93.080 32.360 ;
        RECT 67.680 32.180 70.240 32.200 ;
        RECT 69.840 32.160 70.150 32.180 ;
        RECT 75.420 32.110 76.960 32.200 ;
        RECT 83.800 32.110 85.340 32.200 ;
        RECT 90.520 32.180 93.080 32.200 ;
        RECT 90.610 32.160 90.920 32.180 ;
        RECT 69.840 31.930 70.150 31.940 ;
        RECT 90.610 31.930 90.920 31.940 ;
        RECT 67.680 31.760 77.740 31.930 ;
        RECT 83.020 31.760 93.080 31.930 ;
        RECT 67.680 31.750 70.150 31.760 ;
        RECT 47.760 31.730 48.080 31.740 ;
        RECT 47.760 31.530 49.390 31.730 ;
        RECT 69.840 31.610 70.150 31.750 ;
        RECT 90.610 31.750 93.080 31.760 ;
        RECT 90.610 31.610 90.920 31.750 ;
        RECT 47.760 31.480 48.080 31.530 ;
        RECT 60.430 31.350 60.770 31.420 ;
        RECT 70.320 31.360 70.470 31.550 ;
        RECT 90.320 31.360 90.450 31.540 ;
        RECT 40.660 30.840 41.120 31.160 ;
        RECT 49.160 31.130 49.270 31.330 ;
        RECT 49.560 31.100 49.940 31.300 ;
        RECT 60.290 31.120 60.770 31.350 ;
        RECT 49.560 31.070 49.930 31.100 ;
        RECT 42.830 30.800 45.270 31.020 ;
        RECT 49.560 30.800 49.760 31.070 ;
        RECT 56.060 30.970 57.820 31.070 ;
        RECT 40.470 30.440 40.560 30.760 ;
        RECT 42.930 30.000 43.190 30.800 ;
        RECT 44.930 30.740 45.270 30.800 ;
        RECT 49.370 30.600 49.760 30.800 ;
        RECT 55.460 30.890 57.820 30.970 ;
        RECT 55.460 30.790 56.340 30.890 ;
        RECT 61.530 30.830 61.850 30.910 ;
        RECT 64.010 30.880 65.960 31.020 ;
        RECT 70.320 30.930 70.450 31.110 ;
        RECT 90.310 30.930 90.450 31.110 ;
        RECT 63.940 30.860 65.960 30.880 ;
        RECT 63.940 30.830 64.260 30.860 ;
        RECT 64.740 30.850 65.960 30.860 ;
        RECT 65.440 30.840 65.960 30.850 ;
        RECT 61.530 30.640 64.260 30.830 ;
        RECT 61.530 30.590 61.850 30.640 ;
        RECT 63.940 30.620 64.260 30.640 ;
        RECT 47.760 30.180 48.080 30.190 ;
        RECT 47.760 29.980 49.390 30.180 ;
        RECT 61.530 30.070 61.850 30.120 ;
        RECT 63.940 30.070 64.260 30.090 ;
        RECT 47.760 29.930 48.080 29.980 ;
        RECT 56.070 29.820 57.820 29.920 ;
        RECT 40.660 29.290 41.120 29.610 ;
        RECT 49.160 29.580 49.270 29.780 ;
        RECT 55.460 29.740 57.820 29.820 ;
        RECT 61.530 29.880 64.260 30.070 ;
        RECT 61.530 29.800 61.850 29.880 ;
        RECT 63.940 29.870 64.260 29.880 ;
        RECT 63.940 29.830 65.960 29.870 ;
        RECT 55.460 29.640 56.340 29.740 ;
        RECT 64.050 29.710 65.960 29.830 ;
        RECT 70.320 29.780 70.390 29.960 ;
        RECT 90.360 29.780 90.450 29.960 ;
        RECT 64.770 29.690 65.960 29.710 ;
        RECT 42.830 29.250 45.270 29.470 ;
        RECT 49.770 29.250 49.970 29.530 ;
        RECT 60.290 29.360 60.770 29.590 ;
        RECT 60.430 29.290 60.770 29.360 ;
        RECT 70.320 29.350 70.390 29.530 ;
        RECT 90.360 29.350 90.450 29.530 ;
        RECT 40.470 28.890 40.560 29.210 ;
        RECT 42.930 28.450 43.190 29.250 ;
        RECT 44.930 29.190 45.270 29.250 ;
        RECT 49.370 29.050 49.970 29.250 ;
        RECT 77.020 28.800 83.780 28.980 ;
        RECT 47.760 28.630 48.080 28.640 ;
        RECT 47.760 28.430 49.390 28.630 ;
        RECT 47.760 28.380 48.080 28.430 ;
        RECT 60.430 28.420 60.770 28.490 ;
        RECT 40.660 27.740 41.120 28.060 ;
        RECT 49.160 28.030 49.270 28.230 ;
        RECT 42.830 27.700 45.270 27.920 ;
        RECT 49.770 27.700 49.970 28.370 ;
        RECT 60.290 28.190 60.770 28.420 ;
        RECT 70.320 28.360 70.390 28.540 ;
        RECT 90.360 28.360 90.450 28.540 ;
        RECT 56.040 27.960 57.820 28.070 ;
        RECT 64.710 28.000 65.960 28.010 ;
        RECT 55.460 27.890 57.820 27.960 ;
        RECT 61.530 27.900 61.850 27.980 ;
        RECT 64.020 27.950 65.960 28.000 ;
        RECT 63.940 27.900 65.960 27.950 ;
        RECT 70.320 27.930 70.390 28.110 ;
        RECT 90.360 27.930 90.450 28.110 ;
        RECT 55.460 27.780 56.340 27.890 ;
        RECT 61.530 27.840 65.960 27.900 ;
        RECT 40.470 27.340 40.560 27.660 ;
        RECT 42.930 26.900 43.190 27.700 ;
        RECT 44.930 27.640 45.270 27.700 ;
        RECT 49.370 27.500 49.970 27.700 ;
        RECT 61.530 27.710 64.260 27.840 ;
        RECT 64.710 27.830 65.960 27.840 ;
        RECT 61.530 27.660 61.850 27.710 ;
        RECT 63.940 27.690 64.260 27.710 ;
        RECT 47.760 27.080 48.080 27.090 ;
        RECT 47.760 26.880 49.390 27.080 ;
        RECT 57.140 26.970 57.450 27.110 ;
        RECT 47.760 26.830 48.080 26.880 ;
        RECT 54.980 26.790 57.550 26.970 ;
        RECT 57.140 26.780 57.450 26.790 ;
        RECT 49.160 26.480 49.270 26.680 ;
        RECT 57.140 23.960 57.450 24.100 ;
        RECT 54.970 23.950 57.450 23.960 ;
        RECT 54.970 23.780 57.570 23.950 ;
        RECT 57.140 23.770 57.450 23.780 ;
        RECT 55.310 22.970 57.640 23.150 ;
        RECT 58.170 22.940 58.490 23.000 ;
        RECT 62.190 22.940 62.520 22.970 ;
        RECT 40.660 22.620 41.120 22.940 ;
        RECT 42.830 22.580 45.270 22.800 ;
        RECT 58.170 22.770 62.520 22.940 ;
        RECT 58.170 22.720 58.490 22.770 ;
        RECT 62.190 22.710 62.520 22.770 ;
        RECT 40.470 22.220 40.560 22.540 ;
        RECT 42.930 21.780 43.190 22.580 ;
        RECT 44.930 22.520 45.270 22.580 ;
        RECT 49.350 22.380 50.000 22.580 ;
        RECT 47.760 21.960 48.080 21.970 ;
        RECT 47.760 21.760 49.390 21.960 ;
        RECT 47.760 21.710 48.080 21.760 ;
        RECT 40.660 21.070 41.120 21.390 ;
        RECT 49.160 21.360 49.270 21.560 ;
        RECT 49.730 21.330 49.980 21.560 ;
        RECT 42.830 21.030 45.270 21.250 ;
        RECT 49.730 21.030 49.930 21.330 ;
        RECT 40.470 20.670 40.560 20.990 ;
        RECT 42.930 20.230 43.190 21.030 ;
        RECT 44.930 20.970 45.270 21.030 ;
        RECT 49.370 20.830 49.930 21.030 ;
        RECT 55.310 21.110 57.650 21.290 ;
        RECT 55.310 21.010 55.490 21.110 ;
        RECT 47.760 20.410 48.080 20.420 ;
        RECT 47.760 20.210 49.390 20.410 ;
        RECT 47.760 20.160 48.080 20.210 ;
        RECT 40.660 19.520 41.120 19.840 ;
        RECT 49.160 19.810 49.270 20.010 ;
        RECT 55.320 19.960 57.640 20.140 ;
        RECT 57.090 19.950 57.250 19.960 ;
        RECT 49.740 19.770 49.940 19.780 ;
        RECT 42.830 19.480 45.270 19.700 ;
        RECT 49.740 19.500 50.030 19.770 ;
        RECT 49.740 19.480 49.940 19.500 ;
        RECT 40.470 19.120 40.560 19.440 ;
        RECT 42.930 18.680 43.190 19.480 ;
        RECT 44.930 19.420 45.270 19.480 ;
        RECT 49.330 19.280 49.940 19.480 ;
        RECT 70.760 19.190 71.090 19.280 ;
        RECT 64.410 19.020 71.090 19.190 ;
        RECT 70.760 18.990 71.090 19.020 ;
        RECT 47.760 18.860 48.080 18.870 ;
        RECT 47.760 18.660 49.390 18.860 ;
        RECT 47.760 18.610 48.080 18.660 ;
        RECT 49.720 18.620 50.020 18.660 ;
        RECT 19.470 18.030 20.080 18.360 ;
        RECT 19.480 17.540 20.080 18.030 ;
        RECT 40.660 17.970 41.120 18.290 ;
        RECT 49.160 18.260 49.270 18.460 ;
        RECT 49.710 18.380 50.020 18.620 ;
        RECT 57.040 18.470 57.350 18.800 ;
        RECT 60.430 18.660 60.770 18.730 ;
        RECT 60.290 18.430 60.770 18.660 ;
        RECT 42.830 17.930 45.270 18.150 ;
        RECT 49.710 17.930 49.910 18.380 ;
        RECT 57.110 18.290 57.270 18.300 ;
        RECT 55.320 18.110 57.640 18.290 ;
        RECT 64.710 18.240 65.960 18.250 ;
        RECT 61.530 18.140 61.850 18.220 ;
        RECT 64.020 18.190 65.960 18.240 ;
        RECT 63.940 18.140 65.960 18.190 ;
        RECT 61.530 18.110 65.960 18.140 ;
        RECT 68.480 18.120 68.790 18.180 ;
        RECT 67.930 18.110 68.790 18.120 ;
        RECT 40.470 17.570 40.560 17.890 ;
        RECT 42.930 17.130 43.190 17.930 ;
        RECT 44.930 17.870 45.270 17.930 ;
        RECT 49.360 17.730 49.910 17.930 ;
        RECT 57.090 17.830 57.400 17.950 ;
        RECT 60.350 17.890 68.790 18.110 ;
        RECT 60.350 17.880 67.940 17.890 ;
        RECT 60.350 17.870 61.120 17.880 ;
        RECT 60.350 17.830 60.590 17.870 ;
        RECT 68.480 17.850 68.790 17.890 ;
        RECT 57.090 17.630 60.590 17.830 ;
        RECT 57.090 17.620 59.780 17.630 ;
        RECT 57.090 17.340 57.410 17.430 ;
        RECT 67.710 17.340 68.120 17.450 ;
        RECT 47.760 17.310 48.080 17.320 ;
        RECT 47.760 17.110 49.390 17.310 ;
        RECT 57.090 17.180 68.120 17.340 ;
        RECT 57.090 17.150 57.410 17.180 ;
        RECT 47.760 17.060 48.080 17.110 ;
        RECT 67.710 17.080 68.120 17.180 ;
        RECT 73.750 15.880 74.050 15.900 ;
        RECT 67.410 15.300 68.070 15.660 ;
        RECT 73.040 15.540 74.060 15.880 ;
        RECT 73.750 15.520 74.060 15.540 ;
        RECT 69.160 14.580 69.610 15.010 ;
        RECT 117.910 10.800 117.920 10.810 ;
        RECT 19.510 10.470 20.120 10.800 ;
        RECT 19.520 9.980 20.120 10.470 ;
        RECT 48.240 6.400 48.840 6.890 ;
        RECT 48.240 6.070 48.850 6.400 ;
        RECT 104.800 3.500 105.090 3.560 ;
        RECT 104.630 3.190 105.090 3.500 ;
        RECT 104.800 3.150 105.090 3.190 ;
        RECT 104.810 2.830 105.090 3.150 ;
        RECT 104.630 2.520 105.090 2.830 ;
        RECT 104.810 2.400 105.090 2.520 ;
        RECT 2.770 -2.960 4.040 -1.080 ;
        RECT 2.840 -7.710 4.110 -5.830 ;
        RECT 101.540 -10.040 101.860 -9.720 ;
        RECT 102.480 -10.040 102.800 -9.720 ;
      LAYER via2 ;
        RECT 80.590 43.820 80.930 44.160 ;
        RECT 80.610 37.770 80.950 38.130 ;
  END
END sky130_hilas_TopLevelTextStructure

MACRO sky130_hilas_pFETLarge
  CLASS CORE ;
  FOREIGN sky130_hilas_pFETLarge ;
  ORIGIN 0.750 0.000 ;
  SIZE 5.390 BY 6.100 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA 5.457400 ;
    ANTENNADIFFAREA 1.079500 ;
    PORT
      LAYER met2 ;
        RECT 0.000 0.340 0.600 0.830 ;
        RECT 0.000 0.010 0.610 0.340 ;
    END
  END GATE
  PIN SOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 2.724600 ;
    PORT
      LAYER met2 ;
        RECT 0.330 5.600 3.390 5.610 ;
        RECT 0.240 5.270 3.390 5.600 ;
        RECT 0.240 2.820 0.560 5.270 ;
        RECT 3.060 5.260 3.370 5.270 ;
        RECT 0.240 2.490 3.400 2.820 ;
        RECT 0.240 1.450 0.560 2.490 ;
        RECT 0.240 1.130 3.400 1.450 ;
        RECT 0.860 1.120 1.170 1.130 ;
        RECT 1.960 1.120 2.270 1.130 ;
        RECT 3.060 1.120 3.370 1.130 ;
    END
  END SOURCE
  PIN DRAIN
    USE ANALOG ;
    ANTENNADIFFAREA 1.386200 ;
    PORT
      LAYER met2 ;
        RECT 1.420 4.890 1.730 4.920 ;
        RECT 2.510 4.890 2.820 4.900 ;
        RECT 1.420 4.590 4.370 4.890 ;
        RECT 2.510 4.570 2.820 4.590 ;
        RECT 3.620 4.550 4.370 4.590 ;
        RECT 3.990 4.420 4.370 4.550 ;
        RECT 4.020 3.550 4.370 4.420 ;
        RECT 1.420 3.220 4.370 3.550 ;
        RECT 4.020 0.780 4.370 3.220 ;
        RECT 1.430 0.770 4.370 0.780 ;
        RECT 1.420 0.460 4.370 0.770 ;
        RECT 1.420 0.450 4.140 0.460 ;
        RECT 1.420 0.440 1.730 0.450 ;
        RECT 2.510 0.440 2.820 0.450 ;
    END
  END DRAIN
  PIN WELL
    USE ANALOG ;
    ANTENNADIFFAREA 0.213200 ;
    PORT
      LAYER nwell ;
        RECT 4.020 0.180 4.640 5.880 ;
      LAYER met1 ;
        RECT 4.140 5.790 4.400 5.990 ;
        RECT 4.140 4.980 4.450 5.790 ;
        RECT 4.140 0.000 4.400 4.980 ;
    END
  END WELL
  OBS
      LAYER nwell ;
        RECT -0.750 0.400 2.640 6.100 ;
        RECT 3.640 3.060 3.650 3.100 ;
      LAYER li1 ;
        RECT -0.510 3.380 -0.340 5.870 ;
        RECT 0.040 3.370 0.210 5.870 ;
        RECT 0.590 3.370 0.760 5.870 ;
        RECT 1.140 5.560 1.310 5.870 ;
        RECT 0.880 5.300 1.310 5.560 ;
        RECT 1.140 3.370 1.310 5.300 ;
        RECT 1.690 4.880 1.860 5.870 ;
        RECT 2.240 5.560 2.410 5.870 ;
        RECT 1.970 5.300 2.410 5.560 ;
        RECT 1.430 4.620 1.860 4.880 ;
        RECT 1.690 3.510 1.860 4.620 ;
        RECT 1.430 3.370 1.860 3.510 ;
        RECT 2.240 3.370 2.410 5.300 ;
        RECT 3.070 5.510 3.390 5.550 ;
        RECT 3.070 5.320 3.400 5.510 ;
        RECT 3.070 5.290 3.390 5.320 ;
        RECT 4.250 4.920 4.420 5.680 ;
        RECT 2.520 4.820 2.840 4.860 ;
        RECT 2.520 4.630 2.850 4.820 ;
        RECT 3.630 4.810 3.950 4.850 ;
        RECT 2.520 4.600 2.840 4.630 ;
        RECT 3.630 4.620 3.960 4.810 ;
        RECT 3.630 4.590 3.950 4.620 ;
        RECT 2.520 3.470 2.840 3.510 ;
        RECT 3.620 3.470 3.940 3.510 ;
        RECT 1.430 3.280 1.760 3.370 ;
        RECT 2.520 3.280 2.850 3.470 ;
        RECT 3.620 3.280 3.950 3.470 ;
        RECT 1.430 3.250 1.750 3.280 ;
        RECT 2.520 3.250 2.840 3.280 ;
        RECT 3.620 3.250 3.940 3.280 ;
        RECT 0.960 3.160 1.120 3.190 ;
        RECT -0.510 0.550 -0.340 3.040 ;
        RECT 0.040 1.020 0.210 3.040 ;
        RECT 0.590 1.020 0.760 3.040 ;
        RECT 0.960 2.820 1.130 3.160 ;
        RECT 1.510 3.150 1.670 3.190 ;
        RECT 0.960 2.810 1.120 2.820 ;
        RECT 1.140 2.780 1.310 3.040 ;
        RECT 1.510 2.820 1.680 3.150 ;
        RECT 1.510 2.810 1.670 2.820 ;
        RECT 0.870 2.520 1.310 2.780 ;
        RECT 1.140 1.410 1.310 2.520 ;
        RECT 0.870 1.150 1.310 1.410 ;
        RECT 0.040 0.540 0.760 1.020 ;
        RECT 1.140 0.540 1.310 1.150 ;
        RECT 1.690 0.730 1.860 3.040 ;
        RECT 2.060 2.820 2.230 3.220 ;
        RECT 2.610 3.150 2.770 3.190 ;
        RECT 3.160 3.150 3.320 3.190 ;
        RECT 3.710 3.170 3.870 3.190 ;
        RECT 2.060 2.810 2.220 2.820 ;
        RECT 2.240 2.780 2.410 3.040 ;
        RECT 2.610 2.820 2.780 3.150 ;
        RECT 3.160 2.820 3.330 3.150 ;
        RECT 3.710 2.820 3.880 3.170 ;
        RECT 2.610 2.810 2.770 2.820 ;
        RECT 3.160 2.810 3.320 2.820 ;
        RECT 3.710 2.810 3.870 2.820 ;
        RECT 1.970 2.520 2.410 2.780 ;
        RECT 3.070 2.740 3.390 2.780 ;
        RECT 3.070 2.550 3.400 2.740 ;
        RECT 3.070 2.520 3.390 2.550 ;
        RECT 2.240 1.410 2.410 2.520 ;
        RECT 1.970 1.150 2.410 1.410 ;
        RECT 3.070 1.370 3.390 1.410 ;
        RECT 3.070 1.180 3.400 1.370 ;
        RECT 3.070 1.150 3.390 1.180 ;
        RECT 1.430 0.540 1.860 0.730 ;
        RECT 2.240 0.540 2.410 1.150 ;
        RECT 2.520 0.690 2.840 0.730 ;
        RECT 3.620 0.700 3.940 0.740 ;
        RECT 0.200 0.010 0.710 0.540 ;
        RECT 1.430 0.500 1.760 0.540 ;
        RECT 2.520 0.500 2.850 0.690 ;
        RECT 3.620 0.510 3.950 0.700 ;
        RECT 1.430 0.470 1.750 0.500 ;
        RECT 2.520 0.470 2.840 0.500 ;
        RECT 3.620 0.480 3.940 0.510 ;
      LAYER mcon ;
        RECT 0.940 5.340 1.110 5.510 ;
        RECT 2.030 5.340 2.200 5.510 ;
        RECT 1.490 4.660 1.660 4.830 ;
        RECT 1.490 3.290 1.660 3.460 ;
        RECT 4.250 5.510 4.420 5.680 ;
        RECT 3.130 5.330 3.300 5.500 ;
        RECT 4.250 5.170 4.420 5.340 ;
        RECT 2.580 4.640 2.750 4.810 ;
        RECT 3.690 4.630 3.860 4.800 ;
        RECT 2.580 3.290 2.750 3.460 ;
        RECT 3.680 3.290 3.850 3.460 ;
        RECT 0.930 2.560 1.100 2.730 ;
        RECT 0.930 1.190 1.100 1.360 ;
        RECT 0.360 0.550 0.530 0.720 ;
        RECT 2.030 2.560 2.200 2.730 ;
        RECT 3.130 2.560 3.300 2.730 ;
        RECT 2.030 1.190 2.200 1.360 ;
        RECT 3.130 1.190 3.300 1.360 ;
        RECT 1.490 0.510 1.660 0.680 ;
        RECT 2.580 0.510 2.750 0.680 ;
        RECT 3.680 0.520 3.850 0.690 ;
        RECT 0.370 0.080 0.540 0.250 ;
      LAYER met1 ;
        RECT 0.870 5.270 1.190 5.590 ;
        RECT 1.960 5.270 2.280 5.590 ;
        RECT 3.060 5.260 3.380 5.580 ;
        RECT 1.420 4.590 1.740 4.910 ;
        RECT 2.510 4.570 2.830 4.890 ;
        RECT 3.620 4.560 3.940 4.880 ;
        RECT 1.420 3.220 1.740 3.540 ;
        RECT 2.510 3.220 2.830 3.540 ;
        RECT 3.610 3.220 3.930 3.540 ;
        RECT 0.860 2.490 1.180 2.810 ;
        RECT 1.960 2.490 2.280 2.810 ;
        RECT 3.060 2.490 3.380 2.810 ;
        RECT 0.860 1.120 1.180 1.440 ;
        RECT 1.960 1.120 2.280 1.440 ;
        RECT 3.060 1.120 3.380 1.440 ;
        RECT 0.290 0.480 0.610 0.800 ;
        RECT 1.420 0.440 1.740 0.760 ;
        RECT 2.510 0.440 2.830 0.760 ;
        RECT 3.610 0.450 3.930 0.770 ;
        RECT 0.300 0.010 0.620 0.330 ;
      LAYER via ;
        RECT 0.900 5.300 1.160 5.560 ;
        RECT 1.990 5.300 2.250 5.560 ;
        RECT 3.090 5.290 3.350 5.550 ;
        RECT 1.450 4.620 1.710 4.880 ;
        RECT 2.540 4.600 2.800 4.860 ;
        RECT 3.650 4.590 3.910 4.850 ;
        RECT 1.450 3.250 1.710 3.510 ;
        RECT 2.540 3.250 2.800 3.510 ;
        RECT 3.640 3.250 3.900 3.510 ;
        RECT 0.890 2.520 1.150 2.780 ;
        RECT 1.990 2.520 2.250 2.780 ;
        RECT 3.090 2.520 3.350 2.780 ;
        RECT 0.890 1.150 1.150 1.410 ;
        RECT 1.990 1.150 2.250 1.410 ;
        RECT 3.090 1.150 3.350 1.410 ;
        RECT 0.320 0.510 0.580 0.770 ;
        RECT 1.450 0.470 1.710 0.730 ;
        RECT 2.540 0.470 2.800 0.730 ;
        RECT 3.640 0.480 3.900 0.740 ;
        RECT 0.330 0.040 0.590 0.300 ;
  END
END sky130_hilas_pFETLarge

MACRO sky130_hilas_VinjInv2
  CLASS BLOCK ;
  FOREIGN sky130_hilas_VinjInv2 ;
  ORIGIN 3.360 -1.440 ;
  SIZE 3.610 BY 1.640 ;
  OBS
      LAYER nwell ;
        RECT -3.360 1.440 -1.380 3.080 ;
      LAYER li1 ;
        RECT -2.740 2.650 -2.570 2.790 ;
        RECT -2.740 2.480 -2.550 2.650 ;
        RECT -2.740 2.380 -2.570 2.480 ;
        RECT -3.170 2.000 -3.000 2.100 ;
        RECT -3.190 1.830 -3.000 2.000 ;
        RECT -3.170 1.770 -3.000 1.830 ;
        RECT -2.750 2.040 -2.580 2.100 ;
        RECT -2.750 1.770 -2.500 2.040 ;
        RECT -2.010 2.020 -1.760 2.100 ;
        RECT -2.010 1.850 -0.710 2.020 ;
        RECT -0.150 2.010 0.020 2.640 ;
        RECT -2.740 1.750 -2.500 1.770 ;
        RECT -1.930 1.760 -1.760 1.850 ;
        RECT -0.230 1.840 0.100 2.010 ;
      LAYER mcon ;
        RECT -2.720 2.480 -2.550 2.650 ;
        RECT -0.150 2.120 0.020 2.290 ;
        RECT -2.710 1.800 -2.540 1.970 ;
        RECT -1.370 1.850 -1.200 2.020 ;
      LAYER met1 ;
        RECT -2.750 2.700 -2.530 3.040 ;
        RECT -2.750 2.440 -2.520 2.700 ;
        RECT -3.280 1.760 -2.970 2.110 ;
        RECT -2.750 2.040 -2.530 2.440 ;
        RECT -2.750 1.730 -2.500 2.040 ;
        RECT -1.450 1.800 -1.130 2.060 ;
        RECT -2.750 1.530 -2.530 1.730 ;
        RECT -0.180 1.530 0.050 3.040 ;
      LAYER via ;
        RECT -3.250 1.790 -2.990 2.050 ;
        RECT -1.420 1.800 -1.160 2.060 ;
      LAYER met2 ;
        RECT -3.360 2.470 0.250 2.650 ;
        RECT -3.280 1.950 -2.960 2.050 ;
        RECT -3.290 1.790 -2.960 1.950 ;
        RECT -1.450 1.980 -1.130 2.060 ;
        RECT -1.450 1.800 0.250 1.980 ;
  END
END sky130_hilas_VinjInv2

MACRO sky130_hilas_capacitorSize03
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize03 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.790 BY 5.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 4.960 2.630 5.620 3.290 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 2.570 4.530 3.020 4.540 ;
        RECT 2.550 4.040 3.070 4.530 ;
        RECT 0.110 3.190 0.770 3.250 ;
        RECT 2.580 3.200 3.020 4.040 ;
        RECT 1.160 3.190 2.170 3.200 ;
        RECT 2.570 3.190 3.030 3.200 ;
        RECT 0.110 2.690 3.030 3.190 ;
        RECT 0.110 2.680 1.520 2.690 ;
        RECT 0.110 2.590 0.770 2.680 ;
        RECT 2.570 2.030 3.030 2.690 ;
        RECT 2.570 1.520 3.050 2.030 ;
        RECT 2.550 1.030 3.070 1.520 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 0.000 5.270 5.780 5.450 ;
        RECT 0.000 4.840 5.780 5.020 ;
        RECT 0.030 3.840 5.780 4.020 ;
        RECT 0.030 3.410 5.780 3.590 ;
        RECT 0.240 3.070 0.610 3.130 ;
        RECT 0.020 2.790 0.610 3.070 ;
        RECT 0.240 2.730 0.610 2.790 ;
        RECT 5.090 3.110 5.460 3.170 ;
        RECT 5.090 2.830 5.790 3.110 ;
        RECT 5.090 2.770 5.460 2.830 ;
        RECT 0.030 2.260 5.780 2.430 ;
        RECT 0.030 1.840 5.780 2.010 ;
        RECT 0.030 0.860 5.780 1.030 ;
        RECT 0.030 0.420 5.780 0.590 ;
      LAYER via2 ;
        RECT 0.290 2.790 0.570 3.070 ;
        RECT 5.140 2.830 5.420 3.110 ;
      LAYER met3 ;
        RECT 1.450 3.320 4.290 5.870 ;
        RECT 0.020 2.530 0.810 3.280 ;
        RECT 1.450 2.570 5.660 3.320 ;
        RECT 1.450 0.000 4.290 2.570 ;
      LAYER via3 ;
        RECT 0.210 2.680 0.640 3.160 ;
        RECT 5.060 2.720 5.490 3.200 ;
  END
END sky130_hilas_capacitorSize03

MACRO sky130_hilas_swc4x1BiasCell
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x1BiasCell ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.110 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN ROW1
    USE ANALOG ;
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 7.630 5.120 7.940 5.140 ;
        RECT 0.020 4.940 10.100 5.120 ;
        RECT 0.020 4.930 0.170 4.940 ;
        RECT 7.630 4.810 7.940 4.940 ;
    END
  END ROW1
  PIN ROW2
    USE ANALOG ;
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 0.000 4.120 0.140 4.140 ;
        RECT 7.630 4.120 7.940 4.250 ;
        RECT 0.000 3.940 10.110 4.120 ;
        RECT 7.630 3.920 7.940 3.940 ;
    END
  END ROW2
  PIN ROW3
    USE ANALOG ;
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 7.630 2.110 7.940 2.130 ;
        RECT 0.030 1.950 10.100 2.110 ;
        RECT 0.040 1.940 10.100 1.950 ;
        RECT 7.540 1.930 10.100 1.940 ;
        RECT 7.630 1.800 7.940 1.930 ;
    END
  END ROW3
  PIN ROW4
    USE ANALOG ;
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 7.630 1.130 7.940 1.250 ;
        RECT 0.030 1.120 7.940 1.130 ;
        RECT 0.030 0.960 10.100 1.120 ;
        RECT 0.820 0.870 2.360 0.960 ;
        RECT 7.540 0.940 10.100 0.960 ;
        RECT 7.630 0.920 7.940 0.940 ;
    END
  END ROW4
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 1.978000 ;
    PORT
      LAYER nwell ;
        RECT 0.030 5.420 1.760 6.050 ;
        RECT 0.020 2.350 1.760 5.420 ;
        RECT 0.030 0.000 1.760 2.350 ;
      LAYER met1 ;
        RECT 0.380 0.000 0.780 6.050 ;
    END
  END VTUN
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 2.743300 ;
    PORT
      LAYER nwell ;
        RECT 3.780 0.000 6.010 6.050 ;
      LAYER met1 ;
        RECT 4.430 4.130 4.810 6.050 ;
        RECT 4.420 2.270 4.810 4.130 ;
        RECT 4.430 0.000 4.810 2.270 ;
    END
  END GATE1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 7.540 6.040 10.090 6.050 ;
        RECT 7.540 0.020 10.100 6.040 ;
        RECT 7.540 0.010 10.090 0.020 ;
      LAYER met1 ;
        RECT 9.580 5.400 9.740 6.050 ;
        RECT 9.470 4.850 9.740 5.400 ;
        RECT 9.470 4.800 9.750 4.850 ;
        RECT 9.580 4.710 9.750 4.800 ;
        RECT 9.580 4.350 9.740 4.710 ;
        RECT 9.580 4.260 9.750 4.350 ;
        RECT 9.470 4.210 9.750 4.260 ;
        RECT 9.470 3.660 9.740 4.210 ;
        RECT 9.580 2.390 9.740 3.660 ;
        RECT 9.470 1.840 9.740 2.390 ;
        RECT 9.470 1.790 9.750 1.840 ;
        RECT 9.580 1.700 9.750 1.790 ;
        RECT 9.580 1.350 9.740 1.700 ;
        RECT 9.580 1.260 9.750 1.350 ;
        RECT 9.470 1.210 9.750 1.260 ;
        RECT 9.470 0.660 9.740 1.210 ;
        RECT 9.580 0.010 9.740 0.660 ;
    END
  END VINJ
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 8.770 5.370 8.930 6.050 ;
        RECT 8.770 5.350 8.970 5.370 ;
        RECT 8.750 5.110 8.980 5.350 ;
        RECT 8.770 4.890 8.970 5.110 ;
        RECT 8.770 4.170 8.930 4.890 ;
        RECT 8.770 3.950 8.970 4.170 ;
        RECT 8.750 3.710 8.980 3.950 ;
        RECT 8.770 3.690 8.970 3.710 ;
        RECT 8.770 2.360 8.930 3.690 ;
        RECT 8.770 2.340 8.970 2.360 ;
        RECT 8.750 2.100 8.980 2.340 ;
        RECT 8.770 1.880 8.970 2.100 ;
        RECT 8.770 1.170 8.930 1.880 ;
        RECT 8.770 0.950 8.970 1.170 ;
        RECT 8.750 0.710 8.980 0.950 ;
        RECT 8.770 0.690 8.970 0.710 ;
        RECT 8.770 0.010 8.930 0.690 ;
    END
  END VPWR
  PIN COLSEL1
    USE ANALOG ;
    ANTENNAGATEAREA 0.620000 ;
    PORT
      LAYER met1 ;
        RECT 9.140 5.060 9.330 6.050 ;
        RECT 9.160 4.940 9.330 5.060 ;
        RECT 9.170 4.120 9.330 4.940 ;
        RECT 9.160 4.000 9.330 4.120 ;
        RECT 9.140 3.140 9.330 4.000 ;
        RECT 9.120 2.910 9.360 3.140 ;
        RECT 9.140 2.050 9.330 2.910 ;
        RECT 9.160 1.930 9.330 2.050 ;
        RECT 9.170 1.120 9.330 1.930 ;
        RECT 9.160 1.000 9.330 1.120 ;
        RECT 9.140 0.010 9.330 1.000 ;
    END
  END COLSEL1
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER met2 ;
        RECT 7.630 5.550 7.940 5.690 ;
        RECT 7.530 5.370 10.100 5.550 ;
        RECT 7.630 5.360 7.940 5.370 ;
    END
  END DRAIN1
  PIN DRAIN2
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER met2 ;
        RECT 7.630 3.690 7.940 3.700 ;
        RECT 7.630 3.650 10.100 3.690 ;
        RECT 7.540 3.510 10.100 3.650 ;
        RECT 7.630 3.370 7.940 3.510 ;
    END
  END DRAIN2
  PIN DRAIN3
    USE ANALOG ;
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER met2 ;
        RECT 7.630 2.540 7.940 2.680 ;
        RECT 7.630 2.530 10.110 2.540 ;
        RECT 7.510 2.360 10.110 2.530 ;
        RECT 7.630 2.350 7.940 2.360 ;
    END
  END DRAIN3
  PIN DRAIN4
    USE ANALOG ;
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER met2 ;
        RECT 7.630 0.690 7.940 0.700 ;
        RECT 7.530 0.520 10.100 0.690 ;
        RECT 7.630 0.510 10.100 0.520 ;
        RECT 7.630 0.370 7.940 0.510 ;
    END
  END DRAIN4
  PIN VGND
    ANTENNADIFFAREA 1.053100 ;
    PORT
      LAYER met2 ;
        RECT 2.560 1.520 2.890 1.550 ;
        RECT 6.590 1.520 6.910 1.580 ;
        RECT 2.560 1.350 6.910 1.520 ;
        RECT 2.560 1.290 2.890 1.350 ;
        RECT 6.590 1.300 6.910 1.350 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.620 1.610 6.870 6.050 ;
        RECT 6.610 1.580 6.890 1.610 ;
        RECT 6.600 1.300 6.900 1.580 ;
        RECT 6.610 1.280 6.890 1.300 ;
        RECT 6.620 0.000 6.870 1.280 ;
      LAYER via ;
        RECT 6.620 1.310 6.880 1.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.590 1.580 2.860 6.050 ;
        RECT 2.570 1.270 2.880 1.580 ;
        RECT 2.590 0.000 2.860 1.270 ;
      LAYER via ;
        RECT 2.590 1.290 2.860 1.550 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 7.640 5.640 7.960 5.650 ;
        RECT 7.640 5.470 8.220 5.640 ;
        RECT 7.640 5.420 7.970 5.470 ;
        RECT 7.640 5.390 7.960 5.420 ;
        RECT 9.500 5.370 9.700 5.720 ;
        RECT 7.640 5.060 7.960 5.100 ;
        RECT 7.640 5.020 7.970 5.060 ;
        RECT 7.640 4.850 8.220 5.020 ;
        RECT 7.640 4.840 7.960 4.850 ;
        RECT 2.640 4.300 2.810 4.810 ;
        RECT 8.770 4.780 8.970 5.350 ;
        RECT 9.500 5.340 9.710 5.370 ;
        RECT 6.660 4.270 6.830 4.780 ;
        RECT 9.490 4.750 9.710 5.340 ;
        RECT 7.640 4.210 7.960 4.220 ;
        RECT 7.640 4.040 8.220 4.210 ;
        RECT 7.640 4.000 7.970 4.040 ;
        RECT 7.640 3.960 7.960 4.000 ;
        RECT 8.770 3.710 8.970 4.280 ;
        RECT 9.490 3.720 9.710 4.310 ;
        RECT 9.500 3.690 9.710 3.720 ;
        RECT 7.640 3.640 7.960 3.670 ;
        RECT 0.450 2.800 1.000 3.230 ;
        RECT 2.650 2.350 2.820 3.540 ;
        RECT 4.480 2.730 5.030 3.160 ;
        RECT 6.670 2.410 6.840 3.600 ;
        RECT 7.640 3.590 7.970 3.640 ;
        RECT 7.640 3.420 8.220 3.590 ;
        RECT 7.640 3.410 7.960 3.420 ;
        RECT 9.500 3.340 9.700 3.690 ;
        RECT 8.890 2.940 9.330 3.110 ;
        RECT 7.640 2.630 7.960 2.640 ;
        RECT 7.640 2.460 8.220 2.630 ;
        RECT 7.640 2.410 7.970 2.460 ;
        RECT 7.640 2.380 7.960 2.410 ;
        RECT 9.500 2.360 9.700 2.710 ;
        RECT 7.640 2.050 7.960 2.090 ;
        RECT 7.640 2.010 7.970 2.050 ;
        RECT 7.640 1.840 8.220 2.010 ;
        RECT 7.640 1.830 7.960 1.840 ;
        RECT 8.770 1.770 8.970 2.340 ;
        RECT 9.500 2.330 9.710 2.360 ;
        RECT 9.490 1.740 9.710 2.330 ;
        RECT 7.640 1.210 7.960 1.220 ;
        RECT 7.640 1.040 8.220 1.210 ;
        RECT 7.640 1.000 7.970 1.040 ;
        RECT 7.640 0.960 7.960 1.000 ;
        RECT 8.770 0.710 8.970 1.280 ;
        RECT 9.490 0.720 9.710 1.310 ;
        RECT 9.500 0.690 9.710 0.720 ;
        RECT 7.640 0.640 7.960 0.670 ;
        RECT 7.640 0.590 7.970 0.640 ;
        RECT 7.640 0.420 8.220 0.590 ;
        RECT 7.640 0.410 7.960 0.420 ;
        RECT 9.500 0.340 9.700 0.690 ;
      LAYER mcon ;
        RECT 7.700 5.430 7.870 5.600 ;
        RECT 8.780 5.140 8.950 5.310 ;
        RECT 7.700 4.880 7.870 5.050 ;
        RECT 2.640 4.640 2.810 4.810 ;
        RECT 9.510 5.170 9.680 5.340 ;
        RECT 6.660 4.610 6.830 4.780 ;
        RECT 7.700 4.010 7.870 4.180 ;
        RECT 8.780 3.750 8.950 3.920 ;
        RECT 9.510 3.720 9.680 3.890 ;
        RECT 2.650 3.370 2.820 3.540 ;
        RECT 0.450 2.880 0.720 3.150 ;
        RECT 2.650 3.030 2.820 3.200 ;
        RECT 6.670 3.430 6.840 3.600 ;
        RECT 7.700 3.460 7.870 3.630 ;
        RECT 2.650 2.690 2.820 2.860 ;
        RECT 4.480 2.810 4.750 3.080 ;
        RECT 6.670 3.090 6.840 3.260 ;
        RECT 9.150 2.940 9.330 3.110 ;
        RECT 6.670 2.750 6.840 2.920 ;
        RECT 7.700 2.420 7.870 2.590 ;
        RECT 8.780 2.130 8.950 2.300 ;
        RECT 7.700 1.870 7.870 2.040 ;
        RECT 9.510 2.160 9.680 2.330 ;
        RECT 7.700 1.010 7.870 1.180 ;
        RECT 8.780 0.750 8.950 0.920 ;
        RECT 9.510 0.720 9.680 0.890 ;
        RECT 7.700 0.460 7.870 0.630 ;
      LAYER met1 ;
        RECT 7.630 5.360 7.950 5.680 ;
        RECT 7.630 4.810 7.950 5.130 ;
        RECT 7.630 3.930 7.950 4.250 ;
        RECT 7.630 3.380 7.950 3.700 ;
        RECT 7.630 2.350 7.950 2.670 ;
        RECT 7.630 1.800 7.950 2.120 ;
        RECT 7.630 0.930 7.950 1.250 ;
        RECT 7.630 0.380 7.950 0.700 ;
      LAYER via ;
        RECT 7.660 5.390 7.920 5.650 ;
        RECT 7.660 4.840 7.920 5.100 ;
        RECT 7.660 3.960 7.920 4.220 ;
        RECT 7.660 3.410 7.920 3.670 ;
        RECT 7.660 2.380 7.920 2.640 ;
        RECT 7.660 1.830 7.920 2.090 ;
        RECT 7.660 0.960 7.920 1.220 ;
        RECT 7.660 0.410 7.920 0.670 ;
  END
END sky130_hilas_swc4x1BiasCell

MACRO sky130_hilas_FGtrans2x1cell
  CLASS CORE ;
  FOREIGN sky130_hilas_FGtrans2x1cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.520 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN COLSEL1
    USE ANALOG ;
    ANTENNAGATEAREA 0.310000 ;
    PORT
      LAYER met1 ;
        RECT 10.560 4.590 10.750 6.050 ;
        RECT 10.560 4.560 10.780 4.590 ;
        RECT 10.540 4.290 10.790 4.560 ;
        RECT 10.550 4.280 10.790 4.290 ;
        RECT 10.550 4.040 10.780 4.280 ;
        RECT 10.590 2.010 10.750 4.040 ;
        RECT 10.550 1.770 10.780 2.010 ;
        RECT 10.550 1.760 10.790 1.770 ;
        RECT 10.540 1.490 10.790 1.760 ;
        RECT 10.560 1.460 10.780 1.490 ;
        RECT 10.560 0.000 10.750 1.460 ;
    END
  END COLSEL1
  PIN VINJ
    USE ANALOG ;
    ANTENNADIFFAREA 0.510000 ;
    PORT
      LAYER nwell ;
        RECT 8.210 0.010 11.520 6.040 ;
      LAYER met1 ;
        RECT 11.000 5.400 11.160 6.050 ;
        RECT 10.890 4.850 11.160 5.400 ;
        RECT 10.890 4.800 11.170 4.850 ;
        RECT 11.000 4.710 11.170 4.800 ;
        RECT 11.000 1.340 11.160 4.710 ;
        RECT 11.000 1.250 11.170 1.340 ;
        RECT 10.890 1.200 11.170 1.250 ;
        RECT 10.890 0.650 11.160 1.200 ;
        RECT 11.000 0.000 11.160 0.650 ;
    END
  END VINJ
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.105400 ;
    PORT
      LAYER met2 ;
        RECT 8.790 5.560 9.110 5.570 ;
        RECT 8.790 5.550 9.350 5.560 ;
        RECT 0.000 5.370 11.520 5.550 ;
        RECT 9.040 5.230 9.350 5.370 ;
    END
  END DRAIN1
  PIN DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.105400 ;
    PORT
      LAYER met2 ;
        RECT 9.040 0.680 9.350 0.820 ;
        RECT 9.040 0.670 11.520 0.680 ;
        RECT 0.000 0.520 11.520 0.670 ;
        RECT 9.040 0.500 11.520 0.520 ;
        RECT 9.040 0.490 9.350 0.500 ;
    END
  END DRAIN2
  PIN PROG
    USE ANALOG ;
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER met1 ;
        RECT 7.790 3.330 8.000 6.050 ;
        RECT 7.790 2.820 8.030 3.330 ;
        RECT 7.790 0.000 8.000 2.820 ;
    END
  END PROG
  PIN RUN
    USE ANALOG ;
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER met1 ;
        RECT 6.740 1.520 6.920 6.050 ;
        RECT 6.690 1.180 6.980 1.520 ;
        RECT 6.740 0.000 6.920 1.180 ;
    END
  END RUN
  PIN VIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.217200 ;
    PORT
      LAYER met1 ;
        RECT 8.670 2.620 8.860 2.750 ;
        RECT 8.650 2.330 8.880 2.620 ;
        RECT 8.670 0.710 8.860 2.330 ;
        RECT 8.630 0.500 8.860 0.710 ;
        RECT 8.630 0.420 8.870 0.500 ;
        RECT 8.640 0.000 8.870 0.420 ;
    END
  END VIN2
  PIN VIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.217200 ;
    PORT
      LAYER met1 ;
        RECT 8.670 5.680 8.880 6.050 ;
        RECT 8.660 5.390 8.890 5.680 ;
        RECT 8.670 3.690 8.880 5.390 ;
        RECT 8.660 3.400 8.890 3.690 ;
        RECT 8.670 3.260 8.880 3.400 ;
    END
  END VIN1
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 0.434600 ;
    PORT
      LAYER met1 ;
        RECT 8.220 5.120 8.410 6.050 ;
        RECT 8.190 4.830 8.420 5.120 ;
        RECT 8.220 2.800 8.410 4.830 ;
        RECT 8.190 2.510 8.420 2.800 ;
        RECT 8.220 1.220 8.410 2.510 ;
        RECT 8.200 0.930 8.430 1.220 ;
        RECT 8.220 0.000 8.410 0.930 ;
    END
  END GATE1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2.820 0.000 3.050 6.050 ;
    END
  END VGND
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 2.516100 ;
    PORT
      LAYER nwell ;
        RECT 0.000 5.300 1.730 6.050 ;
        RECT 0.000 1.730 1.740 5.300 ;
        RECT 0.000 0.010 1.730 1.730 ;
      LAYER met1 ;
        RECT 0.340 0.000 0.760 6.050 ;
    END
  END VTUN
  PIN COL1
    ANTENNADIFFAREA 1.030400 ;
    PORT
      LAYER met2 ;
        RECT 10.140 3.130 10.460 3.160 ;
        RECT 0.000 2.900 10.460 3.130 ;
    END
  END COL1
  PIN ROW1
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 9.430 4.010 9.740 4.030 ;
        RECT 0.000 3.820 9.740 4.010 ;
        RECT 9.430 3.700 9.740 3.820 ;
    END
  END ROW1
  PIN ROW2
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 9.440 2.150 9.750 2.340 ;
        RECT 0.000 2.010 9.750 2.150 ;
        RECT 0.000 1.960 9.720 2.010 ;
    END
  END ROW2
  OBS
      LAYER nwell ;
        RECT 3.760 3.660 6.480 5.310 ;
        RECT 3.770 3.620 6.480 3.660 ;
        RECT 3.770 2.290 6.480 2.330 ;
        RECT 3.760 0.640 6.480 2.290 ;
      LAYER li1 ;
        RECT 8.680 5.620 8.870 5.650 ;
        RECT 7.810 5.450 8.870 5.620 ;
        RECT 9.110 5.470 9.640 5.640 ;
        RECT 7.810 5.060 7.980 5.450 ;
        RECT 8.680 5.420 8.870 5.450 ;
        RECT 10.920 5.370 11.120 5.720 ;
        RECT 10.920 5.340 11.130 5.370 ;
        RECT 7.240 4.890 7.980 5.060 ;
        RECT 8.210 5.060 8.400 5.090 ;
        RECT 8.210 4.890 8.940 5.060 ;
        RECT 8.210 4.860 8.400 4.890 ;
        RECT 0.430 3.910 0.980 4.340 ;
        RECT 5.950 4.270 6.180 4.790 ;
        RECT 5.950 4.100 8.940 4.270 ;
        RECT 9.360 3.990 9.530 5.080 ;
        RECT 9.360 3.950 9.760 3.990 ;
        RECT 9.360 3.760 9.770 3.950 ;
        RECT 9.360 3.730 9.760 3.760 ;
        RECT 8.680 3.480 8.870 3.660 ;
        RECT 3.030 3.080 3.220 3.480 ;
        RECT 7.250 3.310 7.590 3.480 ;
        RECT 2.840 3.070 3.220 3.080 ;
        RECT 2.840 2.890 6.580 3.070 ;
        RECT 2.840 2.850 3.220 2.890 ;
        RECT 0.430 2.180 0.980 2.610 ;
        RECT 3.030 2.470 3.220 2.850 ;
        RECT 7.330 2.740 7.500 3.310 ;
        RECT 7.810 2.900 8.020 3.330 ;
        RECT 8.590 3.310 8.940 3.480 ;
        RECT 9.360 3.390 9.530 3.730 ;
        RECT 10.190 3.480 10.360 5.090 ;
        RECT 10.910 4.760 11.130 5.340 ;
        RECT 10.920 4.750 11.130 4.760 ;
        RECT 10.560 4.580 10.750 4.590 ;
        RECT 10.560 4.290 10.760 4.580 ;
        RECT 10.550 3.960 10.790 4.290 ;
        RECT 10.190 3.290 10.370 3.480 ;
        RECT 7.830 2.880 8.000 2.900 ;
        RECT 7.250 2.710 7.590 2.740 ;
        RECT 8.210 2.720 8.400 2.770 ;
        RECT 8.170 2.710 8.400 2.720 ;
        RECT 7.250 2.570 8.400 2.710 ;
        RECT 8.590 2.570 8.940 2.740 ;
        RECT 7.420 2.540 8.400 2.570 ;
        RECT 7.420 2.510 8.260 2.540 ;
        RECT 8.670 2.360 8.860 2.570 ;
        RECT 9.360 2.300 9.530 2.660 ;
        RECT 10.190 2.570 10.370 2.760 ;
        RECT 9.360 2.260 9.770 2.300 ;
        RECT 9.360 2.070 9.780 2.260 ;
        RECT 9.360 2.040 9.770 2.070 ;
        RECT 6.010 1.850 8.940 1.950 ;
        RECT 5.950 1.780 8.940 1.850 ;
        RECT 5.950 1.160 6.180 1.780 ;
        RECT 6.750 1.460 6.920 1.520 ;
        RECT 6.730 1.250 6.940 1.460 ;
        RECT 6.750 1.180 6.920 1.250 ;
        RECT 8.220 1.160 8.410 1.190 ;
        RECT 7.240 0.990 8.050 1.160 ;
        RECT 7.860 0.650 8.050 0.990 ;
        RECT 8.220 0.990 8.940 1.160 ;
        RECT 8.220 0.960 8.410 0.990 ;
        RECT 9.360 0.970 9.530 2.040 ;
        RECT 10.190 0.960 10.360 2.570 ;
        RECT 10.550 1.760 10.790 2.090 ;
        RECT 10.560 1.470 10.760 1.760 ;
        RECT 10.560 1.460 10.750 1.470 ;
        RECT 10.920 1.290 11.130 1.300 ;
        RECT 10.910 0.710 11.130 1.290 ;
        RECT 10.920 0.680 11.130 0.710 ;
        RECT 8.650 0.650 8.840 0.680 ;
        RECT 7.860 0.470 8.840 0.650 ;
        RECT 8.650 0.450 8.840 0.470 ;
        RECT 9.110 0.410 9.640 0.580 ;
        RECT 10.920 0.330 11.120 0.680 ;
      LAYER mcon ;
        RECT 8.690 5.450 8.860 5.620 ;
        RECT 10.930 5.170 11.100 5.340 ;
        RECT 8.220 4.890 8.390 5.060 ;
        RECT 5.980 4.590 6.150 4.760 ;
        RECT 0.430 3.990 0.700 4.260 ;
        RECT 5.980 4.140 6.150 4.310 ;
        RECT 9.500 3.770 9.670 3.940 ;
        RECT 8.690 3.460 8.860 3.630 ;
        RECT 2.850 2.880 3.020 3.050 ;
        RECT 0.430 2.260 0.700 2.530 ;
        RECT 10.570 4.330 10.750 4.520 ;
        RECT 8.220 2.570 8.390 2.740 ;
        RECT 8.680 2.390 8.850 2.560 ;
        RECT 9.510 2.080 9.680 2.250 ;
        RECT 5.980 1.640 6.150 1.810 ;
        RECT 5.980 1.190 6.150 1.360 ;
        RECT 8.230 0.990 8.400 1.160 ;
        RECT 10.570 1.530 10.750 1.720 ;
        RECT 10.930 0.710 11.100 0.880 ;
        RECT 8.660 0.480 8.830 0.650 ;
      LAYER met1 ;
        RECT 9.040 5.230 9.350 5.670 ;
        RECT 5.940 4.050 6.200 4.840 ;
        RECT 9.430 3.700 9.750 4.020 ;
        RECT 10.160 3.190 10.400 3.610 ;
        RECT 10.160 2.870 10.430 3.190 ;
        RECT 10.160 2.440 10.400 2.870 ;
        RECT 9.440 2.010 9.760 2.330 ;
        RECT 5.940 1.110 6.200 1.900 ;
        RECT 9.040 0.380 9.350 0.820 ;
      LAYER via ;
        RECT 9.070 5.260 9.330 5.520 ;
        RECT 9.460 3.730 9.720 3.990 ;
        RECT 10.170 2.900 10.430 3.160 ;
        RECT 9.470 2.040 9.730 2.300 ;
        RECT 9.070 0.530 9.330 0.790 ;
  END
END sky130_hilas_FGtrans2x1cell

MACRO sky130_hilas_capacitorSize01
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.420 BY 5.830 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 9.600 2.610 10.260 3.270 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 0.110 3.200 0.770 3.260 ;
        RECT 1.160 3.200 2.170 3.210 ;
        RECT 0.110 2.700 3.800 3.200 ;
        RECT 0.110 2.690 1.520 2.700 ;
        RECT 0.110 2.600 0.770 2.690 ;
        RECT 3.160 1.580 3.790 2.700 ;
        RECT 3.160 1.570 5.310 1.580 ;
        RECT 2.350 1.100 5.390 1.570 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 0.000 5.280 10.420 5.460 ;
        RECT 0.000 4.850 10.420 5.030 ;
        RECT 0.030 3.850 10.420 4.030 ;
        RECT 8.510 3.600 10.420 3.610 ;
        RECT 0.030 3.420 10.420 3.600 ;
        RECT 0.240 3.080 0.610 3.140 ;
        RECT 0.020 2.800 0.610 3.080 ;
        RECT 0.240 2.740 0.610 2.800 ;
        RECT 9.730 3.090 10.100 3.150 ;
        RECT 9.730 2.810 10.420 3.090 ;
        RECT 9.730 2.750 10.100 2.810 ;
        RECT 0.030 2.270 10.420 2.440 ;
        RECT 0.030 1.850 10.420 2.020 ;
        RECT 0.030 0.870 10.420 1.040 ;
        RECT 0.030 0.430 10.420 0.600 ;
      LAYER via2 ;
        RECT 0.290 2.800 0.570 3.080 ;
        RECT 9.780 2.810 10.060 3.090 ;
      LAYER met3 ;
        RECT 1.460 5.800 4.280 5.830 ;
        RECT 1.460 3.300 8.660 5.800 ;
        RECT 0.020 2.540 0.810 3.290 ;
        RECT 1.460 2.550 10.300 3.300 ;
        RECT 1.460 0.020 8.660 2.550 ;
        RECT 4.250 0.000 8.660 0.020 ;
      LAYER via3 ;
        RECT 0.210 2.690 0.640 3.170 ;
        RECT 9.700 2.700 10.130 3.180 ;
  END
END sky130_hilas_capacitorSize01

MACRO sky130_hilas_Tgate4Double01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_Tgate4Double01 ;
  ORIGIN 0.360 1.410 ;
  SIZE 7.080 BY 6.050 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER nwell ;
        RECT -0.240 -1.410 3.230 4.640 ;
      LAYER met1 ;
        RECT 0.380 3.770 0.580 4.640 ;
        RECT 0.370 3.480 0.600 3.770 ;
        RECT 0.380 2.770 0.580 3.480 ;
        RECT 0.370 2.480 0.600 2.770 ;
        RECT 0.380 0.750 0.580 2.480 ;
        RECT 0.370 0.460 0.600 0.750 ;
        RECT 0.380 -0.250 0.580 0.460 ;
        RECT 0.370 -0.540 0.600 -0.250 ;
        RECT 0.380 -1.410 0.580 -0.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.210 3.770 6.400 4.640 ;
        RECT 6.190 3.480 6.420 3.770 ;
        RECT 6.210 2.770 6.400 3.480 ;
        RECT 6.190 2.480 6.420 2.770 ;
        RECT 6.210 0.750 6.400 2.480 ;
        RECT 6.190 0.460 6.420 0.750 ;
        RECT 6.210 -0.250 6.400 0.460 ;
        RECT 6.190 -0.540 6.420 -0.250 ;
        RECT 6.210 -1.410 6.400 -0.540 ;
    END
  END VGND
  PIN INPUT1_1
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.090 4.530 2.400 4.540 ;
        RECT -0.360 4.330 5.480 4.530 ;
        RECT 2.090 4.210 2.400 4.330 ;
        RECT 5.170 4.200 5.480 4.330 ;
    END
  END INPUT1_1
  PIN SELECT1
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER met2 ;
        RECT -0.360 3.350 0.250 3.550 ;
        RECT -0.070 3.260 0.250 3.350 ;
    END
  END SELECT1
  PIN SELECT2
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER met2 ;
        RECT -0.070 2.900 0.250 2.990 ;
        RECT -0.360 2.700 0.250 2.900 ;
    END
  END SELECT2
  PIN INPUT2_2
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 0.740 2.400 1.050 2.410 ;
        RECT 3.660 2.400 3.970 2.410 ;
        RECT -0.360 2.200 4.010 2.400 ;
        RECT 0.740 2.080 1.050 2.200 ;
        RECT 3.660 2.080 3.970 2.200 ;
    END
  END INPUT2_2
  PIN INPUT1_2
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.090 1.920 2.400 2.040 ;
        RECT 5.170 1.920 5.480 2.050 ;
        RECT -0.360 1.720 5.480 1.920 ;
        RECT 2.090 1.710 2.400 1.720 ;
    END
  END INPUT1_2
  PIN SELECT3
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER met2 ;
        RECT -0.360 0.330 0.250 0.530 ;
        RECT -0.070 0.240 0.250 0.330 ;
    END
  END SELECT3
  PIN INPUT2_3
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 0.740 1.030 1.050 1.150 ;
        RECT 3.660 1.030 3.970 1.150 ;
        RECT -0.360 0.830 4.010 1.030 ;
        RECT 0.740 0.820 1.050 0.830 ;
        RECT 3.660 0.820 3.970 0.830 ;
    END
  END INPUT2_3
  PIN SELECT4
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER met2 ;
        RECT -0.070 -0.120 0.250 -0.030 ;
        RECT -0.360 -0.320 0.250 -0.120 ;
    END
  END SELECT4
  PIN INPUT2_4
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 0.740 -0.620 1.050 -0.610 ;
        RECT 3.660 -0.620 3.970 -0.610 ;
        RECT -0.360 -0.820 4.010 -0.620 ;
        RECT 0.740 -0.940 1.050 -0.820 ;
        RECT 3.660 -0.940 3.970 -0.820 ;
    END
  END INPUT2_4
  PIN INPUT1_4
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.090 -1.100 2.400 -0.980 ;
        RECT 5.170 -1.100 5.480 -0.970 ;
        RECT -0.360 -1.300 5.480 -1.100 ;
        RECT 2.090 -1.310 2.400 -1.300 ;
    END
  END INPUT1_4
  PIN OUTPUT4
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER met2 ;
        RECT 1.320 -0.120 1.640 -0.110 ;
        RECT 2.740 -0.120 3.060 -0.100 ;
        RECT 4.490 -0.120 4.810 -0.080 ;
        RECT 5.530 -0.120 5.850 -0.090 ;
        RECT 1.320 -0.320 6.720 -0.120 ;
        RECT 1.320 -0.370 1.640 -0.320 ;
        RECT 2.740 -0.360 3.060 -0.320 ;
        RECT 4.490 -0.340 4.810 -0.320 ;
        RECT 5.530 -0.350 5.850 -0.320 ;
    END
  END OUTPUT4
  PIN OUTPUT3
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER met2 ;
        RECT 1.320 0.530 1.640 0.580 ;
        RECT 2.740 0.530 3.060 0.570 ;
        RECT 4.490 0.530 4.810 0.550 ;
        RECT 5.530 0.530 5.850 0.560 ;
        RECT 1.320 0.330 6.720 0.530 ;
        RECT 1.320 0.320 1.640 0.330 ;
        RECT 2.740 0.310 3.060 0.330 ;
        RECT 4.490 0.290 4.810 0.330 ;
        RECT 5.530 0.300 5.850 0.330 ;
    END
  END OUTPUT3
  PIN OUTPUT2
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER met2 ;
        RECT 1.320 2.900 1.640 2.910 ;
        RECT 2.740 2.900 3.060 2.920 ;
        RECT 4.490 2.900 4.810 2.940 ;
        RECT 5.530 2.900 5.850 2.930 ;
        RECT 1.320 2.700 6.720 2.900 ;
        RECT 1.320 2.650 1.640 2.700 ;
        RECT 2.740 2.660 3.060 2.700 ;
        RECT 4.490 2.680 4.810 2.700 ;
        RECT 5.530 2.670 5.850 2.700 ;
    END
  END OUTPUT2
  PIN OUTPUT1
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER met2 ;
        RECT 1.320 3.550 1.640 3.600 ;
        RECT 2.740 3.550 3.060 3.590 ;
        RECT 4.490 3.550 4.810 3.570 ;
        RECT 5.530 3.550 5.850 3.580 ;
        RECT 1.320 3.350 6.720 3.550 ;
        RECT 1.320 3.340 1.640 3.350 ;
        RECT 2.740 3.330 3.060 3.350 ;
        RECT 4.490 3.310 4.810 3.350 ;
        RECT 5.530 3.320 5.850 3.350 ;
    END
  END OUTPUT1
  PIN INPUT2_1
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 0.740 4.050 1.050 4.170 ;
        RECT 3.660 4.050 3.970 4.170 ;
        RECT -0.360 3.850 4.010 4.050 ;
        RECT 0.740 3.840 1.050 3.850 ;
        RECT 3.660 3.840 3.970 3.850 ;
    END
  END INPUT2_1
  PIN INPUT1_3
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.090 1.510 2.400 1.520 ;
        RECT -0.360 1.310 5.480 1.510 ;
        RECT 2.090 1.190 2.400 1.310 ;
        RECT 5.170 1.180 5.480 1.310 ;
    END
  END INPUT1_3
  OBS
      LAYER li1 ;
        RECT 2.100 4.480 2.420 4.510 ;
        RECT 0.070 4.130 0.240 4.410 ;
        RECT 0.580 4.170 0.930 4.340 ;
        RECT 0.750 4.140 0.930 4.170 ;
        RECT 1.350 4.150 1.520 4.420 ;
        RECT 2.100 4.290 2.430 4.480 ;
        RECT 5.180 4.470 5.500 4.500 ;
        RECT 2.100 4.250 2.420 4.290 ;
        RECT 0.070 4.090 0.280 4.130 ;
        RECT 0.750 4.110 1.070 4.140 ;
        RECT 0.070 4.070 0.300 4.090 ;
        RECT 0.070 4.050 0.330 4.070 ;
        RECT 0.070 4.000 0.410 4.050 ;
        RECT 0.070 3.940 0.560 4.000 ;
        RECT 0.070 3.910 0.580 3.940 ;
        RECT 0.110 3.880 0.580 3.910 ;
        RECT 0.750 3.920 1.080 4.110 ;
        RECT 1.350 3.930 1.550 4.150 ;
        RECT 2.130 4.080 2.300 4.250 ;
        RECT 2.820 4.130 2.990 4.420 ;
        RECT 3.780 4.140 3.950 4.420 ;
        RECT 4.520 4.140 4.690 4.430 ;
        RECT 5.180 4.280 5.510 4.470 ;
        RECT 5.750 4.330 5.940 4.360 ;
        RECT 5.180 4.240 5.500 4.280 ;
        RECT 1.360 3.920 1.550 3.930 ;
        RECT 0.750 3.880 1.070 3.920 ;
        RECT 2.810 3.900 3.000 4.130 ;
        RECT 3.670 4.110 3.990 4.140 ;
        RECT 3.670 3.920 4.000 4.110 ;
        RECT 3.670 3.880 3.990 3.920 ;
        RECT 4.520 3.910 4.710 4.140 ;
        RECT 5.240 4.080 5.410 4.240 ;
        RECT 5.750 4.160 6.190 4.330 ;
        RECT 5.750 4.130 5.940 4.160 ;
        RECT 0.240 3.830 0.580 3.880 ;
        RECT 0.360 3.820 0.580 3.830 ;
        RECT 0.370 3.790 0.580 3.820 ;
        RECT 0.390 3.710 0.580 3.790 ;
        RECT 1.750 3.710 2.080 3.830 ;
        RECT 6.470 3.740 6.640 4.420 ;
        RECT -0.100 3.660 0.070 3.680 ;
        RECT -0.120 3.230 0.090 3.660 ;
        RECT 0.390 3.540 0.910 3.710 ;
        RECT 0.390 3.510 0.580 3.540 ;
        RECT 1.260 3.530 5.480 3.710 ;
        RECT 6.210 3.700 6.640 3.740 ;
        RECT 5.860 3.540 6.640 3.700 ;
        RECT 5.860 3.530 6.400 3.540 ;
        RECT 6.210 3.510 6.400 3.530 ;
        RECT -0.120 2.590 0.090 3.020 ;
        RECT 0.390 2.710 0.580 2.740 ;
        RECT 6.210 2.720 6.400 2.740 ;
        RECT -0.100 2.570 0.070 2.590 ;
        RECT 0.390 2.540 0.910 2.710 ;
        RECT 1.260 2.540 5.480 2.720 ;
        RECT 5.860 2.710 6.400 2.720 ;
        RECT 5.860 2.550 6.640 2.710 ;
        RECT 0.390 2.460 0.580 2.540 ;
        RECT 0.370 2.430 0.580 2.460 ;
        RECT 0.360 2.420 0.580 2.430 ;
        RECT 1.750 2.420 2.080 2.540 ;
        RECT 6.210 2.510 6.640 2.550 ;
        RECT 0.240 2.370 0.580 2.420 ;
        RECT 0.110 2.340 0.580 2.370 ;
        RECT 0.070 2.310 0.580 2.340 ;
        RECT 0.750 2.330 1.070 2.370 ;
        RECT 0.070 2.250 0.560 2.310 ;
        RECT 0.070 2.200 0.410 2.250 ;
        RECT 0.070 2.180 0.330 2.200 ;
        RECT 0.070 2.160 0.300 2.180 ;
        RECT 0.070 2.120 0.280 2.160 ;
        RECT 0.750 2.140 1.080 2.330 ;
        RECT 1.360 2.320 1.550 2.330 ;
        RECT 0.070 1.840 0.240 2.120 ;
        RECT 0.750 2.110 1.070 2.140 ;
        RECT 0.750 2.080 0.930 2.110 ;
        RECT 0.580 1.910 0.930 2.080 ;
        RECT 1.350 2.100 1.550 2.320 ;
        RECT 1.350 1.830 1.520 2.100 ;
        RECT 2.130 2.000 2.300 2.170 ;
        RECT 2.810 2.120 3.000 2.350 ;
        RECT 3.670 2.330 3.990 2.370 ;
        RECT 3.670 2.140 4.000 2.330 ;
        RECT 2.100 1.960 2.420 2.000 ;
        RECT 2.100 1.770 2.430 1.960 ;
        RECT 2.820 1.830 2.990 2.120 ;
        RECT 3.670 2.110 3.990 2.140 ;
        RECT 4.520 2.110 4.710 2.340 ;
        RECT 3.780 1.830 3.950 2.110 ;
        RECT 4.520 1.820 4.690 2.110 ;
        RECT 5.240 2.010 5.410 2.170 ;
        RECT 5.750 2.090 5.940 2.120 ;
        RECT 5.180 1.970 5.500 2.010 ;
        RECT 5.180 1.780 5.510 1.970 ;
        RECT 5.750 1.920 6.190 2.090 ;
        RECT 5.750 1.890 5.940 1.920 ;
        RECT 6.470 1.830 6.640 2.510 ;
        RECT 2.100 1.740 2.420 1.770 ;
        RECT 5.180 1.750 5.500 1.780 ;
        RECT 2.100 1.460 2.420 1.490 ;
        RECT 0.070 1.110 0.240 1.390 ;
        RECT 0.580 1.150 0.930 1.320 ;
        RECT 0.750 1.120 0.930 1.150 ;
        RECT 1.350 1.130 1.520 1.400 ;
        RECT 2.100 1.270 2.430 1.460 ;
        RECT 5.180 1.450 5.500 1.480 ;
        RECT 2.100 1.230 2.420 1.270 ;
        RECT 0.070 1.070 0.280 1.110 ;
        RECT 0.750 1.090 1.070 1.120 ;
        RECT 0.070 1.050 0.300 1.070 ;
        RECT 0.070 1.030 0.330 1.050 ;
        RECT 0.070 0.980 0.410 1.030 ;
        RECT 0.070 0.920 0.560 0.980 ;
        RECT 0.070 0.890 0.580 0.920 ;
        RECT 0.110 0.860 0.580 0.890 ;
        RECT 0.750 0.900 1.080 1.090 ;
        RECT 1.350 0.910 1.550 1.130 ;
        RECT 2.130 1.060 2.300 1.230 ;
        RECT 2.820 1.110 2.990 1.400 ;
        RECT 3.780 1.120 3.950 1.400 ;
        RECT 4.520 1.120 4.690 1.410 ;
        RECT 5.180 1.260 5.510 1.450 ;
        RECT 5.750 1.310 5.940 1.340 ;
        RECT 5.180 1.220 5.500 1.260 ;
        RECT 1.360 0.900 1.550 0.910 ;
        RECT 0.750 0.860 1.070 0.900 ;
        RECT 2.810 0.880 3.000 1.110 ;
        RECT 3.670 1.090 3.990 1.120 ;
        RECT 3.670 0.900 4.000 1.090 ;
        RECT 3.670 0.860 3.990 0.900 ;
        RECT 4.520 0.890 4.710 1.120 ;
        RECT 5.240 1.060 5.410 1.220 ;
        RECT 5.750 1.140 6.190 1.310 ;
        RECT 5.750 1.110 5.940 1.140 ;
        RECT 0.240 0.810 0.580 0.860 ;
        RECT 0.360 0.800 0.580 0.810 ;
        RECT 0.370 0.770 0.580 0.800 ;
        RECT 0.390 0.690 0.580 0.770 ;
        RECT 1.750 0.690 2.080 0.810 ;
        RECT 6.470 0.720 6.640 1.400 ;
        RECT -0.100 0.640 0.070 0.660 ;
        RECT -0.120 0.210 0.090 0.640 ;
        RECT 0.390 0.520 0.910 0.690 ;
        RECT 0.390 0.490 0.580 0.520 ;
        RECT 1.260 0.510 5.480 0.690 ;
        RECT 6.210 0.680 6.640 0.720 ;
        RECT 5.860 0.520 6.640 0.680 ;
        RECT 5.860 0.510 6.400 0.520 ;
        RECT 6.210 0.490 6.400 0.510 ;
        RECT -0.120 -0.430 0.090 0.000 ;
        RECT 0.390 -0.310 0.580 -0.280 ;
        RECT 6.210 -0.300 6.400 -0.280 ;
        RECT -0.100 -0.450 0.070 -0.430 ;
        RECT 0.390 -0.480 0.910 -0.310 ;
        RECT 1.260 -0.480 5.480 -0.300 ;
        RECT 5.860 -0.310 6.400 -0.300 ;
        RECT 5.860 -0.470 6.640 -0.310 ;
        RECT 0.390 -0.560 0.580 -0.480 ;
        RECT 0.370 -0.590 0.580 -0.560 ;
        RECT 0.360 -0.600 0.580 -0.590 ;
        RECT 1.750 -0.600 2.080 -0.480 ;
        RECT 6.210 -0.510 6.640 -0.470 ;
        RECT 0.240 -0.650 0.580 -0.600 ;
        RECT 0.110 -0.680 0.580 -0.650 ;
        RECT 0.070 -0.710 0.580 -0.680 ;
        RECT 0.750 -0.690 1.070 -0.650 ;
        RECT 0.070 -0.770 0.560 -0.710 ;
        RECT 0.070 -0.820 0.410 -0.770 ;
        RECT 0.070 -0.840 0.330 -0.820 ;
        RECT 0.070 -0.860 0.300 -0.840 ;
        RECT 0.070 -0.900 0.280 -0.860 ;
        RECT 0.750 -0.880 1.080 -0.690 ;
        RECT 1.360 -0.700 1.550 -0.690 ;
        RECT 0.070 -1.180 0.240 -0.900 ;
        RECT 0.750 -0.910 1.070 -0.880 ;
        RECT 0.750 -0.940 0.930 -0.910 ;
        RECT 0.580 -1.110 0.930 -0.940 ;
        RECT 1.350 -0.920 1.550 -0.700 ;
        RECT 1.350 -1.190 1.520 -0.920 ;
        RECT 2.130 -1.020 2.300 -0.850 ;
        RECT 2.810 -0.900 3.000 -0.670 ;
        RECT 3.670 -0.690 3.990 -0.650 ;
        RECT 3.670 -0.880 4.000 -0.690 ;
        RECT 2.100 -1.060 2.420 -1.020 ;
        RECT 2.100 -1.250 2.430 -1.060 ;
        RECT 2.820 -1.190 2.990 -0.900 ;
        RECT 3.670 -0.910 3.990 -0.880 ;
        RECT 4.520 -0.910 4.710 -0.680 ;
        RECT 3.780 -1.190 3.950 -0.910 ;
        RECT 4.520 -1.200 4.690 -0.910 ;
        RECT 5.240 -1.010 5.410 -0.850 ;
        RECT 5.750 -0.930 5.940 -0.900 ;
        RECT 5.180 -1.050 5.500 -1.010 ;
        RECT 5.180 -1.240 5.510 -1.050 ;
        RECT 5.750 -1.100 6.190 -0.930 ;
        RECT 5.750 -1.130 5.940 -1.100 ;
        RECT 6.470 -1.190 6.640 -0.510 ;
        RECT 2.100 -1.280 2.420 -1.250 ;
        RECT 5.180 -1.270 5.500 -1.240 ;
      LAYER mcon ;
        RECT 2.160 4.300 2.330 4.470 ;
        RECT 0.810 3.930 0.980 4.100 ;
        RECT 1.370 3.950 1.540 4.120 ;
        RECT 5.240 4.290 5.410 4.460 ;
        RECT 2.820 3.930 2.990 4.100 ;
        RECT 3.730 3.930 3.900 4.100 ;
        RECT 4.530 3.940 4.700 4.110 ;
        RECT 5.760 4.160 5.930 4.330 ;
        RECT -0.100 3.510 0.070 3.680 ;
        RECT 0.400 3.540 0.570 3.710 ;
        RECT 6.220 3.540 6.390 3.710 ;
        RECT 0.400 2.540 0.570 2.710 ;
        RECT 6.220 2.540 6.390 2.710 ;
        RECT 0.810 2.150 0.980 2.320 ;
        RECT 1.370 2.130 1.540 2.300 ;
        RECT 2.820 2.150 2.990 2.320 ;
        RECT 3.730 2.150 3.900 2.320 ;
        RECT 4.530 2.140 4.700 2.310 ;
        RECT 2.160 1.780 2.330 1.950 ;
        RECT 5.240 1.790 5.410 1.960 ;
        RECT 5.760 1.920 5.930 2.090 ;
        RECT 2.160 1.280 2.330 1.450 ;
        RECT 0.810 0.910 0.980 1.080 ;
        RECT 1.370 0.930 1.540 1.100 ;
        RECT 5.240 1.270 5.410 1.440 ;
        RECT 2.820 0.910 2.990 1.080 ;
        RECT 3.730 0.910 3.900 1.080 ;
        RECT 4.530 0.920 4.700 1.090 ;
        RECT 5.760 1.140 5.930 1.310 ;
        RECT -0.100 0.490 0.070 0.660 ;
        RECT 0.400 0.520 0.570 0.690 ;
        RECT 6.220 0.520 6.390 0.690 ;
        RECT 0.400 -0.480 0.570 -0.310 ;
        RECT 6.220 -0.480 6.390 -0.310 ;
        RECT 0.810 -0.870 0.980 -0.700 ;
        RECT 1.370 -0.890 1.540 -0.720 ;
        RECT 2.820 -0.870 2.990 -0.700 ;
        RECT 3.730 -0.870 3.900 -0.700 ;
        RECT 4.530 -0.880 4.700 -0.710 ;
        RECT 2.160 -1.240 2.330 -1.070 ;
        RECT 5.240 -1.230 5.410 -1.060 ;
        RECT 5.760 -1.100 5.930 -0.930 ;
      LAYER met1 ;
        RECT 2.090 4.220 2.410 4.540 ;
        RECT 5.170 4.210 5.490 4.530 ;
        RECT 0.740 3.850 1.060 4.170 ;
        RECT 1.340 3.890 1.570 4.180 ;
        RECT -0.130 3.550 0.100 3.740 ;
        RECT 1.360 3.630 1.530 3.890 ;
        RECT 2.790 3.870 3.020 4.160 ;
        RECT -0.130 3.450 0.220 3.550 ;
        RECT -0.120 3.230 0.220 3.450 ;
        RECT 1.350 3.310 1.610 3.630 ;
        RECT 2.810 3.620 2.980 3.870 ;
        RECT 3.660 3.850 3.980 4.170 ;
        RECT 4.500 3.880 4.730 4.170 ;
        RECT 5.730 4.100 5.960 4.390 ;
        RECT 2.770 3.300 3.030 3.620 ;
        RECT 4.530 3.600 4.700 3.880 ;
        RECT 5.730 3.610 5.920 4.100 ;
        RECT 4.520 3.280 4.780 3.600 ;
        RECT 5.560 3.360 5.920 3.610 ;
        RECT 5.560 3.290 5.820 3.360 ;
        RECT -0.120 2.800 0.220 3.020 ;
        RECT -0.130 2.700 0.220 2.800 ;
        RECT -0.130 2.510 0.100 2.700 ;
        RECT 1.350 2.620 1.610 2.940 ;
        RECT 2.770 2.630 3.030 2.950 ;
        RECT 4.520 2.650 4.780 2.970 ;
        RECT 5.560 2.890 5.820 2.960 ;
        RECT 0.740 2.080 1.060 2.400 ;
        RECT 1.360 2.360 1.530 2.620 ;
        RECT 2.810 2.380 2.980 2.630 ;
        RECT 1.340 2.070 1.570 2.360 ;
        RECT 2.790 2.090 3.020 2.380 ;
        RECT 3.660 2.080 3.980 2.400 ;
        RECT 4.530 2.370 4.700 2.650 ;
        RECT 5.560 2.640 5.920 2.890 ;
        RECT 4.500 2.080 4.730 2.370 ;
        RECT 5.730 2.150 5.920 2.640 ;
        RECT 2.090 1.710 2.410 2.030 ;
        RECT 5.170 1.720 5.490 2.040 ;
        RECT 5.730 1.860 5.960 2.150 ;
        RECT 2.090 1.200 2.410 1.520 ;
        RECT 5.170 1.190 5.490 1.510 ;
        RECT 0.740 0.830 1.060 1.150 ;
        RECT 1.340 0.870 1.570 1.160 ;
        RECT -0.130 0.530 0.100 0.720 ;
        RECT 1.360 0.610 1.530 0.870 ;
        RECT 2.790 0.850 3.020 1.140 ;
        RECT -0.130 0.430 0.220 0.530 ;
        RECT -0.120 0.210 0.220 0.430 ;
        RECT 1.350 0.290 1.610 0.610 ;
        RECT 2.810 0.600 2.980 0.850 ;
        RECT 3.660 0.830 3.980 1.150 ;
        RECT 4.500 0.860 4.730 1.150 ;
        RECT 5.730 1.080 5.960 1.370 ;
        RECT 2.770 0.280 3.030 0.600 ;
        RECT 4.530 0.580 4.700 0.860 ;
        RECT 5.730 0.590 5.920 1.080 ;
        RECT 4.520 0.260 4.780 0.580 ;
        RECT 5.560 0.340 5.920 0.590 ;
        RECT 5.560 0.270 5.820 0.340 ;
        RECT -0.120 -0.220 0.220 0.000 ;
        RECT -0.130 -0.320 0.220 -0.220 ;
        RECT -0.130 -0.510 0.100 -0.320 ;
        RECT 1.350 -0.400 1.610 -0.080 ;
        RECT 2.770 -0.390 3.030 -0.070 ;
        RECT 4.520 -0.370 4.780 -0.050 ;
        RECT 5.560 -0.130 5.820 -0.060 ;
        RECT 0.740 -0.940 1.060 -0.620 ;
        RECT 1.360 -0.660 1.530 -0.400 ;
        RECT 2.810 -0.640 2.980 -0.390 ;
        RECT 1.340 -0.950 1.570 -0.660 ;
        RECT 2.790 -0.930 3.020 -0.640 ;
        RECT 3.660 -0.940 3.980 -0.620 ;
        RECT 4.530 -0.650 4.700 -0.370 ;
        RECT 5.560 -0.380 5.920 -0.130 ;
        RECT 4.500 -0.940 4.730 -0.650 ;
        RECT 5.730 -0.870 5.920 -0.380 ;
        RECT 2.090 -1.310 2.410 -0.990 ;
        RECT 5.170 -1.300 5.490 -0.980 ;
        RECT 5.730 -1.160 5.960 -0.870 ;
      LAYER via ;
        RECT 2.120 4.250 2.380 4.510 ;
        RECT 5.200 4.240 5.460 4.500 ;
        RECT 0.770 3.880 1.030 4.140 ;
        RECT 3.690 3.880 3.950 4.140 ;
        RECT -0.040 3.260 0.220 3.520 ;
        RECT 1.350 3.340 1.610 3.600 ;
        RECT 2.770 3.330 3.030 3.590 ;
        RECT 4.520 3.310 4.780 3.570 ;
        RECT 5.560 3.320 5.820 3.580 ;
        RECT -0.040 2.730 0.220 2.990 ;
        RECT 1.350 2.650 1.610 2.910 ;
        RECT 2.770 2.660 3.030 2.920 ;
        RECT 4.520 2.680 4.780 2.940 ;
        RECT 5.560 2.670 5.820 2.930 ;
        RECT 0.770 2.110 1.030 2.370 ;
        RECT 3.690 2.110 3.950 2.370 ;
        RECT 2.120 1.740 2.380 2.000 ;
        RECT 5.200 1.750 5.460 2.010 ;
        RECT 2.120 1.230 2.380 1.490 ;
        RECT 5.200 1.220 5.460 1.480 ;
        RECT 0.770 0.860 1.030 1.120 ;
        RECT 3.690 0.860 3.950 1.120 ;
        RECT -0.040 0.240 0.220 0.500 ;
        RECT 1.350 0.320 1.610 0.580 ;
        RECT 2.770 0.310 3.030 0.570 ;
        RECT 4.520 0.290 4.780 0.550 ;
        RECT 5.560 0.300 5.820 0.560 ;
        RECT -0.040 -0.290 0.220 -0.030 ;
        RECT 1.350 -0.370 1.610 -0.110 ;
        RECT 2.770 -0.360 3.030 -0.100 ;
        RECT 4.520 -0.340 4.780 -0.080 ;
        RECT 5.560 -0.350 5.820 -0.090 ;
        RECT 0.770 -0.910 1.030 -0.650 ;
        RECT 3.690 -0.910 3.950 -0.650 ;
        RECT 2.120 -1.280 2.380 -1.020 ;
        RECT 5.200 -1.270 5.460 -1.010 ;
  END
END sky130_hilas_Tgate4Double01

MACRO sky130_hilas_cellAttempt01
  CLASS CORE ;
  FOREIGN sky130_hilas_cellAttempt01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VTUN
    ANTENNADIFFAREA 1.978000 ;
    PORT
      LAYER nwell ;
        RECT 0.010 4.190 1.740 6.050 ;
        RECT 0.000 2.350 1.740 4.190 ;
        RECT 0.010 0.000 1.740 2.350 ;
      LAYER met1 ;
        RECT 0.360 0.000 0.760 6.050 ;
    END
  END VTUN
  PIN VINJ
    ANTENNADIFFAREA 1.020000 ;
    PORT
      LAYER nwell ;
        RECT 7.520 6.040 10.070 6.050 ;
        RECT 7.520 0.020 10.080 6.040 ;
        RECT 7.520 0.010 10.070 0.020 ;
      LAYER met1 ;
        RECT 9.560 5.400 9.720 6.050 ;
        RECT 9.450 4.850 9.720 5.400 ;
        RECT 9.450 4.800 9.730 4.850 ;
        RECT 9.560 4.710 9.730 4.800 ;
        RECT 9.560 4.350 9.720 4.710 ;
        RECT 9.560 4.260 9.730 4.350 ;
        RECT 9.450 4.210 9.730 4.260 ;
        RECT 9.450 3.660 9.720 4.210 ;
        RECT 9.560 2.390 9.720 3.660 ;
        RECT 9.450 1.840 9.720 2.390 ;
        RECT 9.450 1.790 9.730 1.840 ;
        RECT 9.560 1.700 9.730 1.790 ;
        RECT 9.560 1.350 9.720 1.700 ;
        RECT 9.560 1.260 9.730 1.350 ;
        RECT 9.450 1.210 9.730 1.260 ;
        RECT 9.450 0.660 9.720 1.210 ;
        RECT 9.560 0.010 9.720 0.660 ;
    END
  END VINJ
  PIN COLSEL1
    ANTENNAGATEAREA 0.620000 ;
    PORT
      LAYER met1 ;
        RECT 9.120 5.060 9.310 6.050 ;
        RECT 9.140 4.940 9.310 5.060 ;
        RECT 9.150 4.120 9.310 4.940 ;
        RECT 9.140 4.000 9.310 4.120 ;
        RECT 9.120 3.140 9.310 4.000 ;
        RECT 9.100 2.910 9.340 3.140 ;
        RECT 9.120 2.050 9.310 2.910 ;
        RECT 9.140 1.930 9.310 2.050 ;
        RECT 9.150 1.120 9.310 1.930 ;
        RECT 9.140 1.000 9.310 1.120 ;
        RECT 9.120 0.010 9.310 1.000 ;
    END
  END COLSEL1
  PIN COL1
    ANTENNADIFFAREA 0.372000 ;
    PORT
      LAYER met1 ;
        RECT 8.750 5.370 8.910 6.050 ;
        RECT 8.750 5.350 8.950 5.370 ;
        RECT 8.730 5.110 8.960 5.350 ;
        RECT 8.750 4.890 8.950 5.110 ;
        RECT 8.750 4.170 8.910 4.890 ;
        RECT 8.750 3.950 8.950 4.170 ;
        RECT 8.730 3.710 8.960 3.950 ;
        RECT 8.750 3.690 8.950 3.710 ;
        RECT 8.750 2.360 8.910 3.690 ;
        RECT 8.750 2.340 8.950 2.360 ;
        RECT 8.730 2.100 8.960 2.340 ;
        RECT 8.750 1.880 8.950 2.100 ;
        RECT 8.750 1.170 8.910 1.880 ;
        RECT 8.750 0.950 8.950 1.170 ;
        RECT 8.730 0.710 8.960 0.950 ;
        RECT 8.750 0.690 8.950 0.710 ;
        RECT 8.750 0.010 8.910 0.690 ;
    END
  END COL1
  PIN GATE1
    ANTENNADIFFAREA 2.743300 ;
    PORT
      LAYER nwell ;
        RECT 3.760 0.000 5.990 6.050 ;
      LAYER met1 ;
        RECT 4.410 4.130 4.790 6.050 ;
        RECT 4.400 2.270 4.790 4.130 ;
        RECT 4.410 0.000 4.790 2.270 ;
    END
  END GATE1
  PIN DRAIN1
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER met2 ;
        RECT 7.610 5.550 7.920 5.690 ;
        RECT 0.010 5.370 10.080 5.550 ;
        RECT 7.610 5.360 7.920 5.370 ;
    END
  END DRAIN1
  PIN ROW3
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 7.610 2.110 7.920 2.130 ;
        RECT 0.020 1.940 10.080 2.110 ;
        RECT 7.520 1.930 10.080 1.940 ;
        RECT 7.610 1.800 7.920 1.930 ;
    END
  END ROW3
  PIN DRAIN2
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER met2 ;
        RECT 7.610 3.690 7.920 3.700 ;
        RECT 0.000 3.510 10.080 3.690 ;
        RECT 7.610 3.370 7.920 3.510 ;
    END
  END DRAIN2
  PIN ROW2
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 7.610 4.120 7.920 4.250 ;
        RECT 0.000 3.940 10.080 4.120 ;
        RECT 7.610 3.920 7.920 3.940 ;
    END
  END ROW2
  PIN DRAIN3
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER met2 ;
        RECT 7.610 2.540 7.920 2.680 ;
        RECT 7.610 2.530 10.080 2.540 ;
        RECT 0.020 2.360 10.080 2.530 ;
        RECT 7.610 2.350 7.920 2.360 ;
    END
  END DRAIN3
  PIN ROW4
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 7.610 1.130 7.920 1.250 ;
        RECT 0.020 1.120 7.920 1.130 ;
        RECT 0.020 0.960 10.080 1.120 ;
        RECT 0.800 0.870 2.340 0.960 ;
        RECT 7.520 0.940 10.080 0.960 ;
        RECT 7.610 0.920 7.920 0.940 ;
    END
  END ROW4
  PIN DRAIN4
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER met2 ;
        RECT 7.610 0.690 7.920 0.700 ;
        RECT 0.020 0.520 10.080 0.690 ;
        RECT 7.610 0.510 10.080 0.520 ;
        RECT 7.610 0.370 7.920 0.510 ;
    END
  END DRAIN4
  PIN ROW1
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 7.610 5.120 7.920 5.140 ;
        RECT 0.010 4.940 10.080 5.120 ;
        RECT 7.610 4.810 7.920 4.940 ;
    END
  END ROW1
  PIN VGND
    ANTENNADIFFAREA 1.012300 ;
    PORT
      LAYER met2 ;
        RECT 2.760 1.560 3.080 1.570 ;
        RECT 6.690 1.560 7.010 1.640 ;
        RECT 2.760 1.380 7.010 1.560 ;
        RECT 2.760 1.310 3.080 1.380 ;
        RECT 6.690 1.320 7.010 1.380 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.730 4.890 6.970 6.050 ;
        RECT 6.710 4.230 6.980 4.890 ;
        RECT 6.730 1.640 6.970 4.230 ;
        RECT 6.720 1.320 6.980 1.640 ;
        RECT 6.730 0.000 6.970 1.320 ;
      LAYER via ;
        RECT 6.720 1.350 6.980 1.610 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.800 4.870 3.040 6.050 ;
        RECT 2.790 4.210 3.050 4.870 ;
        RECT 2.800 1.600 3.040 4.210 ;
        RECT 2.790 1.280 3.050 1.600 ;
        RECT 2.800 0.000 3.040 1.280 ;
      LAYER via ;
        RECT 2.790 1.310 3.050 1.570 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 7.620 5.640 7.940 5.650 ;
        RECT 7.620 5.470 8.200 5.640 ;
        RECT 7.620 5.420 7.950 5.470 ;
        RECT 7.620 5.390 7.940 5.420 ;
        RECT 9.480 5.370 9.680 5.720 ;
        RECT 7.620 5.060 7.940 5.100 ;
        RECT 7.620 5.020 7.950 5.060 ;
        RECT 7.620 4.850 8.200 5.020 ;
        RECT 7.620 4.840 7.940 4.850 ;
        RECT 2.830 4.300 3.000 4.810 ;
        RECT 6.770 4.290 6.940 4.800 ;
        RECT 8.750 4.780 8.950 5.350 ;
        RECT 9.480 5.340 9.690 5.370 ;
        RECT 9.470 4.750 9.690 5.340 ;
        RECT 7.620 4.210 7.940 4.220 ;
        RECT 7.620 4.040 8.200 4.210 ;
        RECT 7.620 4.000 7.950 4.040 ;
        RECT 7.620 3.960 7.940 4.000 ;
        RECT 8.750 3.710 8.950 4.280 ;
        RECT 9.470 3.720 9.690 4.310 ;
        RECT 9.480 3.690 9.690 3.720 ;
        RECT 7.620 3.640 7.940 3.670 ;
        RECT 0.430 2.800 0.980 3.230 ;
        RECT 2.840 2.590 3.010 3.600 ;
        RECT 7.620 3.590 7.950 3.640 ;
        RECT 4.460 2.730 5.010 3.160 ;
        RECT 6.770 2.450 6.940 3.460 ;
        RECT 7.620 3.420 8.200 3.590 ;
        RECT 7.620 3.410 7.940 3.420 ;
        RECT 9.480 3.340 9.680 3.690 ;
        RECT 8.870 2.940 9.310 3.110 ;
        RECT 7.620 2.630 7.940 2.640 ;
        RECT 7.620 2.460 8.200 2.630 ;
        RECT 7.620 2.410 7.950 2.460 ;
        RECT 7.620 2.380 7.940 2.410 ;
        RECT 9.480 2.360 9.680 2.710 ;
        RECT 7.620 2.050 7.940 2.090 ;
        RECT 7.620 2.010 7.950 2.050 ;
        RECT 7.620 1.840 8.200 2.010 ;
        RECT 7.620 1.830 7.940 1.840 ;
        RECT 8.750 1.770 8.950 2.340 ;
        RECT 9.480 2.330 9.690 2.360 ;
        RECT 9.470 1.740 9.690 2.330 ;
        RECT 7.620 1.210 7.940 1.220 ;
        RECT 7.620 1.040 8.200 1.210 ;
        RECT 7.620 1.000 7.950 1.040 ;
        RECT 7.620 0.960 7.940 1.000 ;
        RECT 8.750 0.710 8.950 1.280 ;
        RECT 9.470 0.720 9.690 1.310 ;
        RECT 9.480 0.690 9.690 0.720 ;
        RECT 7.620 0.640 7.940 0.670 ;
        RECT 7.620 0.590 7.950 0.640 ;
        RECT 7.620 0.420 8.200 0.590 ;
        RECT 7.620 0.410 7.940 0.420 ;
        RECT 9.480 0.340 9.680 0.690 ;
      LAYER mcon ;
        RECT 7.680 5.430 7.850 5.600 ;
        RECT 8.760 5.140 8.930 5.310 ;
        RECT 7.680 4.880 7.850 5.050 ;
        RECT 2.830 4.640 3.000 4.810 ;
        RECT 6.770 4.630 6.940 4.800 ;
        RECT 9.490 5.170 9.660 5.340 ;
        RECT 7.680 4.010 7.850 4.180 ;
        RECT 8.760 3.750 8.930 3.920 ;
        RECT 9.490 3.720 9.660 3.890 ;
        RECT 7.680 3.460 7.850 3.630 ;
        RECT 0.430 2.880 0.700 3.150 ;
        RECT 2.840 3.180 3.010 3.350 ;
        RECT 2.840 2.840 3.010 3.010 ;
        RECT 4.460 2.810 4.730 3.080 ;
        RECT 6.770 3.040 6.940 3.210 ;
        RECT 9.130 2.940 9.310 3.110 ;
        RECT 6.770 2.700 6.940 2.870 ;
        RECT 7.680 2.420 7.850 2.590 ;
        RECT 8.760 2.130 8.930 2.300 ;
        RECT 7.680 1.870 7.850 2.040 ;
        RECT 9.490 2.160 9.660 2.330 ;
        RECT 7.680 1.010 7.850 1.180 ;
        RECT 8.760 0.750 8.930 0.920 ;
        RECT 9.490 0.720 9.660 0.890 ;
        RECT 7.680 0.460 7.850 0.630 ;
      LAYER met1 ;
        RECT 7.610 5.360 7.930 5.680 ;
        RECT 7.610 4.810 7.930 5.130 ;
        RECT 7.610 3.930 7.930 4.250 ;
        RECT 7.610 3.380 7.930 3.700 ;
        RECT 7.610 2.350 7.930 2.670 ;
        RECT 7.610 1.800 7.930 2.120 ;
        RECT 7.610 0.930 7.930 1.250 ;
        RECT 7.610 0.380 7.930 0.700 ;
      LAYER via ;
        RECT 7.640 5.390 7.900 5.650 ;
        RECT 7.640 4.840 7.900 5.100 ;
        RECT 7.640 3.960 7.900 4.220 ;
        RECT 7.640 3.410 7.900 3.670 ;
        RECT 7.640 2.380 7.900 2.640 ;
        RECT 7.640 1.830 7.900 2.090 ;
        RECT 7.640 0.960 7.900 1.220 ;
        RECT 7.640 0.410 7.900 0.670 ;
  END
END sky130_hilas_cellAttempt01

MACRO sky130_hilas_StepUpDigital
  CLASS CORE ;
  FOREIGN sky130_hilas_StepUpDigital ;
  ORIGIN 0.000 0.800 ;
  SIZE 8.800 BY 1.590 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 0.000 -0.800 2.510 0.790 ;
        RECT 6.470 -0.800 8.240 0.790 ;
      LAYER li1 ;
        RECT 1.280 0.400 3.510 0.550 ;
        RECT 0.340 0.220 0.670 0.390 ;
        RECT 1.130 0.380 3.510 0.400 ;
        RECT 1.130 0.230 1.730 0.380 ;
        RECT 3.330 0.370 3.510 0.380 ;
        RECT 3.330 0.350 3.970 0.370 ;
        RECT 0.410 -0.240 0.590 0.220 ;
        RECT 2.060 0.030 2.390 0.200 ;
        RECT 3.330 0.180 4.010 0.350 ;
        RECT 4.460 0.320 4.920 0.350 ;
        RECT 6.230 0.320 6.580 0.420 ;
        RECT 4.460 0.180 5.570 0.320 ;
        RECT 3.330 0.120 3.510 0.180 ;
        RECT 4.750 0.150 5.570 0.180 ;
        RECT 5.810 0.150 6.980 0.320 ;
        RECT 7.230 0.150 7.990 0.320 ;
        RECT 2.060 -0.220 2.310 0.030 ;
        RECT 4.750 0.010 5.010 0.150 ;
        RECT 0.410 -0.410 1.370 -0.240 ;
        RECT 1.840 -0.320 2.310 -0.220 ;
        RECT 3.830 -0.160 5.010 0.010 ;
        RECT 7.760 0.140 7.990 0.150 ;
        RECT 1.840 -0.330 2.480 -0.320 ;
        RECT 1.840 -0.390 3.280 -0.330 ;
        RECT 1.920 -0.500 3.280 -0.390 ;
        RECT 3.830 -0.600 4.010 -0.160 ;
        RECT 4.750 -0.300 5.010 -0.160 ;
        RECT 6.220 -0.300 6.550 -0.040 ;
        RECT 7.760 -0.300 8.030 0.140 ;
        RECT 4.250 -0.660 4.460 -0.330 ;
        RECT 4.750 -0.470 5.080 -0.300 ;
        RECT 5.320 -0.470 7.480 -0.300 ;
        RECT 4.750 -0.520 4.920 -0.470 ;
        RECT 7.730 -0.480 8.060 -0.300 ;
        RECT 8.410 -0.440 8.580 -0.380 ;
        RECT 8.390 -0.660 8.610 -0.440 ;
        RECT 8.410 -0.710 8.580 -0.660 ;
      LAYER mcon ;
        RECT 1.450 0.300 1.620 0.470 ;
        RECT 0.410 -0.050 0.580 0.120 ;
        RECT 6.290 0.190 6.500 0.400 ;
        RECT 0.410 -0.400 0.580 -0.230 ;
        RECT 7.800 -0.180 7.970 -0.010 ;
      LAYER met1 ;
        RECT 0.340 -0.800 0.630 0.790 ;
        RECT 1.380 0.250 1.700 0.550 ;
        RECT 4.220 -0.600 4.500 -0.270 ;
        RECT 4.750 -0.800 5.060 0.790 ;
        RECT 6.230 0.150 6.580 0.440 ;
        RECT 6.380 0.130 6.580 0.150 ;
        RECT 7.760 -0.800 8.000 0.790 ;
        RECT 8.330 -0.710 8.740 -0.380 ;
      LAYER via ;
        RECT 1.410 0.260 1.670 0.520 ;
        RECT 4.230 -0.560 4.490 -0.300 ;
        RECT 6.270 0.160 6.530 0.420 ;
        RECT 8.370 -0.680 8.630 -0.420 ;
      LAYER met2 ;
        RECT 1.380 0.470 1.700 0.520 ;
        RECT 0.070 0.270 1.700 0.470 ;
        RECT 1.380 0.260 1.700 0.270 ;
        RECT 4.190 -0.350 4.530 -0.290 ;
        RECT 6.270 -0.350 6.530 0.450 ;
        RECT 4.190 -0.570 6.630 -0.350 ;
        RECT 8.340 -0.710 8.800 -0.390 ;
  END
END sky130_hilas_StepUpDigital

MACRO sky130_hilas_VinjNOR3
  CLASS BLOCK ;
  FOREIGN sky130_hilas_VinjNOR3 ;
  ORIGIN 3.370 -1.440 ;
  SIZE 6.880 BY 1.640 ;
  OBS
      LAYER nwell ;
        RECT -3.360 1.440 0.080 3.080 ;
      LAYER li1 ;
        RECT -2.740 2.650 -2.570 2.790 ;
        RECT -2.010 2.670 -1.840 2.750 ;
        RECT -1.200 2.670 -1.030 2.750 ;
        RECT 0.340 2.710 0.510 2.830 ;
        RECT -2.740 2.480 -2.550 2.650 ;
        RECT -2.740 2.380 -2.570 2.480 ;
        RECT -2.010 2.100 -1.800 2.670 ;
        RECT -1.240 2.420 -1.030 2.670 ;
        RECT -0.640 2.490 -0.470 2.590 ;
        RECT 0.300 2.540 0.510 2.710 ;
        RECT 2.230 2.640 2.490 2.710 ;
        RECT 3.030 2.640 3.210 2.770 ;
        RECT 0.340 2.500 0.510 2.540 ;
        RECT -1.240 2.100 -1.070 2.420 ;
        RECT -0.670 2.320 -0.470 2.490 ;
        RECT -0.640 2.220 -0.470 2.320 ;
        RECT 0.900 2.460 1.770 2.630 ;
        RECT 2.230 2.460 3.210 2.640 ;
        RECT -3.170 2.000 -3.000 2.100 ;
        RECT -3.190 1.830 -3.000 2.000 ;
        RECT -3.170 1.770 -3.000 1.830 ;
        RECT -2.750 2.040 -2.580 2.100 ;
        RECT -2.750 1.770 -2.500 2.040 ;
        RECT -2.010 1.850 -1.760 2.100 ;
        RECT -2.740 1.750 -2.500 1.770 ;
        RECT -1.930 1.760 -1.760 1.850 ;
        RECT -1.280 1.850 -1.070 2.100 ;
        RECT 0.900 2.020 1.070 2.460 ;
        RECT 2.230 2.020 2.490 2.460 ;
        RECT 3.030 2.350 3.210 2.460 ;
        RECT -0.560 1.850 1.070 2.020 ;
        RECT 1.520 1.850 2.490 2.020 ;
        RECT 2.940 1.850 3.280 2.020 ;
        RECT -1.280 1.770 -1.110 1.850 ;
        RECT 0.210 1.810 0.380 1.850 ;
      LAYER mcon ;
        RECT -2.720 2.480 -2.550 2.650 ;
        RECT -2.710 1.800 -2.540 1.970 ;
        RECT 2.260 2.140 2.440 2.320 ;
      LAYER met1 ;
        RECT -2.750 2.700 -2.530 3.040 ;
        RECT -2.750 2.440 -2.520 2.700 ;
        RECT -3.280 1.760 -2.970 2.110 ;
        RECT -2.750 2.040 -2.530 2.440 ;
        RECT -0.730 2.280 -0.400 2.540 ;
        RECT 0.240 2.500 0.670 2.790 ;
        RECT -2.750 1.730 -2.500 2.040 ;
        RECT 0.110 1.750 0.500 2.020 ;
        RECT -2.750 1.530 -2.530 1.730 ;
        RECT 2.220 1.530 2.490 3.050 ;
        RECT 3.040 1.760 3.350 2.080 ;
      LAYER via ;
        RECT -3.250 1.790 -2.990 2.050 ;
        RECT -0.690 2.280 -0.430 2.540 ;
        RECT 0.300 2.530 0.560 2.790 ;
        RECT 0.170 1.750 0.430 2.010 ;
        RECT 3.070 1.790 3.330 2.050 ;
      LAYER met2 ;
        RECT -3.370 2.730 0.670 2.890 ;
        RECT -0.730 2.460 -0.400 2.540 ;
        RECT 0.250 2.500 0.670 2.730 ;
        RECT -1.000 2.440 -0.400 2.460 ;
        RECT -3.360 2.280 -0.400 2.440 ;
        RECT -3.280 1.950 -2.960 2.050 ;
        RECT -3.360 1.790 -2.960 1.950 ;
        RECT 0.130 1.930 0.500 2.010 ;
        RECT 0.130 1.920 1.160 1.930 ;
        RECT 3.040 1.920 3.350 2.080 ;
        RECT 0.130 1.750 3.510 1.920 ;
  END
END sky130_hilas_VinjNOR3

MACRO sky130_hilas_VinjDiodeProtect01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_VinjDiodeProtect01 ;
  ORIGIN 7.450 2.290 ;
  SIZE 28.590 BY 10.870 ;
  PIN OUTPUT 
    ANTENNADIFFAREA 58.900799 ;
    PORT
      LAYER met1 ;
        RECT 6.900 7.960 7.250 8.110 ;
        RECT 6.890 7.010 7.260 7.960 ;
        RECT 5.110 6.640 9.010 7.010 ;
        RECT 5.100 5.180 9.010 6.640 ;
        RECT -4.610 5.170 9.010 5.180 ;
        RECT -5.280 4.610 9.010 5.170 ;
        RECT -5.280 0.310 18.070 4.610 ;
        RECT -5.280 0.030 9.010 0.310 ;
        RECT 5.100 -1.520 9.010 0.030 ;
        RECT 5.080 -2.290 9.030 -1.520 ;
    END
  END OUTPUT 
  PIN VGND
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met2 ;
        RECT -7.450 5.090 21.140 6.490 ;
        RECT -6.980 5.080 -6.050 5.090 ;
        RECT -6.730 3.970 -6.560 5.080 ;
    END
    PORT
      LAYER met1 ;
        RECT -7.010 5.840 -4.640 6.470 ;
        RECT 16.330 5.990 20.460 6.390 ;
        RECT 16.330 5.900 20.470 5.990 ;
        RECT -6.980 3.880 -6.030 5.840 ;
        RECT -5.280 5.820 -4.700 5.840 ;
        RECT 19.940 5.000 20.470 5.900 ;
        RECT -6.750 -1.790 -6.030 3.880 ;
      LAYER via ;
        RECT -6.790 5.990 -4.760 6.320 ;
        RECT 16.600 5.990 19.590 6.340 ;
        RECT -6.850 5.130 -6.150 5.750 ;
        RECT 20.030 5.190 20.380 5.950 ;
    END
  END VGND
  PIN VINJ
    ANTENNADIFFAREA 9.088799 ;
    PORT
      LAYER nwell ;
        RECT 7.420 -0.380 19.470 5.560 ;
      LAYER met2 ;
        RECT 18.890 0.190 19.530 3.200 ;
        RECT -7.450 -1.210 21.140 0.190 ;
        RECT 17.990 -1.340 20.620 -1.210 ;
        RECT 17.990 -1.850 20.540 -1.340 ;
        RECT 17.990 -1.920 18.610 -1.850 ;
    END
  END VINJ
  PIN INPUT
    PORT
      LAYER met1 ;
        RECT 0.260 7.990 4.160 8.580 ;
        RECT 0.260 6.640 0.550 7.990 ;
    END
  END INPUT
  OBS
      LAYER li1 ;
        RECT 0.280 6.640 0.530 8.100 ;
        RECT 0.320 6.630 0.490 6.640 ;
        RECT 6.960 6.610 7.210 8.080 ;
        RECT -6.900 5.890 20.480 6.400 ;
        RECT -6.900 3.960 -6.100 5.890 ;
        RECT -5.520 5.440 -5.350 5.520 ;
        RECT 5.720 5.440 5.950 5.530 ;
        RECT -5.520 5.430 5.950 5.440 ;
        RECT -6.900 -0.620 -6.390 3.960 ;
        RECT -5.530 -0.040 5.950 5.430 ;
        RECT -5.600 -0.210 5.950 -0.040 ;
        RECT -5.530 -0.270 -5.340 -0.210 ;
        RECT 5.720 -0.450 5.950 -0.210 ;
        RECT -5.650 -0.620 -3.850 -0.610 ;
        RECT 6.510 -0.620 7.020 5.890 ;
        RECT 7.780 5.000 19.030 5.170 ;
        RECT 7.780 0.130 7.950 5.000 ;
        RECT 8.340 4.670 18.450 4.690 ;
        RECT 8.340 4.630 18.470 4.670 ;
        RECT 8.290 4.460 18.470 4.630 ;
        RECT 8.340 0.440 18.470 4.460 ;
        RECT 18.860 3.240 19.030 5.000 ;
        RECT 8.340 0.360 18.450 0.440 ;
        RECT 7.770 0.060 7.950 0.130 ;
        RECT 18.860 0.060 19.470 3.240 ;
        RECT 7.770 -0.110 19.470 0.060 ;
        RECT 18.930 -0.220 19.470 -0.110 ;
        RECT 19.930 -0.460 20.480 5.890 ;
        RECT 19.920 -0.620 20.480 -0.460 ;
        RECT -6.900 -0.960 20.480 -0.620 ;
        RECT -6.870 -1.130 20.480 -0.960 ;
        RECT -6.870 -1.150 -6.180 -1.130 ;
        RECT -5.670 -1.140 -3.870 -1.130 ;
      LAYER mcon ;
        RECT 0.320 7.900 0.490 8.070 ;
        RECT 0.320 7.560 0.490 7.730 ;
        RECT 0.320 7.220 0.490 7.390 ;
        RECT 0.320 6.880 0.490 7.050 ;
        RECT 7.000 7.880 7.170 8.050 ;
        RECT 7.000 7.540 7.170 7.710 ;
        RECT 7.000 7.200 7.170 7.370 ;
        RECT 7.000 6.860 7.170 7.030 ;
        RECT -6.820 6.230 -4.960 6.240 ;
        RECT -6.820 6.060 -4.950 6.230 ;
        RECT 16.540 6.050 19.700 6.230 ;
        RECT -6.740 5.100 -6.560 5.890 ;
        RECT -6.730 3.970 -6.560 5.100 ;
        RECT -6.380 3.960 -6.200 5.880 ;
        RECT -5.190 4.930 5.790 5.100 ;
        RECT -5.190 4.310 5.790 4.480 ;
        RECT -5.180 3.690 5.800 3.860 ;
        RECT -5.160 3.110 5.820 3.280 ;
        RECT -5.150 2.520 5.830 2.690 ;
        RECT -5.150 1.920 5.830 2.090 ;
        RECT -5.200 1.320 5.780 1.490 ;
        RECT -5.190 0.710 5.790 0.880 ;
        RECT -5.200 0.110 5.780 0.280 ;
        RECT 8.540 4.170 17.990 4.340 ;
        RECT 8.530 3.420 17.920 3.590 ;
        RECT 8.560 2.700 17.960 2.870 ;
        RECT 8.570 2.040 17.940 2.210 ;
        RECT 8.560 1.390 18.010 1.560 ;
        RECT 8.570 0.750 17.960 0.920 ;
        RECT 20.110 5.070 20.310 6.000 ;
        RECT 19.040 -0.170 19.390 3.130 ;
      LAYER met1 ;
        RECT 18.840 3.190 19.410 3.200 ;
        RECT 18.840 -0.230 19.460 3.190 ;
        RECT 18.840 -0.240 19.410 -0.230 ;
        RECT 18.010 -1.870 18.570 -1.370 ;
        RECT 18.020 -2.090 18.570 -1.870 ;
      LAYER via ;
        RECT 19.000 -0.100 19.420 3.070 ;
        RECT 18.030 -1.920 18.550 -1.400 ;
  END
END sky130_hilas_VinjDiodeProtect01

MACRO sky130_hilas_LevelShift4InputUp
  CLASS CORE ;
  FOREIGN sky130_hilas_LevelShift4InputUp ;
  ORIGIN 0.190 0.400 ;
  SIZE 8.990 BY 6.640 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN INPUT1
    PORT
      LAYER met2 ;
        RECT 8.710 4.740 8.800 5.060 ;
    END
  END INPUT1
  PIN INPUT2
    PORT
      LAYER met2 ;
        RECT 8.710 3.190 8.800 3.510 ;
    END
  END INPUT2
  PIN INPUT3
    PORT
      LAYER met2 ;
        RECT 8.710 1.640 8.800 1.960 ;
    END
  END INPUT3
  PIN INPUT4
    PORT
      LAYER met2 ;
        RECT 8.710 0.090 8.800 0.410 ;
    END
  END INPUT4
  PIN VPWR
    PORT
      LAYER met1 ;
        RECT 7.760 6.190 8.000 6.240 ;
    END
    PORT
      LAYER nwell ;
        RECT 6.280 -0.400 8.050 5.840 ;
      LAYER met1 ;
        RECT 7.570 0.050 7.810 5.840 ;
        RECT 7.570 0.000 8.000 0.050 ;
        RECT 7.570 -0.400 7.810 0.000 ;
    END
  END VPWR
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 0.340 6.190 0.630 6.240 ;
    END
    PORT
      LAYER nwell ;
        RECT -0.190 -0.400 2.320 5.840 ;
      LAYER met1 ;
        RECT 0.150 0.050 0.440 5.840 ;
        RECT 0.150 0.000 0.630 0.050 ;
        RECT 0.150 -0.400 0.440 0.000 ;
    END
  END VINJ
  PIN OUTPUT1
    PORT
      LAYER met2 ;
        RECT 0.000 5.720 0.110 5.920 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    PORT
      LAYER met2 ;
        RECT 0.000 4.170 0.110 4.370 ;
    END
  END OUTPUT2
  PIN OUTPUT3
    PORT
      LAYER met2 ;
        RECT 0.000 2.620 0.110 2.820 ;
    END
  END OUTPUT3
  PIN OUTPUT4
    PORT
      LAYER met2 ;
        RECT 0.000 1.070 0.110 1.270 ;
    END
  END OUTPUT4
  PIN VGND
    PORT
      LAYER met1 ;
        RECT 4.750 6.170 5.060 6.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.560 0.060 4.870 5.840 ;
        RECT 4.560 0.000 5.060 0.060 ;
        RECT 4.560 -0.400 4.870 0.000 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.090 5.450 3.320 5.600 ;
        RECT 0.150 5.270 0.480 5.440 ;
        RECT 0.940 5.430 3.320 5.450 ;
        RECT 0.940 5.280 1.540 5.430 ;
        RECT 3.140 5.420 3.320 5.430 ;
        RECT 3.140 5.400 3.780 5.420 ;
        RECT 0.220 4.810 0.400 5.270 ;
        RECT 1.870 5.080 2.200 5.250 ;
        RECT 3.140 5.230 3.820 5.400 ;
        RECT 4.270 5.370 4.730 5.400 ;
        RECT 6.040 5.370 6.390 5.470 ;
        RECT 4.270 5.230 5.380 5.370 ;
        RECT 3.140 5.170 3.320 5.230 ;
        RECT 4.560 5.200 5.380 5.230 ;
        RECT 5.620 5.200 6.790 5.370 ;
        RECT 7.040 5.200 7.800 5.370 ;
        RECT 1.870 4.830 2.120 5.080 ;
        RECT 4.560 5.060 4.820 5.200 ;
        RECT 0.220 4.640 1.180 4.810 ;
        RECT 1.650 4.730 2.120 4.830 ;
        RECT 3.640 4.890 4.820 5.060 ;
        RECT 7.570 5.190 7.800 5.200 ;
        RECT 1.650 4.720 2.290 4.730 ;
        RECT 1.650 4.660 3.090 4.720 ;
        RECT 1.730 4.550 3.090 4.660 ;
        RECT 3.640 4.450 3.820 4.890 ;
        RECT 4.560 4.750 4.820 4.890 ;
        RECT 6.030 4.750 6.360 5.010 ;
        RECT 7.570 4.750 7.840 5.190 ;
        RECT 4.060 4.390 4.270 4.720 ;
        RECT 4.560 4.580 4.890 4.750 ;
        RECT 5.130 4.580 7.290 4.750 ;
        RECT 4.560 4.530 4.730 4.580 ;
        RECT 7.540 4.570 7.870 4.750 ;
        RECT 8.220 4.610 8.390 4.670 ;
        RECT 8.200 4.390 8.420 4.610 ;
        RECT 8.220 4.340 8.390 4.390 ;
        RECT 1.090 3.900 3.320 4.050 ;
        RECT 0.150 3.720 0.480 3.890 ;
        RECT 0.940 3.880 3.320 3.900 ;
        RECT 0.940 3.730 1.540 3.880 ;
        RECT 3.140 3.870 3.320 3.880 ;
        RECT 3.140 3.850 3.780 3.870 ;
        RECT 0.220 3.260 0.400 3.720 ;
        RECT 1.870 3.530 2.200 3.700 ;
        RECT 3.140 3.680 3.820 3.850 ;
        RECT 4.270 3.820 4.730 3.850 ;
        RECT 6.040 3.820 6.390 3.920 ;
        RECT 4.270 3.680 5.380 3.820 ;
        RECT 3.140 3.620 3.320 3.680 ;
        RECT 4.560 3.650 5.380 3.680 ;
        RECT 5.620 3.650 6.790 3.820 ;
        RECT 7.040 3.650 7.800 3.820 ;
        RECT 1.870 3.280 2.120 3.530 ;
        RECT 4.560 3.510 4.820 3.650 ;
        RECT 0.220 3.090 1.180 3.260 ;
        RECT 1.650 3.180 2.120 3.280 ;
        RECT 3.640 3.340 4.820 3.510 ;
        RECT 7.570 3.640 7.800 3.650 ;
        RECT 1.650 3.170 2.290 3.180 ;
        RECT 1.650 3.110 3.090 3.170 ;
        RECT 1.730 3.000 3.090 3.110 ;
        RECT 3.640 2.900 3.820 3.340 ;
        RECT 4.560 3.200 4.820 3.340 ;
        RECT 6.030 3.200 6.360 3.460 ;
        RECT 7.570 3.200 7.840 3.640 ;
        RECT 4.060 2.840 4.270 3.170 ;
        RECT 4.560 3.030 4.890 3.200 ;
        RECT 5.130 3.030 7.290 3.200 ;
        RECT 4.560 2.980 4.730 3.030 ;
        RECT 7.540 3.020 7.870 3.200 ;
        RECT 8.220 3.060 8.390 3.120 ;
        RECT 8.200 2.840 8.420 3.060 ;
        RECT 8.220 2.790 8.390 2.840 ;
        RECT 1.090 2.350 3.320 2.500 ;
        RECT 0.150 2.170 0.480 2.340 ;
        RECT 0.940 2.330 3.320 2.350 ;
        RECT 0.940 2.180 1.540 2.330 ;
        RECT 3.140 2.320 3.320 2.330 ;
        RECT 3.140 2.300 3.780 2.320 ;
        RECT 0.220 1.710 0.400 2.170 ;
        RECT 1.870 1.980 2.200 2.150 ;
        RECT 3.140 2.130 3.820 2.300 ;
        RECT 4.270 2.270 4.730 2.300 ;
        RECT 6.040 2.270 6.390 2.370 ;
        RECT 4.270 2.130 5.380 2.270 ;
        RECT 3.140 2.070 3.320 2.130 ;
        RECT 4.560 2.100 5.380 2.130 ;
        RECT 5.620 2.100 6.790 2.270 ;
        RECT 7.040 2.100 7.800 2.270 ;
        RECT 1.870 1.730 2.120 1.980 ;
        RECT 4.560 1.960 4.820 2.100 ;
        RECT 0.220 1.540 1.180 1.710 ;
        RECT 1.650 1.630 2.120 1.730 ;
        RECT 3.640 1.790 4.820 1.960 ;
        RECT 7.570 2.090 7.800 2.100 ;
        RECT 1.650 1.620 2.290 1.630 ;
        RECT 1.650 1.560 3.090 1.620 ;
        RECT 1.730 1.450 3.090 1.560 ;
        RECT 3.640 1.350 3.820 1.790 ;
        RECT 4.560 1.650 4.820 1.790 ;
        RECT 6.030 1.650 6.360 1.910 ;
        RECT 7.570 1.650 7.840 2.090 ;
        RECT 4.060 1.290 4.270 1.620 ;
        RECT 4.560 1.480 4.890 1.650 ;
        RECT 5.130 1.480 7.290 1.650 ;
        RECT 4.560 1.430 4.730 1.480 ;
        RECT 7.540 1.470 7.870 1.650 ;
        RECT 8.220 1.510 8.390 1.570 ;
        RECT 8.200 1.290 8.420 1.510 ;
        RECT 8.220 1.240 8.390 1.290 ;
        RECT 1.090 0.800 3.320 0.950 ;
        RECT 0.150 0.620 0.480 0.790 ;
        RECT 0.940 0.780 3.320 0.800 ;
        RECT 0.940 0.630 1.540 0.780 ;
        RECT 3.140 0.770 3.320 0.780 ;
        RECT 3.140 0.750 3.780 0.770 ;
        RECT 0.220 0.160 0.400 0.620 ;
        RECT 1.870 0.430 2.200 0.600 ;
        RECT 3.140 0.580 3.820 0.750 ;
        RECT 4.270 0.720 4.730 0.750 ;
        RECT 6.040 0.720 6.390 0.820 ;
        RECT 4.270 0.580 5.380 0.720 ;
        RECT 3.140 0.520 3.320 0.580 ;
        RECT 4.560 0.550 5.380 0.580 ;
        RECT 5.620 0.550 6.790 0.720 ;
        RECT 7.040 0.550 7.800 0.720 ;
        RECT 1.870 0.180 2.120 0.430 ;
        RECT 4.560 0.410 4.820 0.550 ;
        RECT 0.220 -0.010 1.180 0.160 ;
        RECT 1.650 0.080 2.120 0.180 ;
        RECT 3.640 0.240 4.820 0.410 ;
        RECT 7.570 0.540 7.800 0.550 ;
        RECT 1.650 0.070 2.290 0.080 ;
        RECT 1.650 0.010 3.090 0.070 ;
        RECT 1.730 -0.100 3.090 0.010 ;
        RECT 3.640 -0.200 3.820 0.240 ;
        RECT 4.560 0.100 4.820 0.240 ;
        RECT 6.030 0.100 6.360 0.360 ;
        RECT 7.570 0.100 7.840 0.540 ;
        RECT 4.060 -0.260 4.270 0.070 ;
        RECT 4.560 -0.070 4.890 0.100 ;
        RECT 5.130 -0.070 7.290 0.100 ;
        RECT 4.560 -0.120 4.730 -0.070 ;
        RECT 7.540 -0.080 7.870 0.100 ;
        RECT 8.220 -0.040 8.390 0.020 ;
        RECT 8.200 -0.260 8.420 -0.040 ;
        RECT 8.220 -0.310 8.390 -0.260 ;
      LAYER mcon ;
        RECT 1.260 5.350 1.430 5.520 ;
        RECT 0.220 5.000 0.390 5.170 ;
        RECT 6.100 5.240 6.310 5.450 ;
        RECT 0.220 4.650 0.390 4.820 ;
        RECT 7.610 4.870 7.780 5.040 ;
        RECT 1.260 3.800 1.430 3.970 ;
        RECT 0.220 3.450 0.390 3.620 ;
        RECT 6.100 3.690 6.310 3.900 ;
        RECT 0.220 3.100 0.390 3.270 ;
        RECT 7.610 3.320 7.780 3.490 ;
        RECT 1.260 2.250 1.430 2.420 ;
        RECT 0.220 1.900 0.390 2.070 ;
        RECT 6.100 2.140 6.310 2.350 ;
        RECT 0.220 1.550 0.390 1.720 ;
        RECT 7.610 1.770 7.780 1.940 ;
        RECT 1.260 0.700 1.430 0.870 ;
        RECT 0.220 0.350 0.390 0.520 ;
        RECT 6.100 0.590 6.310 0.800 ;
        RECT 0.220 0.000 0.390 0.170 ;
        RECT 7.610 0.220 7.780 0.390 ;
      LAYER met1 ;
        RECT 1.190 5.300 1.510 5.600 ;
        RECT 6.040 5.200 6.390 5.490 ;
        RECT 6.190 5.180 6.390 5.200 ;
        RECT 4.030 4.450 4.310 4.780 ;
        RECT 8.140 4.340 8.550 4.670 ;
        RECT 1.190 3.750 1.510 4.050 ;
        RECT 6.040 3.650 6.390 3.940 ;
        RECT 6.190 3.630 6.390 3.650 ;
        RECT 4.030 2.900 4.310 3.230 ;
        RECT 8.140 2.790 8.550 3.120 ;
        RECT 1.190 2.200 1.510 2.500 ;
        RECT 6.040 2.100 6.390 2.390 ;
        RECT 6.190 2.080 6.390 2.100 ;
        RECT 4.030 1.350 4.310 1.680 ;
        RECT 8.140 1.240 8.550 1.570 ;
        RECT 1.190 0.650 1.510 0.950 ;
        RECT 6.040 0.550 6.390 0.840 ;
        RECT 6.190 0.530 6.390 0.550 ;
        RECT 4.030 -0.200 4.310 0.130 ;
        RECT 8.140 -0.310 8.550 0.020 ;
      LAYER via ;
        RECT 1.220 5.310 1.480 5.570 ;
        RECT 6.080 5.210 6.340 5.470 ;
        RECT 4.040 4.490 4.300 4.750 ;
        RECT 8.180 4.370 8.440 4.630 ;
        RECT 1.220 3.760 1.480 4.020 ;
        RECT 6.080 3.660 6.340 3.920 ;
        RECT 4.040 2.940 4.300 3.200 ;
        RECT 8.180 2.820 8.440 3.080 ;
        RECT 1.220 2.210 1.480 2.470 ;
        RECT 6.080 2.110 6.340 2.370 ;
        RECT 4.040 1.390 4.300 1.650 ;
        RECT 8.180 1.270 8.440 1.530 ;
        RECT 1.220 0.660 1.480 0.920 ;
        RECT 6.080 0.560 6.340 0.820 ;
        RECT 4.040 -0.160 4.300 0.100 ;
        RECT 8.180 -0.280 8.440 -0.020 ;
      LAYER met2 ;
        RECT 1.190 5.520 1.510 5.570 ;
        RECT -0.120 5.320 1.510 5.520 ;
        RECT 1.190 5.310 1.510 5.320 ;
        RECT 4.000 4.700 4.340 4.760 ;
        RECT 6.080 4.700 6.340 5.500 ;
        RECT 4.000 4.480 6.440 4.700 ;
        RECT 8.150 4.340 8.610 4.660 ;
        RECT 1.190 3.970 1.510 4.020 ;
        RECT -0.120 3.770 1.510 3.970 ;
        RECT 1.190 3.760 1.510 3.770 ;
        RECT 4.000 3.150 4.340 3.210 ;
        RECT 6.080 3.150 6.340 3.950 ;
        RECT 4.000 2.930 6.440 3.150 ;
        RECT 8.150 2.790 8.610 3.110 ;
        RECT 1.190 2.420 1.510 2.470 ;
        RECT -0.120 2.220 1.510 2.420 ;
        RECT 1.190 2.210 1.510 2.220 ;
        RECT 4.000 1.600 4.340 1.660 ;
        RECT 6.080 1.600 6.340 2.400 ;
        RECT 4.000 1.380 6.440 1.600 ;
        RECT 8.150 1.240 8.610 1.560 ;
        RECT 1.190 0.870 1.510 0.920 ;
        RECT -0.120 0.670 1.510 0.870 ;
        RECT 1.190 0.660 1.510 0.670 ;
        RECT 4.000 0.050 4.340 0.110 ;
        RECT 6.080 0.050 6.340 0.850 ;
        RECT 4.000 -0.170 6.440 0.050 ;
        RECT 8.150 -0.310 8.610 0.010 ;
  END
END sky130_hilas_LevelShift4InputUp

MACRO sky130_hilas_WTA4Stage01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_WTA4Stage01 ;
  ORIGIN 13.280 0.430 ;
  SIZE 16.240 BY 9.870 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 2.510 1.160 2.840 1.250 ;
        RECT -3.840 0.990 2.840 1.160 ;
        RECT 2.510 0.960 2.840 0.990 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.570 1.270 2.800 5.620 ;
        RECT 2.530 1.260 2.810 1.270 ;
        RECT 2.530 0.940 2.830 1.260 ;
        RECT 2.570 -0.430 2.800 0.940 ;
      LAYER via ;
        RECT 2.540 0.970 2.810 1.240 ;
    END
  END VGND
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT -0.540 4.570 -0.500 4.660 ;
        RECT -0.650 4.480 0.560 4.570 ;
        RECT -0.650 4.420 0.690 4.480 ;
        RECT -0.650 4.370 2.960 4.420 ;
        RECT 0.380 4.260 2.960 4.370 ;
        RECT 0.380 4.150 0.690 4.260 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT -0.550 3.600 0.660 3.710 ;
        RECT -0.550 3.510 0.690 3.600 ;
        RECT 0.380 3.490 0.690 3.510 ;
        RECT 0.380 3.330 2.960 3.490 ;
        RECT 0.380 3.270 0.690 3.330 ;
    END
  END OUTPUT2
  PIN OUTPUT3
    USE ANALOG ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 0.380 1.680 0.690 1.710 ;
        RECT -0.560 1.650 0.690 1.680 ;
        RECT -0.560 1.520 2.960 1.650 ;
        RECT 0.380 1.490 2.960 1.520 ;
        RECT 0.380 1.380 0.690 1.490 ;
    END
  END OUTPUT3
  PIN OUTPUT4
    USE ANALOG ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 0.380 0.720 0.690 0.830 ;
        RECT 0.380 0.710 2.960 0.720 ;
        RECT -0.550 0.560 2.960 0.710 ;
        RECT -0.550 0.530 0.690 0.560 ;
        RECT 0.380 0.500 0.690 0.530 ;
    END
  END OUTPUT4
  PIN INPUT1
    USE ANALOG ;
    ANTENNAGATEAREA 0.236000 ;
    ANTENNADIFFAREA 4.378700 ;
    PORT
      LAYER nwell ;
        RECT -13.260 9.430 -10.710 9.440 ;
        RECT -13.270 5.620 -10.710 9.430 ;
        RECT -9.180 5.620 -6.950 9.440 ;
        RECT -13.270 5.610 -6.950 5.620 ;
        RECT -13.270 5.460 -10.600 5.610 ;
        RECT -13.270 5.450 -10.420 5.460 ;
        RECT -13.270 3.410 -10.600 5.450 ;
        RECT -13.260 3.400 -10.600 3.410 ;
        RECT -11.120 2.540 -10.600 3.400 ;
        RECT -9.180 3.390 -6.950 5.610 ;
        RECT -11.010 -0.420 -10.600 2.540 ;
      LAYER met2 ;
        RECT -11.110 5.500 -10.800 5.520 ;
        RECT -13.270 5.340 -3.200 5.500 ;
        RECT -13.270 5.330 -3.210 5.340 ;
        RECT -13.270 5.320 -10.710 5.330 ;
        RECT -11.110 5.190 -10.800 5.320 ;
        RECT -7.850 5.310 -7.530 5.330 ;
        RECT -7.850 5.120 0.070 5.310 ;
        RECT 0.230 5.120 0.540 5.160 ;
        RECT -7.850 5.100 0.540 5.120 ;
        RECT -7.850 5.070 -7.530 5.100 ;
        RECT -0.140 4.910 0.540 5.100 ;
        RECT 0.230 4.830 0.540 4.910 ;
        RECT -11.120 4.640 -10.970 4.690 ;
        RECT -11.120 4.520 -10.800 4.640 ;
        RECT -11.120 4.510 -3.200 4.520 ;
        RECT -13.270 4.350 -3.200 4.510 ;
        RECT -13.270 4.330 -10.710 4.350 ;
        RECT -11.120 4.310 -10.800 4.330 ;
        RECT -11.120 4.180 -10.970 4.310 ;
        RECT -7.870 4.180 -7.550 4.280 ;
        RECT -5.530 4.260 -3.990 4.350 ;
        RECT -11.120 4.080 -7.550 4.180 ;
        RECT -13.270 4.020 -7.550 4.080 ;
        RECT -13.270 3.910 -10.700 4.020 ;
        RECT -13.270 3.900 -10.800 3.910 ;
        RECT -11.110 3.780 -10.800 3.900 ;
        RECT -11.140 3.760 -10.800 3.780 ;
        RECT -11.140 3.520 -10.820 3.760 ;
        RECT -11.070 3.510 -10.900 3.520 ;
        RECT -7.910 3.040 -7.680 3.050 ;
        RECT -7.910 3.010 -0.340 3.040 ;
        RECT -7.910 2.840 -0.280 3.010 ;
        RECT 0.230 2.840 0.540 2.920 ;
        RECT -11.160 2.740 -10.840 2.770 ;
        RECT -7.910 2.740 -7.670 2.840 ;
        RECT -11.160 2.560 -7.670 2.740 ;
        RECT -0.470 2.640 0.540 2.840 ;
        RECT 0.130 2.630 0.540 2.640 ;
        RECT 0.230 2.590 0.540 2.630 ;
        RECT -11.160 2.540 -7.750 2.560 ;
        RECT -11.160 2.510 -10.840 2.540 ;
    END
  END INPUT1
  PIN INPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER met1 ;
        RECT -11.120 3.770 -10.800 4.090 ;
        RECT -11.110 3.690 -10.850 3.770 ;
        RECT -11.120 3.490 -10.850 3.690 ;
        RECT -11.120 2.800 -10.910 3.490 ;
        RECT -11.130 2.480 -10.870 2.800 ;
      LAYER via ;
        RECT -11.090 3.800 -10.830 4.060 ;
        RECT -11.110 3.520 -10.850 3.780 ;
        RECT -11.130 2.510 -10.870 2.770 ;
    END
  END INPUT2
  PIN INPUT3
    USE ANALOG ;
    ANTENNAGATEAREA 0.118000 ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT -7.870 2.360 -7.550 2.400 ;
        RECT -7.870 2.340 -0.320 2.360 ;
        RECT 0.230 2.350 0.540 2.390 ;
        RECT 0.130 2.340 0.540 2.350 ;
        RECT -7.870 2.140 0.540 2.340 ;
        RECT -7.770 2.130 -7.450 2.140 ;
        RECT 0.230 2.060 0.540 2.140 ;
        RECT -11.180 1.180 -10.980 1.680 ;
        RECT -8.030 1.180 -7.710 1.220 ;
        RECT -11.180 0.980 -7.630 1.180 ;
        RECT -8.030 0.960 -7.710 0.980 ;
    END
  END INPUT3
  PIN INPUT4
    USE ANALOG ;
    ANTENNAGATEAREA 0.118000 ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT -11.210 0.440 -10.900 0.770 ;
        RECT 0.230 0.090 0.540 0.150 ;
        RECT -0.320 0.080 0.540 0.090 ;
        RECT -11.160 -0.200 -10.850 -0.080 ;
        RECT -7.900 -0.140 0.540 0.080 ;
        RECT -7.900 -0.150 -0.310 -0.140 ;
        RECT -7.900 -0.160 -7.130 -0.150 ;
        RECT -7.900 -0.200 -7.660 -0.160 ;
        RECT 0.230 -0.180 0.540 -0.140 ;
        RECT -11.160 -0.400 -7.660 -0.200 ;
        RECT -11.160 -0.410 -8.470 -0.400 ;
    END
  END INPUT4
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT -11.160 4.940 -10.610 5.120 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT -11.180 3.080 -10.610 3.260 ;
    END
  END DRAIN2
  PIN DRAIN3
    PORT
      LAYER met2 ;
        RECT -11.160 1.930 -10.610 2.110 ;
        RECT -11.160 1.920 -11.000 1.930 ;
    END
  END DRAIN3
  PIN DRAIN4
    PORT
      LAYER met2 ;
        RECT -11.140 0.260 -10.980 0.270 ;
        RECT -11.140 0.080 -10.610 0.260 ;
    END
  END DRAIN4
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT -5.320 5.520 -4.940 5.620 ;
    END
  END GATE1
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT -1.290 5.480 -0.890 5.620 ;
    END
  END VTUN
  PIN WTAMIDDLENODE
    ANTENNAGATEAREA 0.472000 ;
    ANTENNADIFFAREA 0.708000 ;
    PORT
      LAYER met1 ;
        RECT 1.310 -0.430 1.540 5.620 ;
    END
  END WTAMIDDLENODE
  PIN COLSEL1
    ANTENNADIFFAREA 1.053100 ;
    PORT
      LAYER met2 ;
        RECT -10.080 4.910 -9.760 4.970 ;
        RECT -6.060 4.910 -5.730 4.940 ;
        RECT -10.080 4.740 -5.730 4.910 ;
        RECT -10.080 4.690 -9.760 4.740 ;
        RECT -6.060 4.680 -5.730 4.740 ;
    END
  END COLSEL1
  PIN VPWR
    PORT
      LAYER met1 ;
        RECT -9.440 5.550 -9.280 5.620 ;
    END
  END VPWR
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT -10.250 5.550 -10.090 5.620 ;
    END
  END VINJ
  OBS
      LAYER nwell ;
        RECT -4.930 8.810 -3.200 9.440 ;
        RECT -4.930 5.740 -3.190 8.810 ;
        RECT -5.320 5.520 -4.940 5.620 ;
        RECT -4.930 3.390 -3.200 5.740 ;
        RECT -1.290 5.480 -0.890 5.620 ;
      LAYER li1 ;
        RECT -12.870 8.760 -12.670 9.110 ;
        RECT -11.130 9.030 -10.810 9.040 ;
        RECT -11.390 8.860 -10.810 9.030 ;
        RECT -11.140 8.810 -10.810 8.860 ;
        RECT -11.130 8.780 -10.810 8.810 ;
        RECT -12.880 8.730 -12.670 8.760 ;
        RECT -12.880 8.140 -12.660 8.730 ;
        RECT -12.140 8.170 -11.940 8.740 ;
        RECT -11.130 8.450 -10.810 8.490 ;
        RECT -11.140 8.410 -10.810 8.450 ;
        RECT -11.390 8.240 -10.810 8.410 ;
        RECT -11.130 8.230 -10.810 8.240 ;
        RECT -12.880 7.110 -12.660 7.700 ;
        RECT -12.880 7.080 -12.670 7.110 ;
        RECT -12.140 7.100 -11.940 7.670 ;
        RECT -10.000 7.660 -9.830 8.170 ;
        RECT -5.980 7.690 -5.810 8.200 ;
        RECT -11.130 7.600 -10.810 7.610 ;
        RECT -11.390 7.430 -10.810 7.600 ;
        RECT -11.140 7.390 -10.810 7.430 ;
        RECT -11.130 7.350 -10.810 7.390 ;
        RECT -12.870 6.730 -12.670 7.080 ;
        RECT -11.130 7.030 -10.810 7.060 ;
        RECT -11.140 6.980 -10.810 7.030 ;
        RECT -11.390 6.810 -10.810 6.980 ;
        RECT -11.130 6.800 -10.810 6.810 ;
        RECT -12.500 6.330 -12.060 6.500 ;
        RECT -12.870 5.750 -12.670 6.100 ;
        RECT -11.130 6.020 -10.810 6.030 ;
        RECT -11.390 5.850 -10.810 6.020 ;
        RECT -11.140 5.800 -10.810 5.850 ;
        RECT -10.010 5.800 -9.840 6.990 ;
        RECT -8.200 6.120 -7.650 6.550 ;
        RECT -11.130 5.770 -10.810 5.800 ;
        RECT -12.880 5.720 -12.670 5.750 ;
        RECT -5.990 5.740 -5.820 6.930 ;
        RECT -4.170 6.190 -3.620 6.620 ;
        RECT -12.880 5.130 -12.660 5.720 ;
        RECT -12.140 5.160 -11.940 5.730 ;
        RECT -11.130 5.440 -10.810 5.480 ;
        RECT -11.140 5.400 -10.810 5.440 ;
        RECT -11.390 5.230 -10.810 5.400 ;
        RECT -11.130 5.220 -10.810 5.230 ;
        RECT 0.240 5.100 0.560 5.130 ;
        RECT 0.240 4.930 2.030 5.100 ;
        RECT 0.240 4.910 0.570 4.930 ;
        RECT 0.240 4.870 0.560 4.910 ;
        RECT 1.860 4.700 2.030 4.930 ;
        RECT -12.880 4.110 -12.660 4.700 ;
        RECT -12.880 4.080 -12.670 4.110 ;
        RECT -12.140 4.100 -11.940 4.670 ;
        RECT -11.130 4.600 -10.810 4.610 ;
        RECT -11.390 4.430 -10.810 4.600 ;
        RECT 0.710 4.450 1.050 4.700 ;
        RECT 1.220 4.530 1.550 4.700 ;
        RECT 1.770 4.530 2.110 4.700 ;
        RECT -11.140 4.390 -10.810 4.430 ;
        RECT -11.130 4.350 -10.810 4.390 ;
        RECT 0.390 4.190 1.050 4.450 ;
        RECT 1.300 4.360 1.470 4.530 ;
        RECT 1.860 4.360 2.030 4.530 ;
        RECT 1.220 4.190 1.550 4.360 ;
        RECT 1.770 4.190 2.110 4.360 ;
        RECT -12.870 3.730 -12.670 4.080 ;
        RECT -11.130 4.030 -10.810 4.060 ;
        RECT -11.140 3.980 -10.810 4.030 ;
        RECT -11.390 3.810 -10.810 3.980 ;
        RECT -11.130 3.800 -10.810 3.810 ;
        RECT 1.300 3.960 1.550 4.190 ;
        RECT 2.430 4.110 2.940 4.780 ;
        RECT 1.300 3.790 1.970 3.960 ;
        RECT 1.300 3.560 1.550 3.790 ;
        RECT 0.390 3.300 1.050 3.560 ;
        RECT 1.220 3.390 1.550 3.560 ;
        RECT 1.770 3.390 2.110 3.560 ;
        RECT 0.710 3.050 1.050 3.300 ;
        RECT 1.300 3.220 1.470 3.390 ;
        RECT 1.860 3.220 2.030 3.390 ;
        RECT 1.220 3.050 1.550 3.220 ;
        RECT 1.770 3.050 2.110 3.220 ;
        RECT 0.240 2.840 0.560 2.880 ;
        RECT 0.240 2.820 0.570 2.840 ;
        RECT 1.860 2.820 2.030 3.050 ;
        RECT 2.430 2.970 2.940 3.640 ;
        RECT 0.240 2.650 2.030 2.820 ;
        RECT 0.240 2.620 0.560 2.650 ;
        RECT 0.240 2.330 0.560 2.360 ;
        RECT 0.240 2.160 2.030 2.330 ;
        RECT 0.240 2.140 0.570 2.160 ;
        RECT 0.240 2.100 0.560 2.140 ;
        RECT 1.860 1.930 2.030 2.160 ;
        RECT 0.710 1.680 1.050 1.930 ;
        RECT 1.220 1.760 1.550 1.930 ;
        RECT 1.770 1.760 2.110 1.930 ;
        RECT 0.390 1.420 1.050 1.680 ;
        RECT 1.300 1.590 1.470 1.760 ;
        RECT 1.860 1.590 2.030 1.760 ;
        RECT 1.220 1.420 1.550 1.590 ;
        RECT 1.770 1.420 2.110 1.590 ;
        RECT 1.300 1.190 1.550 1.420 ;
        RECT 2.430 1.340 2.940 2.010 ;
        RECT 1.300 1.020 1.970 1.190 ;
        RECT 1.300 0.790 1.550 1.020 ;
        RECT -11.200 0.690 -10.880 0.730 ;
        RECT -11.200 0.500 -10.870 0.690 ;
        RECT 0.390 0.530 1.050 0.790 ;
        RECT 1.220 0.620 1.550 0.790 ;
        RECT 1.770 0.620 2.110 0.790 ;
        RECT -11.200 0.470 -10.880 0.500 ;
        RECT -11.150 -0.120 -10.970 0.470 ;
        RECT 0.710 0.280 1.050 0.530 ;
        RECT 1.300 0.450 1.470 0.620 ;
        RECT 1.860 0.450 2.030 0.620 ;
        RECT 1.220 0.280 1.550 0.450 ;
        RECT 1.770 0.280 2.110 0.450 ;
        RECT 0.240 0.070 0.560 0.110 ;
        RECT 0.240 0.050 0.570 0.070 ;
        RECT 1.860 0.050 2.030 0.280 ;
        RECT 2.430 0.200 2.940 0.870 ;
        RECT 0.240 -0.120 2.030 0.050 ;
        RECT -11.150 -0.160 -10.830 -0.120 ;
        RECT 0.240 -0.150 0.560 -0.120 ;
        RECT -11.150 -0.350 -10.820 -0.160 ;
        RECT -11.150 -0.380 -10.830 -0.350 ;
      LAYER mcon ;
        RECT -11.040 8.820 -10.870 8.990 ;
        RECT -12.850 8.560 -12.680 8.730 ;
        RECT -12.120 8.530 -11.950 8.700 ;
        RECT -11.040 8.270 -10.870 8.440 ;
        RECT -10.000 8.000 -9.830 8.170 ;
        RECT -12.850 7.110 -12.680 7.280 ;
        RECT -5.980 8.030 -5.810 8.200 ;
        RECT -11.040 7.400 -10.870 7.570 ;
        RECT -12.120 7.140 -11.950 7.310 ;
        RECT -11.040 6.850 -10.870 7.020 ;
        RECT -10.010 6.820 -9.840 6.990 ;
        RECT -10.010 6.480 -9.840 6.650 ;
        RECT -5.990 6.760 -5.820 6.930 ;
        RECT -10.010 6.140 -9.840 6.310 ;
        RECT -11.040 5.810 -10.870 5.980 ;
        RECT -7.920 6.200 -7.650 6.470 ;
        RECT -5.990 6.420 -5.820 6.590 ;
        RECT -5.990 6.080 -5.820 6.250 ;
        RECT -3.890 6.270 -3.620 6.540 ;
        RECT -12.850 5.550 -12.680 5.720 ;
        RECT -12.120 5.520 -11.950 5.690 ;
        RECT -11.040 5.260 -10.870 5.430 ;
        RECT 0.300 4.920 0.470 5.090 ;
        RECT -12.850 4.110 -12.680 4.280 ;
        RECT -11.040 4.400 -10.870 4.570 ;
        RECT -12.120 4.140 -11.950 4.310 ;
        RECT 0.450 4.240 0.620 4.410 ;
        RECT 2.600 4.360 2.770 4.530 ;
        RECT -11.040 3.850 -10.870 4.020 ;
        RECT 1.340 3.790 1.510 3.960 ;
        RECT 0.450 3.340 0.620 3.510 ;
        RECT 2.600 3.220 2.770 3.390 ;
        RECT 0.300 2.660 0.470 2.830 ;
        RECT 0.300 2.150 0.470 2.320 ;
        RECT 0.450 1.470 0.620 1.640 ;
        RECT 2.600 1.590 2.770 1.760 ;
        RECT 1.340 1.020 1.510 1.190 ;
        RECT -11.140 0.510 -10.970 0.680 ;
        RECT 0.450 0.570 0.620 0.740 ;
        RECT 2.600 0.450 2.770 0.620 ;
        RECT 0.300 -0.110 0.470 0.060 ;
        RECT -11.090 -0.340 -10.920 -0.170 ;
      LAYER met1 ;
        RECT -12.910 8.790 -12.750 9.440 ;
        RECT -12.910 8.240 -12.640 8.790 ;
        RECT -12.920 8.190 -12.640 8.240 ;
        RECT -12.500 8.450 -12.310 9.440 ;
        RECT -12.100 8.760 -11.940 9.440 ;
        RECT -12.140 8.740 -11.940 8.760 ;
        RECT -11.120 8.750 -10.800 9.070 ;
        RECT -12.150 8.500 -11.920 8.740 ;
        RECT -12.500 8.330 -12.330 8.450 ;
        RECT -12.920 8.100 -12.750 8.190 ;
        RECT -12.910 7.740 -12.750 8.100 ;
        RECT -12.920 7.650 -12.750 7.740 ;
        RECT -12.920 7.600 -12.640 7.650 ;
        RECT -12.910 7.050 -12.640 7.600 ;
        RECT -12.500 7.510 -12.340 8.330 ;
        RECT -12.140 8.280 -11.940 8.500 ;
        RECT -12.100 7.560 -11.940 8.280 ;
        RECT -11.120 8.200 -10.800 8.520 ;
        RECT -12.500 7.390 -12.330 7.510 ;
        RECT -12.910 5.780 -12.750 7.050 ;
        RECT -12.500 6.530 -12.310 7.390 ;
        RECT -12.140 7.340 -11.940 7.560 ;
        RECT -12.150 7.100 -11.920 7.340 ;
        RECT -11.120 7.320 -10.800 7.640 ;
        RECT -12.140 7.080 -11.940 7.100 ;
        RECT -12.530 6.300 -12.290 6.530 ;
        RECT -12.910 5.230 -12.640 5.780 ;
        RECT -12.920 5.180 -12.640 5.230 ;
        RECT -12.500 5.440 -12.310 6.300 ;
        RECT -12.100 5.750 -11.940 7.080 ;
        RECT -11.120 6.770 -10.800 7.090 ;
        RECT -12.140 5.730 -11.940 5.750 ;
        RECT -11.120 5.740 -10.800 6.060 ;
        RECT -12.150 5.490 -11.920 5.730 ;
        RECT -10.040 5.620 -9.790 9.440 ;
        RECT -7.980 7.520 -7.600 9.440 ;
        RECT -7.980 5.660 -7.590 7.520 ;
        RECT -10.040 5.550 -9.650 5.620 ;
        RECT -12.500 5.320 -12.330 5.440 ;
        RECT -12.920 5.090 -12.750 5.180 ;
        RECT -12.910 4.740 -12.750 5.090 ;
        RECT -12.920 4.650 -12.750 4.740 ;
        RECT -12.920 4.600 -12.640 4.650 ;
        RECT -12.910 4.050 -12.640 4.600 ;
        RECT -12.500 4.510 -12.340 5.320 ;
        RECT -12.140 5.270 -11.940 5.490 ;
        RECT -12.100 4.560 -11.940 5.270 ;
        RECT -11.120 5.190 -10.800 5.510 ;
        RECT -10.040 5.000 -9.790 5.550 ;
        RECT -7.980 5.360 -7.600 5.660 ;
        RECT -7.980 5.040 -7.560 5.360 ;
        RECT -10.060 4.970 -9.780 5.000 ;
        RECT -10.070 4.690 -9.770 4.970 ;
        RECT -10.060 4.670 -9.780 4.690 ;
        RECT -12.500 4.390 -12.330 4.510 ;
        RECT -12.910 3.400 -12.750 4.050 ;
        RECT -12.500 3.400 -12.310 4.390 ;
        RECT -12.140 4.340 -11.940 4.560 ;
        RECT -12.150 4.100 -11.920 4.340 ;
        RECT -11.120 4.320 -10.800 4.640 ;
        RECT -12.140 4.080 -11.940 4.100 ;
        RECT -12.100 3.400 -11.940 4.080 ;
        RECT -10.040 3.390 -9.790 4.670 ;
        RECT -7.980 4.310 -7.600 5.040 ;
        RECT -6.030 4.970 -5.760 9.440 ;
        RECT -6.050 4.660 -5.740 4.970 ;
        RECT -7.980 3.990 -7.580 4.310 ;
        RECT -7.980 3.390 -7.600 3.990 ;
        RECT -6.030 3.390 -5.760 4.660 ;
        RECT -3.950 3.390 -3.550 9.440 ;
        RECT 0.230 4.840 0.550 5.160 ;
        RECT 0.380 4.160 0.700 4.480 ;
        RECT 0.380 3.270 0.700 3.590 ;
        RECT 0.230 2.590 0.550 2.910 ;
        RECT -7.840 2.110 -7.580 2.430 ;
        RECT -7.840 1.250 -7.680 2.110 ;
        RECT 0.230 2.070 0.550 2.390 ;
        RECT 0.380 1.390 0.700 1.710 ;
        RECT -8.000 0.930 -7.680 1.250 ;
        RECT -11.210 0.440 -10.890 0.760 ;
        RECT 0.380 0.500 0.700 0.820 ;
        RECT -11.160 -0.410 -10.840 -0.090 ;
        RECT 0.230 -0.180 0.550 0.140 ;
        RECT -5.320 -0.430 -4.940 -0.330 ;
      LAYER via ;
        RECT -11.090 8.780 -10.830 9.040 ;
        RECT -11.090 8.230 -10.830 8.490 ;
        RECT -11.090 7.350 -10.830 7.610 ;
        RECT -11.090 6.800 -10.830 7.060 ;
        RECT -11.090 5.770 -10.830 6.030 ;
        RECT -11.090 5.220 -10.830 5.480 ;
        RECT -7.820 5.070 -7.560 5.330 ;
        RECT -10.050 4.700 -9.790 4.960 ;
        RECT -11.090 4.350 -10.830 4.610 ;
        RECT -6.030 4.680 -5.760 4.940 ;
        RECT -7.840 4.020 -7.580 4.280 ;
        RECT 0.260 4.870 0.520 5.130 ;
        RECT 0.410 4.190 0.670 4.450 ;
        RECT 0.410 3.300 0.670 3.560 ;
        RECT 0.260 2.620 0.520 2.880 ;
        RECT -7.840 2.140 -7.580 2.400 ;
        RECT 0.260 2.100 0.520 2.360 ;
        RECT 0.410 1.420 0.670 1.680 ;
        RECT -8.000 0.960 -7.740 1.220 ;
        RECT -11.180 0.470 -10.920 0.730 ;
        RECT 0.410 0.530 0.670 0.790 ;
        RECT -11.130 -0.380 -10.870 -0.120 ;
        RECT 0.260 -0.150 0.520 0.110 ;
      LAYER met2 ;
        RECT -11.110 8.940 -10.800 9.080 ;
        RECT -13.270 8.760 -10.700 8.940 ;
        RECT -11.110 8.750 -10.800 8.760 ;
        RECT -11.110 8.510 -10.800 8.530 ;
        RECT -13.270 8.330 -3.190 8.510 ;
        RECT -11.110 8.200 -10.800 8.330 ;
        RECT -3.340 8.320 -3.190 8.330 ;
        RECT -11.110 7.510 -10.800 7.640 ;
        RECT -3.310 7.510 -3.170 7.530 ;
        RECT -13.280 7.330 -3.170 7.510 ;
        RECT -11.110 7.310 -10.800 7.330 ;
        RECT -11.110 7.080 -10.800 7.090 ;
        RECT -13.270 7.040 -10.800 7.080 ;
        RECT -13.270 6.900 -10.710 7.040 ;
        RECT -11.110 6.760 -10.800 6.900 ;
        RECT -11.110 5.930 -10.800 6.070 ;
        RECT -13.280 5.920 -10.800 5.930 ;
        RECT -13.280 5.750 -10.680 5.920 ;
        RECT -11.110 5.740 -10.800 5.750 ;
  END
END sky130_hilas_WTA4Stage01

MACRO sky130_hilas_Trans4small
  CLASS BLOCK ;
  FOREIGN sky130_hilas_Trans4small ;
  ORIGIN -1.910 1.500 ;
  SIZE 2.800 BY 5.880 ;
  PIN NFET_SOURCE1
    USE ANALOG ;
    ANTENNADIFFAREA 0.108500 ;
    PORT
      LAYER met2 ;
        RECT 2.510 4.150 2.820 4.240 ;
        RECT 1.910 3.980 2.820 4.150 ;
        RECT 2.510 3.910 2.820 3.980 ;
    END
  END NFET_SOURCE1
  PIN NFET_GATE1
    USE ANALOG ;
    ANTENNAGATEAREA 0.094500 ;
    PORT
      LAYER met2 ;
        RECT 2.040 3.740 2.360 3.820 ;
        RECT 1.910 3.570 2.360 3.740 ;
        RECT 2.040 3.500 2.360 3.570 ;
    END
  END NFET_GATE1
  PIN NFET_SOURCE2
    USE ANALOG ;
    ANTENNADIFFAREA 0.108500 ;
    PORT
      LAYER met2 ;
        RECT 2.510 3.230 2.820 3.320 ;
        RECT 1.910 3.060 2.820 3.230 ;
        RECT 2.510 2.990 2.820 3.060 ;
    END
  END NFET_SOURCE2
  PIN NFET_GATE2
    USE ANALOG ;
    ANTENNAGATEAREA 0.094500 ;
    PORT
      LAYER met2 ;
        RECT 2.040 2.820 2.360 2.900 ;
        RECT 1.910 2.650 2.360 2.820 ;
        RECT 2.040 2.580 2.360 2.650 ;
    END
  END NFET_GATE2
  PIN NFET_SOURCE3
    USE ANALOG ;
    ANTENNADIFFAREA 0.108500 ;
    PORT
      LAYER met2 ;
        RECT 2.510 2.310 2.820 2.400 ;
        RECT 1.910 2.140 2.820 2.310 ;
        RECT 2.510 2.070 2.820 2.140 ;
    END
  END NFET_SOURCE3
  PIN NFET_GATE3
    USE ANALOG ;
    ANTENNAGATEAREA 0.094500 ;
    PORT
      LAYER met2 ;
        RECT 2.040 1.900 2.360 1.980 ;
        RECT 1.910 1.730 2.360 1.900 ;
        RECT 2.040 1.660 2.360 1.730 ;
    END
  END NFET_GATE3
  PIN PFET_SOURCE1
    USE ANALOG ;
    ANTENNADIFFAREA 0.109200 ;
    PORT
      LAYER met2 ;
        RECT 2.320 1.310 2.630 1.420 ;
        RECT 1.910 1.120 2.630 1.310 ;
        RECT 2.320 1.090 2.630 1.120 ;
    END
  END PFET_SOURCE1
  PIN PFET_GATE1
    USE ANALOG ;
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER met2 ;
        RECT 2.320 0.890 2.640 0.950 ;
        RECT 1.910 0.700 2.640 0.890 ;
        RECT 2.320 0.630 2.640 0.700 ;
    END
  END PFET_GATE1
  PIN PFET_SOURCE2
    USE ANALOG ;
    ANTENNADIFFAREA 0.109200 ;
    PORT
      LAYER met2 ;
        RECT 2.320 0.350 2.630 0.460 ;
        RECT 1.910 0.160 2.630 0.350 ;
        RECT 2.320 0.130 2.630 0.160 ;
    END
  END PFET_SOURCE2
  PIN PFET_GATE2
    USE ANALOG ;
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER met2 ;
        RECT 2.320 -0.070 2.640 -0.010 ;
        RECT 1.910 -0.260 2.640 -0.070 ;
        RECT 2.320 -0.330 2.640 -0.260 ;
    END
  END PFET_GATE2
  PIN PFET_SOURCE3
    USE ANALOG ;
    ANTENNADIFFAREA 0.109200 ;
    PORT
      LAYER met2 ;
        RECT 2.320 -0.610 2.630 -0.500 ;
        RECT 1.910 -0.800 2.630 -0.610 ;
        RECT 2.320 -0.830 2.630 -0.800 ;
    END
  END PFET_SOURCE3
  PIN PFET_GATE3
    USE ANALOG ;
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER met2 ;
        RECT 2.320 -1.030 2.640 -0.970 ;
        RECT 1.910 -1.220 2.640 -1.030 ;
        RECT 2.320 -1.290 2.640 -1.220 ;
    END
  END PFET_GATE3
  PIN WELL
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 1.980 -1.500 4.550 1.590 ;
      LAYER met1 ;
        RECT 4.090 -1.100 4.310 4.380 ;
        RECT 4.030 -1.330 4.320 -1.100 ;
        RECT 4.090 -1.500 4.310 -1.330 ;
    END
  END WELL
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 4.490 3.750 4.710 4.380 ;
        RECT 4.480 3.460 4.710 3.750 ;
        RECT 4.490 -1.500 4.710 3.460 ;
    END
  END VGND
  PIN PFET_DRAIN3
    USE ANALOG ;
    ANTENNADIFFAREA 0.105300 ;
    PORT
      LAYER met2 ;
        RECT 3.620 -0.670 3.930 -0.600 ;
        RECT 3.620 -0.870 4.710 -0.670 ;
        RECT 3.620 -0.930 3.930 -0.870 ;
    END
  END PFET_DRAIN3
  PIN PFET_DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.105300 ;
    PORT
      LAYER met2 ;
        RECT 3.620 0.290 3.930 0.360 ;
        RECT 3.620 0.090 4.710 0.290 ;
        RECT 3.620 0.030 3.930 0.090 ;
    END
  END PFET_DRAIN2
  PIN PFET_DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.105300 ;
    PORT
      LAYER met2 ;
        RECT 3.620 1.250 3.930 1.320 ;
        RECT 3.620 1.050 4.710 1.250 ;
        RECT 3.620 0.990 3.930 1.050 ;
    END
  END PFET_DRAIN1
  PIN NFET_DRAIN3
    USE ANALOG ;
    ANTENNADIFFAREA 0.108500 ;
    PORT
      LAYER met2 ;
        RECT 3.600 2.320 3.910 2.410 ;
        RECT 3.600 2.150 4.710 2.320 ;
        RECT 3.600 2.080 3.910 2.150 ;
    END
  END NFET_DRAIN3
  PIN NFET_DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.108500 ;
    PORT
      LAYER met2 ;
        RECT 3.600 3.240 3.910 3.330 ;
        RECT 3.600 3.070 4.710 3.240 ;
        RECT 3.600 3.000 3.910 3.070 ;
    END
  END NFET_DRAIN2
  PIN NFET_DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.108500 ;
    PORT
      LAYER met2 ;
        RECT 3.600 4.160 3.910 4.250 ;
        RECT 3.600 3.990 4.710 4.160 ;
        RECT 3.600 3.920 3.910 3.990 ;
    END
  END NFET_DRAIN1
  OBS
      LAYER li1 ;
        RECT 2.830 4.200 3.030 4.240 ;
        RECT 2.520 3.940 3.030 4.200 ;
        RECT 2.830 3.910 3.030 3.940 ;
        RECT 3.420 4.210 3.620 4.240 ;
        RECT 3.420 4.170 3.930 4.210 ;
        RECT 3.420 3.980 3.940 4.170 ;
        RECT 3.420 3.950 3.930 3.980 ;
        RECT 3.420 3.910 3.620 3.950 ;
        RECT 4.110 3.760 4.280 3.810 ;
        RECT 2.080 3.740 2.510 3.760 ;
        RECT 2.080 3.570 2.530 3.740 ;
        RECT 4.100 3.730 4.280 3.760 ;
        RECT 4.100 3.720 4.530 3.730 ;
        RECT 2.080 3.550 2.510 3.570 ;
        RECT 4.100 3.490 4.690 3.720 ;
        RECT 4.100 3.480 4.530 3.490 ;
        RECT 4.100 3.420 4.270 3.480 ;
        RECT 2.830 3.280 3.030 3.320 ;
        RECT 2.520 3.020 3.030 3.280 ;
        RECT 2.830 2.990 3.030 3.020 ;
        RECT 3.420 3.290 3.620 3.320 ;
        RECT 3.420 3.250 3.930 3.290 ;
        RECT 3.420 3.060 3.940 3.250 ;
        RECT 3.420 3.030 3.930 3.060 ;
        RECT 3.420 2.990 3.620 3.030 ;
        RECT 2.080 2.820 2.510 2.840 ;
        RECT 2.080 2.650 2.530 2.820 ;
        RECT 2.080 2.630 2.510 2.650 ;
        RECT 2.830 2.360 3.030 2.400 ;
        RECT 2.520 2.100 3.030 2.360 ;
        RECT 2.830 2.070 3.030 2.100 ;
        RECT 3.420 2.370 3.620 2.400 ;
        RECT 3.420 2.330 3.930 2.370 ;
        RECT 3.420 2.140 3.940 2.330 ;
        RECT 3.420 2.110 3.930 2.140 ;
        RECT 3.420 2.070 3.620 2.110 ;
        RECT 2.080 1.900 2.510 1.920 ;
        RECT 2.080 1.730 2.530 1.900 ;
        RECT 2.080 1.710 2.510 1.730 ;
        RECT 2.330 1.340 2.650 1.380 ;
        RECT 2.330 1.320 2.660 1.340 ;
        RECT 2.330 1.120 2.950 1.320 ;
        RECT 2.780 0.990 2.950 1.120 ;
        RECT 3.460 1.280 3.630 1.320 ;
        RECT 3.460 1.240 3.950 1.280 ;
        RECT 3.460 1.050 3.960 1.240 ;
        RECT 3.460 1.020 3.950 1.050 ;
        RECT 3.460 0.990 3.630 1.020 ;
        RECT 2.170 0.880 2.600 0.900 ;
        RECT 2.150 0.710 2.600 0.880 ;
        RECT 2.170 0.690 2.600 0.710 ;
        RECT 2.330 0.380 2.650 0.420 ;
        RECT 2.330 0.360 2.660 0.380 ;
        RECT 2.330 0.160 2.950 0.360 ;
        RECT 2.780 0.030 2.950 0.160 ;
        RECT 3.460 0.320 3.630 0.360 ;
        RECT 3.460 0.280 3.950 0.320 ;
        RECT 3.460 0.090 3.960 0.280 ;
        RECT 3.460 0.060 3.950 0.090 ;
        RECT 3.460 0.030 3.630 0.060 ;
        RECT 2.170 -0.080 2.600 -0.060 ;
        RECT 2.150 -0.250 2.600 -0.080 ;
        RECT 2.170 -0.270 2.600 -0.250 ;
        RECT 2.330 -0.580 2.650 -0.540 ;
        RECT 2.330 -0.600 2.660 -0.580 ;
        RECT 2.330 -0.800 2.950 -0.600 ;
        RECT 2.780 -0.930 2.950 -0.800 ;
        RECT 3.460 -0.640 3.630 -0.600 ;
        RECT 3.460 -0.680 3.950 -0.640 ;
        RECT 3.460 -0.870 3.960 -0.680 ;
        RECT 3.460 -0.900 3.950 -0.870 ;
        RECT 3.460 -0.930 3.630 -0.900 ;
        RECT 2.170 -1.040 2.600 -1.020 ;
        RECT 2.150 -1.210 2.600 -1.040 ;
        RECT 2.170 -1.230 2.600 -1.210 ;
        RECT 3.960 -1.270 4.380 -1.100 ;
        RECT 4.060 -1.310 4.290 -1.270 ;
      LAYER mcon ;
        RECT 2.580 3.980 2.750 4.150 ;
        RECT 3.670 3.990 3.840 4.160 ;
        RECT 2.360 3.570 2.530 3.740 ;
        RECT 4.510 3.520 4.680 3.690 ;
        RECT 2.580 3.060 2.750 3.230 ;
        RECT 3.670 3.070 3.840 3.240 ;
        RECT 2.360 2.650 2.530 2.820 ;
        RECT 2.580 2.140 2.750 2.310 ;
        RECT 3.670 2.150 3.840 2.320 ;
        RECT 2.360 1.730 2.530 1.900 ;
        RECT 2.390 1.160 2.560 1.330 ;
        RECT 3.690 1.060 3.860 1.230 ;
        RECT 2.390 0.200 2.560 0.370 ;
        RECT 3.690 0.100 3.860 0.270 ;
        RECT 2.390 -0.760 2.560 -0.590 ;
        RECT 3.690 -0.860 3.860 -0.690 ;
        RECT 4.090 -1.300 4.260 -1.130 ;
      LAYER met1 ;
        RECT 2.510 3.910 2.830 4.230 ;
        RECT 3.600 3.920 3.920 4.240 ;
        RECT 2.040 3.770 2.360 3.820 ;
        RECT 2.040 3.540 2.590 3.770 ;
        RECT 2.040 3.500 2.360 3.540 ;
        RECT 2.510 2.990 2.830 3.310 ;
        RECT 3.600 3.000 3.920 3.320 ;
        RECT 2.040 2.850 2.360 2.900 ;
        RECT 2.040 2.620 2.590 2.850 ;
        RECT 2.040 2.580 2.360 2.620 ;
        RECT 2.510 2.070 2.830 2.390 ;
        RECT 3.600 2.080 3.920 2.400 ;
        RECT 2.040 1.930 2.360 1.980 ;
        RECT 2.040 1.700 2.590 1.930 ;
        RECT 2.040 1.660 2.360 1.700 ;
        RECT 2.320 1.090 2.640 1.410 ;
        RECT 3.620 0.990 3.940 1.310 ;
        RECT 2.320 0.910 2.640 0.950 ;
        RECT 2.090 0.680 2.640 0.910 ;
        RECT 2.320 0.630 2.640 0.680 ;
        RECT 2.320 0.130 2.640 0.450 ;
        RECT 3.620 0.030 3.940 0.350 ;
        RECT 2.320 -0.050 2.640 -0.010 ;
        RECT 2.090 -0.280 2.640 -0.050 ;
        RECT 2.320 -0.330 2.640 -0.280 ;
        RECT 2.320 -0.830 2.640 -0.510 ;
        RECT 3.620 -0.930 3.940 -0.610 ;
        RECT 2.320 -1.010 2.640 -0.970 ;
        RECT 2.090 -1.240 2.640 -1.010 ;
        RECT 2.320 -1.290 2.640 -1.240 ;
      LAYER via ;
        RECT 2.540 3.940 2.800 4.200 ;
        RECT 3.630 3.950 3.890 4.210 ;
        RECT 2.070 3.530 2.330 3.790 ;
        RECT 2.540 3.020 2.800 3.280 ;
        RECT 3.630 3.030 3.890 3.290 ;
        RECT 2.070 2.610 2.330 2.870 ;
        RECT 2.540 2.100 2.800 2.360 ;
        RECT 3.630 2.110 3.890 2.370 ;
        RECT 2.070 1.690 2.330 1.950 ;
        RECT 2.350 1.120 2.610 1.380 ;
        RECT 3.650 1.020 3.910 1.280 ;
        RECT 2.350 0.660 2.610 0.920 ;
        RECT 2.350 0.160 2.610 0.420 ;
        RECT 3.650 0.060 3.910 0.320 ;
        RECT 2.350 -0.300 2.610 -0.040 ;
        RECT 2.350 -0.800 2.610 -0.540 ;
        RECT 3.650 -0.900 3.910 -0.640 ;
        RECT 2.350 -1.260 2.610 -1.000 ;
  END
END sky130_hilas_Trans4small

MACRO sky130_hilas_FGBiasWeakGate2x1cell
  CLASS CORE ;
  FOREIGN sky130_hilas_FGBiasWeakGate2x1cell ;
  ORIGIN -0.010 0.000 ;
  SIZE 11.530 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.105400 ;
    PORT
      LAYER met2 ;
        RECT 9.060 5.550 9.370 5.560 ;
        RECT 0.010 5.370 11.540 5.550 ;
        RECT 9.060 5.230 9.370 5.370 ;
    END
  END DRAIN1
  PIN VIN11
    PORT
      LAYER met2 ;
        RECT 1.950 4.960 2.260 5.010 ;
        RECT 1.800 4.950 2.260 4.960 ;
        RECT 0.010 4.770 2.260 4.950 ;
        RECT 1.950 4.680 2.260 4.770 ;
    END
  END VIN11
  PIN ROW1
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 9.210 4.530 9.520 4.600 ;
        RECT 9.210 4.520 11.540 4.530 ;
        RECT 0.010 4.310 11.540 4.520 ;
        RECT 0.010 4.300 10.230 4.310 ;
        RECT 9.210 4.270 9.520 4.300 ;
    END
  END ROW1
  PIN ROW2
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 9.210 1.770 9.520 1.840 ;
        RECT 0.010 1.560 11.540 1.770 ;
        RECT 0.010 1.550 10.230 1.560 ;
        RECT 9.210 1.510 9.520 1.550 ;
    END
  END ROW2
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 8.230 0.010 11.540 6.040 ;
      LAYER met1 ;
        RECT 11.020 5.400 11.300 6.050 ;
        RECT 10.910 4.800 11.300 5.400 ;
        RECT 11.020 1.250 11.300 4.800 ;
        RECT 10.910 0.650 11.300 1.250 ;
        RECT 11.020 0.000 11.300 0.650 ;
    END
  END VINJ
  PIN COLSEL1
    USE ANALOG ;
    ANTENNAGATEAREA 0.310000 ;
    PORT
      LAYER met1 ;
        RECT 10.580 4.590 10.770 6.050 ;
        RECT 10.580 4.560 10.800 4.590 ;
        RECT 10.560 4.290 10.810 4.560 ;
        RECT 10.570 4.280 10.810 4.290 ;
        RECT 10.570 4.040 10.800 4.280 ;
        RECT 10.610 2.010 10.770 4.040 ;
        RECT 10.570 1.770 10.800 2.010 ;
        RECT 10.570 1.760 10.810 1.770 ;
        RECT 10.560 1.490 10.810 1.760 ;
        RECT 10.580 1.460 10.800 1.490 ;
        RECT 10.580 0.000 10.770 1.460 ;
    END
  END COLSEL1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2.840 5.080 3.070 6.050 ;
        RECT 2.840 4.830 3.080 5.080 ;
        RECT 2.840 0.000 3.070 4.830 ;
    END
  END VGND
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT 3.780 3.660 6.500 5.310 ;
        RECT 3.780 3.620 6.490 3.660 ;
        RECT 3.780 2.290 6.490 2.330 ;
        RECT 3.780 0.640 6.500 2.290 ;
      LAYER met1 ;
        RECT 4.060 4.840 4.290 6.050 ;
        RECT 4.060 4.050 4.320 4.840 ;
        RECT 4.060 1.900 4.290 4.050 ;
        RECT 4.060 1.110 4.320 1.900 ;
        RECT 4.060 0.000 4.290 1.110 ;
    END
  END GATE1
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 2.516100 ;
    PORT
      LAYER nwell ;
        RECT 0.020 5.300 1.750 6.050 ;
        RECT 0.020 1.730 1.760 5.300 ;
        RECT 0.020 0.010 1.750 1.730 ;
      LAYER met1 ;
        RECT 0.360 0.010 0.780 6.050 ;
    END
  END VTUN
  PIN DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.105400 ;
    PORT
      LAYER met2 ;
        RECT 9.060 0.680 9.370 0.820 ;
        RECT 9.060 0.670 11.540 0.680 ;
        RECT 0.010 0.520 11.540 0.670 ;
        RECT 9.060 0.500 11.540 0.520 ;
        RECT 9.060 0.490 9.370 0.500 ;
    END
  END DRAIN2
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.920 1.240 2.230 1.320 ;
        RECT 0.010 1.030 2.230 1.240 ;
        RECT 1.920 0.990 2.230 1.030 ;
    END
  END VIN12
  PIN COMMONSOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 1.030400 ;
    PORT
      LAYER met2 ;
        RECT 0.010 3.330 10.470 3.550 ;
        RECT 10.150 3.190 10.470 3.330 ;
        RECT 10.190 2.850 10.450 3.190 ;
        RECT 10.150 2.590 10.470 2.850 ;
    END
  END COMMONSOURCE
  OBS
      LAYER li1 ;
        RECT 1.880 5.040 6.940 5.870 ;
        RECT 9.130 5.470 9.660 5.640 ;
        RECT 10.940 5.370 11.140 5.720 ;
        RECT 10.940 5.340 11.150 5.370 ;
        RECT 1.950 4.960 2.430 5.040 ;
        RECT 1.960 4.710 2.430 4.960 ;
        RECT 7.260 4.890 7.610 5.060 ;
        RECT 8.630 4.890 8.960 5.060 ;
        RECT 0.450 3.910 1.000 4.340 ;
        RECT 4.080 4.100 4.310 4.790 ;
        RECT 9.380 4.560 9.550 5.080 ;
        RECT 9.220 4.300 9.550 4.560 ;
        RECT 7.260 4.100 7.610 4.270 ;
        RECT 8.630 4.100 8.960 4.270 ;
        RECT 3.050 3.080 3.240 3.480 ;
        RECT 7.270 3.310 7.610 3.480 ;
        RECT 8.630 3.310 8.960 3.480 ;
        RECT 9.380 3.390 9.550 4.300 ;
        RECT 10.210 3.480 10.380 5.090 ;
        RECT 10.930 4.760 11.150 5.340 ;
        RECT 10.940 4.750 11.150 4.760 ;
        RECT 10.580 4.580 10.770 4.590 ;
        RECT 10.580 4.290 10.780 4.580 ;
        RECT 10.570 3.960 10.810 4.290 ;
        RECT 2.860 3.070 3.240 3.080 ;
        RECT 2.860 2.890 6.600 3.070 ;
        RECT 2.860 2.850 3.240 2.890 ;
        RECT 0.450 2.180 1.000 2.610 ;
        RECT 3.050 2.470 3.240 2.850 ;
        RECT 8.710 2.740 8.880 3.310 ;
        RECT 10.210 3.290 10.390 3.480 ;
        RECT 7.270 2.570 7.610 2.740 ;
        RECT 8.630 2.570 8.960 2.740 ;
        RECT 1.930 1.030 2.270 1.280 ;
        RECT 4.080 1.160 4.310 1.890 ;
        RECT 7.260 1.780 7.610 1.950 ;
        RECT 8.630 1.780 8.960 1.950 ;
        RECT 9.380 1.800 9.550 2.660 ;
        RECT 9.220 1.540 9.550 1.800 ;
        RECT 1.920 0.950 2.270 1.030 ;
        RECT 7.260 0.990 7.610 1.160 ;
        RECT 8.630 0.990 8.960 1.160 ;
        RECT 9.380 0.970 9.550 1.540 ;
        RECT 10.210 2.570 10.390 2.760 ;
        RECT 10.210 0.960 10.380 2.570 ;
        RECT 10.570 1.760 10.810 2.090 ;
        RECT 10.580 1.470 10.780 1.760 ;
        RECT 10.580 1.460 10.770 1.470 ;
        RECT 10.940 1.290 11.150 1.300 ;
        RECT 1.920 0.100 6.970 0.950 ;
        RECT 10.930 0.710 11.150 1.290 ;
        RECT 10.940 0.680 11.150 0.710 ;
        RECT 9.130 0.410 9.660 0.580 ;
        RECT 10.940 0.330 11.140 0.680 ;
      LAYER mcon ;
        RECT 10.950 5.170 11.120 5.340 ;
        RECT 2.020 4.750 2.190 4.920 ;
        RECT 4.110 4.590 4.280 4.760 ;
        RECT 0.450 3.990 0.720 4.260 ;
        RECT 4.110 4.140 4.280 4.310 ;
        RECT 9.280 4.340 9.450 4.510 ;
        RECT 10.590 4.330 10.770 4.520 ;
        RECT 2.870 2.880 3.040 3.050 ;
        RECT 0.450 2.260 0.720 2.530 ;
        RECT 4.110 1.640 4.280 1.810 ;
        RECT 9.280 1.580 9.450 1.750 ;
        RECT 1.990 1.060 2.160 1.230 ;
        RECT 4.110 1.190 4.280 1.360 ;
        RECT 10.590 1.530 10.770 1.720 ;
        RECT 10.950 0.710 11.120 0.880 ;
      LAYER met1 ;
        RECT 9.060 5.230 9.370 5.670 ;
        RECT 1.950 4.680 2.270 5.000 ;
        RECT 9.210 4.270 9.530 4.590 ;
        RECT 10.180 3.480 10.420 3.610 ;
        RECT 10.180 3.160 10.440 3.480 ;
        RECT 10.180 2.560 10.440 2.880 ;
        RECT 10.180 2.440 10.420 2.560 ;
        RECT 9.210 1.510 9.530 1.830 ;
        RECT 1.920 0.990 2.240 1.310 ;
        RECT 9.060 0.380 9.370 0.820 ;
      LAYER via ;
        RECT 9.090 5.260 9.350 5.520 ;
        RECT 1.980 4.710 2.240 4.970 ;
        RECT 9.240 4.300 9.500 4.560 ;
        RECT 10.180 3.190 10.440 3.450 ;
        RECT 10.180 2.590 10.440 2.850 ;
        RECT 9.240 1.540 9.500 1.800 ;
        RECT 1.950 1.020 2.210 1.280 ;
        RECT 9.090 0.530 9.350 0.790 ;
  END
END sky130_hilas_FGBiasWeakGate2x1cell

MACRO sky130_hilas_swc4x2cell
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x2cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.400 BY 9.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 17.090 5.950 17.470 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.090 0.000 17.470 0.150 ;
    END
  END GATE2
  PIN VTUN
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 11.960 0.000 12.360 0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.040 0.000 13.440 0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.040 5.950 13.440 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.960 5.920 12.360 6.050 ;
    END
  END VTUN
  PIN GATE1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 7.930 5.950 8.310 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 7.930 0.000 8.310 0.090 ;
    END
  END GATE1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 22.240 0.010 22.400 0.070 ;
    END
  END VINJ
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 2.160 5.930 2.470 5.950 ;
        RECT 2.840 5.930 5.690 6.010 ;
        RECT 19.730 5.930 22.560 6.010 ;
        RECT 22.930 5.930 23.240 5.950 ;
        RECT 0.000 5.910 10.060 5.930 ;
        RECT 15.340 5.910 25.400 5.930 ;
        RECT 0.000 5.760 25.400 5.910 ;
        RECT 0.000 5.750 2.560 5.760 ;
        RECT 2.160 5.620 2.470 5.750 ;
        RECT 2.840 5.710 3.260 5.760 ;
        RECT 5.250 5.730 19.930 5.760 ;
        RECT 22.240 5.710 22.560 5.760 ;
        RECT 22.840 5.750 25.400 5.760 ;
        RECT 22.930 5.620 23.240 5.750 ;
        RECT 3.070 5.380 3.390 5.460 ;
        RECT 7.000 5.380 7.320 5.390 ;
        RECT 3.070 5.200 7.320 5.380 ;
        RECT 3.070 5.140 3.390 5.200 ;
        RECT 7.000 5.130 7.320 5.200 ;
        RECT 18.080 5.380 18.400 5.390 ;
        RECT 22.010 5.380 22.330 5.460 ;
        RECT 18.080 5.200 22.330 5.380 ;
        RECT 18.080 5.130 18.400 5.200 ;
        RECT 22.010 5.140 22.330 5.200 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.110 8.710 3.350 9.870 ;
        RECT 3.100 8.050 3.370 8.710 ;
        RECT 3.110 6.050 3.350 8.050 ;
        RECT 3.000 6.010 3.350 6.050 ;
        RECT 2.840 5.710 3.350 6.010 ;
        RECT 3.110 5.460 3.350 5.710 ;
        RECT 3.100 5.140 3.360 5.460 ;
        RECT 3.110 3.820 3.350 5.140 ;
      LAYER via ;
        RECT 2.870 5.730 3.130 5.990 ;
        RECT 3.100 5.170 3.360 5.430 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.000 0.000 3.160 0.060 ;
    END
  END VINJ
  PIN GATESELECT1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 3.410 6.000 3.600 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.410 0.010 3.600 0.070 ;
    END
  END GATESELECT1
  PIN GATESELECT2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 21.800 0.010 21.990 0.070 ;
    END
  END GATESELECT2
  PIN COL1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 3.810 6.000 3.970 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.810 0.010 3.970 0.070 ;
    END
  END COL1
  PIN COL2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 21.430 0.010 21.590 0.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.430 6.000 21.590 6.050 ;
    END
  END COL2
  PIN ROW1
    USE ANALOG ;
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 2.160 4.950 2.470 5.070 ;
        RECT 2.640 4.950 2.780 5.130 ;
        RECT 2.160 4.940 10.060 4.950 ;
        RECT 0.000 4.780 10.060 4.940 ;
        RECT 0.000 4.760 2.560 4.780 ;
        RECT 2.160 4.740 2.470 4.760 ;
        RECT 7.740 4.690 9.280 4.780 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.670 4.950 22.760 5.120 ;
        RECT 22.930 4.950 23.240 5.070 ;
        RECT 15.340 4.940 23.240 4.950 ;
        RECT 15.340 4.780 25.400 4.940 ;
        RECT 16.120 4.690 17.660 4.780 ;
        RECT 22.840 4.760 25.400 4.780 ;
        RECT 22.930 4.740 23.240 4.760 ;
    END
  END ROW1
  PIN ROW2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 2.640 3.940 2.790 4.130 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.640 3.940 22.770 4.120 ;
    END
  END ROW2
  PIN DRAIN1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 2.640 5.370 2.780 5.560 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.670 5.370 22.760 5.550 ;
    END
  END DRAIN1
  PIN DRAIN2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 2.640 3.510 2.770 3.690 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.630 3.510 22.770 3.690 ;
    END
  END DRAIN2
  PIN DRAIN3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 2.640 2.360 2.710 2.540 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.680 2.360 22.770 2.540 ;
    END
  END DRAIN3
  PIN ROW3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 2.640 1.930 2.710 2.110 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.680 1.930 22.770 2.110 ;
    END
  END ROW3
  PIN ROW4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 2.640 0.940 2.710 1.120 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.680 0.940 22.770 1.120 ;
    END
  END ROW4
  PIN DRAIN4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 2.640 0.510 2.710 0.690 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.680 0.510 22.770 0.690 ;
    END
  END DRAIN4
  PIN VGND
    PORT
      LAYER met1 ;
        RECT 5.750 5.960 5.990 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.750 0.000 5.990 0.080 ;
    END
    PORT
      LAYER met1 ;
        RECT 9.680 0.000 9.920 0.070 ;
    END
    PORT
      LAYER nwell ;
        RECT 8.340 8.010 10.070 9.870 ;
        RECT 8.340 6.170 10.080 8.010 ;
        RECT 8.340 3.820 10.070 6.170 ;
      LAYER met1 ;
        RECT 9.320 6.050 9.720 9.870 ;
        RECT 9.320 5.990 9.920 6.050 ;
        RECT 9.320 3.820 9.720 5.990 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.480 0.000 15.720 0.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.410 0.000 19.650 0.060 ;
    END
    PORT
      LAYER nwell ;
        RECT 15.330 8.010 17.060 9.870 ;
        RECT 15.320 6.170 17.060 8.010 ;
        RECT 15.330 3.820 17.060 6.170 ;
      LAYER met1 ;
        RECT 15.680 6.050 16.080 9.870 ;
        RECT 15.480 6.000 16.080 6.050 ;
        RECT 15.680 3.820 16.080 6.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.410 5.980 19.650 6.050 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 0.010 9.860 2.560 9.870 ;
        RECT 0.000 3.840 2.560 9.860 ;
        RECT 0.010 3.830 2.560 3.840 ;
        RECT 4.090 3.820 6.320 9.870 ;
        RECT 19.080 3.820 21.310 9.870 ;
        RECT 22.840 9.860 25.390 9.870 ;
        RECT 22.840 3.840 25.400 9.860 ;
        RECT 22.840 3.830 25.390 3.840 ;
      LAYER li1 ;
        RECT 0.400 9.190 0.600 9.540 ;
        RECT 2.140 9.460 2.460 9.470 ;
        RECT 1.880 9.290 2.460 9.460 ;
        RECT 2.130 9.240 2.460 9.290 ;
        RECT 2.140 9.210 2.460 9.240 ;
        RECT 22.940 9.460 23.260 9.470 ;
        RECT 22.940 9.290 23.520 9.460 ;
        RECT 22.940 9.240 23.270 9.290 ;
        RECT 22.940 9.210 23.260 9.240 ;
        RECT 0.390 9.160 0.600 9.190 ;
        RECT 24.800 9.190 25.000 9.540 ;
        RECT 0.390 8.570 0.610 9.160 ;
        RECT 1.130 8.600 1.330 9.170 ;
        RECT 2.140 8.880 2.460 8.920 ;
        RECT 2.130 8.840 2.460 8.880 ;
        RECT 1.880 8.670 2.460 8.840 ;
        RECT 2.140 8.660 2.460 8.670 ;
        RECT 22.940 8.880 23.260 8.920 ;
        RECT 22.940 8.840 23.270 8.880 ;
        RECT 22.940 8.670 23.520 8.840 ;
        RECT 22.940 8.660 23.260 8.670 ;
        RECT 0.390 7.540 0.610 8.130 ;
        RECT 3.140 8.110 3.310 8.620 ;
        RECT 7.080 8.120 7.250 8.630 ;
        RECT 18.150 8.120 18.320 8.630 ;
        RECT 22.090 8.110 22.260 8.620 ;
        RECT 24.070 8.600 24.270 9.170 ;
        RECT 24.800 9.160 25.010 9.190 ;
        RECT 24.790 8.570 25.010 9.160 ;
        RECT 0.390 7.510 0.600 7.540 ;
        RECT 1.130 7.530 1.330 8.100 ;
        RECT 2.140 8.030 2.460 8.040 ;
        RECT 1.880 7.860 2.460 8.030 ;
        RECT 2.130 7.820 2.460 7.860 ;
        RECT 2.140 7.780 2.460 7.820 ;
        RECT 22.940 8.030 23.260 8.040 ;
        RECT 22.940 7.860 23.520 8.030 ;
        RECT 22.940 7.820 23.270 7.860 ;
        RECT 22.940 7.780 23.260 7.820 ;
        RECT 24.070 7.530 24.270 8.100 ;
        RECT 24.790 7.540 25.010 8.130 ;
        RECT 0.400 7.160 0.600 7.510 ;
        RECT 24.800 7.510 25.010 7.540 ;
        RECT 2.140 7.460 2.460 7.490 ;
        RECT 2.130 7.410 2.460 7.460 ;
        RECT 22.940 7.460 23.260 7.490 ;
        RECT 1.880 7.240 2.460 7.410 ;
        RECT 2.140 7.230 2.460 7.240 ;
        RECT 0.770 6.760 1.210 6.930 ;
        RECT 0.400 6.180 0.600 6.530 ;
        RECT 2.140 6.450 2.460 6.460 ;
        RECT 1.880 6.280 2.460 6.450 ;
        RECT 2.130 6.230 2.460 6.280 ;
        RECT 3.140 6.270 3.310 7.280 ;
        RECT 5.070 6.550 5.620 6.980 ;
        RECT 7.070 6.410 7.240 7.420 ;
        RECT 9.100 6.620 9.650 7.050 ;
        RECT 15.750 6.620 16.300 7.050 ;
        RECT 18.160 6.410 18.330 7.420 ;
        RECT 22.940 7.410 23.270 7.460 ;
        RECT 19.780 6.550 20.330 6.980 ;
        RECT 22.090 6.270 22.260 7.280 ;
        RECT 22.940 7.240 23.520 7.410 ;
        RECT 22.940 7.230 23.260 7.240 ;
        RECT 24.800 7.160 25.000 7.510 ;
        RECT 24.190 6.760 24.630 6.930 ;
        RECT 22.940 6.450 23.260 6.460 ;
        RECT 22.940 6.280 23.520 6.450 ;
        RECT 2.140 6.200 2.460 6.230 ;
        RECT 22.940 6.230 23.270 6.280 ;
        RECT 22.940 6.200 23.260 6.230 ;
        RECT 0.390 6.150 0.600 6.180 ;
        RECT 24.800 6.180 25.000 6.530 ;
        RECT 0.390 5.560 0.610 6.150 ;
        RECT 1.130 5.590 1.330 6.160 ;
        RECT 2.140 5.870 2.460 5.910 ;
        RECT 2.130 5.830 2.460 5.870 ;
        RECT 1.880 5.660 2.460 5.830 ;
        RECT 2.140 5.650 2.460 5.660 ;
        RECT 22.940 5.870 23.260 5.910 ;
        RECT 22.940 5.830 23.270 5.870 ;
        RECT 22.940 5.660 23.520 5.830 ;
        RECT 22.940 5.650 23.260 5.660 ;
        RECT 24.070 5.590 24.270 6.160 ;
        RECT 24.800 6.150 25.010 6.180 ;
        RECT 24.790 5.560 25.010 6.150 ;
        RECT 0.390 4.540 0.610 5.130 ;
        RECT 0.390 4.510 0.600 4.540 ;
        RECT 1.130 4.530 1.330 5.100 ;
        RECT 2.140 5.030 2.460 5.040 ;
        RECT 1.880 4.860 2.460 5.030 ;
        RECT 2.130 4.820 2.460 4.860 ;
        RECT 2.140 4.780 2.460 4.820 ;
        RECT 22.940 5.030 23.260 5.040 ;
        RECT 22.940 4.860 23.520 5.030 ;
        RECT 22.940 4.820 23.270 4.860 ;
        RECT 22.940 4.780 23.260 4.820 ;
        RECT 24.070 4.530 24.270 5.100 ;
        RECT 24.790 4.540 25.010 5.130 ;
        RECT 0.400 4.160 0.600 4.510 ;
        RECT 24.800 4.510 25.010 4.540 ;
        RECT 2.140 4.460 2.460 4.490 ;
        RECT 2.130 4.410 2.460 4.460 ;
        RECT 1.880 4.240 2.460 4.410 ;
        RECT 2.140 4.230 2.460 4.240 ;
        RECT 22.940 4.460 23.260 4.490 ;
        RECT 22.940 4.410 23.270 4.460 ;
        RECT 22.940 4.240 23.520 4.410 ;
        RECT 22.940 4.230 23.260 4.240 ;
        RECT 24.800 4.160 25.000 4.510 ;
      LAYER mcon ;
        RECT 2.230 9.250 2.400 9.420 ;
        RECT 23.000 9.250 23.170 9.420 ;
        RECT 0.420 8.990 0.590 9.160 ;
        RECT 1.150 8.960 1.320 9.130 ;
        RECT 24.080 8.960 24.250 9.130 ;
        RECT 2.230 8.700 2.400 8.870 ;
        RECT 23.000 8.700 23.170 8.870 ;
        RECT 3.140 8.450 3.310 8.620 ;
        RECT 7.080 8.460 7.250 8.630 ;
        RECT 18.150 8.460 18.320 8.630 ;
        RECT 22.090 8.450 22.260 8.620 ;
        RECT 24.810 8.990 24.980 9.160 ;
        RECT 0.420 7.540 0.590 7.710 ;
        RECT 2.230 7.830 2.400 8.000 ;
        RECT 23.000 7.830 23.170 8.000 ;
        RECT 1.150 7.570 1.320 7.740 ;
        RECT 24.080 7.570 24.250 7.740 ;
        RECT 24.810 7.540 24.980 7.710 ;
        RECT 2.230 7.280 2.400 7.450 ;
        RECT 3.140 6.860 3.310 7.030 ;
        RECT 7.070 7.000 7.240 7.170 ;
        RECT 23.000 7.280 23.170 7.450 ;
        RECT 3.140 6.520 3.310 6.690 ;
        RECT 5.350 6.630 5.620 6.900 ;
        RECT 7.070 6.660 7.240 6.830 ;
        RECT 2.230 6.240 2.400 6.410 ;
        RECT 9.380 6.700 9.650 6.970 ;
        RECT 15.750 6.700 16.020 6.970 ;
        RECT 18.160 7.000 18.330 7.170 ;
        RECT 18.160 6.660 18.330 6.830 ;
        RECT 19.780 6.630 20.050 6.900 ;
        RECT 22.090 6.860 22.260 7.030 ;
        RECT 24.450 6.760 24.630 6.930 ;
        RECT 22.090 6.520 22.260 6.690 ;
        RECT 23.000 6.240 23.170 6.410 ;
        RECT 0.420 5.980 0.590 6.150 ;
        RECT 1.150 5.950 1.320 6.120 ;
        RECT 24.080 5.950 24.250 6.120 ;
        RECT 2.230 5.690 2.400 5.860 ;
        RECT 23.000 5.690 23.170 5.860 ;
        RECT 24.810 5.980 24.980 6.150 ;
        RECT 0.420 4.540 0.590 4.710 ;
        RECT 2.230 4.830 2.400 5.000 ;
        RECT 23.000 4.830 23.170 5.000 ;
        RECT 1.150 4.570 1.320 4.740 ;
        RECT 24.080 4.570 24.250 4.740 ;
        RECT 24.810 4.540 24.980 4.710 ;
        RECT 2.230 4.280 2.400 4.450 ;
        RECT 23.000 4.280 23.170 4.450 ;
      LAYER met1 ;
        RECT 0.360 9.220 0.520 9.870 ;
        RECT 0.360 8.670 0.630 9.220 ;
        RECT 0.350 8.620 0.630 8.670 ;
        RECT 0.770 8.880 0.960 9.870 ;
        RECT 1.170 9.190 1.330 9.870 ;
        RECT 1.130 9.170 1.330 9.190 ;
        RECT 2.150 9.180 2.470 9.500 ;
        RECT 1.120 8.930 1.350 9.170 ;
        RECT 0.770 8.760 0.940 8.880 ;
        RECT 0.350 8.530 0.520 8.620 ;
        RECT 0.360 8.170 0.520 8.530 ;
        RECT 0.350 8.080 0.520 8.170 ;
        RECT 0.350 8.030 0.630 8.080 ;
        RECT 0.360 7.480 0.630 8.030 ;
        RECT 0.770 7.940 0.930 8.760 ;
        RECT 1.130 8.710 1.330 8.930 ;
        RECT 1.170 7.990 1.330 8.710 ;
        RECT 2.150 8.630 2.470 8.950 ;
        RECT 0.770 7.820 0.940 7.940 ;
        RECT 0.360 6.210 0.520 7.480 ;
        RECT 0.770 6.960 0.960 7.820 ;
        RECT 1.130 7.770 1.330 7.990 ;
        RECT 1.120 7.530 1.350 7.770 ;
        RECT 2.150 7.750 2.470 8.070 ;
        RECT 5.290 7.950 5.670 9.870 ;
        RECT 7.040 8.690 7.280 9.870 ;
        RECT 18.120 8.690 18.360 9.870 ;
        RECT 7.030 8.030 7.290 8.690 ;
        RECT 18.110 8.030 18.370 8.690 ;
        RECT 1.130 7.510 1.330 7.530 ;
        RECT 0.740 6.730 0.980 6.960 ;
        RECT 0.360 5.660 0.630 6.210 ;
        RECT 0.350 5.610 0.630 5.660 ;
        RECT 0.770 5.870 0.960 6.730 ;
        RECT 1.170 6.180 1.330 7.510 ;
        RECT 2.150 7.200 2.470 7.520 ;
        RECT 1.130 6.160 1.330 6.180 ;
        RECT 2.150 6.170 2.470 6.490 ;
        RECT 1.120 5.920 1.350 6.160 ;
        RECT 5.290 6.090 5.680 7.950 ;
        RECT 0.770 5.750 0.940 5.870 ;
        RECT 0.350 5.520 0.520 5.610 ;
        RECT 0.360 5.170 0.520 5.520 ;
        RECT 0.350 5.080 0.520 5.170 ;
        RECT 0.350 5.030 0.630 5.080 ;
        RECT 0.360 4.480 0.630 5.030 ;
        RECT 0.770 4.940 0.930 5.750 ;
        RECT 1.130 5.700 1.330 5.920 ;
        RECT 1.170 4.990 1.330 5.700 ;
        RECT 2.150 5.620 2.470 5.940 ;
        RECT 0.770 4.820 0.940 4.940 ;
        RECT 0.360 3.830 0.520 4.480 ;
        RECT 0.770 3.830 0.960 4.820 ;
        RECT 1.130 4.770 1.330 4.990 ;
        RECT 1.120 4.530 1.350 4.770 ;
        RECT 2.150 4.750 2.470 5.070 ;
        RECT 1.130 4.510 1.330 4.530 ;
        RECT 1.170 3.830 1.330 4.510 ;
        RECT 2.150 4.200 2.470 4.520 ;
        RECT 5.290 3.820 5.670 6.090 ;
        RECT 7.040 5.420 7.280 8.030 ;
        RECT 12.360 5.690 13.040 5.910 ;
        RECT 18.120 5.420 18.360 8.030 ;
        RECT 19.730 7.950 20.110 9.870 ;
        RECT 22.050 8.710 22.290 9.870 ;
        RECT 22.930 9.180 23.250 9.500 ;
        RECT 24.070 9.190 24.230 9.870 ;
        RECT 24.070 9.170 24.270 9.190 ;
        RECT 22.030 8.050 22.300 8.710 ;
        RECT 22.930 8.630 23.250 8.950 ;
        RECT 24.050 8.930 24.280 9.170 ;
        RECT 24.070 8.710 24.270 8.930 ;
        RECT 24.440 8.880 24.630 9.870 ;
        RECT 24.880 9.220 25.040 9.870 ;
        RECT 24.460 8.760 24.630 8.880 ;
        RECT 19.720 6.090 20.110 7.950 ;
        RECT 7.030 5.100 7.290 5.420 ;
        RECT 18.110 5.100 18.370 5.420 ;
        RECT 7.040 3.820 7.280 5.100 ;
        RECT 18.120 3.820 18.360 5.100 ;
        RECT 19.730 3.820 20.110 6.090 ;
        RECT 22.050 6.050 22.290 8.050 ;
        RECT 22.930 7.750 23.250 8.070 ;
        RECT 24.070 7.990 24.230 8.710 ;
        RECT 24.070 7.770 24.270 7.990 ;
        RECT 24.470 7.940 24.630 8.760 ;
        RECT 24.770 8.670 25.040 9.220 ;
        RECT 24.770 8.620 25.050 8.670 ;
        RECT 24.880 8.530 25.050 8.620 ;
        RECT 24.880 8.170 25.040 8.530 ;
        RECT 24.880 8.080 25.050 8.170 ;
        RECT 24.460 7.820 24.630 7.940 ;
        RECT 24.050 7.530 24.280 7.770 ;
        RECT 22.930 7.200 23.250 7.520 ;
        RECT 24.070 7.510 24.270 7.530 ;
        RECT 22.930 6.170 23.250 6.490 ;
        RECT 24.070 6.180 24.230 7.510 ;
        RECT 24.440 6.960 24.630 7.820 ;
        RECT 24.770 8.030 25.050 8.080 ;
        RECT 24.770 7.480 25.040 8.030 ;
        RECT 24.420 6.730 24.660 6.960 ;
        RECT 24.070 6.160 24.270 6.180 ;
        RECT 21.800 6.000 21.990 6.050 ;
        RECT 22.050 6.010 22.400 6.050 ;
        RECT 22.050 5.710 22.560 6.010 ;
        RECT 22.050 5.460 22.290 5.710 ;
        RECT 22.930 5.620 23.250 5.940 ;
        RECT 24.050 5.920 24.280 6.160 ;
        RECT 24.070 5.700 24.270 5.920 ;
        RECT 24.440 5.870 24.630 6.730 ;
        RECT 24.880 6.210 25.040 7.480 ;
        RECT 24.460 5.750 24.630 5.870 ;
        RECT 22.040 5.140 22.300 5.460 ;
        RECT 22.050 3.820 22.290 5.140 ;
        RECT 22.930 4.750 23.250 5.070 ;
        RECT 24.070 4.990 24.230 5.700 ;
        RECT 24.070 4.770 24.270 4.990 ;
        RECT 24.470 4.940 24.630 5.750 ;
        RECT 24.770 5.660 25.040 6.210 ;
        RECT 24.770 5.610 25.050 5.660 ;
        RECT 24.880 5.520 25.050 5.610 ;
        RECT 24.880 5.170 25.040 5.520 ;
        RECT 24.880 5.080 25.050 5.170 ;
        RECT 24.460 4.820 24.630 4.940 ;
        RECT 24.050 4.530 24.280 4.770 ;
        RECT 22.930 4.200 23.250 4.520 ;
        RECT 24.070 4.510 24.270 4.530 ;
        RECT 24.070 3.830 24.230 4.510 ;
        RECT 24.440 3.830 24.630 4.820 ;
        RECT 24.770 5.030 25.050 5.080 ;
        RECT 24.770 4.480 25.040 5.030 ;
        RECT 24.880 3.830 25.040 4.480 ;
      LAYER via ;
        RECT 2.180 9.210 2.440 9.470 ;
        RECT 2.180 8.660 2.440 8.920 ;
        RECT 2.180 7.780 2.440 8.040 ;
        RECT 2.180 7.230 2.440 7.490 ;
        RECT 2.180 6.200 2.440 6.460 ;
        RECT 2.180 5.650 2.440 5.910 ;
        RECT 2.180 4.780 2.440 5.040 ;
        RECT 2.180 4.230 2.440 4.490 ;
        RECT 22.960 9.210 23.220 9.470 ;
        RECT 22.960 8.660 23.220 8.920 ;
        RECT 7.030 5.130 7.290 5.390 ;
        RECT 18.110 5.130 18.370 5.390 ;
        RECT 22.960 7.780 23.220 8.040 ;
        RECT 22.960 7.230 23.220 7.490 ;
        RECT 22.960 6.200 23.220 6.460 ;
        RECT 22.270 5.730 22.530 5.990 ;
        RECT 22.960 5.650 23.220 5.910 ;
        RECT 22.040 5.170 22.300 5.430 ;
        RECT 22.960 4.780 23.220 5.040 ;
        RECT 22.960 4.230 23.220 4.490 ;
      LAYER met2 ;
        RECT 2.160 9.370 2.470 9.510 ;
        RECT 22.930 9.370 23.240 9.510 ;
        RECT 0.000 9.190 10.070 9.370 ;
        RECT 15.330 9.190 25.400 9.370 ;
        RECT 2.160 9.180 2.470 9.190 ;
        RECT 22.930 9.180 23.240 9.190 ;
        RECT 2.160 8.940 2.470 8.960 ;
        RECT 22.930 8.940 23.240 8.960 ;
        RECT 0.000 8.760 10.070 8.940 ;
        RECT 15.330 8.760 25.400 8.940 ;
        RECT 2.160 8.630 2.470 8.760 ;
        RECT 22.930 8.630 23.240 8.760 ;
        RECT 2.160 7.940 2.470 8.070 ;
        RECT 22.930 7.940 23.240 8.070 ;
        RECT 0.000 7.760 10.080 7.940 ;
        RECT 15.320 7.760 25.400 7.940 ;
        RECT 2.160 7.740 2.470 7.760 ;
        RECT 22.930 7.740 23.240 7.760 ;
        RECT 2.160 7.510 2.470 7.520 ;
        RECT 22.930 7.510 23.240 7.520 ;
        RECT 0.000 7.330 10.080 7.510 ;
        RECT 15.320 7.330 25.400 7.510 ;
        RECT 2.160 7.190 2.470 7.330 ;
        RECT 22.930 7.190 23.240 7.330 ;
        RECT 2.160 6.360 2.470 6.500 ;
        RECT 0.000 6.350 2.470 6.360 ;
        RECT 22.930 6.360 23.240 6.500 ;
        RECT 22.930 6.350 25.400 6.360 ;
        RECT 0.000 6.180 10.060 6.350 ;
        RECT 15.340 6.180 25.400 6.350 ;
        RECT 2.160 6.170 2.470 6.180 ;
        RECT 22.930 6.170 23.240 6.180 ;
        RECT 2.160 4.510 2.470 4.520 ;
        RECT 22.930 4.510 23.240 4.520 ;
        RECT 0.000 4.340 10.060 4.510 ;
        RECT 15.340 4.340 25.400 4.510 ;
        RECT 0.000 4.330 2.470 4.340 ;
        RECT 2.160 4.190 2.470 4.330 ;
        RECT 22.930 4.330 25.400 4.340 ;
        RECT 22.930 4.190 23.240 4.330 ;
        RECT 9.340 1.380 16.100 1.560 ;
  END
END sky130_hilas_swc4x2cell

MACRO sky130_hilas_polyresistorGND
  CLASS CORE ;
  FOREIGN sky130_hilas_polyresistorGND ;
  ORIGIN 0.000 0.000 ;
  SIZE 55.470 BY 10.890 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN INPUT
    PORT
      LAYER met1 ;
        RECT 21.060 10.250 23.470 10.890 ;
        RECT 21.080 8.900 21.490 10.250 ;
    END
  END INPUT
  PIN OUTPUT
    ANTENNADIFFAREA 16.454399 ;
    PORT
      LAYER met2 ;
        RECT 0.000 7.380 55.470 8.770 ;
    END
  END OUTPUT
  PIN VGND
    ANTENNADIFFAREA 16.454399 ;
    PORT
      LAYER met1 ;
        RECT 27.810 9.320 28.220 10.360 ;
        RECT 0.330 8.710 24.700 8.730 ;
        RECT 0.270 8.320 24.700 8.710 ;
        RECT 0.270 0.070 0.680 8.320 ;
        RECT 26.870 0.820 29.230 9.320 ;
        RECT 33.500 8.720 53.790 8.730 ;
        RECT 33.440 8.710 53.790 8.720 ;
        RECT 33.440 8.330 54.730 8.710 ;
        RECT 33.440 8.320 54.700 8.330 ;
        RECT 26.750 0.000 29.230 0.820 ;
      LAYER via ;
        RECT 0.820 8.410 24.620 8.670 ;
        RECT 33.500 8.410 54.360 8.670 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 21.140 9.120 21.360 10.240 ;
        RECT 21.090 8.930 21.420 9.120 ;
        RECT 27.880 8.930 28.120 10.280 ;
        RECT 0.380 8.460 55.120 8.730 ;
        RECT 0.380 8.330 24.720 8.460 ;
        RECT 33.410 8.330 55.120 8.460 ;
        RECT 0.380 0.730 0.550 8.330 ;
        RECT 54.950 1.250 55.120 8.330 ;
        RECT 26.820 0.390 29.030 0.560 ;
      LAYER mcon ;
        RECT 21.170 9.820 21.340 9.990 ;
        RECT 21.170 9.480 21.340 9.650 ;
        RECT 21.170 9.140 21.340 9.310 ;
        RECT 27.920 9.860 28.090 10.030 ;
        RECT 27.920 9.520 28.090 9.690 ;
        RECT 27.920 9.180 28.090 9.350 ;
        RECT 0.720 8.350 24.620 8.520 ;
        RECT 33.500 8.350 54.670 8.520 ;
        RECT 27.160 0.390 27.330 0.560 ;
        RECT 27.500 0.390 27.670 0.560 ;
        RECT 27.840 0.390 28.010 0.560 ;
        RECT 28.180 0.390 28.350 0.560 ;
        RECT 28.520 0.390 28.690 0.560 ;
        RECT 28.860 0.390 29.030 0.560 ;
      LAYER met2 ;
        RECT 0.000 1.080 55.470 2.480 ;
  END
END sky130_hilas_polyresistorGND

MACRO sky130_hilas_swc4x2cellOverlap
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc4x2cellOverlap ;
  ORIGIN 11.920 -7.280 ;
  SIZE 21.790 BY 9.870 ;
  PIN VERT1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT -8.840 13.270 -8.680 13.330 ;
    END
    PORT
      LAYER met1 ;
        RECT -8.840 7.290 -8.680 7.360 ;
    END
  END VERT1
  PIN HORIZ1
    USE ANALOG ;
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT -10.010 12.220 -9.930 12.400 ;
        RECT -9.760 12.230 -9.450 12.350 ;
        RECT -9.760 12.220 -2.570 12.230 ;
        RECT -11.920 12.060 -2.570 12.220 ;
        RECT -11.920 12.040 -9.360 12.060 ;
        RECT -9.760 12.020 -9.450 12.040 ;
    END
    PORT
      LAYER met2 ;
        RECT 7.400 12.230 7.710 12.350 ;
        RECT 0.520 12.220 7.710 12.230 ;
        RECT 7.860 12.220 7.970 12.400 ;
        RECT 0.520 12.060 9.870 12.220 ;
        RECT 7.310 12.040 9.870 12.060 ;
        RECT 7.400 12.020 7.710 12.040 ;
    END
  END HORIZ1
  PIN DRAIN1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -10.010 12.650 -9.930 12.830 ;
    END
    PORT
      LAYER met2 ;
        RECT 7.850 12.650 7.960 12.830 ;
    END
  END DRAIN1
  PIN HORIZ2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -10.010 11.220 -9.930 11.400 ;
    END
    PORT
      LAYER met2 ;
        RECT 7.860 11.220 7.970 11.400 ;
    END
  END HORIZ2
  PIN DRAIN2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -10.010 10.790 -9.930 10.970 ;
    END
    PORT
      LAYER met2 ;
        RECT 7.860 10.790 7.970 10.970 ;
    END
  END DRAIN2
  PIN DRAIN3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -10.010 9.640 -9.940 9.820 ;
    END
    PORT
      LAYER met2 ;
        RECT 7.850 9.640 7.960 9.820 ;
    END
  END DRAIN3
  PIN HORIZ3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -10.010 9.210 -9.940 9.390 ;
    END
    PORT
      LAYER met2 ;
        RECT 7.850 9.210 7.960 9.390 ;
    END
  END HORIZ3
  PIN HORIZ4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -10.010 8.220 -9.940 8.400 ;
    END
    PORT
      LAYER met2 ;
        RECT 7.850 8.220 7.960 8.400 ;
    END
  END HORIZ4
  PIN DRAIN4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -10.010 7.790 -9.940 7.970 ;
    END
  END DRAIN4
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT -9.650 13.270 -9.490 13.330 ;
    END
    PORT
      LAYER met1 ;
        RECT -9.650 7.290 -9.490 7.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 7.440 7.290 7.600 7.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 7.440 13.260 7.600 13.330 ;
    END
  END VINJ
  PIN GATESELECT1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT -9.240 13.270 -9.050 13.330 ;
    END
    PORT
      LAYER met1 ;
        RECT -9.240 7.290 -9.050 7.360 ;
    END
  END GATESELECT1
  PIN VERT2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 6.630 13.260 6.790 13.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.630 7.290 6.790 7.360 ;
    END
  END VERT2
  PIN GATESELECT2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 7.000 13.260 7.190 13.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 7.000 7.290 7.190 7.360 ;
    END
  END GATESELECT2
  PIN DRAIN
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 7.850 7.790 7.960 7.970 ;
    END
  END DRAIN
  PIN GATE2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 3.280 7.280 3.520 13.330 ;
    END
  END GATE2
  PIN GATE1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT -5.570 7.280 -5.320 13.330 ;
    END
  END GATE1
  PIN VTUN
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT -1.960 7.280 -1.660 13.330 ;
    END
    PORT
      LAYER met1 ;
        RECT -0.380 7.280 -0.080 13.330 ;
    END
  END VTUN
  OBS
      LAYER nwell ;
        RECT -11.910 17.140 -5.360 17.150 ;
        RECT -11.920 11.120 -5.360 17.140 ;
        RECT -11.910 11.110 -5.360 11.120 ;
        RECT -9.360 11.100 -5.360 11.110 ;
        RECT 3.310 17.140 9.860 17.150 ;
        RECT 3.310 11.120 9.870 17.140 ;
        RECT 3.310 11.110 9.860 11.120 ;
        RECT 3.310 11.100 7.310 11.110 ;
      LAYER li1 ;
        RECT -11.520 16.470 -11.320 16.820 ;
        RECT -9.780 16.740 -9.460 16.750 ;
        RECT -10.040 16.570 -9.460 16.740 ;
        RECT -9.790 16.520 -9.460 16.570 ;
        RECT -9.780 16.490 -9.460 16.520 ;
        RECT -11.530 16.440 -11.320 16.470 ;
        RECT -11.530 15.850 -11.310 16.440 ;
        RECT -10.790 15.880 -10.590 16.450 ;
        RECT -9.780 16.160 -9.460 16.200 ;
        RECT -9.790 16.120 -9.460 16.160 ;
        RECT -10.040 15.950 -9.460 16.120 ;
        RECT -9.780 15.940 -9.460 15.950 ;
        RECT -9.020 15.840 -5.710 16.820 ;
        RECT -3.800 15.940 -3.630 16.830 ;
        RECT 1.580 15.940 1.750 16.830 ;
        RECT 3.660 15.840 6.970 16.820 ;
        RECT 7.410 16.740 7.730 16.750 ;
        RECT 7.410 16.570 7.990 16.740 ;
        RECT 7.410 16.520 7.740 16.570 ;
        RECT 7.410 16.490 7.730 16.520 ;
        RECT 9.270 16.470 9.470 16.820 ;
        RECT 7.410 16.160 7.730 16.200 ;
        RECT 7.410 16.120 7.740 16.160 ;
        RECT 7.410 15.950 7.990 16.120 ;
        RECT 7.410 15.940 7.730 15.950 ;
        RECT 8.540 15.880 8.740 16.450 ;
        RECT 9.270 16.440 9.480 16.470 ;
        RECT 9.260 15.850 9.480 16.440 ;
        RECT -11.530 14.820 -11.310 15.410 ;
        RECT -11.530 14.790 -11.320 14.820 ;
        RECT -10.790 14.810 -10.590 15.380 ;
        RECT -9.780 15.310 -9.460 15.320 ;
        RECT -10.040 15.140 -9.460 15.310 ;
        RECT -9.790 15.100 -9.460 15.140 ;
        RECT -9.780 15.060 -9.460 15.100 ;
        RECT -11.520 14.440 -11.320 14.790 ;
        RECT -9.780 14.740 -9.460 14.770 ;
        RECT -9.790 14.690 -9.460 14.740 ;
        RECT -10.040 14.520 -9.460 14.690 ;
        RECT -9.780 14.510 -9.460 14.520 ;
        RECT -9.020 14.370 -5.710 15.350 ;
        RECT -3.800 14.420 -3.630 15.310 ;
        RECT 1.580 14.420 1.750 15.310 ;
        RECT 3.660 14.370 6.970 15.350 ;
        RECT 7.410 15.310 7.730 15.320 ;
        RECT 7.410 15.140 7.990 15.310 ;
        RECT 7.410 15.100 7.740 15.140 ;
        RECT 7.410 15.060 7.730 15.100 ;
        RECT 8.540 14.810 8.740 15.380 ;
        RECT 9.260 14.820 9.480 15.410 ;
        RECT 9.270 14.790 9.480 14.820 ;
        RECT 7.410 14.740 7.730 14.770 ;
        RECT 7.410 14.690 7.740 14.740 ;
        RECT 7.410 14.520 7.990 14.690 ;
        RECT 7.410 14.510 7.730 14.520 ;
        RECT 9.270 14.440 9.470 14.790 ;
        RECT -11.150 14.040 -10.710 14.210 ;
        RECT 8.660 14.040 9.100 14.210 ;
        RECT -11.520 13.460 -11.320 13.810 ;
        RECT -9.780 13.730 -9.460 13.740 ;
        RECT -10.040 13.560 -9.460 13.730 ;
        RECT -9.790 13.510 -9.460 13.560 ;
        RECT -9.780 13.480 -9.460 13.510 ;
        RECT -11.530 13.430 -11.320 13.460 ;
        RECT -11.530 12.840 -11.310 13.430 ;
        RECT -10.790 12.870 -10.590 13.440 ;
        RECT -9.780 13.150 -9.460 13.190 ;
        RECT -9.790 13.110 -9.460 13.150 ;
        RECT -10.040 12.940 -9.460 13.110 ;
        RECT -9.780 12.930 -9.460 12.940 ;
        RECT -9.020 12.900 -5.710 13.880 ;
        RECT -3.800 12.970 -3.630 13.860 ;
        RECT 1.580 12.970 1.750 13.860 ;
        RECT 3.660 12.900 6.970 13.880 ;
        RECT 7.410 13.730 7.730 13.740 ;
        RECT 7.410 13.560 7.990 13.730 ;
        RECT 7.410 13.510 7.740 13.560 ;
        RECT 7.410 13.480 7.730 13.510 ;
        RECT 9.270 13.460 9.470 13.810 ;
        RECT 7.410 13.150 7.730 13.190 ;
        RECT 7.410 13.110 7.740 13.150 ;
        RECT 7.410 12.940 7.990 13.110 ;
        RECT 7.410 12.930 7.730 12.940 ;
        RECT 8.540 12.870 8.740 13.440 ;
        RECT 9.270 13.430 9.480 13.460 ;
        RECT 9.260 12.840 9.480 13.430 ;
        RECT -11.530 11.820 -11.310 12.410 ;
        RECT -11.530 11.790 -11.320 11.820 ;
        RECT -10.790 11.810 -10.590 12.380 ;
        RECT -9.780 12.310 -9.460 12.320 ;
        RECT -10.040 12.140 -9.460 12.310 ;
        RECT -9.790 12.100 -9.460 12.140 ;
        RECT -9.780 12.060 -9.460 12.100 ;
        RECT -11.520 11.440 -11.320 11.790 ;
        RECT -9.780 11.740 -9.460 11.770 ;
        RECT -9.790 11.690 -9.460 11.740 ;
        RECT -10.040 11.520 -9.460 11.690 ;
        RECT -9.780 11.510 -9.460 11.520 ;
        RECT -9.020 11.430 -5.710 12.410 ;
        RECT -3.800 11.430 -3.630 12.320 ;
        RECT 1.580 11.430 1.750 12.320 ;
        RECT 3.660 11.430 6.970 12.410 ;
        RECT 7.410 12.310 7.730 12.320 ;
        RECT 7.410 12.140 7.990 12.310 ;
        RECT 7.410 12.100 7.740 12.140 ;
        RECT 7.410 12.060 7.730 12.100 ;
        RECT 8.540 11.810 8.740 12.380 ;
        RECT 9.260 11.820 9.480 12.410 ;
        RECT 9.270 11.790 9.480 11.820 ;
        RECT 7.410 11.740 7.730 11.770 ;
        RECT 7.410 11.690 7.740 11.740 ;
        RECT 7.410 11.520 7.990 11.690 ;
        RECT 7.410 11.510 7.730 11.520 ;
        RECT 9.270 11.440 9.470 11.790 ;
      LAYER mcon ;
        RECT -9.690 16.530 -9.520 16.700 ;
        RECT -7.450 16.590 -7.280 16.760 ;
        RECT -11.500 16.270 -11.330 16.440 ;
        RECT -10.770 16.240 -10.600 16.410 ;
        RECT -7.450 16.240 -7.280 16.410 ;
        RECT -9.690 15.980 -9.520 16.150 ;
        RECT -7.450 15.900 -7.280 16.070 ;
        RECT -3.800 16.630 -3.630 16.800 ;
        RECT 1.580 16.630 1.750 16.800 ;
        RECT 5.230 16.590 5.400 16.760 ;
        RECT 7.470 16.530 7.640 16.700 ;
        RECT 5.230 16.240 5.400 16.410 ;
        RECT 8.550 16.240 8.720 16.410 ;
        RECT 5.230 15.900 5.400 16.070 ;
        RECT 7.470 15.980 7.640 16.150 ;
        RECT 9.280 16.270 9.450 16.440 ;
        RECT -11.500 14.820 -11.330 14.990 ;
        RECT -9.690 15.110 -9.520 15.280 ;
        RECT -7.450 15.120 -7.280 15.290 ;
        RECT -10.770 14.850 -10.600 15.020 ;
        RECT -7.450 14.770 -7.280 14.940 ;
        RECT -9.690 14.560 -9.520 14.730 ;
        RECT -7.450 14.430 -7.280 14.600 ;
        RECT -3.800 15.110 -3.630 15.280 ;
        RECT 1.580 15.110 1.750 15.280 ;
        RECT 5.230 15.120 5.400 15.290 ;
        RECT 7.470 15.110 7.640 15.280 ;
        RECT 5.230 14.770 5.400 14.940 ;
        RECT 8.550 14.850 8.720 15.020 ;
        RECT 9.280 14.820 9.450 14.990 ;
        RECT 5.230 14.430 5.400 14.600 ;
        RECT 7.470 14.560 7.640 14.730 ;
        RECT 8.920 14.040 9.100 14.210 ;
        RECT -9.690 13.520 -9.520 13.690 ;
        RECT -7.450 13.650 -7.280 13.820 ;
        RECT -11.500 13.260 -11.330 13.430 ;
        RECT -10.770 13.230 -10.600 13.400 ;
        RECT -7.450 13.300 -7.280 13.470 ;
        RECT -9.690 12.970 -9.520 13.140 ;
        RECT -7.450 12.960 -7.280 13.130 ;
        RECT -3.800 13.660 -3.630 13.830 ;
        RECT 1.580 13.660 1.750 13.830 ;
        RECT 5.230 13.650 5.400 13.820 ;
        RECT 7.470 13.520 7.640 13.690 ;
        RECT 5.230 13.300 5.400 13.470 ;
        RECT 8.550 13.230 8.720 13.400 ;
        RECT 5.230 12.960 5.400 13.130 ;
        RECT 7.470 12.970 7.640 13.140 ;
        RECT 9.280 13.260 9.450 13.430 ;
        RECT -11.500 11.820 -11.330 11.990 ;
        RECT -9.690 12.110 -9.520 12.280 ;
        RECT -7.450 12.180 -7.280 12.350 ;
        RECT -10.770 11.850 -10.600 12.020 ;
        RECT -7.450 11.830 -7.280 12.000 ;
        RECT -9.690 11.560 -9.520 11.730 ;
        RECT -7.450 11.490 -7.280 11.660 ;
        RECT -3.800 12.120 -3.630 12.290 ;
        RECT 1.580 12.120 1.750 12.290 ;
        RECT 5.230 12.180 5.400 12.350 ;
        RECT 7.470 12.110 7.640 12.280 ;
        RECT 5.230 11.830 5.400 12.000 ;
        RECT 8.550 11.850 8.720 12.020 ;
        RECT 9.280 11.820 9.450 11.990 ;
        RECT 5.230 11.490 5.400 11.660 ;
        RECT 7.470 11.560 7.640 11.730 ;
      LAYER met1 ;
        RECT -11.560 16.500 -11.400 17.150 ;
        RECT -11.560 15.950 -11.290 16.500 ;
        RECT -11.570 15.900 -11.290 15.950 ;
        RECT -11.150 16.160 -10.960 17.150 ;
        RECT -10.750 16.470 -10.590 17.150 ;
        RECT -10.790 16.450 -10.590 16.470 ;
        RECT -9.770 16.460 -9.450 16.780 ;
        RECT -10.800 16.210 -10.570 16.450 ;
        RECT -11.150 16.040 -10.980 16.160 ;
        RECT -11.570 15.810 -11.400 15.900 ;
        RECT -11.560 15.450 -11.400 15.810 ;
        RECT -11.570 15.360 -11.400 15.450 ;
        RECT -11.570 15.310 -11.290 15.360 ;
        RECT -11.560 14.760 -11.290 15.310 ;
        RECT -11.150 15.220 -10.990 16.040 ;
        RECT -10.790 15.990 -10.590 16.210 ;
        RECT -10.750 15.270 -10.590 15.990 ;
        RECT -9.770 15.910 -9.450 16.230 ;
        RECT -7.480 16.180 -7.240 16.820 ;
        RECT -7.480 15.920 -7.250 16.180 ;
        RECT -7.490 15.700 -7.250 15.920 ;
        RECT -11.150 15.100 -10.980 15.220 ;
        RECT -11.560 13.490 -11.400 14.760 ;
        RECT -11.150 14.240 -10.960 15.100 ;
        RECT -10.790 15.050 -10.590 15.270 ;
        RECT -10.800 14.810 -10.570 15.050 ;
        RECT -9.770 15.030 -9.450 15.350 ;
        RECT -10.790 14.790 -10.590 14.810 ;
        RECT -11.180 14.010 -10.940 14.240 ;
        RECT -11.560 12.940 -11.290 13.490 ;
        RECT -11.570 12.890 -11.290 12.940 ;
        RECT -11.150 13.150 -10.960 14.010 ;
        RECT -10.750 13.460 -10.590 14.790 ;
        RECT -9.770 14.480 -9.450 14.800 ;
        RECT -7.480 14.710 -7.240 15.350 ;
        RECT -7.480 14.450 -7.250 14.710 ;
        RECT -7.490 14.230 -7.250 14.450 ;
        RECT -10.790 13.440 -10.590 13.460 ;
        RECT -9.770 13.450 -9.450 13.770 ;
        RECT -10.800 13.200 -10.570 13.440 ;
        RECT -7.480 13.240 -7.240 13.880 ;
        RECT -11.150 13.030 -10.980 13.150 ;
        RECT -11.570 12.800 -11.400 12.890 ;
        RECT -11.560 12.450 -11.400 12.800 ;
        RECT -11.570 12.360 -11.400 12.450 ;
        RECT -11.570 12.310 -11.290 12.360 ;
        RECT -11.560 11.760 -11.290 12.310 ;
        RECT -11.150 12.220 -10.990 13.030 ;
        RECT -10.790 12.980 -10.590 13.200 ;
        RECT -10.750 12.270 -10.590 12.980 ;
        RECT -9.770 12.900 -9.450 13.220 ;
        RECT -7.480 12.980 -7.250 13.240 ;
        RECT -7.490 12.760 -7.250 12.980 ;
        RECT -11.150 12.100 -10.980 12.220 ;
        RECT -11.560 11.110 -11.400 11.760 ;
        RECT -11.150 11.110 -10.960 12.100 ;
        RECT -10.790 12.050 -10.590 12.270 ;
        RECT -10.800 11.810 -10.570 12.050 ;
        RECT -9.770 12.030 -9.450 12.350 ;
        RECT -10.790 11.790 -10.590 11.810 ;
        RECT -10.750 11.110 -10.590 11.790 ;
        RECT -9.770 11.480 -9.450 11.800 ;
        RECT -7.480 11.770 -7.240 12.410 ;
        RECT -7.480 11.510 -7.250 11.770 ;
        RECT -7.490 11.290 -7.250 11.510 ;
        RECT -3.850 11.100 -3.580 17.150 ;
        RECT 1.530 11.100 1.800 17.150 ;
        RECT 5.190 16.180 5.430 16.820 ;
        RECT 7.400 16.460 7.720 16.780 ;
        RECT 8.540 16.470 8.700 17.150 ;
        RECT 8.540 16.450 8.740 16.470 ;
        RECT 5.200 15.920 5.430 16.180 ;
        RECT 5.200 15.700 5.440 15.920 ;
        RECT 7.400 15.910 7.720 16.230 ;
        RECT 8.520 16.210 8.750 16.450 ;
        RECT 8.540 15.990 8.740 16.210 ;
        RECT 8.910 16.160 9.100 17.150 ;
        RECT 9.350 16.500 9.510 17.150 ;
        RECT 8.930 16.040 9.100 16.160 ;
        RECT 5.190 14.710 5.430 15.350 ;
        RECT 7.400 15.030 7.720 15.350 ;
        RECT 8.540 15.270 8.700 15.990 ;
        RECT 8.540 15.050 8.740 15.270 ;
        RECT 8.940 15.220 9.100 16.040 ;
        RECT 9.240 15.950 9.510 16.500 ;
        RECT 9.240 15.900 9.520 15.950 ;
        RECT 9.350 15.810 9.520 15.900 ;
        RECT 9.350 15.450 9.510 15.810 ;
        RECT 9.350 15.360 9.520 15.450 ;
        RECT 8.930 15.100 9.100 15.220 ;
        RECT 8.520 14.810 8.750 15.050 ;
        RECT 5.200 14.450 5.430 14.710 ;
        RECT 7.400 14.480 7.720 14.800 ;
        RECT 8.540 14.790 8.740 14.810 ;
        RECT 5.200 14.230 5.440 14.450 ;
        RECT 5.190 13.240 5.430 13.880 ;
        RECT 7.400 13.450 7.720 13.770 ;
        RECT 8.540 13.460 8.700 14.790 ;
        RECT 8.910 14.240 9.100 15.100 ;
        RECT 9.240 15.310 9.520 15.360 ;
        RECT 9.240 14.760 9.510 15.310 ;
        RECT 8.890 14.010 9.130 14.240 ;
        RECT 8.540 13.440 8.740 13.460 ;
        RECT 5.200 12.980 5.430 13.240 ;
        RECT 5.200 12.760 5.440 12.980 ;
        RECT 7.400 12.900 7.720 13.220 ;
        RECT 8.520 13.200 8.750 13.440 ;
        RECT 8.540 12.980 8.740 13.200 ;
        RECT 8.910 13.150 9.100 14.010 ;
        RECT 9.350 13.490 9.510 14.760 ;
        RECT 8.930 13.030 9.100 13.150 ;
        RECT 5.190 11.770 5.430 12.410 ;
        RECT 7.400 12.030 7.720 12.350 ;
        RECT 8.540 12.270 8.700 12.980 ;
        RECT 8.540 12.050 8.740 12.270 ;
        RECT 8.940 12.220 9.100 13.030 ;
        RECT 9.240 12.940 9.510 13.490 ;
        RECT 9.240 12.890 9.520 12.940 ;
        RECT 9.350 12.800 9.520 12.890 ;
        RECT 9.350 12.450 9.510 12.800 ;
        RECT 9.350 12.360 9.520 12.450 ;
        RECT 8.930 12.100 9.100 12.220 ;
        RECT 8.520 11.810 8.750 12.050 ;
        RECT 5.200 11.510 5.430 11.770 ;
        RECT 5.200 11.290 5.440 11.510 ;
        RECT 7.400 11.480 7.720 11.800 ;
        RECT 8.540 11.790 8.740 11.810 ;
        RECT 8.540 11.110 8.700 11.790 ;
        RECT 8.910 11.110 9.100 12.100 ;
        RECT 9.240 12.310 9.520 12.360 ;
        RECT 9.240 11.760 9.510 12.310 ;
        RECT 9.350 11.110 9.510 11.760 ;
      LAYER via ;
        RECT -9.740 16.490 -9.480 16.750 ;
        RECT -9.740 15.940 -9.480 16.200 ;
        RECT -9.740 15.060 -9.480 15.320 ;
        RECT -9.740 14.510 -9.480 14.770 ;
        RECT -9.740 13.480 -9.480 13.740 ;
        RECT -9.740 12.930 -9.480 13.190 ;
        RECT -9.740 12.060 -9.480 12.320 ;
        RECT -9.740 11.510 -9.480 11.770 ;
        RECT 7.430 16.490 7.690 16.750 ;
        RECT 7.430 15.940 7.690 16.200 ;
        RECT 7.430 15.060 7.690 15.320 ;
        RECT 7.430 14.510 7.690 14.770 ;
        RECT 7.430 13.480 7.690 13.740 ;
        RECT 7.430 12.930 7.690 13.190 ;
        RECT 7.430 12.060 7.690 12.320 ;
        RECT 7.430 11.510 7.690 11.770 ;
      LAYER met2 ;
        RECT -9.760 16.650 -9.450 16.790 ;
        RECT 7.400 16.650 7.710 16.790 ;
        RECT -11.920 16.470 -2.570 16.650 ;
        RECT 0.520 16.470 9.870 16.650 ;
        RECT -9.760 16.460 -9.450 16.470 ;
        RECT 7.400 16.460 7.710 16.470 ;
        RECT -9.760 16.220 -9.450 16.240 ;
        RECT 7.400 16.220 7.710 16.240 ;
        RECT -11.920 16.040 -2.570 16.220 ;
        RECT 0.520 16.040 9.870 16.220 ;
        RECT -9.760 15.910 -9.450 16.040 ;
        RECT 7.400 15.910 7.710 16.040 ;
        RECT -9.760 15.220 -9.450 15.350 ;
        RECT 7.400 15.220 7.710 15.350 ;
        RECT -11.920 15.040 -2.570 15.220 ;
        RECT 0.520 15.040 9.870 15.220 ;
        RECT -9.760 15.020 -9.450 15.040 ;
        RECT 7.400 15.020 7.710 15.040 ;
        RECT -9.760 14.790 -9.450 14.800 ;
        RECT 7.400 14.790 7.710 14.800 ;
        RECT -11.920 14.720 -9.450 14.790 ;
        RECT -9.440 14.720 -2.570 14.790 ;
        RECT -11.920 14.610 -2.570 14.720 ;
        RECT 0.520 14.720 7.390 14.790 ;
        RECT 7.400 14.720 9.870 14.790 ;
        RECT 0.520 14.610 9.870 14.720 ;
        RECT -9.760 14.470 -9.450 14.610 ;
        RECT 7.400 14.470 7.710 14.610 ;
        RECT -9.760 13.640 -9.450 13.780 ;
        RECT -11.920 13.630 -9.450 13.640 ;
        RECT 7.400 13.640 7.710 13.780 ;
        RECT 7.400 13.630 9.870 13.640 ;
        RECT -11.920 13.460 -2.570 13.630 ;
        RECT 0.520 13.460 9.870 13.630 ;
        RECT -9.760 13.450 -9.450 13.460 ;
        RECT 7.400 13.450 7.710 13.460 ;
        RECT -9.760 13.210 -9.450 13.230 ;
        RECT 7.400 13.210 7.710 13.230 ;
        RECT -11.920 13.040 -2.570 13.210 ;
        RECT 0.520 13.040 9.870 13.210 ;
        RECT -11.920 13.030 -9.360 13.040 ;
        RECT 7.310 13.030 9.870 13.040 ;
        RECT -9.760 12.900 -9.450 13.030 ;
        RECT 7.400 12.900 7.710 13.030 ;
        RECT -9.760 11.790 -9.450 11.800 ;
        RECT 7.400 11.790 7.710 11.800 ;
        RECT -11.920 11.620 -2.570 11.790 ;
        RECT 0.520 11.620 9.870 11.790 ;
        RECT -11.920 11.610 -9.450 11.620 ;
        RECT -9.760 11.470 -9.450 11.610 ;
        RECT 7.400 11.610 9.870 11.620 ;
        RECT 7.400 11.470 7.710 11.610 ;
        RECT -7.610 10.890 -7.490 10.970 ;
        RECT 5.480 10.830 5.600 10.970 ;
  END
END sky130_hilas_swc4x2cellOverlap

MACRO sky130_hilas_FGBias2x1cell
  CLASS CORE ;
  FOREIGN sky130_hilas_FGBias2x1cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.530 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 2.516100 ;
    PORT
      LAYER nwell ;
        RECT 0.010 5.300 1.740 6.050 ;
        RECT 0.010 1.730 1.750 5.300 ;
        RECT 0.010 0.010 1.740 1.730 ;
      LAYER met1 ;
        RECT 0.350 0.000 0.770 6.050 ;
    END
  END VTUN
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2.830 0.000 3.060 6.050 ;
    END
  END VGND
  PIN GATE_CONTROL
    USE ANALOG ;
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT 3.770 3.660 6.490 5.310 ;
        RECT 3.770 3.620 6.480 3.660 ;
        RECT 3.770 2.290 6.480 2.330 ;
        RECT 3.770 0.640 6.490 2.290 ;
      LAYER met1 ;
        RECT 4.050 4.840 4.280 6.050 ;
        RECT 4.050 4.050 4.310 4.840 ;
        RECT 4.050 1.900 4.280 4.050 ;
        RECT 4.050 1.110 4.310 1.900 ;
        RECT 4.050 0.000 4.280 1.110 ;
    END
  END GATE_CONTROL
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.105400 ;
    PORT
      LAYER met2 ;
        RECT 9.050 5.550 9.360 5.560 ;
        RECT 0.000 5.370 11.530 5.550 ;
        RECT 9.050 5.230 9.360 5.370 ;
    END
  END DRAIN1
  PIN DRAIN4
    USE ANALOG ;
    ANTENNADIFFAREA 0.105400 ;
    PORT
      LAYER met2 ;
        RECT 9.050 0.680 9.360 0.820 ;
        RECT 9.050 0.670 11.530 0.680 ;
        RECT 0.000 0.520 11.530 0.670 ;
        RECT 9.050 0.500 11.530 0.520 ;
        RECT 9.050 0.490 9.360 0.500 ;
    END
  END DRAIN4
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 8.220 0.010 11.530 6.050 ;
      LAYER met2 ;
        RECT 10.140 3.190 10.460 3.450 ;
        RECT 10.180 3.170 11.360 3.190 ;
        RECT 10.180 2.910 11.400 3.170 ;
        RECT 10.180 2.850 11.360 2.910 ;
        RECT 10.140 2.840 11.360 2.850 ;
        RECT 10.140 2.590 10.460 2.840 ;
    END
  END VINJ
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 9.200 4.530 9.510 4.600 ;
        RECT 9.200 4.310 11.530 4.530 ;
        RECT 9.200 4.270 9.510 4.310 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 9.200 1.770 9.510 1.840 ;
        RECT 9.200 1.560 11.530 1.770 ;
        RECT 9.200 1.510 9.510 1.560 ;
    END
  END OUTPUT2
  PIN GATECOL
    ANTENNAGATEAREA 0.310000 ;
    PORT
      LAYER met1 ;
        RECT 10.570 4.590 10.760 6.050 ;
        RECT 10.570 4.560 10.790 4.590 ;
        RECT 10.550 4.290 10.800 4.560 ;
        RECT 10.560 4.280 10.800 4.290 ;
        RECT 10.560 4.040 10.790 4.280 ;
        RECT 10.600 2.010 10.760 4.040 ;
        RECT 10.560 1.770 10.790 2.010 ;
        RECT 10.560 1.760 10.800 1.770 ;
        RECT 10.550 1.490 10.800 1.760 ;
        RECT 10.570 1.460 10.790 1.490 ;
        RECT 10.570 0.000 10.760 1.460 ;
    END
  END GATECOL
  PIN VINJ
    ANTENNADIFFAREA 0.510000 ;
    PORT
      LAYER met1 ;
        RECT 11.010 5.400 11.290 6.050 ;
        RECT 10.900 4.800 11.290 5.400 ;
        RECT 11.010 3.200 11.290 4.800 ;
        RECT 11.010 2.880 11.370 3.200 ;
        RECT 11.010 1.250 11.290 2.880 ;
        RECT 10.900 0.650 11.290 1.250 ;
        RECT 11.010 0.000 11.290 0.650 ;
      LAYER via ;
        RECT 11.110 2.910 11.370 3.170 ;
    END
  END VINJ
  OBS
      LAYER li1 ;
        RECT 9.120 5.470 9.650 5.640 ;
        RECT 10.930 5.370 11.130 5.720 ;
        RECT 10.930 5.340 11.140 5.370 ;
        RECT 7.250 4.890 7.600 5.060 ;
        RECT 8.620 4.890 8.950 5.060 ;
        RECT 0.440 3.910 0.990 4.340 ;
        RECT 4.070 4.100 4.300 4.790 ;
        RECT 9.370 4.560 9.540 5.080 ;
        RECT 9.210 4.300 9.540 4.560 ;
        RECT 7.250 4.100 7.600 4.270 ;
        RECT 8.620 4.100 8.950 4.270 ;
        RECT 3.040 3.080 3.230 3.480 ;
        RECT 7.260 3.310 7.600 3.480 ;
        RECT 8.620 3.310 8.950 3.480 ;
        RECT 9.370 3.390 9.540 4.300 ;
        RECT 10.200 3.480 10.370 5.090 ;
        RECT 10.920 4.760 11.140 5.340 ;
        RECT 10.930 4.750 11.140 4.760 ;
        RECT 10.570 4.580 10.760 4.590 ;
        RECT 10.570 4.290 10.770 4.580 ;
        RECT 10.560 3.960 10.800 4.290 ;
        RECT 2.850 3.070 3.230 3.080 ;
        RECT 2.850 2.890 6.590 3.070 ;
        RECT 2.850 2.850 3.230 2.890 ;
        RECT 0.440 2.180 0.990 2.610 ;
        RECT 3.040 2.470 3.230 2.850 ;
        RECT 8.700 2.740 8.870 3.310 ;
        RECT 10.200 3.290 10.380 3.480 ;
        RECT 7.260 2.570 7.600 2.740 ;
        RECT 8.620 2.570 8.950 2.740 ;
        RECT 4.070 1.160 4.300 1.890 ;
        RECT 7.250 1.780 7.600 1.950 ;
        RECT 8.620 1.780 8.950 1.950 ;
        RECT 9.370 1.800 9.540 2.660 ;
        RECT 9.210 1.540 9.540 1.800 ;
        RECT 7.250 0.990 7.600 1.160 ;
        RECT 8.620 0.990 8.950 1.160 ;
        RECT 9.370 0.970 9.540 1.540 ;
        RECT 10.200 2.570 10.380 2.760 ;
        RECT 10.200 0.960 10.370 2.570 ;
        RECT 10.560 1.760 10.800 2.090 ;
        RECT 10.570 1.470 10.770 1.760 ;
        RECT 10.570 1.460 10.760 1.470 ;
        RECT 10.930 1.290 11.140 1.300 ;
        RECT 10.920 0.710 11.140 1.290 ;
        RECT 10.930 0.680 11.140 0.710 ;
        RECT 9.120 0.410 9.650 0.580 ;
        RECT 10.930 0.330 11.130 0.680 ;
      LAYER mcon ;
        RECT 10.940 5.170 11.110 5.340 ;
        RECT 4.100 4.590 4.270 4.760 ;
        RECT 0.440 3.990 0.710 4.260 ;
        RECT 4.100 4.140 4.270 4.310 ;
        RECT 9.270 4.340 9.440 4.510 ;
        RECT 10.580 4.330 10.760 4.520 ;
        RECT 2.860 2.880 3.030 3.050 ;
        RECT 0.440 2.260 0.710 2.530 ;
        RECT 4.100 1.640 4.270 1.810 ;
        RECT 9.270 1.580 9.440 1.750 ;
        RECT 4.100 1.190 4.270 1.360 ;
        RECT 10.580 1.530 10.760 1.720 ;
        RECT 10.940 0.710 11.110 0.880 ;
      LAYER met1 ;
        RECT 9.050 5.230 9.360 5.670 ;
        RECT 9.200 4.270 9.520 4.590 ;
        RECT 10.170 3.480 10.410 3.610 ;
        RECT 10.170 3.160 10.430 3.480 ;
        RECT 10.170 2.560 10.430 2.880 ;
        RECT 10.170 2.440 10.410 2.560 ;
        RECT 9.200 1.510 9.520 1.830 ;
        RECT 9.050 0.380 9.360 0.820 ;
      LAYER via ;
        RECT 9.080 5.260 9.340 5.520 ;
        RECT 9.230 4.300 9.490 4.560 ;
        RECT 10.170 3.190 10.430 3.450 ;
        RECT 10.170 2.590 10.430 2.850 ;
        RECT 9.230 1.540 9.490 1.800 ;
        RECT 9.080 0.530 9.340 0.790 ;
  END
END sky130_hilas_FGBias2x1cell

MACRO sky130_hilas_drainSelect01
  CLASS CORE ;
  FOREIGN sky130_hilas_drainSelect01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.720 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DRAIN4
    ANTENNADIFFAREA 0.275800 ;
    PORT
      LAYER met2 ;
        RECT 0.050 0.690 0.570 0.700 ;
        RECT 0.050 0.620 2.030 0.690 ;
        RECT 0.050 0.570 2.070 0.620 ;
        RECT 4.160 0.570 4.480 0.650 ;
        RECT 0.050 0.520 4.480 0.570 ;
        RECT 1.750 0.380 4.480 0.520 ;
        RECT 1.750 0.360 2.070 0.380 ;
        RECT 4.160 0.330 4.480 0.380 ;
    END
  END DRAIN4
  PIN DRAIN3
    ANTENNADIFFAREA 0.275800 ;
    PORT
      LAYER met2 ;
        RECT 1.750 2.740 2.070 2.760 ;
        RECT 4.160 2.740 4.480 2.790 ;
        RECT 1.750 2.550 4.480 2.740 ;
        RECT 0.050 2.530 0.570 2.540 ;
        RECT 0.050 2.520 1.270 2.530 ;
        RECT 1.750 2.520 2.070 2.550 ;
        RECT 0.050 2.500 2.070 2.520 ;
        RECT 0.050 2.360 2.000 2.500 ;
        RECT 4.160 2.470 4.480 2.550 ;
    END
  END DRAIN3
  PIN DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.275800 ;
    PORT
      LAYER met2 ;
        RECT 0.050 3.670 1.240 3.690 ;
        RECT 0.050 3.550 1.960 3.670 ;
        RECT 0.050 3.510 2.070 3.550 ;
        RECT 1.750 3.500 2.070 3.510 ;
        RECT 4.160 3.500 4.480 3.580 ;
        RECT 1.750 3.310 4.480 3.500 ;
        RECT 1.750 3.290 2.070 3.310 ;
        RECT 4.160 3.260 4.480 3.310 ;
    END
  END DRAIN2
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.275800 ;
    PORT
      LAYER met2 ;
        RECT 1.750 5.670 2.070 5.690 ;
        RECT 4.160 5.670 4.480 5.720 ;
        RECT 0.050 5.540 1.300 5.550 ;
        RECT 1.750 5.540 4.480 5.670 ;
        RECT 0.050 5.480 4.480 5.540 ;
        RECT 0.050 5.430 2.070 5.480 ;
        RECT 0.050 5.380 1.990 5.430 ;
        RECT 4.160 5.400 4.480 5.480 ;
        RECT 0.050 5.370 1.300 5.380 ;
    END
  END DRAIN1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.000 0.000 3.420 6.050 ;
      LAYER met1 ;
        RECT 0.580 5.830 0.830 6.050 ;
        RECT 0.190 4.760 0.830 5.830 ;
        RECT 0.580 4.220 0.830 4.760 ;
        RECT 0.190 3.150 0.830 4.220 ;
        RECT 0.580 2.900 0.830 3.150 ;
        RECT 0.190 1.830 0.830 2.900 ;
        RECT 0.580 1.290 0.830 1.830 ;
        RECT 0.190 0.220 0.830 1.290 ;
        RECT 0.580 0.000 0.830 0.220 ;
    END
  END VINJ
  PIN DRAIN_MUX
    USE ANALOG ;
    ANTENNADIFFAREA 0.719200 ;
    PORT
      LAYER met1 ;
        RECT 3.570 0.000 3.800 6.050 ;
    END
  END DRAIN_MUX
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 4.920 5.830 5.110 6.050 ;
        RECT 4.920 5.340 5.390 5.830 ;
        RECT 4.920 5.080 5.110 5.340 ;
        RECT 4.880 4.790 5.110 5.080 ;
        RECT 4.920 4.190 5.110 4.790 ;
        RECT 4.880 3.900 5.110 4.190 ;
        RECT 4.920 3.640 5.110 3.900 ;
        RECT 4.920 3.150 5.390 3.640 ;
        RECT 4.920 2.900 5.110 3.150 ;
        RECT 4.920 2.410 5.390 2.900 ;
        RECT 4.920 2.150 5.110 2.410 ;
        RECT 4.880 1.860 5.110 2.150 ;
        RECT 4.920 1.260 5.110 1.860 ;
        RECT 4.880 0.970 5.110 1.260 ;
        RECT 4.920 0.710 5.110 0.970 ;
        RECT 4.920 0.220 5.390 0.710 ;
        RECT 4.920 0.000 5.110 0.220 ;
    END
  END VGND
  PIN SELECT4
    ANTENNAGATEAREA 0.625000 ;
    PORT
      LAYER met2 ;
        RECT 5.240 1.090 5.580 1.160 ;
        RECT 5.240 0.860 5.720 1.090 ;
    END
  END SELECT4
  PIN SELECT3
    ANTENNAGATEAREA 0.625000 ;
    PORT
      LAYER met2 ;
        RECT 5.240 2.030 5.720 2.260 ;
        RECT 5.240 1.960 5.580 2.030 ;
    END
  END SELECT3
  PIN SELECT2
    ANTENNAGATEAREA 0.625000 ;
    PORT
      LAYER met2 ;
        RECT 5.240 4.020 5.580 4.090 ;
        RECT 5.240 3.790 5.720 4.020 ;
    END
  END SELECT2
  PIN SELECT1
    ANTENNAGATEAREA 0.625000 ;
    PORT
      LAYER met2 ;
        RECT 5.240 4.960 5.720 5.190 ;
        RECT 5.240 4.890 5.580 4.960 ;
    END
  END SELECT1
  OBS
      LAYER li1 ;
        RECT 0.220 4.920 0.390 5.770 ;
        RECT 0.620 4.790 0.790 5.720 ;
        RECT 4.310 5.650 4.550 5.680 ;
        RECT 1.320 5.480 2.280 5.650 ;
        RECT 2.730 5.480 4.070 5.650 ;
        RECT 4.310 5.480 4.880 5.650 ;
        RECT 1.600 5.470 1.770 5.480 ;
        RECT 4.310 5.440 4.550 5.480 ;
        RECT 5.190 5.350 5.360 5.770 ;
        RECT 1.760 5.030 2.090 5.210 ;
        RECT 5.260 5.130 5.430 5.170 ;
        RECT 4.900 5.030 5.090 5.050 ;
        RECT 1.320 4.860 4.070 5.030 ;
        RECT 4.530 4.860 5.090 5.030 ;
        RECT 4.900 4.820 5.090 4.860 ;
        RECT 5.260 4.960 5.490 5.130 ;
        RECT 5.260 4.610 5.430 4.960 ;
        RECT 0.220 3.210 0.390 4.060 ;
        RECT 0.620 3.260 0.790 4.190 ;
        RECT 4.900 4.120 5.090 4.160 ;
        RECT 1.320 3.950 4.070 4.120 ;
        RECT 4.530 3.950 5.090 4.120 ;
        RECT 1.760 3.770 2.090 3.950 ;
        RECT 4.900 3.930 5.090 3.950 ;
        RECT 5.260 4.020 5.430 4.370 ;
        RECT 5.260 3.850 5.490 4.020 ;
        RECT 5.260 3.810 5.430 3.850 ;
        RECT 1.600 3.500 1.770 3.510 ;
        RECT 4.310 3.500 4.550 3.540 ;
        RECT 1.320 3.330 2.280 3.500 ;
        RECT 2.730 3.330 4.070 3.500 ;
        RECT 4.310 3.330 4.880 3.500 ;
        RECT 4.310 3.300 4.550 3.330 ;
        RECT 5.190 3.210 5.360 3.630 ;
        RECT 0.220 1.990 0.390 2.840 ;
        RECT 0.620 1.860 0.790 2.790 ;
        RECT 4.310 2.720 4.550 2.750 ;
        RECT 1.320 2.550 2.280 2.720 ;
        RECT 2.730 2.550 4.070 2.720 ;
        RECT 4.310 2.550 4.880 2.720 ;
        RECT 1.600 2.540 1.770 2.550 ;
        RECT 4.310 2.510 4.550 2.550 ;
        RECT 5.190 2.420 5.360 2.840 ;
        RECT 1.760 2.100 2.090 2.280 ;
        RECT 5.260 2.200 5.430 2.240 ;
        RECT 4.900 2.100 5.090 2.120 ;
        RECT 1.320 1.930 4.070 2.100 ;
        RECT 4.530 1.930 5.090 2.100 ;
        RECT 4.900 1.890 5.090 1.930 ;
        RECT 5.260 2.030 5.490 2.200 ;
        RECT 5.260 1.680 5.430 2.030 ;
        RECT 0.220 0.280 0.390 1.130 ;
        RECT 0.620 0.330 0.790 1.260 ;
        RECT 4.900 1.190 5.090 1.230 ;
        RECT 1.320 1.020 4.070 1.190 ;
        RECT 4.530 1.020 5.090 1.190 ;
        RECT 1.760 0.840 2.090 1.020 ;
        RECT 4.900 1.000 5.090 1.020 ;
        RECT 5.260 1.090 5.430 1.440 ;
        RECT 5.260 0.920 5.490 1.090 ;
        RECT 5.260 0.880 5.430 0.920 ;
        RECT 1.600 0.570 1.770 0.580 ;
        RECT 4.310 0.570 4.550 0.610 ;
        RECT 1.320 0.400 2.280 0.570 ;
        RECT 2.730 0.400 4.070 0.570 ;
        RECT 4.310 0.400 4.880 0.570 ;
        RECT 4.310 0.370 4.550 0.400 ;
        RECT 5.190 0.280 5.360 0.700 ;
      LAYER mcon ;
        RECT 0.220 5.600 0.390 5.770 ;
        RECT 0.220 5.260 0.390 5.430 ;
        RECT 3.600 5.480 3.770 5.650 ;
        RECT 4.350 5.480 4.520 5.650 ;
        RECT 5.190 5.600 5.360 5.770 ;
        RECT 0.620 5.150 0.790 5.320 ;
        RECT 4.910 4.850 5.080 5.020 ;
        RECT 5.320 4.960 5.490 5.130 ;
        RECT 0.220 3.890 0.390 4.060 ;
        RECT 0.220 3.550 0.390 3.720 ;
        RECT 4.910 3.960 5.080 4.130 ;
        RECT 0.620 3.660 0.790 3.830 ;
        RECT 5.320 3.850 5.490 4.020 ;
        RECT 1.600 3.340 1.770 3.510 ;
        RECT 3.600 3.330 3.770 3.500 ;
        RECT 4.350 3.330 4.520 3.500 ;
        RECT 0.220 2.670 0.390 2.840 ;
        RECT 0.220 2.330 0.390 2.500 ;
        RECT 3.600 2.550 3.770 2.720 ;
        RECT 4.350 2.550 4.520 2.720 ;
        RECT 5.190 2.670 5.360 2.840 ;
        RECT 0.620 2.220 0.790 2.390 ;
        RECT 4.910 1.920 5.080 2.090 ;
        RECT 5.320 2.030 5.490 2.200 ;
        RECT 0.220 0.960 0.390 1.130 ;
        RECT 0.220 0.620 0.390 0.790 ;
        RECT 4.910 1.030 5.080 1.200 ;
        RECT 0.620 0.730 0.790 0.900 ;
        RECT 5.320 0.920 5.490 1.090 ;
        RECT 1.600 0.410 1.770 0.580 ;
        RECT 3.600 0.400 3.770 0.570 ;
        RECT 4.350 0.400 4.520 0.570 ;
      LAYER met1 ;
        RECT 1.730 5.670 2.070 5.720 ;
        RECT 1.510 5.650 2.070 5.670 ;
        RECT 4.160 5.690 4.530 5.710 ;
        RECT 1.510 5.480 2.190 5.650 ;
        RECT 1.510 5.440 2.070 5.480 ;
        RECT 1.730 5.400 2.070 5.440 ;
        RECT 4.160 5.430 4.580 5.690 ;
        RECT 4.160 5.420 4.530 5.430 ;
        RECT 5.250 4.900 5.570 5.180 ;
        RECT 5.250 3.800 5.570 4.080 ;
        RECT 1.730 3.540 2.070 3.580 ;
        RECT 1.510 3.500 2.070 3.540 ;
        RECT 4.160 3.550 4.530 3.560 ;
        RECT 1.510 3.330 2.190 3.500 ;
        RECT 1.510 3.310 2.070 3.330 ;
        RECT 1.730 3.260 2.070 3.310 ;
        RECT 4.160 3.290 4.580 3.550 ;
        RECT 4.160 3.270 4.530 3.290 ;
        RECT 1.730 2.740 2.070 2.790 ;
        RECT 1.510 2.720 2.070 2.740 ;
        RECT 4.160 2.760 4.530 2.780 ;
        RECT 1.510 2.550 2.190 2.720 ;
        RECT 1.510 2.510 2.070 2.550 ;
        RECT 1.730 2.470 2.070 2.510 ;
        RECT 4.160 2.500 4.580 2.760 ;
        RECT 4.160 2.490 4.530 2.500 ;
        RECT 5.250 1.970 5.570 2.250 ;
        RECT 5.250 0.870 5.570 1.150 ;
        RECT 1.730 0.610 2.070 0.650 ;
        RECT 1.510 0.570 2.070 0.610 ;
        RECT 4.160 0.620 4.530 0.630 ;
        RECT 1.510 0.400 2.190 0.570 ;
        RECT 1.510 0.380 2.070 0.400 ;
        RECT 1.730 0.330 2.070 0.380 ;
        RECT 4.160 0.360 4.580 0.620 ;
        RECT 4.160 0.340 4.530 0.360 ;
      LAYER via ;
        RECT 1.780 5.430 2.040 5.690 ;
        RECT 4.190 5.430 4.450 5.690 ;
        RECT 5.280 4.910 5.540 5.170 ;
        RECT 5.280 3.810 5.540 4.070 ;
        RECT 1.780 3.290 2.040 3.550 ;
        RECT 4.190 3.290 4.450 3.550 ;
        RECT 1.780 2.500 2.040 2.760 ;
        RECT 4.190 2.500 4.450 2.760 ;
        RECT 5.280 1.980 5.540 2.240 ;
        RECT 5.280 0.880 5.540 1.140 ;
        RECT 1.780 0.360 2.040 0.620 ;
        RECT 4.190 0.360 4.450 0.620 ;
  END
END sky130_hilas_drainSelect01

MACRO sky130_hilas_DAC5bit01
  CLASS CORE ;
  FOREIGN sky130_hilas_DAC5bit01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.580 BY 5.970 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    USE ANALOG ;
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER met2 ;
        RECT 8.260 0.990 8.580 1.020 ;
        RECT 0.000 0.790 8.580 0.990 ;
        RECT 8.260 0.760 8.580 0.790 ;
    END
  END A0
  PIN A1
    USE ANALOG ;
    ANTENNAGATEAREA 0.456300 ;
    PORT
      LAYER met2 ;
        RECT 11.590 5.630 11.910 5.950 ;
        RECT 11.710 2.110 11.860 5.630 ;
        RECT 0.000 1.910 11.870 2.110 ;
        RECT 0.000 1.900 0.140 1.910 ;
    END
  END A1
  PIN A2
    USE ANALOG ;
    ANTENNAGATEAREA 0.608400 ;
    PORT
      LAYER met2 ;
        RECT 9.980 5.650 10.300 5.950 ;
        RECT 9.980 5.630 10.310 5.650 ;
        RECT 10.110 3.090 10.310 5.630 ;
        RECT 0.000 2.880 10.310 3.090 ;
    END
  END A2
  PIN A3
    USE ANALOG ;
    ANTENNAGATEAREA 2.281500 ;
    PORT
      LAYER met2 ;
        RECT 8.370 5.620 8.690 5.940 ;
        RECT 3.540 5.420 3.860 5.570 ;
        RECT 3.480 5.250 3.860 5.420 ;
        RECT 0.000 4.960 2.060 5.020 ;
        RECT 3.480 4.960 3.700 5.250 ;
        RECT 8.400 4.970 8.650 5.620 ;
        RECT 8.400 4.960 8.680 4.970 ;
        RECT 0.000 4.810 8.680 4.960 ;
        RECT 0.260 4.630 0.460 4.810 ;
        RECT 1.900 4.660 8.680 4.810 ;
        RECT 0.210 4.310 0.530 4.630 ;
    END
  END A3
  PIN A4
    USE ANALOG ;
    ANTENNAGATEAREA 3.650400 ;
    PORT
      LAYER met2 ;
        RECT 0.000 5.940 7.050 5.970 ;
        RECT 0.000 5.780 7.070 5.940 ;
        RECT 0.000 5.760 0.150 5.780 ;
        RECT 0.350 5.620 0.670 5.780 ;
        RECT 1.940 5.630 2.260 5.780 ;
        RECT 5.140 5.620 5.460 5.780 ;
        RECT 6.750 5.620 7.070 5.780 ;
    END
  END A4
  PIN VPWR
    USE ANALOG ;
    ANTENNADIFFAREA 3.264300 ;
    PORT
      LAYER met2 ;
        RECT 12.710 5.690 13.870 5.970 ;
        RECT 12.830 5.510 13.140 5.690 ;
        RECT 13.460 5.680 13.870 5.690 ;
        RECT 13.500 5.510 13.810 5.680 ;
    END
  END VPWR
  PIN OUT
    USE ANALOG ;
    ANTENNADIFFAREA 3.264300 ;
    PORT
      LAYER met1 ;
        RECT 3.010 0.240 3.240 0.290 ;
        RECT 4.630 0.240 4.860 0.290 ;
        RECT 6.230 0.240 6.460 0.290 ;
        RECT 7.850 0.240 8.080 0.290 ;
        RECT 9.450 0.240 9.680 0.290 ;
        RECT 11.070 0.240 11.300 0.290 ;
        RECT 12.670 0.240 12.900 0.290 ;
        RECT 14.280 0.240 14.510 0.290 ;
        RECT 3.010 0.010 16.580 0.240 ;
        RECT 3.010 0.000 3.240 0.010 ;
        RECT 4.630 0.000 4.860 0.010 ;
        RECT 6.230 0.000 6.460 0.010 ;
        RECT 7.850 0.000 8.080 0.010 ;
        RECT 9.450 0.000 9.680 0.010 ;
        RECT 11.070 0.000 11.300 0.010 ;
        RECT 12.670 0.000 12.900 0.010 ;
        RECT 14.280 0.000 14.510 0.010 ;
    END
  END OUT
  OBS
      LAYER nwell ;
        RECT 0.370 0.030 16.470 5.680 ;
      LAYER li1 ;
        RECT 0.400 5.470 0.610 5.900 ;
        RECT 1.990 5.480 2.200 5.910 ;
        RECT 3.390 5.500 3.820 5.520 ;
        RECT 0.420 5.450 0.590 5.470 ;
        RECT 2.010 5.460 2.180 5.480 ;
        RECT 3.370 5.330 3.820 5.500 ;
        RECT 5.190 5.470 5.400 5.900 ;
        RECT 6.800 5.470 7.010 5.900 ;
        RECT 8.420 5.470 8.630 5.900 ;
        RECT 10.030 5.480 10.240 5.910 ;
        RECT 11.640 5.480 11.850 5.910 ;
        RECT 12.950 5.800 13.160 5.810 ;
        RECT 12.840 5.760 13.160 5.800 ;
        RECT 13.510 5.760 13.830 5.800 ;
        RECT 12.840 5.570 13.170 5.760 ;
        RECT 13.510 5.570 13.840 5.760 ;
        RECT 12.840 5.540 13.160 5.570 ;
        RECT 13.510 5.540 13.830 5.570 ;
        RECT 5.210 5.450 5.380 5.470 ;
        RECT 6.820 5.450 6.990 5.470 ;
        RECT 8.440 5.450 8.610 5.470 ;
        RECT 10.050 5.460 10.220 5.480 ;
        RECT 11.660 5.460 11.830 5.480 ;
        RECT 3.390 5.310 3.820 5.330 ;
        RECT 3.980 5.030 4.150 5.040 ;
        RECT 12.950 5.030 13.160 5.540 ;
        RECT 13.620 5.030 13.790 5.540 ;
        RECT 2.370 4.800 13.800 5.030 ;
        RECT 0.260 4.160 0.470 4.590 ;
        RECT 2.370 4.460 2.540 4.800 ;
        RECT 0.280 4.140 0.450 4.160 ;
        RECT 2.360 4.130 2.540 4.460 ;
        RECT 0.320 3.210 0.530 3.640 ;
        RECT 2.370 3.500 2.540 4.130 ;
        RECT 0.340 3.190 0.510 3.210 ;
        RECT 2.360 3.170 2.540 3.500 ;
        RECT 0.320 2.270 0.530 2.700 ;
        RECT 2.370 2.540 2.540 3.170 ;
        RECT 0.340 2.250 0.510 2.270 ;
        RECT 2.360 2.210 2.540 2.540 ;
        RECT 2.370 1.580 2.540 2.210 ;
        RECT 2.360 1.250 2.540 1.580 ;
        RECT 2.370 1.240 2.540 1.250 ;
        RECT 3.030 4.460 3.200 4.470 ;
        RECT 3.980 4.460 4.150 4.800 ;
        RECT 5.570 4.460 5.740 4.800 ;
        RECT 3.030 4.130 3.210 4.460 ;
        RECT 3.970 4.130 4.150 4.460 ;
        RECT 4.650 4.430 4.820 4.460 ;
        RECT 4.650 4.130 4.830 4.430 ;
        RECT 3.030 3.500 3.200 4.130 ;
        RECT 3.980 3.500 4.150 4.130 ;
        RECT 4.660 3.500 4.830 4.130 ;
        RECT 3.030 3.170 3.210 3.500 ;
        RECT 3.970 3.170 4.150 3.500 ;
        RECT 4.650 3.170 4.830 3.500 ;
        RECT 3.030 2.540 3.200 3.170 ;
        RECT 3.980 2.540 4.150 3.170 ;
        RECT 4.660 2.540 4.830 3.170 ;
        RECT 3.030 2.210 3.210 2.540 ;
        RECT 3.970 2.210 4.150 2.540 ;
        RECT 4.650 2.210 4.830 2.540 ;
        RECT 3.030 1.580 3.200 2.210 ;
        RECT 3.980 1.580 4.150 2.210 ;
        RECT 4.660 1.580 4.830 2.210 ;
        RECT 3.030 1.250 3.210 1.580 ;
        RECT 3.970 1.250 4.150 1.580 ;
        RECT 4.650 1.250 4.830 1.580 ;
        RECT 3.030 0.260 3.200 1.250 ;
        RECT 3.980 1.240 4.150 1.250 ;
        RECT 4.660 0.260 4.830 1.250 ;
        RECT 5.570 4.130 5.750 4.460 ;
        RECT 5.570 3.500 5.740 4.130 ;
        RECT 5.570 3.170 5.750 3.500 ;
        RECT 5.570 2.540 5.740 3.170 ;
        RECT 5.570 2.210 5.750 2.540 ;
        RECT 5.570 1.580 5.740 2.210 ;
        RECT 5.570 1.250 5.750 1.580 ;
        RECT 5.570 1.240 5.740 1.250 ;
        RECT 6.260 0.260 6.430 4.510 ;
        RECT 6.740 3.220 6.950 3.650 ;
        RECT 6.760 3.200 6.930 3.220 ;
        RECT 7.190 1.240 7.360 4.800 ;
        RECT 8.810 4.460 8.980 4.800 ;
        RECT 7.870 4.130 8.050 4.460 ;
        RECT 8.800 4.130 8.980 4.460 ;
        RECT 7.880 3.500 8.050 4.130 ;
        RECT 8.810 3.500 8.980 4.130 ;
        RECT 7.870 3.170 8.050 3.500 ;
        RECT 8.800 3.170 8.980 3.500 ;
        RECT 7.880 2.540 8.050 3.170 ;
        RECT 8.270 2.740 8.440 2.760 ;
        RECT 7.870 2.210 8.050 2.540 ;
        RECT 8.250 2.310 8.460 2.740 ;
        RECT 7.880 1.580 8.050 2.210 ;
        RECT 8.810 1.580 8.980 3.170 ;
        RECT 7.870 1.250 8.050 1.580 ;
        RECT 8.800 1.260 8.980 1.580 ;
        RECT 8.800 1.250 8.970 1.260 ;
        RECT 7.880 0.260 8.050 1.250 ;
        RECT 9.480 0.260 9.650 4.510 ;
        RECT 9.990 1.310 10.200 1.740 ;
        RECT 10.010 1.290 10.180 1.310 ;
        RECT 10.410 1.250 10.580 4.800 ;
        RECT 11.100 4.460 11.270 4.510 ;
        RECT 11.090 4.130 11.270 4.460 ;
        RECT 11.100 3.500 11.270 4.130 ;
        RECT 11.090 3.170 11.270 3.500 ;
        RECT 11.100 2.540 11.270 3.170 ;
        RECT 11.090 2.210 11.270 2.540 ;
        RECT 11.100 1.580 11.270 2.210 ;
        RECT 11.090 1.250 11.270 1.580 ;
        RECT 12.020 1.250 12.190 4.800 ;
        RECT 11.100 0.260 11.270 1.250 ;
        RECT 12.700 0.260 12.870 4.490 ;
        RECT 13.630 1.230 13.800 4.800 ;
        RECT 14.310 0.260 14.480 4.670 ;
        RECT 3.030 0.030 3.220 0.260 ;
        RECT 4.650 0.030 4.840 0.260 ;
        RECT 6.250 0.030 6.440 0.260 ;
        RECT 7.870 0.030 8.060 0.260 ;
        RECT 9.470 0.030 9.660 0.260 ;
        RECT 11.090 0.030 11.280 0.260 ;
        RECT 12.690 0.030 12.880 0.260 ;
        RECT 14.300 0.030 14.490 0.260 ;
        RECT 3.030 0.010 3.200 0.030 ;
        RECT 4.660 0.010 4.830 0.030 ;
        RECT 6.260 0.010 6.430 0.030 ;
        RECT 7.880 0.010 8.050 0.030 ;
        RECT 9.480 0.010 9.650 0.030 ;
        RECT 11.100 0.010 11.270 0.030 ;
        RECT 12.700 0.010 12.870 0.030 ;
        RECT 14.310 0.010 14.480 0.030 ;
      LAYER mcon ;
        RECT 12.900 5.580 13.070 5.750 ;
        RECT 13.570 5.580 13.740 5.750 ;
        RECT 8.270 2.590 8.440 2.760 ;
        RECT 3.040 0.060 3.210 0.230 ;
        RECT 4.660 0.060 4.830 0.230 ;
        RECT 6.260 0.060 6.430 0.230 ;
        RECT 7.880 0.060 8.050 0.230 ;
        RECT 9.480 0.060 9.650 0.230 ;
        RECT 11.100 0.060 11.270 0.230 ;
        RECT 12.700 0.060 12.870 0.230 ;
        RECT 14.310 0.060 14.480 0.230 ;
      LAYER met1 ;
        RECT 0.350 5.620 0.670 5.940 ;
        RECT 1.940 5.630 2.260 5.950 ;
        RECT 0.390 5.390 0.620 5.620 ;
        RECT 1.980 5.400 2.210 5.630 ;
        RECT 5.140 5.620 5.460 5.940 ;
        RECT 6.750 5.620 7.070 5.940 ;
        RECT 8.370 5.620 8.690 5.940 ;
        RECT 9.980 5.630 10.300 5.950 ;
        RECT 11.590 5.630 11.910 5.950 ;
        RECT 3.540 5.530 3.860 5.570 ;
        RECT 3.310 5.300 3.860 5.530 ;
        RECT 5.180 5.390 5.410 5.620 ;
        RECT 6.790 5.390 7.020 5.620 ;
        RECT 8.410 5.390 8.640 5.620 ;
        RECT 10.020 5.400 10.250 5.630 ;
        RECT 11.630 5.400 11.860 5.630 ;
        RECT 12.830 5.510 13.150 5.830 ;
        RECT 13.500 5.510 13.820 5.830 ;
        RECT 3.540 5.250 3.860 5.300 ;
        RECT 0.210 4.310 0.530 4.630 ;
        RECT 0.250 4.080 0.480 4.310 ;
        RECT 0.270 3.360 0.590 3.680 ;
        RECT 6.740 3.560 10.190 3.730 ;
        RECT 6.740 3.430 6.960 3.560 ;
        RECT 0.310 3.130 0.540 3.360 ;
        RECT 6.730 3.140 6.960 3.430 ;
        RECT 0.270 2.420 0.590 2.740 ;
        RECT 8.240 2.530 8.470 2.820 ;
        RECT 0.310 2.190 0.540 2.420 ;
        RECT 8.250 2.310 8.470 2.530 ;
        RECT 8.290 1.050 8.470 2.310 ;
        RECT 9.990 1.740 10.190 3.560 ;
        RECT 9.990 1.520 10.210 1.740 ;
        RECT 9.980 1.230 10.210 1.520 ;
        RECT 8.290 0.730 8.550 1.050 ;
      LAYER via ;
        RECT 0.380 5.650 0.640 5.910 ;
        RECT 1.970 5.660 2.230 5.920 ;
        RECT 5.170 5.650 5.430 5.910 ;
        RECT 6.780 5.650 7.040 5.910 ;
        RECT 8.400 5.650 8.660 5.910 ;
        RECT 10.010 5.660 10.270 5.920 ;
        RECT 11.620 5.660 11.880 5.920 ;
        RECT 3.570 5.280 3.830 5.540 ;
        RECT 12.860 5.540 13.120 5.800 ;
        RECT 13.530 5.540 13.790 5.800 ;
        RECT 0.240 4.340 0.500 4.600 ;
        RECT 0.300 3.390 0.560 3.650 ;
        RECT 0.300 2.450 0.560 2.710 ;
        RECT 8.290 0.760 8.550 1.020 ;
      LAYER met2 ;
        RECT 0.270 3.360 0.590 3.680 ;
        RECT 0.270 2.420 0.590 2.740 ;
  END
END sky130_hilas_DAC5bit01

MACRO sky130_hilas_capacitorSize04
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize04 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.780 BY 5.290 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAP1TERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 4.960 3.830 5.620 4.490 ;
    END
  END CAP1TERM02
  PIN CAP2TERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 4.960 0.830 5.620 1.490 ;
    END
  END CAP2TERM02
  PIN CAP2TERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 0.120 1.230 0.780 1.490 ;
        RECT 2.560 1.230 3.010 1.240 ;
        RECT 0.120 0.830 3.060 1.230 ;
        RECT 0.570 0.820 3.060 0.830 ;
        RECT 2.540 0.740 3.060 0.820 ;
    END
  END CAP2TERM01
  PIN CAP1TERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 0.090 4.240 0.750 4.490 ;
        RECT 2.560 4.240 3.010 4.250 ;
        RECT 0.090 3.830 3.060 4.240 ;
        RECT 2.540 3.750 3.060 3.830 ;
    END
  END CAP1TERM01
  OBS
      LAYER met2 ;
        RECT 0.020 4.980 5.770 5.160 ;
        RECT 0.020 4.550 5.770 4.730 ;
        RECT 0.220 4.310 0.590 4.370 ;
        RECT 0.020 4.030 0.590 4.310 ;
        RECT 0.220 3.970 0.590 4.030 ;
        RECT 5.090 4.310 5.460 4.370 ;
        RECT 5.090 4.030 5.770 4.310 ;
        RECT 5.090 3.970 5.460 4.030 ;
        RECT 0.020 3.550 5.770 3.730 ;
        RECT 0.020 3.120 5.770 3.300 ;
        RECT 0.020 1.970 5.770 2.140 ;
        RECT 0.020 1.550 5.770 1.720 ;
        RECT 0.250 1.310 0.620 1.370 ;
        RECT 0.020 1.030 0.620 1.310 ;
        RECT 0.250 0.970 0.620 1.030 ;
        RECT 5.090 1.310 5.460 1.370 ;
        RECT 5.090 1.030 5.780 1.310 ;
        RECT 5.090 0.970 5.460 1.030 ;
        RECT 0.020 0.570 5.770 0.740 ;
        RECT 0.020 0.130 5.770 0.300 ;
      LAYER via2 ;
        RECT 0.270 4.030 0.550 4.310 ;
        RECT 5.140 4.030 5.420 4.310 ;
        RECT 0.300 1.030 0.580 1.310 ;
        RECT 5.140 1.030 5.420 1.310 ;
      LAYER met3 ;
        RECT 1.710 4.520 4.010 5.290 ;
        RECT 0.000 3.770 0.790 4.520 ;
        RECT 1.710 3.770 5.660 4.520 ;
        RECT 1.710 3.010 4.010 3.770 ;
        RECT 0.030 0.770 0.820 1.520 ;
        RECT 1.710 1.510 4.010 2.280 ;
        RECT 4.870 1.510 5.660 1.520 ;
        RECT 1.710 0.780 5.660 1.510 ;
        RECT 1.710 0.000 4.010 0.780 ;
        RECT 4.870 0.770 5.660 0.780 ;
      LAYER via3 ;
        RECT 0.190 3.920 0.620 4.400 ;
        RECT 5.060 3.920 5.490 4.400 ;
        RECT 0.220 0.920 0.650 1.400 ;
        RECT 5.060 0.920 5.490 1.400 ;
  END
END sky130_hilas_capacitorSize04

MACRO sky130_hilas_capacitorArray01
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorArray01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.700 BY 9.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM2
    USE ANALOG ;
    PORT
      LAYER met3 ;
        RECT 35.230 2.200 36.380 3.840 ;
        RECT 35.680 2.190 36.380 2.200 ;
    END
  END CAPTERM2
  PIN CAPTERM1
    USE ANALOG ;
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met3 ;
        RECT 11.250 5.740 11.630 6.030 ;
        RECT 11.170 4.490 11.710 5.740 ;
    END
  END CAPTERM1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 5.400 5.380 5.720 5.390 ;
        RECT 8.980 5.380 36.700 5.550 ;
        RECT 5.400 5.370 36.700 5.380 ;
        RECT 5.400 5.200 9.650 5.370 ;
        RECT 5.400 5.130 5.720 5.200 ;
        RECT 9.330 5.140 9.650 5.200 ;
    END
  END VINJ
  PIN GATESELECT
    PORT
      LAYER met1 ;
        RECT 9.120 6.000 9.310 6.050 ;
    END
  END GATESELECT
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 0.360 5.910 0.760 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.360 0.000 0.750 0.120 ;
    END
  END VTUN
  PIN GATE
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 4.420 5.970 4.790 6.050 ;
        RECT 4.410 5.920 4.790 5.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.400 0.130 4.410 0.150 ;
        RECT 4.400 0.010 4.790 0.130 ;
        RECT 4.400 0.000 4.410 0.010 ;
    END
  END GATE
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 0.000 3.510 0.120 3.690 ;
    END
    PORT
      LAYER met2 ;
        RECT 35.690 3.690 36.700 3.700 ;
        RECT 8.940 3.510 36.700 3.690 ;
    END
  END DRAIN2
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 0.010 5.370 0.120 5.550 ;
    END
  END DRAIN1
  PIN DRAIN4
    PORT
      LAYER met2 ;
        RECT 8.810 0.520 36.700 0.690 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.020 0.520 0.120 0.690 ;
    END
  END DRAIN4
  PIN DRAIN3
    PORT
      LAYER met2 ;
        RECT 8.770 2.360 36.700 2.530 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.020 2.360 0.120 2.530 ;
    END
  END DRAIN3
  PIN VGND
    ANTENNADIFFAREA 1.978000 ;
    PORT
      LAYER nwell ;
        RECT 2.650 8.010 4.380 9.870 ;
        RECT 2.640 6.170 4.380 8.010 ;
        RECT 2.650 3.820 4.380 6.170 ;
      LAYER met1 ;
        RECT 3.000 6.050 3.400 9.870 ;
        RECT 2.800 5.990 3.400 6.050 ;
        RECT 3.000 3.820 3.400 5.990 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.730 5.980 6.970 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.800 0.000 3.040 0.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.730 0.000 6.970 0.070 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 0.010 5.370 0.120 5.550 ;
        RECT 6.400 3.820 8.630 9.870 ;
        RECT 10.160 9.860 12.710 9.870 ;
        RECT 10.160 6.050 12.720 9.860 ;
        RECT 10.070 6.040 35.420 6.050 ;
        RECT 10.080 5.970 35.420 6.040 ;
        RECT 0.000 3.510 0.120 3.690 ;
        RECT 0.020 0.520 0.120 0.690 ;
        RECT 10.060 0.060 35.420 5.970 ;
        RECT 10.070 0.010 35.420 0.060 ;
        RECT 12.000 0.000 35.420 0.010 ;
      LAYER li1 ;
        RECT 10.260 9.460 10.580 9.470 ;
        RECT 10.260 9.290 10.840 9.460 ;
        RECT 10.260 9.240 10.590 9.290 ;
        RECT 10.260 9.210 10.580 9.240 ;
        RECT 12.120 9.190 12.320 9.540 ;
        RECT 10.260 8.880 10.580 8.920 ;
        RECT 10.260 8.840 10.590 8.880 ;
        RECT 10.260 8.670 10.840 8.840 ;
        RECT 10.260 8.660 10.580 8.670 ;
        RECT 5.470 8.120 5.640 8.630 ;
        RECT 9.410 8.110 9.580 8.620 ;
        RECT 11.390 8.600 11.590 9.170 ;
        RECT 12.120 9.160 12.330 9.190 ;
        RECT 12.110 8.570 12.330 9.160 ;
        RECT 10.260 8.030 10.580 8.040 ;
        RECT 10.260 7.860 10.840 8.030 ;
        RECT 10.260 7.820 10.590 7.860 ;
        RECT 10.260 7.780 10.580 7.820 ;
        RECT 11.390 7.530 11.590 8.100 ;
        RECT 12.110 7.540 12.330 8.130 ;
        RECT 12.120 7.510 12.330 7.540 ;
        RECT 10.260 7.460 10.580 7.490 ;
        RECT 3.070 6.620 3.620 7.050 ;
        RECT 5.480 6.410 5.650 7.420 ;
        RECT 10.260 7.410 10.590 7.460 ;
        RECT 7.100 6.550 7.650 6.980 ;
        RECT 9.410 6.270 9.580 7.280 ;
        RECT 10.260 7.240 10.840 7.410 ;
        RECT 10.260 7.230 10.580 7.240 ;
        RECT 12.120 7.160 12.320 7.510 ;
        RECT 11.510 6.760 11.950 6.930 ;
        RECT 10.260 6.450 10.580 6.460 ;
        RECT 10.260 6.280 10.840 6.450 ;
        RECT 10.260 6.230 10.590 6.280 ;
        RECT 10.260 6.200 10.580 6.230 ;
        RECT 12.120 6.180 12.320 6.530 ;
        RECT 10.260 5.870 10.580 5.910 ;
        RECT 10.260 5.830 10.590 5.870 ;
        RECT 10.260 5.660 10.840 5.830 ;
        RECT 10.260 5.650 10.580 5.660 ;
        RECT 11.390 5.590 11.590 6.160 ;
        RECT 12.120 6.150 12.330 6.180 ;
        RECT 12.110 5.560 12.330 6.150 ;
        RECT 10.260 5.030 10.580 5.040 ;
        RECT 10.260 4.860 10.840 5.030 ;
        RECT 10.260 4.820 10.590 4.860 ;
        RECT 10.260 4.780 10.580 4.820 ;
        RECT 11.390 4.530 11.590 5.100 ;
        RECT 12.110 4.540 12.330 5.130 ;
        RECT 12.120 4.510 12.330 4.540 ;
        RECT 10.260 4.460 10.580 4.490 ;
        RECT 10.260 4.410 10.590 4.460 ;
        RECT 10.260 4.240 10.840 4.410 ;
        RECT 10.260 4.230 10.580 4.240 ;
        RECT 12.120 4.160 12.320 4.510 ;
      LAYER mcon ;
        RECT 10.320 9.250 10.490 9.420 ;
        RECT 11.400 8.960 11.570 9.130 ;
        RECT 10.320 8.700 10.490 8.870 ;
        RECT 5.470 8.460 5.640 8.630 ;
        RECT 9.410 8.450 9.580 8.620 ;
        RECT 12.130 8.990 12.300 9.160 ;
        RECT 10.320 7.830 10.490 8.000 ;
        RECT 11.400 7.570 11.570 7.740 ;
        RECT 12.130 7.540 12.300 7.710 ;
        RECT 10.320 7.280 10.490 7.450 ;
        RECT 3.070 6.700 3.340 6.970 ;
        RECT 5.480 7.000 5.650 7.170 ;
        RECT 5.480 6.660 5.650 6.830 ;
        RECT 7.100 6.630 7.370 6.900 ;
        RECT 9.410 6.860 9.580 7.030 ;
        RECT 11.770 6.760 11.950 6.930 ;
        RECT 9.410 6.520 9.580 6.690 ;
        RECT 10.320 6.240 10.490 6.410 ;
        RECT 11.400 5.950 11.570 6.120 ;
        RECT 10.320 5.690 10.490 5.860 ;
        RECT 12.130 5.980 12.300 6.150 ;
        RECT 10.320 4.830 10.490 5.000 ;
        RECT 11.400 4.570 11.570 4.740 ;
        RECT 12.130 4.540 12.300 4.710 ;
        RECT 10.320 4.280 10.490 4.450 ;
      LAYER met1 ;
        RECT 5.440 8.690 5.680 9.870 ;
        RECT 5.430 8.030 5.690 8.690 ;
        RECT 5.440 5.420 5.680 8.030 ;
        RECT 7.050 7.950 7.430 9.870 ;
        RECT 9.370 8.710 9.610 9.870 ;
        RECT 10.250 9.180 10.570 9.500 ;
        RECT 11.390 9.190 11.550 9.870 ;
        RECT 11.390 9.170 11.590 9.190 ;
        RECT 9.350 8.050 9.620 8.710 ;
        RECT 10.250 8.630 10.570 8.950 ;
        RECT 11.370 8.930 11.600 9.170 ;
        RECT 11.390 8.710 11.590 8.930 ;
        RECT 11.760 8.880 11.950 9.870 ;
        RECT 12.200 9.220 12.360 9.870 ;
        RECT 11.780 8.760 11.950 8.880 ;
        RECT 7.040 6.090 7.430 7.950 ;
        RECT 5.430 5.100 5.690 5.420 ;
        RECT 5.440 3.820 5.680 5.100 ;
        RECT 7.050 3.820 7.430 6.090 ;
        RECT 9.370 6.050 9.610 8.050 ;
        RECT 10.250 7.750 10.570 8.070 ;
        RECT 11.390 7.990 11.550 8.710 ;
        RECT 11.390 7.770 11.590 7.990 ;
        RECT 11.790 7.940 11.950 8.760 ;
        RECT 12.090 8.670 12.360 9.220 ;
        RECT 12.090 8.620 12.370 8.670 ;
        RECT 12.200 8.530 12.370 8.620 ;
        RECT 12.200 8.170 12.360 8.530 ;
        RECT 12.200 8.080 12.370 8.170 ;
        RECT 11.780 7.820 11.950 7.940 ;
        RECT 11.370 7.530 11.600 7.770 ;
        RECT 10.250 7.200 10.570 7.520 ;
        RECT 11.390 7.510 11.590 7.530 ;
        RECT 10.250 6.170 10.570 6.490 ;
        RECT 11.390 6.180 11.550 7.510 ;
        RECT 11.760 6.960 11.950 7.820 ;
        RECT 12.090 8.030 12.370 8.080 ;
        RECT 12.090 7.480 12.360 8.030 ;
        RECT 11.740 6.730 11.980 6.960 ;
        RECT 11.390 6.160 11.590 6.180 ;
        RECT 8.700 5.710 8.960 6.030 ;
        RECT 9.370 6.000 9.720 6.050 ;
        RECT 9.370 5.460 9.610 6.000 ;
        RECT 10.250 5.620 10.570 5.940 ;
        RECT 11.370 5.920 11.600 6.160 ;
        RECT 11.390 5.700 11.590 5.920 ;
        RECT 11.760 5.870 11.950 6.730 ;
        RECT 12.200 6.210 12.360 7.480 ;
        RECT 11.780 5.750 11.950 5.870 ;
        RECT 9.360 5.140 9.620 5.460 ;
        RECT 9.370 3.820 9.610 5.140 ;
        RECT 10.250 4.750 10.570 5.070 ;
        RECT 11.390 4.990 11.550 5.700 ;
        RECT 11.390 4.770 11.590 4.990 ;
        RECT 11.790 4.940 11.950 5.750 ;
        RECT 12.090 5.660 12.360 6.210 ;
        RECT 12.090 5.610 12.370 5.660 ;
        RECT 12.200 5.520 12.370 5.610 ;
        RECT 12.200 5.170 12.360 5.520 ;
        RECT 12.200 5.080 12.370 5.170 ;
        RECT 11.780 4.820 11.950 4.940 ;
        RECT 11.370 4.530 11.600 4.770 ;
        RECT 10.250 4.200 10.570 4.520 ;
        RECT 11.390 4.510 11.590 4.530 ;
        RECT 11.390 3.830 11.550 4.510 ;
        RECT 11.760 3.830 11.950 4.820 ;
        RECT 12.090 5.030 12.370 5.080 ;
        RECT 12.090 4.480 12.360 5.030 ;
        RECT 12.200 3.830 12.360 4.480 ;
        RECT 8.750 0.010 8.910 0.070 ;
        RECT 9.120 0.010 9.310 0.070 ;
        RECT 9.560 0.010 9.720 0.070 ;
      LAYER via ;
        RECT 10.280 9.210 10.540 9.470 ;
        RECT 10.280 8.660 10.540 8.920 ;
        RECT 5.430 5.130 5.690 5.390 ;
        RECT 10.280 7.780 10.540 8.040 ;
        RECT 10.280 7.230 10.540 7.490 ;
        RECT 10.280 6.200 10.540 6.460 ;
        RECT 8.700 5.740 8.960 6.000 ;
        RECT 10.280 5.650 10.540 5.910 ;
        RECT 9.360 5.170 9.620 5.430 ;
        RECT 10.280 4.780 10.540 5.040 ;
        RECT 10.280 4.230 10.540 4.490 ;
      LAYER met2 ;
        RECT 10.250 9.370 10.560 9.510 ;
        RECT 2.650 9.190 12.720 9.370 ;
        RECT 10.250 9.180 10.560 9.190 ;
        RECT 10.250 8.940 10.560 8.960 ;
        RECT 2.650 8.760 12.720 8.940 ;
        RECT 10.250 8.630 10.560 8.760 ;
        RECT 10.250 7.940 10.560 8.070 ;
        RECT 2.640 7.760 12.720 7.940 ;
        RECT 10.250 7.740 10.560 7.760 ;
        RECT 10.250 7.510 10.560 7.520 ;
        RECT 2.640 7.330 12.720 7.510 ;
        RECT 10.250 7.190 10.560 7.330 ;
        RECT 10.250 6.360 10.560 6.500 ;
        RECT 10.250 6.350 12.720 6.360 ;
        RECT 2.660 6.180 12.720 6.350 ;
        RECT 10.250 6.170 10.560 6.180 ;
        RECT 10.740 6.020 11.250 6.050 ;
        RECT 8.670 5.930 8.990 6.000 ;
        RECT 10.250 5.930 10.560 5.950 ;
        RECT 10.740 5.930 11.670 6.020 ;
        RECT 2.660 5.760 12.720 5.930 ;
        RECT 8.670 5.750 12.720 5.760 ;
        RECT 8.670 5.740 11.670 5.750 ;
        RECT 10.250 5.620 10.560 5.740 ;
        RECT 11.170 5.720 11.670 5.740 ;
        RECT 8.920 4.950 36.700 5.120 ;
        RECT 2.660 4.940 36.700 4.950 ;
        RECT 2.660 4.780 12.720 4.940 ;
        RECT 3.440 4.690 4.980 4.780 ;
        RECT 10.160 4.760 12.720 4.780 ;
        RECT 10.250 4.740 10.560 4.760 ;
        RECT 10.250 4.510 10.560 4.520 ;
        RECT 2.660 4.340 12.720 4.510 ;
        RECT 10.250 4.330 12.720 4.340 ;
        RECT 10.250 4.290 10.560 4.330 ;
        RECT 9.880 4.190 10.560 4.290 ;
        RECT 9.880 4.120 10.250 4.190 ;
        RECT 8.980 3.940 36.700 4.120 ;
        RECT 9.880 3.890 10.250 3.940 ;
        RECT 36.010 2.790 36.700 3.200 ;
        RECT 9.840 2.110 10.210 2.200 ;
        RECT 8.870 1.940 36.700 2.110 ;
        RECT 9.840 1.800 10.210 1.940 ;
        RECT 10.930 1.130 11.300 1.330 ;
        RECT 8.850 0.960 36.700 1.130 ;
        RECT 10.930 0.930 11.300 0.960 ;
      LAYER via2 ;
        RECT 11.300 5.720 11.580 6.000 ;
        RECT 9.930 3.950 10.210 4.230 ;
        RECT 36.080 2.850 36.370 3.130 ;
        RECT 9.890 1.860 10.170 2.140 ;
        RECT 10.980 0.990 11.260 1.270 ;
      LAYER met3 ;
        RECT 9.660 3.690 10.450 4.440 ;
        RECT 9.620 2.300 10.410 2.350 ;
        RECT 9.620 2.000 10.550 2.300 ;
        RECT 9.620 1.600 10.410 2.000 ;
        RECT 10.710 1.090 11.500 1.480 ;
        RECT 10.710 0.790 11.640 1.090 ;
        RECT 10.710 0.730 11.500 0.790 ;
      LAYER via3 ;
        RECT 9.850 3.840 10.280 4.320 ;
        RECT 9.810 1.750 10.240 2.230 ;
        RECT 10.900 0.880 11.330 1.360 ;
      LAYER met4 ;
        RECT 12.790 5.380 16.890 5.680 ;
        RECT 11.100 4.770 13.800 4.880 ;
        RECT 11.100 4.470 14.010 4.770 ;
        RECT 9.750 4.050 10.410 4.410 ;
        RECT 13.500 4.130 14.010 4.470 ;
        RECT 16.510 4.180 16.890 5.380 ;
        RECT 19.350 4.210 22.630 4.510 ;
        RECT 9.750 3.750 11.770 4.050 ;
        RECT 11.470 3.190 11.770 3.750 ;
        RECT 19.350 3.190 19.650 4.210 ;
        RECT 22.330 3.190 22.630 4.210 ;
        RECT 11.470 2.890 22.630 3.190 ;
        RECT 25.030 4.190 33.920 4.490 ;
        RECT 9.710 2.300 10.370 2.320 ;
        RECT 13.710 2.300 16.900 2.330 ;
        RECT 19.350 2.300 19.650 2.330 ;
        RECT 9.710 2.000 22.570 2.300 ;
        RECT 9.710 1.660 10.370 2.000 ;
        RECT 13.710 1.630 14.010 2.000 ;
        RECT 16.600 1.660 16.900 2.000 ;
        RECT 19.350 1.660 19.650 2.000 ;
        RECT 16.600 1.630 19.650 1.660 ;
        RECT 22.270 1.630 22.570 2.000 ;
        RECT 10.800 1.090 11.460 1.450 ;
        RECT 13.710 1.330 22.570 1.630 ;
        RECT 25.030 1.670 25.330 4.190 ;
        RECT 27.860 4.160 30.970 4.190 ;
        RECT 27.860 1.670 28.160 4.160 ;
        RECT 30.670 1.670 30.970 4.160 ;
        RECT 33.620 1.670 33.920 4.190 ;
        RECT 25.030 1.370 33.980 1.670 ;
        RECT 30.670 1.360 33.980 1.370 ;
        RECT 10.800 0.790 11.850 1.090 ;
        RECT 11.550 0.550 11.850 0.790 ;
        RECT 33.680 0.550 33.980 1.360 ;
        RECT 11.550 0.250 33.980 0.550 ;
  END
END sky130_hilas_capacitorArray01

MACRO sky130_hilas_pFETmed
  CLASS CORE ;
  FOREIGN sky130_hilas_pFETmed ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.190 BY 2.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 0.000 0.000 1.190 2.870 ;
      LAYER li1 ;
        RECT 0.240 0.150 0.410 2.640 ;
        RECT 0.790 0.140 0.960 2.640 ;
  END
END sky130_hilas_pFETmed

MACRO sky130_hilas_swc4x1cellOverlap2
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x1cellOverlap2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.350 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 2.790 6.040 9.340 6.050 ;
        RECT 2.790 0.020 9.350 6.040 ;
        RECT 2.790 0.010 9.340 0.020 ;
        RECT 2.790 0.000 6.790 0.010 ;
      LAYER li1 ;
        RECT 1.060 4.840 1.230 5.730 ;
        RECT 3.140 4.740 6.450 5.720 ;
        RECT 6.890 5.640 7.210 5.650 ;
        RECT 6.890 5.470 7.470 5.640 ;
        RECT 6.890 5.420 7.220 5.470 ;
        RECT 6.890 5.390 7.210 5.420 ;
        RECT 8.750 5.370 8.950 5.720 ;
        RECT 6.890 5.060 7.210 5.100 ;
        RECT 6.890 5.020 7.220 5.060 ;
        RECT 6.890 4.850 7.470 5.020 ;
        RECT 6.890 4.840 7.210 4.850 ;
        RECT 8.020 4.780 8.220 5.350 ;
        RECT 8.750 5.340 8.960 5.370 ;
        RECT 8.740 4.750 8.960 5.340 ;
        RECT 1.060 3.320 1.230 4.210 ;
        RECT 3.140 3.270 6.450 4.250 ;
        RECT 6.890 4.210 7.210 4.220 ;
        RECT 6.890 4.040 7.470 4.210 ;
        RECT 6.890 4.000 7.220 4.040 ;
        RECT 6.890 3.960 7.210 4.000 ;
        RECT 8.020 3.710 8.220 4.280 ;
        RECT 8.740 3.720 8.960 4.310 ;
        RECT 8.750 3.690 8.960 3.720 ;
        RECT 6.890 3.640 7.210 3.670 ;
        RECT 6.890 3.590 7.220 3.640 ;
        RECT 6.890 3.420 7.470 3.590 ;
        RECT 6.890 3.410 7.210 3.420 ;
        RECT 8.750 3.340 8.950 3.690 ;
        RECT 8.140 2.940 8.580 3.110 ;
        RECT 1.060 1.870 1.230 2.760 ;
        RECT 3.140 1.800 6.450 2.780 ;
        RECT 6.890 2.630 7.210 2.640 ;
        RECT 6.890 2.460 7.470 2.630 ;
        RECT 6.890 2.410 7.220 2.460 ;
        RECT 6.890 2.380 7.210 2.410 ;
        RECT 8.750 2.360 8.950 2.710 ;
        RECT 6.890 2.050 7.210 2.090 ;
        RECT 6.890 2.010 7.220 2.050 ;
        RECT 6.890 1.840 7.470 2.010 ;
        RECT 6.890 1.830 7.210 1.840 ;
        RECT 8.020 1.770 8.220 2.340 ;
        RECT 8.750 2.330 8.960 2.360 ;
        RECT 8.740 1.740 8.960 2.330 ;
        RECT 1.060 0.330 1.230 1.220 ;
        RECT 3.140 0.330 6.450 1.310 ;
        RECT 6.890 1.210 7.210 1.220 ;
        RECT 6.890 1.040 7.470 1.210 ;
        RECT 6.890 1.000 7.220 1.040 ;
        RECT 6.890 0.960 7.210 1.000 ;
        RECT 8.020 0.710 8.220 1.280 ;
        RECT 8.740 0.720 8.960 1.310 ;
        RECT 8.750 0.690 8.960 0.720 ;
        RECT 6.890 0.640 7.210 0.670 ;
        RECT 6.890 0.590 7.220 0.640 ;
        RECT 6.890 0.420 7.470 0.590 ;
        RECT 6.890 0.410 7.210 0.420 ;
        RECT 8.750 0.340 8.950 0.690 ;
      LAYER mcon ;
        RECT 1.060 5.530 1.230 5.700 ;
        RECT 4.710 5.490 4.880 5.660 ;
        RECT 6.950 5.430 7.120 5.600 ;
        RECT 4.710 5.140 4.880 5.310 ;
        RECT 8.030 5.140 8.200 5.310 ;
        RECT 4.710 4.800 4.880 4.970 ;
        RECT 6.950 4.880 7.120 5.050 ;
        RECT 8.760 5.170 8.930 5.340 ;
        RECT 1.060 4.010 1.230 4.180 ;
        RECT 4.710 4.020 4.880 4.190 ;
        RECT 6.950 4.010 7.120 4.180 ;
        RECT 4.710 3.670 4.880 3.840 ;
        RECT 8.030 3.750 8.200 3.920 ;
        RECT 8.760 3.720 8.930 3.890 ;
        RECT 4.710 3.330 4.880 3.500 ;
        RECT 6.950 3.460 7.120 3.630 ;
        RECT 8.400 2.940 8.580 3.110 ;
        RECT 1.060 2.560 1.230 2.730 ;
        RECT 4.710 2.550 4.880 2.720 ;
        RECT 6.950 2.420 7.120 2.590 ;
        RECT 4.710 2.200 4.880 2.370 ;
        RECT 8.030 2.130 8.200 2.300 ;
        RECT 4.710 1.860 4.880 2.030 ;
        RECT 6.950 1.870 7.120 2.040 ;
        RECT 8.760 2.160 8.930 2.330 ;
        RECT 1.060 1.020 1.230 1.190 ;
        RECT 4.710 1.080 4.880 1.250 ;
        RECT 6.950 1.010 7.120 1.180 ;
        RECT 4.710 0.730 4.880 0.900 ;
        RECT 8.030 0.750 8.200 0.920 ;
        RECT 8.760 0.720 8.930 0.890 ;
        RECT 4.710 0.390 4.880 0.560 ;
        RECT 6.950 0.460 7.120 0.630 ;
      LAYER met1 ;
        RECT 1.010 0.000 1.280 6.050 ;
        RECT 4.670 5.080 4.910 5.720 ;
        RECT 6.880 5.360 7.200 5.680 ;
        RECT 8.020 5.370 8.180 6.050 ;
        RECT 8.020 5.350 8.220 5.370 ;
        RECT 4.680 4.820 4.910 5.080 ;
        RECT 4.680 4.600 4.920 4.820 ;
        RECT 6.880 4.810 7.200 5.130 ;
        RECT 8.000 5.110 8.230 5.350 ;
        RECT 8.020 4.890 8.220 5.110 ;
        RECT 8.390 5.060 8.580 6.050 ;
        RECT 8.830 5.400 8.990 6.050 ;
        RECT 8.410 4.940 8.580 5.060 ;
        RECT 4.670 3.610 4.910 4.250 ;
        RECT 6.880 3.930 7.200 4.250 ;
        RECT 8.020 4.170 8.180 4.890 ;
        RECT 8.020 3.950 8.220 4.170 ;
        RECT 8.420 4.120 8.580 4.940 ;
        RECT 8.720 4.850 8.990 5.400 ;
        RECT 8.720 4.800 9.000 4.850 ;
        RECT 8.830 4.710 9.000 4.800 ;
        RECT 8.830 4.350 8.990 4.710 ;
        RECT 8.830 4.260 9.000 4.350 ;
        RECT 8.410 4.000 8.580 4.120 ;
        RECT 8.000 3.710 8.230 3.950 ;
        RECT 4.680 3.350 4.910 3.610 ;
        RECT 6.880 3.380 7.200 3.700 ;
        RECT 8.020 3.690 8.220 3.710 ;
        RECT 4.680 3.130 4.920 3.350 ;
        RECT 4.670 2.140 4.910 2.780 ;
        RECT 6.880 2.350 7.200 2.670 ;
        RECT 8.020 2.360 8.180 3.690 ;
        RECT 8.390 3.140 8.580 4.000 ;
        RECT 8.720 4.210 9.000 4.260 ;
        RECT 8.720 3.660 8.990 4.210 ;
        RECT 8.370 2.910 8.610 3.140 ;
        RECT 8.020 2.340 8.220 2.360 ;
        RECT 4.680 1.880 4.910 2.140 ;
        RECT 4.680 1.660 4.920 1.880 ;
        RECT 6.880 1.800 7.200 2.120 ;
        RECT 8.000 2.100 8.230 2.340 ;
        RECT 8.020 1.880 8.220 2.100 ;
        RECT 8.390 2.050 8.580 2.910 ;
        RECT 8.830 2.390 8.990 3.660 ;
        RECT 8.410 1.930 8.580 2.050 ;
        RECT 4.670 0.670 4.910 1.310 ;
        RECT 6.880 0.930 7.200 1.250 ;
        RECT 8.020 1.170 8.180 1.880 ;
        RECT 8.020 0.950 8.220 1.170 ;
        RECT 8.420 1.120 8.580 1.930 ;
        RECT 8.720 1.840 8.990 2.390 ;
        RECT 8.720 1.790 9.000 1.840 ;
        RECT 8.830 1.700 9.000 1.790 ;
        RECT 8.830 1.350 8.990 1.700 ;
        RECT 8.830 1.260 9.000 1.350 ;
        RECT 8.410 1.000 8.580 1.120 ;
        RECT 8.000 0.710 8.230 0.950 ;
        RECT 4.680 0.410 4.910 0.670 ;
        RECT 4.680 0.190 4.920 0.410 ;
        RECT 6.880 0.380 7.200 0.700 ;
        RECT 8.020 0.690 8.220 0.710 ;
        RECT 8.020 0.010 8.180 0.690 ;
        RECT 8.390 0.010 8.580 1.000 ;
        RECT 8.720 1.210 9.000 1.260 ;
        RECT 8.720 0.660 8.990 1.210 ;
        RECT 8.830 0.010 8.990 0.660 ;
      LAYER via ;
        RECT 6.910 5.390 7.170 5.650 ;
        RECT 6.910 4.840 7.170 5.100 ;
        RECT 6.910 3.960 7.170 4.220 ;
        RECT 6.910 3.410 7.170 3.670 ;
        RECT 6.910 2.380 7.170 2.640 ;
        RECT 6.910 1.830 7.170 2.090 ;
        RECT 6.910 0.960 7.170 1.220 ;
        RECT 6.910 0.410 7.170 0.670 ;
      LAYER met2 ;
        RECT 6.880 5.550 7.190 5.690 ;
        RECT 0.000 5.370 9.350 5.550 ;
        RECT 6.880 5.360 7.190 5.370 ;
        RECT 6.880 5.120 7.190 5.140 ;
        RECT 0.000 4.940 9.350 5.120 ;
        RECT 6.880 4.810 7.190 4.940 ;
        RECT 6.880 4.120 7.190 4.250 ;
        RECT 0.000 3.940 9.350 4.120 ;
        RECT 6.880 3.920 7.190 3.940 ;
        RECT 6.880 3.690 7.190 3.700 ;
        RECT 0.000 3.620 6.870 3.690 ;
        RECT 6.880 3.620 9.350 3.690 ;
        RECT 0.000 3.510 9.350 3.620 ;
        RECT 6.880 3.370 7.190 3.510 ;
        RECT 6.880 2.540 7.190 2.680 ;
        RECT 6.880 2.530 9.350 2.540 ;
        RECT 0.000 2.360 9.350 2.530 ;
        RECT 6.880 2.350 7.190 2.360 ;
        RECT 6.880 2.110 7.190 2.130 ;
        RECT 0.000 1.940 9.350 2.110 ;
        RECT 6.790 1.930 9.350 1.940 ;
        RECT 6.880 1.800 7.190 1.930 ;
        RECT 6.880 1.130 7.190 1.250 ;
        RECT 0.000 1.120 7.190 1.130 ;
        RECT 0.000 0.960 9.350 1.120 ;
        RECT 6.790 0.940 9.350 0.960 ;
        RECT 6.880 0.920 7.190 0.940 ;
        RECT 6.880 0.690 7.190 0.700 ;
        RECT 0.000 0.520 9.350 0.690 ;
        RECT 6.880 0.510 9.350 0.520 ;
        RECT 6.880 0.370 7.190 0.510 ;
  END
END sky130_hilas_swc4x1cellOverlap2

MACRO sky130_hilas_TA2SignalBiasCell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TA2SignalBiasCell ;
  ORIGIN 5.690 -1.400 ;
  SIZE 8.880 BY 6.050 ;
  PIN VOUT_AMP2
    USE ANALOG ;
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER met2 ;
        RECT 0.270 4.970 0.580 5.020 ;
        RECT 2.570 4.970 2.880 4.990 ;
        RECT 0.270 4.740 3.190 4.970 ;
        RECT 0.270 4.690 0.580 4.740 ;
        RECT 2.570 4.660 2.880 4.740 ;
    END
  END VOUT_AMP2
  PIN VOUT_AMP1
    USE ANALOG ;
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER met2 ;
        RECT 0.270 4.140 0.580 4.200 ;
        RECT 2.560 4.140 2.870 4.270 ;
        RECT 0.270 3.920 3.190 4.140 ;
        RECT 0.270 3.870 0.580 3.920 ;
    END
  END VOUT_AMP1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 1.230 1.400 1.570 7.450 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -5.690 7.440 -1.650 7.450 ;
        RECT -5.690 1.410 -0.090 7.440 ;
        RECT -1.950 1.400 -0.090 1.410 ;
        RECT 1.910 1.400 3.190 7.450 ;
      LAYER met2 ;
        RECT -4.900 7.270 -4.660 7.450 ;
        RECT -4.940 6.980 -4.630 7.270 ;
        RECT -5.420 6.940 -4.630 6.980 ;
        RECT -5.420 6.630 -4.660 6.940 ;
        RECT -5.420 6.400 -0.880 6.630 ;
        RECT -5.420 6.160 -4.660 6.400 ;
        RECT -5.420 6.150 -4.970 6.160 ;
        RECT -1.110 6.040 -0.880 6.400 ;
        RECT 1.910 6.040 2.240 6.190 ;
        RECT -1.110 5.840 2.240 6.040 ;
        RECT -0.850 5.830 2.240 5.840 ;
        RECT 1.910 5.260 2.240 5.830 ;
        RECT -4.980 2.780 -4.670 3.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.900 6.190 2.170 7.450 ;
        RECT 1.900 5.260 2.250 6.190 ;
        RECT 1.900 3.280 2.170 5.260 ;
        RECT 1.900 2.990 2.180 3.280 ;
        RECT 1.900 1.400 2.170 2.990 ;
      LAYER via ;
        RECT 1.940 5.290 2.200 6.150 ;
    END
  END VPWR
  PIN VIN22
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -1.300 7.430 -1.050 7.440 ;
        RECT -0.700 7.430 -0.390 7.440 ;
        RECT -1.300 7.180 -0.390 7.430 ;
        RECT -0.700 7.110 -0.390 7.180 ;
    END
  END VIN22
  PIN VIN21
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -0.940 4.750 -0.630 4.790 ;
        RECT -1.030 4.740 -0.600 4.750 ;
        RECT -1.260 4.510 -0.160 4.740 ;
        RECT -0.940 4.460 -0.630 4.510 ;
    END
  END VIN21
  PIN VIN11
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -2.500 4.340 -2.190 4.390 ;
        RECT -2.820 4.110 -1.720 4.340 ;
        RECT -2.820 4.100 -2.160 4.110 ;
        RECT -2.500 4.060 -2.190 4.100 ;
    END
  END VIN11
  PIN VIN12
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -2.260 1.670 -1.950 1.740 ;
        RECT -2.860 1.420 -1.950 1.670 ;
        RECT -2.260 1.410 -1.950 1.420 ;
    END
  END VIN12
  PIN VBIAS2
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -4.010 1.670 -3.700 1.740 ;
        RECT -4.580 1.660 -3.700 1.670 ;
        RECT -5.640 1.430 -3.700 1.660 ;
        RECT -4.580 1.420 -3.700 1.430 ;
        RECT -4.010 1.410 -3.700 1.420 ;
    END
  END VBIAS2
  PIN VBIAS1
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -4.250 4.340 -3.940 4.390 ;
        RECT -5.680 4.110 -3.470 4.340 ;
        RECT -5.680 4.100 -3.910 4.110 ;
        RECT -5.680 4.090 -5.040 4.100 ;
        RECT -4.250 4.060 -3.940 4.100 ;
    END
  END VBIAS1
  OBS
      LAYER li1 ;
        RECT -0.960 7.400 -0.790 7.450 ;
        RECT -4.930 7.190 -4.610 7.230 ;
        RECT -4.930 7.000 -4.600 7.190 ;
        RECT -0.960 7.140 -0.400 7.400 ;
        RECT -0.960 7.120 -0.790 7.140 ;
        RECT 0.510 7.120 0.710 7.160 ;
        RECT -4.930 6.980 -4.610 7.000 ;
        RECT -5.020 6.970 -4.610 6.980 ;
        RECT -5.270 6.780 -4.670 6.970 ;
        RECT -5.440 6.240 -4.670 6.780 ;
        RECT -5.440 4.910 -5.270 6.240 ;
        RECT -5.430 1.970 -5.260 3.750 ;
        RECT -4.850 3.070 -4.670 6.240 ;
        RECT -4.040 5.950 -3.870 6.970 ;
        RECT -4.090 5.910 -3.770 5.950 ;
        RECT -4.090 5.720 -3.760 5.910 ;
        RECT -4.090 5.690 -3.770 5.720 ;
        RECT -4.040 5.190 -3.870 5.690 ;
        RECT -4.120 5.130 -3.580 5.190 ;
        RECT -4.120 5.020 -3.570 5.130 ;
        RECT -3.760 4.900 -3.570 5.020 ;
        RECT -4.290 4.600 -4.120 4.760 ;
        RECT -4.290 4.430 -4.070 4.600 ;
        RECT -4.240 4.350 -4.070 4.430 ;
        RECT -4.240 4.310 -3.920 4.350 ;
        RECT -4.240 4.120 -3.910 4.310 ;
        RECT -4.240 4.090 -3.920 4.120 ;
        RECT -4.970 3.030 -4.650 3.070 ;
        RECT -4.970 2.840 -4.640 3.030 ;
        RECT -4.970 2.810 -4.650 2.840 ;
        RECT -4.850 1.880 -4.670 2.810 ;
        RECT -4.040 2.540 -3.870 3.920 ;
        RECT -3.100 3.070 -2.920 6.980 ;
        RECT -2.290 5.190 -2.120 6.970 ;
        RECT -1.540 6.040 -1.360 6.970 ;
        RECT -0.810 6.710 -0.480 6.880 ;
        RECT 0.280 6.860 0.710 7.120 ;
        RECT 0.510 6.830 0.710 6.860 ;
        RECT -0.730 6.570 -0.480 6.710 ;
        RECT -0.730 6.310 -0.250 6.570 ;
        RECT 0.100 6.470 0.270 6.510 ;
        RECT 0.510 6.470 0.710 6.500 ;
        RECT -1.660 6.010 -1.340 6.040 ;
        RECT -1.660 5.820 -1.330 6.010 ;
        RECT -1.660 5.780 -1.340 5.820 ;
        RECT -2.370 5.130 -1.830 5.190 ;
        RECT -2.370 5.020 -1.820 5.130 ;
        RECT -2.010 4.900 -1.820 5.020 ;
        RECT -2.540 4.600 -2.370 4.760 ;
        RECT -2.540 4.430 -2.320 4.600 ;
        RECT -2.490 4.350 -2.320 4.430 ;
        RECT -2.490 4.310 -2.170 4.350 ;
        RECT -2.490 4.120 -2.160 4.310 ;
        RECT -2.490 4.090 -2.170 4.120 ;
        RECT -3.220 3.030 -2.900 3.070 ;
        RECT -3.220 2.840 -2.890 3.030 ;
        RECT -3.220 2.810 -2.900 2.840 ;
        RECT -4.040 2.280 -3.560 2.540 ;
        RECT -4.040 2.140 -3.790 2.280 ;
        RECT -4.120 1.970 -3.790 2.140 ;
        RECT -3.100 1.880 -2.920 2.810 ;
        RECT -2.290 2.540 -2.120 3.920 ;
        RECT -2.290 2.280 -1.810 2.540 ;
        RECT -2.290 2.140 -2.040 2.280 ;
        RECT -2.370 1.970 -2.040 2.140 ;
        RECT -1.540 1.870 -1.360 5.780 ;
        RECT -0.730 4.930 -0.560 6.310 ;
        RECT 0.100 6.210 0.710 6.470 ;
        RECT 0.100 6.180 0.270 6.210 ;
        RECT 0.510 6.170 0.710 6.210 ;
        RECT 1.100 6.170 1.650 7.160 ;
        RECT 2.470 7.040 3.050 7.210 ;
        RECT 2.470 6.940 2.860 7.040 ;
        RECT 2.470 6.910 2.850 6.940 ;
        RECT 2.470 6.760 2.830 6.910 ;
        RECT 2.120 6.590 2.830 6.760 ;
        RECT 0.100 5.640 0.270 5.670 ;
        RECT 0.510 5.640 0.710 5.680 ;
        RECT 0.100 5.380 0.710 5.640 ;
        RECT 0.100 5.340 0.270 5.380 ;
        RECT 0.510 5.350 0.710 5.380 ;
        RECT 0.510 4.990 0.710 5.020 ;
        RECT -0.930 4.730 -0.610 4.760 ;
        RECT 0.280 4.730 0.710 4.990 ;
        RECT -0.930 4.540 -0.600 4.730 ;
        RECT 0.510 4.690 0.710 4.730 ;
        RECT 1.100 4.690 1.650 5.680 ;
        RECT 1.960 5.270 2.820 6.150 ;
        RECT 1.960 5.260 2.170 5.270 ;
        RECT 2.580 4.910 2.900 4.950 ;
        RECT 2.580 4.850 2.910 4.910 ;
        RECT 2.110 4.720 2.910 4.850 ;
        RECT 2.110 4.690 2.900 4.720 ;
        RECT 2.110 4.670 2.810 4.690 ;
        RECT -0.930 4.500 -0.610 4.540 ;
        RECT -0.930 4.420 -0.760 4.500 ;
        RECT -0.980 4.250 -0.760 4.420 ;
        RECT -0.980 4.090 -0.810 4.250 ;
        RECT 0.510 4.160 0.710 4.200 ;
        RECT -0.450 3.830 -0.260 3.950 ;
        RECT 0.280 3.900 0.710 4.160 ;
        RECT 0.510 3.870 0.710 3.900 ;
        RECT -0.810 3.720 -0.260 3.830 ;
        RECT -0.810 3.660 -0.270 3.720 ;
        RECT -0.730 1.880 -0.560 3.660 ;
        RECT 0.100 3.510 0.270 3.550 ;
        RECT 0.510 3.510 0.710 3.540 ;
        RECT 0.100 3.250 0.710 3.510 ;
        RECT 0.100 3.220 0.270 3.250 ;
        RECT 0.510 3.210 0.710 3.250 ;
        RECT 1.100 3.210 1.650 4.200 ;
        RECT 2.570 4.190 2.890 4.230 ;
        RECT 2.110 4.010 2.900 4.190 ;
        RECT 2.570 4.000 2.900 4.010 ;
        RECT 2.570 3.970 2.890 4.000 ;
        RECT 2.120 3.250 2.820 3.590 ;
        RECT 1.970 3.020 2.820 3.250 ;
        RECT 0.100 2.680 0.270 2.710 ;
        RECT 0.510 2.680 0.710 2.720 ;
        RECT 0.100 2.420 0.710 2.680 ;
        RECT 0.100 2.380 0.270 2.420 ;
        RECT 0.510 2.390 0.710 2.420 ;
        RECT 0.510 2.030 0.710 2.060 ;
        RECT 0.280 1.770 0.710 2.030 ;
        RECT 0.510 1.730 0.710 1.770 ;
        RECT 1.100 1.730 1.650 2.720 ;
        RECT 2.120 2.710 2.820 3.020 ;
        RECT 2.120 2.100 2.830 2.270 ;
        RECT 2.470 1.820 2.830 2.100 ;
        RECT -4.270 1.710 -4.100 1.730 ;
        RECT -2.520 1.710 -2.350 1.730 ;
        RECT -4.270 1.450 -3.710 1.710 ;
        RECT -2.520 1.450 -1.960 1.710 ;
        RECT 2.470 1.650 3.050 1.820 ;
        RECT -4.270 1.400 -4.100 1.450 ;
        RECT -2.520 1.400 -2.350 1.450 ;
      LAYER mcon ;
        RECT -4.870 7.010 -4.700 7.180 ;
        RECT -0.630 7.180 -0.460 7.350 ;
        RECT -5.440 6.610 -5.270 6.780 ;
        RECT -4.850 6.560 -4.680 6.730 ;
        RECT -5.440 6.270 -5.270 6.440 ;
        RECT -5.440 5.930 -5.270 6.100 ;
        RECT -5.440 5.590 -5.270 5.760 ;
        RECT -5.440 5.250 -5.270 5.420 ;
        RECT -4.850 6.220 -4.680 6.390 ;
        RECT -5.430 3.580 -5.260 3.750 ;
        RECT -5.430 3.240 -5.260 3.410 ;
        RECT -4.030 5.730 -3.860 5.900 ;
        RECT -3.750 4.930 -3.580 5.100 ;
        RECT -4.180 4.130 -4.010 4.300 ;
        RECT -5.430 2.900 -5.260 3.070 ;
        RECT -4.910 2.850 -4.740 3.020 ;
        RECT -5.430 2.560 -5.260 2.730 ;
        RECT -5.430 2.220 -5.260 2.390 ;
        RECT 0.340 6.900 0.510 7.070 ;
        RECT 2.590 6.950 2.760 7.120 ;
        RECT 1.320 6.580 1.490 6.750 ;
        RECT -0.480 6.350 -0.310 6.520 ;
        RECT -1.600 5.830 -1.430 6.000 ;
        RECT -2.000 4.930 -1.830 5.100 ;
        RECT -2.430 4.130 -2.260 4.300 ;
        RECT -3.160 2.850 -2.990 3.020 ;
        RECT -3.790 2.330 -3.620 2.500 ;
        RECT -2.040 2.330 -1.870 2.500 ;
        RECT 0.290 6.250 0.460 6.420 ;
        RECT 1.980 5.980 2.150 6.150 ;
        RECT 0.290 5.430 0.460 5.600 ;
        RECT 1.320 5.100 1.490 5.270 ;
        RECT 1.980 5.640 2.150 5.810 ;
        RECT 1.980 5.280 2.150 5.450 ;
        RECT 0.340 4.780 0.510 4.950 ;
        RECT -0.870 4.550 -0.700 4.720 ;
        RECT 2.640 4.730 2.810 4.900 ;
        RECT -0.440 3.750 -0.270 3.920 ;
        RECT 0.340 3.940 0.510 4.110 ;
        RECT 2.630 4.010 2.800 4.180 ;
        RECT 1.320 3.620 1.490 3.790 ;
        RECT 0.290 3.290 0.460 3.460 ;
        RECT 1.980 3.050 2.150 3.220 ;
        RECT 0.290 2.470 0.460 2.640 ;
        RECT 1.320 2.140 1.490 2.310 ;
        RECT 0.340 1.820 0.510 1.990 ;
        RECT 2.550 1.760 2.720 1.930 ;
        RECT -3.940 1.500 -3.770 1.670 ;
        RECT -2.190 1.500 -2.020 1.670 ;
      LAYER met1 ;
        RECT -4.940 6.990 -4.620 7.260 ;
        RECT -0.710 7.110 -0.390 7.430 ;
        RECT -5.470 6.940 -4.620 6.990 ;
        RECT -5.470 6.670 -4.650 6.940 ;
        RECT 0.270 6.830 0.590 7.150 ;
        RECT 2.520 6.880 2.840 7.200 ;
        RECT -5.470 6.380 -4.620 6.670 ;
        RECT -5.470 6.130 -4.650 6.380 ;
        RECT -0.560 6.280 -0.240 6.600 ;
        RECT 0.220 6.180 0.540 6.500 ;
        RECT -5.470 3.100 -4.830 6.130 ;
        RECT -4.100 5.660 -3.780 5.980 ;
        RECT -1.670 5.750 -1.350 6.070 ;
        RECT -0.450 5.590 -0.240 5.700 ;
        RECT -0.470 5.270 -0.210 5.590 ;
        RECT 0.220 5.350 0.540 5.670 ;
        RECT -3.780 4.870 -3.550 5.160 ;
        RECT -2.030 4.870 -1.800 5.160 ;
        RECT -4.250 4.060 -3.930 4.380 ;
        RECT -3.760 3.580 -3.550 4.870 ;
        RECT -2.500 4.060 -2.180 4.380 ;
        RECT -2.010 3.580 -1.800 4.870 ;
        RECT -0.940 4.470 -0.620 4.790 ;
        RECT -0.450 3.980 -0.240 5.270 ;
        RECT 0.270 4.700 0.590 5.020 ;
        RECT 2.570 4.660 2.890 4.980 ;
        RECT -0.470 3.690 -0.240 3.980 ;
        RECT 0.270 3.870 0.590 4.190 ;
        RECT 2.560 3.940 2.880 4.260 ;
        RECT -3.780 3.260 -3.520 3.580 ;
        RECT -2.030 3.260 -1.770 3.580 ;
        RECT -3.760 3.150 -3.550 3.260 ;
        RECT -2.010 3.150 -1.800 3.260 ;
        RECT 0.220 3.220 0.540 3.540 ;
        RECT -5.470 2.780 -4.660 3.100 ;
        RECT -3.230 2.780 -2.910 3.100 ;
        RECT -5.470 1.950 -4.830 2.780 ;
        RECT -3.870 2.250 -3.550 2.570 ;
        RECT -2.120 2.250 -1.800 2.570 ;
        RECT 0.220 2.390 0.540 2.710 ;
        RECT -5.250 1.940 -4.830 1.950 ;
        RECT 0.270 1.740 0.590 2.060 ;
        RECT -4.020 1.420 -3.700 1.740 ;
        RECT -2.270 1.420 -1.950 1.740 ;
        RECT 2.480 1.690 2.800 2.010 ;
      LAYER via ;
        RECT -4.910 6.970 -4.650 7.230 ;
        RECT -0.680 7.140 -0.420 7.400 ;
        RECT -5.350 6.190 -4.760 6.910 ;
        RECT 0.300 6.860 0.560 7.120 ;
        RECT 2.550 6.910 2.810 7.170 ;
        RECT -0.530 6.310 -0.270 6.570 ;
        RECT 0.250 6.210 0.510 6.470 ;
        RECT -4.070 5.690 -3.810 5.950 ;
        RECT -1.640 5.780 -1.380 6.040 ;
        RECT -0.470 5.300 -0.210 5.560 ;
        RECT 0.250 5.380 0.510 5.640 ;
        RECT -4.220 4.090 -3.960 4.350 ;
        RECT -2.470 4.090 -2.210 4.350 ;
        RECT -0.910 4.500 -0.650 4.760 ;
        RECT 0.300 4.730 0.560 4.990 ;
        RECT 2.600 4.690 2.860 4.950 ;
        RECT 0.300 3.900 0.560 4.160 ;
        RECT 2.590 3.970 2.850 4.230 ;
        RECT -3.780 3.290 -3.520 3.550 ;
        RECT -2.030 3.290 -1.770 3.550 ;
        RECT 0.250 3.250 0.510 3.510 ;
        RECT -4.950 2.810 -4.690 3.070 ;
        RECT -3.200 2.810 -2.940 3.070 ;
        RECT -3.840 2.280 -3.580 2.540 ;
        RECT -2.090 2.280 -1.830 2.540 ;
        RECT 0.250 2.420 0.510 2.680 ;
        RECT 0.300 1.770 0.560 2.030 ;
        RECT -3.990 1.450 -3.730 1.710 ;
        RECT -2.240 1.450 -1.980 1.710 ;
        RECT 2.510 1.720 2.770 1.980 ;
      LAYER met2 ;
        RECT 0.270 7.110 0.580 7.160 ;
        RECT 2.520 7.110 2.830 7.210 ;
        RECT 0.270 6.880 2.830 7.110 ;
        RECT 0.270 6.830 0.580 6.880 ;
        RECT -0.550 6.570 -0.240 6.610 ;
        RECT -0.730 6.430 0.010 6.570 ;
        RECT 0.220 6.430 0.530 6.510 ;
        RECT -0.730 6.320 0.530 6.430 ;
        RECT -0.550 6.280 0.530 6.320 ;
        RECT -0.240 6.220 0.530 6.280 ;
        RECT -0.240 6.200 0.010 6.220 ;
        RECT 0.220 6.180 0.530 6.220 ;
        RECT -4.100 5.930 -3.790 5.990 ;
        RECT -1.670 5.930 -1.360 6.070 ;
        RECT -4.100 5.740 -1.360 5.930 ;
        RECT -4.100 5.710 -1.620 5.740 ;
        RECT -4.100 5.660 -3.790 5.710 ;
        RECT -0.210 5.630 0.000 5.640 ;
        RECT 0.220 5.630 0.530 5.670 ;
        RECT -0.210 5.560 0.530 5.630 ;
        RECT -0.500 5.540 0.530 5.560 ;
        RECT -0.550 5.420 0.530 5.540 ;
        RECT -0.550 5.350 0.000 5.420 ;
        RECT -0.550 5.290 -0.080 5.350 ;
        RECT 0.220 5.340 0.530 5.420 ;
        RECT -3.860 3.310 -3.390 3.560 ;
        RECT -2.110 3.470 -1.640 3.560 ;
        RECT 0.220 3.470 0.530 3.550 ;
        RECT -2.110 3.310 0.530 3.470 ;
        RECT -3.810 3.290 -3.490 3.310 ;
        RECT -2.060 3.290 0.530 3.310 ;
        RECT -1.770 3.270 0.530 3.290 ;
        RECT -0.080 3.260 0.530 3.270 ;
        RECT 0.220 3.220 0.530 3.260 ;
        RECT -3.230 3.100 -2.920 3.110 ;
        RECT -3.340 2.920 -2.920 3.100 ;
        RECT -3.360 2.910 -2.920 2.920 ;
        RECT -3.580 2.780 -2.920 2.910 ;
        RECT -3.580 2.570 -3.220 2.780 ;
        RECT 0.220 2.670 0.530 2.710 ;
        RECT -2.060 2.570 0.530 2.670 ;
        RECT -3.860 2.530 -3.220 2.570 ;
        RECT -2.110 2.530 0.530 2.570 ;
        RECT -4.040 2.290 -3.220 2.530 ;
        RECT -2.290 2.460 0.530 2.530 ;
        RECT -4.040 2.280 -3.490 2.290 ;
        RECT -2.290 2.280 -1.740 2.460 ;
        RECT 0.220 2.380 0.530 2.460 ;
        RECT -3.860 2.240 -3.550 2.280 ;
        RECT -2.110 2.240 -1.800 2.280 ;
        RECT 0.270 1.980 0.580 2.060 ;
        RECT 2.480 1.980 2.790 2.020 ;
        RECT 0.270 1.750 2.980 1.980 ;
        RECT 0.270 1.730 0.580 1.750 ;
        RECT 2.480 1.690 2.790 1.750 ;
  END
END sky130_hilas_TA2SignalBiasCell

MACRO sky130_hilas_Tgate4Single01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_Tgate4Single01 ;
  ORIGIN 0.360 1.410 ;
  SIZE 4.760 BY 6.050 ;
  PIN INPUT1_4
    USE ANALOG ;
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 1.280 -1.090 1.590 -0.970 ;
        RECT 0.510 -1.100 1.630 -1.090 ;
        RECT 2.850 -1.100 3.160 -0.970 ;
        RECT -0.360 -1.300 3.160 -1.100 ;
        RECT 0.510 -1.310 1.630 -1.300 ;
    END
  END INPUT1_4
  PIN VPWR
    USE ANALOG ;
    ANTENNADIFFAREA 0.908800 ;
    PORT
      LAYER nwell ;
        RECT -0.240 -1.410 2.520 4.640 ;
      LAYER met1 ;
        RECT 0.380 3.770 0.580 4.640 ;
        RECT 0.370 3.480 0.600 3.770 ;
        RECT 0.380 2.770 0.580 3.480 ;
        RECT 0.370 2.480 0.600 2.770 ;
        RECT 0.380 0.750 0.580 2.480 ;
        RECT 0.370 0.460 0.600 0.750 ;
        RECT 0.380 -0.250 0.580 0.460 ;
        RECT 0.370 -0.540 0.600 -0.250 ;
        RECT 0.380 -1.410 0.580 -0.540 ;
    END
  END VPWR
  PIN SELECT4
    USE ANALOG ;
    ANTENNAGATEAREA 0.372000 ;
    PORT
      LAYER met2 ;
        RECT -0.070 -0.120 0.250 -0.030 ;
        RECT -0.360 -0.320 0.250 -0.120 ;
    END
  END SELECT4
  PIN SELECT3
    USE ANALOG ;
    ANTENNAGATEAREA 0.372000 ;
    PORT
      LAYER met2 ;
        RECT -0.360 0.330 0.250 0.530 ;
        RECT -0.070 0.240 0.250 0.330 ;
    END
  END SELECT3
  PIN INPUT1_3
    USE ANALOG ;
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 0.510 1.510 1.630 1.520 ;
        RECT -0.360 1.310 3.160 1.510 ;
        RECT 0.510 1.300 1.630 1.310 ;
        RECT 1.280 1.180 1.590 1.300 ;
        RECT 2.850 1.180 3.160 1.310 ;
    END
  END INPUT1_3
  PIN INPUT1_2
    USE ANALOG ;
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 1.280 1.930 1.590 2.050 ;
        RECT 0.510 1.920 1.630 1.930 ;
        RECT 2.850 1.920 3.160 2.050 ;
        RECT -0.360 1.720 3.160 1.920 ;
        RECT 0.510 1.710 1.630 1.720 ;
    END
  END INPUT1_2
  PIN SELECT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.372000 ;
    PORT
      LAYER met2 ;
        RECT -0.070 2.900 0.250 2.990 ;
        RECT -0.360 2.700 0.250 2.900 ;
    END
  END SELECT2
  PIN SELECT1
    USE ANALOG ;
    ANTENNAGATEAREA 0.372000 ;
    PORT
      LAYER met2 ;
        RECT -0.360 3.350 0.250 3.550 ;
        RECT -0.070 3.260 0.250 3.350 ;
    END
  END SELECT1
  PIN INPUT1_1
    USE ANALOG ;
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 0.510 4.530 1.630 4.540 ;
        RECT -0.360 4.330 3.160 4.530 ;
        RECT 0.510 4.320 1.630 4.330 ;
        RECT 1.280 4.200 1.590 4.320 ;
        RECT 2.850 4.200 3.160 4.330 ;
    END
  END INPUT1_1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 3.890 3.770 4.080 4.640 ;
        RECT 3.870 3.480 4.100 3.770 ;
        RECT 3.890 2.770 4.080 3.480 ;
        RECT 3.870 2.480 4.100 2.770 ;
        RECT 3.890 0.750 4.080 2.480 ;
        RECT 3.870 0.460 4.100 0.750 ;
        RECT 3.890 -0.250 4.080 0.460 ;
        RECT 3.870 -0.540 4.100 -0.250 ;
        RECT 3.890 -1.410 4.080 -0.540 ;
    END
  END VGND
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.182900 ;
    PORT
      LAYER met2 ;
        RECT 2.200 3.550 2.520 3.590 ;
        RECT 3.210 3.550 3.530 3.580 ;
        RECT 2.150 3.350 4.400 3.550 ;
        RECT 2.200 3.330 2.520 3.350 ;
        RECT 3.210 3.320 3.530 3.350 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.182900 ;
    PORT
      LAYER met2 ;
        RECT 2.200 2.900 2.520 2.920 ;
        RECT 3.210 2.900 3.530 2.930 ;
        RECT 2.150 2.700 4.400 2.900 ;
        RECT 2.200 2.660 2.520 2.700 ;
        RECT 3.210 2.670 3.530 2.700 ;
    END
  END OUTPUT2
  PIN OUTPUT3
    USE ANALOG ;
    ANTENNADIFFAREA 0.182900 ;
    PORT
      LAYER met2 ;
        RECT 2.200 0.530 2.520 0.570 ;
        RECT 3.210 0.530 3.530 0.560 ;
        RECT 2.150 0.330 4.400 0.530 ;
        RECT 2.200 0.310 2.520 0.330 ;
        RECT 3.210 0.300 3.530 0.330 ;
    END
  END OUTPUT3
  PIN OUTPUT4
    USE ANALOG ;
    ANTENNADIFFAREA 0.182900 ;
    PORT
      LAYER met2 ;
        RECT 2.200 -0.120 2.520 -0.100 ;
        RECT 3.210 -0.120 3.530 -0.090 ;
        RECT 2.150 -0.320 4.400 -0.120 ;
        RECT 2.200 -0.360 2.520 -0.320 ;
        RECT 3.210 -0.350 3.530 -0.320 ;
    END
  END OUTPUT4
  OBS
      LAYER li1 ;
        RECT 1.290 4.470 1.610 4.500 ;
        RECT 2.860 4.470 3.180 4.500 ;
        RECT 0.070 4.130 0.240 4.410 ;
        RECT 1.290 4.280 1.620 4.470 ;
        RECT 2.300 4.330 2.490 4.350 ;
        RECT 1.290 4.240 1.610 4.280 ;
        RECT 0.070 4.090 0.280 4.130 ;
        RECT 0.070 4.070 0.300 4.090 ;
        RECT 1.420 4.080 1.590 4.240 ;
        RECT 2.030 4.160 2.490 4.330 ;
        RECT 2.860 4.280 3.190 4.470 ;
        RECT 3.430 4.330 3.620 4.360 ;
        RECT 2.860 4.240 3.180 4.280 ;
        RECT 2.280 4.150 2.490 4.160 ;
        RECT 2.300 4.120 2.490 4.150 ;
        RECT 2.920 4.080 3.090 4.240 ;
        RECT 3.430 4.160 3.870 4.330 ;
        RECT 3.430 4.130 3.620 4.160 ;
        RECT 0.070 4.050 0.330 4.070 ;
        RECT 0.070 4.000 0.410 4.050 ;
        RECT 0.070 3.940 0.560 4.000 ;
        RECT 0.070 3.910 0.580 3.940 ;
        RECT 0.110 3.880 0.580 3.910 ;
        RECT 0.240 3.830 0.580 3.880 ;
        RECT 0.360 3.820 0.580 3.830 ;
        RECT 0.370 3.790 0.580 3.820 ;
        RECT 0.390 3.710 0.580 3.790 ;
        RECT 1.750 3.710 2.080 3.830 ;
        RECT 4.150 3.740 4.320 4.420 ;
        RECT -0.100 3.660 0.070 3.680 ;
        RECT -0.120 3.230 0.090 3.660 ;
        RECT 0.390 3.540 0.910 3.710 ;
        RECT 0.390 3.510 0.580 3.540 ;
        RECT 1.260 3.530 3.160 3.710 ;
        RECT 3.890 3.700 4.320 3.740 ;
        RECT 3.540 3.540 4.320 3.700 ;
        RECT 3.540 3.530 4.080 3.540 ;
        RECT 3.890 3.510 4.080 3.530 ;
        RECT -0.120 2.590 0.090 3.020 ;
        RECT 0.390 2.710 0.580 2.740 ;
        RECT 3.890 2.720 4.080 2.740 ;
        RECT -0.100 2.570 0.070 2.590 ;
        RECT 0.390 2.540 0.910 2.710 ;
        RECT 1.260 2.540 3.160 2.720 ;
        RECT 3.540 2.710 4.080 2.720 ;
        RECT 3.540 2.550 4.320 2.710 ;
        RECT 0.390 2.460 0.580 2.540 ;
        RECT 0.370 2.430 0.580 2.460 ;
        RECT 0.360 2.420 0.580 2.430 ;
        RECT 1.750 2.420 2.080 2.540 ;
        RECT 3.890 2.510 4.320 2.550 ;
        RECT 0.240 2.370 0.580 2.420 ;
        RECT 0.110 2.340 0.580 2.370 ;
        RECT 0.070 2.310 0.580 2.340 ;
        RECT 0.070 2.250 0.560 2.310 ;
        RECT 0.070 2.200 0.410 2.250 ;
        RECT 0.070 2.180 0.330 2.200 ;
        RECT 0.070 2.160 0.300 2.180 ;
        RECT 0.070 2.120 0.280 2.160 ;
        RECT 0.070 1.840 0.240 2.120 ;
        RECT 1.420 2.010 1.590 2.170 ;
        RECT 2.300 2.100 2.490 2.130 ;
        RECT 2.280 2.090 2.490 2.100 ;
        RECT 1.290 1.970 1.610 2.010 ;
        RECT 1.290 1.780 1.620 1.970 ;
        RECT 2.030 1.920 2.490 2.090 ;
        RECT 2.920 2.010 3.090 2.170 ;
        RECT 3.430 2.090 3.620 2.120 ;
        RECT 2.300 1.900 2.490 1.920 ;
        RECT 2.860 1.970 3.180 2.010 ;
        RECT 2.860 1.780 3.190 1.970 ;
        RECT 3.430 1.920 3.870 2.090 ;
        RECT 3.430 1.890 3.620 1.920 ;
        RECT 4.150 1.830 4.320 2.510 ;
        RECT 1.290 1.750 1.610 1.780 ;
        RECT 2.860 1.750 3.180 1.780 ;
        RECT 1.290 1.450 1.610 1.480 ;
        RECT 2.860 1.450 3.180 1.480 ;
        RECT 0.070 1.110 0.240 1.390 ;
        RECT 1.290 1.260 1.620 1.450 ;
        RECT 2.300 1.310 2.490 1.330 ;
        RECT 1.290 1.220 1.610 1.260 ;
        RECT 0.070 1.070 0.280 1.110 ;
        RECT 0.070 1.050 0.300 1.070 ;
        RECT 1.420 1.060 1.590 1.220 ;
        RECT 2.030 1.140 2.490 1.310 ;
        RECT 2.860 1.260 3.190 1.450 ;
        RECT 3.430 1.310 3.620 1.340 ;
        RECT 2.860 1.220 3.180 1.260 ;
        RECT 2.280 1.130 2.490 1.140 ;
        RECT 2.300 1.100 2.490 1.130 ;
        RECT 2.920 1.060 3.090 1.220 ;
        RECT 3.430 1.140 3.870 1.310 ;
        RECT 3.430 1.110 3.620 1.140 ;
        RECT 0.070 1.030 0.330 1.050 ;
        RECT 0.070 0.980 0.410 1.030 ;
        RECT 0.070 0.920 0.560 0.980 ;
        RECT 0.070 0.890 0.580 0.920 ;
        RECT 0.110 0.860 0.580 0.890 ;
        RECT 0.240 0.810 0.580 0.860 ;
        RECT 0.360 0.800 0.580 0.810 ;
        RECT 0.370 0.770 0.580 0.800 ;
        RECT 0.390 0.690 0.580 0.770 ;
        RECT 1.750 0.690 2.080 0.810 ;
        RECT 4.150 0.720 4.320 1.400 ;
        RECT -0.100 0.640 0.070 0.660 ;
        RECT -0.120 0.210 0.090 0.640 ;
        RECT 0.390 0.520 0.910 0.690 ;
        RECT 0.390 0.490 0.580 0.520 ;
        RECT 1.260 0.510 3.160 0.690 ;
        RECT 3.890 0.680 4.320 0.720 ;
        RECT 3.540 0.520 4.320 0.680 ;
        RECT 3.540 0.510 4.080 0.520 ;
        RECT 3.890 0.490 4.080 0.510 ;
        RECT -0.120 -0.430 0.090 0.000 ;
        RECT 0.390 -0.310 0.580 -0.280 ;
        RECT 3.890 -0.300 4.080 -0.280 ;
        RECT -0.100 -0.450 0.070 -0.430 ;
        RECT 0.390 -0.480 0.910 -0.310 ;
        RECT 1.260 -0.480 3.160 -0.300 ;
        RECT 3.540 -0.310 4.080 -0.300 ;
        RECT 3.540 -0.470 4.320 -0.310 ;
        RECT 0.390 -0.560 0.580 -0.480 ;
        RECT 0.370 -0.590 0.580 -0.560 ;
        RECT 0.360 -0.600 0.580 -0.590 ;
        RECT 1.750 -0.600 2.080 -0.480 ;
        RECT 3.890 -0.510 4.320 -0.470 ;
        RECT 0.240 -0.650 0.580 -0.600 ;
        RECT 0.110 -0.680 0.580 -0.650 ;
        RECT 0.070 -0.710 0.580 -0.680 ;
        RECT 0.070 -0.770 0.560 -0.710 ;
        RECT 0.070 -0.820 0.410 -0.770 ;
        RECT 0.070 -0.840 0.330 -0.820 ;
        RECT 0.070 -0.860 0.300 -0.840 ;
        RECT 0.070 -0.900 0.280 -0.860 ;
        RECT 0.070 -1.180 0.240 -0.900 ;
        RECT 1.420 -1.010 1.590 -0.850 ;
        RECT 2.300 -0.920 2.490 -0.890 ;
        RECT 2.280 -0.930 2.490 -0.920 ;
        RECT 1.290 -1.050 1.610 -1.010 ;
        RECT 1.290 -1.240 1.620 -1.050 ;
        RECT 2.030 -1.100 2.490 -0.930 ;
        RECT 2.920 -1.010 3.090 -0.850 ;
        RECT 3.430 -0.930 3.620 -0.900 ;
        RECT 2.300 -1.120 2.490 -1.100 ;
        RECT 2.860 -1.050 3.180 -1.010 ;
        RECT 2.860 -1.240 3.190 -1.050 ;
        RECT 3.430 -1.100 3.870 -0.930 ;
        RECT 3.430 -1.130 3.620 -1.100 ;
        RECT 4.150 -1.190 4.320 -0.510 ;
        RECT 1.290 -1.270 1.610 -1.240 ;
        RECT 2.860 -1.270 3.180 -1.240 ;
      LAYER mcon ;
        RECT 1.350 4.290 1.520 4.460 ;
        RECT 2.310 4.150 2.480 4.320 ;
        RECT 2.920 4.290 3.090 4.460 ;
        RECT 3.440 4.160 3.610 4.330 ;
        RECT -0.100 3.510 0.070 3.680 ;
        RECT 0.400 3.540 0.570 3.710 ;
        RECT 3.900 3.540 4.070 3.710 ;
        RECT 0.400 2.540 0.570 2.710 ;
        RECT 3.900 2.540 4.070 2.710 ;
        RECT 1.350 1.790 1.520 1.960 ;
        RECT 2.310 1.930 2.480 2.100 ;
        RECT 2.920 1.790 3.090 1.960 ;
        RECT 3.440 1.920 3.610 2.090 ;
        RECT 1.350 1.270 1.520 1.440 ;
        RECT 2.310 1.130 2.480 1.300 ;
        RECT 2.920 1.270 3.090 1.440 ;
        RECT 3.440 1.140 3.610 1.310 ;
        RECT -0.100 0.490 0.070 0.660 ;
        RECT 0.400 0.520 0.570 0.690 ;
        RECT 3.900 0.520 4.070 0.690 ;
        RECT 0.400 -0.480 0.570 -0.310 ;
        RECT 3.900 -0.480 4.070 -0.310 ;
        RECT 1.350 -1.230 1.520 -1.060 ;
        RECT 2.310 -1.090 2.480 -0.920 ;
        RECT 2.920 -1.230 3.090 -1.060 ;
        RECT 3.440 -1.100 3.610 -0.930 ;
      LAYER met1 ;
        RECT 1.280 4.210 1.600 4.530 ;
        RECT 2.280 4.090 2.510 4.380 ;
        RECT 2.850 4.210 3.170 4.530 ;
        RECT 3.410 4.100 3.640 4.390 ;
        RECT -0.130 3.550 0.100 3.740 ;
        RECT 2.300 3.620 2.490 4.090 ;
        RECT -0.130 3.450 0.220 3.550 ;
        RECT -0.120 3.230 0.220 3.450 ;
        RECT 2.230 3.300 2.490 3.620 ;
        RECT 3.410 3.610 3.600 4.100 ;
        RECT 3.240 3.360 3.600 3.610 ;
        RECT 3.240 3.290 3.500 3.360 ;
        RECT -0.120 2.800 0.220 3.020 ;
        RECT -0.130 2.700 0.220 2.800 ;
        RECT -0.130 2.510 0.100 2.700 ;
        RECT 2.230 2.630 2.490 2.950 ;
        RECT 3.240 2.890 3.500 2.960 ;
        RECT 3.240 2.640 3.600 2.890 ;
        RECT 2.300 2.160 2.490 2.630 ;
        RECT 1.280 1.720 1.600 2.040 ;
        RECT 2.280 1.870 2.510 2.160 ;
        RECT 3.410 2.150 3.600 2.640 ;
        RECT 2.850 1.720 3.170 2.040 ;
        RECT 3.410 1.860 3.640 2.150 ;
        RECT 1.280 1.190 1.600 1.510 ;
        RECT 2.280 1.070 2.510 1.360 ;
        RECT 2.850 1.190 3.170 1.510 ;
        RECT 3.410 1.080 3.640 1.370 ;
        RECT -0.130 0.530 0.100 0.720 ;
        RECT 2.300 0.600 2.490 1.070 ;
        RECT -0.130 0.430 0.220 0.530 ;
        RECT -0.120 0.210 0.220 0.430 ;
        RECT 2.230 0.280 2.490 0.600 ;
        RECT 3.410 0.590 3.600 1.080 ;
        RECT 3.240 0.340 3.600 0.590 ;
        RECT 3.240 0.270 3.500 0.340 ;
        RECT -0.120 -0.220 0.220 0.000 ;
        RECT -0.130 -0.320 0.220 -0.220 ;
        RECT -0.130 -0.510 0.100 -0.320 ;
        RECT 2.230 -0.390 2.490 -0.070 ;
        RECT 3.240 -0.130 3.500 -0.060 ;
        RECT 3.240 -0.380 3.600 -0.130 ;
        RECT 2.300 -0.860 2.490 -0.390 ;
        RECT 1.280 -1.300 1.600 -0.980 ;
        RECT 2.280 -1.150 2.510 -0.860 ;
        RECT 3.410 -0.870 3.600 -0.380 ;
        RECT 2.850 -1.300 3.170 -0.980 ;
        RECT 3.410 -1.160 3.640 -0.870 ;
      LAYER via ;
        RECT 1.310 4.240 1.570 4.500 ;
        RECT 2.880 4.240 3.140 4.500 ;
        RECT -0.040 3.260 0.220 3.520 ;
        RECT 2.230 3.330 2.490 3.590 ;
        RECT 3.240 3.320 3.500 3.580 ;
        RECT -0.040 2.730 0.220 2.990 ;
        RECT 2.230 2.660 2.490 2.920 ;
        RECT 3.240 2.670 3.500 2.930 ;
        RECT 1.310 1.750 1.570 2.010 ;
        RECT 2.880 1.750 3.140 2.010 ;
        RECT 1.310 1.220 1.570 1.480 ;
        RECT 2.880 1.220 3.140 1.480 ;
        RECT -0.040 0.240 0.220 0.500 ;
        RECT 2.230 0.310 2.490 0.570 ;
        RECT 3.240 0.300 3.500 0.560 ;
        RECT -0.040 -0.290 0.220 -0.030 ;
        RECT 2.230 -0.360 2.490 -0.100 ;
        RECT 3.240 -0.350 3.500 -0.090 ;
        RECT 1.310 -1.270 1.570 -1.010 ;
        RECT 2.880 -1.270 3.140 -1.010 ;
  END
END sky130_hilas_Tgate4Single01

MACRO sky130_hilas_VinjDecode2to4
  CLASS BLOCK ;
  FOREIGN sky130_hilas_VinjDecode2to4 ;
  ORIGIN 6.370 -0.540 ;
  SIZE 12.950 BY 6.160 ;
  PIN OUTPUT00
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 3.200 5.550 3.570 5.630 ;
        RECT 3.200 5.540 4.230 5.550 ;
        RECT 6.110 5.540 6.420 5.700 ;
        RECT 3.200 5.370 6.580 5.540 ;
    END
  END OUTPUT00
  PIN OUTPUT01
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 3.200 4.040 3.570 4.120 ;
        RECT 3.200 4.030 4.230 4.040 ;
        RECT 6.110 4.030 6.420 4.190 ;
        RECT 3.200 3.860 6.580 4.030 ;
    END
  END OUTPUT01
  PIN OUTPUT10
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 3.200 2.530 3.570 2.610 ;
        RECT 3.200 2.520 4.230 2.530 ;
        RECT 6.110 2.520 6.420 2.680 ;
        RECT 3.200 2.350 6.580 2.520 ;
    END
  END OUTPUT10
  PIN OUTPUT11
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 3.200 1.030 3.570 1.110 ;
        RECT 3.200 1.020 4.230 1.030 ;
        RECT 6.110 1.020 6.420 1.180 ;
        RECT 3.200 0.850 6.580 1.020 ;
    END
  END OUTPUT11
  PIN VGND
    ANTENNADIFFAREA 1.564800 ;
    PORT
      LAYER met1 ;
        RECT 5.290 0.630 5.560 6.670 ;
    END
    PORT
      LAYER met1 ;
        RECT -3.190 2.130 -2.960 6.660 ;
    END
  END VGND
  PIN VINJ
    ANTENNADIFFAREA 0.914000 ;
    PORT
      LAYER nwell ;
        RECT -0.290 0.540 3.150 6.700 ;
      LAYER met1 ;
        RECT 0.320 6.320 0.540 6.660 ;
        RECT 0.320 6.060 0.550 6.320 ;
        RECT 0.320 5.660 0.540 6.060 ;
        RECT 0.320 5.350 0.570 5.660 ;
        RECT 0.320 4.810 0.540 5.350 ;
        RECT 0.320 4.550 0.550 4.810 ;
        RECT 0.320 4.150 0.540 4.550 ;
        RECT 0.320 3.840 0.570 4.150 ;
        RECT 0.320 3.300 0.540 3.840 ;
        RECT 0.320 3.040 0.550 3.300 ;
        RECT 0.320 2.640 0.540 3.040 ;
        RECT 0.320 2.330 0.570 2.640 ;
        RECT 0.320 1.800 0.540 2.330 ;
        RECT 0.320 1.540 0.550 1.800 ;
        RECT 0.320 1.140 0.540 1.540 ;
        RECT 0.320 0.830 0.570 1.140 ;
        RECT 0.320 0.630 0.540 0.830 ;
    END
    PORT
      LAYER nwell ;
        RECT -6.370 2.040 -4.390 6.700 ;
      LAYER met1 ;
        RECT -5.760 6.320 -5.540 6.660 ;
        RECT -5.760 6.060 -5.530 6.320 ;
        RECT -5.760 5.660 -5.540 6.060 ;
        RECT -5.760 5.350 -5.510 5.660 ;
        RECT -5.760 4.810 -5.540 5.350 ;
        RECT -5.760 4.550 -5.530 4.810 ;
        RECT -5.760 4.150 -5.540 4.550 ;
        RECT -5.760 3.840 -5.510 4.150 ;
        RECT -5.760 3.300 -5.540 3.840 ;
        RECT -5.760 3.040 -5.530 3.300 ;
        RECT -5.760 2.640 -5.540 3.040 ;
        RECT -5.760 2.330 -5.510 2.640 ;
        RECT -5.760 2.130 -5.540 2.330 ;
    END
  END VINJ
  PIN IN2
    ANTENNAGATEAREA 0.642800 ;
    PORT
      LAYER met2 ;
        RECT -1.810 6.060 -1.480 6.120 ;
        RECT 2.340 6.080 2.670 6.160 ;
        RECT 2.070 6.060 2.670 6.080 ;
        RECT -1.810 5.900 2.670 6.060 ;
        RECT -1.810 5.850 -1.480 5.900 ;
        RECT -6.370 4.740 -1.580 4.760 ;
        RECT -6.370 4.580 -1.530 4.740 ;
        RECT -1.800 4.550 -1.530 4.580 ;
        RECT -1.800 4.410 -1.520 4.550 ;
        RECT -1.750 4.390 -1.520 4.410 ;
        RECT -1.830 3.040 -1.500 3.100 ;
        RECT 2.340 3.060 2.670 3.140 ;
        RECT 2.070 3.040 2.670 3.060 ;
        RECT -1.830 2.880 2.670 3.040 ;
        RECT -1.830 2.830 -1.500 2.880 ;
    END
  END IN2
  PIN IN1
    ANTENNAGATEAREA 0.673600 ;
    PORT
      LAYER met2 ;
        RECT -2.660 6.500 3.740 6.510 ;
        RECT -2.680 6.350 3.740 6.500 ;
        RECT -2.680 6.340 -2.410 6.350 ;
        RECT -2.710 6.270 -2.410 6.340 ;
        RECT -6.370 6.090 -2.410 6.270 ;
        RECT 3.320 6.120 3.740 6.350 ;
        RECT -2.710 6.010 -2.440 6.090 ;
        RECT -2.740 5.170 -2.410 5.230 ;
        RECT -2.740 5.010 -1.100 5.170 ;
        RECT -2.740 4.960 -2.410 5.010 ;
        RECT -1.260 5.000 -1.100 5.010 ;
        RECT -1.260 4.840 3.740 5.000 ;
        RECT 3.320 4.610 3.740 4.840 ;
    END
  END IN1
  PIN ENABLE
    PORT
      LAYER met2 ;
        RECT -6.370 3.070 -2.760 3.250 ;
    END
  END ENABLE
  OBS
      LAYER li1 ;
        RECT -5.750 6.270 -5.580 6.410 ;
        RECT 0.330 6.270 0.500 6.410 ;
        RECT 1.060 6.290 1.230 6.370 ;
        RECT 1.870 6.290 2.040 6.370 ;
        RECT 3.410 6.330 3.580 6.450 ;
        RECT -5.750 6.100 -5.560 6.270 ;
        RECT -5.750 6.000 -5.580 6.100 ;
        RECT -6.180 5.620 -6.010 5.720 ;
        RECT -6.200 5.450 -6.010 5.620 ;
        RECT -6.180 5.390 -6.010 5.450 ;
        RECT -5.760 5.660 -5.590 5.720 ;
        RECT -5.760 5.390 -5.510 5.660 ;
        RECT -5.020 5.640 -4.770 5.720 ;
        RECT -5.020 5.470 -3.720 5.640 ;
        RECT -3.160 5.630 -2.990 6.260 ;
        RECT 0.330 6.100 0.520 6.270 ;
        RECT 0.330 6.000 0.500 6.100 ;
        RECT 1.060 5.720 1.270 6.290 ;
        RECT 1.830 6.040 2.040 6.290 ;
        RECT 2.430 6.110 2.600 6.210 ;
        RECT 3.370 6.160 3.580 6.330 ;
        RECT 5.300 6.260 5.560 6.330 ;
        RECT 6.100 6.260 6.280 6.390 ;
        RECT 3.410 6.120 3.580 6.160 ;
        RECT 1.830 5.720 2.000 6.040 ;
        RECT 2.400 5.940 2.600 6.110 ;
        RECT 2.430 5.840 2.600 5.940 ;
        RECT 3.970 6.080 4.840 6.250 ;
        RECT 5.300 6.080 6.280 6.260 ;
        RECT -5.750 5.370 -5.510 5.390 ;
        RECT -4.940 5.380 -4.770 5.470 ;
        RECT -3.240 5.460 -2.910 5.630 ;
        RECT -0.100 5.620 0.070 5.720 ;
        RECT -0.120 5.450 0.070 5.620 ;
        RECT -0.100 5.390 0.070 5.450 ;
        RECT 0.320 5.660 0.490 5.720 ;
        RECT 0.320 5.390 0.570 5.660 ;
        RECT 1.060 5.470 1.310 5.720 ;
        RECT 0.330 5.370 0.570 5.390 ;
        RECT 1.140 5.380 1.310 5.470 ;
        RECT 1.790 5.470 2.000 5.720 ;
        RECT 3.970 5.640 4.140 6.080 ;
        RECT 5.300 5.640 5.560 6.080 ;
        RECT 6.100 5.970 6.280 6.080 ;
        RECT 2.510 5.470 4.140 5.640 ;
        RECT 4.590 5.470 5.560 5.640 ;
        RECT 6.010 5.470 6.350 5.640 ;
        RECT 1.790 5.390 1.960 5.470 ;
        RECT 3.280 5.430 3.450 5.470 ;
        RECT -5.750 4.760 -5.580 4.900 ;
        RECT 0.330 4.760 0.500 4.900 ;
        RECT 1.060 4.780 1.230 4.860 ;
        RECT 1.870 4.780 2.040 4.860 ;
        RECT 3.410 4.820 3.580 4.940 ;
        RECT -5.750 4.590 -5.560 4.760 ;
        RECT -5.750 4.490 -5.580 4.590 ;
        RECT -6.180 4.110 -6.010 4.210 ;
        RECT -6.200 3.940 -6.010 4.110 ;
        RECT -6.180 3.880 -6.010 3.940 ;
        RECT -5.760 4.150 -5.590 4.210 ;
        RECT -5.760 3.880 -5.510 4.150 ;
        RECT -5.020 4.130 -4.770 4.210 ;
        RECT -5.020 3.960 -3.720 4.130 ;
        RECT -3.160 4.120 -2.990 4.750 ;
        RECT 0.330 4.590 0.520 4.760 ;
        RECT 0.330 4.490 0.500 4.590 ;
        RECT 1.060 4.210 1.270 4.780 ;
        RECT 1.830 4.530 2.040 4.780 ;
        RECT 2.430 4.600 2.600 4.700 ;
        RECT 3.370 4.650 3.580 4.820 ;
        RECT 5.300 4.750 5.560 4.820 ;
        RECT 6.100 4.750 6.280 4.880 ;
        RECT 3.410 4.610 3.580 4.650 ;
        RECT 1.830 4.210 2.000 4.530 ;
        RECT 2.400 4.430 2.600 4.600 ;
        RECT 2.430 4.330 2.600 4.430 ;
        RECT 3.970 4.570 4.840 4.740 ;
        RECT 5.300 4.570 6.280 4.750 ;
        RECT -5.750 3.860 -5.510 3.880 ;
        RECT -4.940 3.870 -4.770 3.960 ;
        RECT -3.240 3.950 -2.910 4.120 ;
        RECT -0.100 4.110 0.070 4.210 ;
        RECT -0.120 3.940 0.070 4.110 ;
        RECT -0.100 3.880 0.070 3.940 ;
        RECT 0.320 4.150 0.490 4.210 ;
        RECT 0.320 3.880 0.570 4.150 ;
        RECT 1.060 3.960 1.310 4.210 ;
        RECT 0.330 3.860 0.570 3.880 ;
        RECT 1.140 3.870 1.310 3.960 ;
        RECT 1.790 3.960 2.000 4.210 ;
        RECT 3.970 4.130 4.140 4.570 ;
        RECT 5.300 4.130 5.560 4.570 ;
        RECT 6.100 4.460 6.280 4.570 ;
        RECT 2.510 3.960 4.140 4.130 ;
        RECT 4.590 3.960 5.560 4.130 ;
        RECT 6.010 3.960 6.350 4.130 ;
        RECT 1.790 3.880 1.960 3.960 ;
        RECT 3.280 3.920 3.450 3.960 ;
        RECT -5.750 3.250 -5.580 3.390 ;
        RECT 0.330 3.250 0.500 3.390 ;
        RECT 1.060 3.270 1.230 3.350 ;
        RECT 1.870 3.270 2.040 3.350 ;
        RECT 3.410 3.310 3.580 3.430 ;
        RECT -5.750 3.080 -5.560 3.250 ;
        RECT -5.750 2.980 -5.580 3.080 ;
        RECT -6.180 2.600 -6.010 2.700 ;
        RECT -6.200 2.430 -6.010 2.600 ;
        RECT -6.180 2.370 -6.010 2.430 ;
        RECT -5.760 2.640 -5.590 2.700 ;
        RECT -5.760 2.370 -5.510 2.640 ;
        RECT -5.020 2.620 -4.770 2.700 ;
        RECT -5.020 2.450 -3.720 2.620 ;
        RECT -3.160 2.610 -2.990 3.240 ;
        RECT 0.330 3.080 0.520 3.250 ;
        RECT 0.330 2.980 0.500 3.080 ;
        RECT 1.060 2.700 1.270 3.270 ;
        RECT 1.830 3.020 2.040 3.270 ;
        RECT 2.430 3.090 2.600 3.190 ;
        RECT 3.370 3.140 3.580 3.310 ;
        RECT 5.300 3.240 5.560 3.310 ;
        RECT 6.100 3.240 6.280 3.370 ;
        RECT 3.410 3.100 3.580 3.140 ;
        RECT 1.830 2.700 2.000 3.020 ;
        RECT 2.400 2.920 2.600 3.090 ;
        RECT 2.430 2.820 2.600 2.920 ;
        RECT 3.970 3.060 4.840 3.230 ;
        RECT 5.300 3.060 6.280 3.240 ;
        RECT -5.750 2.350 -5.510 2.370 ;
        RECT -4.940 2.360 -4.770 2.450 ;
        RECT -3.240 2.440 -2.910 2.610 ;
        RECT -0.100 2.600 0.070 2.700 ;
        RECT -0.120 2.430 0.070 2.600 ;
        RECT -0.100 2.370 0.070 2.430 ;
        RECT 0.320 2.640 0.490 2.700 ;
        RECT 0.320 2.370 0.570 2.640 ;
        RECT 1.060 2.450 1.310 2.700 ;
        RECT 0.330 2.350 0.570 2.370 ;
        RECT 1.140 2.360 1.310 2.450 ;
        RECT 1.790 2.450 2.000 2.700 ;
        RECT 3.970 2.620 4.140 3.060 ;
        RECT 5.300 2.620 5.560 3.060 ;
        RECT 6.100 2.950 6.280 3.060 ;
        RECT 2.510 2.450 4.140 2.620 ;
        RECT 4.590 2.450 5.560 2.620 ;
        RECT 6.010 2.450 6.350 2.620 ;
        RECT 1.790 2.370 1.960 2.450 ;
        RECT 3.280 2.410 3.450 2.450 ;
        RECT 0.330 1.750 0.500 1.890 ;
        RECT 1.060 1.770 1.230 1.850 ;
        RECT 1.870 1.770 2.040 1.850 ;
        RECT 3.410 1.810 3.580 1.930 ;
        RECT 0.330 1.580 0.520 1.750 ;
        RECT 0.330 1.480 0.500 1.580 ;
        RECT 1.060 1.200 1.270 1.770 ;
        RECT 1.830 1.520 2.040 1.770 ;
        RECT 2.430 1.590 2.600 1.690 ;
        RECT 3.370 1.640 3.580 1.810 ;
        RECT 5.300 1.740 5.560 1.810 ;
        RECT 6.100 1.740 6.280 1.870 ;
        RECT 3.410 1.600 3.580 1.640 ;
        RECT 1.830 1.200 2.000 1.520 ;
        RECT 2.400 1.420 2.600 1.590 ;
        RECT 2.430 1.320 2.600 1.420 ;
        RECT 3.970 1.560 4.840 1.730 ;
        RECT 5.300 1.560 6.280 1.740 ;
        RECT -0.100 1.100 0.070 1.200 ;
        RECT -0.120 0.930 0.070 1.100 ;
        RECT -0.100 0.870 0.070 0.930 ;
        RECT 0.320 1.140 0.490 1.200 ;
        RECT 0.320 0.870 0.570 1.140 ;
        RECT 1.060 0.950 1.310 1.200 ;
        RECT 0.330 0.850 0.570 0.870 ;
        RECT 1.140 0.860 1.310 0.950 ;
        RECT 1.790 0.950 2.000 1.200 ;
        RECT 3.970 1.120 4.140 1.560 ;
        RECT 5.300 1.120 5.560 1.560 ;
        RECT 6.100 1.450 6.280 1.560 ;
        RECT 2.510 0.950 4.140 1.120 ;
        RECT 4.590 0.950 5.560 1.120 ;
        RECT 6.010 0.950 6.350 1.120 ;
        RECT 1.790 0.870 1.960 0.950 ;
        RECT 3.280 0.910 3.450 0.950 ;
      LAYER mcon ;
        RECT -5.730 6.100 -5.560 6.270 ;
        RECT 0.350 6.100 0.520 6.270 ;
        RECT -3.160 5.740 -2.990 5.910 ;
        RECT -5.720 5.420 -5.550 5.590 ;
        RECT -4.380 5.470 -4.210 5.640 ;
        RECT 0.360 5.420 0.530 5.590 ;
        RECT 5.330 5.760 5.510 5.940 ;
        RECT -5.730 4.590 -5.560 4.760 ;
        RECT 0.350 4.590 0.520 4.760 ;
        RECT -3.160 4.230 -2.990 4.400 ;
        RECT -5.720 3.910 -5.550 4.080 ;
        RECT -4.380 3.960 -4.210 4.130 ;
        RECT 0.360 3.910 0.530 4.080 ;
        RECT 5.330 4.250 5.510 4.430 ;
        RECT -5.730 3.080 -5.560 3.250 ;
        RECT 0.350 3.080 0.520 3.250 ;
        RECT -3.160 2.720 -2.990 2.890 ;
        RECT -5.720 2.400 -5.550 2.570 ;
        RECT -4.380 2.450 -4.210 2.620 ;
        RECT 0.360 2.400 0.530 2.570 ;
        RECT 5.330 2.740 5.510 2.920 ;
        RECT 0.350 1.580 0.520 1.750 ;
        RECT 0.360 0.900 0.530 1.070 ;
        RECT 5.330 1.240 5.510 1.420 ;
      LAYER met1 ;
        RECT -2.700 6.310 -2.430 6.600 ;
        RECT -2.740 6.040 -2.410 6.310 ;
        RECT -6.290 5.380 -5.980 5.730 ;
        RECT -4.460 5.420 -4.140 5.680 ;
        RECT -2.700 5.260 -2.430 6.040 ;
        RECT -2.710 4.930 -2.430 5.260 ;
        RECT -2.700 4.900 -2.430 4.930 ;
        RECT -6.290 3.870 -5.980 4.220 ;
        RECT -4.460 3.910 -4.140 4.170 ;
        RECT -2.240 3.580 -1.970 5.700 ;
        RECT -1.780 4.710 -1.510 6.170 ;
        RECT 2.340 5.900 2.670 6.160 ;
        RECT 3.310 6.120 3.740 6.410 ;
        RECT -0.830 5.670 -0.540 5.720 ;
        RECT -0.850 5.320 -0.540 5.670 ;
        RECT -0.210 5.380 0.100 5.730 ;
        RECT 3.180 5.370 3.570 5.640 ;
        RECT 6.110 5.380 6.420 5.700 ;
        RECT -1.830 4.440 -1.500 4.710 ;
        RECT -2.250 3.250 -1.970 3.580 ;
        RECT -6.290 2.360 -5.980 2.710 ;
        RECT -4.460 2.400 -4.140 2.660 ;
        RECT -2.240 2.080 -1.970 3.250 ;
        RECT -1.780 3.130 -1.510 4.440 ;
        RECT -1.800 2.800 -1.510 3.130 ;
        RECT -1.780 2.780 -1.510 2.800 ;
        RECT -1.310 4.170 -1.040 4.230 ;
        RECT -1.310 3.840 -1.030 4.170 ;
        RECT -2.240 1.750 -1.940 2.080 ;
        RECT -2.240 1.700 -1.970 1.750 ;
        RECT -1.310 1.630 -1.040 3.840 ;
        RECT -1.330 1.300 -1.040 1.630 ;
        RECT -1.310 1.270 -1.040 1.300 ;
        RECT -0.830 2.670 -0.540 5.320 ;
        RECT 2.340 4.390 2.670 4.650 ;
        RECT 3.310 4.610 3.740 4.900 ;
        RECT -0.210 3.870 0.100 4.220 ;
        RECT 3.180 3.860 3.570 4.130 ;
        RECT 6.110 3.870 6.420 4.190 ;
        RECT 2.340 2.880 2.670 3.140 ;
        RECT 3.310 3.100 3.740 3.390 ;
        RECT -0.830 2.320 -0.530 2.670 ;
        RECT -0.210 2.360 0.100 2.710 ;
        RECT 3.180 2.350 3.570 2.620 ;
        RECT 6.110 2.360 6.420 2.680 ;
        RECT -0.830 0.780 -0.540 2.320 ;
        RECT 2.340 1.380 2.670 1.640 ;
        RECT 3.310 1.600 3.740 1.890 ;
        RECT -0.210 0.860 0.100 1.210 ;
        RECT 3.180 0.850 3.570 1.120 ;
        RECT 6.110 0.860 6.420 1.180 ;
      LAYER via ;
        RECT -2.710 6.040 -2.440 6.310 ;
        RECT -6.260 5.410 -6.000 5.670 ;
        RECT -4.430 5.420 -4.170 5.680 ;
        RECT -1.780 5.850 -1.510 6.120 ;
        RECT 2.380 5.900 2.640 6.160 ;
        RECT 3.370 6.150 3.630 6.410 ;
        RECT -2.710 4.960 -2.440 5.230 ;
        RECT -2.240 5.360 -1.970 5.630 ;
        RECT -6.260 3.900 -6.000 4.160 ;
        RECT -4.430 3.910 -4.170 4.170 ;
        RECT -0.850 5.350 -0.560 5.640 ;
        RECT -0.180 5.410 0.080 5.670 ;
        RECT 3.240 5.370 3.500 5.630 ;
        RECT 6.140 5.410 6.400 5.670 ;
        RECT -1.800 4.440 -1.530 4.710 ;
        RECT -2.250 3.280 -1.980 3.550 ;
        RECT -6.260 2.390 -6.000 2.650 ;
        RECT -4.430 2.400 -4.170 2.660 ;
        RECT -1.800 2.830 -1.530 3.100 ;
        RECT -1.300 3.870 -1.030 4.140 ;
        RECT 2.380 4.390 2.640 4.650 ;
        RECT 3.370 4.640 3.630 4.900 ;
        RECT -0.810 3.840 -0.550 4.100 ;
        RECT -0.180 3.900 0.080 4.160 ;
        RECT 3.240 3.860 3.500 4.120 ;
        RECT 6.140 3.900 6.400 4.160 ;
        RECT -2.210 1.780 -1.940 2.050 ;
        RECT -1.330 1.330 -1.060 1.600 ;
        RECT 2.380 2.880 2.640 3.140 ;
        RECT 3.370 3.130 3.630 3.390 ;
        RECT -0.820 2.350 -0.530 2.640 ;
        RECT -0.180 2.390 0.080 2.650 ;
        RECT 3.240 2.350 3.500 2.610 ;
        RECT 6.140 2.390 6.400 2.650 ;
        RECT 2.380 1.380 2.640 1.640 ;
        RECT 3.370 1.630 3.630 1.890 ;
        RECT -0.830 0.810 -0.540 1.100 ;
        RECT -0.180 0.890 0.080 1.150 ;
        RECT 3.240 0.850 3.500 1.110 ;
        RECT 6.140 0.890 6.400 1.150 ;
      LAYER met2 ;
        RECT -6.290 5.570 -5.970 5.670 ;
        RECT -6.300 5.410 -5.970 5.570 ;
        RECT -4.460 5.600 -4.140 5.680 ;
        RECT -2.270 5.600 -1.940 5.630 ;
        RECT -4.460 5.420 -1.920 5.600 ;
        RECT -2.270 5.410 -1.920 5.420 ;
        RECT -0.880 5.570 -0.530 5.640 ;
        RECT -0.210 5.570 0.110 5.670 ;
        RECT -0.880 5.410 0.110 5.570 ;
        RECT -2.270 5.360 -1.940 5.410 ;
        RECT -0.880 5.350 -0.530 5.410 ;
        RECT 2.340 4.570 2.670 4.650 ;
        RECT 2.070 4.550 2.670 4.570 ;
        RECT -1.250 4.390 2.670 4.550 ;
        RECT -6.290 4.060 -5.970 4.160 ;
        RECT -6.300 3.900 -5.970 4.060 ;
        RECT -4.460 4.090 -4.140 4.170 ;
        RECT -1.250 4.140 -1.090 4.390 ;
        RECT -1.330 4.090 -1.000 4.140 ;
        RECT -4.460 3.910 -1.000 4.090 ;
        RECT -1.330 3.870 -1.000 3.910 ;
        RECT -0.840 4.060 -0.520 4.100 ;
        RECT -0.210 4.060 0.110 4.160 ;
        RECT -0.840 3.900 0.110 4.060 ;
        RECT -0.840 3.840 -0.520 3.900 ;
        RECT -2.280 3.490 -1.950 3.550 ;
        RECT -2.280 3.330 3.740 3.490 ;
        RECT -2.280 3.280 -1.950 3.330 ;
        RECT 3.320 3.100 3.740 3.330 ;
        RECT -6.290 2.550 -5.970 2.650 ;
        RECT -6.300 2.390 -5.970 2.550 ;
        RECT -4.460 2.580 -4.140 2.660 ;
        RECT -0.850 2.580 -0.500 2.640 ;
        RECT -4.460 2.550 -0.360 2.580 ;
        RECT -0.210 2.550 0.110 2.650 ;
        RECT -4.460 2.400 0.110 2.550 ;
        RECT -0.850 2.390 0.110 2.400 ;
        RECT -0.850 2.350 -0.500 2.390 ;
        RECT -2.240 1.990 -1.910 2.050 ;
        RECT -2.240 1.830 3.740 1.990 ;
        RECT -2.240 1.780 -1.910 1.830 ;
        RECT -1.360 1.540 -1.030 1.600 ;
        RECT 2.340 1.560 2.670 1.640 ;
        RECT 3.320 1.600 3.740 1.830 ;
        RECT 2.070 1.540 2.670 1.560 ;
        RECT -1.360 1.380 2.670 1.540 ;
        RECT -1.360 1.330 -1.030 1.380 ;
        RECT -0.860 1.050 -0.510 1.100 ;
        RECT -0.210 1.050 0.110 1.150 ;
        RECT -0.860 0.890 0.110 1.050 ;
        RECT -0.860 0.810 -0.510 0.890 ;
  END
END sky130_hilas_VinjDecode2to4

MACRO sky130_hilas_TA2Cell_1FG
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TA2Cell_1FG ;
  ORIGIN 30.130 -1.400 ;
  SIZE 32.060 BY 9.870 ;
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -17.310 2.650 -16.830 2.660 ;
        RECT -17.310 2.410 -16.420 2.650 ;
    END
  END VIN12
  PIN VIN11
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -17.260 6.170 -16.420 6.370 ;
    END
  END VIN11
  PIN VIN21
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -2.200 4.750 -1.890 4.790 ;
        RECT -2.520 4.740 -1.860 4.750 ;
        RECT -2.520 4.510 -1.420 4.740 ;
        RECT -2.200 4.460 -1.890 4.510 ;
    END
  END VIN21
  PIN VIN22
    USE ANALOG ;
    ANTENNAGATEAREA 4.342100 ;
    ANTENNADIFFAREA 8.158800 ;
    PORT
      LAYER nwell ;
        RECT -2.550 7.450 0.760 11.270 ;
        RECT -3.200 7.440 1.930 7.450 ;
        RECT -3.210 5.230 1.930 7.440 ;
        RECT -3.210 1.400 -1.350 5.230 ;
        RECT 0.650 1.400 1.930 5.230 ;
      LAYER met2 ;
        RECT -0.630 8.410 -0.310 8.670 ;
        RECT -0.590 8.390 0.590 8.410 ;
        RECT -0.590 8.130 0.630 8.390 ;
        RECT -0.590 8.070 0.590 8.130 ;
        RECT -0.630 8.060 0.590 8.070 ;
        RECT -0.630 7.810 -0.310 8.060 ;
        RECT -1.960 7.430 -1.650 7.440 ;
        RECT -2.530 7.420 -1.650 7.430 ;
        RECT -2.600 7.180 -1.650 7.420 ;
        RECT -1.960 7.110 -1.650 7.180 ;
        RECT -0.990 7.110 -0.680 7.160 ;
        RECT 1.260 7.110 1.570 7.210 ;
        RECT -1.570 6.990 -1.260 7.060 ;
        RECT -0.990 6.990 1.570 7.110 ;
        RECT -1.570 6.880 1.570 6.990 ;
        RECT -1.570 6.780 0.760 6.880 ;
        RECT -1.570 6.730 -1.260 6.780 ;
        RECT -1.810 6.570 -1.500 6.610 ;
        RECT -1.990 6.430 -1.270 6.570 ;
        RECT -1.040 6.430 -0.730 6.510 ;
        RECT -1.990 6.320 -0.730 6.430 ;
        RECT -1.810 6.280 -0.730 6.320 ;
        RECT -1.540 6.220 -0.730 6.280 ;
        RECT -1.540 6.210 -1.270 6.220 ;
        RECT -1.040 6.180 -0.730 6.220 ;
        RECT -2.930 5.930 -2.620 6.070 ;
        RECT -16.810 5.890 -6.670 5.920 ;
        RECT -3.280 5.890 -2.620 5.930 ;
        RECT -1.720 5.900 -1.410 6.040 ;
        RECT -1.720 5.890 0.760 5.900 ;
        RECT -16.810 5.740 0.760 5.890 ;
        RECT -16.810 5.700 -6.670 5.740 ;
        RECT -3.280 5.710 -2.930 5.740 ;
        RECT -1.720 5.720 0.760 5.740 ;
        RECT -1.720 5.710 -1.410 5.720 ;
        RECT -6.890 4.500 -6.670 5.700 ;
        RECT -1.470 5.640 -1.270 5.650 ;
        RECT -1.470 5.630 -1.250 5.640 ;
        RECT -1.040 5.630 -0.730 5.670 ;
        RECT -1.470 5.560 -0.730 5.630 ;
        RECT -1.760 5.540 -0.730 5.560 ;
        RECT -1.810 5.420 -0.730 5.540 ;
        RECT -1.810 5.300 -1.250 5.420 ;
        RECT -1.040 5.340 -0.730 5.420 ;
        RECT -1.810 5.290 -1.340 5.300 ;
        RECT -6.920 4.460 -6.670 4.500 ;
        RECT -6.920 3.820 -6.660 4.460 ;
        RECT -6.920 3.610 -2.790 3.820 ;
        RECT -3.000 3.470 -2.790 3.610 ;
        RECT -1.040 3.470 -0.730 3.550 ;
        RECT -3.000 3.260 -0.730 3.470 ;
        RECT -1.040 3.220 -0.730 3.260 ;
        RECT -11.980 1.750 -11.660 1.760 ;
        RECT -1.540 1.750 -1.210 1.890 ;
        RECT -11.980 1.590 -1.210 1.750 ;
        RECT -11.980 1.580 -11.290 1.590 ;
        RECT -11.980 1.460 -11.660 1.580 ;
    END
  END VIN22
  PIN VPWR
    USE ANALOG ;
    ANTENNADIFFAREA 1.373600 ;
    PORT
      LAYER met1 ;
        RECT 0.630 7.300 0.910 7.450 ;
        RECT 0.640 5.870 0.910 7.300 ;
        RECT 0.640 5.580 0.920 5.870 ;
        RECT 0.640 3.280 0.910 5.580 ;
        RECT 0.640 2.990 0.920 3.280 ;
        RECT 0.640 1.400 0.910 2.990 ;
    END
  END VPWR
  PIN VGND
    USE ANALOG ;
    ANTENNAGATEAREA 3.745100 ;
    ANTENNADIFFAREA 3.678400 ;
    PORT
      LAYER met1 ;
        RECT -0.200 9.810 -0.010 11.270 ;
        RECT 0.240 10.620 0.520 11.270 ;
        RECT 0.130 10.020 0.520 10.620 ;
        RECT -0.200 9.780 0.020 9.810 ;
        RECT -0.220 9.510 0.030 9.780 ;
        RECT -0.210 9.500 0.030 9.510 ;
        RECT -0.210 9.260 0.020 9.500 ;
        RECT -0.600 7.780 -0.340 8.100 ;
        RECT -0.600 7.660 -0.360 7.780 ;
        RECT -0.170 7.450 -0.010 9.260 ;
        RECT 0.240 8.420 0.520 10.020 ;
        RECT 0.240 8.100 0.600 8.420 ;
        RECT 0.240 7.450 0.520 8.100 ;
        RECT -1.970 7.110 -1.650 7.430 ;
        RECT -0.170 7.230 0.520 7.450 ;
        RECT -0.990 6.830 -0.670 7.150 ;
        RECT -0.210 6.980 0.520 7.230 ;
        RECT -0.220 6.710 0.520 6.980 ;
        RECT -1.040 6.180 -0.720 6.500 ;
        RECT -1.720 5.600 -1.410 6.040 ;
        RECT -1.710 5.590 -1.500 5.600 ;
        RECT -1.730 5.270 -1.470 5.590 ;
        RECT -1.040 5.350 -0.720 5.670 ;
        RECT -1.710 3.980 -1.500 5.270 ;
        RECT -0.200 5.220 0.520 6.710 ;
        RECT -1.730 3.690 -1.500 3.980 ;
        RECT -1.540 1.600 -1.210 1.890 ;
        RECT -0.030 1.600 0.310 5.220 ;
        RECT -1.550 1.460 0.310 1.600 ;
        RECT -0.030 1.400 0.310 1.460 ;
      LAYER via ;
        RECT -0.600 7.810 -0.340 8.070 ;
        RECT 0.340 8.130 0.600 8.390 ;
        RECT -1.940 7.140 -1.680 7.400 ;
        RECT -0.960 6.860 -0.700 7.120 ;
        RECT -1.010 6.210 -0.750 6.470 ;
        RECT -1.690 5.750 -1.430 6.010 ;
        RECT -1.730 5.300 -1.470 5.560 ;
        RECT -1.010 5.380 -0.750 5.640 ;
        RECT -1.510 1.610 -1.240 1.870 ;
    END
    PORT
      LAYER met1 ;
        RECT -17.690 7.360 -17.460 7.440 ;
    END
    PORT
      LAYER met1 ;
        RECT -11.900 7.360 -11.670 7.450 ;
    END
  END VGND
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT -25.920 7.280 -25.600 7.400 ;
        RECT -3.720 7.280 -3.400 7.400 ;
        RECT -25.920 7.100 -3.400 7.280 ;
    END
    PORT
      LAYER met1 ;
        RECT -3.720 1.400 -3.440 1.450 ;
    END
    PORT
      LAYER met1 ;
        RECT -25.920 7.400 -25.640 7.450 ;
        RECT -25.920 7.120 -25.600 7.400 ;
      LAYER via ;
        RECT -25.890 7.130 -25.630 7.390 ;
    END
  END VINJ
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER met2 ;
        RECT -0.990 4.970 -0.680 5.020 ;
        RECT 1.310 4.970 1.620 4.990 ;
        RECT -0.990 4.740 1.930 4.970 ;
        RECT -0.990 4.690 -0.680 4.740 ;
        RECT 1.310 4.660 1.620 4.740 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER met2 ;
        RECT -0.990 4.140 -0.680 4.200 ;
        RECT 1.300 4.140 1.610 4.270 ;
        RECT -0.990 3.920 1.930 4.140 ;
        RECT -0.990 3.870 -0.680 3.920 ;
    END
  END OUTPUT2
  PIN DRAIN1
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT -28.110 6.990 -27.800 7.060 ;
        RECT -30.130 6.780 -18.600 6.990 ;
        RECT -28.820 6.770 -18.600 6.780 ;
        RECT -28.110 6.730 -27.800 6.770 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT -26.160 1.900 -26.080 2.080 ;
    END
  END DRAIN2
  PIN COLSEL2
    PORT
      LAYER met1 ;
        RECT -25.390 7.390 -25.200 7.450 ;
    END
  END COLSEL2
  PIN GATE2
    PORT
      LAYER met1 ;
        RECT -18.910 7.360 -18.680 7.440 ;
    END
  END GATE2
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT -10.680 7.370 -10.450 7.450 ;
    END
  END GATE1
  PIN COLSEL1
    PORT
      LAYER met1 ;
        RECT -4.160 7.370 -3.970 7.450 ;
    END
    PORT
      LAYER met1 ;
        RECT -4.160 1.400 -3.970 1.450 ;
    END
  END COLSEL1
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT -15.400 7.290 -13.960 7.450 ;
    END
  END VTUN
  OBS
      LAYER nwell ;
        RECT -30.130 5.230 -26.820 11.260 ;
        RECT -25.090 8.880 -22.370 10.530 ;
        RECT -20.340 10.520 -18.610 11.270 ;
        RECT -25.080 8.840 -22.370 8.880 ;
        RECT -25.080 7.510 -22.370 7.550 ;
        RECT -25.090 7.450 -22.370 7.510 ;
        RECT -26.160 7.440 -22.370 7.450 ;
        RECT -26.160 6.770 -26.090 6.950 ;
        RECT -25.090 5.860 -22.370 7.440 ;
        RECT -20.350 6.950 -18.610 10.520 ;
        RECT -20.340 5.230 -18.610 6.950 ;
        RECT -10.760 10.520 -9.030 11.270 ;
        RECT -10.760 6.950 -9.020 10.520 ;
        RECT -7.000 8.880 -4.280 10.530 ;
        RECT -7.000 8.840 -4.290 8.880 ;
        RECT -7.000 7.510 -4.290 7.550 ;
        RECT -10.760 5.230 -9.030 6.950 ;
        RECT -7.000 5.860 -4.280 7.510 ;
        RECT -26.160 1.900 -26.080 2.080 ;
      LAYER li1 ;
        RECT -29.730 10.590 -29.530 10.940 ;
        RECT -28.250 10.690 -27.720 10.860 ;
        RECT -29.740 10.560 -29.530 10.590 ;
        RECT -29.740 9.980 -29.520 10.560 ;
        RECT -29.740 9.970 -29.530 9.980 ;
        RECT -29.360 9.800 -29.170 9.810 ;
        RECT -29.370 9.510 -29.170 9.800 ;
        RECT -29.400 9.180 -29.160 9.510 ;
        RECT -28.970 8.700 -28.800 10.310 ;
        RECT -28.980 8.510 -28.800 8.700 ;
        RECT -28.140 9.780 -27.970 10.300 ;
        RECT -27.550 10.110 -27.220 10.280 ;
        RECT -26.200 10.110 -25.850 10.280 ;
        RECT -25.530 10.260 -20.470 11.090 ;
        RECT -1.650 10.690 -1.120 10.860 ;
        RECT 0.160 10.590 0.360 10.940 ;
        RECT 0.160 10.560 0.370 10.590 ;
        RECT -21.020 10.180 -20.540 10.260 ;
        RECT -28.140 9.520 -27.810 9.780 ;
        RECT -28.140 8.610 -27.970 9.520 ;
        RECT -27.550 9.320 -27.220 9.490 ;
        RECT -26.200 9.320 -25.850 9.490 ;
        RECT -22.900 9.320 -22.670 10.010 ;
        RECT -21.020 9.930 -20.550 10.180 ;
        RECT -3.520 10.110 -3.170 10.280 ;
        RECT -2.150 10.110 -1.820 10.280 ;
        RECT -19.590 9.130 -19.040 9.560 ;
        RECT -10.330 9.130 -9.780 9.560 ;
        RECT -6.700 9.320 -6.470 10.010 ;
        RECT -1.400 9.780 -1.230 10.300 ;
        RECT -1.560 9.520 -1.230 9.780 ;
        RECT -3.520 9.320 -3.170 9.490 ;
        RECT -2.150 9.320 -1.820 9.490 ;
        RECT -27.550 8.530 -27.220 8.700 ;
        RECT -26.200 8.530 -25.860 8.700 ;
        RECT -28.980 7.790 -28.800 7.980 ;
        RECT -27.470 7.960 -27.300 8.530 ;
        RECT -21.830 8.300 -21.640 8.700 ;
        RECT -7.730 8.300 -7.540 8.700 ;
        RECT -3.510 8.530 -3.170 8.700 ;
        RECT -2.150 8.530 -1.820 8.700 ;
        RECT -1.400 8.610 -1.230 9.520 ;
        RECT -0.570 8.700 -0.400 10.310 ;
        RECT 0.150 9.980 0.370 10.560 ;
        RECT 0.160 9.970 0.370 9.980 ;
        RECT -0.200 9.800 -0.010 9.810 ;
        RECT -0.200 9.510 0.000 9.800 ;
        RECT -0.210 9.180 0.030 9.510 ;
        RECT -21.830 8.290 -21.450 8.300 ;
        RECT -25.190 8.110 -21.450 8.290 ;
        RECT -21.830 8.070 -21.450 8.110 ;
        RECT -7.920 8.290 -7.540 8.300 ;
        RECT -7.920 8.110 -4.180 8.290 ;
        RECT -7.920 8.070 -7.540 8.110 ;
        RECT -29.400 6.980 -29.160 7.310 ;
        RECT -29.370 6.690 -29.170 6.980 ;
        RECT -29.360 6.680 -29.170 6.690 ;
        RECT -29.740 6.510 -29.530 6.520 ;
        RECT -29.740 5.930 -29.520 6.510 ;
        RECT -28.970 6.180 -28.800 7.790 ;
        RECT -28.140 7.020 -27.970 7.880 ;
        RECT -27.550 7.790 -27.220 7.960 ;
        RECT -26.200 7.790 -25.860 7.960 ;
        RECT -21.830 7.690 -21.640 8.070 ;
        RECT -19.590 7.400 -19.040 7.830 ;
        RECT -10.330 7.400 -9.780 7.830 ;
        RECT -7.730 7.690 -7.540 8.070 ;
        RECT -2.070 7.960 -1.900 8.530 ;
        RECT -0.570 8.510 -0.390 8.700 ;
        RECT -3.510 7.790 -3.170 7.960 ;
        RECT -2.150 7.790 -1.820 7.960 ;
        RECT -2.220 7.400 -2.050 7.450 ;
        RECT -28.140 6.760 -27.810 7.020 ;
        RECT -27.550 7.000 -27.220 7.170 ;
        RECT -26.200 7.000 -25.850 7.170 ;
        RECT -28.140 6.190 -27.970 6.760 ;
        RECT -22.900 6.380 -22.670 7.110 ;
        RECT -27.550 6.210 -27.220 6.380 ;
        RECT -26.200 6.210 -25.850 6.380 ;
        RECT -20.860 6.250 -20.520 6.500 ;
        RECT -6.700 6.380 -6.470 7.110 ;
        RECT -3.520 7.000 -3.170 7.170 ;
        RECT -2.220 7.140 -1.660 7.400 ;
        RECT -2.220 7.120 -1.820 7.140 ;
        RECT -2.150 7.000 -1.820 7.120 ;
        RECT -1.400 7.020 -1.230 7.880 ;
        RECT -0.570 7.790 -0.390 7.980 ;
        RECT -0.570 7.160 -0.400 7.790 ;
        RECT -0.750 7.120 -0.400 7.160 ;
        RECT -20.860 6.170 -20.510 6.250 ;
        RECT -3.520 6.210 -3.170 6.380 ;
        RECT -29.740 5.900 -29.530 5.930 ;
        RECT -29.730 5.550 -29.530 5.900 ;
        RECT -28.250 5.630 -27.720 5.800 ;
        RECT -25.560 5.320 -20.510 6.170 ;
        RECT -2.800 6.040 -2.620 6.970 ;
        RECT -2.070 6.710 -1.740 6.880 ;
        RECT -1.560 6.760 -1.230 7.020 ;
        RECT -0.980 6.860 -0.400 7.120 ;
        RECT -0.210 7.160 0.030 7.310 ;
        RECT -0.210 6.980 0.390 7.160 ;
        RECT -0.750 6.830 -0.400 6.860 ;
        RECT -1.990 6.570 -1.740 6.710 ;
        RECT -1.990 6.380 -1.510 6.570 ;
        RECT -2.150 6.310 -1.510 6.380 ;
        RECT -2.150 6.210 -1.820 6.310 ;
        RECT -2.920 6.010 -2.600 6.040 ;
        RECT -2.920 5.820 -2.590 6.010 ;
        RECT -2.920 5.780 -2.600 5.820 ;
        RECT -17.670 3.870 -17.470 4.880 ;
        RECT -11.920 3.870 -11.630 4.880 ;
        RECT -2.800 1.870 -2.620 5.780 ;
        RECT -1.990 4.930 -1.820 6.210 ;
        RECT -1.400 6.190 -1.230 6.760 ;
        RECT -1.160 6.470 -0.990 6.510 ;
        RECT -0.570 6.500 -0.400 6.830 ;
        RECT -0.200 6.680 0.390 6.980 ;
        RECT 1.210 7.040 1.790 7.210 ;
        RECT 1.210 6.940 1.600 7.040 ;
        RECT 1.210 6.910 1.590 6.940 ;
        RECT 1.210 6.760 1.570 6.910 ;
        RECT -0.750 6.470 -0.400 6.500 ;
        RECT -1.160 6.210 -0.400 6.470 ;
        RECT -1.160 6.180 -0.990 6.210 ;
        RECT -0.750 6.180 -0.400 6.210 ;
        RECT -0.750 6.170 -0.550 6.180 ;
        RECT -0.160 6.170 0.390 6.680 ;
        RECT 0.860 6.590 1.570 6.760 ;
        RECT 0.150 5.930 0.370 6.170 ;
        RECT 0.160 5.900 0.370 5.930 ;
        RECT -1.650 5.670 -1.120 5.800 ;
        RECT 0.160 5.680 0.360 5.900 ;
        RECT 0.860 5.840 1.560 6.150 ;
        RECT -1.650 5.640 -0.990 5.670 ;
        RECT -0.750 5.640 -0.550 5.680 ;
        RECT -1.650 5.630 -0.550 5.640 ;
        RECT -1.160 5.380 -0.550 5.630 ;
        RECT -1.160 5.340 -0.990 5.380 ;
        RECT -0.750 5.350 -0.550 5.380 ;
        RECT -0.750 4.990 -0.550 5.020 ;
        RECT -2.190 4.730 -1.870 4.760 ;
        RECT -0.980 4.730 -0.550 4.990 ;
        RECT -2.190 4.540 -1.860 4.730 ;
        RECT -0.750 4.690 -0.550 4.730 ;
        RECT -0.160 4.690 0.390 5.680 ;
        RECT 0.710 5.610 1.560 5.840 ;
        RECT 0.860 5.270 1.560 5.610 ;
        RECT 1.320 4.910 1.640 4.950 ;
        RECT 1.320 4.850 1.650 4.910 ;
        RECT 0.850 4.720 1.650 4.850 ;
        RECT 0.850 4.690 1.640 4.720 ;
        RECT 0.850 4.670 1.550 4.690 ;
        RECT -2.190 4.500 -1.870 4.540 ;
        RECT -2.190 4.420 -2.020 4.500 ;
        RECT -2.240 4.250 -2.020 4.420 ;
        RECT -2.240 4.090 -2.070 4.250 ;
        RECT -0.750 4.160 -0.550 4.200 ;
        RECT -1.710 3.830 -1.520 3.950 ;
        RECT -0.980 3.900 -0.550 4.160 ;
        RECT -0.750 3.870 -0.550 3.900 ;
        RECT -2.070 3.720 -1.520 3.830 ;
        RECT -2.070 3.660 -1.530 3.720 ;
        RECT -1.990 1.880 -1.820 3.660 ;
        RECT -1.160 3.510 -0.990 3.550 ;
        RECT -0.750 3.510 -0.550 3.540 ;
        RECT -1.160 3.250 -0.550 3.510 ;
        RECT -1.160 3.220 -0.990 3.250 ;
        RECT -0.750 3.210 -0.550 3.250 ;
        RECT -0.160 3.210 0.390 4.200 ;
        RECT 1.310 4.190 1.630 4.230 ;
        RECT 0.850 4.010 1.640 4.190 ;
        RECT 1.310 4.000 1.640 4.010 ;
        RECT 1.310 3.970 1.630 4.000 ;
        RECT 0.860 3.250 1.560 3.590 ;
        RECT 0.710 3.020 1.560 3.250 ;
        RECT -1.160 2.680 -0.990 2.710 ;
        RECT -0.750 2.680 -0.550 2.720 ;
        RECT -1.160 2.420 -0.550 2.680 ;
        RECT -1.160 2.380 -0.990 2.420 ;
        RECT -0.750 2.390 -0.550 2.420 ;
        RECT -0.750 2.030 -0.550 2.060 ;
        RECT -0.980 1.770 -0.550 2.030 ;
        RECT -0.750 1.730 -0.550 1.770 ;
        RECT -0.160 1.730 0.390 2.720 ;
        RECT 0.860 2.710 1.560 3.020 ;
        RECT 0.860 2.100 1.570 2.270 ;
        RECT 1.210 1.820 1.570 2.100 ;
        RECT 1.210 1.650 1.790 1.820 ;
      LAYER mcon ;
        RECT -27.900 10.690 -27.720 10.860 ;
        RECT -29.710 10.390 -29.540 10.560 ;
        RECT -29.360 9.550 -29.180 9.740 ;
        RECT 0.170 10.390 0.340 10.560 ;
        RECT -22.870 9.810 -22.700 9.980 ;
        RECT -20.780 9.970 -20.610 10.140 ;
        RECT -28.040 9.560 -27.870 9.730 ;
        RECT -6.670 9.810 -6.500 9.980 ;
        RECT -22.870 9.360 -22.700 9.530 ;
        RECT -19.310 9.210 -19.040 9.480 ;
        RECT -10.330 9.210 -10.060 9.480 ;
        RECT -6.670 9.360 -6.500 9.530 ;
        RECT -1.500 9.560 -1.330 9.730 ;
        RECT -0.190 9.550 -0.010 9.740 ;
        RECT -21.630 8.100 -21.460 8.270 ;
        RECT -7.910 8.100 -7.740 8.270 ;
        RECT -29.360 6.750 -29.180 6.940 ;
        RECT -19.310 7.480 -19.040 7.750 ;
        RECT -10.330 7.480 -10.060 7.750 ;
        RECT -1.890 7.180 -1.720 7.350 ;
        RECT -28.040 6.800 -27.870 6.970 ;
        RECT -22.870 6.860 -22.700 7.030 ;
        RECT -22.870 6.410 -22.700 6.580 ;
        RECT -6.670 6.860 -6.500 7.030 ;
        RECT -20.750 6.280 -20.580 6.450 ;
        RECT -6.670 6.410 -6.500 6.580 ;
        RECT -29.710 5.930 -29.540 6.100 ;
        RECT -27.900 5.630 -27.720 5.800 ;
        RECT -1.500 6.800 -1.330 6.970 ;
        RECT -0.920 6.900 -0.750 7.070 ;
        RECT -1.740 6.350 -1.570 6.520 ;
        RECT -2.860 5.830 -2.690 6.000 ;
        RECT -17.660 4.630 -17.490 4.800 ;
        RECT -17.650 3.940 -17.480 4.110 ;
        RECT -11.870 4.630 -11.700 4.800 ;
        RECT -11.870 3.950 -11.700 4.120 ;
        RECT -0.190 6.750 -0.010 6.940 ;
        RECT 1.330 6.950 1.500 7.120 ;
        RECT -0.970 6.250 -0.800 6.420 ;
        RECT 0.060 6.580 0.230 6.750 ;
        RECT 0.170 5.930 0.340 6.100 ;
        RECT -0.970 5.430 -0.800 5.600 ;
        RECT 0.720 5.640 0.890 5.810 ;
        RECT 0.060 5.100 0.230 5.270 ;
        RECT -0.920 4.780 -0.750 4.950 ;
        RECT -2.130 4.550 -1.960 4.720 ;
        RECT 1.380 4.730 1.550 4.900 ;
        RECT -1.700 3.750 -1.530 3.920 ;
        RECT -0.920 3.940 -0.750 4.110 ;
        RECT 1.370 4.010 1.540 4.180 ;
        RECT 0.060 3.620 0.230 3.790 ;
        RECT -0.970 3.290 -0.800 3.460 ;
        RECT 0.720 3.050 0.890 3.220 ;
        RECT -0.970 2.470 -0.800 2.640 ;
        RECT 0.060 2.140 0.230 2.310 ;
        RECT -0.920 1.820 -0.750 1.990 ;
        RECT 1.290 1.760 1.460 1.930 ;
      LAYER met1 ;
        RECT -29.890 10.620 -29.610 11.270 ;
        RECT -29.890 10.020 -29.500 10.620 ;
        RECT -29.890 6.470 -29.610 10.020 ;
        RECT -29.360 9.810 -29.170 11.270 ;
        RECT -27.960 10.450 -27.650 10.890 ;
        RECT -22.880 10.060 -22.650 11.270 ;
        RECT -21.660 10.300 -21.430 11.270 ;
        RECT -29.390 9.780 -29.170 9.810 ;
        RECT -29.400 9.510 -29.150 9.780 ;
        RECT -29.400 9.500 -29.160 9.510 ;
        RECT -29.390 9.260 -29.160 9.500 ;
        RECT -28.120 9.490 -27.800 9.810 ;
        RECT -22.910 9.270 -22.650 10.060 ;
        RECT -21.670 10.050 -21.430 10.300 ;
        RECT -29.360 7.230 -29.200 9.260 ;
        RECT -29.010 8.700 -28.770 8.830 ;
        RECT -29.030 8.380 -28.770 8.700 ;
        RECT -29.030 7.780 -28.770 8.100 ;
        RECT -29.010 7.660 -28.770 7.780 ;
        RECT -29.390 6.990 -29.160 7.230 ;
        RECT -22.880 7.120 -22.650 9.270 ;
        RECT -29.400 6.980 -29.160 6.990 ;
        RECT -29.400 6.710 -29.150 6.980 ;
        RECT -28.120 6.730 -27.800 7.050 ;
        RECT -29.390 6.680 -29.170 6.710 ;
        RECT -29.890 5.870 -29.500 6.470 ;
        RECT -29.890 5.220 -29.610 5.870 ;
        RECT -29.360 5.220 -29.170 6.680 ;
        RECT -22.910 6.330 -22.650 7.120 ;
        RECT -27.960 5.600 -27.650 6.040 ;
        RECT -22.880 5.220 -22.650 6.330 ;
        RECT -21.660 5.220 -21.430 10.050 ;
        RECT -20.860 9.900 -20.540 10.220 ;
        RECT -20.830 6.210 -20.510 6.530 ;
        RECT -19.370 5.230 -18.950 11.270 ;
        RECT -10.420 5.220 -10.000 11.270 ;
        RECT -7.940 5.220 -7.710 11.270 ;
        RECT -6.720 10.060 -6.490 11.270 ;
        RECT -1.720 10.450 -1.410 10.890 ;
        RECT -6.720 9.270 -6.460 10.060 ;
        RECT -1.570 9.490 -1.250 9.810 ;
        RECT -6.720 7.120 -6.490 9.270 ;
        RECT -0.600 8.700 -0.360 8.830 ;
        RECT -0.600 8.380 -0.340 8.700 ;
        RECT -3.720 7.400 -3.440 7.450 ;
        RECT -6.720 6.330 -6.460 7.120 ;
        RECT -3.720 7.100 -3.400 7.400 ;
        RECT -1.570 6.730 -1.250 7.050 ;
        RECT 1.260 6.880 1.580 7.200 ;
        RECT -6.720 5.220 -6.490 6.330 ;
        RECT -1.820 6.280 -1.500 6.600 ;
        RECT -2.930 5.750 -2.610 6.070 ;
        RECT -17.660 4.630 -17.490 4.800 ;
        RECT -11.870 4.630 -11.700 4.800 ;
        RECT -2.200 4.470 -1.880 4.790 ;
        RECT -0.990 4.700 -0.670 5.020 ;
        RECT 1.310 4.660 1.630 4.980 ;
        RECT -17.680 4.040 -17.360 4.340 ;
        RECT -17.650 3.940 -17.480 4.040 ;
        RECT -11.980 3.970 -11.660 4.290 ;
        RECT -11.870 3.950 -11.700 3.970 ;
        RECT -0.990 3.870 -0.670 4.190 ;
        RECT 1.300 3.940 1.620 4.260 ;
        RECT -1.040 3.220 -0.720 3.540 ;
        RECT -1.040 2.390 -0.720 2.710 ;
        RECT -11.980 1.460 -11.660 1.760 ;
        RECT -0.990 1.740 -0.670 2.060 ;
        RECT 1.220 1.690 1.540 2.010 ;
      LAYER via ;
        RECT -27.940 10.480 -27.680 10.740 ;
        RECT -28.090 9.520 -27.830 9.780 ;
        RECT -29.030 8.410 -28.770 8.670 ;
        RECT -29.030 7.810 -28.770 8.070 ;
        RECT -28.090 6.760 -27.830 7.020 ;
        RECT -27.940 5.750 -27.680 6.010 ;
        RECT -20.830 9.930 -20.570 10.190 ;
        RECT -20.800 6.240 -20.540 6.500 ;
        RECT -1.690 10.480 -1.430 10.740 ;
        RECT -1.540 9.520 -1.280 9.780 ;
        RECT -0.600 8.410 -0.340 8.670 ;
        RECT -3.690 7.120 -3.430 7.380 ;
        RECT -1.540 6.760 -1.280 7.020 ;
        RECT 1.290 6.910 1.550 7.170 ;
        RECT -1.790 6.310 -1.530 6.570 ;
        RECT -2.900 5.780 -2.640 6.040 ;
        RECT -2.170 4.500 -1.910 4.760 ;
        RECT -0.960 4.730 -0.700 4.990 ;
        RECT 1.340 4.690 1.600 4.950 ;
        RECT -17.650 4.060 -17.390 4.320 ;
        RECT -11.950 4.000 -11.690 4.260 ;
        RECT -0.960 3.900 -0.700 4.160 ;
        RECT 1.330 3.970 1.590 4.230 ;
        RECT -1.010 3.250 -0.750 3.510 ;
        RECT -1.010 2.420 -0.750 2.680 ;
        RECT -0.960 1.770 -0.700 2.030 ;
        RECT -11.950 1.480 -11.690 1.740 ;
        RECT 1.250 1.720 1.510 1.980 ;
      LAYER met2 ;
        RECT -27.960 10.770 -27.650 10.780 ;
        RECT -1.720 10.770 -1.410 10.780 ;
        RECT -30.130 10.590 -18.600 10.770 ;
        RECT -10.770 10.590 0.760 10.770 ;
        RECT -27.960 10.450 -27.650 10.590 ;
        RECT -1.720 10.450 -1.410 10.590 ;
        RECT -20.850 10.180 -20.540 10.230 ;
        RECT -20.850 10.170 -20.390 10.180 ;
        RECT -20.850 9.990 -18.600 10.170 ;
        RECT -20.850 9.900 -20.540 9.990 ;
        RECT -28.110 9.750 -27.800 9.820 ;
        RECT -30.130 9.740 -27.800 9.750 ;
        RECT -1.570 9.750 -1.260 9.820 ;
        RECT -30.130 9.530 -18.600 9.740 ;
        RECT -28.820 9.520 -18.600 9.530 ;
        RECT -1.570 9.530 0.760 9.750 ;
        RECT -28.110 9.490 -27.800 9.520 ;
        RECT -1.570 9.490 -1.260 9.530 ;
        RECT -29.060 8.550 -18.600 8.770 ;
        RECT -29.060 8.410 -28.740 8.550 ;
        RECT -29.040 8.070 -28.780 8.410 ;
        RECT -29.060 7.810 -28.740 8.070 ;
        RECT -20.820 6.460 -20.510 6.540 ;
        RECT -20.820 6.250 -18.600 6.460 ;
        RECT -20.820 6.210 -20.510 6.250 ;
        RECT -27.960 5.900 -27.650 6.040 ;
        RECT -30.130 5.890 -27.650 5.900 ;
        RECT -30.130 5.740 -18.600 5.890 ;
        RECT -30.130 5.720 -27.650 5.740 ;
        RECT -27.960 5.710 -27.650 5.720 ;
        RECT -16.860 4.730 -7.850 4.950 ;
        RECT -17.680 4.290 -17.360 4.340 ;
        RECT -17.680 4.040 -11.660 4.290 ;
        RECT -11.980 3.970 -11.660 4.040 ;
        RECT -16.810 2.950 -11.150 3.170 ;
        RECT -11.370 2.620 -11.150 2.950 ;
        RECT -8.070 3.120 -7.850 4.730 ;
        RECT -8.070 2.900 -5.220 3.120 ;
        RECT -1.040 2.670 -0.730 2.710 ;
        RECT -7.000 2.620 -0.730 2.670 ;
        RECT -11.370 2.460 -0.730 2.620 ;
        RECT -11.370 2.400 -6.610 2.460 ;
        RECT -1.040 2.380 -0.730 2.460 ;
        RECT -0.990 1.980 -0.680 2.060 ;
        RECT 1.220 1.980 1.530 2.020 ;
        RECT -0.990 1.750 1.720 1.980 ;
        RECT -0.990 1.730 -0.680 1.750 ;
        RECT 1.220 1.690 1.530 1.750 ;
  END
END sky130_hilas_TA2Cell_1FG

MACRO sky130_hilas_swc4x1cellOverlap
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x1cellOverlap ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 6.710 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 4.870 6.360 7.590 6.650 ;
        RECT 0.010 4.500 1.740 6.360 ;
        RECT 0.000 2.660 1.740 4.500 ;
        RECT 4.870 6.350 10.070 6.360 ;
        RECT 4.870 3.560 10.080 6.350 ;
        RECT 0.010 0.310 1.740 2.660 ;
        RECT 4.860 0.330 10.080 3.560 ;
        RECT 4.860 0.320 10.070 0.330 ;
        RECT 4.860 0.060 7.580 0.320 ;
      LAYER li1 ;
        RECT 5.270 5.080 7.220 6.250 ;
        RECT 7.620 5.950 7.940 5.960 ;
        RECT 7.620 5.780 8.200 5.950 ;
        RECT 7.620 5.730 7.950 5.780 ;
        RECT 7.620 5.700 7.940 5.730 ;
        RECT 9.480 5.680 9.680 6.030 ;
        RECT 7.620 5.370 7.940 5.410 ;
        RECT 7.620 5.330 7.950 5.370 ;
        RECT 7.620 5.160 8.200 5.330 ;
        RECT 7.620 5.150 7.940 5.160 ;
        RECT 8.750 5.090 8.950 5.660 ;
        RECT 9.480 5.650 9.690 5.680 ;
        RECT 9.470 5.060 9.690 5.650 ;
        RECT 5.270 3.550 7.220 4.720 ;
        RECT 7.620 4.520 7.940 4.530 ;
        RECT 7.620 4.350 8.200 4.520 ;
        RECT 7.620 4.310 7.950 4.350 ;
        RECT 7.620 4.270 7.940 4.310 ;
        RECT 8.750 4.020 8.950 4.590 ;
        RECT 9.470 4.030 9.690 4.620 ;
        RECT 9.480 4.000 9.690 4.030 ;
        RECT 7.620 3.950 7.940 3.980 ;
        RECT 7.620 3.900 7.950 3.950 ;
        RECT 7.620 3.730 8.200 3.900 ;
        RECT 7.620 3.720 7.940 3.730 ;
        RECT 9.480 3.650 9.680 4.000 ;
        RECT 0.430 3.110 0.980 3.540 ;
        RECT 8.870 3.250 9.310 3.420 ;
        RECT 5.260 1.990 7.210 3.160 ;
        RECT 7.620 2.940 7.940 2.950 ;
        RECT 7.620 2.770 8.200 2.940 ;
        RECT 7.620 2.720 7.950 2.770 ;
        RECT 7.620 2.690 7.940 2.720 ;
        RECT 9.480 2.670 9.680 3.020 ;
        RECT 7.620 2.360 7.940 2.400 ;
        RECT 7.620 2.320 7.950 2.360 ;
        RECT 7.620 2.150 8.200 2.320 ;
        RECT 7.620 2.140 7.940 2.150 ;
        RECT 8.750 2.080 8.950 2.650 ;
        RECT 9.480 2.640 9.690 2.670 ;
        RECT 9.470 2.050 9.690 2.640 ;
        RECT 5.260 0.450 7.210 1.620 ;
        RECT 7.620 1.520 7.940 1.530 ;
        RECT 7.620 1.350 8.200 1.520 ;
        RECT 7.620 1.310 7.950 1.350 ;
        RECT 7.620 1.270 7.940 1.310 ;
        RECT 8.750 1.020 8.950 1.590 ;
        RECT 9.470 1.030 9.690 1.620 ;
        RECT 9.480 1.000 9.690 1.030 ;
        RECT 7.620 0.950 7.940 0.980 ;
        RECT 7.620 0.900 7.950 0.950 ;
        RECT 7.620 0.730 8.200 0.900 ;
        RECT 7.620 0.720 7.940 0.730 ;
        RECT 9.480 0.650 9.680 1.000 ;
      LAYER mcon ;
        RECT 5.750 5.910 5.920 6.080 ;
        RECT 5.750 5.570 5.920 5.740 ;
        RECT 7.680 5.740 7.850 5.910 ;
        RECT 8.760 5.450 8.930 5.620 ;
        RECT 5.750 5.230 5.920 5.400 ;
        RECT 7.680 5.190 7.850 5.360 ;
        RECT 9.490 5.480 9.660 5.650 ;
        RECT 5.750 4.380 5.920 4.550 ;
        RECT 7.680 4.320 7.850 4.490 ;
        RECT 5.750 4.040 5.920 4.210 ;
        RECT 8.760 4.060 8.930 4.230 ;
        RECT 9.490 4.030 9.660 4.200 ;
        RECT 5.750 3.700 5.920 3.870 ;
        RECT 7.680 3.770 7.850 3.940 ;
        RECT 0.430 3.190 0.700 3.460 ;
        RECT 9.130 3.250 9.310 3.420 ;
        RECT 5.740 2.820 5.910 2.990 ;
        RECT 7.680 2.730 7.850 2.900 ;
        RECT 5.740 2.480 5.910 2.650 ;
        RECT 8.760 2.440 8.930 2.610 ;
        RECT 5.740 2.140 5.910 2.310 ;
        RECT 7.680 2.180 7.850 2.350 ;
        RECT 9.490 2.470 9.660 2.640 ;
        RECT 5.740 1.280 5.910 1.450 ;
        RECT 7.680 1.320 7.850 1.490 ;
        RECT 5.740 0.940 5.910 1.110 ;
        RECT 8.760 1.060 8.930 1.230 ;
        RECT 9.490 1.030 9.660 1.200 ;
        RECT 5.740 0.600 5.910 0.770 ;
        RECT 7.680 0.770 7.850 0.940 ;
      LAYER met1 ;
        RECT 0.360 0.310 0.760 6.300 ;
        RECT 5.710 5.660 5.970 6.140 ;
        RECT 7.610 5.670 7.930 5.990 ;
        RECT 8.750 5.680 8.910 6.360 ;
        RECT 8.750 5.660 8.950 5.680 ;
        RECT 5.700 5.140 5.970 5.660 ;
        RECT 5.700 4.690 5.960 5.140 ;
        RECT 7.610 5.120 7.930 5.440 ;
        RECT 8.730 5.420 8.960 5.660 ;
        RECT 8.750 5.200 8.950 5.420 ;
        RECT 9.120 5.370 9.310 6.360 ;
        RECT 9.560 5.710 9.720 6.360 ;
        RECT 9.140 5.250 9.310 5.370 ;
        RECT 5.710 4.130 5.970 4.610 ;
        RECT 7.610 4.240 7.930 4.560 ;
        RECT 8.750 4.480 8.910 5.200 ;
        RECT 8.750 4.260 8.950 4.480 ;
        RECT 9.150 4.430 9.310 5.250 ;
        RECT 9.450 5.160 9.720 5.710 ;
        RECT 9.450 5.110 9.730 5.160 ;
        RECT 9.560 5.020 9.730 5.110 ;
        RECT 9.560 4.660 9.720 5.020 ;
        RECT 9.560 4.570 9.730 4.660 ;
        RECT 9.140 4.310 9.310 4.430 ;
        RECT 5.700 3.610 5.970 4.130 ;
        RECT 8.730 4.020 8.960 4.260 ;
        RECT 7.610 3.690 7.930 4.010 ;
        RECT 8.750 4.000 8.950 4.020 ;
        RECT 5.700 3.160 5.960 3.610 ;
        RECT 5.700 2.570 5.960 3.050 ;
        RECT 7.610 2.660 7.930 2.980 ;
        RECT 8.750 2.670 8.910 4.000 ;
        RECT 9.120 3.450 9.310 4.310 ;
        RECT 9.450 4.520 9.730 4.570 ;
        RECT 9.450 3.970 9.720 4.520 ;
        RECT 9.100 3.220 9.340 3.450 ;
        RECT 8.750 2.650 8.950 2.670 ;
        RECT 5.690 2.050 5.960 2.570 ;
        RECT 7.610 2.110 7.930 2.430 ;
        RECT 8.730 2.410 8.960 2.650 ;
        RECT 8.750 2.190 8.950 2.410 ;
        RECT 9.120 2.360 9.310 3.220 ;
        RECT 9.560 2.700 9.720 3.970 ;
        RECT 9.140 2.240 9.310 2.360 ;
        RECT 5.690 1.600 5.950 2.050 ;
        RECT 5.700 1.030 5.960 1.510 ;
        RECT 7.610 1.240 7.930 1.560 ;
        RECT 8.750 1.480 8.910 2.190 ;
        RECT 8.750 1.260 8.950 1.480 ;
        RECT 9.150 1.430 9.310 2.240 ;
        RECT 9.450 2.150 9.720 2.700 ;
        RECT 9.450 2.100 9.730 2.150 ;
        RECT 9.560 2.010 9.730 2.100 ;
        RECT 9.560 1.660 9.720 2.010 ;
        RECT 9.560 1.570 9.730 1.660 ;
        RECT 9.140 1.310 9.310 1.430 ;
        RECT 5.690 0.510 5.960 1.030 ;
        RECT 8.730 1.020 8.960 1.260 ;
        RECT 7.610 0.690 7.930 1.010 ;
        RECT 8.750 1.000 8.950 1.020 ;
        RECT 5.690 0.060 5.950 0.510 ;
        RECT 8.750 0.320 8.910 1.000 ;
        RECT 9.120 0.320 9.310 1.310 ;
        RECT 9.450 1.520 9.730 1.570 ;
        RECT 9.450 0.970 9.720 1.520 ;
        RECT 9.560 0.320 9.720 0.970 ;
      LAYER via ;
        RECT 7.640 5.700 7.900 5.960 ;
        RECT 7.640 5.150 7.900 5.410 ;
        RECT 7.640 4.270 7.900 4.530 ;
        RECT 7.640 3.720 7.900 3.980 ;
        RECT 7.640 2.690 7.900 2.950 ;
        RECT 7.640 2.140 7.900 2.400 ;
        RECT 7.640 1.270 7.900 1.530 ;
        RECT 7.640 0.720 7.900 0.980 ;
      LAYER met2 ;
        RECT 7.610 5.860 7.920 6.000 ;
        RECT 0.000 5.680 10.080 5.860 ;
        RECT 7.610 5.670 7.920 5.680 ;
        RECT 7.610 5.430 7.920 5.450 ;
        RECT 0.000 5.250 10.080 5.430 ;
        RECT 7.610 5.120 7.920 5.250 ;
        RECT 7.610 4.430 7.920 4.560 ;
        RECT 0.000 4.250 10.080 4.430 ;
        RECT 7.610 4.230 7.920 4.250 ;
        RECT 7.610 4.000 7.920 4.010 ;
        RECT 0.000 3.930 7.600 4.000 ;
        RECT 7.610 3.930 10.080 4.000 ;
        RECT 0.000 3.820 10.080 3.930 ;
        RECT 7.610 3.680 7.920 3.820 ;
        RECT 7.610 2.850 7.920 2.990 ;
        RECT 7.610 2.840 10.080 2.850 ;
        RECT 0.020 2.670 10.080 2.840 ;
        RECT 7.610 2.660 7.920 2.670 ;
        RECT 7.610 2.420 7.920 2.440 ;
        RECT 0.020 2.250 10.080 2.420 ;
        RECT 7.520 2.240 10.080 2.250 ;
        RECT 7.610 2.110 7.920 2.240 ;
        RECT 7.610 1.440 7.920 1.560 ;
        RECT 0.020 1.430 7.920 1.440 ;
        RECT 0.020 1.270 10.080 1.430 ;
        RECT 0.800 1.180 2.340 1.270 ;
        RECT 7.520 1.250 10.080 1.270 ;
        RECT 7.610 1.230 7.920 1.250 ;
        RECT 7.610 1.000 7.920 1.010 ;
        RECT 0.020 0.830 10.080 1.000 ;
        RECT 7.610 0.820 10.080 0.830 ;
        RECT 7.610 0.680 7.920 0.820 ;
  END
END sky130_hilas_swc4x1cellOverlap

MACRO sky130_hilas_capacitorSize02
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize02 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.970 BY 5.830 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 7.230 2.620 7.890 3.280 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 0.110 3.200 0.770 3.260 ;
        RECT 1.160 3.200 2.170 3.210 ;
        RECT 0.110 2.700 3.800 3.200 ;
        RECT 0.110 2.690 1.520 2.700 ;
        RECT 0.110 2.600 0.770 2.690 ;
        RECT 3.160 1.580 3.790 2.700 ;
        RECT 3.160 1.570 5.310 1.580 ;
        RECT 1.840 1.270 5.310 1.570 ;
        RECT 1.840 1.100 4.850 1.270 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 0.000 5.280 7.970 5.460 ;
        RECT 0.000 4.850 7.970 5.030 ;
        RECT 0.030 3.850 7.970 4.030 ;
        RECT 0.030 3.420 7.970 3.600 ;
        RECT 0.240 3.080 0.610 3.140 ;
        RECT 0.020 2.800 0.610 3.080 ;
        RECT 0.240 2.740 0.610 2.800 ;
        RECT 7.360 3.100 7.730 3.160 ;
        RECT 7.360 2.820 7.970 3.100 ;
        RECT 7.360 2.760 7.730 2.820 ;
        RECT 0.030 2.270 7.970 2.440 ;
        RECT 0.030 1.850 7.970 2.020 ;
        RECT 0.030 0.870 7.970 1.040 ;
        RECT 0.030 0.430 7.970 0.600 ;
      LAYER via2 ;
        RECT 0.290 2.800 0.570 3.080 ;
        RECT 7.410 2.820 7.690 3.100 ;
      LAYER met3 ;
        RECT 1.460 5.800 3.770 5.830 ;
        RECT 1.460 3.310 5.690 5.800 ;
        RECT 0.020 2.540 0.810 3.290 ;
        RECT 1.460 2.560 7.930 3.310 ;
        RECT 1.460 0.020 5.690 2.560 ;
        RECT 3.740 0.000 5.690 0.020 ;
      LAYER via3 ;
        RECT 0.210 2.690 0.640 3.170 ;
        RECT 7.330 2.710 7.760 3.190 ;
  END
END sky130_hilas_capacitorSize02

MACRO sky130_hilas_TopProtectStructure
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TopProtectStructure ;
  ORIGIN 154.680 243.370 ;
  SIZE 372.850 BY 389.100 ;
  PIN IO07
    PORT
      LAYER met1 ;
        RECT 215.620 -58.690 216.210 -58.680 ;
        RECT 215.620 -62.290 218.170 -58.690 ;
        RECT 214.270 -62.580 218.170 -62.290 ;
    END
  END IO07
  PIN IO08
    PORT
      LAYER met1 ;
        RECT 216.920 -30.090 218.170 -30.080 ;
        RECT 215.620 -33.700 218.170 -30.090 ;
        RECT 214.270 -33.970 218.170 -33.700 ;
        RECT 214.270 -33.980 216.920 -33.970 ;
        RECT 214.270 -33.990 216.210 -33.980 ;
    END
  END IO08
  PIN IO09
    PORT
      LAYER met1 ;
        RECT 215.620 -5.110 218.150 -1.500 ;
        RECT 214.270 -5.390 218.150 -5.110 ;
        RECT 214.270 -5.400 216.210 -5.390 ;
    END
  END IO09
  PIN IO10
    PORT
      LAYER met1 ;
        RECT 216.920 27.100 218.170 27.110 ;
        RECT 216.200 27.090 218.170 27.100 ;
        RECT 215.620 23.480 218.170 27.090 ;
        RECT 214.270 23.220 218.170 23.480 ;
        RECT 214.270 23.210 216.920 23.220 ;
        RECT 214.270 23.190 216.210 23.210 ;
    END
  END IO10
  PIN IO11
    PORT
      LAYER met1 ;
        RECT 215.620 55.670 216.210 55.680 ;
        RECT 215.620 52.070 218.160 55.670 ;
        RECT 214.270 51.780 218.160 52.070 ;
    END
  END IO11
  PIN IO12
    PORT
      LAYER met1 ;
        RECT 215.620 80.660 218.160 84.270 ;
        RECT 214.270 80.380 218.160 80.660 ;
        RECT 214.270 80.370 216.210 80.380 ;
    END
  END IO12
  PIN IO13
    PORT
      LAYER met1 ;
        RECT 216.920 112.860 218.170 112.870 ;
        RECT 215.620 109.250 218.170 112.860 ;
        RECT 214.270 108.980 218.170 109.250 ;
        RECT 214.270 108.970 216.920 108.980 ;
        RECT 214.270 108.960 216.210 108.970 ;
    END
  END IO13
  PIN IO25
    PORT
      LAYER met1 ;
        RECT -153.430 113.570 -152.030 113.580 ;
        RECT -154.680 109.970 -152.030 113.570 ;
        RECT -154.680 109.680 -150.680 109.970 ;
    END
  END IO25
  PIN IO26
    PORT
      LAYER met1 ;
        RECT -154.670 81.380 -152.030 84.990 ;
        RECT -154.670 81.100 -150.680 81.380 ;
        RECT -153.430 81.090 -150.680 81.100 ;
    END
  END IO26
  PIN IO27
    PORT
      LAYER met1 ;
        RECT -153.430 56.390 -152.030 56.400 ;
        RECT -154.680 52.790 -152.030 56.390 ;
        RECT -154.680 52.500 -150.680 52.790 ;
    END
  END IO27
  PIN IO28
    PORT
      LAYER met1 ;
        RECT -153.420 27.800 -152.030 27.810 ;
        RECT -154.660 24.200 -152.030 27.800 ;
        RECT -154.660 23.910 -150.680 24.200 ;
    END
  END IO28
  PIN IO29
    PORT
      LAYER met1 ;
        RECT -154.670 -4.390 -152.030 -0.780 ;
        RECT -154.670 -4.670 -150.680 -4.390 ;
        RECT -153.430 -4.680 -150.680 -4.670 ;
    END
  END IO29
  PIN IO30
    PORT
      LAYER met1 ;
        RECT -153.430 -29.380 -152.030 -29.370 ;
        RECT -154.680 -32.980 -152.030 -29.380 ;
        RECT -154.680 -33.270 -150.680 -32.980 ;
    END
  END IO30
  PIN IO31
    PORT
      LAYER met1 ;
        RECT -153.430 -57.960 -152.620 -57.950 ;
        RECT -154.670 -61.570 -152.030 -57.960 ;
        RECT -154.670 -61.850 -150.680 -61.570 ;
        RECT -152.620 -61.860 -150.680 -61.850 ;
    END
  END IO31
  PIN IO32
    PORT
      LAYER met1 ;
        RECT -154.640 -86.550 -152.600 -86.540 ;
        RECT -154.640 -90.160 -152.030 -86.550 ;
        RECT -154.640 -90.430 -150.680 -90.160 ;
        RECT -153.410 -90.440 -150.680 -90.430 ;
        RECT -152.620 -90.450 -150.680 -90.440 ;
    END
  END IO32
  PIN IO33
    PORT
      LAYER met1 ;
        RECT -153.420 -115.150 -152.030 -115.140 ;
        RECT -154.660 -118.750 -152.030 -115.150 ;
        RECT -154.660 -119.040 -150.680 -118.750 ;
    END
  END IO33
  PIN IO34
    PORT
      LAYER met1 ;
        RECT -153.420 -143.740 -152.030 -143.730 ;
        RECT -154.670 -147.340 -152.030 -143.740 ;
        RECT -154.670 -147.630 -150.680 -147.340 ;
    END
  END IO34
  PIN IO35
    PORT
      LAYER met1 ;
        RECT -153.420 -172.330 -152.030 -172.320 ;
        RECT -154.670 -175.930 -152.030 -172.330 ;
        RECT -154.670 -176.220 -150.680 -175.930 ;
    END
  END IO35
  PIN IO36
    PORT
      LAYER met1 ;
        RECT -153.410 -200.920 -152.030 -200.910 ;
        RECT -154.660 -204.520 -152.030 -200.920 ;
        RECT -154.660 -204.810 -150.680 -204.520 ;
    END
  END IO36
  PIN IO37
    PORT
      LAYER met1 ;
        RECT -154.660 -233.110 -152.030 -229.500 ;
        RECT -154.660 -233.390 -150.680 -233.110 ;
        RECT -153.430 -233.400 -150.680 -233.390 ;
    END
  END IO37
  PIN VSSA1
    ANTENNADIFFAREA 783.889587 ;
    PORT
      LAYER met2 ;
        RECT -151.260 141.640 -53.000 141.650 ;
        RECT -151.390 140.250 -53.000 141.640 ;
        RECT -151.390 138.730 -149.100 140.250 ;
        RECT -138.300 140.240 -137.370 140.250 ;
        RECT -109.710 140.240 -108.780 140.250 ;
        RECT -81.120 140.240 -80.190 140.250 ;
        RECT -138.050 139.130 -137.880 140.240 ;
        RECT -109.460 139.130 -109.290 140.240 ;
        RECT -80.870 139.130 -80.700 140.240 ;
        RECT -150.940 138.690 -149.100 138.730 ;
        RECT -150.500 130.560 -149.100 138.690 ;
        RECT -150.530 130.170 -149.100 130.560 ;
        RECT -150.530 103.370 -149.130 130.170 ;
        RECT -150.530 102.860 -149.120 103.370 ;
        RECT -150.530 102.690 -148.010 102.860 ;
        RECT -150.530 102.440 -149.120 102.690 ;
        RECT -150.530 74.780 -149.130 102.440 ;
        RECT -150.530 74.270 -149.120 74.780 ;
        RECT -150.530 74.100 -148.010 74.270 ;
        RECT -150.530 73.850 -149.120 74.100 ;
        RECT -150.530 46.190 -149.130 73.850 ;
        RECT -150.530 45.680 -149.120 46.190 ;
        RECT -150.530 45.510 -148.010 45.680 ;
        RECT -150.530 45.260 -149.120 45.510 ;
        RECT -150.530 17.600 -149.130 45.260 ;
        RECT -150.530 17.090 -149.120 17.600 ;
        RECT -150.530 16.920 -148.010 17.090 ;
        RECT -150.530 16.670 -149.120 16.920 ;
        RECT -150.530 -10.990 -149.130 16.670 ;
        RECT -150.530 -11.500 -149.120 -10.990 ;
        RECT -150.530 -11.670 -148.010 -11.500 ;
        RECT -150.530 -11.920 -149.120 -11.670 ;
        RECT -150.530 -39.580 -149.130 -11.920 ;
        RECT -150.530 -40.090 -149.120 -39.580 ;
        RECT -150.530 -40.260 -148.010 -40.090 ;
        RECT -150.530 -40.510 -149.120 -40.260 ;
        RECT -150.530 -68.170 -149.130 -40.510 ;
        RECT -150.530 -68.680 -149.120 -68.170 ;
        RECT -150.530 -68.850 -148.010 -68.680 ;
        RECT -150.530 -69.100 -149.120 -68.850 ;
        RECT -150.530 -96.760 -149.130 -69.100 ;
        RECT -150.530 -97.270 -149.120 -96.760 ;
        RECT -150.530 -97.440 -148.010 -97.270 ;
        RECT -150.530 -97.690 -149.120 -97.440 ;
        RECT -150.530 -125.350 -149.130 -97.690 ;
        RECT -150.530 -125.860 -149.120 -125.350 ;
        RECT -150.530 -126.030 -148.010 -125.860 ;
        RECT -150.530 -126.280 -149.120 -126.030 ;
        RECT -150.530 -153.940 -149.130 -126.280 ;
        RECT -150.530 -154.450 -149.120 -153.940 ;
        RECT -150.530 -154.620 -148.010 -154.450 ;
        RECT -150.530 -154.870 -149.120 -154.620 ;
        RECT -150.530 -182.530 -149.130 -154.870 ;
        RECT -150.530 -183.040 -149.120 -182.530 ;
        RECT -150.530 -183.210 -148.010 -183.040 ;
        RECT -150.530 -183.460 -149.120 -183.210 ;
        RECT -150.530 -211.120 -149.130 -183.460 ;
        RECT -150.530 -211.630 -149.120 -211.120 ;
        RECT -150.530 -211.800 -148.010 -211.630 ;
        RECT -150.530 -212.050 -149.120 -211.800 ;
        RECT -150.530 -239.710 -149.130 -212.050 ;
        RECT -150.530 -240.220 -149.120 -239.710 ;
        RECT -150.530 -240.390 -148.010 -240.220 ;
        RECT -150.530 -240.640 -149.120 -240.390 ;
        RECT -150.530 -243.040 -149.130 -240.640 ;
    END
  END VSSA1
  PIN ANALOG10
    PORT
      LAYER met1 ;
        RECT -131.060 143.740 -127.170 145.710 ;
        RECT -131.060 143.150 -127.160 143.740 ;
        RECT -131.060 141.800 -130.770 143.150 ;
    END
  END ANALOG10
  PIN ANALOG09
    PORT
      LAYER met1 ;
        RECT -102.470 143.740 -98.580 145.700 ;
        RECT -102.470 143.150 -98.570 143.740 ;
        RECT -102.470 141.800 -102.180 143.150 ;
    END
  END ANALOG09
  PIN ANALOG08
    PORT
      LAYER met1 ;
        RECT -73.880 143.740 -69.990 145.700 ;
        RECT -73.880 143.150 -69.980 143.740 ;
        RECT -73.880 141.800 -73.590 143.150 ;
    END
  END ANALOG08
  PIN ANALOG07
    PORT
      LAYER met1 ;
        RECT -31.980 143.760 -28.090 145.730 ;
    END
  END ANALOG07
  PIN ANALOG06
    ANTENNAGATEAREA 62.701500 ;
    ANTENNADIFFAREA 1693.265747 ;
    PORT
      LAYER nwell ;
        RECT -123.900 134.780 -111.850 140.720 ;
        RECT -95.310 134.780 -83.260 140.720 ;
        RECT -66.720 134.780 -54.670 140.720 ;
        RECT -149.600 116.840 -143.660 128.890 ;
        RECT -23.810 124.410 -21.070 127.910 ;
        RECT -1.370 127.900 1.340 127.940 ;
        RECT -6.930 121.910 -2.930 127.900 ;
        RECT -1.380 126.250 1.340 127.900 ;
        RECT -1.370 124.910 1.340 124.950 ;
        RECT -1.380 122.250 1.340 124.910 ;
        RECT 11.320 110.490 13.090 116.730 ;
        RECT 52.460 110.840 55.770 115.460 ;
        RECT 62.250 114.720 63.980 115.470 ;
        RECT 62.240 111.150 63.980 114.720 ;
        RECT 75.580 113.080 78.300 114.730 ;
        RECT 75.580 113.040 78.290 113.080 ;
        RECT -10.540 107.330 -7.970 110.420 ;
        RECT 32.120 110.090 33.850 110.840 ;
        RECT 32.110 109.690 33.850 110.090 ;
        RECT 32.110 106.520 36.110 109.690 ;
        RECT 49.910 109.430 55.770 110.840 ;
        RECT 62.250 109.430 63.980 111.150 ;
        RECT 75.580 111.710 78.290 111.750 ;
        RECT 75.580 110.350 78.300 111.710 ;
        RECT 80.030 111.650 83.340 115.470 ;
        RECT 79.380 111.640 84.510 111.650 ;
        RECT 79.370 110.350 84.510 111.640 ;
        RECT 75.580 110.060 84.510 110.350 ;
        RECT 77.660 109.430 84.510 110.060 ;
        RECT 49.910 107.020 53.220 109.430 ;
        RECT 49.260 107.010 54.390 107.020 ;
        RECT 32.120 104.800 36.110 106.520 ;
        RECT 32.690 103.640 36.110 104.800 ;
        RECT 49.250 104.800 54.390 107.010 ;
        RECT 49.250 100.970 51.110 104.800 ;
        RECT 53.110 103.530 54.390 104.800 ;
        RECT 77.660 105.600 81.230 109.430 ;
        RECT 83.230 105.600 84.510 109.430 ;
        RECT 77.660 104.300 80.420 105.600 ;
        RECT 53.110 101.670 54.840 103.530 ;
        RECT -149.600 88.250 -143.660 100.300 ;
        RECT 53.100 99.830 54.840 101.670 ;
        RECT 25.090 93.700 27.640 93.710 ;
        RECT 25.080 89.890 27.640 93.700 ;
        RECT 29.170 89.890 31.400 93.710 ;
        RECT 32.690 93.570 36.110 99.620 ;
        RECT 53.110 97.480 54.840 99.830 ;
        RECT 60.620 103.520 63.170 103.530 ;
        RECT 60.620 97.500 63.180 103.520 ;
        RECT 60.620 97.490 63.170 97.500 ;
        RECT 33.420 93.080 35.150 93.570 ;
        RECT 33.420 90.010 35.160 93.080 ;
        RECT 25.080 89.880 31.400 89.890 ;
        RECT 25.080 89.730 27.750 89.880 ;
        RECT 25.080 89.720 27.930 89.730 ;
        RECT -10.000 85.530 -9.440 87.500 ;
        RECT 11.320 83.030 13.090 89.270 ;
        RECT 17.050 83.030 19.560 89.270 ;
        RECT 25.080 87.680 27.750 89.720 ;
        RECT 25.090 87.670 27.750 87.680 ;
        RECT 25.600 83.850 27.750 87.670 ;
        RECT 29.170 87.660 31.400 89.880 ;
        RECT 33.030 89.860 33.410 89.890 ;
        RECT 33.420 89.860 35.150 90.010 ;
        RECT 25.600 83.830 27.350 83.850 ;
        RECT 32.690 83.810 36.110 89.860 ;
        RECT -149.600 59.660 -143.660 71.710 ;
        RECT 80.140 60.580 81.490 76.050 ;
        RECT 80.130 60.110 81.490 60.580 ;
        RECT -149.600 31.070 -143.660 43.120 ;
        RECT -149.600 2.480 -143.660 14.530 ;
        RECT -149.600 -26.110 -143.660 -14.060 ;
        RECT -149.600 -54.700 -143.660 -42.650 ;
        RECT -149.600 -83.290 -143.660 -71.240 ;
        RECT -149.600 -111.880 -143.660 -99.830 ;
        RECT -149.600 -140.470 -143.660 -128.420 ;
        RECT -149.600 -169.060 -143.660 -157.010 ;
        RECT -149.600 -197.650 -143.660 -185.600 ;
        RECT -149.600 -226.240 -143.660 -214.190 ;
      LAYER met3 ;
        RECT 49.510 113.180 49.960 113.930 ;
        RECT 49.510 107.020 49.880 113.180 ;
        RECT 50.550 113.170 51.000 113.920 ;
        RECT 50.630 110.530 51.000 113.170 ;
        RECT 50.630 109.930 51.070 110.530 ;
        RECT 49.510 106.690 50.000 107.020 ;
        RECT 49.560 106.530 50.000 106.690 ;
        RECT 50.630 104.820 51.000 109.930 ;
        RECT 50.620 103.950 51.090 104.820 ;
    END
  END ANALOG06
  PIN ANALOG05
    PORT
      LAYER met1 ;
        RECT 38.730 143.740 42.620 145.710 ;
        RECT 38.730 143.150 42.630 143.740 ;
        RECT 38.730 141.800 39.020 143.150 ;
    END
  END ANALOG05
  PIN ANALOG04
    PORT
      LAYER met1 ;
        RECT 67.330 143.740 71.220 145.710 ;
        RECT 67.320 143.150 71.220 143.740 ;
        RECT 67.320 141.800 67.610 143.150 ;
    END
  END ANALOG04
  PIN ANALOG03
    PORT
      LAYER met1 ;
        RECT 95.920 143.740 99.810 145.710 ;
        RECT 95.910 143.150 99.810 143.740 ;
        RECT 95.910 141.800 96.200 143.150 ;
    END
  END ANALOG03
  PIN ANALOG02
    PORT
      LAYER met1 ;
        RECT 124.510 144.540 128.400 145.710 ;
        RECT 124.500 143.740 128.390 144.540 ;
        RECT 124.500 143.150 128.400 143.740 ;
        RECT 124.500 141.800 124.790 143.150 ;
    END
  END ANALOG02
  PIN ANALOG01
    PORT
      LAYER met1 ;
        RECT 153.100 144.540 156.990 145.700 ;
        RECT 153.090 144.530 156.990 144.540 ;
        RECT 153.090 143.740 156.980 144.530 ;
        RECT 153.090 143.150 156.990 143.740 ;
        RECT 153.090 141.800 153.380 143.150 ;
    END
  END ANALOG01
  PIN ANALOG00
    PORT
      LAYER met1 ;
        RECT 181.690 143.740 185.580 145.700 ;
        RECT 181.680 143.150 185.580 143.740 ;
        RECT 181.680 141.800 181.970 143.150 ;
    END
  END ANALOG00
  PIN VSSA1
    ANTENNAGATEAREA 60.628899 ;
    ANTENNADIFFAREA 1678.220215 ;
    PORT
      LAYER met2 ;
        RECT -25.550 141.650 29.920 142.210 ;
        RECT 213.810 141.650 215.000 141.660 ;
        RECT -25.550 140.820 215.000 141.650 ;
        RECT 2.430 140.370 215.000 140.820 ;
        RECT 2.430 140.250 202.560 140.370 ;
        RECT 2.900 140.240 3.830 140.250 ;
        RECT 31.490 140.240 32.420 140.250 ;
        RECT 60.080 140.240 61.010 140.250 ;
        RECT 88.670 140.240 89.600 140.250 ;
        RECT 117.260 140.240 118.190 140.250 ;
        RECT 145.850 140.240 146.780 140.250 ;
        RECT 174.440 140.240 175.370 140.250 ;
        RECT 3.150 139.130 3.320 140.240 ;
        RECT 31.740 139.130 31.910 140.240 ;
        RECT 60.330 139.130 60.500 140.240 ;
        RECT 88.920 139.130 89.090 140.240 ;
        RECT 117.510 139.130 117.680 140.240 ;
        RECT 146.100 139.130 146.270 140.240 ;
        RECT 174.690 139.130 174.860 140.240 ;
        RECT 212.840 139.050 215.000 140.370 ;
        RECT -112.430 135.350 -111.790 138.360 ;
        RECT -83.840 135.350 -83.200 138.360 ;
        RECT -55.250 135.350 -54.610 138.360 ;
        RECT -138.770 135.280 -53.000 135.350 ;
        RECT -144.230 133.950 -53.000 135.280 ;
        RECT -144.230 133.880 -138.480 133.950 ;
        RECT -144.230 130.040 -142.830 133.880 ;
        RECT -113.330 133.820 -110.700 133.950 ;
        RECT -84.740 133.820 -82.110 133.950 ;
        RECT -56.150 133.820 -53.520 133.950 ;
        RECT -113.330 133.310 -110.780 133.820 ;
        RECT -84.740 133.310 -82.190 133.820 ;
        RECT -56.150 133.310 -53.600 133.820 ;
        RECT -113.330 133.240 -112.710 133.310 ;
        RECT -84.740 133.240 -84.120 133.310 ;
        RECT -56.150 133.240 -55.530 133.310 ;
        RECT -144.230 129.960 -142.700 130.040 ;
        RECT -144.230 128.950 -142.190 129.960 ;
        RECT -147.240 128.310 -142.190 128.950 ;
        RECT -144.230 128.030 -142.190 128.310 ;
        RECT -68.920 129.870 -64.830 130.120 ;
        RECT -26.950 129.870 -26.270 129.920 ;
        RECT -68.920 128.700 -26.270 129.870 ;
        RECT 212.840 129.840 214.120 139.050 ;
        RECT -25.720 128.700 -25.270 128.800 ;
        RECT -68.920 128.470 -25.270 128.700 ;
        RECT -144.230 127.410 -142.120 128.030 ;
        RECT -68.920 127.620 -26.270 128.470 ;
        RECT -25.720 128.370 -25.270 128.470 ;
        RECT -144.230 101.450 -142.830 127.410 ;
        RECT -68.920 127.020 -64.830 127.620 ;
        RECT -26.950 127.600 -26.270 127.620 ;
        RECT -56.220 126.510 -55.600 126.530 ;
        RECT -56.220 126.500 -24.620 126.510 ;
        RECT -23.310 126.500 -22.990 126.700 ;
        RECT -22.580 126.500 -22.270 126.710 ;
        RECT -21.900 126.500 -21.580 126.710 ;
        RECT -21.240 126.500 -6.590 126.630 ;
        RECT -56.220 126.420 -6.590 126.500 ;
        RECT -56.220 126.250 -21.100 126.420 ;
        RECT -7.170 126.410 -6.420 126.420 ;
        RECT -56.220 126.140 -21.240 126.250 ;
        RECT -56.220 126.070 -55.600 126.140 ;
        RECT -27.100 126.110 -21.240 126.140 ;
        RECT -24.830 125.740 -21.240 126.110 ;
        RECT -20.750 125.950 -20.430 126.270 ;
        RECT -7.170 126.110 -5.550 126.410 ;
        RECT 17.280 126.240 17.730 126.260 ;
        RECT 17.270 126.180 17.750 126.240 ;
        RECT -7.170 125.970 -6.930 126.110 ;
        RECT -5.850 126.050 -5.550 126.110 ;
        RECT -23.310 125.570 -22.990 125.740 ;
        RECT -22.580 125.540 -22.270 125.740 ;
        RECT -21.880 125.590 -21.560 125.740 ;
        RECT -25.620 124.900 -25.190 125.370 ;
        RECT -20.730 124.910 -20.460 125.950 ;
        RECT -7.190 125.640 -6.880 125.970 ;
        RECT -5.850 125.730 -5.520 126.050 ;
        RECT -5.120 126.040 17.750 126.180 ;
        RECT -5.830 125.720 -5.520 125.730 ;
        RECT -5.140 125.880 17.750 126.040 ;
        RECT -5.140 125.720 -4.820 125.880 ;
        RECT 17.270 125.820 17.750 125.880 ;
        RECT 17.280 125.800 17.730 125.820 ;
        RECT -5.140 125.710 -4.830 125.720 ;
        RECT -23.250 124.900 -20.460 124.910 ;
        RECT -25.620 124.890 -20.460 124.900 ;
        RECT -25.530 124.680 -20.460 124.890 ;
        RECT -25.530 124.670 -20.980 124.680 ;
        RECT -22.600 122.860 -22.290 123.070 ;
        RECT -21.170 122.860 -20.860 123.090 ;
        RECT -24.950 122.700 -20.030 122.860 ;
        RECT -26.760 122.530 -20.030 122.700 ;
        RECT 14.520 122.850 15.020 122.870 ;
        RECT 20.260 122.850 20.700 122.900 ;
        RECT 34.630 122.850 35.130 122.870 ;
        RECT -26.760 122.480 -20.020 122.530 ;
        RECT -26.760 122.370 -20.000 122.480 ;
        RECT 14.520 122.430 41.030 122.850 ;
        RECT 14.670 122.410 41.030 122.430 ;
        RECT 20.260 122.400 20.700 122.410 ;
        RECT 40.430 122.390 40.930 122.410 ;
        RECT -26.760 122.300 -24.490 122.370 ;
        RECT -52.870 122.090 -52.390 122.120 ;
        RECT -26.760 122.100 -26.360 122.300 ;
        RECT -23.390 122.160 -23.080 122.370 ;
        RECT -22.460 122.160 -22.150 122.370 ;
        RECT -21.760 122.160 -21.450 122.370 ;
        RECT -21.020 122.190 -20.000 122.370 ;
        RECT -7.910 122.190 -7.600 122.310 ;
        RECT 1.950 122.190 2.260 122.330 ;
        RECT -21.020 122.160 2.260 122.190 ;
        RECT -27.110 122.090 -26.360 122.100 ;
        RECT -52.870 121.710 -26.360 122.090 ;
        RECT -21.000 122.000 2.260 122.160 ;
        RECT -21.000 121.980 2.230 122.000 ;
        RECT -52.870 121.690 -52.390 121.710 ;
        RECT -27.110 121.700 -26.360 121.710 ;
        RECT 11.770 119.640 12.070 119.700 ;
        RECT 53.090 119.640 53.390 119.670 ;
        RECT 11.770 119.410 53.460 119.640 ;
        RECT 11.770 119.380 12.070 119.410 ;
        RECT 53.090 119.330 53.390 119.410 ;
        RECT 4.690 118.980 5.000 119.000 ;
        RECT -5.100 118.900 -4.780 118.910 ;
        RECT 4.690 118.900 5.010 118.980 ;
        RECT 28.870 118.910 29.190 118.930 ;
        RECT 28.870 118.900 29.200 118.910 ;
        RECT 35.640 118.900 35.960 118.930 ;
        RECT 50.410 118.900 50.730 118.920 ;
        RECT 65.070 118.900 65.630 119.040 ;
        RECT -5.100 118.670 65.630 118.900 ;
        RECT -5.100 118.590 -4.780 118.670 ;
        RECT 4.690 118.660 5.000 118.670 ;
        RECT 28.870 118.650 29.200 118.670 ;
        RECT 35.640 118.650 35.960 118.670 ;
        RECT 50.410 118.660 50.730 118.670 ;
        RECT 65.070 118.530 65.630 118.670 ;
        RECT 0.690 118.450 1.060 118.510 ;
        RECT 63.890 118.450 64.430 118.470 ;
        RECT -56.340 118.220 -55.720 118.310 ;
        RECT 0.690 118.220 64.430 118.450 ;
        RECT -56.340 118.100 -26.890 118.220 ;
        RECT 0.690 118.160 1.060 118.220 ;
        RECT -56.340 117.810 -24.300 118.100 ;
        RECT 32.490 118.000 32.770 118.010 ;
        RECT -56.340 117.720 -55.720 117.810 ;
        RECT -26.890 117.800 -24.300 117.810 ;
        RECT 3.520 117.990 3.830 118.000 ;
        RECT 32.470 117.990 32.790 118.000 ;
        RECT 35.200 117.990 35.520 118.020 ;
        RECT 49.520 117.990 49.840 118.050 ;
        RECT 62.810 117.990 63.350 118.000 ;
        RECT 3.520 117.760 63.350 117.990 ;
        RECT 63.890 117.910 64.430 118.220 ;
        RECT 3.520 117.730 3.850 117.760 ;
        RECT 32.470 117.740 32.790 117.760 ;
        RECT 35.200 117.740 35.520 117.760 ;
        RECT 32.490 117.730 32.770 117.740 ;
        RECT 3.520 117.710 3.830 117.730 ;
        RECT -2.560 117.530 -2.240 117.540 ;
        RECT 61.870 117.530 62.400 117.560 ;
        RECT -52.870 117.320 -52.330 117.350 ;
        RECT -52.870 117.300 -26.930 117.320 ;
        RECT -7.800 117.300 -7.400 117.310 ;
        RECT -52.870 116.950 -7.400 117.300 ;
        RECT -2.560 117.300 62.400 117.530 ;
        RECT 62.810 117.440 63.350 117.760 ;
        RECT -2.560 117.240 -2.240 117.300 ;
        RECT 61.870 116.950 62.400 117.300 ;
        RECT -52.870 116.910 -26.930 116.950 ;
        RECT -7.800 116.920 -7.400 116.950 ;
        RECT -52.870 116.870 -52.330 116.910 ;
        RECT 187.060 116.890 190.560 117.430 ;
        RECT 41.760 116.370 42.040 116.390 ;
        RECT 41.740 116.340 42.060 116.370 ;
        RECT 73.880 116.340 75.220 116.880 ;
        RECT 88.580 116.870 190.650 116.890 ;
        RECT 41.740 116.130 75.220 116.340 ;
        RECT 41.740 116.110 42.060 116.130 ;
        RECT 41.760 116.090 42.040 116.110 ;
        RECT 73.880 115.600 75.220 116.130 ;
        RECT 54.870 114.980 55.190 114.990 ;
        RECT 54.630 114.970 55.190 114.980 ;
        RECT 80.860 114.970 81.170 114.980 ;
        RECT 52.460 114.890 63.980 114.970 ;
        RECT 71.810 114.890 83.340 114.970 ;
        RECT 87.740 114.890 190.650 116.870 ;
        RECT 52.460 114.840 190.650 114.890 ;
        RECT 52.460 114.790 88.600 114.840 ;
        RECT 54.630 114.650 54.940 114.790 ;
        RECT 59.390 114.770 88.600 114.790 ;
        RECT 59.390 114.520 88.490 114.770 ;
        RECT 59.390 114.490 59.800 114.520 ;
        RECT -7.420 114.290 -7.130 114.310 ;
        RECT -19.870 113.890 -7.110 114.290 ;
        RECT -130.950 112.070 -27.430 112.110 ;
        RECT -130.950 111.200 -26.160 112.070 ;
        RECT -19.870 111.200 -19.470 113.890 ;
        RECT -7.420 113.880 -7.130 113.890 ;
        RECT 49.460 113.580 50.040 114.020 ;
        RECT 49.460 113.390 50.100 113.580 ;
        RECT -8.920 112.990 -8.610 113.080 ;
        RECT -7.410 112.990 -7.090 113.040 ;
        RECT -8.920 112.820 -7.030 112.990 ;
        RECT -8.920 112.750 -8.610 112.820 ;
        RECT -7.410 112.780 -7.090 112.820 ;
        RECT 49.860 112.780 50.100 113.390 ;
        RECT 50.480 113.380 51.060 114.010 ;
        RECT 81.010 113.950 81.320 114.020 ;
        RECT 53.300 113.870 53.770 113.930 ;
        RECT 78.200 113.880 78.490 113.890 ;
        RECT 78.200 113.870 78.500 113.880 ;
        RECT 81.010 113.870 83.340 113.950 ;
        RECT 88.730 113.870 89.180 113.890 ;
        RECT 53.300 113.440 112.090 113.870 ;
        RECT 54.240 113.430 54.550 113.440 ;
        RECT 78.200 113.430 78.500 113.440 ;
        RECT 54.240 113.240 63.980 113.430 ;
        RECT 78.200 113.410 78.490 113.430 ;
        RECT 54.240 113.120 54.550 113.240 ;
        RECT -11.180 112.570 -10.860 112.620 ;
        RECT -10.480 112.570 -10.160 112.650 ;
        RECT 81.950 112.610 82.270 112.870 ;
        RECT 198.760 112.820 204.470 118.460 ;
        RECT 198.320 112.780 204.470 112.820 ;
        RECT 88.580 112.770 204.470 112.780 ;
        RECT 88.230 112.760 204.470 112.770 ;
        RECT 74.380 112.580 74.680 112.600 ;
        RECT 81.990 112.590 83.170 112.610 ;
        RECT 81.990 112.580 83.210 112.590 ;
        RECT 87.670 112.580 204.470 112.760 ;
        RECT -11.180 112.400 -10.160 112.570 ;
        RECT -11.180 112.360 -10.860 112.400 ;
        RECT -10.480 112.330 -10.160 112.400 ;
        RECT 53.520 112.550 53.840 112.580 ;
        RECT 53.520 112.320 63.980 112.550 ;
        RECT 74.370 112.320 204.470 112.580 ;
        RECT 74.370 112.160 204.310 112.320 ;
        RECT -8.920 112.070 -8.610 112.160 ;
        RECT 74.380 112.140 74.680 112.160 ;
        RECT -7.410 112.070 -7.090 112.120 ;
        RECT -8.920 111.900 -7.030 112.070 ;
        RECT 81.950 112.010 82.270 112.160 ;
        RECT -8.920 111.830 -8.610 111.900 ;
        RECT -7.410 111.860 -7.090 111.900 ;
        RECT 87.670 111.820 204.310 112.160 ;
        RECT -11.210 111.650 -10.890 111.700 ;
        RECT -10.480 111.650 -10.160 111.730 ;
        RECT -11.210 111.480 -10.160 111.650 ;
        RECT 80.620 111.630 80.930 111.640 ;
        RECT 80.050 111.620 80.930 111.630 ;
        RECT -11.210 111.440 -10.890 111.480 ;
        RECT -10.480 111.410 -10.160 111.480 ;
        RECT 79.980 111.380 80.930 111.620 ;
        RECT 80.620 111.310 80.930 111.380 ;
        RECT 81.590 111.310 81.900 111.360 ;
        RECT 83.840 111.310 84.150 111.410 ;
        RECT -130.950 110.800 -19.470 111.200 ;
        RECT -8.920 111.150 -8.610 111.240 ;
        RECT -7.440 111.150 -7.120 111.200 ;
        RECT 81.010 111.190 81.320 111.260 ;
        RECT 81.590 111.190 84.150 111.310 ;
        RECT -8.920 110.980 -7.030 111.150 ;
        RECT 81.010 111.080 84.150 111.190 ;
        RECT 81.010 110.980 83.340 111.080 ;
        RECT -8.920 110.910 -8.610 110.980 ;
        RECT -7.440 110.940 -7.120 110.980 ;
        RECT 81.010 110.930 81.320 110.980 ;
        RECT -130.950 110.190 -26.160 110.800 ;
        RECT -11.200 110.730 -10.880 110.780 ;
        RECT -10.480 110.730 -10.160 110.810 ;
        RECT 80.770 110.770 81.080 110.810 ;
        RECT -11.200 110.560 -10.160 110.730 ;
        RECT 80.590 110.630 81.310 110.770 ;
        RECT 81.540 110.630 81.850 110.710 ;
        RECT -11.200 110.520 -10.880 110.560 ;
        RECT -10.480 110.490 -10.160 110.560 ;
        RECT 59.760 110.340 68.910 110.570 ;
        RECT 80.590 110.520 81.850 110.630 ;
        RECT 80.770 110.480 81.850 110.520 ;
        RECT 81.040 110.420 81.850 110.480 ;
        RECT 81.040 110.410 81.310 110.420 ;
        RECT 81.540 110.380 81.850 110.420 ;
        RECT 87.730 110.420 204.310 111.820 ;
        RECT 87.730 110.390 88.630 110.420 ;
        RECT 68.620 110.240 68.910 110.340 ;
        RECT 78.410 110.240 79.530 110.250 ;
        RECT 79.650 110.240 79.960 110.270 ;
        RECT -130.950 110.030 -27.430 110.190 ;
        RECT 68.620 110.100 81.170 110.240 ;
        RECT 68.620 110.040 83.340 110.100 ;
        RECT 68.620 110.030 68.910 110.040 ;
        RECT -144.230 101.370 -142.700 101.450 ;
        RECT -144.230 100.360 -142.190 101.370 ;
        RECT -147.240 99.720 -142.190 100.360 ;
        RECT -144.230 99.440 -142.190 99.720 ;
        RECT -144.230 98.820 -142.120 99.440 ;
        RECT -144.230 72.860 -142.830 98.820 ;
        RECT -130.950 89.920 -128.870 110.030 ;
        RECT 71.810 109.940 83.340 110.040 ;
        RECT 79.180 109.910 79.650 109.940 ;
        RECT 80.750 109.920 83.340 109.940 ;
        RECT 80.750 109.910 81.170 109.920 ;
        RECT 81.110 109.840 81.310 109.850 ;
        RECT 81.110 109.830 81.330 109.840 ;
        RECT 81.540 109.830 81.850 109.870 ;
        RECT -11.850 109.720 -11.530 109.760 ;
        RECT -10.200 109.720 -9.880 109.780 ;
        RECT 81.110 109.760 81.850 109.830 ;
        RECT 80.820 109.740 81.850 109.760 ;
        RECT -11.850 109.530 -9.880 109.720 ;
        RECT -11.850 109.500 -11.530 109.530 ;
        RECT -10.200 109.460 -9.880 109.530 ;
        RECT 59.760 109.620 67.970 109.740 ;
        RECT 80.770 109.620 81.850 109.740 ;
        RECT 59.760 109.520 75.910 109.620 ;
        RECT 67.750 109.420 75.910 109.520 ;
        RECT 80.770 109.500 81.330 109.620 ;
        RECT 81.540 109.540 81.850 109.620 ;
        RECT 80.770 109.490 81.240 109.500 ;
        RECT -11.890 108.760 -11.570 108.800 ;
        RECT -10.200 108.760 -9.880 108.820 ;
        RECT -11.890 108.570 -9.880 108.760 ;
        RECT -11.890 108.540 -11.570 108.570 ;
        RECT -10.200 108.500 -9.880 108.570 ;
        RECT 67.750 108.740 67.970 109.420 ;
        RECT 70.370 109.260 70.830 109.390 ;
        RECT 75.690 109.260 75.910 109.420 ;
        RECT 80.100 109.260 80.420 109.300 ;
        RECT 81.110 109.260 81.430 109.290 ;
        RECT 70.370 109.060 78.150 109.260 ;
        RECT 80.050 109.170 83.810 109.260 ;
        RECT 83.890 109.170 84.200 109.190 ;
        RECT 80.050 109.060 84.510 109.170 ;
        RECT 70.370 108.940 70.830 109.060 ;
        RECT 74.510 108.740 74.730 108.750 ;
        RECT 67.750 108.610 74.760 108.740 ;
        RECT 75.690 108.700 75.910 109.060 ;
        RECT 77.830 108.970 78.150 109.060 ;
        RECT 80.100 109.040 80.420 109.060 ;
        RECT 81.110 109.030 81.430 109.060 ;
        RECT 80.380 108.950 80.690 108.990 ;
        RECT 80.060 108.940 80.720 108.950 ;
        RECT 81.590 108.940 84.510 109.060 ;
        RECT 80.060 108.710 81.160 108.940 ;
        RECT 81.590 108.890 81.900 108.940 ;
        RECT 75.660 108.660 75.910 108.700 ;
        RECT 75.660 108.610 75.920 108.660 ;
        RECT 77.830 108.610 78.150 108.700 ;
        RECT 80.380 108.660 80.690 108.710 ;
        RECT 80.100 108.610 80.420 108.630 ;
        RECT 81.110 108.610 81.430 108.640 ;
        RECT 83.610 108.610 83.810 108.940 ;
        RECT 83.890 108.860 84.200 108.940 ;
        RECT 67.750 108.490 78.150 108.610 ;
        RECT 51.830 107.980 52.150 108.240 ;
        RECT 51.870 107.960 53.050 107.980 ;
        RECT -11.850 107.800 -11.530 107.840 ;
        RECT -10.200 107.800 -9.880 107.860 ;
        RECT -11.850 107.610 -9.880 107.800 ;
        RECT 51.870 107.700 53.090 107.960 ;
        RECT 67.750 107.760 67.970 108.490 ;
        RECT 71.380 108.410 78.150 108.490 ;
        RECT 80.050 108.410 83.810 108.610 ;
        RECT 71.380 108.290 71.740 108.410 ;
        RECT 51.870 107.640 53.050 107.700 ;
        RECT -11.850 107.580 -11.530 107.610 ;
        RECT -10.200 107.540 -9.880 107.610 ;
        RECT 51.830 107.630 53.050 107.640 ;
        RECT 67.750 107.630 71.440 107.760 ;
        RECT 74.470 107.630 74.760 108.410 ;
        RECT 75.660 108.020 75.920 108.410 ;
        RECT 80.100 108.370 80.420 108.410 ;
        RECT 81.110 108.380 81.430 108.410 ;
        RECT 81.590 108.340 81.900 108.400 ;
        RECT 83.610 108.340 83.810 108.410 ;
        RECT 83.880 108.340 84.190 108.470 ;
        RECT 81.590 108.120 84.510 108.340 ;
        RECT 81.590 108.070 81.900 108.120 ;
        RECT 75.660 107.810 79.790 108.020 ;
        RECT 79.180 107.640 79.490 107.760 ;
        RECT 79.580 107.670 79.790 107.810 ;
        RECT 80.750 107.670 81.060 107.760 ;
        RECT 81.540 107.670 81.850 107.750 ;
        RECT 78.410 107.630 79.530 107.640 ;
        RECT 79.580 107.630 81.850 107.670 ;
        RECT 51.830 107.380 52.150 107.630 ;
        RECT 67.750 107.460 81.850 107.630 ;
        RECT 67.750 107.430 81.060 107.460 ;
        RECT 67.750 107.420 69.350 107.430 ;
        RECT 32.470 107.330 32.780 107.340 ;
        RECT 32.460 107.270 32.790 107.330 ;
        RECT 32.110 107.220 32.790 107.270 ;
        RECT 28.880 107.140 32.790 107.220 ;
        RECT 34.110 107.190 36.060 107.330 ;
        RECT 71.210 107.220 71.440 107.430 ;
        RECT 74.470 107.320 74.760 107.430 ;
        RECT 78.410 107.420 79.530 107.430 ;
        RECT 81.540 107.420 81.850 107.460 ;
        RECT 83.610 107.360 83.810 108.120 ;
        RECT 192.980 108.040 195.070 108.220 ;
        RECT 88.580 108.030 195.070 108.040 ;
        RECT 87.700 107.360 195.070 108.030 ;
        RECT 74.470 107.220 77.360 107.320 ;
        RECT 78.410 107.220 79.530 107.230 ;
        RECT 34.040 107.170 36.060 107.190 ;
        RECT 34.040 107.140 34.360 107.170 ;
        RECT 34.840 107.160 36.060 107.170 ;
        RECT 35.540 107.150 36.060 107.160 ;
        RECT 28.880 107.000 34.360 107.140 ;
        RECT 59.760 107.020 81.060 107.220 ;
        RECT 31.630 106.950 34.360 107.000 ;
        RECT 31.630 106.900 31.950 106.950 ;
        RECT 34.040 106.930 34.360 106.950 ;
        RECT 49.500 107.000 50.060 107.020 ;
        RECT 50.500 107.000 50.810 107.010 ;
        RECT 49.500 106.750 50.810 107.000 ;
        RECT 71.210 106.970 71.440 107.020 ;
        RECT 78.410 107.010 79.530 107.020 ;
        RECT 71.210 106.820 71.430 106.970 ;
        RECT 79.180 106.890 79.490 107.010 ;
        RECT 80.750 106.890 81.060 107.020 ;
        RECT 83.610 106.930 195.070 107.360 ;
        RECT 81.540 106.870 81.850 106.910 ;
        RECT 75.580 106.820 81.850 106.870 ;
        RECT 49.500 106.480 50.060 106.750 ;
        RECT 50.500 106.680 50.810 106.750 ;
        RECT 51.470 106.680 51.780 106.730 ;
        RECT 53.720 106.680 54.030 106.780 ;
        RECT 50.890 106.560 51.200 106.630 ;
        RECT 51.470 106.560 54.030 106.680 ;
        RECT 71.210 106.660 81.850 106.820 ;
        RECT 71.210 106.600 75.970 106.660 ;
        RECT 81.540 106.580 81.850 106.660 ;
        RECT 50.890 106.450 54.030 106.560 ;
        RECT 50.890 106.350 53.220 106.450 ;
        RECT 72.300 106.350 72.690 106.370 ;
        RECT 50.890 106.300 51.200 106.350 ;
        RECT 72.290 106.240 72.700 106.350 ;
        RECT 80.100 106.240 80.420 106.280 ;
        RECT 81.110 106.240 81.430 106.270 ;
        RECT 81.590 106.240 81.900 106.260 ;
        RECT 83.610 106.240 83.810 106.930 ;
        RECT 50.650 106.140 50.960 106.180 ;
        RECT 50.470 106.000 51.190 106.140 ;
        RECT 51.420 106.000 51.730 106.080 ;
        RECT 50.470 105.890 51.730 106.000 ;
        RECT 72.290 106.040 78.150 106.240 ;
        RECT 80.050 106.220 83.810 106.240 ;
        RECT 80.050 106.180 84.110 106.220 ;
        RECT 80.050 106.040 84.300 106.180 ;
        RECT 72.290 105.950 72.700 106.040 ;
        RECT 77.830 105.950 78.150 106.040 ;
        RECT 80.100 106.020 80.420 106.040 ;
        RECT 81.020 106.010 81.430 106.040 ;
        RECT 81.020 105.950 81.340 106.010 ;
        RECT 50.650 105.850 51.730 105.890 ;
        RECT 50.920 105.790 51.730 105.850 ;
        RECT 50.920 105.780 51.190 105.790 ;
        RECT 51.420 105.750 51.730 105.790 ;
        RECT 64.830 105.800 81.340 105.950 ;
        RECT 81.590 105.950 84.300 106.040 ;
        RECT 87.700 105.950 195.070 106.930 ;
        RECT 81.590 105.930 81.900 105.950 ;
        RECT 83.610 105.890 84.110 105.950 ;
        RECT 87.700 105.940 88.600 105.950 ;
        RECT 64.830 105.650 65.150 105.800 ;
        RECT 70.630 105.650 70.950 105.800 ;
        RECT 73.120 105.650 73.520 105.660 ;
        RECT 49.530 105.500 49.840 105.640 ;
        RECT 35.650 105.460 45.790 105.490 ;
        RECT 49.180 105.460 49.840 105.500 ;
        RECT 50.740 105.470 51.050 105.610 ;
        RECT 73.100 105.590 73.540 105.650 ;
        RECT 77.830 105.590 78.150 105.680 ;
        RECT 80.100 105.590 80.420 105.610 ;
        RECT 81.110 105.590 81.430 105.620 ;
        RECT 83.610 105.590 83.810 105.890 ;
        RECT 50.740 105.460 53.220 105.470 ;
        RECT 35.650 105.310 53.220 105.460 ;
        RECT 73.100 105.390 78.150 105.590 ;
        RECT 80.050 105.470 83.810 105.590 ;
        RECT 80.050 105.390 83.780 105.470 ;
        RECT 73.120 105.380 73.520 105.390 ;
        RECT 80.100 105.350 80.420 105.390 ;
        RECT 81.110 105.360 81.430 105.390 ;
        RECT 35.650 105.270 45.790 105.310 ;
        RECT 49.180 105.280 49.530 105.310 ;
        RECT 50.740 105.290 53.220 105.310 ;
        RECT 50.740 105.280 51.050 105.290 ;
        RECT 45.570 104.070 45.790 105.270 ;
        RECT 50.990 105.210 51.190 105.220 ;
        RECT 50.990 105.200 51.210 105.210 ;
        RECT 51.420 105.200 51.730 105.240 ;
        RECT 50.990 105.130 51.730 105.200 ;
        RECT 50.700 105.110 51.730 105.130 ;
        RECT 50.650 104.990 51.730 105.110 ;
        RECT 50.650 104.870 51.210 104.990 ;
        RECT 51.420 104.910 51.730 104.990 ;
        RECT 50.650 104.860 51.120 104.870 ;
        RECT 45.540 104.030 45.790 104.070 ;
        RECT 45.540 103.390 45.800 104.030 ;
        RECT 45.540 103.180 49.670 103.390 ;
        RECT 49.460 103.040 49.670 103.180 ;
        RECT 51.420 103.040 51.730 103.120 ;
        RECT 49.460 102.830 51.730 103.040 ;
        RECT 51.420 102.790 51.730 102.830 ;
        RECT 40.480 101.320 40.800 101.330 ;
        RECT 50.920 101.320 51.250 101.460 ;
        RECT 39.940 101.170 40.250 101.180 ;
        RECT 40.480 101.170 51.250 101.320 ;
        RECT 37.780 101.160 51.250 101.170 ;
        RECT 37.780 100.990 47.860 101.160 ;
        RECT 39.940 100.850 40.250 100.990 ;
        RECT 39.940 99.590 40.250 99.610 ;
        RECT 40.620 99.590 43.470 99.670 ;
        RECT 57.510 99.590 60.340 99.670 ;
        RECT 60.710 99.590 61.020 99.610 ;
        RECT 37.780 99.570 47.840 99.590 ;
        RECT 53.120 99.570 63.180 99.590 ;
        RECT 37.780 99.420 63.180 99.570 ;
        RECT 37.780 99.410 40.340 99.420 ;
        RECT 39.940 99.280 40.250 99.410 ;
        RECT 40.620 99.370 41.040 99.420 ;
        RECT 43.030 99.390 57.710 99.420 ;
        RECT 60.020 99.370 60.340 99.420 ;
        RECT 60.620 99.410 63.180 99.420 ;
        RECT 60.710 99.280 61.020 99.410 ;
        RECT 40.850 99.040 41.170 99.120 ;
        RECT 44.780 99.040 45.100 99.050 ;
        RECT 40.850 98.860 45.100 99.040 ;
        RECT 40.850 98.800 41.170 98.860 ;
        RECT 44.780 98.790 45.100 98.860 ;
        RECT 55.860 99.040 56.180 99.050 ;
        RECT 59.790 99.040 60.110 99.120 ;
        RECT 55.860 98.860 60.110 99.040 ;
        RECT 55.860 98.790 56.180 98.860 ;
        RECT 59.790 98.800 60.110 98.860 ;
        RECT 87.700 97.760 88.600 97.770 ;
        RECT 64.980 96.740 65.580 96.800 ;
        RECT 87.700 96.740 186.850 97.760 ;
        RECT 64.980 96.270 186.850 96.740 ;
        RECT 64.980 96.220 65.580 96.270 ;
        RECT 87.700 95.680 186.850 96.270 ;
        RECT 88.580 95.670 186.850 95.680 ;
        RECT -11.890 92.770 -11.580 92.790 ;
        RECT -11.230 92.770 -10.920 92.790 ;
        RECT 27.240 92.780 27.550 92.800 ;
        RECT -11.890 92.300 -4.570 92.770 ;
        RECT -11.890 92.280 -11.580 92.300 ;
        RECT -11.230 92.280 -10.920 92.300 ;
        RECT -5.040 91.620 -4.570 92.300 ;
        RECT 21.730 92.630 22.040 92.650 ;
        RECT 25.080 92.630 35.160 92.780 ;
        RECT 59.370 92.630 59.820 92.660 ;
        RECT 21.730 92.220 59.820 92.630 ;
        RECT 21.730 92.200 22.040 92.220 ;
        RECT 59.370 92.200 59.820 92.220 ;
        RECT 87.730 92.560 88.630 92.590 ;
        RECT 27.240 91.780 27.550 91.910 ;
        RECT 35.040 91.780 35.180 91.800 ;
        RECT 25.070 91.620 35.180 91.780 ;
        RECT 87.730 91.620 182.760 92.560 ;
        RECT -13.220 91.490 -12.960 91.560 ;
        RECT -11.170 91.490 -10.850 91.510 ;
        RECT -9.410 91.490 -9.080 91.530 ;
        RECT -13.220 91.300 -9.080 91.490 ;
        RECT -13.220 91.240 -12.960 91.300 ;
        RECT -11.170 91.250 -10.850 91.300 ;
        RECT -9.410 91.260 -9.080 91.300 ;
        RECT -5.040 91.150 182.760 91.620 ;
        RECT -13.770 91.090 -13.450 91.130 ;
        RECT -11.830 91.090 -11.510 91.150 ;
        RECT -8.910 91.090 -8.590 91.130 ;
        RECT -13.770 90.900 -8.590 91.090 ;
        RECT 27.240 91.030 27.550 91.150 ;
        RECT 63.890 91.030 64.460 91.150 ;
        RECT -13.770 90.870 -13.450 90.900 ;
        RECT -11.830 90.890 -11.510 90.900 ;
        RECT -8.910 90.870 -8.590 90.900 ;
        RECT -10.430 90.510 -10.120 90.580 ;
        RECT -7.430 90.530 -7.130 90.550 ;
        RECT -7.440 90.510 -7.120 90.530 ;
        RECT -10.430 90.300 -7.120 90.510 ;
        RECT 87.730 90.500 182.760 91.150 ;
        RECT 88.580 90.470 182.760 90.500 ;
        RECT -10.430 90.250 -10.120 90.300 ;
        RECT -9.660 90.290 -7.120 90.300 ;
        RECT -11.600 90.070 -11.290 90.140 ;
        RECT -9.660 90.070 -9.440 90.290 ;
        RECT -7.440 90.270 -7.120 90.290 ;
        RECT -7.430 90.250 -7.130 90.270 ;
        RECT -131.020 86.550 -128.680 89.920 ;
        RECT -11.600 89.850 -9.440 90.070 ;
        RECT -11.600 89.810 -11.290 89.850 ;
        RECT 27.240 89.770 27.550 89.790 ;
        RECT 25.080 89.610 35.150 89.770 ;
        RECT 25.080 89.600 35.140 89.610 ;
        RECT 25.080 89.590 27.640 89.600 ;
        RECT 27.240 89.460 27.550 89.590 ;
        RECT 30.500 89.580 30.820 89.600 ;
        RECT -9.920 89.350 -9.600 89.410 ;
        RECT -8.050 89.380 -7.760 89.400 ;
        RECT 30.500 89.390 38.420 89.580 ;
        RECT 38.580 89.390 38.890 89.430 ;
        RECT -9.920 89.340 -9.440 89.350 ;
        RECT -8.060 89.340 -7.740 89.380 ;
        RECT 30.500 89.370 38.890 89.390 ;
        RECT 30.500 89.340 30.820 89.370 ;
        RECT 31.630 89.340 34.360 89.370 ;
        RECT -9.920 89.150 -7.740 89.340 ;
        RECT 31.630 89.290 36.060 89.340 ;
        RECT 31.630 89.210 31.950 89.290 ;
        RECT 34.040 89.240 36.060 89.290 ;
        RECT 34.080 89.170 36.060 89.240 ;
        RECT 38.210 89.180 38.890 89.370 ;
        RECT 35.540 89.160 36.060 89.170 ;
        RECT -9.920 89.140 -9.440 89.150 ;
        RECT -9.920 89.090 -9.600 89.140 ;
        RECT -8.060 89.120 -7.740 89.150 ;
        RECT -8.050 89.100 -7.760 89.120 ;
        RECT 38.580 89.100 38.890 89.180 ;
        RECT 27.230 88.950 27.380 88.960 ;
        RECT 26.210 88.910 27.380 88.950 ;
        RECT 26.210 88.800 27.550 88.910 ;
        RECT 26.150 88.780 26.430 88.800 ;
        RECT 27.230 88.790 27.550 88.800 ;
        RECT 30.390 88.790 30.870 89.000 ;
        RECT 27.230 88.780 35.150 88.790 ;
        RECT -12.750 88.740 -12.430 88.760 ;
        RECT -12.970 88.520 -12.430 88.740 ;
        RECT 25.080 88.620 35.150 88.780 ;
        RECT 25.080 88.600 27.640 88.620 ;
        RECT -12.750 88.500 -12.430 88.520 ;
        RECT 26.150 88.470 26.430 88.600 ;
        RECT 27.230 88.580 27.550 88.600 ;
        RECT 27.230 88.450 27.380 88.580 ;
        RECT 30.480 88.450 30.800 88.550 ;
        RECT 32.820 88.530 34.360 88.620 ;
        RECT 27.230 88.350 30.800 88.450 ;
        RECT 25.080 88.290 30.800 88.350 ;
        RECT -10.000 88.160 -9.680 88.280 ;
        RECT 25.080 88.180 27.650 88.290 ;
        RECT 25.080 88.170 27.550 88.180 ;
        RECT -12.970 87.960 -9.680 88.160 ;
        RECT 27.240 88.050 27.550 88.170 ;
        RECT 27.210 88.030 27.550 88.050 ;
        RECT -12.970 87.950 -9.990 87.960 ;
        RECT 27.210 87.790 27.530 88.030 ;
        RECT 30.530 87.830 30.870 87.900 ;
        RECT 27.280 87.780 27.450 87.790 ;
        RECT -12.970 87.740 -9.990 87.760 ;
        RECT -12.970 87.550 -9.670 87.740 ;
        RECT 30.390 87.600 30.870 87.830 ;
        RECT -9.990 87.420 -9.670 87.550 ;
        RECT 88.580 87.510 178.630 87.520 ;
        RECT 30.440 87.310 30.670 87.320 ;
        RECT 31.630 87.310 31.950 87.390 ;
        RECT 34.110 87.360 36.060 87.500 ;
        RECT 34.040 87.340 36.060 87.360 ;
        RECT 34.040 87.310 34.360 87.340 ;
        RECT 34.840 87.330 36.060 87.340 ;
        RECT 35.540 87.320 36.060 87.330 ;
        RECT 30.440 87.280 38.010 87.310 ;
        RECT -13.740 87.220 -13.450 87.230 ;
        RECT -13.750 87.200 -13.430 87.220 ;
        RECT -12.750 87.200 -12.430 87.210 ;
        RECT -13.750 86.980 -12.430 87.200 ;
        RECT 30.440 87.110 38.070 87.280 ;
        RECT 38.580 87.110 38.890 87.190 ;
        RECT -13.750 86.960 -13.430 86.980 ;
        RECT -13.740 86.940 -13.450 86.960 ;
        RECT -12.750 86.950 -12.430 86.980 ;
        RECT 27.190 87.010 27.510 87.040 ;
        RECT 30.440 87.010 30.680 87.110 ;
        RECT 31.630 87.070 31.950 87.110 ;
        RECT 34.040 87.100 34.360 87.110 ;
        RECT 27.190 86.830 30.680 87.010 ;
        RECT 37.880 86.910 38.890 87.110 ;
        RECT 38.480 86.900 38.890 86.910 ;
        RECT 38.580 86.860 38.890 86.900 ;
        RECT 27.190 86.810 30.600 86.830 ;
        RECT -9.940 86.740 -9.620 86.790 ;
        RECT -8.480 86.740 -8.160 86.790 ;
        RECT 27.190 86.780 27.510 86.810 ;
        RECT -130.950 85.680 -128.870 86.550 ;
        RECT -9.940 86.530 -8.160 86.740 ;
        RECT -9.940 86.470 -9.620 86.530 ;
        RECT -8.480 86.490 -8.160 86.530 ;
        RECT 30.480 86.630 30.800 86.670 ;
        RECT 30.480 86.610 38.030 86.630 ;
        RECT 38.580 86.620 38.890 86.660 ;
        RECT 38.480 86.610 38.890 86.620 ;
        RECT 30.480 86.410 38.890 86.610 ;
        RECT 30.580 86.400 30.900 86.410 ;
        RECT 31.630 86.360 34.360 86.410 ;
        RECT 31.630 86.280 31.950 86.360 ;
        RECT 34.040 86.350 34.360 86.360 ;
        RECT 34.040 86.310 36.060 86.350 ;
        RECT 38.580 86.330 38.890 86.410 ;
        RECT 62.770 86.380 63.320 86.390 ;
        RECT 62.770 86.360 63.330 86.380 ;
        RECT 87.700 86.360 178.630 87.510 ;
        RECT 34.150 86.190 36.060 86.310 ;
        RECT 34.870 86.170 36.060 86.190 ;
        RECT 26.760 85.950 27.080 86.000 ;
        RECT 26.760 85.680 27.370 85.950 ;
        RECT 30.390 85.840 30.870 86.070 ;
        RECT 62.770 85.890 178.630 86.360 ;
        RECT 62.770 85.880 63.330 85.890 ;
        RECT 62.770 85.860 63.320 85.880 ;
        RECT 30.530 85.770 30.870 85.840 ;
        RECT 27.170 85.450 27.370 85.680 ;
        RECT 30.320 85.450 30.640 85.490 ;
        RECT 27.170 85.250 30.720 85.450 ;
        RECT 87.700 85.430 178.630 85.890 ;
        RECT 87.700 85.420 88.600 85.430 ;
        RECT 30.320 85.230 30.640 85.250 ;
        RECT 109.550 84.210 114.080 84.290 ;
        RECT 88.860 84.190 114.150 84.210 ;
        RECT -12.640 84.160 -12.330 84.170 ;
        RECT -11.550 84.160 -11.240 84.170 ;
        RECT -13.960 84.150 -11.240 84.160 ;
        RECT -14.190 83.840 -11.240 84.150 ;
        RECT -14.190 83.830 -11.250 83.840 ;
        RECT -56.240 82.220 -55.640 82.270 ;
        RECT -56.240 82.210 -26.900 82.220 ;
        RECT -14.190 82.210 -13.840 83.830 ;
        RECT 19.550 83.580 19.870 83.630 ;
        RECT 26.160 83.580 26.480 83.680 ;
        RECT -13.190 83.480 -12.880 83.490 ;
        RECT -12.090 83.480 -11.780 83.490 ;
        RECT -10.990 83.480 -10.680 83.490 ;
        RECT -13.220 83.160 -10.060 83.480 ;
        RECT 19.550 83.420 26.480 83.580 ;
        RECT 19.550 83.370 19.870 83.420 ;
        RECT 26.160 83.400 26.480 83.420 ;
        RECT 67.960 83.550 68.520 83.620 ;
        RECT 80.680 83.550 81.360 83.610 ;
        RECT 88.210 83.550 114.150 84.190 ;
        RECT 26.750 83.340 27.030 83.350 ;
        RECT 19.020 83.290 19.350 83.310 ;
        RECT -10.380 82.210 -10.060 83.160 ;
        RECT 19.010 83.210 19.360 83.290 ;
        RECT 24.760 83.210 25.080 83.270 ;
        RECT 26.730 83.250 27.050 83.340 ;
        RECT 28.970 83.250 29.290 83.280 ;
        RECT 19.010 83.050 25.080 83.210 ;
        RECT 26.700 83.090 29.290 83.250 ;
        RECT 67.960 83.140 114.150 83.550 ;
        RECT 67.960 83.090 68.520 83.140 ;
        RECT 26.730 83.080 27.050 83.090 ;
        RECT 26.750 83.070 27.030 83.080 ;
        RECT 19.010 82.980 19.370 83.050 ;
        RECT 24.760 83.000 25.080 83.050 ;
        RECT 28.970 83.020 29.290 83.090 ;
        RECT 80.680 83.080 81.360 83.140 ;
        RECT 88.210 83.060 114.150 83.140 ;
        RECT 88.210 83.040 88.870 83.060 ;
        RECT 109.550 83.040 114.080 83.060 ;
        RECT 28.990 83.010 29.270 83.020 ;
        RECT 19.260 82.950 19.370 82.980 ;
        RECT 14.590 82.590 14.920 82.830 ;
        RECT 20.450 82.720 20.750 82.730 ;
        RECT 20.440 82.590 20.760 82.720 ;
        RECT 30.980 82.590 31.260 82.890 ;
        RECT 35.010 82.590 35.310 82.870 ;
        RECT 14.590 82.570 35.310 82.590 ;
        RECT 14.590 82.540 35.300 82.570 ;
        RECT 14.590 82.430 35.240 82.540 ;
        RECT 18.400 82.210 18.840 82.220 ;
        RECT -56.240 82.200 18.840 82.210 ;
        RECT -56.240 81.790 18.860 82.200 ;
        RECT -56.240 81.780 -26.900 81.790 ;
        RECT -56.240 81.710 -55.640 81.780 ;
        RECT -14.190 81.390 -13.840 81.790 ;
        RECT -52.810 81.240 -52.350 81.250 ;
        RECT -14.190 81.240 -11.240 81.390 ;
        RECT -10.380 81.240 -10.060 81.790 ;
        RECT 11.550 81.780 12.030 81.790 ;
        RECT 18.380 81.780 18.860 81.790 ;
        RECT 18.400 81.770 18.840 81.780 ;
        RECT 27.770 81.740 28.150 82.130 ;
        RECT 28.920 81.700 29.320 82.040 ;
        RECT 88.900 82.000 174.390 82.010 ;
        RECT -52.810 80.820 15.040 81.240 ;
        RECT -52.810 80.800 -26.940 80.820 ;
        RECT -52.810 80.780 -52.350 80.800 ;
        RECT -14.190 80.190 -13.840 80.820 ;
        RECT -14.190 80.060 -13.810 80.190 ;
        RECT -14.190 80.020 -13.440 80.060 ;
        RECT -12.640 80.020 -12.330 80.040 ;
        RECT -14.190 79.720 -11.240 80.020 ;
        RECT -12.640 79.710 -12.330 79.720 ;
        RECT -11.550 79.690 -11.240 79.720 ;
        RECT -13.190 79.340 -12.880 79.350 ;
        RECT -10.380 79.340 -10.060 80.820 ;
        RECT -3.890 80.320 -3.060 80.820 ;
        RECT 19.070 80.700 19.450 81.080 ;
        RECT 61.720 81.060 62.320 81.110 ;
        RECT 88.130 81.060 174.390 82.000 ;
        RECT 61.720 80.590 174.390 81.060 ;
        RECT 61.720 80.550 62.320 80.590 ;
        RECT 88.130 79.920 174.390 80.590 ;
        RECT 88.150 79.910 88.920 79.920 ;
        RECT -13.210 79.010 -10.060 79.340 ;
        RECT -13.210 79.000 -10.150 79.010 ;
        RECT -10.300 78.800 -10.010 78.820 ;
        RECT -8.070 78.800 -7.760 78.820 ;
        RECT -10.310 78.440 -7.760 78.800 ;
        RECT -10.300 78.420 -10.010 78.440 ;
        RECT -8.070 78.420 -7.760 78.440 ;
        RECT 28.480 77.930 31.540 77.940 ;
        RECT 28.390 77.910 31.540 77.930 ;
        RECT 18.670 77.900 21.730 77.910 ;
        RECT 18.580 77.570 21.730 77.900 ;
        RECT 25.510 77.600 31.540 77.910 ;
        RECT 35.320 77.930 38.380 77.940 ;
        RECT 35.320 77.600 38.470 77.930 ;
        RECT 25.510 77.570 28.710 77.600 ;
        RECT 31.210 77.590 31.520 77.600 ;
        RECT 35.340 77.590 35.650 77.600 ;
        RECT -12.600 76.600 -12.290 76.610 ;
        RECT -11.510 76.600 -11.200 76.610 ;
        RECT -13.920 76.590 -11.200 76.600 ;
        RECT -14.150 76.280 -11.200 76.590 ;
        RECT -14.150 76.270 -11.210 76.280 ;
        RECT -14.150 73.830 -13.800 76.270 ;
        RECT -13.150 75.920 -12.840 75.930 ;
        RECT -12.050 75.920 -11.740 75.930 ;
        RECT -10.950 75.920 -10.640 75.930 ;
        RECT -13.180 75.600 -10.020 75.920 ;
        RECT -10.340 75.140 -10.020 75.600 ;
        RECT -7.440 75.140 -7.160 75.150 ;
        RECT -11.030 74.810 -7.140 75.140 ;
        RECT 18.580 75.120 18.900 77.570 ;
        RECT 21.400 77.560 21.710 77.570 ;
        RECT 25.530 77.560 25.840 77.570 ;
        RECT 19.760 77.190 20.070 77.220 ;
        RECT 20.850 77.190 21.160 77.200 ;
        RECT 26.080 77.190 26.390 77.200 ;
        RECT 27.170 77.190 27.480 77.220 ;
        RECT 19.760 76.890 22.710 77.190 ;
        RECT 20.850 76.870 21.160 76.890 ;
        RECT 21.960 76.850 22.710 76.890 ;
        RECT 22.330 76.720 22.710 76.850 ;
        RECT 22.360 75.850 22.710 76.720 ;
        RECT 24.530 76.890 27.480 77.190 ;
        RECT 24.530 76.850 25.280 76.890 ;
        RECT 26.080 76.870 26.390 76.890 ;
        RECT 24.530 76.720 24.910 76.850 ;
        RECT 24.530 76.290 24.880 76.720 ;
        RECT 28.340 76.290 28.710 77.570 ;
        RECT 29.570 77.220 29.880 77.250 ;
        RECT 30.660 77.220 30.970 77.230 ;
        RECT 35.890 77.220 36.200 77.230 ;
        RECT 36.980 77.220 37.290 77.250 ;
        RECT 29.570 76.920 32.520 77.220 ;
        RECT 30.660 76.900 30.970 76.920 ;
        RECT 31.770 76.880 32.520 76.920 ;
        RECT 32.140 76.750 32.520 76.880 ;
        RECT 32.170 76.290 32.520 76.750 ;
        RECT 34.340 76.920 37.290 77.220 ;
        RECT 34.340 76.880 35.090 76.920 ;
        RECT 35.890 76.900 36.200 76.920 ;
        RECT 34.340 76.750 34.720 76.880 ;
        RECT 23.090 76.260 33.990 76.290 ;
        RECT 23.080 76.010 33.990 76.260 ;
        RECT 23.080 75.980 23.420 76.010 ;
        RECT 23.820 76.000 24.160 76.010 ;
        RECT 19.760 75.520 22.710 75.850 ;
        RECT 19.160 75.470 19.660 75.480 ;
        RECT 22.360 75.470 22.710 75.520 ;
        RECT 24.530 75.850 24.880 76.010 ;
        RECT 24.530 75.520 27.480 75.850 ;
        RECT 24.530 75.470 24.880 75.520 ;
        RECT 28.340 75.470 28.710 76.010 ;
        RECT 32.170 75.880 32.520 76.010 ;
        RECT 32.890 75.980 33.230 76.010 ;
        RECT 29.570 75.550 32.520 75.880 ;
        RECT 32.170 75.470 32.520 75.550 ;
        RECT 34.340 75.880 34.690 76.750 ;
        RECT 34.340 75.550 37.290 75.880 ;
        RECT 34.340 75.470 34.690 75.550 ;
        RECT 38.150 75.470 38.470 77.600 ;
        RECT 41.060 77.910 44.120 77.920 ;
        RECT 41.060 77.580 44.210 77.910 ;
        RECT 41.080 77.570 41.390 77.580 ;
        RECT 41.630 77.200 41.940 77.210 ;
        RECT 42.720 77.200 43.030 77.230 ;
        RECT 40.080 76.900 43.030 77.200 ;
        RECT 40.080 76.860 40.830 76.900 ;
        RECT 41.630 76.880 41.940 76.900 ;
        RECT 40.080 76.730 40.460 76.860 ;
        RECT 40.080 75.860 40.430 76.730 ;
        RECT 40.080 75.530 43.030 75.860 ;
        RECT 40.080 75.470 40.430 75.530 ;
        RECT 43.890 75.470 44.210 77.580 ;
        RECT 65.090 75.470 65.650 75.490 ;
        RECT 19.160 75.120 65.650 75.470 ;
        RECT 18.580 75.010 65.650 75.120 ;
        RECT -10.340 74.560 -10.020 74.810 ;
        RECT -7.440 74.790 -7.160 74.810 ;
        RECT 18.580 74.790 21.740 75.010 ;
        RECT -13.180 74.230 -10.020 74.560 ;
        RECT -14.150 73.500 -11.200 73.830 ;
        RECT -14.860 73.460 -14.510 73.490 ;
        RECT -14.150 73.460 -13.800 73.500 ;
        RECT -10.340 73.460 -10.020 74.230 ;
        RECT 18.580 73.750 18.900 74.790 ;
        RECT -8.480 73.480 -8.150 73.520 ;
        RECT -8.490 73.460 -8.140 73.480 ;
        RECT -14.860 73.200 -4.830 73.460 ;
        RECT 18.580 73.430 21.740 73.750 ;
        RECT 19.200 73.420 19.510 73.430 ;
        RECT 20.300 73.420 20.610 73.430 ;
        RECT 21.400 73.420 21.710 73.430 ;
        RECT -14.820 73.170 -4.830 73.200 ;
        RECT -144.230 72.780 -142.700 72.860 ;
        RECT -144.230 71.770 -142.190 72.780 ;
        RECT -14.150 72.630 -13.800 73.170 ;
        RECT -10.340 72.830 -10.020 73.170 ;
        RECT -8.480 73.150 -8.150 73.170 ;
        RECT -14.150 72.500 -13.770 72.630 ;
        RECT -14.150 72.460 -13.400 72.500 ;
        RECT -11.020 72.490 -8.680 72.830 ;
        RECT -12.600 72.460 -12.290 72.480 ;
        RECT -14.150 72.160 -11.200 72.460 ;
        RECT -11.020 72.250 -8.640 72.490 ;
        RECT -11.020 72.230 -8.680 72.250 ;
        RECT -12.600 72.150 -12.290 72.160 ;
        RECT -11.510 72.130 -11.200 72.160 ;
        RECT -13.150 71.780 -12.840 71.790 ;
        RECT -10.340 71.780 -10.020 72.230 ;
        RECT -9.650 72.160 -8.990 72.230 ;
        RECT -9.620 72.150 -9.020 72.160 ;
        RECT -147.240 71.130 -142.190 71.770 ;
        RECT -13.170 71.450 -10.020 71.780 ;
        RECT -13.170 71.440 -10.110 71.450 ;
        RECT -144.230 70.850 -142.190 71.130 ;
        RECT -5.130 71.090 -4.840 73.170 ;
        RECT 22.360 73.080 22.710 75.010 ;
        RECT 19.770 73.070 22.710 73.080 ;
        RECT 19.760 72.760 22.710 73.070 ;
        RECT 24.530 73.080 24.880 75.010 ;
        RECT 25.500 74.820 31.550 75.010 ;
        RECT 25.500 74.790 28.710 74.820 ;
        RECT 28.340 74.560 28.710 74.790 ;
        RECT 32.170 74.560 32.520 75.010 ;
        RECT 34.340 74.560 34.690 75.010 ;
        RECT 35.310 74.820 38.470 75.010 ;
        RECT 38.150 74.560 38.470 74.820 ;
        RECT 40.080 74.560 40.430 75.010 ;
        RECT 41.050 74.800 44.210 75.010 ;
        RECT 65.090 74.990 65.650 75.010 ;
        RECT 43.890 74.560 44.210 74.800 ;
        RECT 27.470 74.100 64.550 74.560 ;
        RECT 27.540 74.000 28.060 74.100 ;
        RECT 28.340 73.780 28.710 74.100 ;
        RECT 28.340 73.750 31.550 73.780 ;
        RECT 25.500 73.650 31.550 73.750 ;
        RECT 32.170 73.650 32.520 74.100 ;
        RECT 34.340 73.650 34.690 74.100 ;
        RECT 38.150 73.780 38.470 74.100 ;
        RECT 35.310 73.650 38.470 73.780 ;
        RECT 40.080 73.650 40.430 74.100 ;
        RECT 43.890 73.760 44.210 74.100 ;
        RECT 63.900 74.040 64.460 74.100 ;
        RECT 41.050 73.650 44.210 73.760 ;
        RECT 25.500 73.460 63.460 73.650 ;
        RECT 25.500 73.430 28.660 73.460 ;
        RECT 25.530 73.420 25.840 73.430 ;
        RECT 26.630 73.420 26.940 73.430 ;
        RECT 27.730 73.420 28.040 73.430 ;
        RECT 28.900 73.190 63.460 73.460 ;
        RECT 28.150 73.130 28.750 73.160 ;
        RECT 28.900 73.130 29.550 73.190 ;
        RECT 24.530 73.070 27.470 73.080 ;
        RECT 24.530 72.760 27.480 73.070 ;
        RECT 19.760 72.750 22.480 72.760 ;
        RECT 24.760 72.750 27.480 72.760 ;
        RECT 19.760 72.740 20.070 72.750 ;
        RECT 20.850 72.740 21.160 72.750 ;
        RECT 26.080 72.740 26.390 72.750 ;
        RECT 27.170 72.740 27.480 72.750 ;
        RECT 28.150 73.060 29.550 73.130 ;
        RECT 32.170 73.110 32.520 73.190 ;
        RECT 29.580 73.100 32.520 73.110 ;
        RECT 28.150 72.340 28.900 73.060 ;
        RECT 29.570 72.790 32.520 73.100 ;
        RECT 34.340 73.110 34.690 73.190 ;
        RECT 34.340 73.100 37.280 73.110 ;
        RECT 34.340 72.790 37.290 73.100 ;
        RECT 29.570 72.780 32.290 72.790 ;
        RECT 34.570 72.780 37.290 72.790 ;
        RECT 29.570 72.770 29.880 72.780 ;
        RECT 30.660 72.770 30.970 72.780 ;
        RECT 35.890 72.770 36.200 72.780 ;
        RECT 36.980 72.770 37.290 72.780 ;
        RECT 28.290 72.310 28.900 72.340 ;
        RECT 37.350 72.710 37.870 72.730 ;
        RECT 38.110 72.710 38.710 73.160 ;
        RECT 40.080 73.090 40.430 73.190 ;
        RECT 62.770 73.170 63.330 73.190 ;
        RECT 40.080 73.080 43.020 73.090 ;
        RECT 40.080 72.770 43.030 73.080 ;
        RECT 40.310 72.760 43.030 72.770 ;
        RECT 41.630 72.750 41.940 72.760 ;
        RECT 42.720 72.750 43.030 72.760 ;
        RECT 43.850 72.710 44.450 73.140 ;
        RECT 61.840 72.710 62.400 72.720 ;
        RECT 37.350 72.250 62.490 72.710 ;
        RECT 37.350 72.200 37.880 72.250 ;
        RECT 37.350 72.150 37.870 72.200 ;
        RECT 11.290 71.090 11.610 71.110 ;
        RECT 67.290 71.090 68.450 71.120 ;
        RECT -144.230 70.230 -142.120 70.850 ;
        RECT -144.230 44.270 -142.830 70.230 ;
        RECT -5.320 69.970 68.450 71.090 ;
        RECT 11.290 69.950 11.610 69.970 ;
        RECT 22.660 69.890 24.580 69.970 ;
        RECT 32.470 69.860 34.400 69.970 ;
        RECT 67.290 69.940 68.450 69.970 ;
        RECT 71.130 67.790 71.330 67.800 ;
        RECT 74.850 67.790 75.170 67.840 ;
        RECT 71.130 67.640 75.170 67.790 ;
        RECT -25.790 66.640 -25.290 66.750 ;
        RECT 43.180 66.670 43.570 66.680 ;
        RECT 43.170 66.640 43.570 66.670 ;
        RECT -25.790 66.360 43.570 66.640 ;
        RECT -25.790 66.280 -25.290 66.360 ;
        RECT 43.170 66.340 43.570 66.360 ;
        RECT 43.180 66.330 43.570 66.340 ;
        RECT 70.450 65.550 70.880 65.570 ;
        RECT 51.950 65.520 53.910 65.550 ;
        RECT 70.430 65.520 70.890 65.550 ;
        RECT 51.950 65.170 70.890 65.520 ;
        RECT 51.950 59.070 53.910 65.170 ;
        RECT 70.430 65.150 70.890 65.170 ;
        RECT 70.450 65.140 70.880 65.150 ;
        RECT 71.130 64.730 71.330 67.640 ;
        RECT 74.850 67.520 75.170 67.640 ;
        RECT 72.100 66.230 74.870 66.240 ;
        RECT 72.100 66.040 75.170 66.230 ;
        RECT 71.350 64.740 71.780 64.760 ;
        RECT 71.340 64.730 71.790 64.740 ;
        RECT 55.880 64.350 71.790 64.730 ;
        RECT 51.920 58.430 53.950 59.070 ;
        RECT 55.880 59.050 57.840 64.350 ;
        RECT 69.980 64.190 70.240 64.350 ;
        RECT 70.010 63.910 70.210 64.190 ;
        RECT 71.130 63.910 71.330 64.350 ;
        RECT 71.350 64.330 71.780 64.350 ;
        RECT 72.100 63.920 72.310 66.040 ;
        RECT 74.850 65.910 75.170 66.040 ;
        RECT 73.880 64.580 74.190 64.610 ;
        RECT 74.840 64.580 75.160 64.620 ;
        RECT 73.880 64.330 75.160 64.580 ;
        RECT 72.100 63.910 72.720 63.920 ;
        RECT 60.030 63.530 72.720 63.910 ;
        RECT 60.030 59.070 62.010 63.530 ;
        RECT 70.010 63.120 70.210 63.530 ;
        RECT 71.130 63.120 71.330 63.530 ;
        RECT 72.100 63.120 72.310 63.530 ;
        RECT 73.110 63.120 73.530 63.150 ;
        RECT 64.140 62.740 73.530 63.120 ;
        RECT 51.910 58.420 53.950 58.430 ;
        RECT -144.230 44.190 -142.700 44.270 ;
        RECT -144.230 43.180 -142.190 44.190 ;
        RECT -147.240 42.540 -142.190 43.180 ;
        RECT -144.230 42.260 -142.190 42.540 ;
        RECT -144.230 41.640 -142.120 42.260 ;
        RECT -144.230 15.680 -142.830 41.640 ;
        RECT -144.230 15.600 -142.700 15.680 ;
        RECT -144.230 14.590 -142.190 15.600 ;
        RECT -147.240 13.950 -142.190 14.590 ;
        RECT -144.230 13.670 -142.190 13.950 ;
        RECT -144.230 13.050 -142.120 13.670 ;
        RECT -144.230 -12.910 -142.830 13.050 ;
        RECT -144.230 -12.990 -142.700 -12.910 ;
        RECT -144.230 -14.000 -142.190 -12.990 ;
        RECT -147.240 -14.640 -142.190 -14.000 ;
        RECT -144.230 -14.920 -142.190 -14.640 ;
        RECT -144.230 -15.540 -142.120 -14.920 ;
        RECT -144.230 -41.500 -142.830 -15.540 ;
        RECT -144.230 -41.580 -142.700 -41.500 ;
        RECT -144.230 -42.590 -142.190 -41.580 ;
        RECT -147.240 -43.230 -142.190 -42.590 ;
        RECT -144.230 -43.510 -142.190 -43.230 ;
        RECT -144.230 -44.130 -142.120 -43.510 ;
        RECT -144.230 -70.090 -142.830 -44.130 ;
        RECT -144.230 -70.170 -142.700 -70.090 ;
        RECT -144.230 -71.180 -142.190 -70.170 ;
        RECT -147.240 -71.820 -142.190 -71.180 ;
        RECT -144.230 -72.100 -142.190 -71.820 ;
        RECT -144.230 -72.720 -142.120 -72.100 ;
        RECT -144.230 -98.680 -142.830 -72.720 ;
        RECT -144.230 -98.760 -142.700 -98.680 ;
        RECT -144.230 -99.770 -142.190 -98.760 ;
        RECT -147.240 -100.410 -142.190 -99.770 ;
        RECT -144.230 -100.690 -142.190 -100.410 ;
        RECT -144.230 -101.310 -142.120 -100.690 ;
        RECT -144.230 -127.270 -142.830 -101.310 ;
        RECT -144.230 -127.350 -142.700 -127.270 ;
        RECT -144.230 -128.360 -142.190 -127.350 ;
        RECT -147.240 -129.000 -142.190 -128.360 ;
        RECT -144.230 -129.280 -142.190 -129.000 ;
        RECT -144.230 -129.900 -142.120 -129.280 ;
        RECT -144.230 -155.860 -142.830 -129.900 ;
        RECT -144.230 -155.940 -142.700 -155.860 ;
        RECT -144.230 -156.950 -142.190 -155.940 ;
        RECT -147.240 -157.590 -142.190 -156.950 ;
        RECT -144.230 -157.870 -142.190 -157.590 ;
        RECT -144.230 -158.490 -142.120 -157.870 ;
        RECT -144.230 -184.450 -142.830 -158.490 ;
        RECT -144.230 -184.530 -142.700 -184.450 ;
        RECT -144.230 -185.540 -142.190 -184.530 ;
        RECT -147.240 -186.180 -142.190 -185.540 ;
        RECT -144.230 -186.460 -142.190 -186.180 ;
        RECT -144.230 -187.080 -142.120 -186.460 ;
        RECT -144.230 -213.040 -142.830 -187.080 ;
        RECT -144.230 -213.120 -142.700 -213.040 ;
        RECT -144.230 -214.130 -142.190 -213.120 ;
        RECT -147.240 -214.770 -142.190 -214.130 ;
        RECT -144.230 -215.050 -142.190 -214.770 ;
        RECT -144.230 -215.670 -142.120 -215.050 ;
        RECT -144.230 -243.370 -142.830 -215.670 ;
        RECT 51.910 -238.160 53.930 58.420 ;
        RECT 55.870 58.400 57.900 59.050 ;
        RECT 59.990 58.420 62.020 59.070 ;
        RECT 64.140 59.040 66.120 62.740 ;
        RECT 70.010 59.950 70.210 62.740 ;
        RECT 71.130 59.950 71.330 62.740 ;
        RECT 72.100 59.950 72.310 62.740 ;
        RECT 73.110 62.710 73.530 62.740 ;
        RECT 73.880 59.950 74.180 64.330 ;
        RECT 74.840 64.300 75.160 64.330 ;
        RECT 74.840 62.980 75.160 63.000 ;
        RECT 74.840 62.680 75.190 62.980 ;
        RECT 75.000 61.390 75.190 62.680 ;
        RECT 74.840 61.070 75.190 61.390 ;
        RECT 75.000 59.950 75.190 61.070 ;
        RECT 69.210 59.750 75.450 59.950 ;
        RECT 69.210 59.070 69.410 59.750 ;
        RECT 70.010 59.070 70.210 59.750 ;
        RECT 55.880 -238.160 57.900 58.400 ;
        RECT 60.000 -238.160 62.020 58.420 ;
        RECT 64.130 58.390 66.160 59.040 ;
        RECT 68.120 58.420 70.210 59.070 ;
        RECT 64.130 -238.170 66.150 58.390 ;
        RECT 68.140 55.930 70.210 58.420 ;
        RECT 71.130 56.070 71.330 59.750 ;
        RECT 71.120 55.930 71.330 56.070 ;
        RECT 72.100 59.070 72.310 59.750 ;
        RECT 73.880 59.630 74.180 59.750 ;
        RECT 74.470 59.630 74.790 59.750 ;
        RECT 73.880 59.540 74.790 59.630 ;
        RECT 75.000 59.540 75.190 59.750 ;
        RECT 76.370 59.540 76.570 59.950 ;
        RECT 73.880 59.340 76.570 59.540 ;
        RECT 73.880 59.070 74.340 59.340 ;
        RECT 72.100 58.770 74.340 59.070 ;
        RECT 72.100 57.990 74.180 58.770 ;
        RECT 75.000 58.190 75.190 59.340 ;
        RECT 72.100 55.930 74.240 57.990 ;
        RECT 74.850 57.870 75.190 58.190 ;
        RECT 75.000 56.600 75.190 57.870 ;
        RECT 74.840 56.280 75.190 56.600 ;
        RECT 75.000 56.080 75.190 56.280 ;
        RECT 74.980 55.930 75.190 56.080 ;
        RECT 68.140 -238.160 70.160 55.930 ;
        RECT 72.150 -236.480 74.170 55.930 ;
        RECT 172.300 -51.510 174.390 79.920 ;
        RECT 176.540 -25.040 178.630 85.430 ;
        RECT 180.670 3.440 182.760 90.470 ;
        RECT 184.760 32.210 186.850 95.670 ;
        RECT 192.980 89.270 195.070 105.950 ;
        RECT 212.720 102.650 214.120 129.840 ;
        RECT 212.710 102.140 214.120 102.650 ;
        RECT 211.600 101.970 214.120 102.140 ;
        RECT 212.710 101.720 214.120 101.970 ;
        RECT 192.780 85.730 195.210 89.270 ;
        RECT 192.980 85.060 195.070 85.730 ;
        RECT 212.720 74.060 214.120 101.720 ;
        RECT 212.710 73.550 214.120 74.060 ;
        RECT 211.600 73.380 214.120 73.550 ;
        RECT 212.710 73.130 214.120 73.380 ;
        RECT 212.720 45.470 214.120 73.130 ;
        RECT 212.710 44.960 214.120 45.470 ;
        RECT 211.600 44.790 214.120 44.960 ;
        RECT 212.710 44.540 214.120 44.790 ;
        RECT 184.560 28.500 187.080 32.210 ;
        RECT 184.760 28.470 186.850 28.500 ;
        RECT 212.720 16.880 214.120 44.540 ;
        RECT 212.710 16.370 214.120 16.880 ;
        RECT 211.600 16.200 214.120 16.370 ;
        RECT 212.710 15.950 214.120 16.200 ;
        RECT 180.400 0.020 182.760 3.440 ;
        RECT 180.670 -0.690 182.760 0.020 ;
        RECT 212.720 -11.710 214.120 15.950 ;
        RECT 212.710 -12.220 214.120 -11.710 ;
        RECT 211.600 -12.390 214.120 -12.220 ;
        RECT 212.710 -12.640 214.120 -12.390 ;
        RECT 176.370 -28.750 178.800 -25.040 ;
        RECT 212.720 -40.300 214.120 -12.640 ;
        RECT 212.710 -40.810 214.120 -40.300 ;
        RECT 211.600 -40.980 214.120 -40.810 ;
        RECT 212.710 -41.230 214.120 -40.980 ;
        RECT 172.310 -53.410 174.390 -51.510 ;
        RECT 172.310 -53.530 174.400 -53.410 ;
        RECT 172.200 -53.590 174.400 -53.530 ;
        RECT 171.940 -57.270 174.470 -53.590 ;
        RECT 172.200 -57.290 174.290 -57.270 ;
        RECT 212.720 -68.890 214.120 -41.230 ;
        RECT 212.710 -69.400 214.120 -68.890 ;
        RECT 211.600 -69.570 214.120 -69.400 ;
        RECT 212.710 -69.820 214.120 -69.570 ;
        RECT 212.720 -69.980 214.120 -69.820 ;
        RECT 212.720 -70.380 214.130 -69.980 ;
        RECT 212.740 -71.070 214.120 -70.380 ;
        RECT 212.730 -72.240 214.130 -71.070 ;
        RECT 108.710 -79.140 113.310 -78.360 ;
        RECT 108.710 -80.820 207.860 -79.140 ;
        RECT 108.710 -82.110 207.990 -80.820 ;
        RECT 108.710 -82.930 113.310 -82.110 ;
        RECT 72.150 -238.140 74.190 -236.480 ;
      LAYER via2 ;
        RECT 49.580 113.550 49.900 113.870 ;
        RECT 50.610 113.540 50.930 113.860 ;
        RECT 49.620 106.580 49.950 106.930 ;
    END
  END VSSA1
  PIN VDDA1
    ANTENNADIFFAREA 125.345993 ;
    PORT
      LAYER nwell ;
        RECT 17.300 134.780 29.350 140.720 ;
        RECT 45.890 134.780 57.940 140.720 ;
        RECT 74.480 134.780 86.530 140.720 ;
        RECT 103.070 134.780 115.120 140.720 ;
        RECT 131.660 134.780 143.710 140.720 ;
        RECT 160.250 134.780 172.300 140.720 ;
        RECT 188.840 134.780 200.890 140.720 ;
        RECT 17.050 110.490 19.560 116.730 ;
        RECT 207.250 116.120 213.190 128.170 ;
        RECT 207.250 87.530 213.190 99.580 ;
        RECT 207.250 58.940 213.190 70.990 ;
        RECT 207.250 30.350 213.190 42.400 ;
        RECT 207.250 1.760 213.190 13.810 ;
        RECT 207.250 -26.830 213.190 -14.780 ;
        RECT 207.250 -55.420 213.190 -43.370 ;
      LAYER met2 ;
        RECT 28.770 135.920 29.410 138.360 ;
        RECT -25.550 135.350 29.920 135.920 ;
        RECT 57.360 135.350 58.000 138.360 ;
        RECT 85.950 135.350 86.590 138.360 ;
        RECT 114.540 135.350 115.180 138.360 ;
        RECT 143.130 135.350 143.770 138.360 ;
        RECT 171.720 135.350 172.360 138.360 ;
        RECT 200.310 135.350 200.950 138.360 ;
        RECT -25.550 134.520 207.830 135.350 ;
        RECT 2.430 133.950 207.830 134.520 ;
        RECT 27.870 133.820 30.500 133.950 ;
        RECT 56.460 133.820 59.090 133.950 ;
        RECT 85.050 133.820 87.680 133.950 ;
        RECT 113.640 133.820 116.270 133.950 ;
        RECT 142.230 133.820 144.860 133.950 ;
        RECT 170.820 133.820 173.450 133.950 ;
        RECT 199.410 133.820 202.040 133.950 ;
        RECT 27.870 133.310 30.420 133.820 ;
        RECT 56.460 133.310 59.010 133.820 ;
        RECT 85.050 133.310 87.600 133.820 ;
        RECT 113.640 133.310 116.190 133.820 ;
        RECT 142.230 133.310 144.780 133.820 ;
        RECT 170.820 133.310 173.370 133.820 ;
        RECT 199.410 133.310 201.960 133.820 ;
        RECT 27.870 133.240 28.490 133.310 ;
        RECT 56.460 133.240 57.080 133.310 ;
        RECT 85.050 133.240 85.670 133.310 ;
        RECT 113.640 133.240 114.260 133.310 ;
        RECT 142.230 133.240 142.850 133.310 ;
        RECT 170.820 133.240 171.440 133.310 ;
        RECT 199.410 133.240 200.030 133.310 ;
        RECT 206.420 129.320 207.820 133.950 ;
        RECT 206.290 129.240 207.820 129.320 ;
        RECT 205.780 128.230 207.820 129.240 ;
        RECT 205.780 127.590 210.830 128.230 ;
        RECT 205.780 127.310 207.820 127.590 ;
        RECT 205.710 126.690 207.820 127.310 ;
        RECT 18.940 123.860 19.440 123.890 ;
        RECT 24.660 123.860 25.160 123.890 ;
        RECT 18.940 123.450 49.100 123.860 ;
        RECT 19.090 123.420 49.100 123.450 ;
        RECT 26.210 112.380 26.500 112.560 ;
        RECT 24.500 110.340 24.810 110.350 ;
        RECT 26.210 110.340 26.390 112.380 ;
        RECT 22.330 110.160 33.860 110.340 ;
        RECT 24.500 110.020 24.810 110.160 ;
        RECT 24.350 109.320 24.660 109.390 ;
        RECT 22.330 109.310 24.660 109.320 ;
        RECT 26.210 109.310 26.390 110.160 ;
        RECT 31.630 109.310 31.950 109.360 ;
        RECT 34.040 109.310 34.360 109.330 ;
        RECT 22.330 109.170 34.360 109.310 ;
        RECT 22.330 109.120 36.060 109.170 ;
        RECT 22.330 109.100 33.860 109.120 ;
        RECT 23.640 109.090 33.860 109.100 ;
        RECT 24.350 109.060 24.660 109.090 ;
        RECT 25.380 108.940 26.390 109.090 ;
        RECT 31.630 109.040 31.950 109.090 ;
        RECT 34.040 109.070 36.060 109.120 ;
        RECT 34.080 109.000 36.060 109.070 ;
        RECT 35.540 108.990 36.060 109.000 ;
        RECT 206.420 100.730 207.820 126.690 ;
        RECT 206.290 100.650 207.820 100.730 ;
        RECT 205.780 99.640 207.820 100.650 ;
        RECT 205.780 99.000 210.830 99.640 ;
        RECT 205.780 98.720 207.820 99.000 ;
        RECT 205.710 98.100 207.820 98.720 ;
        RECT 206.420 72.140 207.820 98.100 ;
        RECT 206.290 72.060 207.820 72.140 ;
        RECT 205.780 71.050 207.820 72.060 ;
        RECT 205.780 70.410 210.830 71.050 ;
        RECT 205.780 70.130 207.820 70.410 ;
        RECT 205.710 69.510 207.820 70.130 ;
        RECT 206.420 43.550 207.820 69.510 ;
        RECT 206.290 43.470 207.820 43.550 ;
        RECT 205.780 42.460 207.820 43.470 ;
        RECT 205.780 41.820 210.830 42.460 ;
        RECT 205.780 41.540 207.820 41.820 ;
        RECT 205.710 40.920 207.820 41.540 ;
        RECT 206.420 14.960 207.820 40.920 ;
        RECT 206.290 14.880 207.820 14.960 ;
        RECT 205.780 13.870 207.820 14.880 ;
        RECT 205.780 13.230 210.830 13.870 ;
        RECT 205.780 12.950 207.820 13.230 ;
        RECT 205.710 12.330 207.820 12.950 ;
        RECT 206.420 -13.630 207.820 12.330 ;
        RECT 206.290 -13.710 207.820 -13.630 ;
        RECT 205.780 -14.720 207.820 -13.710 ;
        RECT 205.780 -15.360 210.830 -14.720 ;
        RECT 205.780 -15.640 207.820 -15.360 ;
        RECT 205.710 -16.260 207.820 -15.640 ;
        RECT 206.420 -42.220 207.820 -16.260 ;
        RECT 206.290 -42.300 207.820 -42.220 ;
        RECT 205.780 -43.310 207.820 -42.300 ;
        RECT 205.780 -43.950 210.830 -43.310 ;
        RECT 205.780 -44.230 207.820 -43.950 ;
        RECT 205.710 -44.850 207.820 -44.230 ;
        RECT 206.420 -70.230 207.820 -44.850 ;
        RECT 206.400 -70.290 207.820 -70.230 ;
        RECT 206.400 -71.010 207.800 -70.290 ;
        RECT 206.390 -71.130 207.800 -71.010 ;
        RECT 206.380 -71.280 207.800 -71.130 ;
        RECT 206.380 -72.180 207.790 -71.280 ;
    END
  END VDDA1
  PIN LADATAOUT01
    PORT
      LAYER met2 ;
        RECT 0.940 86.560 1.310 86.570 ;
        RECT 0.940 86.390 11.040 86.560 ;
        RECT 0.940 86.180 1.310 86.390 ;
        RECT 0.850 60.520 1.390 60.590 ;
        RECT -8.580 60.090 1.390 60.520 ;
        RECT -8.580 59.080 -6.600 60.090 ;
        RECT -8.630 58.420 -6.600 59.080 ;
        RECT -8.630 -236.590 -6.610 58.420 ;
        RECT -8.630 -238.150 -6.600 -236.590 ;
        RECT -8.630 -238.160 -6.610 -238.150 ;
    END
  END LADATAOUT01
  PIN LADATAOUT00
    PORT
      LAYER met2 ;
        RECT 0.250 85.020 0.640 85.120 ;
        RECT 0.250 84.850 11.040 85.020 ;
        RECT 0.250 84.750 0.640 84.850 ;
        RECT 0.200 61.360 0.740 61.400 ;
        RECT -12.630 61.320 0.740 61.360 ;
        RECT -12.680 60.930 0.740 61.320 ;
        RECT -12.680 59.050 -10.670 60.930 ;
        RECT 0.200 60.900 0.740 60.930 ;
        RECT -12.700 58.390 -10.670 59.050 ;
        RECT -12.690 -238.160 -10.670 58.390 ;
    END
  END LADATAOUT00
  PIN LADATAOUT02
    PORT
      LAYER met2 ;
        RECT 1.550 88.100 1.940 88.210 ;
        RECT 1.550 87.930 11.040 88.100 ;
        RECT 1.550 87.830 1.940 87.930 ;
        RECT 1.530 59.710 2.020 59.910 ;
        RECT -4.080 59.690 2.020 59.710 ;
        RECT -4.650 59.410 2.020 59.690 ;
        RECT -4.650 59.310 1.930 59.410 ;
        RECT -4.650 59.080 -2.670 59.310 ;
        RECT -4.670 58.420 -2.640 59.080 ;
        RECT -4.660 -236.600 -2.640 58.420 ;
        RECT -4.670 -238.160 -2.640 -236.600 ;
    END
  END LADATAOUT02
  PIN LADATAOUT03
    PORT
      LAYER met2 ;
        RECT 2.210 89.670 2.620 89.770 ;
        RECT 2.210 89.500 11.040 89.670 ;
        RECT 2.210 89.410 2.620 89.500 ;
        RECT 1.360 59.080 2.010 59.090 ;
        RECT -0.670 58.450 2.010 59.080 ;
        RECT -0.670 58.420 1.360 58.450 ;
        RECT -0.660 -236.600 1.360 58.420 ;
        RECT -0.670 -238.160 1.360 -236.600 ;
    END
  END LADATAOUT03
  PIN LADATAOUT04
    PORT
      LAYER met2 ;
        RECT 2.850 94.840 3.270 94.930 ;
        RECT 2.850 94.670 11.040 94.840 ;
        RECT 2.850 94.570 3.270 94.670 ;
        RECT 2.860 59.060 3.410 59.080 ;
        RECT 2.860 58.630 5.410 59.060 ;
        RECT 3.380 58.400 5.410 58.630 ;
        RECT 3.390 -238.160 5.410 58.400 ;
    END
  END LADATAOUT04
  PIN LADATAOUT05
    PORT
      LAYER met2 ;
        RECT 3.460 96.320 3.850 96.400 ;
        RECT 3.460 96.150 11.040 96.320 ;
        RECT 3.460 96.070 3.850 96.150 ;
        RECT 3.470 59.310 9.450 59.650 ;
        RECT 7.440 59.060 9.450 59.310 ;
        RECT 9.110 59.050 9.450 59.060 ;
        RECT 7.410 58.870 9.450 59.050 ;
        RECT 7.410 58.430 9.440 58.870 ;
        RECT 7.400 58.390 9.440 58.430 ;
        RECT 7.400 -236.590 9.420 58.390 ;
        RECT 7.390 -238.150 9.420 -236.590 ;
        RECT 7.400 -238.160 9.420 -238.150 ;
    END
  END LADATAOUT05
  PIN LADATAOUT06
    PORT
      LAYER met2 ;
        RECT 4.080 97.870 4.470 97.960 ;
        RECT 4.080 97.700 11.040 97.870 ;
        RECT 4.080 97.610 4.470 97.700 ;
        RECT 11.370 60.300 13.390 60.320 ;
        RECT 4.210 60.290 13.390 60.300 ;
        RECT 4.110 59.970 13.390 60.290 ;
        RECT 4.110 59.960 4.500 59.970 ;
        RECT 11.350 59.090 13.390 59.970 ;
        RECT 11.350 59.080 13.370 59.090 ;
        RECT 11.350 59.010 13.400 59.080 ;
        RECT 11.370 58.430 13.400 59.010 ;
        RECT 11.370 58.420 13.420 58.430 ;
        RECT 11.400 -238.160 13.420 58.420 ;
    END
  END LADATAOUT06
  PIN LADATAOUT07
    PORT
      LAYER met2 ;
        RECT 4.720 99.460 5.090 99.580 ;
        RECT 4.720 99.290 11.040 99.460 ;
        RECT 4.720 99.180 5.090 99.290 ;
        RECT 4.760 60.600 17.500 60.930 ;
        RECT 15.450 59.070 17.480 60.600 ;
        RECT 15.450 59.060 17.470 59.070 ;
        RECT 15.450 59.010 17.490 59.060 ;
        RECT 15.460 58.430 17.490 59.010 ;
        RECT 15.460 58.400 17.510 58.430 ;
        RECT 15.490 -238.160 17.510 58.400 ;
    END
  END LADATAOUT07
  PIN LADATAOUT08
    PORT
      LAYER met2 ;
        RECT 5.330 104.930 5.720 105.020 ;
        RECT 5.330 104.760 11.340 104.930 ;
        RECT 5.330 104.670 5.720 104.760 ;
        RECT 5.340 61.570 5.730 61.620 ;
        RECT 5.340 61.290 21.700 61.570 ;
        RECT 5.600 61.240 21.700 61.290 ;
        RECT 19.630 58.430 21.660 61.240 ;
        RECT 19.620 58.420 21.660 58.430 ;
        RECT 19.620 -236.600 21.640 58.420 ;
        RECT 19.610 -238.160 21.640 -236.600 ;
    END
  END LADATAOUT08
  PIN LADATAOUT09
    PORT
      LAYER met2 ;
        RECT 5.890 106.500 6.310 106.590 ;
        RECT 5.890 106.330 11.340 106.500 ;
        RECT 5.890 106.240 6.310 106.330 ;
        RECT 5.920 62.180 6.310 62.190 ;
        RECT 5.920 61.860 25.610 62.180 ;
        RECT 6.020 61.850 25.610 61.860 ;
        RECT 23.620 59.140 25.610 61.850 ;
        RECT 23.610 58.390 25.640 59.140 ;
        RECT 23.620 -236.600 25.640 58.390 ;
        RECT 23.610 -238.160 25.640 -236.600 ;
    END
  END LADATAOUT09
  PIN LADATAOUT10
    PORT
      LAYER met2 ;
        RECT 6.520 108.030 6.910 108.130 ;
        RECT 6.520 107.860 11.340 108.030 ;
        RECT 6.520 107.760 6.910 107.860 ;
        RECT 6.520 62.830 6.930 62.840 ;
        RECT 6.520 62.810 29.590 62.830 ;
        RECT 6.520 62.500 29.600 62.810 ;
        RECT 6.520 62.490 6.930 62.500 ;
        RECT 27.600 59.120 29.600 62.500 ;
        RECT 27.570 58.420 29.600 59.120 ;
        RECT 27.580 -236.600 29.600 58.420 ;
        RECT 27.570 -238.160 29.600 -236.600 ;
    END
  END LADATAOUT10
  PIN LADATAOUT11
    PORT
      LAYER met2 ;
        RECT 7.130 109.600 7.520 109.710 ;
        RECT 7.130 109.430 11.340 109.600 ;
        RECT 7.130 109.330 7.520 109.430 ;
        RECT 7.100 63.450 7.510 63.460 ;
        RECT 7.090 63.120 33.610 63.450 ;
        RECT 7.100 63.100 7.510 63.120 ;
        RECT 31.700 59.050 33.610 63.120 ;
        RECT 31.620 58.400 33.650 59.050 ;
        RECT 31.630 -236.590 33.650 58.400 ;
        RECT 31.630 -238.150 33.660 -236.590 ;
        RECT 31.630 -238.160 33.650 -238.150 ;
    END
  END LADATAOUT11
  PIN LADATAOUT12
    PORT
      LAYER met2 ;
        RECT 7.770 110.170 8.160 110.260 ;
        RECT 7.770 110.000 11.340 110.170 ;
        RECT 7.770 109.910 8.160 110.000 ;
        RECT 7.760 64.120 8.160 64.140 ;
        RECT 7.760 63.790 37.700 64.120 ;
        RECT 7.760 63.780 8.160 63.790 ;
        RECT 35.740 59.070 37.690 63.790 ;
        RECT 35.690 58.430 37.720 59.070 ;
        RECT 35.690 58.420 37.740 58.430 ;
        RECT 35.720 -238.160 37.740 58.420 ;
    END
  END LADATAOUT12
  PIN LADATAOUT13
    PORT
      LAYER met2 ;
        RECT 8.410 111.770 8.800 111.870 ;
        RECT 8.410 111.600 11.340 111.770 ;
        RECT 8.410 111.500 8.800 111.600 ;
        RECT 8.350 64.760 8.770 64.770 ;
        RECT 8.350 64.430 41.710 64.760 ;
        RECT 8.350 64.420 8.770 64.430 ;
        RECT 39.720 59.070 41.710 64.430 ;
        RECT 39.720 58.420 41.750 59.070 ;
        RECT 39.730 -236.610 41.750 58.420 ;
        RECT 39.730 -238.160 41.760 -236.610 ;
        RECT 39.740 -238.170 41.760 -238.160 ;
    END
  END LADATAOUT13
  PIN LADATAOUT14
    PORT
      LAYER met2 ;
        RECT 9.010 113.350 9.340 113.360 ;
        RECT 8.990 113.250 9.360 113.350 ;
        RECT 8.990 113.080 11.340 113.250 ;
        RECT 8.990 112.970 9.360 113.080 ;
        RECT 8.990 65.390 9.370 65.400 ;
        RECT 8.990 65.060 45.790 65.390 ;
        RECT 8.990 65.050 9.370 65.060 ;
        RECT 39.720 65.050 45.790 65.060 ;
        RECT 43.830 64.730 45.790 65.050 ;
        RECT 43.830 59.070 45.780 64.730 ;
        RECT 43.770 58.420 45.800 59.070 ;
        RECT 43.770 -236.600 45.790 58.420 ;
        RECT 43.770 -238.160 45.800 -236.600 ;
    END
  END LADATAOUT14
  PIN LADATAOUT15
    PORT
      LAYER met2 ;
        RECT 9.610 114.890 10.000 114.980 ;
        RECT 9.610 114.720 11.340 114.890 ;
        RECT 9.590 66.010 10.010 66.020 ;
        RECT 9.590 65.760 49.860 66.010 ;
        RECT 9.590 65.680 49.870 65.760 ;
        RECT 9.590 65.670 10.010 65.680 ;
        RECT 43.830 65.660 49.870 65.680 ;
        RECT 47.930 65.160 49.870 65.660 ;
        RECT 47.930 59.090 49.860 65.160 ;
        RECT 47.840 58.430 49.870 59.090 ;
        RECT 47.840 58.310 49.880 58.430 ;
        RECT 47.860 -236.620 49.880 58.310 ;
        RECT 47.860 -238.160 49.890 -236.620 ;
        RECT 47.870 -238.180 49.890 -238.160 ;
    END
  END LADATAOUT15
  PIN LADATAOUT22
    PORT
      LAYER met2 ;
        RECT 77.340 59.070 77.550 59.960 ;
        RECT 76.220 58.430 78.250 59.070 ;
        RECT 76.220 58.420 78.260 58.430 ;
        RECT 76.240 -236.500 78.260 58.420 ;
        RECT 76.240 -238.160 78.270 -236.500 ;
    END
  END LADATAOUT22
  PIN LADATAOUT23
    PORT
      LAYER met2 ;
        RECT 79.270 58.980 79.480 59.960 ;
        RECT 80.400 58.980 82.430 59.070 ;
        RECT 79.270 58.770 82.430 58.980 ;
        RECT 80.400 58.420 82.430 58.770 ;
        RECT 80.410 -238.160 82.430 58.420 ;
    END
  END LADATAOUT23
  PIN LADATAOUT24
    PORT
      LAYER met2 ;
        RECT 80.240 59.770 80.430 59.940 ;
        RECT 80.240 59.580 85.240 59.770 ;
        RECT 85.050 59.050 85.240 59.580 ;
        RECT 85.890 59.050 86.080 59.120 ;
        RECT 84.380 58.430 86.410 59.050 ;
        RECT 84.380 58.400 86.430 58.430 ;
        RECT 84.410 -236.500 86.430 58.400 ;
        RECT 84.410 -238.160 86.440 -236.500 ;
    END
  END LADATAOUT24
  PIN LADATAIN00
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 38.730 84.990 39.040 85.100 ;
        RECT 44.520 84.990 44.840 85.040 ;
        RECT 38.730 84.980 44.840 84.990 ;
        RECT 37.800 84.830 44.840 84.980 ;
        RECT 37.800 84.800 39.040 84.830 ;
        RECT 38.730 84.770 39.040 84.800 ;
        RECT 44.520 84.780 44.840 84.830 ;
        RECT 44.500 76.860 90.290 76.870 ;
        RECT 44.500 76.370 90.500 76.860 ;
        RECT 88.490 59.070 90.500 76.370 ;
        RECT 88.430 58.550 90.500 59.070 ;
        RECT 88.430 58.430 90.460 58.550 ;
        RECT 88.420 58.420 90.460 58.430 ;
        RECT 88.420 -236.500 90.440 58.420 ;
        RECT 88.390 -238.160 90.440 -236.500 ;
    END
  END LADATAIN00
  PIN LADATAIN01
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 38.730 85.950 39.040 85.980 ;
        RECT 37.790 85.920 39.040 85.950 ;
        RECT 45.020 85.920 45.340 85.970 ;
        RECT 37.790 85.790 45.340 85.920 ;
        RECT 38.730 85.760 45.340 85.790 ;
        RECT 38.730 85.650 39.040 85.760 ;
        RECT 45.020 85.710 45.340 85.760 ;
        RECT 44.980 77.750 94.250 77.770 ;
        RECT 44.980 77.270 94.360 77.750 ;
        RECT 92.350 59.070 94.360 77.270 ;
        RECT 92.350 58.420 94.420 59.070 ;
        RECT 92.350 58.380 94.400 58.420 ;
        RECT 92.380 -236.500 94.400 58.380 ;
        RECT 92.370 -238.160 94.400 -236.500 ;
    END
  END LADATAIN01
  PIN LADATAIN02
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 37.800 87.870 39.010 87.980 ;
        RECT 37.800 87.780 39.040 87.870 ;
        RECT 38.730 87.760 39.040 87.780 ;
        RECT 45.490 87.760 45.810 87.810 ;
        RECT 38.730 87.600 45.810 87.760 ;
        RECT 38.730 87.540 39.040 87.600 ;
        RECT 45.490 87.550 45.810 87.600 ;
        RECT 96.430 78.670 98.440 78.690 ;
        RECT 45.450 78.170 98.440 78.670 ;
        RECT 96.430 59.050 98.440 78.170 ;
        RECT 96.430 58.400 98.470 59.050 ;
        RECT 96.430 -236.500 98.450 58.400 ;
        RECT 96.430 -238.160 98.470 -236.500 ;
    END
  END LADATAIN02
  PIN LADATAIN03
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 37.810 88.840 37.850 88.930 ;
        RECT 37.700 88.750 38.910 88.840 ;
        RECT 37.700 88.690 39.040 88.750 ;
        RECT 46.010 88.690 46.330 88.740 ;
        RECT 37.700 88.640 46.330 88.690 ;
        RECT 38.730 88.530 46.330 88.640 ;
        RECT 38.730 88.420 39.040 88.530 ;
        RECT 46.010 88.480 46.330 88.530 ;
        RECT 45.990 79.530 101.820 79.570 ;
        RECT 45.990 79.070 102.530 79.530 ;
        RECT 100.520 59.070 102.530 79.070 ;
        RECT 100.490 58.490 102.530 59.070 ;
        RECT 100.490 58.420 102.520 58.490 ;
        RECT 100.490 -236.500 102.510 58.420 ;
        RECT 100.490 -238.160 102.530 -236.500 ;
    END
  END LADATAIN03
  OBS
      LAYER nwell ;
        RECT -18.200 123.320 -8.510 127.920 ;
        RECT 3.820 126.200 6.040 127.890 ;
        RECT -18.800 121.930 -8.510 123.320 ;
        RECT 57.500 113.080 60.220 114.730 ;
        RECT 71.820 114.720 73.550 115.470 ;
        RECT 57.500 113.040 60.210 113.080 ;
        RECT 57.500 111.710 60.210 111.750 ;
        RECT 57.500 111.650 60.220 111.710 ;
        RECT 56.410 111.640 60.220 111.650 ;
        RECT 56.610 111.330 56.930 111.630 ;
        RECT 11.970 109.880 12.210 109.930 ;
        RECT 11.730 109.870 13.200 109.880 ;
        RECT 11.430 109.790 13.200 109.870 ;
        RECT 17.460 109.790 19.670 109.880 ;
        RECT 22.330 109.640 25.640 110.830 ;
        RECT 22.330 109.630 26.290 109.640 ;
        RECT 11.320 102.930 13.090 109.170 ;
        RECT 17.050 102.930 19.560 109.170 ;
        RECT 22.330 107.020 26.300 109.630 ;
        RECT 27.370 108.450 30.090 110.100 ;
        RECT 27.380 108.410 30.090 108.450 ;
        RECT 41.700 110.090 43.430 110.840 ;
        RECT 27.380 107.080 30.090 107.120 ;
        RECT 27.370 107.020 30.090 107.080 ;
        RECT 22.330 107.010 30.090 107.020 ;
        RECT 22.330 106.520 26.300 107.010 ;
        RECT 22.330 106.340 26.370 106.520 ;
        RECT 22.330 104.800 26.300 106.340 ;
        RECT 27.370 105.430 30.090 107.010 ;
        RECT 41.700 106.520 43.440 110.090 ;
        RECT 45.460 108.450 48.180 110.100 ;
        RECT 57.500 110.060 60.220 111.640 ;
        RECT 71.820 111.150 73.560 114.720 ;
        RECT 78.880 111.330 79.200 111.630 ;
        RECT 71.820 109.430 73.550 111.150 ;
        RECT 45.460 108.410 48.170 108.450 ;
        RECT 45.460 107.080 48.170 107.120 ;
        RECT 41.700 104.800 43.430 106.520 ;
        RECT 45.460 105.430 48.180 107.080 ;
        RECT 25.600 103.580 26.300 104.800 ;
        RECT 37.790 103.520 40.340 103.530 ;
        RECT 26.300 101.470 26.380 101.650 ;
        RECT 11.320 92.800 13.090 99.040 ;
        RECT 17.050 92.800 19.560 99.040 ;
        RECT 37.780 97.500 40.340 103.520 ;
        RECT 37.790 97.490 40.340 97.500 ;
        RECT 41.870 97.480 44.100 103.530 ;
        RECT 46.120 101.670 47.850 103.530 ;
        RECT 46.120 99.830 47.860 101.670 ;
        RECT 46.120 97.480 47.850 99.830 ;
        RECT 56.860 97.480 59.090 103.530 ;
        RECT 37.060 89.750 37.460 89.890 ;
        RECT -13.840 84.610 -11.470 87.480 ;
        RECT 27.500 78.430 29.520 82.390 ;
        RECT 27.400 78.400 30.790 78.430 ;
        RECT -14.420 71.170 -13.800 76.870 ;
        RECT -13.430 73.950 -13.420 73.990 ;
        RECT -12.420 70.950 -9.030 76.650 ;
        RECT 17.590 72.700 20.980 78.400 ;
        RECT 21.980 75.360 21.990 75.400 ;
        RECT 22.360 72.480 22.980 78.180 ;
        RECT 24.260 72.480 24.880 78.180 ;
        RECT 25.250 75.360 25.260 75.400 ;
        RECT 26.260 72.730 30.790 78.400 ;
        RECT 31.790 75.390 31.800 75.430 ;
        RECT 26.260 72.700 29.650 72.730 ;
        RECT 32.170 72.510 32.790 78.210 ;
        RECT 34.070 72.510 34.690 78.210 ;
        RECT 35.060 75.390 35.070 75.430 ;
        RECT 36.070 72.730 39.460 78.430 ;
        RECT 69.250 56.300 74.900 72.400 ;
      LAYER li1 ;
        RECT -131.040 141.800 -130.790 143.260 ;
        RECT -131.000 141.790 -130.830 141.800 ;
        RECT -124.360 141.770 -124.110 143.240 ;
        RECT -102.450 141.800 -102.200 143.260 ;
        RECT -102.410 141.790 -102.240 141.800 ;
        RECT -95.770 141.770 -95.520 143.240 ;
        RECT -73.860 141.800 -73.610 143.260 ;
        RECT -73.820 141.790 -73.650 141.800 ;
        RECT -67.180 141.770 -66.930 143.240 ;
        RECT -4.410 142.560 -4.190 143.680 ;
        RECT -4.460 142.370 -4.130 142.560 ;
        RECT 2.330 142.370 2.570 143.720 ;
        RECT 10.160 142.170 10.410 143.260 ;
        RECT 16.840 142.170 17.090 143.240 ;
        RECT -25.170 141.900 29.570 142.170 ;
        RECT -25.170 141.770 -0.830 141.900 ;
        RECT 7.860 141.770 29.570 141.900 ;
        RECT 38.750 141.800 39.000 143.260 ;
        RECT 38.790 141.790 38.960 141.800 ;
        RECT 45.430 141.770 45.680 143.240 ;
        RECT 67.340 141.800 67.590 143.260 ;
        RECT 67.380 141.790 67.550 141.800 ;
        RECT 74.020 141.770 74.270 143.240 ;
        RECT 95.930 141.800 96.180 143.260 ;
        RECT 95.970 141.790 96.140 141.800 ;
        RECT 102.610 141.770 102.860 143.240 ;
        RECT 124.520 141.800 124.770 143.260 ;
        RECT 124.560 141.790 124.730 141.800 ;
        RECT 131.200 141.770 131.450 143.240 ;
        RECT 153.110 141.800 153.360 143.260 ;
        RECT 153.150 141.790 153.320 141.800 ;
        RECT 159.790 141.770 160.040 143.240 ;
        RECT 181.700 141.800 181.950 143.260 ;
        RECT 181.740 141.790 181.910 141.800 ;
        RECT 188.380 141.770 188.630 143.240 ;
        RECT -138.220 141.050 -110.840 141.560 ;
        RECT -138.220 139.120 -137.420 141.050 ;
        RECT -136.840 140.600 -136.670 140.680 ;
        RECT -125.600 140.600 -125.370 140.690 ;
        RECT -136.840 140.590 -125.370 140.600 ;
        RECT -138.220 134.540 -137.710 139.120 ;
        RECT -136.850 135.120 -125.370 140.590 ;
        RECT -136.920 134.950 -125.370 135.120 ;
        RECT -136.850 134.890 -136.660 134.950 ;
        RECT -125.600 134.710 -125.370 134.950 ;
        RECT -136.970 134.540 -135.170 134.550 ;
        RECT -124.810 134.540 -124.300 141.050 ;
        RECT -123.540 140.160 -112.290 140.330 ;
        RECT -123.540 135.290 -123.370 140.160 ;
        RECT -122.980 139.830 -112.870 139.850 ;
        RECT -122.980 139.790 -112.850 139.830 ;
        RECT -123.030 139.620 -112.850 139.790 ;
        RECT -122.980 135.600 -112.850 139.620 ;
        RECT -112.460 138.400 -112.290 140.160 ;
        RECT -122.980 135.520 -112.870 135.600 ;
        RECT -123.550 135.220 -123.370 135.290 ;
        RECT -112.460 135.220 -111.850 138.400 ;
        RECT -123.550 135.050 -111.850 135.220 ;
        RECT -112.390 134.940 -111.850 135.050 ;
        RECT -111.390 134.700 -110.840 141.050 ;
        RECT -111.400 134.540 -110.840 134.700 ;
        RECT -138.220 134.200 -110.840 134.540 ;
        RECT -109.630 141.050 -82.250 141.560 ;
        RECT -109.630 139.120 -108.830 141.050 ;
        RECT -108.250 140.600 -108.080 140.680 ;
        RECT -97.010 140.600 -96.780 140.690 ;
        RECT -108.250 140.590 -96.780 140.600 ;
        RECT -109.630 134.540 -109.120 139.120 ;
        RECT -108.260 135.120 -96.780 140.590 ;
        RECT -108.330 134.950 -96.780 135.120 ;
        RECT -108.260 134.890 -108.070 134.950 ;
        RECT -97.010 134.710 -96.780 134.950 ;
        RECT -108.380 134.540 -106.580 134.550 ;
        RECT -96.220 134.540 -95.710 141.050 ;
        RECT -94.950 140.160 -83.700 140.330 ;
        RECT -94.950 135.290 -94.780 140.160 ;
        RECT -94.390 139.830 -84.280 139.850 ;
        RECT -94.390 139.790 -84.260 139.830 ;
        RECT -94.440 139.620 -84.260 139.790 ;
        RECT -94.390 135.600 -84.260 139.620 ;
        RECT -83.870 138.400 -83.700 140.160 ;
        RECT -94.390 135.520 -84.280 135.600 ;
        RECT -94.960 135.220 -94.780 135.290 ;
        RECT -83.870 135.220 -83.260 138.400 ;
        RECT -94.960 135.050 -83.260 135.220 ;
        RECT -83.800 134.940 -83.260 135.050 ;
        RECT -82.800 134.700 -82.250 141.050 ;
        RECT -82.810 134.540 -82.250 134.700 ;
        RECT -109.630 134.200 -82.250 134.540 ;
        RECT -81.040 141.050 -53.660 141.560 ;
        RECT -81.040 139.120 -80.240 141.050 ;
        RECT -79.660 140.600 -79.490 140.680 ;
        RECT -68.420 140.600 -68.190 140.690 ;
        RECT -79.660 140.590 -68.190 140.600 ;
        RECT -81.040 134.540 -80.530 139.120 ;
        RECT -79.670 135.120 -68.190 140.590 ;
        RECT -79.740 134.950 -68.190 135.120 ;
        RECT -79.670 134.890 -79.480 134.950 ;
        RECT -68.420 134.710 -68.190 134.950 ;
        RECT -79.790 134.540 -77.990 134.550 ;
        RECT -67.630 134.540 -67.120 141.050 ;
        RECT -66.360 140.160 -55.110 140.330 ;
        RECT -66.360 135.290 -66.190 140.160 ;
        RECT -65.800 139.830 -55.690 139.850 ;
        RECT -65.800 139.790 -55.670 139.830 ;
        RECT -65.850 139.620 -55.670 139.790 ;
        RECT -65.800 135.600 -55.670 139.620 ;
        RECT -55.280 138.400 -55.110 140.160 ;
        RECT -65.800 135.520 -55.690 135.600 ;
        RECT -66.370 135.220 -66.190 135.290 ;
        RECT -55.280 135.220 -54.670 138.400 ;
        RECT -66.370 135.050 -54.670 135.220 ;
        RECT -55.210 134.940 -54.670 135.050 ;
        RECT -54.210 134.700 -53.660 141.050 ;
        RECT -54.220 134.540 -53.660 134.700 ;
        RECT -81.040 134.200 -53.660 134.540 ;
        RECT -138.190 134.030 -110.840 134.200 ;
        RECT -109.600 134.030 -82.250 134.200 ;
        RECT -81.010 134.030 -53.660 134.200 ;
        RECT -25.170 134.170 -25.000 141.770 ;
        RECT 29.400 141.560 29.570 141.770 ;
        RECT 2.980 141.050 30.360 141.560 ;
        RECT 2.980 139.120 3.780 141.050 ;
        RECT 4.360 140.600 4.530 140.680 ;
        RECT 15.600 140.600 15.830 140.690 ;
        RECT 4.360 140.590 15.830 140.600 ;
        RECT 2.980 134.540 3.490 139.120 ;
        RECT 4.350 135.120 15.830 140.590 ;
        RECT 4.280 134.950 15.830 135.120 ;
        RECT 4.350 134.890 4.540 134.950 ;
        RECT 15.600 134.710 15.830 134.950 ;
        RECT 4.230 134.540 6.030 134.550 ;
        RECT 16.390 134.540 16.900 141.050 ;
        RECT 17.660 140.160 28.910 140.330 ;
        RECT 17.660 135.290 17.830 140.160 ;
        RECT 18.220 139.830 28.330 139.850 ;
        RECT 18.220 139.790 28.350 139.830 ;
        RECT 18.170 139.620 28.350 139.790 ;
        RECT 18.220 135.600 28.350 139.620 ;
        RECT 28.740 138.400 28.910 140.160 ;
        RECT 18.220 135.520 28.330 135.600 ;
        RECT 17.650 135.220 17.830 135.290 ;
        RECT 28.740 135.220 29.350 138.400 ;
        RECT 17.650 135.050 29.350 135.220 ;
        RECT 28.810 134.940 29.350 135.050 ;
        RECT 29.400 134.690 29.570 141.050 ;
        RECT 29.810 134.700 30.360 141.050 ;
        RECT 29.800 134.540 30.360 134.700 ;
        RECT 2.980 134.200 30.360 134.540 ;
        RECT 31.570 141.050 58.950 141.560 ;
        RECT 31.570 139.120 32.370 141.050 ;
        RECT 32.950 140.600 33.120 140.680 ;
        RECT 44.190 140.600 44.420 140.690 ;
        RECT 32.950 140.590 44.420 140.600 ;
        RECT 31.570 134.540 32.080 139.120 ;
        RECT 32.940 135.120 44.420 140.590 ;
        RECT 32.870 134.950 44.420 135.120 ;
        RECT 32.940 134.890 33.130 134.950 ;
        RECT 44.190 134.710 44.420 134.950 ;
        RECT 32.820 134.540 34.620 134.550 ;
        RECT 44.980 134.540 45.490 141.050 ;
        RECT 46.250 140.160 57.500 140.330 ;
        RECT 46.250 135.290 46.420 140.160 ;
        RECT 46.810 139.830 56.920 139.850 ;
        RECT 46.810 139.790 56.940 139.830 ;
        RECT 46.760 139.620 56.940 139.790 ;
        RECT 46.810 135.600 56.940 139.620 ;
        RECT 57.330 138.400 57.500 140.160 ;
        RECT 46.810 135.520 56.920 135.600 ;
        RECT 46.240 135.220 46.420 135.290 ;
        RECT 57.330 135.220 57.940 138.400 ;
        RECT 46.240 135.050 57.940 135.220 ;
        RECT 57.400 134.940 57.940 135.050 ;
        RECT 58.400 134.700 58.950 141.050 ;
        RECT 58.390 134.540 58.950 134.700 ;
        RECT 31.570 134.200 58.950 134.540 ;
        RECT 60.160 141.050 87.540 141.560 ;
        RECT 60.160 139.120 60.960 141.050 ;
        RECT 61.540 140.600 61.710 140.680 ;
        RECT 72.780 140.600 73.010 140.690 ;
        RECT 61.540 140.590 73.010 140.600 ;
        RECT 60.160 134.540 60.670 139.120 ;
        RECT 61.530 135.120 73.010 140.590 ;
        RECT 61.460 134.950 73.010 135.120 ;
        RECT 61.530 134.890 61.720 134.950 ;
        RECT 72.780 134.710 73.010 134.950 ;
        RECT 61.410 134.540 63.210 134.550 ;
        RECT 73.570 134.540 74.080 141.050 ;
        RECT 74.840 140.160 86.090 140.330 ;
        RECT 74.840 135.290 75.010 140.160 ;
        RECT 75.400 139.830 85.510 139.850 ;
        RECT 75.400 139.790 85.530 139.830 ;
        RECT 75.350 139.620 85.530 139.790 ;
        RECT 75.400 135.600 85.530 139.620 ;
        RECT 85.920 138.400 86.090 140.160 ;
        RECT 75.400 135.520 85.510 135.600 ;
        RECT 74.830 135.220 75.010 135.290 ;
        RECT 85.920 135.220 86.530 138.400 ;
        RECT 74.830 135.050 86.530 135.220 ;
        RECT 85.990 134.940 86.530 135.050 ;
        RECT 86.990 134.700 87.540 141.050 ;
        RECT 86.980 134.540 87.540 134.700 ;
        RECT 60.160 134.200 87.540 134.540 ;
        RECT 88.750 141.050 116.130 141.560 ;
        RECT 88.750 139.120 89.550 141.050 ;
        RECT 90.130 140.600 90.300 140.680 ;
        RECT 101.370 140.600 101.600 140.690 ;
        RECT 90.130 140.590 101.600 140.600 ;
        RECT 88.750 134.540 89.260 139.120 ;
        RECT 90.120 135.120 101.600 140.590 ;
        RECT 90.050 134.950 101.600 135.120 ;
        RECT 90.120 134.890 90.310 134.950 ;
        RECT 101.370 134.710 101.600 134.950 ;
        RECT 90.000 134.540 91.800 134.550 ;
        RECT 102.160 134.540 102.670 141.050 ;
        RECT 103.430 140.160 114.680 140.330 ;
        RECT 103.430 135.290 103.600 140.160 ;
        RECT 103.990 139.830 114.100 139.850 ;
        RECT 103.990 139.790 114.120 139.830 ;
        RECT 103.940 139.620 114.120 139.790 ;
        RECT 103.990 135.600 114.120 139.620 ;
        RECT 114.510 138.400 114.680 140.160 ;
        RECT 103.990 135.520 114.100 135.600 ;
        RECT 103.420 135.220 103.600 135.290 ;
        RECT 114.510 135.220 115.120 138.400 ;
        RECT 103.420 135.050 115.120 135.220 ;
        RECT 114.580 134.940 115.120 135.050 ;
        RECT 115.580 134.700 116.130 141.050 ;
        RECT 115.570 134.540 116.130 134.700 ;
        RECT 88.750 134.200 116.130 134.540 ;
        RECT 117.340 141.050 144.720 141.560 ;
        RECT 117.340 139.120 118.140 141.050 ;
        RECT 118.720 140.600 118.890 140.680 ;
        RECT 129.960 140.600 130.190 140.690 ;
        RECT 118.720 140.590 130.190 140.600 ;
        RECT 117.340 134.540 117.850 139.120 ;
        RECT 118.710 135.120 130.190 140.590 ;
        RECT 118.640 134.950 130.190 135.120 ;
        RECT 118.710 134.890 118.900 134.950 ;
        RECT 129.960 134.710 130.190 134.950 ;
        RECT 118.590 134.540 120.390 134.550 ;
        RECT 130.750 134.540 131.260 141.050 ;
        RECT 132.020 140.160 143.270 140.330 ;
        RECT 132.020 135.290 132.190 140.160 ;
        RECT 132.580 139.830 142.690 139.850 ;
        RECT 132.580 139.790 142.710 139.830 ;
        RECT 132.530 139.620 142.710 139.790 ;
        RECT 132.580 135.600 142.710 139.620 ;
        RECT 143.100 138.400 143.270 140.160 ;
        RECT 132.580 135.520 142.690 135.600 ;
        RECT 132.010 135.220 132.190 135.290 ;
        RECT 143.100 135.220 143.710 138.400 ;
        RECT 132.010 135.050 143.710 135.220 ;
        RECT 143.170 134.940 143.710 135.050 ;
        RECT 144.170 134.700 144.720 141.050 ;
        RECT 144.160 134.540 144.720 134.700 ;
        RECT 117.340 134.200 144.720 134.540 ;
        RECT 145.930 141.050 173.310 141.560 ;
        RECT 145.930 139.120 146.730 141.050 ;
        RECT 147.310 140.600 147.480 140.680 ;
        RECT 158.550 140.600 158.780 140.690 ;
        RECT 147.310 140.590 158.780 140.600 ;
        RECT 145.930 134.540 146.440 139.120 ;
        RECT 147.300 135.120 158.780 140.590 ;
        RECT 147.230 134.950 158.780 135.120 ;
        RECT 147.300 134.890 147.490 134.950 ;
        RECT 158.550 134.710 158.780 134.950 ;
        RECT 147.180 134.540 148.980 134.550 ;
        RECT 159.340 134.540 159.850 141.050 ;
        RECT 160.610 140.160 171.860 140.330 ;
        RECT 160.610 135.290 160.780 140.160 ;
        RECT 161.170 139.830 171.280 139.850 ;
        RECT 161.170 139.790 171.300 139.830 ;
        RECT 161.120 139.620 171.300 139.790 ;
        RECT 161.170 135.600 171.300 139.620 ;
        RECT 171.690 138.400 171.860 140.160 ;
        RECT 161.170 135.520 171.280 135.600 ;
        RECT 160.600 135.220 160.780 135.290 ;
        RECT 171.690 135.220 172.300 138.400 ;
        RECT 160.600 135.050 172.300 135.220 ;
        RECT 171.760 134.940 172.300 135.050 ;
        RECT 172.760 134.700 173.310 141.050 ;
        RECT 172.750 134.540 173.310 134.700 ;
        RECT 145.930 134.200 173.310 134.540 ;
        RECT 174.520 141.050 201.900 141.560 ;
        RECT 174.520 139.120 175.320 141.050 ;
        RECT 175.900 140.600 176.070 140.680 ;
        RECT 187.140 140.600 187.370 140.690 ;
        RECT 175.900 140.590 187.370 140.600 ;
        RECT 174.520 134.540 175.030 139.120 ;
        RECT 175.890 135.120 187.370 140.590 ;
        RECT 175.820 134.950 187.370 135.120 ;
        RECT 175.890 134.890 176.080 134.950 ;
        RECT 187.140 134.710 187.370 134.950 ;
        RECT 175.770 134.540 177.570 134.550 ;
        RECT 187.930 134.540 188.440 141.050 ;
        RECT 189.200 140.160 200.450 140.330 ;
        RECT 189.200 135.290 189.370 140.160 ;
        RECT 189.760 139.830 199.870 139.850 ;
        RECT 189.760 139.790 199.890 139.830 ;
        RECT 189.710 139.620 199.890 139.790 ;
        RECT 189.760 135.600 199.890 139.620 ;
        RECT 200.280 138.400 200.450 140.160 ;
        RECT 189.760 135.520 199.870 135.600 ;
        RECT 189.190 135.220 189.370 135.290 ;
        RECT 200.280 135.220 200.890 138.400 ;
        RECT 189.190 135.050 200.890 135.220 ;
        RECT 200.350 134.940 200.890 135.050 ;
        RECT 201.350 134.700 201.900 141.050 ;
        RECT 201.340 134.540 201.900 134.700 ;
        RECT 174.520 134.200 201.900 134.540 ;
        RECT 3.010 134.030 30.360 134.200 ;
        RECT 31.600 134.030 58.950 134.200 ;
        RECT 60.190 134.030 87.540 134.200 ;
        RECT 88.780 134.030 116.130 134.200 ;
        RECT 117.370 134.030 144.720 134.200 ;
        RECT 145.960 134.030 173.310 134.200 ;
        RECT 174.550 134.030 201.900 134.200 ;
        RECT -138.190 134.010 -137.500 134.030 ;
        RECT -136.990 134.020 -135.190 134.030 ;
        RECT -109.600 134.010 -108.910 134.030 ;
        RECT -108.400 134.020 -106.600 134.030 ;
        RECT -81.010 134.010 -80.320 134.030 ;
        RECT -79.810 134.020 -78.010 134.030 ;
        RECT 3.010 134.010 3.700 134.030 ;
        RECT 4.210 134.020 6.010 134.030 ;
        RECT 31.600 134.010 32.290 134.030 ;
        RECT 32.800 134.020 34.600 134.030 ;
        RECT 60.190 134.010 60.880 134.030 ;
        RECT 61.390 134.020 63.190 134.030 ;
        RECT 88.780 134.010 89.470 134.030 ;
        RECT 89.980 134.020 91.780 134.030 ;
        RECT 117.370 134.010 118.060 134.030 ;
        RECT 118.570 134.020 120.370 134.030 ;
        RECT 145.960 134.010 146.650 134.030 ;
        RECT 147.160 134.020 148.960 134.030 ;
        RECT 174.550 134.010 175.240 134.030 ;
        RECT 175.750 134.020 177.550 134.030 ;
        RECT 1.270 133.830 3.480 134.000 ;
        RECT -150.440 129.350 -142.910 129.900 ;
        RECT -152.120 116.380 -150.650 116.630 ;
        RECT -150.440 116.440 -149.930 129.350 ;
        RECT -143.580 129.340 -142.910 129.350 ;
        RECT -147.280 128.450 -143.820 128.890 ;
        RECT -149.210 128.350 -143.820 128.450 ;
        RECT -149.210 128.280 -143.930 128.350 ;
        RECT -149.210 117.370 -149.040 128.280 ;
        RECT -148.710 127.870 -144.480 127.890 ;
        RECT -148.730 117.760 -144.400 127.870 ;
        RECT -148.670 117.710 -148.500 117.760 ;
        RECT -144.100 117.370 -143.930 128.280 ;
        RECT -149.210 117.200 -143.930 117.370 ;
        RECT -144.170 117.190 -143.930 117.200 ;
        RECT -143.420 116.440 -142.910 129.340 ;
        RECT 206.500 128.630 214.030 129.180 ;
        RECT 206.500 128.620 207.170 128.630 ;
        RECT -23.810 127.490 -23.640 127.790 ;
        RECT -23.810 127.310 -22.810 127.490 ;
        RECT -22.410 127.480 -22.240 127.790 ;
        RECT -20.610 127.520 -19.940 127.690 ;
        RECT -22.410 127.310 -21.400 127.480 ;
        RECT -20.610 126.730 -19.940 126.900 ;
        RECT -22.600 126.630 -22.280 126.670 ;
        RECT -23.480 126.460 -21.400 126.630 ;
        RECT -6.590 126.590 -3.280 127.570 ;
        RECT 0.810 126.770 1.040 127.460 ;
        RECT 5.510 126.720 5.740 127.410 ;
        RECT -22.610 126.440 -22.280 126.460 ;
        RECT -22.600 126.410 -22.280 126.440 ;
        RECT -23.300 126.050 -21.480 126.220 ;
        RECT -22.600 125.810 -22.280 125.830 ;
        RECT -23.480 125.640 -21.400 125.810 ;
        RECT -20.690 125.800 -20.480 126.230 ;
        RECT -6.480 125.930 -6.310 126.280 ;
        RECT -5.760 126.010 -5.590 126.040 ;
        RECT -5.850 125.970 -5.530 126.010 ;
        RECT -5.080 126.000 -4.910 126.040 ;
        RECT -7.210 125.890 -6.310 125.930 ;
        RECT -20.670 125.780 -20.500 125.800 ;
        RECT -7.220 125.700 -6.310 125.890 ;
        RECT -5.860 125.780 -5.530 125.970 ;
        RECT -5.160 125.960 -4.840 126.000 ;
        RECT -5.850 125.750 -5.530 125.780 ;
        RECT -5.170 125.770 -4.840 125.960 ;
        RECT -5.760 125.710 -5.590 125.750 ;
        RECT -5.160 125.740 -4.840 125.770 ;
        RECT -5.080 125.710 -4.910 125.740 ;
        RECT -7.210 125.670 -6.310 125.700 ;
        RECT 2.020 125.690 2.190 125.710 ;
        RECT -22.610 125.600 -22.280 125.640 ;
        RECT -22.600 125.570 -22.280 125.600 ;
        RECT -20.610 125.300 -19.940 125.470 ;
        RECT -23.480 124.800 -22.810 124.970 ;
        RECT -22.080 124.800 -21.400 124.970 ;
        RECT -21.100 124.680 -20.910 124.740 ;
        RECT -21.100 124.510 -19.930 124.680 ;
        RECT -21.170 124.230 -21.000 124.260 ;
        RECT -21.170 124.200 -20.840 124.230 ;
        RECT -21.170 124.010 -20.830 124.200 ;
        RECT -21.170 123.970 -20.840 124.010 ;
        RECT -21.170 123.930 -21.000 123.970 ;
        RECT -22.420 123.850 -22.250 123.910 ;
        RECT -20.600 123.900 -19.930 124.070 ;
        RECT -23.480 123.680 -22.810 123.850 ;
        RECT -22.420 123.680 -21.400 123.850 ;
        RECT -22.420 123.580 -22.250 123.680 ;
        RECT -22.620 123.010 -22.300 123.030 ;
        RECT -21.190 123.010 -20.870 123.050 ;
        RECT -23.490 122.840 -19.910 123.010 ;
        RECT -22.630 122.800 -22.300 122.840 ;
        RECT -21.200 122.820 -20.870 122.840 ;
        RECT -22.620 122.770 -22.300 122.800 ;
        RECT -21.190 122.790 -20.870 122.820 ;
        RECT -23.410 122.410 -23.090 122.450 ;
        RECT -22.480 122.410 -22.160 122.450 ;
        RECT -21.780 122.410 -21.460 122.450 ;
        RECT -21.040 122.410 -20.720 122.450 ;
        RECT -23.420 122.340 -23.090 122.410 ;
        RECT -22.490 122.340 -22.160 122.410 ;
        RECT -21.790 122.340 -21.460 122.410 ;
        RECT -21.050 122.390 -20.720 122.410 ;
        RECT -20.330 122.400 -20.010 122.440 ;
        RECT -20.340 122.390 -20.010 122.400 ;
        RECT -21.050 122.340 -20.010 122.390 ;
        RECT -23.440 122.170 -20.010 122.340 ;
        RECT -18.340 122.230 -18.170 122.900 ;
        RECT -7.850 122.810 -7.680 125.460 ;
        RECT -6.480 125.270 -6.310 125.670 ;
        RECT -0.870 125.520 2.190 125.690 ;
        RECT 2.020 124.870 2.190 125.520 ;
        RECT -6.590 123.790 -3.280 124.770 ;
        RECT 2.020 124.700 3.290 124.870 ;
        RECT 0.810 123.780 1.040 124.470 ;
        RECT -7.850 122.270 -7.670 122.810 ;
        RECT -7.930 122.230 -7.610 122.270 ;
        RECT -6.590 122.240 -3.280 123.220 ;
        RECT 0.810 122.770 1.040 123.460 ;
        RECT 2.020 122.290 2.190 124.700 ;
        RECT 4.760 123.050 4.930 123.940 ;
        RECT 1.930 122.250 2.250 122.290 ;
        RECT -20.860 122.160 -20.010 122.170 ;
        RECT -7.940 122.040 -7.610 122.230 ;
        RECT 1.920 122.060 2.250 122.250 ;
        RECT -7.930 122.010 -7.610 122.040 ;
        RECT 1.930 122.030 2.250 122.060 ;
        RECT -7.900 118.450 -6.380 118.460 ;
        RECT -7.900 117.660 -6.350 118.450 ;
        RECT -150.440 115.930 -142.910 116.440 ;
        RECT 12.980 116.260 13.330 116.360 ;
        RECT 16.050 116.340 18.280 116.490 ;
        RECT 16.050 116.320 18.430 116.340 ;
        RECT 16.050 116.310 16.230 116.320 ;
        RECT 15.590 116.290 16.230 116.310 ;
        RECT 14.640 116.260 15.100 116.290 ;
        RECT 11.570 116.090 12.330 116.260 ;
        RECT 12.580 116.090 13.750 116.260 ;
        RECT 13.990 116.120 15.100 116.260 ;
        RECT 15.550 116.120 16.230 116.290 ;
        RECT 17.830 116.170 18.430 116.320 ;
        RECT 18.890 116.160 19.220 116.330 ;
        RECT 13.990 116.090 14.810 116.120 ;
        RECT 11.570 116.080 11.800 116.090 ;
        RECT -152.140 109.910 -150.680 109.950 ;
        RECT -152.140 109.740 -150.670 109.910 ;
        RECT -152.140 109.700 -150.680 109.740 ;
        RECT -150.440 103.320 -149.930 115.930 ;
        RECT -149.570 115.140 -143.590 115.370 ;
        RECT -149.480 104.080 -143.830 115.140 ;
        RECT -143.420 105.570 -142.910 115.930 ;
        RECT 11.530 115.640 11.800 116.080 ;
        RECT 14.550 115.950 14.810 116.090 ;
        RECT 16.050 116.060 16.230 116.120 ;
        RECT 17.170 115.970 17.500 116.140 ;
        RECT 13.010 115.640 13.340 115.900 ;
        RECT 14.550 115.780 15.730 115.950 ;
        RECT 14.550 115.640 14.810 115.780 ;
        RECT 10.980 115.500 11.150 115.560 ;
        RECT 10.950 115.280 11.170 115.500 ;
        RECT 11.500 115.460 11.830 115.640 ;
        RECT 12.080 115.470 14.240 115.640 ;
        RECT 14.480 115.470 14.810 115.640 ;
        RECT 14.640 115.420 14.810 115.470 ;
        RECT 15.100 115.280 15.310 115.610 ;
        RECT 15.550 115.340 15.730 115.780 ;
        RECT 17.250 115.720 17.500 115.970 ;
        RECT 17.250 115.620 17.720 115.720 ;
        RECT 18.970 115.700 19.150 116.160 ;
        RECT 17.080 115.610 17.720 115.620 ;
        RECT 16.280 115.550 17.720 115.610 ;
        RECT 16.280 115.440 17.640 115.550 ;
        RECT 18.190 115.530 19.150 115.700 ;
        RECT 206.500 115.720 207.010 128.620 ;
        RECT 207.410 127.730 210.870 128.170 ;
        RECT 207.410 127.630 212.800 127.730 ;
        RECT 207.520 127.560 212.800 127.630 ;
        RECT 207.520 116.650 207.690 127.560 ;
        RECT 208.070 127.150 212.300 127.170 ;
        RECT 207.990 117.040 212.320 127.150 ;
        RECT 212.090 116.990 212.260 117.040 ;
        RECT 212.630 116.650 212.800 127.560 ;
        RECT 207.520 116.480 212.800 116.650 ;
        RECT 207.520 116.470 207.760 116.480 ;
        RECT 213.520 115.720 214.030 128.630 ;
        RECT 10.980 115.230 11.150 115.280 ;
        RECT 12.980 114.710 13.330 114.810 ;
        RECT 16.050 114.790 18.280 114.940 ;
        RECT 16.050 114.770 18.430 114.790 ;
        RECT 16.050 114.760 16.230 114.770 ;
        RECT 15.590 114.740 16.230 114.760 ;
        RECT 14.640 114.710 15.100 114.740 ;
        RECT 11.570 114.540 12.330 114.710 ;
        RECT 12.580 114.540 13.750 114.710 ;
        RECT 13.990 114.570 15.100 114.710 ;
        RECT 15.550 114.570 16.230 114.740 ;
        RECT 17.830 114.620 18.430 114.770 ;
        RECT 18.890 114.610 19.220 114.780 ;
        RECT 13.990 114.540 14.810 114.570 ;
        RECT 11.570 114.530 11.800 114.540 ;
        RECT 11.530 114.090 11.800 114.530 ;
        RECT 14.550 114.400 14.810 114.540 ;
        RECT 16.050 114.510 16.230 114.570 ;
        RECT 17.170 114.420 17.500 114.590 ;
        RECT 13.010 114.090 13.340 114.350 ;
        RECT 14.550 114.230 15.730 114.400 ;
        RECT 14.550 114.090 14.810 114.230 ;
        RECT 10.980 113.950 11.150 114.010 ;
        RECT 10.950 113.730 11.170 113.950 ;
        RECT 11.500 113.910 11.830 114.090 ;
        RECT 12.080 113.920 14.240 114.090 ;
        RECT 14.480 113.920 14.810 114.090 ;
        RECT 14.640 113.870 14.810 113.920 ;
        RECT 15.100 113.730 15.310 114.060 ;
        RECT 15.550 113.790 15.730 114.230 ;
        RECT 17.250 114.170 17.500 114.420 ;
        RECT 17.250 114.070 17.720 114.170 ;
        RECT 18.970 114.150 19.150 114.610 ;
        RECT 40.070 114.500 40.740 115.370 ;
        RECT 52.350 115.060 54.450 115.370 ;
        RECT 206.500 115.210 214.030 115.720 ;
        RECT 214.240 115.660 215.710 115.910 ;
        RECT 52.350 114.890 54.870 115.060 ;
        RECT 55.110 115.040 55.300 115.070 ;
        RECT 52.350 114.520 54.450 114.890 ;
        RECT 55.110 114.870 56.170 115.040 ;
        RECT 80.930 114.890 81.460 115.060 ;
        RECT 55.110 114.840 55.300 114.870 ;
        RECT 52.850 114.180 53.070 114.520 ;
        RECT 52.850 114.170 53.060 114.180 ;
        RECT 17.080 114.060 17.720 114.070 ;
        RECT 16.280 114.000 17.720 114.060 ;
        RECT 16.280 113.890 17.640 114.000 ;
        RECT 18.190 113.980 19.150 114.150 ;
        RECT 53.230 114.000 53.420 114.010 ;
        RECT 10.980 113.680 11.150 113.730 ;
        RECT 53.220 113.710 53.420 114.000 ;
        RECT 12.980 113.160 13.330 113.260 ;
        RECT 16.050 113.240 18.280 113.390 ;
        RECT 53.190 113.380 53.430 113.710 ;
        RECT 16.050 113.220 18.430 113.240 ;
        RECT 16.050 113.210 16.230 113.220 ;
        RECT 15.590 113.190 16.230 113.210 ;
        RECT 14.640 113.160 15.100 113.190 ;
        RECT -9.690 113.030 -9.490 113.070 ;
        RECT -10.000 112.770 -9.490 113.030 ;
        RECT -9.690 112.740 -9.490 112.770 ;
        RECT -9.100 113.040 -8.900 113.070 ;
        RECT -9.100 113.000 -8.590 113.040 ;
        RECT -9.100 112.810 -8.580 113.000 ;
        RECT 11.570 112.990 12.330 113.160 ;
        RECT 12.580 112.990 13.750 113.160 ;
        RECT 13.990 113.020 15.100 113.160 ;
        RECT 15.550 113.020 16.230 113.190 ;
        RECT 17.830 113.070 18.430 113.220 ;
        RECT 18.890 113.060 19.220 113.230 ;
        RECT 13.990 112.990 14.810 113.020 ;
        RECT 11.570 112.980 11.800 112.990 ;
        RECT -9.100 112.780 -8.590 112.810 ;
        RECT -9.100 112.740 -8.900 112.780 ;
        RECT -8.410 112.590 -8.240 112.640 ;
        RECT -10.440 112.570 -10.010 112.590 ;
        RECT -10.440 112.400 -9.990 112.570 ;
        RECT -8.420 112.560 -8.240 112.590 ;
        RECT -8.420 112.550 -7.990 112.560 ;
        RECT -10.440 112.380 -10.010 112.400 ;
        RECT -8.420 112.320 -7.830 112.550 ;
        RECT 11.530 112.540 11.800 112.980 ;
        RECT 14.550 112.850 14.810 112.990 ;
        RECT 16.050 112.960 16.230 113.020 ;
        RECT 17.170 112.870 17.500 113.040 ;
        RECT 13.010 112.540 13.340 112.800 ;
        RECT 14.550 112.680 15.730 112.850 ;
        RECT 14.550 112.540 14.810 112.680 ;
        RECT 10.980 112.400 11.150 112.460 ;
        RECT -8.420 112.310 -7.990 112.320 ;
        RECT -8.420 112.250 -8.250 112.310 ;
        RECT 10.950 112.180 11.170 112.400 ;
        RECT 11.500 112.360 11.830 112.540 ;
        RECT 12.080 112.370 14.240 112.540 ;
        RECT 14.480 112.370 14.810 112.540 ;
        RECT 14.640 112.320 14.810 112.370 ;
        RECT 15.100 112.180 15.310 112.510 ;
        RECT 15.550 112.240 15.730 112.680 ;
        RECT 17.250 112.620 17.500 112.870 ;
        RECT 17.250 112.520 17.720 112.620 ;
        RECT 18.970 112.600 19.150 113.060 ;
        RECT 53.620 112.900 53.790 114.510 ;
        RECT 54.450 113.410 54.620 114.500 ;
        RECT 55.580 114.480 55.770 114.510 ;
        RECT 55.040 114.310 55.770 114.480 ;
        RECT 56.000 114.480 56.170 114.870 ;
        RECT 82.740 114.790 82.940 115.140 ;
        RECT 82.740 114.760 82.950 114.790 ;
        RECT 56.000 114.310 56.740 114.480 ;
        RECT 79.060 114.310 79.410 114.480 ;
        RECT 80.430 114.310 80.760 114.480 ;
        RECT 55.580 114.280 55.770 114.310 ;
        RECT 57.800 113.690 58.030 114.210 ;
        RECT 55.040 113.520 58.030 113.690 ;
        RECT 54.220 113.370 54.620 113.410 ;
        RECT 54.210 113.180 54.620 113.370 ;
        RECT 63.000 113.330 63.550 113.760 ;
        RECT 72.250 113.330 72.800 113.760 ;
        RECT 75.880 113.520 76.110 114.210 ;
        RECT 81.180 113.980 81.350 114.500 ;
        RECT 81.020 113.720 81.350 113.980 ;
        RECT 79.060 113.520 79.410 113.690 ;
        RECT 80.430 113.520 80.760 113.690 ;
        RECT 54.220 113.150 54.620 113.180 ;
        RECT 53.610 112.710 53.790 112.900 ;
        RECT 54.450 112.810 54.620 113.150 ;
        RECT 55.110 112.900 55.300 113.080 ;
        RECT 55.040 112.730 55.390 112.900 ;
        RECT 17.080 112.510 17.720 112.520 ;
        RECT 16.280 112.450 17.720 112.510 ;
        RECT 16.280 112.340 17.640 112.450 ;
        RECT 18.190 112.430 19.150 112.600 ;
        RECT 55.960 112.320 56.170 112.750 ;
        RECT 56.390 112.730 56.730 112.900 ;
        RECT 55.980 112.300 56.150 112.320 ;
        RECT -9.690 112.110 -9.490 112.150 ;
        RECT -10.000 111.850 -9.490 112.110 ;
        RECT -9.690 111.820 -9.490 111.850 ;
        RECT -9.100 112.120 -8.900 112.150 ;
        RECT 10.980 112.130 11.150 112.180 ;
        RECT -9.100 112.080 -8.590 112.120 ;
        RECT -9.100 111.890 -8.580 112.080 ;
        RECT 53.610 111.990 53.790 112.180 ;
        RECT -9.100 111.860 -8.590 111.890 ;
        RECT -9.100 111.820 -8.900 111.860 ;
        RECT -10.440 111.650 -10.010 111.670 ;
        RECT -10.440 111.480 -9.990 111.650 ;
        RECT 12.980 111.610 13.330 111.710 ;
        RECT 16.050 111.690 18.280 111.840 ;
        RECT 16.050 111.670 18.430 111.690 ;
        RECT 16.050 111.660 16.230 111.670 ;
        RECT 15.590 111.640 16.230 111.660 ;
        RECT 14.640 111.610 15.100 111.640 ;
        RECT -10.440 111.460 -10.010 111.480 ;
        RECT 11.570 111.440 12.330 111.610 ;
        RECT 12.580 111.440 13.750 111.610 ;
        RECT 13.990 111.470 15.100 111.610 ;
        RECT 15.550 111.470 16.230 111.640 ;
        RECT 17.830 111.520 18.430 111.670 ;
        RECT 18.890 111.510 19.220 111.680 ;
        RECT 13.990 111.440 14.810 111.470 ;
        RECT 11.570 111.430 11.800 111.440 ;
        RECT -9.690 111.190 -9.490 111.230 ;
        RECT -10.000 110.930 -9.490 111.190 ;
        RECT -9.690 110.900 -9.490 110.930 ;
        RECT -9.100 111.200 -8.900 111.230 ;
        RECT -9.100 111.160 -8.590 111.200 ;
        RECT -9.100 110.970 -8.580 111.160 ;
        RECT 11.530 110.990 11.800 111.430 ;
        RECT 14.550 111.300 14.810 111.440 ;
        RECT 16.050 111.410 16.230 111.470 ;
        RECT 17.170 111.320 17.500 111.490 ;
        RECT 13.010 110.990 13.340 111.250 ;
        RECT 14.550 111.130 15.730 111.300 ;
        RECT 14.550 110.990 14.810 111.130 ;
        RECT -9.100 110.940 -8.590 110.970 ;
        RECT -9.100 110.900 -8.900 110.940 ;
        RECT 10.980 110.850 11.150 110.910 ;
        RECT -10.440 110.730 -10.010 110.750 ;
        RECT -10.440 110.560 -9.990 110.730 ;
        RECT 10.950 110.630 11.170 110.850 ;
        RECT 11.500 110.810 11.830 110.990 ;
        RECT 12.080 110.820 14.240 110.990 ;
        RECT 14.480 110.820 14.810 110.990 ;
        RECT 14.640 110.770 14.810 110.820 ;
        RECT 15.100 110.630 15.310 110.960 ;
        RECT 15.550 110.690 15.730 111.130 ;
        RECT 17.250 111.070 17.500 111.320 ;
        RECT 17.250 110.970 17.720 111.070 ;
        RECT 18.970 111.050 19.150 111.510 ;
        RECT 53.190 111.180 53.430 111.510 ;
        RECT 17.080 110.960 17.720 110.970 ;
        RECT 16.280 110.900 17.720 110.960 ;
        RECT 16.280 110.790 17.640 110.900 ;
        RECT 18.190 110.880 19.150 111.050 ;
        RECT 53.220 110.890 53.420 111.180 ;
        RECT 53.230 110.880 53.420 110.890 ;
        RECT 52.850 110.710 53.060 110.720 ;
        RECT 10.980 110.580 11.150 110.630 ;
        RECT -10.440 110.540 -10.010 110.560 ;
        RECT -10.190 110.170 -9.870 110.210 ;
        RECT -10.190 110.150 -9.860 110.170 ;
        RECT 22.730 110.160 22.930 110.510 ;
        RECT 24.210 110.260 24.740 110.430 ;
        RECT -10.190 109.950 -9.570 110.150 ;
        RECT -9.740 109.820 -9.570 109.950 ;
        RECT -9.060 110.110 -8.890 110.150 ;
        RECT 22.720 110.130 22.930 110.160 ;
        RECT -9.060 110.070 -8.570 110.110 ;
        RECT -9.060 109.880 -8.560 110.070 ;
        RECT -9.060 109.850 -8.570 109.880 ;
        RECT -9.060 109.820 -8.890 109.850 ;
        RECT -10.350 109.710 -9.920 109.730 ;
        RECT -10.370 109.540 -9.920 109.710 ;
        RECT 22.720 109.550 22.940 110.130 ;
        RECT 22.720 109.540 22.930 109.550 ;
        RECT -10.350 109.520 -9.920 109.540 ;
        RECT 23.100 109.370 23.290 109.380 ;
        RECT -10.190 109.210 -9.870 109.250 ;
        RECT -10.190 109.190 -9.860 109.210 ;
        RECT -10.190 108.990 -9.570 109.190 ;
        RECT -9.740 108.860 -9.570 108.990 ;
        RECT -9.060 109.150 -8.890 109.190 ;
        RECT -9.060 109.110 -8.570 109.150 ;
        RECT -9.060 108.920 -8.560 109.110 ;
        RECT 23.090 109.080 23.290 109.370 ;
        RECT 10.980 109.030 11.150 109.080 ;
        RECT -9.060 108.890 -8.570 108.920 ;
        RECT -9.060 108.860 -8.890 108.890 ;
        RECT 10.950 108.810 11.170 109.030 ;
        RECT -10.350 108.750 -9.920 108.770 ;
        RECT 10.980 108.750 11.150 108.810 ;
        RECT -10.370 108.580 -9.920 108.750 ;
        RECT 11.500 108.670 11.830 108.850 ;
        RECT 14.640 108.840 14.810 108.890 ;
        RECT 12.080 108.670 14.240 108.840 ;
        RECT 14.480 108.670 14.810 108.840 ;
        RECT 15.100 108.700 15.310 109.030 ;
        RECT -10.350 108.560 -9.920 108.580 ;
        RECT -10.190 108.250 -9.870 108.290 ;
        RECT -10.190 108.230 -9.860 108.250 ;
        RECT 11.530 108.230 11.800 108.670 ;
        RECT 13.010 108.410 13.340 108.670 ;
        RECT 14.550 108.530 14.810 108.670 ;
        RECT 15.550 108.530 15.730 108.970 ;
        RECT 16.280 108.760 17.640 108.870 ;
        RECT 16.280 108.700 17.720 108.760 ;
        RECT 17.080 108.690 17.720 108.700 ;
        RECT -10.190 108.030 -9.570 108.230 ;
        RECT -9.740 107.900 -9.570 108.030 ;
        RECT -9.060 108.190 -8.890 108.230 ;
        RECT 11.570 108.220 11.800 108.230 ;
        RECT 14.550 108.360 15.730 108.530 ;
        RECT 17.250 108.590 17.720 108.690 ;
        RECT 18.190 108.610 19.150 108.780 ;
        RECT 23.060 108.750 23.300 109.080 ;
        RECT 14.550 108.220 14.810 108.360 ;
        RECT 17.250 108.340 17.500 108.590 ;
        RECT -9.060 108.150 -8.570 108.190 ;
        RECT -9.060 107.960 -8.560 108.150 ;
        RECT 11.570 108.050 12.330 108.220 ;
        RECT 12.580 108.050 13.750 108.220 ;
        RECT 13.990 108.190 14.810 108.220 ;
        RECT 16.050 108.190 16.230 108.250 ;
        RECT 13.990 108.050 15.100 108.190 ;
        RECT -9.060 107.930 -8.570 107.960 ;
        RECT 12.980 107.950 13.330 108.050 ;
        RECT 14.640 108.020 15.100 108.050 ;
        RECT 15.550 108.020 16.230 108.190 ;
        RECT 17.170 108.170 17.500 108.340 ;
        RECT 18.970 108.150 19.150 108.610 ;
        RECT 23.490 108.270 23.660 109.880 ;
        RECT 15.590 108.000 16.230 108.020 ;
        RECT 16.050 107.990 16.230 108.000 ;
        RECT 17.830 107.990 18.430 108.140 ;
        RECT 16.050 107.970 18.430 107.990 ;
        RECT 18.890 107.980 19.220 108.150 ;
        RECT 23.480 108.080 23.660 108.270 ;
        RECT 24.320 109.350 24.490 109.870 ;
        RECT 24.910 109.680 25.240 109.850 ;
        RECT 26.260 109.680 26.610 109.850 ;
        RECT 26.930 109.830 31.990 110.660 ;
        RECT 50.810 110.260 51.340 110.430 ;
        RECT 52.620 110.160 52.820 110.510 ;
        RECT 52.620 110.130 52.830 110.160 ;
        RECT 31.440 109.750 31.920 109.830 ;
        RECT 24.320 109.090 24.650 109.350 ;
        RECT 24.320 108.180 24.490 109.090 ;
        RECT 24.910 108.890 25.240 109.060 ;
        RECT 26.260 108.890 26.610 109.060 ;
        RECT 29.560 108.890 29.790 109.580 ;
        RECT 31.440 109.500 31.910 109.750 ;
        RECT 48.940 109.680 49.290 109.850 ;
        RECT 50.310 109.680 50.640 109.850 ;
        RECT 30.750 108.990 30.920 109.410 ;
        RECT 31.560 109.290 31.800 109.320 ;
        RECT 31.230 109.120 31.800 109.290 ;
        RECT 32.040 109.130 33.380 109.290 ;
        RECT 32.040 109.120 33.420 109.130 ;
        RECT 33.830 109.120 34.790 109.290 ;
        RECT 31.560 109.080 31.800 109.120 ;
        RECT 30.680 108.770 30.850 108.810 ;
        RECT 30.620 108.600 30.850 108.770 ;
        RECT 32.870 108.700 33.420 109.120 ;
        RECT 34.340 109.110 34.510 109.120 ;
        RECT 30.680 108.270 30.850 108.600 ;
        RECT 31.020 108.670 31.210 108.690 ;
        RECT 34.020 108.670 34.350 108.850 ;
        RECT 31.020 108.500 31.580 108.670 ;
        RECT 32.040 108.500 34.790 108.670 ;
        RECT 31.020 108.460 31.210 108.500 ;
        RECT 35.320 108.430 35.490 109.360 ;
        RECT 35.720 108.560 35.890 109.410 ;
        RECT 42.130 108.700 42.680 109.130 ;
        RECT 45.760 108.890 45.990 109.580 ;
        RECT 51.060 109.350 51.230 109.870 ;
        RECT 50.900 109.090 51.230 109.350 ;
        RECT 48.940 108.890 49.290 109.060 ;
        RECT 50.310 108.890 50.640 109.060 ;
        RECT 24.910 108.100 25.240 108.270 ;
        RECT 26.260 108.100 26.600 108.270 ;
        RECT 30.630 108.250 30.850 108.270 ;
        RECT -9.060 107.900 -8.890 107.930 ;
        RECT 16.050 107.820 18.280 107.970 ;
        RECT -10.350 107.790 -9.920 107.810 ;
        RECT -10.370 107.620 -9.920 107.790 ;
        RECT -10.350 107.600 -9.920 107.620 ;
        RECT -8.560 107.560 -8.140 107.730 ;
        RECT -8.460 107.520 -8.230 107.560 ;
        RECT 10.980 107.480 11.150 107.530 ;
        RECT 10.950 107.260 11.170 107.480 ;
        RECT 10.980 107.200 11.150 107.260 ;
        RECT 11.500 107.120 11.830 107.300 ;
        RECT 14.640 107.290 14.810 107.340 ;
        RECT 12.080 107.120 14.240 107.290 ;
        RECT 14.480 107.120 14.810 107.290 ;
        RECT 15.100 107.150 15.310 107.480 ;
        RECT 11.530 106.680 11.800 107.120 ;
        RECT 13.010 106.860 13.340 107.120 ;
        RECT 14.550 106.980 14.810 107.120 ;
        RECT 15.550 106.980 15.730 107.420 ;
        RECT 23.480 107.360 23.660 107.550 ;
        RECT 24.990 107.530 25.160 108.100 ;
        RECT 30.630 108.010 30.820 108.250 ;
        RECT 30.630 107.870 30.850 108.010 ;
        RECT 44.730 107.870 44.920 108.270 ;
        RECT 48.950 108.100 49.290 108.270 ;
        RECT 50.310 108.100 50.640 108.270 ;
        RECT 51.060 108.180 51.230 109.090 ;
        RECT 51.890 108.270 52.060 109.880 ;
        RECT 52.610 109.550 52.830 110.130 ;
        RECT 52.850 110.130 53.070 110.710 ;
        RECT 53.620 110.380 53.790 111.990 ;
        RECT 54.450 111.720 54.620 112.080 ;
        RECT 55.040 111.990 55.390 112.160 ;
        RECT 55.580 112.140 55.770 112.190 ;
        RECT 56.480 112.160 56.650 112.730 ;
        RECT 60.760 112.500 60.950 112.900 ;
        RECT 74.850 112.500 75.040 112.900 ;
        RECT 79.070 112.730 79.410 112.900 ;
        RECT 80.430 112.730 80.760 112.900 ;
        RECT 81.180 112.810 81.350 113.720 ;
        RECT 82.010 112.900 82.180 114.510 ;
        RECT 82.730 114.180 82.950 114.760 ;
        RECT 82.740 114.170 82.950 114.180 ;
        RECT 82.380 114.000 82.570 114.010 ;
        RECT 82.380 113.710 82.580 114.000 ;
        RECT 82.370 113.380 82.610 113.710 ;
        RECT 60.760 112.490 61.140 112.500 ;
        RECT 57.400 112.310 61.140 112.490 ;
        RECT 60.760 112.270 61.140 112.310 ;
        RECT 74.660 112.490 75.040 112.500 ;
        RECT 74.660 112.310 78.400 112.490 ;
        RECT 74.660 112.270 75.040 112.310 ;
        RECT 55.580 112.130 55.810 112.140 ;
        RECT 56.390 112.130 56.730 112.160 ;
        RECT 55.580 111.990 56.730 112.130 ;
        RECT 55.120 111.780 55.310 111.990 ;
        RECT 55.580 111.960 56.560 111.990 ;
        RECT 55.720 111.930 56.560 111.960 ;
        RECT 60.760 111.890 60.950 112.270 ;
        RECT 54.210 111.680 54.620 111.720 ;
        RECT 54.200 111.490 54.620 111.680 ;
        RECT 63.000 111.600 63.550 112.030 ;
        RECT 72.250 111.600 72.800 112.030 ;
        RECT 74.850 111.890 75.040 112.270 ;
        RECT 80.510 112.160 80.680 112.730 ;
        RECT 82.010 112.710 82.190 112.900 ;
        RECT 79.070 111.990 79.410 112.160 ;
        RECT 80.430 111.990 80.760 112.160 ;
        RECT 80.360 111.600 80.530 111.650 ;
        RECT 54.210 111.460 54.620 111.490 ;
        RECT 54.450 110.390 54.620 111.460 ;
        RECT 55.040 111.270 57.970 111.370 ;
        RECT 55.040 111.200 58.030 111.270 ;
        RECT 57.060 110.880 57.230 110.940 ;
        RECT 57.040 110.670 57.250 110.880 ;
        RECT 55.570 110.580 55.760 110.610 ;
        RECT 57.060 110.600 57.230 110.670 ;
        RECT 57.800 110.580 58.030 111.200 ;
        RECT 75.880 110.580 76.110 111.310 ;
        RECT 79.060 111.200 79.410 111.370 ;
        RECT 80.360 111.340 80.920 111.600 ;
        RECT 80.360 111.320 80.760 111.340 ;
        RECT 80.430 111.200 80.760 111.320 ;
        RECT 81.180 111.220 81.350 112.080 ;
        RECT 82.010 111.990 82.190 112.180 ;
        RECT 82.010 111.360 82.180 111.990 ;
        RECT 81.830 111.320 82.180 111.360 ;
        RECT 55.040 110.410 55.760 110.580 ;
        RECT 55.570 110.380 55.760 110.410 ;
        RECT 55.930 110.410 56.740 110.580 ;
        RECT 79.060 110.410 79.410 110.580 ;
        RECT 52.850 110.100 53.060 110.130 ;
        RECT 52.860 109.750 53.060 110.100 ;
        RECT 55.140 110.070 55.330 110.100 ;
        RECT 55.930 110.070 56.120 110.410 ;
        RECT 79.780 110.240 79.960 111.170 ;
        RECT 80.510 110.910 80.840 111.080 ;
        RECT 81.020 110.960 81.350 111.220 ;
        RECT 81.600 111.060 82.180 111.320 ;
        RECT 82.370 111.360 82.610 111.510 ;
        RECT 82.370 111.180 82.970 111.360 ;
        RECT 81.830 111.030 82.180 111.060 ;
        RECT 80.590 110.770 80.840 110.910 ;
        RECT 80.590 110.580 81.070 110.770 ;
        RECT 80.430 110.510 81.070 110.580 ;
        RECT 80.430 110.410 80.760 110.510 ;
        RECT 79.660 110.210 79.980 110.240 ;
        RECT 80.590 110.210 80.760 110.410 ;
        RECT 81.180 110.390 81.350 110.960 ;
        RECT 81.420 110.670 81.590 110.710 ;
        RECT 82.010 110.700 82.180 111.030 ;
        RECT 82.380 110.880 82.970 111.180 ;
        RECT 83.790 111.240 84.370 111.410 ;
        RECT 83.790 111.140 84.180 111.240 ;
        RECT 83.790 111.110 84.170 111.140 ;
        RECT 83.790 110.960 84.150 111.110 ;
        RECT 81.830 110.670 82.180 110.700 ;
        RECT 81.420 110.410 82.180 110.670 ;
        RECT 81.420 110.380 81.590 110.410 ;
        RECT 81.830 110.380 82.180 110.410 ;
        RECT 81.830 110.370 82.030 110.380 ;
        RECT 82.420 110.370 82.970 110.880 ;
        RECT 83.440 110.790 84.150 110.960 ;
        RECT 79.190 110.180 79.510 110.210 ;
        RECT 54.340 109.830 54.870 110.000 ;
        RECT 55.140 109.890 56.120 110.070 ;
        RECT 55.140 109.870 55.330 109.890 ;
        RECT 77.970 109.840 78.140 110.120 ;
        RECT 79.190 109.990 79.520 110.180 ;
        RECT 79.660 110.040 79.990 110.210 ;
        RECT 80.590 110.180 81.080 110.210 ;
        RECT 80.200 110.040 80.390 110.060 ;
        RECT 79.190 109.950 79.510 109.990 ;
        RECT 79.660 109.980 80.390 110.040 ;
        RECT 77.970 109.800 78.180 109.840 ;
        RECT 77.970 109.780 78.200 109.800 ;
        RECT 79.320 109.790 79.490 109.950 ;
        RECT 79.780 109.870 80.390 109.980 ;
        RECT 77.970 109.760 78.230 109.780 ;
        RECT 77.970 109.710 78.310 109.760 ;
        RECT 77.970 109.650 78.460 109.710 ;
        RECT 77.970 109.620 78.480 109.650 ;
        RECT 78.010 109.590 78.480 109.620 ;
        RECT 52.620 109.540 52.830 109.550 ;
        RECT 78.140 109.540 78.480 109.590 ;
        RECT 79.780 109.540 79.960 109.870 ;
        RECT 80.180 109.860 80.390 109.870 ;
        RECT 80.200 109.830 80.390 109.860 ;
        RECT 80.590 110.000 81.090 110.180 ;
        RECT 82.730 110.130 82.950 110.370 ;
        RECT 81.330 110.040 81.520 110.070 ;
        RECT 81.330 110.000 81.770 110.040 ;
        RECT 80.590 109.950 81.770 110.000 ;
        RECT 78.260 109.530 78.480 109.540 ;
        RECT 78.270 109.500 78.480 109.530 ;
        RECT 78.290 109.420 78.480 109.500 ;
        RECT 79.650 109.420 79.980 109.540 ;
        RECT 80.590 109.420 80.760 109.950 ;
        RECT 80.820 109.870 81.770 109.950 ;
        RECT 80.820 109.840 81.590 109.870 ;
        RECT 81.830 109.840 82.030 109.880 ;
        RECT 80.820 109.830 82.030 109.840 ;
        RECT 80.820 109.790 80.990 109.830 ;
        RECT 81.420 109.580 82.030 109.830 ;
        RECT 81.420 109.540 81.590 109.580 ;
        RECT 81.830 109.550 82.030 109.580 ;
        RECT 82.050 109.450 82.220 110.130 ;
        RECT 82.740 110.100 82.950 110.130 ;
        RECT 82.740 109.880 82.940 110.100 ;
        RECT 83.440 110.040 84.140 110.350 ;
        RECT 52.260 109.370 52.450 109.380 ;
        RECT 77.800 109.370 77.970 109.390 ;
        RECT 52.260 109.080 52.460 109.370 ;
        RECT 52.250 108.750 52.490 109.080 ;
        RECT 77.780 108.940 77.990 109.370 ;
        RECT 78.290 109.250 78.810 109.420 ;
        RECT 78.290 109.220 78.480 109.250 ;
        RECT 79.160 109.240 81.060 109.420 ;
        RECT 81.790 109.410 82.220 109.450 ;
        RECT 81.440 109.250 82.220 109.410 ;
        RECT 81.440 109.240 81.980 109.250 ;
        RECT 77.780 108.300 77.990 108.730 ;
        RECT 78.290 108.420 78.480 108.450 ;
        RECT 79.780 108.430 79.960 109.240 ;
        RECT 80.590 109.130 80.760 109.240 ;
        RECT 81.790 109.220 81.980 109.240 ;
        RECT 81.830 109.190 82.030 109.220 ;
        RECT 80.390 108.930 80.710 108.960 ;
        RECT 81.600 108.930 82.030 109.190 ;
        RECT 80.390 108.740 80.720 108.930 ;
        RECT 81.830 108.890 82.030 108.930 ;
        RECT 82.420 108.890 82.970 109.880 ;
        RECT 83.290 109.810 84.140 110.040 ;
        RECT 83.440 109.470 84.140 109.810 ;
        RECT 83.900 109.110 84.220 109.150 ;
        RECT 83.900 109.050 84.230 109.110 ;
        RECT 83.430 108.920 84.230 109.050 ;
        RECT 83.430 108.890 84.220 108.920 ;
        RECT 83.430 108.870 84.130 108.890 ;
        RECT 80.390 108.700 80.710 108.740 ;
        RECT 80.390 108.620 80.560 108.700 ;
        RECT 80.340 108.450 80.560 108.620 ;
        RECT 80.340 108.430 80.510 108.450 ;
        RECT 81.790 108.430 81.980 108.450 ;
        RECT 77.800 108.280 77.970 108.300 ;
        RECT 30.630 107.860 31.010 107.870 ;
        RECT 27.270 107.680 31.010 107.860 ;
        RECT 44.540 107.860 44.920 107.870 ;
        RECT 30.630 107.660 31.010 107.680 ;
        RECT 30.620 107.640 31.010 107.660 ;
        RECT 31.020 107.760 31.210 107.800 ;
        RECT 16.280 107.210 17.640 107.320 ;
        RECT 16.280 107.150 17.720 107.210 ;
        RECT 17.080 107.140 17.720 107.150 ;
        RECT 11.570 106.670 11.800 106.680 ;
        RECT 14.550 106.810 15.730 106.980 ;
        RECT 17.250 107.040 17.720 107.140 ;
        RECT 18.190 107.060 19.150 107.230 ;
        RECT 14.550 106.670 14.810 106.810 ;
        RECT 17.250 106.790 17.500 107.040 ;
        RECT 11.570 106.500 12.330 106.670 ;
        RECT 12.580 106.500 13.750 106.670 ;
        RECT 13.990 106.640 14.810 106.670 ;
        RECT 16.050 106.640 16.230 106.700 ;
        RECT 13.990 106.500 15.100 106.640 ;
        RECT 12.980 106.400 13.330 106.500 ;
        RECT 14.640 106.470 15.100 106.500 ;
        RECT 15.550 106.470 16.230 106.640 ;
        RECT 17.170 106.620 17.500 106.790 ;
        RECT 18.970 106.600 19.150 107.060 ;
        RECT 15.590 106.450 16.230 106.470 ;
        RECT 16.050 106.440 16.230 106.450 ;
        RECT 17.830 106.440 18.430 106.590 ;
        RECT 16.050 106.420 18.430 106.440 ;
        RECT 18.890 106.430 19.220 106.600 ;
        RECT 23.060 106.550 23.300 106.880 ;
        RECT 16.050 106.270 18.280 106.420 ;
        RECT 23.090 106.260 23.290 106.550 ;
        RECT 23.100 106.250 23.290 106.260 ;
        RECT 22.720 106.080 22.930 106.090 ;
        RECT 10.980 105.930 11.150 105.980 ;
        RECT 10.950 105.710 11.170 105.930 ;
        RECT 10.980 105.650 11.150 105.710 ;
        RECT 11.500 105.570 11.830 105.750 ;
        RECT 14.640 105.740 14.810 105.790 ;
        RECT 12.080 105.570 14.240 105.740 ;
        RECT 14.480 105.570 14.810 105.740 ;
        RECT 15.100 105.600 15.310 105.930 ;
        RECT -143.430 105.550 -142.910 105.570 ;
        RECT -149.480 104.070 -143.770 104.080 ;
        RECT -149.560 103.900 -143.770 104.070 ;
        RECT -149.470 103.890 -143.770 103.900 ;
        RECT -144.000 103.820 -143.830 103.890 ;
        RECT -143.430 103.770 -142.900 105.550 ;
        RECT 11.530 105.130 11.800 105.570 ;
        RECT 13.010 105.310 13.340 105.570 ;
        RECT 14.550 105.430 14.810 105.570 ;
        RECT 15.550 105.430 15.730 105.870 ;
        RECT 16.280 105.660 17.640 105.770 ;
        RECT 16.280 105.600 17.720 105.660 ;
        RECT 17.080 105.590 17.720 105.600 ;
        RECT 11.570 105.120 11.800 105.130 ;
        RECT 14.550 105.260 15.730 105.430 ;
        RECT 17.250 105.490 17.720 105.590 ;
        RECT 18.190 105.510 19.150 105.680 ;
        RECT 14.550 105.120 14.810 105.260 ;
        RECT 17.250 105.240 17.500 105.490 ;
        RECT 11.570 104.950 12.330 105.120 ;
        RECT 12.580 104.950 13.750 105.120 ;
        RECT 13.990 105.090 14.810 105.120 ;
        RECT 16.050 105.090 16.230 105.150 ;
        RECT 13.990 104.950 15.100 105.090 ;
        RECT 12.980 104.850 13.330 104.950 ;
        RECT 14.640 104.920 15.100 104.950 ;
        RECT 15.550 104.920 16.230 105.090 ;
        RECT 17.170 105.070 17.500 105.240 ;
        RECT 18.970 105.050 19.150 105.510 ;
        RECT 22.720 105.500 22.940 106.080 ;
        RECT 23.490 105.750 23.660 107.360 ;
        RECT 24.320 106.590 24.490 107.450 ;
        RECT 24.910 107.360 25.240 107.530 ;
        RECT 26.260 107.360 26.600 107.530 ;
        RECT 30.620 107.490 30.850 107.640 ;
        RECT 31.020 107.590 31.580 107.760 ;
        RECT 32.040 107.590 34.790 107.760 ;
        RECT 31.020 107.570 31.210 107.590 ;
        RECT 30.630 107.450 30.850 107.490 ;
        RECT 30.630 107.270 30.820 107.450 ;
        RECT 34.020 107.410 34.350 107.590 ;
        RECT 30.630 107.260 30.920 107.270 ;
        RECT 30.750 106.850 30.920 107.260 ;
        RECT 31.560 107.140 31.800 107.180 ;
        RECT 32.870 107.140 33.420 107.400 ;
        RECT 34.340 107.140 34.510 107.150 ;
        RECT 31.230 106.970 31.800 107.140 ;
        RECT 32.040 106.970 33.420 107.140 ;
        RECT 33.830 106.970 34.790 107.140 ;
        RECT 31.560 106.940 31.800 106.970 ;
        RECT 35.320 106.900 35.490 107.830 ;
        RECT 35.720 106.850 35.890 107.700 ;
        RECT 44.540 107.680 48.280 107.860 ;
        RECT 44.540 107.640 44.920 107.680 ;
        RECT 42.130 106.970 42.680 107.400 ;
        RECT 44.730 107.260 44.920 107.640 ;
        RECT 50.390 107.530 50.560 108.100 ;
        RECT 51.890 108.080 52.070 108.270 ;
        RECT 78.290 108.250 78.810 108.420 ;
        RECT 79.160 108.250 81.060 108.430 ;
        RECT 81.440 108.420 81.980 108.430 ;
        RECT 81.440 108.260 82.220 108.420 ;
        RECT 78.290 108.170 78.480 108.250 ;
        RECT 78.270 108.140 78.480 108.170 ;
        RECT 78.260 108.130 78.480 108.140 ;
        RECT 79.650 108.130 79.980 108.250 ;
        RECT 81.600 108.220 82.220 108.260 ;
        RECT 78.140 108.080 78.480 108.130 ;
        RECT 78.010 108.050 78.480 108.080 ;
        RECT 77.970 108.020 78.480 108.050 ;
        RECT 77.970 107.960 78.460 108.020 ;
        RECT 77.970 107.910 78.310 107.960 ;
        RECT 77.970 107.890 78.230 107.910 ;
        RECT 77.970 107.870 78.200 107.890 ;
        RECT 77.970 107.830 78.180 107.870 ;
        RECT 77.970 107.550 78.140 107.830 ;
        RECT 79.320 107.720 79.490 107.880 ;
        RECT 79.780 107.800 79.960 108.130 ;
        RECT 80.870 108.030 81.060 108.150 ;
        RECT 81.600 108.100 82.030 108.220 ;
        RECT 81.830 108.070 82.030 108.100 ;
        RECT 80.510 107.920 81.060 108.030 ;
        RECT 80.510 107.860 81.050 107.920 ;
        RECT 80.200 107.810 80.390 107.840 ;
        RECT 80.180 107.800 80.390 107.810 ;
        RECT 79.190 107.680 79.510 107.720 ;
        RECT 48.950 107.360 49.290 107.530 ;
        RECT 50.310 107.360 50.640 107.530 ;
        RECT 50.240 106.970 50.410 107.020 ;
        RECT 24.320 106.330 24.650 106.590 ;
        RECT 24.910 106.570 25.240 106.740 ;
        RECT 26.260 106.570 26.610 106.740 ;
        RECT 24.320 105.760 24.490 106.330 ;
        RECT 29.560 105.950 29.790 106.680 ;
        RECT 30.750 106.060 30.920 106.480 ;
        RECT 31.560 106.360 31.800 106.390 ;
        RECT 31.230 106.190 31.800 106.360 ;
        RECT 32.040 106.190 33.380 106.360 ;
        RECT 33.830 106.190 34.790 106.360 ;
        RECT 31.560 106.150 31.800 106.190 ;
        RECT 34.340 106.180 34.510 106.190 ;
        RECT 24.910 105.780 25.240 105.950 ;
        RECT 26.260 105.780 26.610 105.950 ;
        RECT 30.680 105.840 30.850 105.880 ;
        RECT 30.620 105.740 30.850 105.840 ;
        RECT 31.600 105.820 31.940 106.070 ;
        RECT 31.020 105.740 31.210 105.760 ;
        RECT 31.600 105.740 31.950 105.820 ;
        RECT 34.020 105.740 34.350 105.920 ;
        RECT 22.720 105.470 22.930 105.500 ;
        RECT 22.730 105.120 22.930 105.470 ;
        RECT 24.210 105.200 24.740 105.370 ;
        RECT 15.590 104.900 16.230 104.920 ;
        RECT 16.050 104.890 16.230 104.900 ;
        RECT 17.830 104.890 18.430 105.040 ;
        RECT 16.050 104.870 18.430 104.890 ;
        RECT 18.890 104.880 19.220 105.050 ;
        RECT 26.900 104.890 31.950 105.740 ;
        RECT 32.040 105.570 34.790 105.740 ;
        RECT 35.320 105.500 35.490 106.430 ;
        RECT 35.720 105.630 35.890 106.480 ;
        RECT 45.760 105.950 45.990 106.680 ;
        RECT 48.940 106.570 49.290 106.740 ;
        RECT 50.240 106.710 50.800 106.970 ;
        RECT 50.240 106.690 50.640 106.710 ;
        RECT 50.310 106.570 50.640 106.690 ;
        RECT 51.060 106.590 51.230 107.450 ;
        RECT 51.890 107.360 52.070 107.550 ;
        RECT 79.190 107.490 79.520 107.680 ;
        RECT 79.780 107.630 80.390 107.800 ;
        RECT 79.190 107.460 79.510 107.490 ;
        RECT 51.890 106.730 52.060 107.360 ;
        RECT 79.190 107.160 79.510 107.190 ;
        RECT 51.710 106.690 52.060 106.730 ;
        RECT 48.940 105.780 49.290 105.950 ;
        RECT 49.660 105.610 49.840 106.540 ;
        RECT 50.390 106.280 50.720 106.450 ;
        RECT 50.900 106.330 51.230 106.590 ;
        RECT 51.480 106.430 52.060 106.690 ;
        RECT 52.250 106.730 52.490 106.880 ;
        RECT 77.970 106.820 78.140 107.100 ;
        RECT 79.190 106.970 79.520 107.160 ;
        RECT 79.780 107.020 79.960 107.630 ;
        RECT 80.200 107.610 80.390 107.630 ;
        RECT 80.590 107.720 80.760 107.860 ;
        RECT 80.820 107.720 80.990 107.860 ;
        RECT 81.330 107.800 81.520 107.830 ;
        RECT 80.590 107.680 81.080 107.720 ;
        RECT 81.330 107.710 81.770 107.800 ;
        RECT 81.830 107.710 82.030 107.740 ;
        RECT 80.590 107.490 81.090 107.680 ;
        RECT 81.330 107.600 82.030 107.710 ;
        RECT 80.590 107.460 81.080 107.490 ;
        RECT 80.590 107.190 80.760 107.460 ;
        RECT 81.420 107.450 82.030 107.600 ;
        RECT 82.050 107.540 82.220 108.220 ;
        RECT 81.420 107.420 81.590 107.450 ;
        RECT 81.830 107.410 82.030 107.450 ;
        RECT 82.420 107.410 82.970 108.400 ;
        RECT 83.890 108.390 84.210 108.430 ;
        RECT 83.430 108.210 84.220 108.390 ;
        RECT 83.890 108.200 84.220 108.210 ;
        RECT 83.890 108.170 84.210 108.200 ;
        RECT 83.440 107.450 84.140 107.790 ;
        RECT 83.290 107.220 84.140 107.450 ;
        RECT 80.590 107.160 81.080 107.190 ;
        RECT 80.200 107.020 80.390 107.040 ;
        RECT 79.190 106.930 79.510 106.970 ;
        RECT 77.970 106.780 78.180 106.820 ;
        RECT 52.250 106.550 52.850 106.730 ;
        RECT 51.710 106.400 52.060 106.430 ;
        RECT 50.470 106.140 50.720 106.280 ;
        RECT 50.470 105.950 50.950 106.140 ;
        RECT 50.310 105.880 50.950 105.950 ;
        RECT 50.310 105.780 50.640 105.880 ;
        RECT 49.540 105.580 49.860 105.610 ;
        RECT 49.540 105.390 49.870 105.580 ;
        RECT 49.540 105.350 49.860 105.390 ;
        RECT 16.050 104.720 18.280 104.870 ;
        RECT 30.680 104.730 30.850 104.890 ;
        RECT 30.620 104.560 30.850 104.730 ;
        RECT 31.020 104.830 31.210 104.870 ;
        RECT 31.020 104.660 31.580 104.830 ;
        RECT 32.040 104.660 34.790 104.830 ;
        RECT 31.020 104.640 31.210 104.660 ;
        RECT 30.680 104.520 30.850 104.560 ;
        RECT 34.020 104.480 34.350 104.660 ;
        RECT 10.980 104.380 11.150 104.430 ;
        RECT 10.950 104.160 11.170 104.380 ;
        RECT 10.980 104.100 11.150 104.160 ;
        RECT 11.500 104.020 11.830 104.200 ;
        RECT 14.640 104.190 14.810 104.240 ;
        RECT 12.080 104.020 14.240 104.190 ;
        RECT 14.480 104.020 14.810 104.190 ;
        RECT 15.100 104.050 15.310 104.380 ;
        RECT -143.420 103.750 -142.900 103.770 ;
        RECT -150.440 103.030 -148.000 103.320 ;
        RECT -143.420 103.240 -142.910 103.750 ;
        RECT 11.530 103.580 11.800 104.020 ;
        RECT 13.010 103.760 13.340 104.020 ;
        RECT 14.550 103.880 14.810 104.020 ;
        RECT 15.550 103.880 15.730 104.320 ;
        RECT 16.280 104.110 17.640 104.220 ;
        RECT 16.280 104.050 17.720 104.110 ;
        RECT 17.080 104.040 17.720 104.050 ;
        RECT 11.570 103.570 11.800 103.580 ;
        RECT 14.550 103.710 15.730 103.880 ;
        RECT 17.250 103.940 17.720 104.040 ;
        RECT 18.190 103.960 19.150 104.130 ;
        RECT 14.550 103.570 14.810 103.710 ;
        RECT 17.250 103.690 17.500 103.940 ;
        RECT 11.570 103.400 12.330 103.570 ;
        RECT 12.580 103.400 13.750 103.570 ;
        RECT 13.990 103.540 14.810 103.570 ;
        RECT 16.050 103.540 16.230 103.600 ;
        RECT 13.990 103.400 15.100 103.540 ;
        RECT 12.980 103.300 13.330 103.400 ;
        RECT 14.640 103.370 15.100 103.400 ;
        RECT 15.550 103.370 16.230 103.540 ;
        RECT 17.170 103.520 17.500 103.690 ;
        RECT 18.970 103.500 19.150 103.960 ;
        RECT 30.750 103.920 30.920 104.340 ;
        RECT 31.560 104.210 31.800 104.250 ;
        RECT 34.340 104.210 34.510 104.220 ;
        RECT 34.790 104.210 34.990 104.450 ;
        RECT 31.230 104.040 31.800 104.210 ;
        RECT 32.040 104.040 33.380 104.210 ;
        RECT 33.830 104.040 34.990 104.210 ;
        RECT 31.560 104.010 31.800 104.040 ;
        RECT 15.590 103.350 16.230 103.370 ;
        RECT 16.050 103.340 16.230 103.350 ;
        RECT 17.830 103.340 18.430 103.490 ;
        RECT 16.050 103.320 18.430 103.340 ;
        RECT 18.890 103.330 19.220 103.500 ;
        RECT 34.790 103.440 34.990 104.040 ;
        RECT 35.320 103.970 35.490 104.900 ;
        RECT 35.720 103.920 35.890 104.770 ;
        RECT 40.540 103.440 40.830 104.450 ;
        RECT -143.420 103.030 -142.890 103.240 ;
        RECT 16.050 103.170 18.280 103.320 ;
        RECT -150.440 102.550 -142.890 103.030 ;
        RECT 38.180 102.850 38.380 103.200 ;
        RECT 39.920 103.120 40.240 103.130 ;
        RECT 39.660 102.950 40.240 103.120 ;
        RECT 39.910 102.900 40.240 102.950 ;
        RECT 39.920 102.870 40.240 102.900 ;
        RECT 38.170 102.820 38.380 102.850 ;
        RECT -150.440 102.520 -143.080 102.550 ;
        RECT 38.170 102.230 38.390 102.820 ;
        RECT 38.910 102.260 39.110 102.830 ;
        RECT 39.920 102.540 40.240 102.580 ;
        RECT 39.910 102.500 40.240 102.540 ;
        RECT 39.660 102.330 40.240 102.500 ;
        RECT 39.920 102.320 40.240 102.330 ;
        RECT -150.440 100.760 -142.910 101.310 ;
        RECT 38.170 101.200 38.390 101.790 ;
        RECT 40.920 101.770 41.090 102.280 ;
        RECT 44.860 101.780 45.030 102.290 ;
        RECT 38.170 101.170 38.380 101.200 ;
        RECT 38.910 101.190 39.110 101.760 ;
        RECT 39.920 101.690 40.240 101.700 ;
        RECT 39.660 101.520 40.240 101.690 ;
        RECT 39.910 101.480 40.240 101.520 ;
        RECT 39.920 101.440 40.240 101.480 ;
        RECT 49.660 101.440 49.840 105.350 ;
        RECT 50.470 104.500 50.640 105.780 ;
        RECT 51.060 105.760 51.230 106.330 ;
        RECT 51.300 106.040 51.470 106.080 ;
        RECT 51.890 106.070 52.060 106.400 ;
        RECT 52.260 106.250 52.850 106.550 ;
        RECT 53.670 106.610 54.250 106.780 ;
        RECT 77.970 106.760 78.200 106.780 ;
        RECT 79.320 106.770 79.490 106.930 ;
        RECT 79.780 106.850 80.390 107.020 ;
        RECT 77.970 106.740 78.230 106.760 ;
        RECT 77.970 106.690 78.310 106.740 ;
        RECT 77.970 106.630 78.460 106.690 ;
        RECT 53.670 106.510 54.060 106.610 ;
        RECT 77.970 106.600 78.480 106.630 ;
        RECT 78.010 106.570 78.480 106.600 ;
        RECT 78.140 106.520 78.480 106.570 ;
        RECT 79.780 106.520 79.960 106.850 ;
        RECT 80.180 106.840 80.390 106.850 ;
        RECT 80.200 106.810 80.390 106.840 ;
        RECT 80.590 106.970 81.090 107.160 ;
        RECT 81.330 107.020 81.520 107.050 ;
        RECT 80.590 106.930 81.080 106.970 ;
        RECT 78.260 106.510 78.480 106.520 ;
        RECT 53.670 106.480 54.050 106.510 ;
        RECT 78.270 106.480 78.480 106.510 ;
        RECT 53.670 106.330 54.030 106.480 ;
        RECT 78.290 106.400 78.480 106.480 ;
        RECT 79.650 106.400 79.980 106.520 ;
        RECT 80.590 106.400 80.760 106.930 ;
        RECT 80.820 106.770 80.990 106.930 ;
        RECT 81.330 106.880 81.770 107.020 ;
        RECT 81.830 106.880 82.030 106.920 ;
        RECT 81.330 106.820 82.030 106.880 ;
        RECT 81.420 106.620 82.030 106.820 ;
        RECT 81.420 106.580 81.590 106.620 ;
        RECT 81.830 106.590 82.030 106.620 ;
        RECT 82.050 106.430 82.220 107.110 ;
        RECT 77.800 106.350 77.970 106.370 ;
        RECT 51.710 106.040 52.060 106.070 ;
        RECT 51.300 105.780 52.060 106.040 ;
        RECT 51.300 105.750 51.470 105.780 ;
        RECT 51.710 105.750 52.060 105.780 ;
        RECT 51.710 105.740 51.910 105.750 ;
        RECT 52.300 105.740 52.850 106.250 ;
        RECT 53.320 106.160 54.030 106.330 ;
        RECT 77.780 105.920 77.990 106.350 ;
        RECT 78.290 106.230 78.810 106.400 ;
        RECT 78.290 106.200 78.480 106.230 ;
        RECT 79.160 106.220 81.060 106.400 ;
        RECT 81.790 106.390 82.220 106.430 ;
        RECT 81.440 106.230 82.220 106.390 ;
        RECT 81.440 106.220 82.030 106.230 ;
        RECT 79.780 106.070 79.960 106.220 ;
        RECT 80.590 106.080 80.760 106.220 ;
        RECT 81.600 105.970 82.030 106.220 ;
        RECT 81.830 105.930 82.030 105.970 ;
        RECT 82.420 105.930 82.970 106.920 ;
        RECT 83.440 106.910 84.140 107.220 ;
        RECT 83.440 106.300 84.150 106.470 ;
        RECT 83.790 106.020 84.150 106.300 ;
        RECT 83.790 105.850 84.370 106.020 ;
        RECT 52.610 105.500 52.830 105.740 ;
        RECT 52.620 105.470 52.830 105.500 ;
        RECT 50.810 105.240 51.340 105.370 ;
        RECT 52.620 105.250 52.820 105.470 ;
        RECT 53.320 105.410 54.020 105.720 ;
        RECT 50.810 105.210 51.470 105.240 ;
        RECT 51.710 105.210 51.910 105.250 ;
        RECT 50.810 105.200 51.910 105.210 ;
        RECT 51.300 104.950 51.910 105.200 ;
        RECT 51.300 104.910 51.470 104.950 ;
        RECT 51.710 104.920 51.910 104.950 ;
        RECT 51.710 104.560 51.910 104.590 ;
        RECT 50.270 104.300 50.590 104.330 ;
        RECT 51.480 104.300 51.910 104.560 ;
        RECT 50.270 104.110 50.600 104.300 ;
        RECT 51.710 104.260 51.910 104.300 ;
        RECT 52.300 104.260 52.850 105.250 ;
        RECT 53.170 105.180 54.020 105.410 ;
        RECT 77.780 105.280 77.990 105.710 ;
        RECT 78.290 105.400 78.480 105.430 ;
        RECT 81.790 105.410 81.980 105.430 ;
        RECT 77.800 105.260 77.970 105.280 ;
        RECT 53.320 104.840 54.020 105.180 ;
        RECT 78.290 105.230 78.810 105.400 ;
        RECT 79.160 105.230 81.060 105.410 ;
        RECT 81.440 105.400 81.980 105.410 ;
        RECT 81.440 105.240 82.220 105.400 ;
        RECT 78.290 105.150 78.480 105.230 ;
        RECT 78.270 105.120 78.480 105.150 ;
        RECT 78.260 105.110 78.480 105.120 ;
        RECT 79.650 105.110 79.980 105.230 ;
        RECT 81.790 105.200 82.220 105.240 ;
        RECT 78.140 105.060 78.480 105.110 ;
        RECT 78.010 105.030 78.480 105.060 ;
        RECT 77.970 105.000 78.480 105.030 ;
        RECT 77.970 104.940 78.460 105.000 ;
        RECT 77.970 104.890 78.310 104.940 ;
        RECT 77.970 104.870 78.230 104.890 ;
        RECT 77.970 104.850 78.200 104.870 ;
        RECT 77.970 104.810 78.180 104.850 ;
        RECT 77.970 104.530 78.140 104.810 ;
        RECT 79.320 104.700 79.490 104.860 ;
        RECT 80.200 104.790 80.390 104.820 ;
        RECT 80.180 104.780 80.390 104.790 ;
        RECT 79.190 104.660 79.510 104.700 ;
        RECT 53.780 104.480 54.100 104.520 ;
        RECT 53.780 104.420 54.110 104.480 ;
        RECT 79.190 104.470 79.520 104.660 ;
        RECT 79.930 104.610 80.390 104.780 ;
        RECT 80.820 104.700 80.990 104.860 ;
        RECT 81.330 104.780 81.520 104.810 ;
        RECT 80.200 104.590 80.390 104.610 ;
        RECT 80.760 104.660 81.080 104.700 ;
        RECT 80.760 104.470 81.090 104.660 ;
        RECT 81.330 104.610 81.770 104.780 ;
        RECT 81.330 104.580 81.520 104.610 ;
        RECT 82.050 104.520 82.220 105.200 ;
        RECT 206.500 104.850 207.010 115.210 ;
        RECT 207.180 114.420 213.160 114.650 ;
        RECT 206.500 104.830 207.020 104.850 ;
        RECT 79.190 104.440 79.510 104.470 ;
        RECT 80.760 104.440 81.080 104.470 ;
        RECT 53.310 104.290 54.110 104.420 ;
        RECT 53.310 104.260 54.100 104.290 ;
        RECT 53.310 104.240 54.010 104.260 ;
        RECT 50.270 104.070 50.590 104.110 ;
        RECT 50.270 103.990 50.440 104.070 ;
        RECT 50.220 103.820 50.440 103.990 ;
        RECT 50.220 103.660 50.390 103.820 ;
        RECT 51.710 103.730 51.910 103.770 ;
        RECT 50.750 103.400 50.940 103.520 ;
        RECT 51.480 103.470 51.910 103.730 ;
        RECT 51.710 103.440 51.910 103.470 ;
        RECT 50.390 103.290 50.940 103.400 ;
        RECT 50.390 103.230 50.930 103.290 ;
        RECT 50.470 101.450 50.640 103.230 ;
        RECT 51.300 103.080 51.470 103.120 ;
        RECT 51.710 103.080 51.910 103.110 ;
        RECT 51.300 102.820 51.910 103.080 ;
        RECT 51.300 102.790 51.470 102.820 ;
        RECT 51.710 102.780 51.910 102.820 ;
        RECT 52.300 102.780 52.850 103.770 ;
        RECT 53.770 103.760 54.090 103.800 ;
        RECT 53.310 103.580 54.100 103.760 ;
        RECT 53.770 103.570 54.100 103.580 ;
        RECT 53.770 103.540 54.090 103.570 ;
        RECT 53.320 102.820 54.020 103.160 ;
        RECT 60.720 103.120 61.040 103.130 ;
        RECT 60.720 102.950 61.300 103.120 ;
        RECT 60.720 102.900 61.050 102.950 ;
        RECT 60.720 102.870 61.040 102.900 ;
        RECT 62.580 102.850 62.780 103.200 ;
        RECT 206.490 103.050 207.020 104.830 ;
        RECT 207.420 103.360 213.070 114.420 ;
        RECT 207.360 103.350 213.070 103.360 ;
        RECT 207.360 103.180 213.150 103.350 ;
        RECT 207.360 103.170 213.060 103.180 ;
        RECT 207.420 103.100 207.590 103.170 ;
        RECT 206.490 103.030 207.010 103.050 ;
        RECT 53.170 102.590 54.020 102.820 ;
        RECT 51.300 102.250 51.470 102.280 ;
        RECT 51.710 102.250 51.910 102.290 ;
        RECT 51.300 101.990 51.910 102.250 ;
        RECT 51.300 101.950 51.470 101.990 ;
        RECT 51.710 101.960 51.910 101.990 ;
        RECT 51.710 101.600 51.910 101.630 ;
        RECT 51.480 101.340 51.910 101.600 ;
        RECT 51.710 101.300 51.910 101.340 ;
        RECT 52.300 101.300 52.850 102.290 ;
        RECT 53.320 102.280 54.020 102.590 ;
        RECT 60.720 102.540 61.040 102.580 ;
        RECT 60.720 102.500 61.050 102.540 ;
        RECT 60.720 102.330 61.300 102.500 ;
        RECT 60.720 102.320 61.040 102.330 ;
        RECT 53.320 101.670 54.030 101.840 ;
        RECT 55.930 101.780 56.100 102.290 ;
        RECT 59.870 101.770 60.040 102.280 ;
        RECT 61.850 102.260 62.050 102.830 ;
        RECT 62.580 102.820 62.790 102.850 ;
        RECT 62.570 102.230 62.790 102.820 ;
        RECT 206.500 102.520 207.010 103.030 ;
        RECT 213.520 102.600 214.030 115.210 ;
        RECT 214.270 109.190 215.730 109.230 ;
        RECT 214.260 109.020 215.730 109.190 ;
        RECT 214.270 108.980 215.730 109.020 ;
        RECT 206.480 102.310 207.010 102.520 ;
        RECT 211.590 102.310 214.030 102.600 ;
        RECT 206.480 101.830 214.030 102.310 ;
        RECT 206.670 101.800 214.030 101.830 ;
        RECT 53.670 101.390 54.030 101.670 ;
        RECT 60.720 101.690 61.040 101.700 ;
        RECT 60.720 101.520 61.300 101.690 ;
        RECT 60.720 101.480 61.050 101.520 ;
        RECT 60.720 101.440 61.040 101.480 ;
        RECT 53.670 101.220 54.250 101.390 ;
        RECT 61.850 101.190 62.050 101.760 ;
        RECT 62.570 101.200 62.790 101.790 ;
        RECT 38.180 100.820 38.380 101.170 ;
        RECT 62.580 101.170 62.790 101.200 ;
        RECT 39.920 101.120 40.240 101.150 ;
        RECT 39.910 101.070 40.240 101.120 ;
        RECT 60.720 101.120 61.040 101.150 ;
        RECT 39.660 100.900 40.240 101.070 ;
        RECT 39.920 100.890 40.240 100.900 ;
        RECT -152.120 87.790 -150.650 88.040 ;
        RECT -150.440 87.850 -149.930 100.760 ;
        RECT -143.580 100.750 -142.910 100.760 ;
        RECT -147.280 99.860 -143.820 100.300 ;
        RECT -149.210 99.760 -143.820 99.860 ;
        RECT -149.210 99.690 -143.930 99.760 ;
        RECT -149.210 88.780 -149.040 99.690 ;
        RECT -148.710 99.280 -144.480 99.300 ;
        RECT -148.730 89.170 -144.400 99.280 ;
        RECT -148.670 89.120 -148.500 89.170 ;
        RECT -144.100 88.780 -143.930 99.690 ;
        RECT -149.210 88.610 -143.930 88.780 ;
        RECT -144.170 88.600 -143.930 88.610 ;
        RECT -143.420 87.850 -142.910 100.750 ;
        RECT 38.550 100.420 38.990 100.590 ;
        RECT 38.180 99.840 38.380 100.190 ;
        RECT 39.920 100.110 40.240 100.120 ;
        RECT 39.660 99.940 40.240 100.110 ;
        RECT 39.910 99.890 40.240 99.940 ;
        RECT 40.920 99.930 41.090 100.940 ;
        RECT 42.850 100.210 43.400 100.640 ;
        RECT 44.850 100.070 45.020 101.080 ;
        RECT 46.880 100.280 47.430 100.710 ;
        RECT 53.530 100.280 54.080 100.710 ;
        RECT 55.940 100.070 56.110 101.080 ;
        RECT 60.720 101.070 61.050 101.120 ;
        RECT 57.560 100.210 58.110 100.640 ;
        RECT 59.870 99.930 60.040 100.940 ;
        RECT 60.720 100.900 61.300 101.070 ;
        RECT 60.720 100.890 61.040 100.900 ;
        RECT 62.580 100.820 62.780 101.170 ;
        RECT 61.970 100.420 62.410 100.590 ;
        RECT 60.720 100.110 61.040 100.120 ;
        RECT 60.720 99.940 61.300 100.110 ;
        RECT 39.920 99.860 40.240 99.890 ;
        RECT 60.720 99.890 61.050 99.940 ;
        RECT 60.720 99.860 61.040 99.890 ;
        RECT 38.170 99.810 38.380 99.840 ;
        RECT 62.580 99.840 62.780 100.190 ;
        RECT 206.500 100.040 214.030 100.590 ;
        RECT 206.500 100.030 207.170 100.040 ;
        RECT 10.980 98.900 11.150 98.950 ;
        RECT 30.750 98.920 30.920 99.340 ;
        RECT 31.560 99.220 31.800 99.250 ;
        RECT 31.230 99.050 31.800 99.220 ;
        RECT 32.040 99.050 33.380 99.220 ;
        RECT 33.830 99.050 34.790 99.220 ;
        RECT 31.560 99.010 31.800 99.050 ;
        RECT 34.340 99.040 34.510 99.050 ;
        RECT 10.950 98.680 11.170 98.900 ;
        RECT 10.980 98.620 11.150 98.680 ;
        RECT 11.500 98.540 11.830 98.720 ;
        RECT 14.640 98.710 14.810 98.760 ;
        RECT 12.080 98.540 14.240 98.710 ;
        RECT 14.480 98.540 14.810 98.710 ;
        RECT 15.100 98.570 15.310 98.900 ;
        RECT 11.530 98.100 11.800 98.540 ;
        RECT 13.010 98.280 13.340 98.540 ;
        RECT 14.550 98.400 14.810 98.540 ;
        RECT 15.550 98.400 15.730 98.840 ;
        RECT 16.280 98.630 17.640 98.740 ;
        RECT 30.680 98.700 30.850 98.740 ;
        RECT 16.280 98.570 17.720 98.630 ;
        RECT 17.080 98.560 17.720 98.570 ;
        RECT 11.570 98.090 11.800 98.100 ;
        RECT 14.550 98.230 15.730 98.400 ;
        RECT 17.250 98.460 17.720 98.560 ;
        RECT 18.190 98.480 19.150 98.650 ;
        RECT 30.620 98.530 30.850 98.700 ;
        RECT 14.550 98.090 14.810 98.230 ;
        RECT 17.250 98.210 17.500 98.460 ;
        RECT 11.570 97.920 12.330 98.090 ;
        RECT 12.580 97.920 13.750 98.090 ;
        RECT 13.990 98.060 14.810 98.090 ;
        RECT 16.050 98.060 16.230 98.120 ;
        RECT 13.990 97.920 15.100 98.060 ;
        RECT 12.980 97.820 13.330 97.920 ;
        RECT 14.640 97.890 15.100 97.920 ;
        RECT 15.550 97.890 16.230 98.060 ;
        RECT 17.170 98.040 17.500 98.210 ;
        RECT 18.970 98.020 19.150 98.480 ;
        RECT 30.680 98.180 30.850 98.530 ;
        RECT 31.020 98.600 31.210 98.620 ;
        RECT 34.020 98.600 34.350 98.780 ;
        RECT 31.020 98.430 31.580 98.600 ;
        RECT 32.040 98.430 34.790 98.600 ;
        RECT 31.020 98.390 31.210 98.430 ;
        RECT 35.320 98.360 35.490 99.290 ;
        RECT 35.720 98.490 35.890 99.340 ;
        RECT 38.170 99.220 38.390 99.810 ;
        RECT 38.910 99.250 39.110 99.820 ;
        RECT 39.920 99.530 40.240 99.570 ;
        RECT 39.910 99.490 40.240 99.530 ;
        RECT 39.660 99.320 40.240 99.490 ;
        RECT 39.920 99.310 40.240 99.320 ;
        RECT 60.720 99.530 61.040 99.570 ;
        RECT 60.720 99.490 61.050 99.530 ;
        RECT 60.720 99.320 61.300 99.490 ;
        RECT 60.720 99.310 61.040 99.320 ;
        RECT 61.850 99.250 62.050 99.820 ;
        RECT 62.580 99.810 62.790 99.840 ;
        RECT 62.570 99.220 62.790 99.810 ;
        RECT 38.170 98.200 38.390 98.790 ;
        RECT 38.170 98.170 38.380 98.200 ;
        RECT 38.910 98.190 39.110 98.760 ;
        RECT 39.920 98.690 40.240 98.700 ;
        RECT 39.660 98.520 40.240 98.690 ;
        RECT 39.910 98.480 40.240 98.520 ;
        RECT 39.920 98.440 40.240 98.480 ;
        RECT 60.720 98.690 61.040 98.700 ;
        RECT 60.720 98.520 61.300 98.690 ;
        RECT 60.720 98.480 61.050 98.520 ;
        RECT 60.720 98.440 61.040 98.480 ;
        RECT 61.850 98.190 62.050 98.760 ;
        RECT 62.570 98.200 62.790 98.790 ;
        RECT 15.590 97.870 16.230 97.890 ;
        RECT 16.050 97.860 16.230 97.870 ;
        RECT 17.830 97.860 18.430 98.010 ;
        RECT 16.050 97.840 18.430 97.860 ;
        RECT 18.890 97.850 19.220 98.020 ;
        RECT 16.050 97.690 18.280 97.840 ;
        RECT 30.680 97.590 30.850 97.940 ;
        RECT 38.180 97.820 38.380 98.170 ;
        RECT 62.580 98.170 62.790 98.200 ;
        RECT 39.920 98.120 40.240 98.150 ;
        RECT 39.910 98.070 40.240 98.120 ;
        RECT 39.660 97.900 40.240 98.070 ;
        RECT 39.920 97.890 40.240 97.900 ;
        RECT 60.720 98.120 61.040 98.150 ;
        RECT 60.720 98.070 61.050 98.120 ;
        RECT 60.720 97.900 61.300 98.070 ;
        RECT 60.720 97.890 61.040 97.900 ;
        RECT 62.580 97.820 62.780 98.170 ;
        RECT 30.620 97.420 30.850 97.590 ;
        RECT 31.020 97.690 31.210 97.730 ;
        RECT 31.020 97.520 31.580 97.690 ;
        RECT 32.040 97.520 34.790 97.690 ;
        RECT 31.020 97.500 31.210 97.520 ;
        RECT 10.980 97.350 11.150 97.400 ;
        RECT 30.680 97.380 30.850 97.420 ;
        RECT 10.950 97.130 11.170 97.350 ;
        RECT 10.980 97.070 11.150 97.130 ;
        RECT 11.500 96.990 11.830 97.170 ;
        RECT 14.640 97.160 14.810 97.210 ;
        RECT 12.080 96.990 14.240 97.160 ;
        RECT 14.480 96.990 14.810 97.160 ;
        RECT 15.100 97.020 15.310 97.350 ;
        RECT 34.020 97.340 34.350 97.520 ;
        RECT 11.530 96.550 11.800 96.990 ;
        RECT 13.010 96.730 13.340 96.990 ;
        RECT 14.550 96.850 14.810 96.990 ;
        RECT 15.550 96.850 15.730 97.290 ;
        RECT 16.280 97.080 17.640 97.190 ;
        RECT 16.280 97.020 17.720 97.080 ;
        RECT 17.080 97.010 17.720 97.020 ;
        RECT 11.570 96.540 11.800 96.550 ;
        RECT 14.550 96.680 15.730 96.850 ;
        RECT 17.250 96.910 17.720 97.010 ;
        RECT 18.190 96.930 19.150 97.100 ;
        RECT 14.550 96.540 14.810 96.680 ;
        RECT 17.250 96.660 17.500 96.910 ;
        RECT 11.570 96.370 12.330 96.540 ;
        RECT 12.580 96.370 13.750 96.540 ;
        RECT 13.990 96.510 14.810 96.540 ;
        RECT 16.050 96.510 16.230 96.570 ;
        RECT 13.990 96.370 15.100 96.510 ;
        RECT 12.980 96.270 13.330 96.370 ;
        RECT 14.640 96.340 15.100 96.370 ;
        RECT 15.550 96.340 16.230 96.510 ;
        RECT 17.170 96.490 17.500 96.660 ;
        RECT 18.970 96.470 19.150 96.930 ;
        RECT 30.750 96.780 30.920 97.200 ;
        RECT 31.560 97.070 31.800 97.110 ;
        RECT 34.340 97.070 34.510 97.080 ;
        RECT 31.230 96.900 31.800 97.070 ;
        RECT 32.040 96.900 33.380 97.070 ;
        RECT 33.830 96.900 34.790 97.070 ;
        RECT 31.560 96.870 31.800 96.900 ;
        RECT 35.320 96.830 35.490 97.760 ;
        RECT 35.720 96.780 35.890 97.630 ;
        RECT 15.590 96.320 16.230 96.340 ;
        RECT 16.050 96.310 16.230 96.320 ;
        RECT 17.830 96.310 18.430 96.460 ;
        RECT 16.050 96.290 18.430 96.310 ;
        RECT 18.890 96.300 19.220 96.470 ;
        RECT 16.050 96.140 18.280 96.290 ;
        RECT 30.750 95.990 30.920 96.410 ;
        RECT 31.560 96.290 31.800 96.320 ;
        RECT 31.230 96.120 31.800 96.290 ;
        RECT 32.040 96.120 33.380 96.290 ;
        RECT 33.830 96.120 34.790 96.290 ;
        RECT 31.560 96.080 31.800 96.120 ;
        RECT 34.340 96.110 34.510 96.120 ;
        RECT 10.980 95.800 11.150 95.850 ;
        RECT 10.950 95.580 11.170 95.800 ;
        RECT 10.980 95.520 11.150 95.580 ;
        RECT 11.500 95.440 11.830 95.620 ;
        RECT 14.640 95.610 14.810 95.660 ;
        RECT 12.080 95.440 14.240 95.610 ;
        RECT 14.480 95.440 14.810 95.610 ;
        RECT 15.100 95.470 15.310 95.800 ;
        RECT 30.680 95.770 30.850 95.810 ;
        RECT 11.530 95.000 11.800 95.440 ;
        RECT 13.010 95.180 13.340 95.440 ;
        RECT 14.550 95.300 14.810 95.440 ;
        RECT 15.550 95.300 15.730 95.740 ;
        RECT 16.280 95.530 17.640 95.640 ;
        RECT 30.620 95.600 30.850 95.770 ;
        RECT 16.280 95.470 17.720 95.530 ;
        RECT 17.080 95.460 17.720 95.470 ;
        RECT 11.570 94.990 11.800 95.000 ;
        RECT 14.550 95.130 15.730 95.300 ;
        RECT 17.250 95.360 17.720 95.460 ;
        RECT 18.190 95.380 19.150 95.550 ;
        RECT 14.550 94.990 14.810 95.130 ;
        RECT 17.250 95.110 17.500 95.360 ;
        RECT 11.570 94.820 12.330 94.990 ;
        RECT 12.580 94.820 13.750 94.990 ;
        RECT 13.990 94.960 14.810 94.990 ;
        RECT 16.050 94.960 16.230 95.020 ;
        RECT 13.990 94.820 15.100 94.960 ;
        RECT 12.980 94.720 13.330 94.820 ;
        RECT 14.640 94.790 15.100 94.820 ;
        RECT 15.550 94.790 16.230 94.960 ;
        RECT 17.170 94.940 17.500 95.110 ;
        RECT 18.970 94.920 19.150 95.380 ;
        RECT 30.680 95.250 30.850 95.600 ;
        RECT 31.020 95.670 31.210 95.690 ;
        RECT 34.020 95.670 34.350 95.850 ;
        RECT 31.020 95.500 31.580 95.670 ;
        RECT 32.040 95.500 34.790 95.670 ;
        RECT 31.020 95.460 31.210 95.500 ;
        RECT 35.320 95.430 35.490 96.360 ;
        RECT 35.720 95.560 35.890 96.410 ;
        RECT 15.590 94.770 16.230 94.790 ;
        RECT 16.050 94.760 16.230 94.770 ;
        RECT 17.830 94.760 18.430 94.910 ;
        RECT 16.050 94.740 18.430 94.760 ;
        RECT 18.890 94.750 19.220 94.920 ;
        RECT 16.050 94.590 18.280 94.740 ;
        RECT 30.680 94.660 30.850 95.010 ;
        RECT 30.620 94.490 30.850 94.660 ;
        RECT 31.020 94.760 31.210 94.800 ;
        RECT 31.020 94.590 31.580 94.760 ;
        RECT 32.040 94.590 34.790 94.760 ;
        RECT 31.020 94.570 31.210 94.590 ;
        RECT 30.680 94.450 30.850 94.490 ;
        RECT 34.020 94.410 34.350 94.590 ;
        RECT 10.980 94.250 11.150 94.300 ;
        RECT 10.950 94.030 11.170 94.250 ;
        RECT 10.980 93.970 11.150 94.030 ;
        RECT 11.500 93.890 11.830 94.070 ;
        RECT 14.640 94.060 14.810 94.110 ;
        RECT 12.080 93.890 14.240 94.060 ;
        RECT 14.480 93.890 14.810 94.060 ;
        RECT 15.100 93.920 15.310 94.250 ;
        RECT 11.530 93.450 11.800 93.890 ;
        RECT 13.010 93.630 13.340 93.890 ;
        RECT 14.550 93.750 14.810 93.890 ;
        RECT 15.550 93.750 15.730 94.190 ;
        RECT 16.280 93.980 17.640 94.090 ;
        RECT 16.280 93.920 17.720 93.980 ;
        RECT 17.080 93.910 17.720 93.920 ;
        RECT 11.570 93.440 11.800 93.450 ;
        RECT 14.550 93.580 15.730 93.750 ;
        RECT 17.250 93.810 17.720 93.910 ;
        RECT 18.190 93.830 19.150 94.000 ;
        RECT 30.750 93.850 30.920 94.270 ;
        RECT 31.560 94.140 31.800 94.180 ;
        RECT 34.340 94.140 34.510 94.150 ;
        RECT 31.230 93.970 31.800 94.140 ;
        RECT 32.040 93.970 33.380 94.140 ;
        RECT 33.830 93.970 34.790 94.140 ;
        RECT 31.560 93.940 31.800 93.970 ;
        RECT 35.320 93.900 35.490 94.830 ;
        RECT 35.720 93.850 35.890 94.700 ;
        RECT 14.550 93.440 14.810 93.580 ;
        RECT 17.250 93.560 17.500 93.810 ;
        RECT 11.570 93.270 12.330 93.440 ;
        RECT 12.580 93.270 13.750 93.440 ;
        RECT 13.990 93.410 14.810 93.440 ;
        RECT 16.050 93.410 16.230 93.470 ;
        RECT 13.990 93.270 15.100 93.410 ;
        RECT 12.980 93.170 13.330 93.270 ;
        RECT 14.640 93.240 15.100 93.270 ;
        RECT 15.550 93.240 16.230 93.410 ;
        RECT 17.170 93.390 17.500 93.560 ;
        RECT 18.970 93.370 19.150 93.830 ;
        RECT 15.590 93.220 16.230 93.240 ;
        RECT 16.050 93.210 16.230 93.220 ;
        RECT 17.830 93.210 18.430 93.360 ;
        RECT 16.050 93.190 18.430 93.210 ;
        RECT 18.890 93.200 19.220 93.370 ;
        RECT 16.050 93.040 18.280 93.190 ;
        RECT 25.480 93.030 25.680 93.380 ;
        RECT 27.220 93.300 27.540 93.310 ;
        RECT 26.960 93.130 27.540 93.300 ;
        RECT 27.210 93.080 27.540 93.130 ;
        RECT 27.220 93.050 27.540 93.080 ;
        RECT 25.470 93.000 25.680 93.030 ;
        RECT 25.470 92.410 25.690 93.000 ;
        RECT 26.210 92.440 26.410 93.010 ;
        RECT 27.220 92.720 27.540 92.760 ;
        RECT 27.210 92.680 27.540 92.720 ;
        RECT 26.960 92.510 27.540 92.680 ;
        RECT 27.220 92.500 27.540 92.510 ;
        RECT 25.470 91.380 25.690 91.970 ;
        RECT 25.470 91.350 25.680 91.380 ;
        RECT 26.210 91.370 26.410 91.940 ;
        RECT 28.350 91.930 28.520 92.440 ;
        RECT 32.370 91.960 32.540 92.470 ;
        RECT 27.220 91.870 27.540 91.880 ;
        RECT 26.960 91.700 27.540 91.870 ;
        RECT 27.210 91.660 27.540 91.700 ;
        RECT 27.220 91.620 27.540 91.660 ;
        RECT 25.480 91.000 25.680 91.350 ;
        RECT 27.220 91.300 27.540 91.330 ;
        RECT 27.210 91.250 27.540 91.300 ;
        RECT 26.960 91.080 27.540 91.250 ;
        RECT 27.220 91.070 27.540 91.080 ;
        RECT 25.850 90.600 26.290 90.770 ;
        RECT -12.140 90.110 -11.970 90.600 ;
        RECT -12.290 90.080 -11.970 90.110 ;
        RECT -11.590 90.110 -11.420 90.600 ;
        RECT -10.950 90.550 -10.780 90.600 ;
        RECT -10.400 90.550 -10.230 90.600 ;
        RECT -11.070 90.520 -10.750 90.550 ;
        RECT -10.420 90.520 -10.100 90.550 ;
        RECT -11.070 90.330 -10.740 90.520 ;
        RECT -10.420 90.330 -10.090 90.520 ;
        RECT -11.070 90.290 -10.750 90.330 ;
        RECT -10.420 90.290 -10.100 90.330 ;
        RECT -11.590 90.080 -11.270 90.110 ;
        RECT -12.290 89.890 -11.960 90.080 ;
        RECT -11.590 89.890 -11.260 90.080 ;
        RECT -12.290 89.850 -11.970 89.890 ;
        RECT -12.680 88.390 -12.510 88.410 ;
        RECT -12.700 87.960 -12.490 88.390 ;
        RECT -12.140 88.200 -11.970 89.850 ;
        RECT -11.590 89.850 -11.270 89.890 ;
        RECT -11.590 88.200 -11.420 89.850 ;
        RECT -10.950 88.200 -10.780 90.290 ;
        RECT -10.400 88.200 -10.230 90.290 ;
        RECT 25.480 90.020 25.680 90.370 ;
        RECT 27.220 90.290 27.540 90.300 ;
        RECT 26.960 90.120 27.540 90.290 ;
        RECT 27.210 90.070 27.540 90.120 ;
        RECT 28.340 90.070 28.510 91.260 ;
        RECT 30.150 90.390 30.700 90.820 ;
        RECT 27.220 90.040 27.540 90.070 ;
        RECT 25.470 89.990 25.680 90.020 ;
        RECT 32.360 90.010 32.530 91.200 ;
        RECT 34.180 90.460 34.730 90.890 ;
        RECT -9.850 88.840 -9.680 89.690 ;
        RECT 25.470 89.400 25.690 89.990 ;
        RECT 26.210 89.430 26.410 90.000 ;
        RECT 27.220 89.710 27.540 89.750 ;
        RECT 27.210 89.670 27.540 89.710 ;
        RECT 26.960 89.500 27.540 89.670 ;
        RECT 27.220 89.490 27.540 89.500 ;
        RECT 10.980 89.130 11.150 89.180 ;
        RECT 30.750 89.160 30.920 89.580 ;
        RECT 31.560 89.460 31.800 89.490 ;
        RECT 31.230 89.290 31.800 89.460 ;
        RECT 32.040 89.290 33.380 89.460 ;
        RECT 33.830 89.290 34.790 89.460 ;
        RECT 31.560 89.250 31.800 89.290 ;
        RECT 34.340 89.280 34.510 89.290 ;
        RECT 10.950 88.910 11.170 89.130 ;
        RECT 10.980 88.850 11.150 88.910 ;
        RECT 11.500 88.770 11.830 88.950 ;
        RECT 14.640 88.940 14.810 88.990 ;
        RECT 12.080 88.770 14.240 88.940 ;
        RECT 14.480 88.770 14.810 88.940 ;
        RECT 15.100 88.800 15.310 89.130 ;
        RECT 11.530 88.330 11.800 88.770 ;
        RECT 13.010 88.510 13.340 88.770 ;
        RECT 14.550 88.630 14.810 88.770 ;
        RECT 15.550 88.630 15.730 89.070 ;
        RECT 16.280 88.860 17.640 88.970 ;
        RECT 16.280 88.800 17.720 88.860 ;
        RECT 17.080 88.790 17.720 88.800 ;
        RECT 11.570 88.320 11.800 88.330 ;
        RECT 14.550 88.460 15.730 88.630 ;
        RECT 17.250 88.690 17.720 88.790 ;
        RECT 18.190 88.710 19.150 88.880 ;
        RECT 14.550 88.320 14.810 88.460 ;
        RECT 17.250 88.440 17.500 88.690 ;
        RECT -9.960 88.210 -9.530 88.230 ;
        RECT -9.960 88.040 -9.510 88.210 ;
        RECT 11.570 88.150 12.330 88.320 ;
        RECT 12.580 88.150 13.750 88.320 ;
        RECT 13.990 88.290 14.810 88.320 ;
        RECT 16.050 88.290 16.230 88.350 ;
        RECT 13.990 88.150 15.100 88.290 ;
        RECT 12.980 88.050 13.330 88.150 ;
        RECT 14.640 88.120 15.100 88.150 ;
        RECT 15.550 88.120 16.230 88.290 ;
        RECT 17.170 88.270 17.500 88.440 ;
        RECT 18.970 88.250 19.150 88.710 ;
        RECT 25.470 88.380 25.690 88.970 ;
        RECT 30.680 88.940 30.850 88.980 ;
        RECT 25.470 88.350 25.680 88.380 ;
        RECT 26.210 88.370 26.410 88.940 ;
        RECT 27.220 88.870 27.540 88.880 ;
        RECT 26.960 88.700 27.540 88.870 ;
        RECT 30.620 88.770 30.850 88.940 ;
        RECT 27.210 88.660 27.540 88.700 ;
        RECT 27.220 88.620 27.540 88.660 ;
        RECT 30.680 88.420 30.850 88.770 ;
        RECT 31.020 88.840 31.210 88.860 ;
        RECT 34.020 88.840 34.350 89.020 ;
        RECT 31.020 88.670 31.580 88.840 ;
        RECT 32.040 88.670 34.790 88.840 ;
        RECT 31.020 88.630 31.210 88.670 ;
        RECT 35.320 88.600 35.490 89.530 ;
        RECT 35.720 88.730 35.890 89.580 ;
        RECT 38.590 89.370 38.910 89.400 ;
        RECT 38.590 89.200 40.380 89.370 ;
        RECT 38.590 89.180 38.920 89.200 ;
        RECT 38.590 89.140 38.910 89.180 ;
        RECT 40.210 88.970 40.380 89.200 ;
        RECT 39.060 88.720 39.400 88.970 ;
        RECT 39.570 88.800 39.900 88.970 ;
        RECT 40.120 88.800 40.460 88.970 ;
        RECT 38.740 88.460 39.400 88.720 ;
        RECT 39.650 88.630 39.820 88.800 ;
        RECT 40.210 88.630 40.380 88.800 ;
        RECT 39.570 88.460 39.900 88.630 ;
        RECT 40.120 88.460 40.460 88.630 ;
        RECT 15.590 88.100 16.230 88.120 ;
        RECT 16.050 88.090 16.230 88.100 ;
        RECT 17.830 88.090 18.430 88.240 ;
        RECT 16.050 88.070 18.430 88.090 ;
        RECT 18.890 88.080 19.220 88.250 ;
        RECT -9.960 88.020 -9.530 88.040 ;
        RECT 16.050 87.920 18.280 88.070 ;
        RECT 25.480 88.000 25.680 88.350 ;
        RECT 27.220 88.300 27.540 88.330 ;
        RECT 27.210 88.250 27.540 88.300 ;
        RECT 26.960 88.080 27.540 88.250 ;
        RECT 39.650 88.230 39.900 88.460 ;
        RECT 40.780 88.380 41.290 89.050 ;
        RECT 27.220 88.070 27.540 88.080 ;
        RECT -150.440 87.340 -142.910 87.850 ;
        RECT 30.680 87.830 30.850 88.180 ;
        RECT 39.650 88.060 40.320 88.230 ;
        RECT -152.140 81.320 -150.680 81.360 ;
        RECT -152.140 81.150 -150.670 81.320 ;
        RECT -152.140 81.110 -150.680 81.150 ;
        RECT -150.440 74.730 -149.930 87.340 ;
        RECT -149.570 86.550 -143.590 86.780 ;
        RECT -149.480 75.490 -143.830 86.550 ;
        RECT -143.420 76.980 -142.910 87.340 ;
        RECT -13.600 84.840 -13.430 87.330 ;
        RECT -13.050 84.840 -12.880 87.340 ;
        RECT -12.690 87.320 -12.480 87.750 ;
        RECT -9.950 87.670 -9.520 87.690 ;
        RECT -9.950 87.500 -9.500 87.670 ;
        RECT 30.620 87.660 30.850 87.830 ;
        RECT 31.020 87.930 31.210 87.970 ;
        RECT 31.020 87.760 31.580 87.930 ;
        RECT 32.040 87.760 34.790 87.930 ;
        RECT 31.020 87.740 31.210 87.760 ;
        RECT 10.980 87.580 11.150 87.630 ;
        RECT 30.680 87.620 30.850 87.660 ;
        RECT 34.020 87.580 34.350 87.760 ;
        RECT -9.950 87.480 -9.520 87.500 ;
        RECT 10.950 87.360 11.170 87.580 ;
        RECT -12.670 87.300 -12.500 87.320 ;
        RECT -12.420 86.230 -12.250 87.330 ;
        RECT -12.420 86.200 -11.940 86.230 ;
        RECT -12.420 86.010 -11.930 86.200 ;
        RECT -12.420 85.970 -11.940 86.010 ;
        RECT -12.420 84.840 -12.250 85.970 ;
        RECT -11.870 84.840 -11.700 87.340 ;
        RECT 10.980 87.300 11.150 87.360 ;
        RECT 11.500 87.220 11.830 87.400 ;
        RECT 14.640 87.390 14.810 87.440 ;
        RECT 12.080 87.220 14.240 87.390 ;
        RECT 14.480 87.220 14.810 87.390 ;
        RECT 15.100 87.250 15.310 87.580 ;
        RECT -9.860 86.290 -9.690 86.960 ;
        RECT 11.530 86.780 11.800 87.220 ;
        RECT 13.010 86.960 13.340 87.220 ;
        RECT 14.550 87.080 14.810 87.220 ;
        RECT 15.550 87.080 15.730 87.520 ;
        RECT 16.280 87.310 17.640 87.420 ;
        RECT 16.280 87.250 17.720 87.310 ;
        RECT 17.080 87.240 17.720 87.250 ;
        RECT 11.570 86.770 11.800 86.780 ;
        RECT 14.550 86.910 15.730 87.080 ;
        RECT 17.250 87.140 17.720 87.240 ;
        RECT 18.190 87.160 19.150 87.330 ;
        RECT 14.550 86.770 14.810 86.910 ;
        RECT 17.250 86.890 17.500 87.140 ;
        RECT 11.570 86.600 12.330 86.770 ;
        RECT 12.580 86.600 13.750 86.770 ;
        RECT 13.990 86.740 14.810 86.770 ;
        RECT 16.050 86.740 16.230 86.800 ;
        RECT 13.990 86.600 15.100 86.740 ;
        RECT 12.980 86.500 13.330 86.600 ;
        RECT 14.640 86.570 15.100 86.600 ;
        RECT 15.550 86.570 16.230 86.740 ;
        RECT 17.170 86.720 17.500 86.890 ;
        RECT 18.970 86.700 19.150 87.160 ;
        RECT 30.750 87.020 30.920 87.440 ;
        RECT 31.560 87.310 31.800 87.350 ;
        RECT 34.340 87.310 34.510 87.320 ;
        RECT 31.230 87.140 31.800 87.310 ;
        RECT 32.040 87.140 33.380 87.310 ;
        RECT 33.830 87.140 34.790 87.310 ;
        RECT 31.560 87.110 31.800 87.140 ;
        RECT 35.320 87.070 35.490 88.000 ;
        RECT 35.720 87.020 35.890 87.870 ;
        RECT 39.650 87.830 39.900 88.060 ;
        RECT 38.740 87.570 39.400 87.830 ;
        RECT 39.570 87.660 39.900 87.830 ;
        RECT 40.120 87.660 40.460 87.830 ;
        RECT 39.060 87.320 39.400 87.570 ;
        RECT 39.650 87.490 39.820 87.660 ;
        RECT 40.210 87.490 40.380 87.660 ;
        RECT 39.570 87.320 39.900 87.490 ;
        RECT 40.120 87.320 40.460 87.490 ;
        RECT 38.590 87.110 38.910 87.150 ;
        RECT 38.590 87.090 38.920 87.110 ;
        RECT 40.210 87.090 40.380 87.320 ;
        RECT 40.780 87.240 41.290 87.910 ;
        RECT 38.590 86.920 40.380 87.090 ;
        RECT 206.500 87.130 207.010 100.030 ;
        RECT 207.410 99.140 210.870 99.580 ;
        RECT 207.410 99.040 212.800 99.140 ;
        RECT 207.520 98.970 212.800 99.040 ;
        RECT 207.520 88.060 207.690 98.970 ;
        RECT 208.070 98.560 212.300 98.580 ;
        RECT 207.990 88.450 212.320 98.560 ;
        RECT 212.090 88.400 212.260 88.450 ;
        RECT 212.630 88.060 212.800 98.970 ;
        RECT 207.520 87.890 212.800 88.060 ;
        RECT 207.520 87.880 207.760 87.890 ;
        RECT 213.520 87.130 214.030 100.040 ;
        RECT 38.590 86.890 38.910 86.920 ;
        RECT 15.590 86.550 16.230 86.570 ;
        RECT 16.050 86.540 16.230 86.550 ;
        RECT 17.830 86.540 18.430 86.690 ;
        RECT 16.050 86.520 18.430 86.540 ;
        RECT 18.890 86.530 19.220 86.700 ;
        RECT 16.050 86.370 18.280 86.520 ;
        RECT 30.750 86.230 30.920 86.650 ;
        RECT 31.560 86.530 31.800 86.560 ;
        RECT 31.230 86.360 31.800 86.530 ;
        RECT 32.040 86.360 33.380 86.530 ;
        RECT 33.830 86.360 34.790 86.530 ;
        RECT 31.560 86.320 31.800 86.360 ;
        RECT 34.340 86.350 34.510 86.360 ;
        RECT -11.570 86.190 -11.250 86.220 ;
        RECT -11.570 86.000 -11.240 86.190 ;
        RECT 10.980 86.030 11.150 86.080 ;
        RECT -11.570 85.960 -11.250 86.000 ;
        RECT 10.950 85.810 11.170 86.030 ;
        RECT 10.980 85.750 11.150 85.810 ;
        RECT 11.500 85.670 11.830 85.850 ;
        RECT 14.640 85.840 14.810 85.890 ;
        RECT 12.080 85.670 14.240 85.840 ;
        RECT 14.480 85.670 14.810 85.840 ;
        RECT 15.100 85.700 15.310 86.030 ;
        RECT 30.680 86.010 30.850 86.050 ;
        RECT -11.090 85.420 -10.770 85.450 ;
        RECT -11.090 85.230 -10.760 85.420 ;
        RECT -10.380 85.360 -10.060 85.390 ;
        RECT -11.090 85.190 -10.770 85.230 ;
        RECT -10.380 85.170 -10.050 85.360 ;
        RECT 11.530 85.230 11.800 85.670 ;
        RECT 13.010 85.410 13.340 85.670 ;
        RECT 14.550 85.530 14.810 85.670 ;
        RECT 15.550 85.530 15.730 85.970 ;
        RECT 16.280 85.760 17.640 85.870 ;
        RECT 30.620 85.840 30.850 86.010 ;
        RECT 16.280 85.700 17.720 85.760 ;
        RECT 17.080 85.690 17.720 85.700 ;
        RECT 11.570 85.220 11.800 85.230 ;
        RECT 14.550 85.360 15.730 85.530 ;
        RECT 17.250 85.590 17.720 85.690 ;
        RECT 18.190 85.610 19.150 85.780 ;
        RECT 14.550 85.220 14.810 85.360 ;
        RECT 17.250 85.340 17.500 85.590 ;
        RECT -10.380 85.130 -10.060 85.170 ;
        RECT 11.570 85.050 12.330 85.220 ;
        RECT 12.580 85.050 13.750 85.220 ;
        RECT 13.990 85.190 14.810 85.220 ;
        RECT 16.050 85.190 16.230 85.250 ;
        RECT 13.990 85.050 15.100 85.190 ;
        RECT 12.980 84.950 13.330 85.050 ;
        RECT 14.640 85.020 15.100 85.050 ;
        RECT 15.550 85.020 16.230 85.190 ;
        RECT 17.170 85.170 17.500 85.340 ;
        RECT 18.970 85.150 19.150 85.610 ;
        RECT 30.680 85.490 30.850 85.840 ;
        RECT 31.020 85.910 31.210 85.930 ;
        RECT 34.020 85.910 34.350 86.090 ;
        RECT 31.020 85.740 31.580 85.910 ;
        RECT 32.040 85.740 34.790 85.910 ;
        RECT 31.020 85.700 31.210 85.740 ;
        RECT 35.320 85.670 35.490 86.600 ;
        RECT 35.720 85.800 35.890 86.650 ;
        RECT 38.590 86.600 38.910 86.630 ;
        RECT 206.500 86.620 214.030 87.130 ;
        RECT 214.240 87.070 215.710 87.320 ;
        RECT 38.590 86.430 40.380 86.600 ;
        RECT 38.590 86.410 38.920 86.430 ;
        RECT 38.590 86.370 38.910 86.410 ;
        RECT 40.210 86.200 40.380 86.430 ;
        RECT 39.060 85.950 39.400 86.200 ;
        RECT 39.570 86.030 39.900 86.200 ;
        RECT 40.120 86.030 40.460 86.200 ;
        RECT 38.740 85.690 39.400 85.950 ;
        RECT 39.650 85.860 39.820 86.030 ;
        RECT 40.210 85.860 40.380 86.030 ;
        RECT 39.570 85.690 39.900 85.860 ;
        RECT 40.120 85.690 40.460 85.860 ;
        RECT 39.650 85.460 39.900 85.690 ;
        RECT 40.780 85.610 41.290 86.280 ;
        RECT 39.650 85.290 40.320 85.460 ;
        RECT 15.590 85.000 16.230 85.020 ;
        RECT 16.050 84.990 16.230 85.000 ;
        RECT 17.830 84.990 18.430 85.140 ;
        RECT 16.050 84.970 18.430 84.990 ;
        RECT 18.890 84.980 19.220 85.150 ;
        RECT 16.050 84.820 18.280 84.970 ;
        RECT 27.150 84.960 27.470 85.000 ;
        RECT 27.150 84.770 27.480 84.960 ;
        RECT 30.680 84.900 30.850 85.250 ;
        RECT 27.150 84.740 27.470 84.770 ;
        RECT -13.690 84.130 -13.520 84.200 ;
        RECT -13.760 84.100 -13.440 84.130 ;
        RECT -13.770 83.910 -13.440 84.100 ;
        RECT -13.760 83.870 -13.440 83.910 ;
        RECT -13.690 81.360 -13.520 83.870 ;
        RECT -13.140 83.460 -12.970 84.200 ;
        RECT -12.590 84.140 -12.420 84.200 ;
        RECT -12.660 84.110 -12.340 84.140 ;
        RECT -12.670 83.920 -12.340 84.110 ;
        RECT -12.660 83.880 -12.340 83.920 ;
        RECT -13.210 83.430 -12.890 83.460 ;
        RECT -13.220 83.240 -12.890 83.430 ;
        RECT -13.210 83.200 -12.890 83.240 ;
        RECT -13.140 82.090 -12.970 83.200 ;
        RECT -13.210 82.060 -12.890 82.090 ;
        RECT -13.220 81.870 -12.890 82.060 ;
        RECT -13.210 81.830 -12.890 81.870 ;
        RECT -13.760 81.330 -13.440 81.360 ;
        RECT -13.770 81.140 -13.440 81.330 ;
        RECT -13.760 81.100 -13.440 81.140 ;
        RECT -13.690 80.020 -13.520 81.100 ;
        RECT -13.770 79.990 -13.450 80.020 ;
        RECT -13.780 79.800 -13.450 79.990 ;
        RECT -13.770 79.760 -13.450 79.800 ;
        RECT -13.690 79.020 -13.520 79.760 ;
        RECT -13.140 79.320 -12.970 81.830 ;
        RECT -12.590 81.360 -12.420 83.880 ;
        RECT -12.040 83.460 -11.870 84.200 ;
        RECT -11.490 84.140 -11.320 84.200 ;
        RECT -11.570 84.110 -11.250 84.140 ;
        RECT -11.580 83.920 -11.250 84.110 ;
        RECT -11.570 83.880 -11.250 83.920 ;
        RECT -12.110 83.430 -11.790 83.460 ;
        RECT -12.120 83.240 -11.790 83.430 ;
        RECT -12.110 83.200 -11.790 83.240 ;
        RECT -12.040 82.090 -11.870 83.200 ;
        RECT -12.110 82.060 -11.790 82.090 ;
        RECT -12.120 81.870 -11.790 82.060 ;
        RECT -12.110 81.830 -11.790 81.870 ;
        RECT -12.660 81.330 -12.340 81.360 ;
        RECT -12.670 81.140 -12.340 81.330 ;
        RECT -12.660 81.100 -12.340 81.140 ;
        RECT -12.590 80.010 -12.420 81.100 ;
        RECT -12.660 79.980 -12.340 80.010 ;
        RECT -12.670 79.790 -12.340 79.980 ;
        RECT -12.660 79.750 -12.340 79.790 ;
        RECT -13.210 79.290 -12.890 79.320 ;
        RECT -13.220 79.100 -12.890 79.290 ;
        RECT -13.210 79.060 -12.890 79.100 ;
        RECT -13.140 79.020 -12.970 79.060 ;
        RECT -12.590 79.020 -12.420 79.750 ;
        RECT -12.040 79.310 -11.870 81.830 ;
        RECT -11.490 81.360 -11.320 83.880 ;
        RECT -10.940 83.460 -10.770 84.200 ;
        RECT -10.530 83.920 -10.020 84.600 ;
        RECT 10.980 84.480 11.150 84.530 ;
        RECT 10.950 84.260 11.170 84.480 ;
        RECT 10.980 84.200 11.150 84.260 ;
        RECT 11.500 84.120 11.830 84.300 ;
        RECT 14.640 84.290 14.810 84.340 ;
        RECT 12.080 84.120 14.240 84.290 ;
        RECT 14.480 84.120 14.810 84.290 ;
        RECT 15.100 84.150 15.310 84.480 ;
        RECT -10.530 83.850 -10.010 83.920 ;
        RECT -10.520 83.590 -10.010 83.850 ;
        RECT 11.530 83.680 11.800 84.120 ;
        RECT 13.010 83.860 13.340 84.120 ;
        RECT 14.550 83.980 14.810 84.120 ;
        RECT 15.550 83.980 15.730 84.420 ;
        RECT 16.280 84.210 17.640 84.320 ;
        RECT 16.280 84.150 17.720 84.210 ;
        RECT 17.080 84.140 17.720 84.150 ;
        RECT 11.570 83.670 11.800 83.680 ;
        RECT 14.550 83.810 15.730 83.980 ;
        RECT 17.250 84.040 17.720 84.140 ;
        RECT 18.190 84.060 19.150 84.230 ;
        RECT 14.550 83.670 14.810 83.810 ;
        RECT 17.250 83.790 17.500 84.040 ;
        RECT 11.570 83.500 12.330 83.670 ;
        RECT 12.580 83.500 13.750 83.670 ;
        RECT 13.990 83.640 14.810 83.670 ;
        RECT 16.050 83.640 16.230 83.700 ;
        RECT 13.990 83.500 15.100 83.640 ;
        RECT -11.010 83.430 -10.690 83.460 ;
        RECT -11.020 83.240 -10.690 83.430 ;
        RECT 12.980 83.400 13.330 83.500 ;
        RECT 14.640 83.470 15.100 83.500 ;
        RECT 15.550 83.470 16.230 83.640 ;
        RECT 17.170 83.620 17.500 83.790 ;
        RECT 18.970 83.600 19.150 84.060 ;
        RECT 27.200 84.150 27.380 84.740 ;
        RECT 30.620 84.730 30.850 84.900 ;
        RECT 31.020 85.000 31.210 85.040 ;
        RECT 31.020 84.830 31.580 85.000 ;
        RECT 32.040 84.830 34.790 85.000 ;
        RECT 31.020 84.810 31.210 84.830 ;
        RECT 30.680 84.690 30.850 84.730 ;
        RECT 34.020 84.650 34.350 84.830 ;
        RECT 27.200 84.110 27.520 84.150 ;
        RECT 27.200 83.920 27.530 84.110 ;
        RECT 30.750 84.090 30.920 84.510 ;
        RECT 31.560 84.380 31.800 84.420 ;
        RECT 34.340 84.380 34.510 84.390 ;
        RECT 31.230 84.210 31.800 84.380 ;
        RECT 32.040 84.210 33.380 84.380 ;
        RECT 33.830 84.210 34.790 84.380 ;
        RECT 31.560 84.180 31.800 84.210 ;
        RECT 35.320 84.140 35.490 85.070 ;
        RECT 39.650 85.060 39.900 85.290 ;
        RECT 35.720 84.090 35.890 84.940 ;
        RECT 38.740 84.800 39.400 85.060 ;
        RECT 39.570 84.890 39.900 85.060 ;
        RECT 40.120 84.890 40.460 85.060 ;
        RECT 39.060 84.550 39.400 84.800 ;
        RECT 39.650 84.720 39.820 84.890 ;
        RECT 40.210 84.720 40.380 84.890 ;
        RECT 39.570 84.550 39.900 84.720 ;
        RECT 40.120 84.550 40.460 84.720 ;
        RECT 38.590 84.340 38.910 84.380 ;
        RECT 38.590 84.320 38.920 84.340 ;
        RECT 40.210 84.320 40.380 84.550 ;
        RECT 40.780 84.470 41.290 85.140 ;
        RECT 38.590 84.150 40.380 84.320 ;
        RECT 38.590 84.120 38.910 84.150 ;
        RECT 27.200 83.890 27.520 83.920 ;
        RECT 15.590 83.450 16.230 83.470 ;
        RECT 16.050 83.440 16.230 83.450 ;
        RECT 17.830 83.440 18.430 83.590 ;
        RECT 16.050 83.420 18.430 83.440 ;
        RECT 18.890 83.430 19.220 83.600 ;
        RECT -11.010 83.200 -10.690 83.240 ;
        RECT -10.940 82.090 -10.770 83.200 ;
        RECT -10.230 82.210 -10.060 83.400 ;
        RECT 16.050 83.270 18.280 83.420 ;
        RECT -11.010 82.060 -10.690 82.090 ;
        RECT -11.020 81.870 -10.690 82.060 ;
        RECT -11.010 81.830 -10.690 81.870 ;
        RECT -11.570 81.330 -11.250 81.360 ;
        RECT -11.580 81.140 -11.250 81.330 ;
        RECT -11.570 81.100 -11.250 81.140 ;
        RECT -11.490 79.990 -11.320 81.100 ;
        RECT -11.570 79.960 -11.250 79.990 ;
        RECT -11.580 79.770 -11.250 79.960 ;
        RECT -11.570 79.730 -11.250 79.770 ;
        RECT -12.110 79.280 -11.790 79.310 ;
        RECT -12.120 79.090 -11.790 79.280 ;
        RECT -12.110 79.050 -11.790 79.090 ;
        RECT -12.040 79.020 -11.870 79.050 ;
        RECT -11.490 79.020 -11.320 79.730 ;
        RECT -10.940 79.310 -10.770 81.830 ;
        RECT -3.900 79.900 -3.140 80.320 ;
        RECT -11.020 79.280 -10.700 79.310 ;
        RECT -11.030 79.090 -10.700 79.280 ;
        RECT -3.880 79.110 -3.140 79.900 ;
        RECT -11.020 79.050 -10.700 79.090 ;
        RECT -10.940 79.020 -10.770 79.050 ;
        RECT 27.640 78.170 27.810 78.200 ;
        RECT 28.190 78.170 28.360 78.200 ;
        RECT 28.740 78.170 28.910 78.200 ;
        RECT 29.290 78.170 29.460 78.200 ;
        RECT -143.430 76.960 -142.910 76.980 ;
        RECT -149.480 75.480 -143.770 75.490 ;
        RECT -149.560 75.310 -143.770 75.480 ;
        RECT -149.470 75.300 -143.770 75.310 ;
        RECT -144.000 75.230 -143.830 75.300 ;
        RECT -143.430 75.180 -142.900 76.960 ;
        RECT -13.720 76.540 -13.400 76.570 ;
        RECT -12.620 76.550 -12.300 76.580 ;
        RECT -11.530 76.550 -11.210 76.580 ;
        RECT -13.730 76.350 -13.400 76.540 ;
        RECT -12.630 76.360 -12.300 76.550 ;
        RECT -11.540 76.510 -11.210 76.550 ;
        RECT -10.490 76.510 -9.980 77.040 ;
        RECT -13.720 76.310 -13.400 76.350 ;
        RECT -12.620 76.320 -12.300 76.360 ;
        RECT -12.190 75.900 -12.020 76.510 ;
        RECT -11.640 76.320 -11.210 76.510 ;
        RECT -13.170 75.870 -12.850 75.900 ;
        RECT -13.180 75.680 -12.850 75.870 ;
        RECT -13.170 75.640 -12.850 75.680 ;
        RECT -12.190 75.640 -11.750 75.900 ;
        RECT -143.420 75.160 -142.900 75.180 ;
        RECT -150.440 74.440 -148.000 74.730 ;
        RECT -143.420 74.650 -142.910 75.160 ;
        RECT -143.420 74.440 -142.890 74.650 ;
        RECT -12.190 74.530 -12.020 75.640 ;
        RECT -13.170 74.500 -12.850 74.530 ;
        RECT -150.440 73.960 -142.890 74.440 ;
        RECT -13.180 74.310 -12.850 74.500 ;
        RECT -13.170 74.270 -12.850 74.310 ;
        RECT -12.190 74.270 -11.750 74.530 ;
        RECT -13.650 74.230 -13.490 74.240 ;
        RECT -13.100 74.230 -12.940 74.240 ;
        RECT -12.550 74.230 -12.390 74.240 ;
        RECT -150.440 73.930 -143.080 73.960 ;
        RECT -13.660 73.880 -13.490 74.230 ;
        RECT -13.110 73.900 -12.940 74.230 ;
        RECT -12.560 73.900 -12.390 74.230 ;
        RECT -12.190 74.010 -12.020 74.270 ;
        RECT -12.000 74.230 -11.840 74.240 ;
        RECT -13.650 73.860 -13.490 73.880 ;
        RECT -13.100 73.860 -12.940 73.900 ;
        RECT -12.550 73.860 -12.390 73.900 ;
        RECT -12.010 73.830 -11.840 74.230 ;
        RECT -11.640 74.010 -11.470 76.320 ;
        RECT -11.090 75.900 -10.920 76.510 ;
        RECT -10.540 76.030 -9.820 76.510 ;
        RECT -11.090 75.640 -10.650 75.900 ;
        RECT -11.090 74.530 -10.920 75.640 ;
        RECT -11.090 74.270 -10.650 74.530 ;
        RECT -11.450 74.230 -11.290 74.240 ;
        RECT -11.460 73.900 -11.290 74.230 ;
        RECT -11.090 74.010 -10.920 74.270 ;
        RECT -10.900 74.230 -10.740 74.240 ;
        RECT -11.450 73.860 -11.290 73.900 ;
        RECT -10.910 73.890 -10.740 74.230 ;
        RECT -10.540 74.010 -10.370 76.030 ;
        RECT -9.990 74.010 -9.820 76.030 ;
        RECT -9.440 74.010 -9.270 76.500 ;
        RECT 17.830 75.680 18.000 78.170 ;
        RECT 18.380 75.670 18.550 78.170 ;
        RECT 18.930 75.670 19.100 78.170 ;
        RECT 19.480 77.860 19.650 78.170 ;
        RECT 19.220 77.600 19.650 77.860 ;
        RECT 19.480 75.670 19.650 77.600 ;
        RECT 20.030 77.180 20.200 78.170 ;
        RECT 20.580 77.860 20.750 78.170 ;
        RECT 20.310 77.600 20.750 77.860 ;
        RECT 19.770 76.920 20.200 77.180 ;
        RECT 20.030 75.810 20.200 76.920 ;
        RECT 19.770 75.670 20.200 75.810 ;
        RECT 20.580 75.670 20.750 77.600 ;
        RECT 21.410 77.810 21.730 77.850 ;
        RECT 21.410 77.620 21.740 77.810 ;
        RECT 21.410 77.590 21.730 77.620 ;
        RECT 22.590 77.220 22.760 77.980 ;
        RECT 24.480 77.220 24.650 77.980 ;
        RECT 26.490 77.860 26.660 78.170 ;
        RECT 25.510 77.810 25.830 77.850 ;
        RECT 25.500 77.620 25.830 77.810 ;
        RECT 25.510 77.590 25.830 77.620 ;
        RECT 26.490 77.600 26.930 77.860 ;
        RECT 20.860 77.120 21.180 77.160 ;
        RECT 20.860 76.930 21.190 77.120 ;
        RECT 21.970 77.110 22.290 77.150 ;
        RECT 24.950 77.110 25.270 77.150 ;
        RECT 26.060 77.120 26.380 77.160 ;
        RECT 20.860 76.900 21.180 76.930 ;
        RECT 21.970 76.920 22.300 77.110 ;
        RECT 24.940 76.920 25.270 77.110 ;
        RECT 26.050 76.930 26.380 77.120 ;
        RECT 21.970 76.890 22.290 76.920 ;
        RECT 24.950 76.890 25.270 76.920 ;
        RECT 26.060 76.900 26.380 76.930 ;
        RECT 20.860 75.770 21.180 75.810 ;
        RECT 21.960 75.770 22.280 75.810 ;
        RECT 24.960 75.770 25.280 75.810 ;
        RECT 26.060 75.770 26.380 75.810 ;
        RECT 19.770 75.580 20.100 75.670 ;
        RECT 20.860 75.580 21.190 75.770 ;
        RECT 21.960 75.580 22.290 75.770 ;
        RECT 24.950 75.580 25.280 75.770 ;
        RECT 26.050 75.580 26.380 75.770 ;
        RECT 26.490 75.670 26.660 77.600 ;
        RECT 27.040 77.180 27.210 78.170 ;
        RECT 27.590 77.860 27.810 78.170 ;
        RECT 27.590 77.600 28.020 77.860 ;
        RECT 27.040 76.920 27.470 77.180 ;
        RECT 27.040 75.810 27.210 76.920 ;
        RECT 27.040 75.670 27.470 75.810 ;
        RECT 27.590 75.710 27.810 77.600 ;
        RECT 27.590 75.670 27.760 75.710 ;
        RECT 28.140 75.700 28.360 78.170 ;
        RECT 28.690 75.700 28.910 78.170 ;
        RECT 29.240 77.890 29.460 78.170 ;
        RECT 29.030 77.630 29.460 77.890 ;
        RECT 29.240 75.700 29.460 77.630 ;
        RECT 29.840 77.210 30.010 78.200 ;
        RECT 30.390 77.890 30.560 78.200 ;
        RECT 30.120 77.630 30.560 77.890 ;
        RECT 29.580 76.950 30.010 77.210 ;
        RECT 29.840 75.840 30.010 76.950 ;
        RECT 29.580 75.700 30.010 75.840 ;
        RECT 30.390 75.700 30.560 77.630 ;
        RECT 31.220 77.840 31.540 77.880 ;
        RECT 31.220 77.650 31.550 77.840 ;
        RECT 31.220 77.620 31.540 77.650 ;
        RECT 32.400 77.250 32.570 78.010 ;
        RECT 34.290 77.250 34.460 78.010 ;
        RECT 36.300 77.890 36.470 78.200 ;
        RECT 35.320 77.840 35.640 77.880 ;
        RECT 35.310 77.650 35.640 77.840 ;
        RECT 35.320 77.620 35.640 77.650 ;
        RECT 36.300 77.630 36.740 77.890 ;
        RECT 30.670 77.150 30.990 77.190 ;
        RECT 30.670 76.960 31.000 77.150 ;
        RECT 31.780 77.140 32.100 77.180 ;
        RECT 34.760 77.140 35.080 77.180 ;
        RECT 35.870 77.150 36.190 77.190 ;
        RECT 30.670 76.930 30.990 76.960 ;
        RECT 31.780 76.950 32.110 77.140 ;
        RECT 34.750 76.950 35.080 77.140 ;
        RECT 35.860 76.960 36.190 77.150 ;
        RECT 31.780 76.920 32.100 76.950 ;
        RECT 34.760 76.920 35.080 76.950 ;
        RECT 35.870 76.930 36.190 76.960 ;
        RECT 30.670 75.800 30.990 75.840 ;
        RECT 31.770 75.800 32.090 75.840 ;
        RECT 34.770 75.800 35.090 75.840 ;
        RECT 35.870 75.800 36.190 75.840 ;
        RECT 28.140 75.670 28.310 75.700 ;
        RECT 28.690 75.670 28.860 75.700 ;
        RECT 29.240 75.680 29.410 75.700 ;
        RECT 27.140 75.580 27.470 75.670 ;
        RECT 29.580 75.610 29.910 75.700 ;
        RECT 30.670 75.610 31.000 75.800 ;
        RECT 31.770 75.610 32.100 75.800 ;
        RECT 34.760 75.610 35.090 75.800 ;
        RECT 35.860 75.610 36.190 75.800 ;
        RECT 36.300 75.700 36.470 77.630 ;
        RECT 36.850 77.210 37.020 78.200 ;
        RECT 37.400 77.890 37.570 78.200 ;
        RECT 37.400 77.630 37.830 77.890 ;
        RECT 36.850 76.950 37.280 77.210 ;
        RECT 36.850 75.840 37.020 76.950 ;
        RECT 36.850 75.700 37.280 75.840 ;
        RECT 37.400 75.700 37.570 77.630 ;
        RECT 37.950 75.700 38.120 78.200 ;
        RECT 38.500 75.700 38.670 78.200 ;
        RECT 39.050 75.710 39.220 78.200 ;
        RECT 40.580 77.160 40.750 77.900 ;
        RECT 41.130 77.860 41.300 77.900 ;
        RECT 41.060 77.820 41.380 77.860 ;
        RECT 41.050 77.630 41.380 77.820 ;
        RECT 41.060 77.600 41.380 77.630 ;
        RECT 40.500 77.120 40.820 77.160 ;
        RECT 40.490 76.930 40.820 77.120 ;
        RECT 40.500 76.900 40.820 76.930 ;
        RECT 40.580 75.820 40.750 76.900 ;
        RECT 40.510 75.780 40.830 75.820 ;
        RECT 36.950 75.610 37.280 75.700 ;
        RECT 29.580 75.580 29.900 75.610 ;
        RECT 30.670 75.580 30.990 75.610 ;
        RECT 31.770 75.580 32.090 75.610 ;
        RECT 34.770 75.580 35.090 75.610 ;
        RECT 35.870 75.580 36.190 75.610 ;
        RECT 36.960 75.580 37.280 75.610 ;
        RECT 40.500 75.590 40.830 75.780 ;
        RECT 19.770 75.550 20.090 75.580 ;
        RECT 20.860 75.550 21.180 75.580 ;
        RECT 21.960 75.550 22.280 75.580 ;
        RECT 24.960 75.550 25.280 75.580 ;
        RECT 26.060 75.550 26.380 75.580 ;
        RECT 27.150 75.550 27.470 75.580 ;
        RECT 40.510 75.560 40.830 75.590 ;
        RECT 19.300 75.460 19.460 75.490 ;
        RECT -10.900 73.860 -10.740 73.890 ;
        RECT -13.720 73.770 -13.400 73.800 ;
        RECT -12.620 73.770 -12.300 73.800 ;
        RECT -11.530 73.770 -11.210 73.800 ;
        RECT -13.730 73.580 -13.400 73.770 ;
        RECT -12.630 73.580 -12.300 73.770 ;
        RECT -11.540 73.680 -11.210 73.770 ;
        RECT -13.720 73.540 -13.400 73.580 ;
        RECT -12.620 73.540 -12.300 73.580 ;
        RECT -150.440 72.170 -142.910 72.720 ;
        RECT -13.730 72.430 -13.410 72.460 ;
        RECT -13.740 72.240 -13.410 72.430 ;
        RECT -12.620 72.420 -12.300 72.450 ;
        RECT -13.730 72.200 -13.410 72.240 ;
        RECT -12.630 72.230 -12.300 72.420 ;
        RECT -12.620 72.190 -12.300 72.230 ;
        RECT -152.120 59.200 -150.650 59.450 ;
        RECT -150.440 59.260 -149.930 72.170 ;
        RECT -143.580 72.160 -142.910 72.170 ;
        RECT -147.280 71.270 -143.820 71.710 ;
        RECT -149.210 71.170 -143.820 71.270 ;
        RECT -149.210 71.100 -143.930 71.170 ;
        RECT -149.210 60.190 -149.040 71.100 ;
        RECT -148.710 70.690 -144.480 70.710 ;
        RECT -148.730 60.580 -144.400 70.690 ;
        RECT -148.670 60.530 -148.500 60.580 ;
        RECT -144.100 60.190 -143.930 71.100 ;
        RECT -149.210 60.020 -143.930 60.190 ;
        RECT -144.170 60.010 -143.930 60.020 ;
        RECT -143.420 59.260 -142.910 72.160 ;
        RECT -14.200 71.370 -14.030 72.130 ;
        RECT -13.170 71.730 -12.850 71.760 ;
        RECT -13.180 71.540 -12.850 71.730 ;
        RECT -13.170 71.500 -12.850 71.540 ;
        RECT -12.190 71.750 -12.020 73.680 ;
        RECT -11.640 73.540 -11.210 73.680 ;
        RECT -11.640 72.430 -11.470 73.540 ;
        RECT -11.640 72.170 -11.210 72.430 ;
        RECT -12.190 71.490 -11.750 71.750 ;
        RECT -12.190 71.180 -12.020 71.490 ;
        RECT -11.640 71.180 -11.470 72.170 ;
        RECT -11.090 71.750 -10.920 73.680 ;
        RECT -11.090 71.490 -10.660 71.750 ;
        RECT -11.090 71.180 -10.920 71.490 ;
        RECT -10.540 71.180 -10.370 73.680 ;
        RECT -9.990 71.180 -9.820 73.680 ;
        RECT -9.440 71.580 -9.270 73.670 ;
        RECT 17.830 72.850 18.000 75.340 ;
        RECT 18.380 73.320 18.550 75.340 ;
        RECT 18.930 73.320 19.100 75.340 ;
        RECT 19.300 75.120 19.470 75.460 ;
        RECT 19.850 75.450 20.010 75.490 ;
        RECT 19.300 75.110 19.460 75.120 ;
        RECT 19.480 75.080 19.650 75.340 ;
        RECT 19.850 75.120 20.020 75.450 ;
        RECT 19.850 75.110 20.010 75.120 ;
        RECT 19.210 74.820 19.650 75.080 ;
        RECT 19.480 73.710 19.650 74.820 ;
        RECT 19.210 73.450 19.650 73.710 ;
        RECT 18.380 72.840 19.100 73.320 ;
        RECT 19.480 72.840 19.650 73.450 ;
        RECT 20.030 73.030 20.200 75.340 ;
        RECT 20.400 75.120 20.570 75.520 ;
        RECT 20.950 75.450 21.110 75.490 ;
        RECT 21.500 75.450 21.660 75.490 ;
        RECT 22.050 75.470 22.210 75.490 ;
        RECT 25.030 75.470 25.190 75.490 ;
        RECT 20.400 75.110 20.560 75.120 ;
        RECT 20.580 75.080 20.750 75.340 ;
        RECT 20.950 75.120 21.120 75.450 ;
        RECT 21.500 75.120 21.670 75.450 ;
        RECT 22.050 75.120 22.220 75.470 ;
        RECT 25.020 75.120 25.190 75.470 ;
        RECT 25.580 75.450 25.740 75.490 ;
        RECT 26.130 75.450 26.290 75.490 ;
        RECT 25.570 75.120 25.740 75.450 ;
        RECT 26.120 75.120 26.290 75.450 ;
        RECT 20.950 75.110 21.110 75.120 ;
        RECT 21.500 75.110 21.660 75.120 ;
        RECT 22.050 75.110 22.210 75.120 ;
        RECT 25.030 75.110 25.190 75.120 ;
        RECT 25.580 75.110 25.740 75.120 ;
        RECT 26.130 75.110 26.290 75.120 ;
        RECT 26.490 75.080 26.660 75.340 ;
        RECT 26.670 75.120 26.840 75.520 ;
        RECT 29.110 75.490 29.270 75.520 ;
        RECT 27.230 75.450 27.390 75.490 ;
        RECT 27.780 75.460 27.940 75.490 ;
        RECT 26.680 75.110 26.840 75.120 ;
        RECT 20.310 74.820 20.750 75.080 ;
        RECT 21.410 75.040 21.730 75.080 ;
        RECT 25.510 75.040 25.830 75.080 ;
        RECT 21.410 74.850 21.740 75.040 ;
        RECT 25.500 74.850 25.830 75.040 ;
        RECT 21.410 74.820 21.730 74.850 ;
        RECT 25.510 74.820 25.830 74.850 ;
        RECT 26.490 74.820 26.930 75.080 ;
        RECT 20.580 73.710 20.750 74.820 ;
        RECT 26.490 73.710 26.660 74.820 ;
        RECT 20.310 73.450 20.750 73.710 ;
        RECT 21.410 73.670 21.730 73.710 ;
        RECT 25.510 73.670 25.830 73.710 ;
        RECT 21.410 73.480 21.740 73.670 ;
        RECT 25.500 73.480 25.830 73.670 ;
        RECT 21.410 73.450 21.730 73.480 ;
        RECT 25.510 73.450 25.830 73.480 ;
        RECT 26.490 73.450 26.930 73.710 ;
        RECT 19.770 72.840 20.200 73.030 ;
        RECT 20.580 72.840 20.750 73.450 ;
        RECT 20.860 72.990 21.180 73.030 ;
        RECT 21.960 73.000 22.280 73.040 ;
        RECT 24.960 73.000 25.280 73.040 ;
        RECT 18.540 72.310 19.050 72.840 ;
        RECT 19.770 72.800 20.100 72.840 ;
        RECT 20.860 72.800 21.190 72.990 ;
        RECT 21.960 72.810 22.290 73.000 ;
        RECT 24.950 72.810 25.280 73.000 ;
        RECT 26.060 72.990 26.380 73.030 ;
        RECT 19.770 72.770 20.090 72.800 ;
        RECT 20.860 72.770 21.180 72.800 ;
        RECT 21.960 72.780 22.280 72.810 ;
        RECT 24.960 72.780 25.280 72.810 ;
        RECT 26.050 72.800 26.380 72.990 ;
        RECT 26.490 72.840 26.660 73.450 ;
        RECT 27.040 73.030 27.210 75.340 ;
        RECT 27.220 75.120 27.390 75.450 ;
        RECT 27.770 75.370 27.940 75.460 ;
        RECT 27.640 75.340 27.940 75.370 ;
        RECT 28.190 75.340 28.360 75.370 ;
        RECT 28.740 75.340 28.910 75.370 ;
        RECT 27.230 75.110 27.390 75.120 ;
        RECT 27.590 75.110 27.940 75.340 ;
        RECT 27.590 75.080 27.810 75.110 ;
        RECT 27.590 74.820 28.030 75.080 ;
        RECT 27.590 73.710 27.810 74.820 ;
        RECT 27.590 73.450 28.030 73.710 ;
        RECT 27.040 72.840 27.470 73.030 ;
        RECT 27.590 72.880 27.810 73.450 ;
        RECT 28.140 73.350 28.360 75.340 ;
        RECT 28.690 73.350 28.910 75.340 ;
        RECT 29.110 75.340 29.280 75.490 ;
        RECT 29.660 75.480 29.820 75.520 ;
        RECT 29.290 75.340 29.460 75.370 ;
        RECT 29.110 75.140 29.460 75.340 ;
        RECT 29.660 75.150 29.830 75.480 ;
        RECT 29.660 75.140 29.820 75.150 ;
        RECT 29.240 75.110 29.460 75.140 ;
        RECT 29.020 74.850 29.460 75.110 ;
        RECT 29.240 73.740 29.460 74.850 ;
        RECT 29.020 73.480 29.460 73.740 ;
        RECT 27.590 72.840 27.760 72.880 ;
        RECT 28.140 72.870 28.910 73.350 ;
        RECT 29.240 72.870 29.460 73.480 ;
        RECT 29.840 73.060 30.010 75.370 ;
        RECT 30.210 75.150 30.380 75.550 ;
        RECT 30.760 75.480 30.920 75.520 ;
        RECT 31.310 75.480 31.470 75.520 ;
        RECT 31.860 75.500 32.020 75.520 ;
        RECT 34.840 75.500 35.000 75.520 ;
        RECT 30.210 75.140 30.370 75.150 ;
        RECT 30.390 75.110 30.560 75.370 ;
        RECT 30.760 75.150 30.930 75.480 ;
        RECT 31.310 75.150 31.480 75.480 ;
        RECT 31.860 75.150 32.030 75.500 ;
        RECT 34.830 75.150 35.000 75.500 ;
        RECT 35.390 75.480 35.550 75.520 ;
        RECT 35.940 75.480 36.100 75.520 ;
        RECT 35.380 75.150 35.550 75.480 ;
        RECT 35.930 75.150 36.100 75.480 ;
        RECT 30.760 75.140 30.920 75.150 ;
        RECT 31.310 75.140 31.470 75.150 ;
        RECT 31.860 75.140 32.020 75.150 ;
        RECT 34.840 75.140 35.000 75.150 ;
        RECT 35.390 75.140 35.550 75.150 ;
        RECT 35.940 75.140 36.100 75.150 ;
        RECT 36.300 75.110 36.470 75.370 ;
        RECT 36.480 75.150 36.650 75.550 ;
        RECT 37.040 75.480 37.200 75.520 ;
        RECT 37.590 75.490 37.750 75.520 ;
        RECT 36.490 75.140 36.650 75.150 ;
        RECT 30.120 74.850 30.560 75.110 ;
        RECT 31.220 75.070 31.540 75.110 ;
        RECT 35.320 75.070 35.640 75.110 ;
        RECT 31.220 74.880 31.550 75.070 ;
        RECT 35.310 74.880 35.640 75.070 ;
        RECT 31.220 74.850 31.540 74.880 ;
        RECT 35.320 74.850 35.640 74.880 ;
        RECT 36.300 74.850 36.740 75.110 ;
        RECT 30.390 73.740 30.560 74.850 ;
        RECT 36.300 73.740 36.470 74.850 ;
        RECT 30.120 73.480 30.560 73.740 ;
        RECT 31.220 73.700 31.540 73.740 ;
        RECT 35.320 73.700 35.640 73.740 ;
        RECT 31.220 73.510 31.550 73.700 ;
        RECT 35.310 73.510 35.640 73.700 ;
        RECT 31.220 73.480 31.540 73.510 ;
        RECT 35.320 73.480 35.640 73.510 ;
        RECT 36.300 73.480 36.740 73.740 ;
        RECT 29.580 72.870 30.010 73.060 ;
        RECT 30.390 72.870 30.560 73.480 ;
        RECT 30.670 73.020 30.990 73.060 ;
        RECT 31.770 73.030 32.090 73.070 ;
        RECT 34.770 73.030 35.090 73.070 ;
        RECT 28.140 72.840 28.860 72.870 ;
        RECT 29.240 72.850 29.410 72.870 ;
        RECT 27.140 72.800 27.470 72.840 ;
        RECT 26.060 72.770 26.380 72.800 ;
        RECT 27.150 72.770 27.470 72.800 ;
        RECT 28.190 72.340 28.860 72.840 ;
        RECT 29.580 72.830 29.910 72.870 ;
        RECT 30.670 72.830 31.000 73.020 ;
        RECT 31.770 72.840 32.100 73.030 ;
        RECT 34.760 72.840 35.090 73.030 ;
        RECT 35.870 73.020 36.190 73.060 ;
        RECT 29.580 72.800 29.900 72.830 ;
        RECT 30.670 72.800 30.990 72.830 ;
        RECT 31.770 72.810 32.090 72.840 ;
        RECT 34.770 72.810 35.090 72.840 ;
        RECT 35.860 72.830 36.190 73.020 ;
        RECT 36.300 72.870 36.470 73.480 ;
        RECT 36.850 73.060 37.020 75.370 ;
        RECT 37.030 75.150 37.200 75.480 ;
        RECT 37.040 75.140 37.200 75.150 ;
        RECT 37.400 75.110 37.570 75.370 ;
        RECT 37.580 75.150 37.750 75.490 ;
        RECT 37.590 75.140 37.750 75.150 ;
        RECT 37.400 74.850 37.840 75.110 ;
        RECT 37.400 73.740 37.570 74.850 ;
        RECT 37.400 73.480 37.840 73.740 ;
        RECT 36.850 72.870 37.280 73.060 ;
        RECT 37.400 72.870 37.570 73.480 ;
        RECT 37.950 73.350 38.120 75.370 ;
        RECT 38.500 73.350 38.670 75.370 ;
        RECT 37.950 72.870 38.670 73.350 ;
        RECT 39.050 72.880 39.220 75.370 ;
        RECT 40.580 73.050 40.750 75.560 ;
        RECT 41.130 75.090 41.300 77.600 ;
        RECT 41.680 77.170 41.850 77.900 ;
        RECT 42.230 77.870 42.400 77.900 ;
        RECT 42.160 77.830 42.480 77.870 ;
        RECT 42.150 77.640 42.480 77.830 ;
        RECT 42.160 77.610 42.480 77.640 ;
        RECT 41.610 77.130 41.930 77.170 ;
        RECT 41.600 76.940 41.930 77.130 ;
        RECT 41.610 76.910 41.930 76.940 ;
        RECT 41.680 75.820 41.850 76.910 ;
        RECT 41.610 75.780 41.930 75.820 ;
        RECT 41.600 75.590 41.930 75.780 ;
        RECT 41.610 75.560 41.930 75.590 ;
        RECT 41.060 75.050 41.380 75.090 ;
        RECT 41.050 74.860 41.380 75.050 ;
        RECT 41.060 74.830 41.380 74.860 ;
        RECT 41.130 73.720 41.300 74.830 ;
        RECT 41.060 73.680 41.380 73.720 ;
        RECT 41.050 73.490 41.380 73.680 ;
        RECT 41.060 73.460 41.380 73.490 ;
        RECT 40.510 73.010 40.830 73.050 ;
        RECT 36.950 72.830 37.280 72.870 ;
        RECT 35.870 72.800 36.190 72.830 ;
        RECT 36.960 72.800 37.280 72.830 ;
        RECT 38.000 72.340 38.510 72.870 ;
        RECT 40.500 72.820 40.830 73.010 ;
        RECT 40.510 72.790 40.830 72.820 ;
        RECT 40.580 72.720 40.750 72.790 ;
        RECT 41.130 72.720 41.300 73.460 ;
        RECT 41.680 73.040 41.850 75.560 ;
        RECT 42.230 75.090 42.400 77.610 ;
        RECT 42.780 77.190 42.950 77.900 ;
        RECT 43.330 77.870 43.500 77.900 ;
        RECT 43.250 77.830 43.570 77.870 ;
        RECT 43.240 77.640 43.570 77.830 ;
        RECT 43.250 77.610 43.570 77.640 ;
        RECT 42.700 77.150 43.020 77.190 ;
        RECT 42.690 76.960 43.020 77.150 ;
        RECT 42.700 76.930 43.020 76.960 ;
        RECT 42.780 75.820 42.950 76.930 ;
        RECT 42.700 75.780 43.020 75.820 ;
        RECT 42.690 75.590 43.020 75.780 ;
        RECT 42.700 75.560 43.020 75.590 ;
        RECT 42.160 75.050 42.480 75.090 ;
        RECT 42.150 74.860 42.480 75.050 ;
        RECT 42.160 74.830 42.480 74.860 ;
        RECT 42.230 73.720 42.400 74.830 ;
        RECT 42.160 73.680 42.480 73.720 ;
        RECT 42.150 73.490 42.480 73.680 ;
        RECT 42.160 73.460 42.480 73.490 ;
        RECT 41.610 73.000 41.930 73.040 ;
        RECT 41.600 72.810 41.930 73.000 ;
        RECT 41.610 72.780 41.930 72.810 ;
        RECT 41.680 72.720 41.850 72.780 ;
        RECT 42.230 72.720 42.400 73.460 ;
        RECT 42.780 73.040 42.950 75.560 ;
        RECT 43.330 75.090 43.500 77.610 ;
        RECT 206.500 76.260 207.010 86.620 ;
        RECT 207.180 85.830 213.160 86.060 ;
        RECT 206.500 76.240 207.020 76.260 ;
        RECT 43.260 75.050 43.580 75.090 ;
        RECT 43.250 74.860 43.580 75.050 ;
        RECT 43.260 74.830 43.580 74.860 ;
        RECT 43.330 73.720 43.500 74.830 ;
        RECT 43.260 73.680 43.580 73.720 ;
        RECT 43.250 73.490 43.580 73.680 ;
        RECT 44.040 73.520 44.210 74.710 ;
        RECT 43.260 73.460 43.580 73.490 ;
        RECT 42.700 73.000 43.020 73.040 ;
        RECT 42.690 72.810 43.020 73.000 ;
        RECT 42.700 72.780 43.020 72.810 ;
        RECT 42.780 72.720 42.950 72.780 ;
        RECT 43.330 72.720 43.500 73.460 ;
        RECT 43.750 73.070 44.260 73.330 ;
        RECT 43.740 73.000 44.260 73.070 ;
        RECT 28.190 72.310 28.700 72.340 ;
        RECT 43.740 72.320 44.250 73.000 ;
        RECT -9.550 71.210 -7.160 71.580 ;
        RECT -9.500 67.950 -7.160 71.210 ;
        RECT 69.250 70.410 69.480 70.420 ;
        RECT 69.230 70.240 73.890 70.410 ;
        RECT 69.250 70.230 69.480 70.240 ;
        RECT 74.790 69.760 74.980 69.770 ;
        RECT 70.450 69.720 74.250 69.730 ;
        RECT 74.760 69.720 75.020 69.760 ;
        RECT 70.450 69.560 75.020 69.720 ;
        RECT 74.020 69.550 75.020 69.560 ;
        RECT 74.020 69.090 74.250 69.550 ;
        RECT 74.760 69.440 75.020 69.550 ;
        RECT 74.790 69.090 74.980 69.100 ;
        RECT 74.020 68.880 75.030 69.090 ;
        RECT 69.250 68.800 69.480 68.810 ;
        RECT 69.230 68.630 73.710 68.800 ;
        RECT 69.250 68.620 69.480 68.630 ;
        RECT 74.020 68.120 74.250 68.880 ;
        RECT 74.760 68.770 75.020 68.880 ;
        RECT 70.470 67.950 74.250 68.120 ;
        RECT -9.500 67.940 -7.170 67.950 ;
        RECT 69.250 67.200 69.480 67.210 ;
        RECT 69.230 67.030 73.730 67.200 ;
        RECT 69.250 67.020 69.480 67.030 ;
        RECT 70.470 67.020 70.800 67.030 ;
        RECT 71.430 67.020 71.760 67.030 ;
        RECT 72.390 67.020 72.720 67.030 ;
        RECT 73.350 67.020 73.680 67.030 ;
        RECT 74.020 66.510 74.250 67.950 ;
        RECT 74.700 67.760 75.130 67.780 ;
        RECT 74.680 67.590 75.130 67.760 ;
        RECT 74.700 67.570 75.130 67.590 ;
        RECT 70.470 66.340 74.250 66.510 ;
        RECT 70.530 66.110 70.960 66.130 ;
        RECT 70.510 65.940 70.960 66.110 ;
        RECT 70.530 65.920 70.960 65.940 ;
        RECT 69.250 65.580 69.480 65.590 ;
        RECT 69.230 65.410 73.730 65.580 ;
        RECT 69.250 65.400 69.480 65.410 ;
        RECT 74.020 64.910 74.250 66.340 ;
        RECT 74.700 66.150 75.130 66.170 ;
        RECT 74.680 65.980 75.130 66.150 ;
        RECT 74.700 65.960 75.130 65.980 ;
        RECT 70.480 64.900 74.250 64.910 ;
        RECT 70.470 64.740 74.250 64.900 ;
        RECT 70.470 64.730 70.800 64.740 ;
        RECT 72.390 64.730 72.720 64.740 ;
        RECT 73.350 64.730 73.680 64.740 ;
        RECT 71.530 64.370 71.960 64.390 ;
        RECT 71.530 64.200 71.980 64.370 ;
        RECT 71.530 64.180 71.960 64.200 ;
        RECT 69.250 63.980 69.480 63.990 ;
        RECT 69.230 63.810 73.680 63.980 ;
        RECT 69.250 63.800 69.480 63.810 ;
        RECT 70.470 63.800 70.800 63.810 ;
        RECT 71.430 63.800 71.760 63.810 ;
        RECT 72.390 63.800 72.720 63.810 ;
        RECT 73.350 63.800 73.680 63.810 ;
        RECT 74.020 63.290 74.250 64.740 ;
        RECT 74.690 64.540 75.120 64.560 ;
        RECT 74.670 64.370 75.120 64.540 ;
        RECT 74.690 64.350 75.120 64.370 ;
        RECT 70.460 63.120 74.250 63.290 ;
        RECT 72.440 62.860 72.870 62.880 ;
        RECT 72.420 62.690 72.870 62.860 ;
        RECT 72.440 62.670 72.870 62.690 ;
        RECT 69.250 62.360 69.480 62.370 ;
        RECT 69.230 62.190 73.730 62.360 ;
        RECT 69.250 62.180 69.480 62.190 ;
        RECT 70.470 61.670 70.800 61.680 ;
        RECT 71.430 61.670 71.760 61.680 ;
        RECT 72.390 61.670 72.720 61.680 ;
        RECT 73.350 61.670 73.680 61.680 ;
        RECT 74.020 61.670 74.250 63.120 ;
        RECT 74.690 62.920 75.120 62.940 ;
        RECT 74.670 62.750 75.120 62.920 ;
        RECT 74.690 62.730 75.120 62.750 ;
        RECT 70.460 61.500 74.250 61.670 ;
        RECT 69.250 60.760 69.480 60.770 ;
        RECT 69.230 60.750 73.650 60.760 ;
        RECT 69.230 60.590 73.680 60.750 ;
        RECT 69.250 60.580 69.480 60.590 ;
        RECT 70.470 60.580 70.800 60.590 ;
        RECT 71.430 60.580 71.760 60.590 ;
        RECT 72.390 60.580 72.720 60.590 ;
        RECT 73.350 60.580 73.680 60.590 ;
        RECT 74.020 60.080 74.250 61.500 ;
        RECT 74.690 61.310 75.120 61.330 ;
        RECT 74.670 61.140 75.120 61.310 ;
        RECT 74.690 61.120 75.120 61.140 ;
        RECT 80.680 60.950 81.050 75.820 ;
        RECT 206.490 74.460 207.020 76.240 ;
        RECT 207.420 74.770 213.070 85.830 ;
        RECT 207.360 74.760 213.070 74.770 ;
        RECT 207.360 74.590 213.150 74.760 ;
        RECT 207.360 74.580 213.060 74.590 ;
        RECT 207.420 74.510 207.590 74.580 ;
        RECT 206.490 74.440 207.010 74.460 ;
        RECT 206.500 73.930 207.010 74.440 ;
        RECT 213.520 74.010 214.030 86.620 ;
        RECT 214.270 80.600 215.730 80.640 ;
        RECT 214.260 80.430 215.730 80.600 ;
        RECT 214.270 80.390 215.730 80.430 ;
        RECT 206.480 73.720 207.010 73.930 ;
        RECT 211.590 73.720 214.030 74.010 ;
        RECT 206.480 73.240 214.030 73.720 ;
        RECT 206.670 73.210 214.030 73.240 ;
        RECT 206.500 71.450 214.030 72.000 ;
        RECT 206.500 71.440 207.170 71.450 ;
        RECT 80.680 60.700 81.060 60.950 ;
        RECT 70.460 59.910 74.260 60.080 ;
        RECT 70.470 59.900 70.800 59.910 ;
        RECT 71.430 59.900 71.760 59.910 ;
        RECT 72.390 59.900 72.720 59.910 ;
        RECT 73.350 59.900 73.680 59.910 ;
        RECT -150.440 58.750 -142.910 59.260 ;
        RECT 69.250 59.130 69.480 59.150 ;
        RECT 70.470 59.130 70.800 59.140 ;
        RECT 71.430 59.130 71.760 59.140 ;
        RECT 72.390 59.130 72.720 59.140 ;
        RECT 73.350 59.130 73.680 59.140 ;
        RECT 69.230 58.960 73.690 59.130 ;
        RECT -152.140 52.730 -150.680 52.770 ;
        RECT -152.140 52.560 -150.670 52.730 ;
        RECT -152.140 52.520 -150.680 52.560 ;
        RECT -150.440 46.140 -149.930 58.750 ;
        RECT -149.570 57.960 -143.590 58.190 ;
        RECT -149.480 46.900 -143.830 57.960 ;
        RECT -143.420 48.390 -142.910 58.750 ;
        RECT 74.020 58.470 74.250 59.910 ;
        RECT 74.530 59.320 74.740 59.750 ;
        RECT 74.550 59.300 74.720 59.320 ;
        RECT 70.460 58.300 74.250 58.470 ;
        RECT 206.500 58.540 207.010 71.440 ;
        RECT 207.410 70.550 210.870 70.990 ;
        RECT 207.410 70.450 212.800 70.550 ;
        RECT 207.520 70.380 212.800 70.450 ;
        RECT 207.520 59.470 207.690 70.380 ;
        RECT 208.070 69.970 212.300 69.990 ;
        RECT 207.990 59.860 212.320 69.970 ;
        RECT 212.090 59.810 212.260 59.860 ;
        RECT 212.630 59.470 212.800 70.380 ;
        RECT 207.520 59.300 212.800 59.470 ;
        RECT 207.520 59.290 207.760 59.300 ;
        RECT 213.520 58.540 214.030 71.450 ;
        RECT 70.470 58.290 70.800 58.300 ;
        RECT 71.430 58.290 71.760 58.300 ;
        RECT 72.390 58.290 72.720 58.300 ;
        RECT 73.350 58.290 73.680 58.300 ;
        RECT 74.700 58.110 75.130 58.130 ;
        RECT 74.680 57.940 75.130 58.110 ;
        RECT 74.700 57.920 75.130 57.940 ;
        RECT 206.500 58.030 214.030 58.540 ;
        RECT 214.240 58.480 215.710 58.730 ;
        RECT 74.690 56.520 75.120 56.540 ;
        RECT 71.490 56.440 71.920 56.460 ;
        RECT 72.430 56.440 72.860 56.460 ;
        RECT 71.470 56.270 71.920 56.440 ;
        RECT 72.410 56.270 72.860 56.440 ;
        RECT 73.380 56.380 73.810 56.400 ;
        RECT 71.490 56.250 71.920 56.270 ;
        RECT 72.430 56.250 72.860 56.270 ;
        RECT 73.360 56.210 73.810 56.380 ;
        RECT 74.670 56.350 75.120 56.520 ;
        RECT 74.690 56.330 75.120 56.350 ;
        RECT 73.380 56.190 73.810 56.210 ;
        RECT -143.430 48.370 -142.910 48.390 ;
        RECT -149.480 46.890 -143.770 46.900 ;
        RECT -149.560 46.720 -143.770 46.890 ;
        RECT -149.470 46.710 -143.770 46.720 ;
        RECT -144.000 46.640 -143.830 46.710 ;
        RECT -143.430 46.590 -142.900 48.370 ;
        RECT 206.500 47.670 207.010 58.030 ;
        RECT 207.180 57.240 213.160 57.470 ;
        RECT 206.500 47.650 207.020 47.670 ;
        RECT -143.420 46.570 -142.900 46.590 ;
        RECT -150.440 45.850 -148.000 46.140 ;
        RECT -143.420 46.060 -142.910 46.570 ;
        RECT -143.420 45.850 -142.890 46.060 ;
        RECT 206.490 45.870 207.020 47.650 ;
        RECT 207.420 46.180 213.070 57.240 ;
        RECT 207.360 46.170 213.070 46.180 ;
        RECT 207.360 46.000 213.150 46.170 ;
        RECT 207.360 45.990 213.060 46.000 ;
        RECT 207.420 45.920 207.590 45.990 ;
        RECT 206.490 45.850 207.010 45.870 ;
        RECT -150.440 45.370 -142.890 45.850 ;
        RECT -150.440 45.340 -143.080 45.370 ;
        RECT 206.500 45.340 207.010 45.850 ;
        RECT 213.520 45.420 214.030 58.030 ;
        RECT 214.270 52.010 215.730 52.050 ;
        RECT 214.260 51.840 215.730 52.010 ;
        RECT 214.270 51.800 215.730 51.840 ;
        RECT 206.480 45.130 207.010 45.340 ;
        RECT 211.590 45.130 214.030 45.420 ;
        RECT 206.480 44.650 214.030 45.130 ;
        RECT 206.670 44.620 214.030 44.650 ;
        RECT -150.440 43.580 -142.910 44.130 ;
        RECT -152.120 30.610 -150.650 30.860 ;
        RECT -150.440 30.670 -149.930 43.580 ;
        RECT -143.580 43.570 -142.910 43.580 ;
        RECT -147.280 42.680 -143.820 43.120 ;
        RECT -149.210 42.580 -143.820 42.680 ;
        RECT -149.210 42.510 -143.930 42.580 ;
        RECT -149.210 31.600 -149.040 42.510 ;
        RECT -148.710 42.100 -144.480 42.120 ;
        RECT -148.730 31.990 -144.400 42.100 ;
        RECT -148.670 31.940 -148.500 31.990 ;
        RECT -144.100 31.600 -143.930 42.510 ;
        RECT -149.210 31.430 -143.930 31.600 ;
        RECT -144.170 31.420 -143.930 31.430 ;
        RECT -143.420 30.670 -142.910 43.570 ;
        RECT -150.440 30.160 -142.910 30.670 ;
        RECT -152.140 24.140 -150.680 24.180 ;
        RECT -152.140 23.970 -150.670 24.140 ;
        RECT -152.140 23.930 -150.680 23.970 ;
        RECT -150.440 17.550 -149.930 30.160 ;
        RECT -149.570 29.370 -143.590 29.600 ;
        RECT -149.480 18.310 -143.830 29.370 ;
        RECT -143.420 19.800 -142.910 30.160 ;
        RECT -143.430 19.780 -142.910 19.800 ;
        RECT 206.500 42.860 214.030 43.410 ;
        RECT 206.500 42.850 207.170 42.860 ;
        RECT 206.500 29.950 207.010 42.850 ;
        RECT 207.410 41.960 210.870 42.400 ;
        RECT 207.410 41.860 212.800 41.960 ;
        RECT 207.520 41.790 212.800 41.860 ;
        RECT 207.520 30.880 207.690 41.790 ;
        RECT 208.070 41.380 212.300 41.400 ;
        RECT 207.990 31.270 212.320 41.380 ;
        RECT 212.090 31.220 212.260 31.270 ;
        RECT 212.630 30.880 212.800 41.790 ;
        RECT 207.520 30.710 212.800 30.880 ;
        RECT 207.520 30.700 207.760 30.710 ;
        RECT 213.520 29.950 214.030 42.860 ;
        RECT 206.500 29.440 214.030 29.950 ;
        RECT 214.240 29.890 215.710 30.140 ;
        RECT -149.480 18.300 -143.770 18.310 ;
        RECT -149.560 18.130 -143.770 18.300 ;
        RECT -149.470 18.120 -143.770 18.130 ;
        RECT -144.000 18.050 -143.830 18.120 ;
        RECT -143.430 18.000 -142.900 19.780 ;
        RECT 206.500 19.080 207.010 29.440 ;
        RECT 207.180 28.650 213.160 28.880 ;
        RECT 206.500 19.060 207.020 19.080 ;
        RECT -143.420 17.980 -142.900 18.000 ;
        RECT -150.440 17.260 -148.000 17.550 ;
        RECT -143.420 17.470 -142.910 17.980 ;
        RECT -143.420 17.260 -142.890 17.470 ;
        RECT 206.490 17.280 207.020 19.060 ;
        RECT 207.420 17.590 213.070 28.650 ;
        RECT 207.360 17.580 213.070 17.590 ;
        RECT 207.360 17.410 213.150 17.580 ;
        RECT 207.360 17.400 213.060 17.410 ;
        RECT 207.420 17.330 207.590 17.400 ;
        RECT 206.490 17.260 207.010 17.280 ;
        RECT -150.440 16.780 -142.890 17.260 ;
        RECT -150.440 16.750 -143.080 16.780 ;
        RECT 206.500 16.750 207.010 17.260 ;
        RECT 213.520 16.830 214.030 29.440 ;
        RECT 214.270 23.420 215.730 23.460 ;
        RECT 214.260 23.250 215.730 23.420 ;
        RECT 214.270 23.210 215.730 23.250 ;
        RECT 206.480 16.540 207.010 16.750 ;
        RECT 211.590 16.540 214.030 16.830 ;
        RECT 206.480 16.060 214.030 16.540 ;
        RECT 206.670 16.030 214.030 16.060 ;
        RECT -150.440 14.990 -142.910 15.540 ;
        RECT -152.120 2.020 -150.650 2.270 ;
        RECT -150.440 2.080 -149.930 14.990 ;
        RECT -143.580 14.980 -142.910 14.990 ;
        RECT -147.280 14.090 -143.820 14.530 ;
        RECT -149.210 13.990 -143.820 14.090 ;
        RECT -149.210 13.920 -143.930 13.990 ;
        RECT -149.210 3.010 -149.040 13.920 ;
        RECT -148.710 13.510 -144.480 13.530 ;
        RECT -148.730 3.400 -144.400 13.510 ;
        RECT -148.670 3.350 -148.500 3.400 ;
        RECT -144.100 3.010 -143.930 13.920 ;
        RECT -149.210 2.840 -143.930 3.010 ;
        RECT -144.170 2.830 -143.930 2.840 ;
        RECT -143.420 2.080 -142.910 14.980 ;
        RECT -150.440 1.570 -142.910 2.080 ;
        RECT -152.140 -4.450 -150.680 -4.410 ;
        RECT -152.140 -4.620 -150.670 -4.450 ;
        RECT -152.140 -4.660 -150.680 -4.620 ;
        RECT -150.440 -11.040 -149.930 1.570 ;
        RECT -149.570 0.780 -143.590 1.010 ;
        RECT -149.480 -10.280 -143.830 0.780 ;
        RECT -143.420 -8.790 -142.910 1.570 ;
        RECT -143.430 -8.810 -142.910 -8.790 ;
        RECT 206.500 14.270 214.030 14.820 ;
        RECT 206.500 14.260 207.170 14.270 ;
        RECT 206.500 1.360 207.010 14.260 ;
        RECT 207.410 13.370 210.870 13.810 ;
        RECT 207.410 13.270 212.800 13.370 ;
        RECT 207.520 13.200 212.800 13.270 ;
        RECT 207.520 2.290 207.690 13.200 ;
        RECT 208.070 12.790 212.300 12.810 ;
        RECT 207.990 2.680 212.320 12.790 ;
        RECT 212.090 2.630 212.260 2.680 ;
        RECT 212.630 2.290 212.800 13.200 ;
        RECT 207.520 2.120 212.800 2.290 ;
        RECT 207.520 2.110 207.760 2.120 ;
        RECT 213.520 1.360 214.030 14.270 ;
        RECT 206.500 0.850 214.030 1.360 ;
        RECT 214.240 1.300 215.710 1.550 ;
        RECT -149.480 -10.290 -143.770 -10.280 ;
        RECT -149.560 -10.460 -143.770 -10.290 ;
        RECT -149.470 -10.470 -143.770 -10.460 ;
        RECT -144.000 -10.540 -143.830 -10.470 ;
        RECT -143.430 -10.590 -142.900 -8.810 ;
        RECT 206.500 -9.510 207.010 0.850 ;
        RECT 207.180 0.060 213.160 0.290 ;
        RECT 206.500 -9.530 207.020 -9.510 ;
        RECT -143.420 -10.610 -142.900 -10.590 ;
        RECT -150.440 -11.330 -148.000 -11.040 ;
        RECT -143.420 -11.120 -142.910 -10.610 ;
        RECT -143.420 -11.330 -142.890 -11.120 ;
        RECT 206.490 -11.310 207.020 -9.530 ;
        RECT 207.420 -11.000 213.070 0.060 ;
        RECT 207.360 -11.010 213.070 -11.000 ;
        RECT 207.360 -11.180 213.150 -11.010 ;
        RECT 207.360 -11.190 213.060 -11.180 ;
        RECT 207.420 -11.260 207.590 -11.190 ;
        RECT 206.490 -11.330 207.010 -11.310 ;
        RECT -150.440 -11.810 -142.890 -11.330 ;
        RECT -150.440 -11.840 -143.080 -11.810 ;
        RECT 206.500 -11.840 207.010 -11.330 ;
        RECT 213.520 -11.760 214.030 0.850 ;
        RECT 214.270 -5.170 215.730 -5.130 ;
        RECT 214.260 -5.340 215.730 -5.170 ;
        RECT 214.270 -5.380 215.730 -5.340 ;
        RECT 206.480 -12.050 207.010 -11.840 ;
        RECT 211.590 -12.050 214.030 -11.760 ;
        RECT 206.480 -12.530 214.030 -12.050 ;
        RECT 206.670 -12.560 214.030 -12.530 ;
        RECT -150.440 -13.600 -142.910 -13.050 ;
        RECT -152.120 -26.570 -150.650 -26.320 ;
        RECT -150.440 -26.510 -149.930 -13.600 ;
        RECT -143.580 -13.610 -142.910 -13.600 ;
        RECT -147.280 -14.500 -143.820 -14.060 ;
        RECT -149.210 -14.600 -143.820 -14.500 ;
        RECT -149.210 -14.670 -143.930 -14.600 ;
        RECT -149.210 -25.580 -149.040 -14.670 ;
        RECT -148.710 -15.080 -144.480 -15.060 ;
        RECT -148.730 -25.190 -144.400 -15.080 ;
        RECT -148.670 -25.240 -148.500 -25.190 ;
        RECT -144.100 -25.580 -143.930 -14.670 ;
        RECT -149.210 -25.750 -143.930 -25.580 ;
        RECT -144.170 -25.760 -143.930 -25.750 ;
        RECT -143.420 -26.510 -142.910 -13.610 ;
        RECT -150.440 -27.020 -142.910 -26.510 ;
        RECT -152.140 -33.040 -150.680 -33.000 ;
        RECT -152.140 -33.210 -150.670 -33.040 ;
        RECT -152.140 -33.250 -150.680 -33.210 ;
        RECT -150.440 -39.630 -149.930 -27.020 ;
        RECT -149.570 -27.810 -143.590 -27.580 ;
        RECT -149.480 -38.870 -143.830 -27.810 ;
        RECT -143.420 -37.380 -142.910 -27.020 ;
        RECT -143.430 -37.400 -142.910 -37.380 ;
        RECT 206.500 -14.320 214.030 -13.770 ;
        RECT 206.500 -14.330 207.170 -14.320 ;
        RECT 206.500 -27.230 207.010 -14.330 ;
        RECT 207.410 -15.220 210.870 -14.780 ;
        RECT 207.410 -15.320 212.800 -15.220 ;
        RECT 207.520 -15.390 212.800 -15.320 ;
        RECT 207.520 -26.300 207.690 -15.390 ;
        RECT 208.070 -15.800 212.300 -15.780 ;
        RECT 207.990 -25.910 212.320 -15.800 ;
        RECT 212.090 -25.960 212.260 -25.910 ;
        RECT 212.630 -26.300 212.800 -15.390 ;
        RECT 207.520 -26.470 212.800 -26.300 ;
        RECT 207.520 -26.480 207.760 -26.470 ;
        RECT 213.520 -27.230 214.030 -14.320 ;
        RECT 206.500 -27.740 214.030 -27.230 ;
        RECT 214.240 -27.290 215.710 -27.040 ;
        RECT -149.480 -38.880 -143.770 -38.870 ;
        RECT -149.560 -39.050 -143.770 -38.880 ;
        RECT -149.470 -39.060 -143.770 -39.050 ;
        RECT -144.000 -39.130 -143.830 -39.060 ;
        RECT -143.430 -39.180 -142.900 -37.400 ;
        RECT 206.500 -38.100 207.010 -27.740 ;
        RECT 207.180 -28.530 213.160 -28.300 ;
        RECT 206.500 -38.120 207.020 -38.100 ;
        RECT -143.420 -39.200 -142.900 -39.180 ;
        RECT -150.440 -39.920 -148.000 -39.630 ;
        RECT -143.420 -39.710 -142.910 -39.200 ;
        RECT -143.420 -39.920 -142.890 -39.710 ;
        RECT 206.490 -39.900 207.020 -38.120 ;
        RECT 207.420 -39.590 213.070 -28.530 ;
        RECT 207.360 -39.600 213.070 -39.590 ;
        RECT 207.360 -39.770 213.150 -39.600 ;
        RECT 207.360 -39.780 213.060 -39.770 ;
        RECT 207.420 -39.850 207.590 -39.780 ;
        RECT 206.490 -39.920 207.010 -39.900 ;
        RECT -150.440 -40.400 -142.890 -39.920 ;
        RECT -150.440 -40.430 -143.080 -40.400 ;
        RECT 206.500 -40.430 207.010 -39.920 ;
        RECT 213.520 -40.350 214.030 -27.740 ;
        RECT 214.270 -33.760 215.730 -33.720 ;
        RECT 214.260 -33.930 215.730 -33.760 ;
        RECT 214.270 -33.970 215.730 -33.930 ;
        RECT 206.480 -40.640 207.010 -40.430 ;
        RECT 211.590 -40.640 214.030 -40.350 ;
        RECT 206.480 -41.120 214.030 -40.640 ;
        RECT 206.670 -41.150 214.030 -41.120 ;
        RECT -150.440 -42.190 -142.910 -41.640 ;
        RECT -152.120 -55.160 -150.650 -54.910 ;
        RECT -150.440 -55.100 -149.930 -42.190 ;
        RECT -143.580 -42.200 -142.910 -42.190 ;
        RECT -147.280 -43.090 -143.820 -42.650 ;
        RECT -149.210 -43.190 -143.820 -43.090 ;
        RECT -149.210 -43.260 -143.930 -43.190 ;
        RECT -149.210 -54.170 -149.040 -43.260 ;
        RECT -148.710 -43.670 -144.480 -43.650 ;
        RECT -148.730 -53.780 -144.400 -43.670 ;
        RECT -148.670 -53.830 -148.500 -53.780 ;
        RECT -144.100 -54.170 -143.930 -43.260 ;
        RECT -149.210 -54.340 -143.930 -54.170 ;
        RECT -144.170 -54.350 -143.930 -54.340 ;
        RECT -143.420 -55.100 -142.910 -42.200 ;
        RECT -150.440 -55.610 -142.910 -55.100 ;
        RECT -152.140 -61.630 -150.680 -61.590 ;
        RECT -152.140 -61.800 -150.670 -61.630 ;
        RECT -152.140 -61.840 -150.680 -61.800 ;
        RECT -150.440 -68.220 -149.930 -55.610 ;
        RECT -149.570 -56.400 -143.590 -56.170 ;
        RECT -149.480 -67.460 -143.830 -56.400 ;
        RECT -143.420 -65.970 -142.910 -55.610 ;
        RECT -143.430 -65.990 -142.910 -65.970 ;
        RECT 206.500 -42.910 214.030 -42.360 ;
        RECT 206.500 -42.920 207.170 -42.910 ;
        RECT 206.500 -55.820 207.010 -42.920 ;
        RECT 207.410 -43.810 210.870 -43.370 ;
        RECT 207.410 -43.910 212.800 -43.810 ;
        RECT 207.520 -43.980 212.800 -43.910 ;
        RECT 207.520 -54.890 207.690 -43.980 ;
        RECT 208.070 -44.390 212.300 -44.370 ;
        RECT 207.990 -54.500 212.320 -44.390 ;
        RECT 212.090 -54.550 212.260 -54.500 ;
        RECT 212.630 -54.890 212.800 -43.980 ;
        RECT 207.520 -55.060 212.800 -54.890 ;
        RECT 207.520 -55.070 207.760 -55.060 ;
        RECT 213.520 -55.820 214.030 -42.910 ;
        RECT 206.500 -56.330 214.030 -55.820 ;
        RECT 214.240 -55.880 215.710 -55.630 ;
        RECT -149.480 -67.470 -143.770 -67.460 ;
        RECT -149.560 -67.640 -143.770 -67.470 ;
        RECT -149.470 -67.650 -143.770 -67.640 ;
        RECT -144.000 -67.720 -143.830 -67.650 ;
        RECT -143.430 -67.770 -142.900 -65.990 ;
        RECT 206.500 -66.690 207.010 -56.330 ;
        RECT 207.180 -57.120 213.160 -56.890 ;
        RECT 206.500 -66.710 207.020 -66.690 ;
        RECT -143.420 -67.790 -142.900 -67.770 ;
        RECT -150.440 -68.510 -148.000 -68.220 ;
        RECT -143.420 -68.300 -142.910 -67.790 ;
        RECT -143.420 -68.510 -142.890 -68.300 ;
        RECT 206.490 -68.490 207.020 -66.710 ;
        RECT 207.420 -68.180 213.070 -57.120 ;
        RECT 207.360 -68.190 213.070 -68.180 ;
        RECT 207.360 -68.360 213.150 -68.190 ;
        RECT 207.360 -68.370 213.060 -68.360 ;
        RECT 207.420 -68.440 207.590 -68.370 ;
        RECT 206.490 -68.510 207.010 -68.490 ;
        RECT -150.440 -68.990 -142.890 -68.510 ;
        RECT -150.440 -69.020 -143.080 -68.990 ;
        RECT 206.500 -69.020 207.010 -68.510 ;
        RECT 213.520 -68.940 214.030 -56.330 ;
        RECT 214.270 -62.350 215.730 -62.310 ;
        RECT 214.260 -62.520 215.730 -62.350 ;
        RECT 214.270 -62.560 215.730 -62.520 ;
        RECT 206.480 -69.230 207.010 -69.020 ;
        RECT 211.590 -69.230 214.030 -68.940 ;
        RECT 206.480 -69.710 214.030 -69.230 ;
        RECT 206.670 -69.740 214.030 -69.710 ;
        RECT -150.440 -70.780 -142.910 -70.230 ;
        RECT -152.120 -83.750 -150.650 -83.500 ;
        RECT -150.440 -83.690 -149.930 -70.780 ;
        RECT -143.580 -70.790 -142.910 -70.780 ;
        RECT -147.280 -71.680 -143.820 -71.240 ;
        RECT -149.210 -71.780 -143.820 -71.680 ;
        RECT -149.210 -71.850 -143.930 -71.780 ;
        RECT -149.210 -82.760 -149.040 -71.850 ;
        RECT -148.710 -72.260 -144.480 -72.240 ;
        RECT -148.730 -82.370 -144.400 -72.260 ;
        RECT -148.670 -82.420 -148.500 -82.370 ;
        RECT -144.100 -82.760 -143.930 -71.850 ;
        RECT -149.210 -82.930 -143.930 -82.760 ;
        RECT -144.170 -82.940 -143.930 -82.930 ;
        RECT -143.420 -83.690 -142.910 -70.790 ;
        RECT -150.440 -84.200 -142.910 -83.690 ;
        RECT -152.140 -90.220 -150.680 -90.180 ;
        RECT -152.140 -90.390 -150.670 -90.220 ;
        RECT -152.140 -90.430 -150.680 -90.390 ;
        RECT -150.440 -96.810 -149.930 -84.200 ;
        RECT -149.570 -84.990 -143.590 -84.760 ;
        RECT -149.480 -96.050 -143.830 -84.990 ;
        RECT -143.420 -94.560 -142.910 -84.200 ;
        RECT -143.430 -94.580 -142.910 -94.560 ;
        RECT -149.480 -96.060 -143.770 -96.050 ;
        RECT -149.560 -96.230 -143.770 -96.060 ;
        RECT -149.470 -96.240 -143.770 -96.230 ;
        RECT -144.000 -96.310 -143.830 -96.240 ;
        RECT -143.430 -96.360 -142.900 -94.580 ;
        RECT -143.420 -96.380 -142.900 -96.360 ;
        RECT -150.440 -97.100 -148.000 -96.810 ;
        RECT -143.420 -96.890 -142.910 -96.380 ;
        RECT -143.420 -97.100 -142.890 -96.890 ;
        RECT -150.440 -97.580 -142.890 -97.100 ;
        RECT -150.440 -97.610 -143.080 -97.580 ;
        RECT -150.440 -99.370 -142.910 -98.820 ;
        RECT -152.120 -112.340 -150.650 -112.090 ;
        RECT -150.440 -112.280 -149.930 -99.370 ;
        RECT -143.580 -99.380 -142.910 -99.370 ;
        RECT -147.280 -100.270 -143.820 -99.830 ;
        RECT -149.210 -100.370 -143.820 -100.270 ;
        RECT -149.210 -100.440 -143.930 -100.370 ;
        RECT -149.210 -111.350 -149.040 -100.440 ;
        RECT -148.710 -100.850 -144.480 -100.830 ;
        RECT -148.730 -110.960 -144.400 -100.850 ;
        RECT -148.670 -111.010 -148.500 -110.960 ;
        RECT -144.100 -111.350 -143.930 -100.440 ;
        RECT -149.210 -111.520 -143.930 -111.350 ;
        RECT -144.170 -111.530 -143.930 -111.520 ;
        RECT -143.420 -112.280 -142.910 -99.380 ;
        RECT -150.440 -112.790 -142.910 -112.280 ;
        RECT -152.140 -118.810 -150.680 -118.770 ;
        RECT -152.140 -118.980 -150.670 -118.810 ;
        RECT -152.140 -119.020 -150.680 -118.980 ;
        RECT -150.440 -125.400 -149.930 -112.790 ;
        RECT -149.570 -113.580 -143.590 -113.350 ;
        RECT -149.480 -124.640 -143.830 -113.580 ;
        RECT -143.420 -123.150 -142.910 -112.790 ;
        RECT -143.430 -123.170 -142.910 -123.150 ;
        RECT -149.480 -124.650 -143.770 -124.640 ;
        RECT -149.560 -124.820 -143.770 -124.650 ;
        RECT -149.470 -124.830 -143.770 -124.820 ;
        RECT -144.000 -124.900 -143.830 -124.830 ;
        RECT -143.430 -124.950 -142.900 -123.170 ;
        RECT -143.420 -124.970 -142.900 -124.950 ;
        RECT -150.440 -125.690 -148.000 -125.400 ;
        RECT -143.420 -125.480 -142.910 -124.970 ;
        RECT -143.420 -125.690 -142.890 -125.480 ;
        RECT -150.440 -126.170 -142.890 -125.690 ;
        RECT -150.440 -126.200 -143.080 -126.170 ;
        RECT -150.440 -127.960 -142.910 -127.410 ;
        RECT -152.120 -140.930 -150.650 -140.680 ;
        RECT -150.440 -140.870 -149.930 -127.960 ;
        RECT -143.580 -127.970 -142.910 -127.960 ;
        RECT -147.280 -128.860 -143.820 -128.420 ;
        RECT -149.210 -128.960 -143.820 -128.860 ;
        RECT -149.210 -129.030 -143.930 -128.960 ;
        RECT -149.210 -139.940 -149.040 -129.030 ;
        RECT -148.710 -129.440 -144.480 -129.420 ;
        RECT -148.730 -139.550 -144.400 -129.440 ;
        RECT -148.670 -139.600 -148.500 -139.550 ;
        RECT -144.100 -139.940 -143.930 -129.030 ;
        RECT -149.210 -140.110 -143.930 -139.940 ;
        RECT -144.170 -140.120 -143.930 -140.110 ;
        RECT -143.420 -140.870 -142.910 -127.970 ;
        RECT -150.440 -141.380 -142.910 -140.870 ;
        RECT -152.140 -147.400 -150.680 -147.360 ;
        RECT -152.140 -147.570 -150.670 -147.400 ;
        RECT -152.140 -147.610 -150.680 -147.570 ;
        RECT -150.440 -153.990 -149.930 -141.380 ;
        RECT -149.570 -142.170 -143.590 -141.940 ;
        RECT -149.480 -153.230 -143.830 -142.170 ;
        RECT -143.420 -151.740 -142.910 -141.380 ;
        RECT -143.430 -151.760 -142.910 -151.740 ;
        RECT -149.480 -153.240 -143.770 -153.230 ;
        RECT -149.560 -153.410 -143.770 -153.240 ;
        RECT -149.470 -153.420 -143.770 -153.410 ;
        RECT -144.000 -153.490 -143.830 -153.420 ;
        RECT -143.430 -153.540 -142.900 -151.760 ;
        RECT -143.420 -153.560 -142.900 -153.540 ;
        RECT -150.440 -154.280 -148.000 -153.990 ;
        RECT -143.420 -154.070 -142.910 -153.560 ;
        RECT -143.420 -154.280 -142.890 -154.070 ;
        RECT -150.440 -154.760 -142.890 -154.280 ;
        RECT -150.440 -154.790 -143.080 -154.760 ;
        RECT -150.440 -156.550 -142.910 -156.000 ;
        RECT -152.120 -169.520 -150.650 -169.270 ;
        RECT -150.440 -169.460 -149.930 -156.550 ;
        RECT -143.580 -156.560 -142.910 -156.550 ;
        RECT -147.280 -157.450 -143.820 -157.010 ;
        RECT -149.210 -157.550 -143.820 -157.450 ;
        RECT -149.210 -157.620 -143.930 -157.550 ;
        RECT -149.210 -168.530 -149.040 -157.620 ;
        RECT -148.710 -158.030 -144.480 -158.010 ;
        RECT -148.730 -168.140 -144.400 -158.030 ;
        RECT -148.670 -168.190 -148.500 -168.140 ;
        RECT -144.100 -168.530 -143.930 -157.620 ;
        RECT -149.210 -168.700 -143.930 -168.530 ;
        RECT -144.170 -168.710 -143.930 -168.700 ;
        RECT -143.420 -169.460 -142.910 -156.560 ;
        RECT -150.440 -169.970 -142.910 -169.460 ;
        RECT -152.140 -175.990 -150.680 -175.950 ;
        RECT -152.140 -176.160 -150.670 -175.990 ;
        RECT -152.140 -176.200 -150.680 -176.160 ;
        RECT -150.440 -182.580 -149.930 -169.970 ;
        RECT -149.570 -170.760 -143.590 -170.530 ;
        RECT -149.480 -181.820 -143.830 -170.760 ;
        RECT -143.420 -180.330 -142.910 -169.970 ;
        RECT -143.430 -180.350 -142.910 -180.330 ;
        RECT -149.480 -181.830 -143.770 -181.820 ;
        RECT -149.560 -182.000 -143.770 -181.830 ;
        RECT -149.470 -182.010 -143.770 -182.000 ;
        RECT -144.000 -182.080 -143.830 -182.010 ;
        RECT -143.430 -182.130 -142.900 -180.350 ;
        RECT -143.420 -182.150 -142.900 -182.130 ;
        RECT -150.440 -182.870 -148.000 -182.580 ;
        RECT -143.420 -182.660 -142.910 -182.150 ;
        RECT -143.420 -182.870 -142.890 -182.660 ;
        RECT -150.440 -183.350 -142.890 -182.870 ;
        RECT -150.440 -183.380 -143.080 -183.350 ;
        RECT -150.440 -185.140 -142.910 -184.590 ;
        RECT -152.120 -198.110 -150.650 -197.860 ;
        RECT -150.440 -198.050 -149.930 -185.140 ;
        RECT -143.580 -185.150 -142.910 -185.140 ;
        RECT -147.280 -186.040 -143.820 -185.600 ;
        RECT -149.210 -186.140 -143.820 -186.040 ;
        RECT -149.210 -186.210 -143.930 -186.140 ;
        RECT -149.210 -197.120 -149.040 -186.210 ;
        RECT -148.710 -186.620 -144.480 -186.600 ;
        RECT -148.730 -196.730 -144.400 -186.620 ;
        RECT -148.670 -196.780 -148.500 -196.730 ;
        RECT -144.100 -197.120 -143.930 -186.210 ;
        RECT -149.210 -197.290 -143.930 -197.120 ;
        RECT -144.170 -197.300 -143.930 -197.290 ;
        RECT -143.420 -198.050 -142.910 -185.150 ;
        RECT -150.440 -198.560 -142.910 -198.050 ;
        RECT -152.140 -204.580 -150.680 -204.540 ;
        RECT -152.140 -204.750 -150.670 -204.580 ;
        RECT -152.140 -204.790 -150.680 -204.750 ;
        RECT -150.440 -211.170 -149.930 -198.560 ;
        RECT -149.570 -199.350 -143.590 -199.120 ;
        RECT -149.480 -210.410 -143.830 -199.350 ;
        RECT -143.420 -208.920 -142.910 -198.560 ;
        RECT -143.430 -208.940 -142.910 -208.920 ;
        RECT -149.480 -210.420 -143.770 -210.410 ;
        RECT -149.560 -210.590 -143.770 -210.420 ;
        RECT -149.470 -210.600 -143.770 -210.590 ;
        RECT -144.000 -210.670 -143.830 -210.600 ;
        RECT -143.430 -210.720 -142.900 -208.940 ;
        RECT -143.420 -210.740 -142.900 -210.720 ;
        RECT -150.440 -211.460 -148.000 -211.170 ;
        RECT -143.420 -211.250 -142.910 -210.740 ;
        RECT -143.420 -211.460 -142.890 -211.250 ;
        RECT -150.440 -211.940 -142.890 -211.460 ;
        RECT -150.440 -211.970 -143.080 -211.940 ;
        RECT -150.440 -213.730 -142.910 -213.180 ;
        RECT -152.120 -226.700 -150.650 -226.450 ;
        RECT -150.440 -226.640 -149.930 -213.730 ;
        RECT -143.580 -213.740 -142.910 -213.730 ;
        RECT -147.280 -214.630 -143.820 -214.190 ;
        RECT -149.210 -214.730 -143.820 -214.630 ;
        RECT -149.210 -214.800 -143.930 -214.730 ;
        RECT -149.210 -225.710 -149.040 -214.800 ;
        RECT -148.710 -215.210 -144.480 -215.190 ;
        RECT -148.730 -225.320 -144.400 -215.210 ;
        RECT -148.670 -225.370 -148.500 -225.320 ;
        RECT -144.100 -225.710 -143.930 -214.800 ;
        RECT -149.210 -225.880 -143.930 -225.710 ;
        RECT -144.170 -225.890 -143.930 -225.880 ;
        RECT -143.420 -226.640 -142.910 -213.740 ;
        RECT -150.440 -227.150 -142.910 -226.640 ;
        RECT -152.140 -233.170 -150.680 -233.130 ;
        RECT -152.140 -233.340 -150.670 -233.170 ;
        RECT -152.140 -233.380 -150.680 -233.340 ;
        RECT -150.440 -239.760 -149.930 -227.150 ;
        RECT -149.570 -227.940 -143.590 -227.710 ;
        RECT -149.480 -239.000 -143.830 -227.940 ;
        RECT -143.420 -237.510 -142.910 -227.150 ;
        RECT -143.430 -237.530 -142.910 -237.510 ;
        RECT -149.480 -239.010 -143.770 -239.000 ;
        RECT -149.560 -239.180 -143.770 -239.010 ;
        RECT -149.470 -239.190 -143.770 -239.180 ;
        RECT -144.000 -239.260 -143.830 -239.190 ;
        RECT -143.430 -239.310 -142.900 -237.530 ;
        RECT -143.420 -239.330 -142.900 -239.310 ;
        RECT -150.440 -240.050 -148.000 -239.760 ;
        RECT -143.420 -239.840 -142.910 -239.330 ;
        RECT -143.420 -240.050 -142.890 -239.840 ;
        RECT -150.440 -240.530 -142.890 -240.050 ;
        RECT -150.440 -240.560 -143.080 -240.530 ;
      LAYER mcon ;
        RECT -4.380 143.260 -4.210 143.430 ;
        RECT -131.000 143.060 -130.830 143.230 ;
        RECT -131.000 142.720 -130.830 142.890 ;
        RECT -131.000 142.380 -130.830 142.550 ;
        RECT -131.000 142.040 -130.830 142.210 ;
        RECT -124.320 143.040 -124.150 143.210 ;
        RECT -124.320 142.700 -124.150 142.870 ;
        RECT -124.320 142.360 -124.150 142.530 ;
        RECT -124.320 142.020 -124.150 142.190 ;
        RECT -102.410 143.060 -102.240 143.230 ;
        RECT -102.410 142.720 -102.240 142.890 ;
        RECT -102.410 142.380 -102.240 142.550 ;
        RECT -102.410 142.040 -102.240 142.210 ;
        RECT -95.730 143.040 -95.560 143.210 ;
        RECT -95.730 142.700 -95.560 142.870 ;
        RECT -95.730 142.360 -95.560 142.530 ;
        RECT -95.730 142.020 -95.560 142.190 ;
        RECT -73.820 143.060 -73.650 143.230 ;
        RECT -73.820 142.720 -73.650 142.890 ;
        RECT -73.820 142.380 -73.650 142.550 ;
        RECT -73.820 142.040 -73.650 142.210 ;
        RECT -67.140 143.040 -66.970 143.210 ;
        RECT -67.140 142.700 -66.970 142.870 ;
        RECT -4.380 142.920 -4.210 143.090 ;
        RECT -4.380 142.580 -4.210 142.750 ;
        RECT 2.370 143.300 2.540 143.470 ;
        RECT 2.370 142.960 2.540 143.130 ;
        RECT 2.370 142.620 2.540 142.790 ;
        RECT -67.140 142.360 -66.970 142.530 ;
        RECT 10.200 143.060 10.370 143.230 ;
        RECT 10.200 142.720 10.370 142.890 ;
        RECT 10.200 142.380 10.370 142.550 ;
        RECT -67.140 142.020 -66.970 142.190 ;
        RECT 10.200 142.040 10.370 142.210 ;
        RECT 16.880 143.040 17.050 143.210 ;
        RECT 16.880 142.700 17.050 142.870 ;
        RECT 16.880 142.360 17.050 142.530 ;
        RECT 16.880 142.020 17.050 142.190 ;
        RECT 38.790 143.060 38.960 143.230 ;
        RECT 38.790 142.720 38.960 142.890 ;
        RECT 38.790 142.380 38.960 142.550 ;
        RECT -24.830 141.790 -0.930 141.960 ;
        RECT 7.950 141.790 29.120 141.960 ;
        RECT 38.790 142.040 38.960 142.210 ;
        RECT 45.470 143.040 45.640 143.210 ;
        RECT 45.470 142.700 45.640 142.870 ;
        RECT 45.470 142.360 45.640 142.530 ;
        RECT 45.470 142.020 45.640 142.190 ;
        RECT 67.380 143.060 67.550 143.230 ;
        RECT 67.380 142.720 67.550 142.890 ;
        RECT 67.380 142.380 67.550 142.550 ;
        RECT 67.380 142.040 67.550 142.210 ;
        RECT 74.060 143.040 74.230 143.210 ;
        RECT 74.060 142.700 74.230 142.870 ;
        RECT 74.060 142.360 74.230 142.530 ;
        RECT 74.060 142.020 74.230 142.190 ;
        RECT 95.970 143.060 96.140 143.230 ;
        RECT 95.970 142.720 96.140 142.890 ;
        RECT 95.970 142.380 96.140 142.550 ;
        RECT 95.970 142.040 96.140 142.210 ;
        RECT 102.650 143.040 102.820 143.210 ;
        RECT 102.650 142.700 102.820 142.870 ;
        RECT 102.650 142.360 102.820 142.530 ;
        RECT 102.650 142.020 102.820 142.190 ;
        RECT 124.560 143.060 124.730 143.230 ;
        RECT 124.560 142.720 124.730 142.890 ;
        RECT 124.560 142.380 124.730 142.550 ;
        RECT 124.560 142.040 124.730 142.210 ;
        RECT 131.240 143.040 131.410 143.210 ;
        RECT 131.240 142.700 131.410 142.870 ;
        RECT 131.240 142.360 131.410 142.530 ;
        RECT 131.240 142.020 131.410 142.190 ;
        RECT 153.150 143.060 153.320 143.230 ;
        RECT 153.150 142.720 153.320 142.890 ;
        RECT 153.150 142.380 153.320 142.550 ;
        RECT 153.150 142.040 153.320 142.210 ;
        RECT 159.830 143.040 160.000 143.210 ;
        RECT 159.830 142.700 160.000 142.870 ;
        RECT 159.830 142.360 160.000 142.530 ;
        RECT 159.830 142.020 160.000 142.190 ;
        RECT 181.740 143.060 181.910 143.230 ;
        RECT 181.740 142.720 181.910 142.890 ;
        RECT 181.740 142.380 181.910 142.550 ;
        RECT 181.740 142.040 181.910 142.210 ;
        RECT 188.420 143.040 188.590 143.210 ;
        RECT 188.420 142.700 188.590 142.870 ;
        RECT 188.420 142.360 188.590 142.530 ;
        RECT 188.420 142.020 188.590 142.190 ;
        RECT -138.140 141.390 -136.280 141.400 ;
        RECT -138.140 141.220 -136.270 141.390 ;
        RECT -114.780 141.210 -111.620 141.390 ;
        RECT -138.060 140.260 -137.880 141.050 ;
        RECT -138.050 139.130 -137.880 140.260 ;
        RECT -137.700 139.120 -137.520 141.040 ;
        RECT -136.510 140.090 -125.530 140.260 ;
        RECT -136.510 139.470 -125.530 139.640 ;
        RECT -136.500 138.850 -125.520 139.020 ;
        RECT -136.480 138.270 -125.500 138.440 ;
        RECT -136.470 137.680 -125.490 137.850 ;
        RECT -136.470 137.080 -125.490 137.250 ;
        RECT -136.520 136.480 -125.540 136.650 ;
        RECT -136.510 135.870 -125.530 136.040 ;
        RECT -136.520 135.270 -125.540 135.440 ;
        RECT -122.780 139.330 -113.330 139.500 ;
        RECT -122.790 138.580 -113.400 138.750 ;
        RECT -122.760 137.860 -113.360 138.030 ;
        RECT -122.750 137.200 -113.380 137.370 ;
        RECT -122.760 136.550 -113.310 136.720 ;
        RECT -122.750 135.910 -113.360 136.080 ;
        RECT -111.210 140.230 -111.010 141.160 ;
        RECT -112.280 134.990 -111.930 138.290 ;
        RECT -109.550 141.390 -107.690 141.400 ;
        RECT -109.550 141.220 -107.680 141.390 ;
        RECT -86.190 141.210 -83.030 141.390 ;
        RECT -109.470 140.260 -109.290 141.050 ;
        RECT -109.460 139.130 -109.290 140.260 ;
        RECT -109.110 139.120 -108.930 141.040 ;
        RECT -107.920 140.090 -96.940 140.260 ;
        RECT -107.920 139.470 -96.940 139.640 ;
        RECT -107.910 138.850 -96.930 139.020 ;
        RECT -107.890 138.270 -96.910 138.440 ;
        RECT -107.880 137.680 -96.900 137.850 ;
        RECT -107.880 137.080 -96.900 137.250 ;
        RECT -107.930 136.480 -96.950 136.650 ;
        RECT -107.920 135.870 -96.940 136.040 ;
        RECT -107.930 135.270 -96.950 135.440 ;
        RECT -94.190 139.330 -84.740 139.500 ;
        RECT -94.200 138.580 -84.810 138.750 ;
        RECT -94.170 137.860 -84.770 138.030 ;
        RECT -94.160 137.200 -84.790 137.370 ;
        RECT -94.170 136.550 -84.720 136.720 ;
        RECT -94.160 135.910 -84.770 136.080 ;
        RECT -82.620 140.230 -82.420 141.160 ;
        RECT -83.690 134.990 -83.340 138.290 ;
        RECT -80.960 141.390 -79.100 141.400 ;
        RECT -80.960 141.220 -79.090 141.390 ;
        RECT -57.600 141.210 -54.440 141.390 ;
        RECT -80.880 140.260 -80.700 141.050 ;
        RECT -80.870 139.130 -80.700 140.260 ;
        RECT -80.520 139.120 -80.340 141.040 ;
        RECT -79.330 140.090 -68.350 140.260 ;
        RECT -79.330 139.470 -68.350 139.640 ;
        RECT -79.320 138.850 -68.340 139.020 ;
        RECT -79.300 138.270 -68.320 138.440 ;
        RECT -79.290 137.680 -68.310 137.850 ;
        RECT -79.290 137.080 -68.310 137.250 ;
        RECT -79.340 136.480 -68.360 136.650 ;
        RECT -79.330 135.870 -68.350 136.040 ;
        RECT -79.340 135.270 -68.360 135.440 ;
        RECT -65.600 139.330 -56.150 139.500 ;
        RECT -65.610 138.580 -56.220 138.750 ;
        RECT -65.580 137.860 -56.180 138.030 ;
        RECT -65.570 137.200 -56.200 137.370 ;
        RECT -65.580 136.550 -56.130 136.720 ;
        RECT -65.570 135.910 -56.180 136.080 ;
        RECT -54.030 140.230 -53.830 141.160 ;
        RECT -55.100 134.990 -54.750 138.290 ;
        RECT 3.060 141.390 4.920 141.400 ;
        RECT 3.060 141.220 4.930 141.390 ;
        RECT 26.420 141.210 29.580 141.390 ;
        RECT 3.140 140.260 3.320 141.050 ;
        RECT 3.150 139.130 3.320 140.260 ;
        RECT 3.500 139.120 3.680 141.040 ;
        RECT 4.690 140.090 15.670 140.260 ;
        RECT 4.690 139.470 15.670 139.640 ;
        RECT 4.700 138.850 15.680 139.020 ;
        RECT 4.720 138.270 15.700 138.440 ;
        RECT 4.730 137.680 15.710 137.850 ;
        RECT 4.730 137.080 15.710 137.250 ;
        RECT 4.680 136.480 15.660 136.650 ;
        RECT 4.690 135.870 15.670 136.040 ;
        RECT 4.680 135.270 15.660 135.440 ;
        RECT 18.420 139.330 27.870 139.500 ;
        RECT 18.410 138.580 27.800 138.750 ;
        RECT 18.440 137.860 27.840 138.030 ;
        RECT 18.450 137.200 27.820 137.370 ;
        RECT 18.440 136.550 27.890 136.720 ;
        RECT 18.450 135.910 27.840 136.080 ;
        RECT 28.920 134.990 29.270 138.290 ;
        RECT 29.990 140.230 30.190 141.160 ;
        RECT 31.650 141.390 33.510 141.400 ;
        RECT 31.650 141.220 33.520 141.390 ;
        RECT 55.010 141.210 58.170 141.390 ;
        RECT 31.730 140.260 31.910 141.050 ;
        RECT 31.740 139.130 31.910 140.260 ;
        RECT 32.090 139.120 32.270 141.040 ;
        RECT 33.280 140.090 44.260 140.260 ;
        RECT 33.280 139.470 44.260 139.640 ;
        RECT 33.290 138.850 44.270 139.020 ;
        RECT 33.310 138.270 44.290 138.440 ;
        RECT 33.320 137.680 44.300 137.850 ;
        RECT 33.320 137.080 44.300 137.250 ;
        RECT 33.270 136.480 44.250 136.650 ;
        RECT 33.280 135.870 44.260 136.040 ;
        RECT 33.270 135.270 44.250 135.440 ;
        RECT 47.010 139.330 56.460 139.500 ;
        RECT 47.000 138.580 56.390 138.750 ;
        RECT 47.030 137.860 56.430 138.030 ;
        RECT 47.040 137.200 56.410 137.370 ;
        RECT 47.030 136.550 56.480 136.720 ;
        RECT 47.040 135.910 56.430 136.080 ;
        RECT 58.580 140.230 58.780 141.160 ;
        RECT 57.510 134.990 57.860 138.290 ;
        RECT 60.240 141.390 62.100 141.400 ;
        RECT 60.240 141.220 62.110 141.390 ;
        RECT 83.600 141.210 86.760 141.390 ;
        RECT 60.320 140.260 60.500 141.050 ;
        RECT 60.330 139.130 60.500 140.260 ;
        RECT 60.680 139.120 60.860 141.040 ;
        RECT 61.870 140.090 72.850 140.260 ;
        RECT 61.870 139.470 72.850 139.640 ;
        RECT 61.880 138.850 72.860 139.020 ;
        RECT 61.900 138.270 72.880 138.440 ;
        RECT 61.910 137.680 72.890 137.850 ;
        RECT 61.910 137.080 72.890 137.250 ;
        RECT 61.860 136.480 72.840 136.650 ;
        RECT 61.870 135.870 72.850 136.040 ;
        RECT 61.860 135.270 72.840 135.440 ;
        RECT 75.600 139.330 85.050 139.500 ;
        RECT 75.590 138.580 84.980 138.750 ;
        RECT 75.620 137.860 85.020 138.030 ;
        RECT 75.630 137.200 85.000 137.370 ;
        RECT 75.620 136.550 85.070 136.720 ;
        RECT 75.630 135.910 85.020 136.080 ;
        RECT 87.170 140.230 87.370 141.160 ;
        RECT 86.100 134.990 86.450 138.290 ;
        RECT 88.830 141.390 90.690 141.400 ;
        RECT 88.830 141.220 90.700 141.390 ;
        RECT 112.190 141.210 115.350 141.390 ;
        RECT 88.910 140.260 89.090 141.050 ;
        RECT 88.920 139.130 89.090 140.260 ;
        RECT 89.270 139.120 89.450 141.040 ;
        RECT 90.460 140.090 101.440 140.260 ;
        RECT 90.460 139.470 101.440 139.640 ;
        RECT 90.470 138.850 101.450 139.020 ;
        RECT 90.490 138.270 101.470 138.440 ;
        RECT 90.500 137.680 101.480 137.850 ;
        RECT 90.500 137.080 101.480 137.250 ;
        RECT 90.450 136.480 101.430 136.650 ;
        RECT 90.460 135.870 101.440 136.040 ;
        RECT 90.450 135.270 101.430 135.440 ;
        RECT 104.190 139.330 113.640 139.500 ;
        RECT 104.180 138.580 113.570 138.750 ;
        RECT 104.210 137.860 113.610 138.030 ;
        RECT 104.220 137.200 113.590 137.370 ;
        RECT 104.210 136.550 113.660 136.720 ;
        RECT 104.220 135.910 113.610 136.080 ;
        RECT 115.760 140.230 115.960 141.160 ;
        RECT 114.690 134.990 115.040 138.290 ;
        RECT 117.420 141.390 119.280 141.400 ;
        RECT 117.420 141.220 119.290 141.390 ;
        RECT 140.780 141.210 143.940 141.390 ;
        RECT 117.500 140.260 117.680 141.050 ;
        RECT 117.510 139.130 117.680 140.260 ;
        RECT 117.860 139.120 118.040 141.040 ;
        RECT 119.050 140.090 130.030 140.260 ;
        RECT 119.050 139.470 130.030 139.640 ;
        RECT 119.060 138.850 130.040 139.020 ;
        RECT 119.080 138.270 130.060 138.440 ;
        RECT 119.090 137.680 130.070 137.850 ;
        RECT 119.090 137.080 130.070 137.250 ;
        RECT 119.040 136.480 130.020 136.650 ;
        RECT 119.050 135.870 130.030 136.040 ;
        RECT 119.040 135.270 130.020 135.440 ;
        RECT 132.780 139.330 142.230 139.500 ;
        RECT 132.770 138.580 142.160 138.750 ;
        RECT 132.800 137.860 142.200 138.030 ;
        RECT 132.810 137.200 142.180 137.370 ;
        RECT 132.800 136.550 142.250 136.720 ;
        RECT 132.810 135.910 142.200 136.080 ;
        RECT 144.350 140.230 144.550 141.160 ;
        RECT 143.280 134.990 143.630 138.290 ;
        RECT 146.010 141.390 147.870 141.400 ;
        RECT 146.010 141.220 147.880 141.390 ;
        RECT 169.370 141.210 172.530 141.390 ;
        RECT 146.090 140.260 146.270 141.050 ;
        RECT 146.100 139.130 146.270 140.260 ;
        RECT 146.450 139.120 146.630 141.040 ;
        RECT 147.640 140.090 158.620 140.260 ;
        RECT 147.640 139.470 158.620 139.640 ;
        RECT 147.650 138.850 158.630 139.020 ;
        RECT 147.670 138.270 158.650 138.440 ;
        RECT 147.680 137.680 158.660 137.850 ;
        RECT 147.680 137.080 158.660 137.250 ;
        RECT 147.630 136.480 158.610 136.650 ;
        RECT 147.640 135.870 158.620 136.040 ;
        RECT 147.630 135.270 158.610 135.440 ;
        RECT 161.370 139.330 170.820 139.500 ;
        RECT 161.360 138.580 170.750 138.750 ;
        RECT 161.390 137.860 170.790 138.030 ;
        RECT 161.400 137.200 170.770 137.370 ;
        RECT 161.390 136.550 170.840 136.720 ;
        RECT 161.400 135.910 170.790 136.080 ;
        RECT 172.940 140.230 173.140 141.160 ;
        RECT 171.870 134.990 172.220 138.290 ;
        RECT 174.600 141.390 176.460 141.400 ;
        RECT 174.600 141.220 176.470 141.390 ;
        RECT 197.960 141.210 201.120 141.390 ;
        RECT 174.680 140.260 174.860 141.050 ;
        RECT 174.690 139.130 174.860 140.260 ;
        RECT 175.040 139.120 175.220 141.040 ;
        RECT 176.230 140.090 187.210 140.260 ;
        RECT 176.230 139.470 187.210 139.640 ;
        RECT 176.240 138.850 187.220 139.020 ;
        RECT 176.260 138.270 187.240 138.440 ;
        RECT 176.270 137.680 187.250 137.850 ;
        RECT 176.270 137.080 187.250 137.250 ;
        RECT 176.220 136.480 187.200 136.650 ;
        RECT 176.230 135.870 187.210 136.040 ;
        RECT 176.220 135.270 187.200 135.440 ;
        RECT 189.960 139.330 199.410 139.500 ;
        RECT 189.950 138.580 199.340 138.750 ;
        RECT 189.980 137.860 199.380 138.030 ;
        RECT 189.990 137.200 199.360 137.370 ;
        RECT 189.980 136.550 199.430 136.720 ;
        RECT 189.990 135.910 199.380 136.080 ;
        RECT 201.530 140.230 201.730 141.160 ;
        RECT 200.460 134.990 200.810 138.290 ;
        RECT 1.610 133.830 1.780 134.000 ;
        RECT 1.950 133.830 2.120 134.000 ;
        RECT 2.290 133.830 2.460 134.000 ;
        RECT 2.630 133.830 2.800 134.000 ;
        RECT 2.970 133.830 3.140 134.000 ;
        RECT 3.310 133.830 3.480 134.000 ;
        RECT -150.040 129.530 -149.110 129.730 ;
        RECT -150.270 125.960 -150.090 129.120 ;
        RECT -147.170 128.460 -143.870 128.810 ;
        RECT -152.090 116.420 -151.920 116.590 ;
        RECT -151.750 116.420 -151.580 116.590 ;
        RECT -151.410 116.420 -151.240 116.590 ;
        RECT -151.070 116.420 -150.900 116.590 ;
        RECT -148.380 117.960 -148.210 127.410 ;
        RECT -147.630 117.950 -147.460 127.340 ;
        RECT -146.910 117.980 -146.740 127.380 ;
        RECT -146.250 117.990 -146.080 127.360 ;
        RECT -145.600 117.980 -145.430 127.430 ;
        RECT -144.960 117.990 -144.790 127.380 ;
        RECT 212.700 128.810 213.630 129.010 ;
        RECT -23.230 127.310 -23.060 127.480 ;
        RECT -20.360 127.520 -20.190 127.690 ;
        RECT -21.820 127.310 -21.650 127.480 ;
        RECT -5.020 127.340 -4.850 127.510 ;
        RECT -5.020 126.990 -4.850 127.160 ;
        RECT -20.360 126.730 -20.190 126.900 ;
        RECT -5.020 126.650 -4.850 126.820 ;
        RECT 0.840 127.250 1.010 127.420 ;
        RECT 0.840 126.800 1.010 126.970 ;
        RECT 5.540 127.200 5.710 127.370 ;
        RECT 5.540 126.750 5.710 126.920 ;
        RECT -23.230 126.460 -23.060 126.630 ;
        RECT -22.510 126.450 -22.340 126.620 ;
        RECT -21.820 126.460 -21.650 126.630 ;
        RECT -23.050 126.050 -22.880 126.220 ;
        RECT -21.990 126.050 -21.820 126.220 ;
        RECT -23.230 125.640 -23.060 125.810 ;
        RECT -22.510 125.610 -22.340 125.780 ;
        RECT -21.820 125.640 -21.650 125.810 ;
        RECT -7.120 125.710 -6.950 125.880 ;
        RECT -5.760 125.790 -5.590 125.960 ;
        RECT -5.070 125.780 -4.900 125.950 ;
        RECT -20.360 125.300 -20.190 125.470 ;
        RECT -23.230 124.800 -23.060 124.970 ;
        RECT -21.820 124.800 -21.650 124.970 ;
        RECT -21.090 124.540 -20.920 124.710 ;
        RECT -21.100 124.020 -20.930 124.190 ;
        RECT -20.350 123.900 -20.180 124.070 ;
        RECT -23.230 123.680 -23.060 123.850 ;
        RECT -21.820 123.680 -21.650 123.850 ;
        RECT -22.530 122.810 -22.360 122.980 ;
        RECT -21.100 122.830 -20.930 123.000 ;
        RECT -18.340 122.480 -18.170 122.650 ;
        RECT -23.320 122.230 -23.150 122.400 ;
        RECT -22.390 122.230 -22.220 122.400 ;
        RECT -21.690 122.230 -21.520 122.400 ;
        RECT -20.950 122.230 -20.780 122.400 ;
        RECT -20.240 122.220 -20.070 122.390 ;
        RECT -5.020 124.540 -4.850 124.710 ;
        RECT -5.020 124.190 -4.850 124.360 ;
        RECT -5.020 123.850 -4.850 124.020 ;
        RECT 0.840 124.260 1.010 124.430 ;
        RECT 0.840 123.810 1.010 123.980 ;
        RECT 0.840 123.250 1.010 123.420 ;
        RECT -5.020 122.990 -4.850 123.160 ;
        RECT -5.020 122.640 -4.850 122.810 ;
        RECT 0.840 122.800 1.010 122.970 ;
        RECT -5.020 122.300 -4.850 122.470 ;
        RECT 4.760 123.740 4.930 123.910 ;
        RECT -7.840 122.050 -7.670 122.220 ;
        RECT 2.020 122.070 2.190 122.240 ;
        RECT -7.830 117.690 -7.400 118.430 ;
        RECT 13.060 116.130 13.270 116.340 ;
        RECT 17.940 116.240 18.110 116.410 ;
        RECT -152.110 109.740 -151.940 109.910 ;
        RECT -151.770 109.740 -151.600 109.910 ;
        RECT -151.430 109.740 -151.260 109.910 ;
        RECT -151.090 109.740 -150.920 109.910 ;
        RECT -150.270 104.460 -150.100 104.470 ;
        RECT -150.280 102.600 -150.100 104.460 ;
        RECT -149.140 104.230 -148.970 115.210 ;
        RECT -148.520 104.230 -148.350 115.210 ;
        RECT -147.900 104.240 -147.730 115.220 ;
        RECT -147.320 104.260 -147.150 115.240 ;
        RECT -146.730 104.270 -146.560 115.250 ;
        RECT -146.130 104.270 -145.960 115.250 ;
        RECT -145.530 104.220 -145.360 115.200 ;
        RECT -144.920 104.230 -144.750 115.210 ;
        RECT -144.320 104.220 -144.150 115.200 ;
        RECT 11.590 115.760 11.760 115.930 ;
        RECT 18.980 115.890 19.150 116.060 ;
        RECT 18.980 115.540 19.150 115.710 ;
        RECT 207.460 127.740 210.760 128.090 ;
        RECT 208.380 117.270 208.550 126.660 ;
        RECT 209.020 117.260 209.190 126.710 ;
        RECT 209.670 117.270 209.840 126.640 ;
        RECT 210.330 117.260 210.500 126.660 ;
        RECT 211.050 117.230 211.220 126.620 ;
        RECT 211.800 117.240 211.970 126.690 ;
        RECT 213.680 125.240 213.860 128.400 ;
        RECT 13.060 114.580 13.270 114.790 ;
        RECT 17.940 114.690 18.110 114.860 ;
        RECT 11.590 114.210 11.760 114.380 ;
        RECT 18.980 114.340 19.150 114.510 ;
        RECT 40.460 114.530 40.720 115.350 ;
        RECT 52.410 114.560 52.730 115.350 ;
        RECT 214.490 115.700 214.660 115.870 ;
        RECT 214.830 115.700 215.000 115.870 ;
        RECT 215.170 115.700 215.340 115.870 ;
        RECT 215.510 115.700 215.680 115.870 ;
        RECT 54.690 114.890 54.870 115.060 ;
        RECT 55.120 114.870 55.290 115.040 ;
        RECT 52.880 114.590 53.050 114.760 ;
        RECT 18.980 113.990 19.150 114.160 ;
        RECT 53.230 113.750 53.410 113.940 ;
        RECT -9.940 112.810 -9.770 112.980 ;
        RECT -8.850 112.820 -8.680 112.990 ;
        RECT 13.060 113.030 13.270 113.240 ;
        RECT 17.940 113.140 18.110 113.310 ;
        RECT 11.590 112.660 11.760 112.830 ;
        RECT -10.160 112.400 -9.990 112.570 ;
        RECT -8.010 112.350 -7.840 112.520 ;
        RECT 18.980 112.790 19.150 112.960 ;
        RECT 55.590 114.310 55.760 114.480 ;
        RECT 82.750 114.590 82.920 114.760 ;
        RECT 57.830 114.010 58.000 114.180 ;
        RECT 75.910 114.010 76.080 114.180 ;
        RECT 57.830 113.560 58.000 113.730 ;
        RECT 54.310 113.190 54.480 113.360 ;
        RECT 63.280 113.410 63.550 113.680 ;
        RECT 72.250 113.410 72.520 113.680 ;
        RECT 75.910 113.560 76.080 113.730 ;
        RECT 81.080 113.760 81.250 113.930 ;
        RECT 55.120 112.880 55.290 113.050 ;
        RECT 18.980 112.440 19.150 112.610 ;
        RECT -9.940 111.890 -9.770 112.060 ;
        RECT -8.850 111.900 -8.680 112.070 ;
        RECT 82.390 113.750 82.570 113.940 ;
        RECT 60.960 112.300 61.130 112.470 ;
        RECT 74.670 112.300 74.840 112.470 ;
        RECT -10.160 111.480 -9.990 111.650 ;
        RECT 13.060 111.480 13.270 111.690 ;
        RECT 17.940 111.590 18.110 111.760 ;
        RECT -9.940 110.970 -9.770 111.140 ;
        RECT -8.850 110.980 -8.680 111.150 ;
        RECT 11.590 111.110 11.760 111.280 ;
        RECT -10.160 110.560 -9.990 110.730 ;
        RECT 18.980 111.240 19.150 111.410 ;
        RECT 18.980 110.890 19.150 111.060 ;
        RECT 53.230 110.950 53.410 111.140 ;
        RECT 24.560 110.260 24.740 110.430 ;
        RECT -10.130 109.990 -9.960 110.160 ;
        RECT -8.830 109.890 -8.660 110.060 ;
        RECT 22.750 109.960 22.920 110.130 ;
        RECT -10.130 109.030 -9.960 109.200 ;
        RECT 23.100 109.120 23.280 109.310 ;
        RECT -8.830 108.930 -8.660 109.100 ;
        RECT 11.590 108.380 11.760 108.550 ;
        RECT -10.130 108.070 -9.960 108.240 ;
        RECT 18.980 108.600 19.150 108.770 ;
        RECT -8.830 107.970 -8.660 108.140 ;
        RECT 13.060 107.970 13.270 108.180 ;
        RECT 18.980 108.250 19.150 108.420 ;
        RECT 17.940 107.900 18.110 108.070 ;
        RECT 55.590 111.990 55.760 112.160 ;
        RECT 55.130 111.810 55.300 111.980 ;
        RECT 54.300 111.500 54.470 111.670 ;
        RECT 63.280 111.680 63.550 111.950 ;
        RECT 72.250 111.680 72.520 111.950 ;
        RECT 80.690 111.380 80.860 111.550 ;
        RECT 57.830 111.060 58.000 111.230 ;
        RECT 57.830 110.610 58.000 110.780 ;
        RECT 75.910 111.060 76.080 111.230 ;
        RECT 75.910 110.610 76.080 110.780 ;
        RECT 55.580 110.410 55.750 110.580 ;
        RECT 52.630 109.960 52.800 110.130 ;
        RECT 52.880 110.130 53.050 110.300 ;
        RECT 29.590 109.380 29.760 109.550 ;
        RECT 31.680 109.540 31.850 109.710 ;
        RECT 24.420 109.130 24.590 109.300 ;
        RECT 29.590 108.930 29.760 109.100 ;
        RECT 30.750 109.240 30.920 109.410 ;
        RECT 31.590 109.120 31.760 109.290 ;
        RECT 32.340 109.120 32.510 109.290 ;
        RECT 33.150 108.780 33.420 109.050 ;
        RECT 35.320 108.790 35.490 108.960 ;
        RECT 31.030 108.490 31.200 108.660 ;
        RECT 35.720 109.240 35.890 109.410 ;
        RECT 45.790 109.380 45.960 109.550 ;
        RECT 35.720 108.900 35.890 109.070 ;
        RECT 42.130 108.780 42.400 109.050 ;
        RECT 45.790 108.930 45.960 109.100 ;
        RECT 50.960 109.130 51.130 109.300 ;
        RECT -8.430 107.530 -8.260 107.700 ;
        RECT 11.590 106.830 11.760 107.000 ;
        RECT 81.080 111.000 81.250 111.170 ;
        RECT 81.660 111.100 81.830 111.270 ;
        RECT 80.840 110.550 81.010 110.720 ;
        RECT 82.390 110.950 82.570 111.140 ;
        RECT 83.910 111.150 84.080 111.320 ;
        RECT 81.610 110.450 81.780 110.620 ;
        RECT 82.640 110.780 82.810 110.950 ;
        RECT 54.690 109.830 54.870 110.000 ;
        RECT 55.150 109.900 55.320 110.070 ;
        RECT 79.250 110.000 79.420 110.170 ;
        RECT 79.720 110.030 79.890 110.200 ;
        RECT 80.210 109.860 80.380 110.030 ;
        RECT 80.820 110.000 80.990 110.170 ;
        RECT 82.750 110.130 82.920 110.300 ;
        RECT 80.930 109.830 81.110 110.000 ;
        RECT 81.340 109.870 81.510 110.040 ;
        RECT 81.610 109.630 81.780 109.800 ;
        RECT 52.270 109.120 52.450 109.310 ;
        RECT 77.800 109.220 77.970 109.390 ;
        RECT 78.300 109.250 78.470 109.420 ;
        RECT 81.800 109.250 81.970 109.420 ;
        RECT 83.300 109.840 83.470 110.010 ;
        RECT 82.640 109.300 82.810 109.470 ;
        RECT 81.660 108.980 81.830 109.150 ;
        RECT 80.450 108.750 80.620 108.920 ;
        RECT 83.960 108.930 84.130 109.100 ;
        RECT 30.830 107.670 31.000 107.840 ;
        RECT 18.980 107.050 19.150 107.220 ;
        RECT 13.060 106.420 13.270 106.630 ;
        RECT 18.980 106.700 19.150 106.870 ;
        RECT 17.940 106.350 18.110 106.520 ;
        RECT 23.100 106.320 23.280 106.510 ;
        RECT 11.590 105.280 11.760 105.450 ;
        RECT 18.980 105.500 19.150 105.670 ;
        RECT 13.060 104.870 13.270 105.080 ;
        RECT 30.620 107.490 30.790 107.660 ;
        RECT 31.030 107.600 31.200 107.770 ;
        RECT 31.590 106.970 31.760 107.140 ;
        RECT 32.340 106.970 32.510 107.140 ;
        RECT 33.150 107.050 33.420 107.320 ;
        RECT 35.320 107.300 35.490 107.470 ;
        RECT 34.340 106.980 34.510 107.150 ;
        RECT 35.720 107.530 35.890 107.700 ;
        RECT 44.550 107.670 44.720 107.840 ;
        RECT 35.720 107.190 35.890 107.360 ;
        RECT 42.130 107.050 42.400 107.320 ;
        RECT 78.300 108.250 78.470 108.420 ;
        RECT 81.800 108.310 81.970 108.420 ;
        RECT 80.880 107.950 81.050 108.120 ;
        RECT 81.660 108.250 81.970 108.310 ;
        RECT 81.660 108.140 81.830 108.250 ;
        RECT 50.570 106.750 50.740 106.920 ;
        RECT 24.420 106.370 24.590 106.540 ;
        RECT 29.590 106.430 29.760 106.600 ;
        RECT 29.590 105.980 29.760 106.150 ;
        RECT 30.750 106.310 30.920 106.480 ;
        RECT 31.590 106.190 31.760 106.360 ;
        RECT 32.340 106.190 32.510 106.360 ;
        RECT 22.750 105.500 22.920 105.670 ;
        RECT 30.620 105.670 30.790 105.840 ;
        RECT 31.710 105.850 31.880 106.020 ;
        RECT 35.320 105.860 35.490 106.030 ;
        RECT 31.030 105.560 31.200 105.730 ;
        RECT 18.980 105.150 19.150 105.320 ;
        RECT 24.560 105.200 24.740 105.370 ;
        RECT 17.940 104.800 18.110 104.970 ;
        RECT 35.720 106.310 35.890 106.480 ;
        RECT 35.720 105.970 35.890 106.140 ;
        RECT 45.790 106.430 45.960 106.600 ;
        RECT 79.250 107.500 79.420 107.670 ;
        RECT 80.210 107.640 80.380 107.810 ;
        RECT 45.790 105.980 45.960 106.150 ;
        RECT 50.960 106.370 51.130 106.540 ;
        RECT 51.540 106.470 51.710 106.640 ;
        RECT 79.250 106.980 79.420 107.150 ;
        RECT 80.820 107.500 80.990 107.670 ;
        RECT 81.340 107.630 81.510 107.800 ;
        RECT 81.610 107.490 81.780 107.660 ;
        RECT 83.950 108.210 84.120 108.380 ;
        RECT 82.640 107.820 82.810 107.990 ;
        RECT 83.300 107.250 83.470 107.420 ;
        RECT 50.720 105.920 50.890 106.090 ;
        RECT 49.600 105.400 49.770 105.570 ;
        RECT 31.030 104.670 31.200 104.840 ;
        RECT -149.920 103.040 -148.000 103.220 ;
        RECT 11.590 103.730 11.760 103.900 ;
        RECT 18.980 103.950 19.150 104.120 ;
        RECT 13.060 103.320 13.270 103.530 ;
        RECT 31.590 104.040 31.760 104.210 ;
        RECT 32.340 104.040 32.510 104.210 ;
        RECT 34.340 104.050 34.510 104.220 ;
        RECT 34.800 104.200 34.970 104.370 ;
        RECT 18.980 103.600 19.150 103.770 ;
        RECT 35.320 104.370 35.490 104.540 ;
        RECT 35.720 104.600 35.890 104.770 ;
        RECT 35.720 104.260 35.890 104.430 ;
        RECT 40.590 104.200 40.760 104.370 ;
        RECT 34.810 103.510 34.980 103.680 ;
        RECT 17.940 103.250 18.110 103.420 ;
        RECT 40.590 103.520 40.760 103.690 ;
        RECT -149.930 102.690 -148.010 102.860 ;
        RECT 40.010 102.910 40.180 103.080 ;
        RECT -149.930 102.680 -149.140 102.690 ;
        RECT 38.200 102.650 38.370 102.820 ;
        RECT 38.930 102.620 39.100 102.790 ;
        RECT 40.010 102.360 40.180 102.530 ;
        RECT 40.920 102.110 41.090 102.280 ;
        RECT 44.860 102.120 45.030 102.290 ;
        RECT 38.200 101.200 38.370 101.370 ;
        RECT 40.010 101.490 40.180 101.660 ;
        RECT 52.270 106.320 52.450 106.510 ;
        RECT 53.790 106.520 53.960 106.690 ;
        RECT 80.210 106.840 80.380 107.010 ;
        RECT 80.820 106.980 80.990 107.150 ;
        RECT 81.340 106.850 81.510 107.020 ;
        RECT 81.610 106.670 81.780 106.840 ;
        RECT 51.490 105.820 51.660 105.990 ;
        RECT 52.520 106.150 52.690 106.320 ;
        RECT 77.800 106.200 77.970 106.370 ;
        RECT 78.300 106.230 78.470 106.400 ;
        RECT 81.800 106.230 81.970 106.400 ;
        RECT 82.640 106.340 82.810 106.510 ;
        RECT 81.660 106.020 81.830 106.190 ;
        RECT 83.870 105.960 84.040 106.130 ;
        RECT 52.630 105.500 52.800 105.670 ;
        RECT 51.490 105.000 51.660 105.170 ;
        RECT 53.180 105.210 53.350 105.380 ;
        RECT 78.300 105.230 78.470 105.400 ;
        RECT 81.800 105.230 81.970 105.400 ;
        RECT 52.520 104.670 52.690 104.840 ;
        RECT 51.540 104.350 51.710 104.520 ;
        RECT 50.330 104.120 50.500 104.290 ;
        RECT 79.250 104.480 79.420 104.650 ;
        RECT 80.210 104.620 80.380 104.790 ;
        RECT 53.840 104.300 54.010 104.470 ;
        RECT 80.820 104.480 80.990 104.650 ;
        RECT 81.340 104.610 81.510 104.780 ;
        RECT 50.760 103.320 50.930 103.490 ;
        RECT 51.540 103.510 51.710 103.680 ;
        RECT 53.830 103.580 54.000 103.750 ;
        RECT 52.520 103.190 52.690 103.360 ;
        RECT 51.490 102.860 51.660 103.030 ;
        RECT 60.780 102.910 60.950 103.080 ;
        RECT 207.740 103.500 207.910 114.480 ;
        RECT 208.340 103.510 208.510 114.490 ;
        RECT 208.950 103.500 209.120 114.480 ;
        RECT 209.550 103.550 209.720 114.530 ;
        RECT 210.150 103.550 210.320 114.530 ;
        RECT 210.740 103.540 210.910 114.520 ;
        RECT 211.320 103.520 211.490 114.500 ;
        RECT 211.940 103.510 212.110 114.490 ;
        RECT 212.560 103.510 212.730 114.490 ;
        RECT 214.510 109.020 214.680 109.190 ;
        RECT 214.850 109.020 215.020 109.190 ;
        RECT 215.190 109.020 215.360 109.190 ;
        RECT 215.530 109.020 215.700 109.190 ;
        RECT 53.180 102.620 53.350 102.790 ;
        RECT 51.490 102.040 51.660 102.210 ;
        RECT 61.860 102.620 62.030 102.790 ;
        RECT 60.780 102.360 60.950 102.530 ;
        RECT 52.520 101.710 52.690 101.880 ;
        RECT 55.930 102.120 56.100 102.290 ;
        RECT 38.930 101.230 39.100 101.400 ;
        RECT 51.540 101.390 51.710 101.560 ;
        RECT 59.870 102.110 60.040 102.280 ;
        RECT 62.590 102.650 62.760 102.820 ;
        RECT 213.690 103.740 213.860 103.750 ;
        RECT 211.590 102.320 213.510 102.500 ;
        RECT 211.600 101.970 213.520 102.140 ;
        RECT 212.730 101.960 213.520 101.970 ;
        RECT 213.690 101.880 213.870 103.740 ;
        RECT 53.750 101.330 53.920 101.500 ;
        RECT 60.780 101.490 60.950 101.660 ;
        RECT 61.860 101.230 62.030 101.400 ;
        RECT 62.590 101.200 62.760 101.370 ;
        RECT -150.040 100.940 -149.110 101.140 ;
        RECT 40.010 100.940 40.180 101.110 ;
        RECT -150.270 97.370 -150.090 100.530 ;
        RECT -147.170 99.870 -143.870 100.220 ;
        RECT -152.090 87.830 -151.920 88.000 ;
        RECT -151.750 87.830 -151.580 88.000 ;
        RECT -151.410 87.830 -151.240 88.000 ;
        RECT -151.070 87.830 -150.900 88.000 ;
        RECT -148.380 89.370 -148.210 98.820 ;
        RECT -147.630 89.360 -147.460 98.750 ;
        RECT -146.910 89.390 -146.740 98.790 ;
        RECT -146.250 89.400 -146.080 98.770 ;
        RECT -145.600 89.390 -145.430 98.840 ;
        RECT -144.960 89.400 -144.790 98.790 ;
        RECT 40.920 100.520 41.090 100.690 ;
        RECT 44.850 100.660 45.020 100.830 ;
        RECT 60.780 100.940 60.950 101.110 ;
        RECT 40.920 100.180 41.090 100.350 ;
        RECT 43.130 100.290 43.400 100.560 ;
        RECT 44.850 100.320 45.020 100.490 ;
        RECT 40.010 99.900 40.180 100.070 ;
        RECT 47.160 100.360 47.430 100.630 ;
        RECT 53.530 100.360 53.800 100.630 ;
        RECT 55.940 100.660 56.110 100.830 ;
        RECT 55.940 100.320 56.110 100.490 ;
        RECT 57.560 100.290 57.830 100.560 ;
        RECT 59.870 100.520 60.040 100.690 ;
        RECT 62.230 100.420 62.410 100.590 ;
        RECT 59.870 100.180 60.040 100.350 ;
        RECT 212.700 100.220 213.630 100.420 ;
        RECT 60.780 99.900 60.950 100.070 ;
        RECT 38.200 99.640 38.370 99.810 ;
        RECT 30.750 99.170 30.920 99.340 ;
        RECT 31.590 99.050 31.760 99.220 ;
        RECT 32.340 99.050 32.510 99.220 ;
        RECT 11.590 98.250 11.760 98.420 ;
        RECT 18.980 98.470 19.150 98.640 ;
        RECT 13.060 97.840 13.270 98.050 ;
        RECT 18.980 98.120 19.150 98.290 ;
        RECT 35.320 98.720 35.490 98.890 ;
        RECT 31.030 98.420 31.200 98.590 ;
        RECT 35.720 99.170 35.890 99.340 ;
        RECT 38.930 99.610 39.100 99.780 ;
        RECT 61.860 99.610 62.030 99.780 ;
        RECT 40.010 99.350 40.180 99.520 ;
        RECT 60.780 99.350 60.950 99.520 ;
        RECT 62.590 99.640 62.760 99.810 ;
        RECT 35.720 98.830 35.890 99.000 ;
        RECT 38.200 98.200 38.370 98.370 ;
        RECT 40.010 98.490 40.180 98.660 ;
        RECT 60.780 98.490 60.950 98.660 ;
        RECT 38.930 98.230 39.100 98.400 ;
        RECT 61.860 98.230 62.030 98.400 ;
        RECT 62.590 98.200 62.760 98.370 ;
        RECT 17.940 97.770 18.110 97.940 ;
        RECT 40.010 97.940 40.180 98.110 ;
        RECT 60.780 97.940 60.950 98.110 ;
        RECT 31.030 97.530 31.200 97.700 ;
        RECT 11.590 96.700 11.760 96.870 ;
        RECT 35.320 97.230 35.490 97.400 ;
        RECT 18.980 96.920 19.150 97.090 ;
        RECT 13.060 96.290 13.270 96.500 ;
        RECT 31.590 96.900 31.760 97.070 ;
        RECT 32.340 96.900 32.510 97.070 ;
        RECT 34.340 96.910 34.510 97.080 ;
        RECT 35.720 97.460 35.890 97.630 ;
        RECT 35.720 97.120 35.890 97.290 ;
        RECT 18.980 96.570 19.150 96.740 ;
        RECT 17.940 96.220 18.110 96.390 ;
        RECT 30.750 96.240 30.920 96.410 ;
        RECT 31.590 96.120 31.760 96.290 ;
        RECT 32.340 96.120 32.510 96.290 ;
        RECT 11.590 95.150 11.760 95.320 ;
        RECT 18.980 95.370 19.150 95.540 ;
        RECT 13.060 94.740 13.270 94.950 ;
        RECT 35.320 95.790 35.490 95.960 ;
        RECT 31.030 95.490 31.200 95.660 ;
        RECT 35.720 96.240 35.890 96.410 ;
        RECT 35.720 95.900 35.890 96.070 ;
        RECT 18.980 95.020 19.150 95.190 ;
        RECT 17.940 94.670 18.110 94.840 ;
        RECT 31.030 94.600 31.200 94.770 ;
        RECT 35.320 94.300 35.490 94.470 ;
        RECT 11.590 93.600 11.760 93.770 ;
        RECT 18.980 93.820 19.150 93.990 ;
        RECT 31.590 93.970 31.760 94.140 ;
        RECT 32.340 93.970 32.510 94.140 ;
        RECT 34.340 93.980 34.510 94.150 ;
        RECT 35.720 94.530 35.890 94.700 ;
        RECT 35.720 94.190 35.890 94.360 ;
        RECT 13.060 93.190 13.270 93.400 ;
        RECT 18.980 93.470 19.150 93.640 ;
        RECT 17.940 93.120 18.110 93.290 ;
        RECT 27.310 93.090 27.480 93.260 ;
        RECT 25.500 92.830 25.670 93.000 ;
        RECT 26.230 92.800 26.400 92.970 ;
        RECT 27.310 92.540 27.480 92.710 ;
        RECT 28.350 92.270 28.520 92.440 ;
        RECT 25.500 91.380 25.670 91.550 ;
        RECT 32.370 92.300 32.540 92.470 ;
        RECT 27.310 91.670 27.480 91.840 ;
        RECT 26.230 91.410 26.400 91.580 ;
        RECT 27.310 91.120 27.480 91.290 ;
        RECT 28.340 91.090 28.510 91.260 ;
        RECT 28.340 90.750 28.510 90.920 ;
        RECT 32.360 91.030 32.530 91.200 ;
        RECT -11.010 90.340 -10.840 90.510 ;
        RECT -10.360 90.340 -10.190 90.510 ;
        RECT 28.340 90.410 28.510 90.580 ;
        RECT -12.230 89.900 -12.060 90.070 ;
        RECT -11.530 89.900 -11.360 90.070 ;
        RECT -12.680 88.240 -12.510 88.410 ;
        RECT 27.310 90.080 27.480 90.250 ;
        RECT 30.430 90.470 30.700 90.740 ;
        RECT 32.360 90.690 32.530 90.860 ;
        RECT 32.360 90.350 32.530 90.520 ;
        RECT 34.460 90.540 34.730 90.810 ;
        RECT 25.500 89.820 25.670 89.990 ;
        RECT -9.850 89.520 -9.680 89.690 ;
        RECT 26.230 89.790 26.400 89.960 ;
        RECT 27.310 89.530 27.480 89.700 ;
        RECT 30.750 89.410 30.920 89.580 ;
        RECT -9.850 89.180 -9.680 89.350 ;
        RECT 31.590 89.290 31.760 89.460 ;
        RECT 32.340 89.290 32.510 89.460 ;
        RECT 11.590 88.480 11.760 88.650 ;
        RECT 18.980 88.700 19.150 88.870 ;
        RECT -9.680 88.040 -9.510 88.210 ;
        RECT 13.060 88.070 13.270 88.280 ;
        RECT 18.980 88.350 19.150 88.520 ;
        RECT 25.500 88.380 25.670 88.550 ;
        RECT 27.310 88.670 27.480 88.840 ;
        RECT 26.230 88.410 26.400 88.580 ;
        RECT 35.320 88.960 35.490 89.130 ;
        RECT 31.030 88.660 31.200 88.830 ;
        RECT 35.720 89.410 35.890 89.580 ;
        RECT 35.720 89.070 35.890 89.240 ;
        RECT 38.650 89.190 38.820 89.360 ;
        RECT 38.800 88.510 38.970 88.680 ;
        RECT 40.950 88.630 41.120 88.800 ;
        RECT 17.940 88.000 18.110 88.170 ;
        RECT 27.310 88.120 27.480 88.290 ;
        RECT 39.690 88.060 39.860 88.230 ;
        RECT -9.670 87.500 -9.500 87.670 ;
        RECT 31.030 87.770 31.200 87.940 ;
        RECT -152.110 81.150 -151.940 81.320 ;
        RECT -151.770 81.150 -151.600 81.320 ;
        RECT -151.430 81.150 -151.260 81.320 ;
        RECT -151.090 81.150 -150.920 81.320 ;
        RECT -150.270 75.870 -150.100 75.880 ;
        RECT -150.280 74.010 -150.100 75.870 ;
        RECT -149.140 75.640 -148.970 86.620 ;
        RECT -148.520 75.640 -148.350 86.620 ;
        RECT -147.900 75.650 -147.730 86.630 ;
        RECT -147.320 75.670 -147.150 86.650 ;
        RECT -146.730 75.680 -146.560 86.660 ;
        RECT -146.130 75.680 -145.960 86.660 ;
        RECT -145.530 75.630 -145.360 86.610 ;
        RECT -144.920 75.640 -144.750 86.620 ;
        RECT -144.320 75.630 -144.150 86.610 ;
        RECT -12.200 86.020 -12.030 86.190 ;
        RECT 11.590 86.930 11.760 87.100 ;
        RECT 35.320 87.470 35.490 87.640 ;
        RECT -9.860 86.540 -9.690 86.710 ;
        RECT 18.980 87.150 19.150 87.320 ;
        RECT 13.060 86.520 13.270 86.730 ;
        RECT 31.590 87.140 31.760 87.310 ;
        RECT 32.340 87.140 32.510 87.310 ;
        RECT 34.340 87.150 34.510 87.320 ;
        RECT 35.720 87.700 35.890 87.870 ;
        RECT 38.800 87.610 38.970 87.780 ;
        RECT 35.720 87.360 35.890 87.530 ;
        RECT 40.950 87.490 41.120 87.660 ;
        RECT 18.980 86.800 19.150 86.970 ;
        RECT 38.650 86.930 38.820 87.100 ;
        RECT 207.460 99.150 210.760 99.500 ;
        RECT 208.380 88.680 208.550 98.070 ;
        RECT 209.020 88.670 209.190 98.120 ;
        RECT 209.670 88.680 209.840 98.050 ;
        RECT 210.330 88.670 210.500 98.070 ;
        RECT 211.050 88.640 211.220 98.030 ;
        RECT 211.800 88.650 211.970 98.100 ;
        RECT 213.680 96.650 213.860 99.810 ;
        RECT 17.940 86.450 18.110 86.620 ;
        RECT 30.750 86.480 30.920 86.650 ;
        RECT 31.590 86.360 31.760 86.530 ;
        RECT 32.340 86.360 32.510 86.530 ;
        RECT -11.510 86.010 -11.340 86.180 ;
        RECT -11.030 85.240 -10.860 85.410 ;
        RECT 11.590 85.380 11.760 85.550 ;
        RECT -10.320 85.180 -10.150 85.350 ;
        RECT 18.980 85.600 19.150 85.770 ;
        RECT 13.060 84.970 13.270 85.180 ;
        RECT 35.320 86.030 35.490 86.200 ;
        RECT 31.030 85.730 31.200 85.900 ;
        RECT 35.720 86.480 35.890 86.650 ;
        RECT 214.490 87.110 214.660 87.280 ;
        RECT 214.830 87.110 215.000 87.280 ;
        RECT 215.170 87.110 215.340 87.280 ;
        RECT 215.510 87.110 215.680 87.280 ;
        RECT 38.650 86.420 38.820 86.590 ;
        RECT 35.720 86.140 35.890 86.310 ;
        RECT 38.800 85.740 38.970 85.910 ;
        RECT 40.950 85.860 41.120 86.030 ;
        RECT 18.980 85.250 19.150 85.420 ;
        RECT 39.690 85.290 39.860 85.460 ;
        RECT 17.940 84.900 18.110 85.070 ;
        RECT 27.210 84.780 27.380 84.950 ;
        RECT -10.360 84.360 -10.190 84.530 ;
        RECT -13.670 83.920 -13.500 84.090 ;
        RECT -12.570 83.930 -12.400 84.100 ;
        RECT -13.120 83.250 -12.950 83.420 ;
        RECT -13.120 81.880 -12.950 82.050 ;
        RECT -13.670 81.150 -13.500 81.320 ;
        RECT -13.680 79.810 -13.510 79.980 ;
        RECT -11.480 83.930 -11.310 84.100 ;
        RECT -12.020 83.250 -11.850 83.420 ;
        RECT -12.020 81.880 -11.850 82.050 ;
        RECT -12.570 81.150 -12.400 81.320 ;
        RECT -12.570 79.800 -12.400 79.970 ;
        RECT -13.120 79.110 -12.950 79.280 ;
        RECT -10.350 83.890 -10.180 84.060 ;
        RECT 11.590 83.830 11.760 84.000 ;
        RECT 18.980 84.050 19.150 84.220 ;
        RECT -10.920 83.250 -10.750 83.420 ;
        RECT 13.060 83.420 13.270 83.630 ;
        RECT 31.030 84.840 31.200 85.010 ;
        RECT 35.320 84.540 35.490 84.710 ;
        RECT 27.260 83.930 27.430 84.100 ;
        RECT 31.590 84.210 31.760 84.380 ;
        RECT 32.340 84.210 32.510 84.380 ;
        RECT 34.340 84.220 34.510 84.390 ;
        RECT 35.720 84.770 35.890 84.940 ;
        RECT 38.800 84.840 38.970 85.010 ;
        RECT 35.720 84.430 35.890 84.600 ;
        RECT 40.950 84.720 41.120 84.890 ;
        RECT 38.650 84.160 38.820 84.330 ;
        RECT 18.980 83.700 19.150 83.870 ;
        RECT -10.230 83.230 -10.060 83.400 ;
        RECT 17.940 83.350 18.110 83.520 ;
        RECT -10.230 82.890 -10.060 83.060 ;
        RECT -10.230 82.550 -10.060 82.720 ;
        RECT -10.920 81.880 -10.750 82.050 ;
        RECT -11.480 81.150 -11.310 81.320 ;
        RECT -11.480 79.780 -11.310 79.950 ;
        RECT -12.020 79.100 -11.850 79.270 ;
        RECT -3.650 79.980 -3.480 80.320 ;
        RECT -3.310 79.980 -3.140 80.320 ;
        RECT -10.930 79.100 -10.760 79.270 ;
        RECT -10.320 76.800 -10.150 76.970 ;
        RECT -13.630 76.360 -13.460 76.530 ;
        RECT -12.530 76.370 -12.360 76.540 ;
        RECT -11.440 76.370 -11.270 76.540 ;
        RECT -13.080 75.690 -12.910 75.860 ;
        RECT -11.980 75.690 -11.810 75.860 ;
        RECT -149.920 74.450 -148.000 74.630 ;
        RECT -13.080 74.320 -12.910 74.490 ;
        RECT -11.980 74.320 -11.810 74.490 ;
        RECT -149.930 74.100 -148.010 74.270 ;
        RECT -149.930 74.090 -149.140 74.100 ;
        RECT -10.310 76.330 -10.140 76.500 ;
        RECT -10.880 75.690 -10.710 75.860 ;
        RECT -10.880 74.320 -10.710 74.490 ;
        RECT 19.280 77.640 19.450 77.810 ;
        RECT 20.370 77.640 20.540 77.810 ;
        RECT 19.830 76.960 20.000 77.130 ;
        RECT 19.830 75.590 20.000 75.760 ;
        RECT 22.590 77.810 22.760 77.980 ;
        RECT 21.470 77.630 21.640 77.800 ;
        RECT 22.590 77.470 22.760 77.640 ;
        RECT 24.480 77.810 24.650 77.980 ;
        RECT 24.480 77.470 24.650 77.640 ;
        RECT 25.600 77.630 25.770 77.800 ;
        RECT 26.700 77.640 26.870 77.810 ;
        RECT 20.920 76.940 21.090 77.110 ;
        RECT 22.030 76.930 22.200 77.100 ;
        RECT 25.040 76.930 25.210 77.100 ;
        RECT 26.150 76.940 26.320 77.110 ;
        RECT 20.920 75.590 21.090 75.760 ;
        RECT 22.020 75.590 22.190 75.760 ;
        RECT 25.050 75.590 25.220 75.760 ;
        RECT 26.150 75.590 26.320 75.760 ;
        RECT 27.790 77.640 27.960 77.810 ;
        RECT 27.240 76.960 27.410 77.130 ;
        RECT 27.240 75.590 27.410 75.760 ;
        RECT 29.090 77.670 29.260 77.840 ;
        RECT 30.180 77.670 30.350 77.840 ;
        RECT 29.640 76.990 29.810 77.160 ;
        RECT 29.640 75.620 29.810 75.790 ;
        RECT 32.400 77.840 32.570 78.010 ;
        RECT 31.280 77.660 31.450 77.830 ;
        RECT 32.400 77.500 32.570 77.670 ;
        RECT 34.290 77.840 34.460 78.010 ;
        RECT 34.290 77.500 34.460 77.670 ;
        RECT 35.410 77.660 35.580 77.830 ;
        RECT 36.510 77.670 36.680 77.840 ;
        RECT 30.730 76.970 30.900 77.140 ;
        RECT 31.840 76.960 32.010 77.130 ;
        RECT 34.850 76.960 35.020 77.130 ;
        RECT 35.960 76.970 36.130 77.140 ;
        RECT 30.730 75.620 30.900 75.790 ;
        RECT 31.830 75.620 32.000 75.790 ;
        RECT 34.860 75.620 35.030 75.790 ;
        RECT 35.960 75.620 36.130 75.790 ;
        RECT 37.600 77.670 37.770 77.840 ;
        RECT 37.050 76.990 37.220 77.160 ;
        RECT 37.050 75.620 37.220 75.790 ;
        RECT 41.150 77.640 41.320 77.810 ;
        RECT 40.590 76.940 40.760 77.110 ;
        RECT 40.600 75.600 40.770 75.770 ;
        RECT -13.630 73.590 -13.460 73.760 ;
        RECT -12.530 73.590 -12.360 73.760 ;
        RECT -150.040 72.350 -149.110 72.550 ;
        RECT -13.640 72.250 -13.470 72.420 ;
        RECT -12.530 72.240 -12.360 72.410 ;
        RECT -150.270 68.780 -150.090 71.940 ;
        RECT -147.170 71.280 -143.870 71.630 ;
        RECT -152.090 59.240 -151.920 59.410 ;
        RECT -151.750 59.240 -151.580 59.410 ;
        RECT -151.410 59.240 -151.240 59.410 ;
        RECT -151.070 59.240 -150.900 59.410 ;
        RECT -148.380 60.780 -148.210 70.230 ;
        RECT -147.630 60.770 -147.460 70.160 ;
        RECT -146.910 60.800 -146.740 70.200 ;
        RECT -146.250 60.810 -146.080 70.180 ;
        RECT -145.600 60.800 -145.430 70.250 ;
        RECT -144.960 60.810 -144.790 70.200 ;
        RECT -14.200 71.710 -14.030 71.880 ;
        RECT -13.080 71.550 -12.910 71.720 ;
        RECT -11.440 73.590 -11.270 73.760 ;
        RECT -11.440 72.220 -11.270 72.390 ;
        RECT -11.980 71.540 -11.810 71.710 ;
        RECT -10.890 71.540 -10.720 71.710 ;
        RECT 19.270 74.860 19.440 75.030 ;
        RECT 19.270 73.490 19.440 73.660 ;
        RECT 18.700 72.850 18.870 73.020 ;
        RECT 20.370 74.860 20.540 75.030 ;
        RECT 21.470 74.860 21.640 75.030 ;
        RECT 25.600 74.860 25.770 75.030 ;
        RECT 26.700 74.860 26.870 75.030 ;
        RECT 20.370 73.490 20.540 73.660 ;
        RECT 21.470 73.490 21.640 73.660 ;
        RECT 25.600 73.490 25.770 73.660 ;
        RECT 26.700 73.490 26.870 73.660 ;
        RECT 19.830 72.810 20.000 72.980 ;
        RECT 20.920 72.810 21.090 72.980 ;
        RECT 22.020 72.820 22.190 72.990 ;
        RECT 25.050 72.820 25.220 72.990 ;
        RECT 26.150 72.810 26.320 72.980 ;
        RECT 27.800 74.860 27.970 75.030 ;
        RECT 27.800 73.490 27.970 73.660 ;
        RECT 27.240 72.810 27.410 72.980 ;
        RECT 29.080 74.890 29.250 75.060 ;
        RECT 29.080 73.520 29.250 73.690 ;
        RECT 28.510 73.020 28.680 73.050 ;
        RECT 28.370 72.880 28.680 73.020 ;
        RECT 28.370 72.850 28.540 72.880 ;
        RECT 30.180 74.890 30.350 75.060 ;
        RECT 31.280 74.890 31.450 75.060 ;
        RECT 35.410 74.890 35.580 75.060 ;
        RECT 36.510 74.890 36.680 75.060 ;
        RECT 30.180 73.520 30.350 73.690 ;
        RECT 31.280 73.520 31.450 73.690 ;
        RECT 35.410 73.520 35.580 73.690 ;
        RECT 36.510 73.520 36.680 73.690 ;
        RECT 18.710 72.380 18.880 72.550 ;
        RECT 29.640 72.840 29.810 73.010 ;
        RECT 30.730 72.840 30.900 73.010 ;
        RECT 31.830 72.850 32.000 73.020 ;
        RECT 34.860 72.850 35.030 73.020 ;
        RECT 35.960 72.840 36.130 73.010 ;
        RECT 37.610 74.890 37.780 75.060 ;
        RECT 37.610 73.520 37.780 73.690 ;
        RECT 37.050 72.840 37.220 73.010 ;
        RECT 38.180 72.880 38.350 73.050 ;
        RECT 42.250 77.650 42.420 77.820 ;
        RECT 41.700 76.950 41.870 77.120 ;
        RECT 41.700 75.600 41.870 75.770 ;
        RECT 41.150 74.870 41.320 75.040 ;
        RECT 41.150 73.500 41.320 73.670 ;
        RECT 28.520 72.550 28.690 72.580 ;
        RECT 28.360 72.410 28.690 72.550 ;
        RECT 28.360 72.380 28.530 72.410 ;
        RECT 40.600 72.830 40.770 73.000 ;
        RECT 43.340 77.650 43.510 77.820 ;
        RECT 42.790 76.970 42.960 77.140 ;
        RECT 42.790 75.600 42.960 75.770 ;
        RECT 42.250 74.870 42.420 75.040 ;
        RECT 42.250 73.500 42.420 73.670 ;
        RECT 41.700 72.820 41.870 72.990 ;
        RECT 43.350 74.870 43.520 75.040 ;
        RECT 44.040 74.540 44.210 74.710 ;
        RECT 44.040 74.200 44.210 74.370 ;
        RECT 44.040 73.860 44.210 74.030 ;
        RECT 43.350 73.500 43.520 73.670 ;
        RECT 42.790 72.820 42.960 72.990 ;
        RECT 43.920 72.860 44.090 73.030 ;
        RECT 38.170 72.410 38.340 72.580 ;
        RECT 43.910 72.390 44.080 72.560 ;
        RECT -9.490 68.010 -9.320 71.530 ;
        RECT -9.120 68.010 -8.950 71.530 ;
        RECT -8.770 68.010 -8.600 71.530 ;
        RECT -8.430 68.010 -8.260 71.530 ;
        RECT -8.080 68.010 -7.910 71.530 ;
        RECT -7.720 68.010 -7.550 71.530 ;
        RECT -7.360 68.010 -7.190 71.530 ;
        RECT 69.280 70.240 69.450 70.410 ;
        RECT 74.800 69.500 74.970 69.670 ;
        RECT 69.280 68.630 69.450 68.800 ;
        RECT 74.800 68.830 74.970 69.000 ;
        RECT 69.280 67.030 69.450 67.200 ;
        RECT 69.280 65.410 69.450 65.580 ;
        RECT 71.810 64.200 71.980 64.370 ;
        RECT 69.280 63.810 69.450 63.980 ;
        RECT 69.280 62.190 69.450 62.360 ;
        RECT 69.280 60.590 69.450 60.760 ;
        RECT 80.880 60.800 81.050 75.750 ;
        RECT 207.740 74.910 207.910 85.890 ;
        RECT 208.340 74.920 208.510 85.900 ;
        RECT 208.950 74.910 209.120 85.890 ;
        RECT 209.550 74.960 209.720 85.940 ;
        RECT 210.150 74.960 210.320 85.940 ;
        RECT 210.740 74.950 210.910 85.930 ;
        RECT 211.320 74.930 211.490 85.910 ;
        RECT 211.940 74.920 212.110 85.900 ;
        RECT 212.560 74.920 212.730 85.900 ;
        RECT 214.510 80.430 214.680 80.600 ;
        RECT 214.850 80.430 215.020 80.600 ;
        RECT 215.190 80.430 215.360 80.600 ;
        RECT 215.530 80.430 215.700 80.600 ;
        RECT 213.690 75.150 213.860 75.160 ;
        RECT 211.590 73.730 213.510 73.910 ;
        RECT 211.600 73.380 213.520 73.550 ;
        RECT 212.730 73.370 213.520 73.380 ;
        RECT 213.690 73.290 213.870 75.150 ;
        RECT 212.700 71.630 213.630 71.830 ;
        RECT 69.280 58.970 69.450 59.140 ;
        RECT -152.110 52.560 -151.940 52.730 ;
        RECT -151.770 52.560 -151.600 52.730 ;
        RECT -151.430 52.560 -151.260 52.730 ;
        RECT -151.090 52.560 -150.920 52.730 ;
        RECT -150.270 47.280 -150.100 47.290 ;
        RECT -150.280 45.420 -150.100 47.280 ;
        RECT -149.140 47.050 -148.970 58.030 ;
        RECT -148.520 47.050 -148.350 58.030 ;
        RECT -147.900 47.060 -147.730 58.040 ;
        RECT -147.320 47.080 -147.150 58.060 ;
        RECT -146.730 47.090 -146.560 58.070 ;
        RECT -146.130 47.090 -145.960 58.070 ;
        RECT -145.530 47.040 -145.360 58.020 ;
        RECT -144.920 47.050 -144.750 58.030 ;
        RECT -144.320 47.040 -144.150 58.020 ;
        RECT 207.460 70.560 210.760 70.910 ;
        RECT 208.380 60.090 208.550 69.480 ;
        RECT 209.020 60.080 209.190 69.530 ;
        RECT 209.670 60.090 209.840 69.460 ;
        RECT 210.330 60.080 210.500 69.480 ;
        RECT 211.050 60.050 211.220 69.440 ;
        RECT 211.800 60.060 211.970 69.510 ;
        RECT 213.680 68.060 213.860 71.220 ;
        RECT 214.490 58.520 214.660 58.690 ;
        RECT 214.830 58.520 215.000 58.690 ;
        RECT 215.170 58.520 215.340 58.690 ;
        RECT 215.510 58.520 215.680 58.690 ;
        RECT -149.920 45.860 -148.000 46.040 ;
        RECT 207.740 46.320 207.910 57.300 ;
        RECT 208.340 46.330 208.510 57.310 ;
        RECT 208.950 46.320 209.120 57.300 ;
        RECT 209.550 46.370 209.720 57.350 ;
        RECT 210.150 46.370 210.320 57.350 ;
        RECT 210.740 46.360 210.910 57.340 ;
        RECT 211.320 46.340 211.490 57.320 ;
        RECT 211.940 46.330 212.110 57.310 ;
        RECT 212.560 46.330 212.730 57.310 ;
        RECT 214.510 51.840 214.680 52.010 ;
        RECT 214.850 51.840 215.020 52.010 ;
        RECT 215.190 51.840 215.360 52.010 ;
        RECT 215.530 51.840 215.700 52.010 ;
        RECT -149.930 45.510 -148.010 45.680 ;
        RECT -149.930 45.500 -149.140 45.510 ;
        RECT 213.690 46.560 213.860 46.570 ;
        RECT 211.590 45.140 213.510 45.320 ;
        RECT 211.600 44.790 213.520 44.960 ;
        RECT 212.730 44.780 213.520 44.790 ;
        RECT 213.690 44.700 213.870 46.560 ;
        RECT -150.040 43.760 -149.110 43.960 ;
        RECT -150.270 40.190 -150.090 43.350 ;
        RECT -147.170 42.690 -143.870 43.040 ;
        RECT -152.090 30.650 -151.920 30.820 ;
        RECT -151.750 30.650 -151.580 30.820 ;
        RECT -151.410 30.650 -151.240 30.820 ;
        RECT -151.070 30.650 -150.900 30.820 ;
        RECT -148.380 32.190 -148.210 41.640 ;
        RECT -147.630 32.180 -147.460 41.570 ;
        RECT -146.910 32.210 -146.740 41.610 ;
        RECT -146.250 32.220 -146.080 41.590 ;
        RECT -145.600 32.210 -145.430 41.660 ;
        RECT -144.960 32.220 -144.790 41.610 ;
        RECT -152.110 23.970 -151.940 24.140 ;
        RECT -151.770 23.970 -151.600 24.140 ;
        RECT -151.430 23.970 -151.260 24.140 ;
        RECT -151.090 23.970 -150.920 24.140 ;
        RECT -150.270 18.690 -150.100 18.700 ;
        RECT -150.280 16.830 -150.100 18.690 ;
        RECT -149.140 18.460 -148.970 29.440 ;
        RECT -148.520 18.460 -148.350 29.440 ;
        RECT -147.900 18.470 -147.730 29.450 ;
        RECT -147.320 18.490 -147.150 29.470 ;
        RECT -146.730 18.500 -146.560 29.480 ;
        RECT -146.130 18.500 -145.960 29.480 ;
        RECT -145.530 18.450 -145.360 29.430 ;
        RECT -144.920 18.460 -144.750 29.440 ;
        RECT -144.320 18.450 -144.150 29.430 ;
        RECT 212.700 43.040 213.630 43.240 ;
        RECT 207.460 41.970 210.760 42.320 ;
        RECT 208.380 31.500 208.550 40.890 ;
        RECT 209.020 31.490 209.190 40.940 ;
        RECT 209.670 31.500 209.840 40.870 ;
        RECT 210.330 31.490 210.500 40.890 ;
        RECT 211.050 31.460 211.220 40.850 ;
        RECT 211.800 31.470 211.970 40.920 ;
        RECT 213.680 39.470 213.860 42.630 ;
        RECT 214.490 29.930 214.660 30.100 ;
        RECT 214.830 29.930 215.000 30.100 ;
        RECT 215.170 29.930 215.340 30.100 ;
        RECT 215.510 29.930 215.680 30.100 ;
        RECT -149.920 17.270 -148.000 17.450 ;
        RECT 207.740 17.730 207.910 28.710 ;
        RECT 208.340 17.740 208.510 28.720 ;
        RECT 208.950 17.730 209.120 28.710 ;
        RECT 209.550 17.780 209.720 28.760 ;
        RECT 210.150 17.780 210.320 28.760 ;
        RECT 210.740 17.770 210.910 28.750 ;
        RECT 211.320 17.750 211.490 28.730 ;
        RECT 211.940 17.740 212.110 28.720 ;
        RECT 212.560 17.740 212.730 28.720 ;
        RECT 214.510 23.250 214.680 23.420 ;
        RECT 214.850 23.250 215.020 23.420 ;
        RECT 215.190 23.250 215.360 23.420 ;
        RECT 215.530 23.250 215.700 23.420 ;
        RECT -149.930 16.920 -148.010 17.090 ;
        RECT -149.930 16.910 -149.140 16.920 ;
        RECT 213.690 17.970 213.860 17.980 ;
        RECT 211.590 16.550 213.510 16.730 ;
        RECT 211.600 16.200 213.520 16.370 ;
        RECT 212.730 16.190 213.520 16.200 ;
        RECT 213.690 16.110 213.870 17.970 ;
        RECT -150.040 15.170 -149.110 15.370 ;
        RECT -150.270 11.600 -150.090 14.760 ;
        RECT -147.170 14.100 -143.870 14.450 ;
        RECT -152.090 2.060 -151.920 2.230 ;
        RECT -151.750 2.060 -151.580 2.230 ;
        RECT -151.410 2.060 -151.240 2.230 ;
        RECT -151.070 2.060 -150.900 2.230 ;
        RECT -148.380 3.600 -148.210 13.050 ;
        RECT -147.630 3.590 -147.460 12.980 ;
        RECT -146.910 3.620 -146.740 13.020 ;
        RECT -146.250 3.630 -146.080 13.000 ;
        RECT -145.600 3.620 -145.430 13.070 ;
        RECT -144.960 3.630 -144.790 13.020 ;
        RECT -152.110 -4.620 -151.940 -4.450 ;
        RECT -151.770 -4.620 -151.600 -4.450 ;
        RECT -151.430 -4.620 -151.260 -4.450 ;
        RECT -151.090 -4.620 -150.920 -4.450 ;
        RECT -150.270 -9.900 -150.100 -9.890 ;
        RECT -150.280 -11.760 -150.100 -9.900 ;
        RECT -149.140 -10.130 -148.970 0.850 ;
        RECT -148.520 -10.130 -148.350 0.850 ;
        RECT -147.900 -10.120 -147.730 0.860 ;
        RECT -147.320 -10.100 -147.150 0.880 ;
        RECT -146.730 -10.090 -146.560 0.890 ;
        RECT -146.130 -10.090 -145.960 0.890 ;
        RECT -145.530 -10.140 -145.360 0.840 ;
        RECT -144.920 -10.130 -144.750 0.850 ;
        RECT -144.320 -10.140 -144.150 0.840 ;
        RECT 212.700 14.450 213.630 14.650 ;
        RECT 207.460 13.380 210.760 13.730 ;
        RECT 208.380 2.910 208.550 12.300 ;
        RECT 209.020 2.900 209.190 12.350 ;
        RECT 209.670 2.910 209.840 12.280 ;
        RECT 210.330 2.900 210.500 12.300 ;
        RECT 211.050 2.870 211.220 12.260 ;
        RECT 211.800 2.880 211.970 12.330 ;
        RECT 213.680 10.880 213.860 14.040 ;
        RECT 214.490 1.340 214.660 1.510 ;
        RECT 214.830 1.340 215.000 1.510 ;
        RECT 215.170 1.340 215.340 1.510 ;
        RECT 215.510 1.340 215.680 1.510 ;
        RECT -149.920 -11.320 -148.000 -11.140 ;
        RECT 207.740 -10.860 207.910 0.120 ;
        RECT 208.340 -10.850 208.510 0.130 ;
        RECT 208.950 -10.860 209.120 0.120 ;
        RECT 209.550 -10.810 209.720 0.170 ;
        RECT 210.150 -10.810 210.320 0.170 ;
        RECT 210.740 -10.820 210.910 0.160 ;
        RECT 211.320 -10.840 211.490 0.140 ;
        RECT 211.940 -10.850 212.110 0.130 ;
        RECT 212.560 -10.850 212.730 0.130 ;
        RECT 214.510 -5.340 214.680 -5.170 ;
        RECT 214.850 -5.340 215.020 -5.170 ;
        RECT 215.190 -5.340 215.360 -5.170 ;
        RECT 215.530 -5.340 215.700 -5.170 ;
        RECT -149.930 -11.670 -148.010 -11.500 ;
        RECT -149.930 -11.680 -149.140 -11.670 ;
        RECT 213.690 -10.620 213.860 -10.610 ;
        RECT 211.590 -12.040 213.510 -11.860 ;
        RECT 211.600 -12.390 213.520 -12.220 ;
        RECT 212.730 -12.400 213.520 -12.390 ;
        RECT 213.690 -12.480 213.870 -10.620 ;
        RECT -150.040 -13.420 -149.110 -13.220 ;
        RECT -150.270 -16.990 -150.090 -13.830 ;
        RECT -147.170 -14.490 -143.870 -14.140 ;
        RECT -152.090 -26.530 -151.920 -26.360 ;
        RECT -151.750 -26.530 -151.580 -26.360 ;
        RECT -151.410 -26.530 -151.240 -26.360 ;
        RECT -151.070 -26.530 -150.900 -26.360 ;
        RECT -148.380 -24.990 -148.210 -15.540 ;
        RECT -147.630 -25.000 -147.460 -15.610 ;
        RECT -146.910 -24.970 -146.740 -15.570 ;
        RECT -146.250 -24.960 -146.080 -15.590 ;
        RECT -145.600 -24.970 -145.430 -15.520 ;
        RECT -144.960 -24.960 -144.790 -15.570 ;
        RECT -152.110 -33.210 -151.940 -33.040 ;
        RECT -151.770 -33.210 -151.600 -33.040 ;
        RECT -151.430 -33.210 -151.260 -33.040 ;
        RECT -151.090 -33.210 -150.920 -33.040 ;
        RECT -150.270 -38.490 -150.100 -38.480 ;
        RECT -150.280 -40.350 -150.100 -38.490 ;
        RECT -149.140 -38.720 -148.970 -27.740 ;
        RECT -148.520 -38.720 -148.350 -27.740 ;
        RECT -147.900 -38.710 -147.730 -27.730 ;
        RECT -147.320 -38.690 -147.150 -27.710 ;
        RECT -146.730 -38.680 -146.560 -27.700 ;
        RECT -146.130 -38.680 -145.960 -27.700 ;
        RECT -145.530 -38.730 -145.360 -27.750 ;
        RECT -144.920 -38.720 -144.750 -27.740 ;
        RECT -144.320 -38.730 -144.150 -27.750 ;
        RECT 212.700 -14.140 213.630 -13.940 ;
        RECT 207.460 -15.210 210.760 -14.860 ;
        RECT 208.380 -25.680 208.550 -16.290 ;
        RECT 209.020 -25.690 209.190 -16.240 ;
        RECT 209.670 -25.680 209.840 -16.310 ;
        RECT 210.330 -25.690 210.500 -16.290 ;
        RECT 211.050 -25.720 211.220 -16.330 ;
        RECT 211.800 -25.710 211.970 -16.260 ;
        RECT 213.680 -17.710 213.860 -14.550 ;
        RECT 214.490 -27.250 214.660 -27.080 ;
        RECT 214.830 -27.250 215.000 -27.080 ;
        RECT 215.170 -27.250 215.340 -27.080 ;
        RECT 215.510 -27.250 215.680 -27.080 ;
        RECT -149.920 -39.910 -148.000 -39.730 ;
        RECT 207.740 -39.450 207.910 -28.470 ;
        RECT 208.340 -39.440 208.510 -28.460 ;
        RECT 208.950 -39.450 209.120 -28.470 ;
        RECT 209.550 -39.400 209.720 -28.420 ;
        RECT 210.150 -39.400 210.320 -28.420 ;
        RECT 210.740 -39.410 210.910 -28.430 ;
        RECT 211.320 -39.430 211.490 -28.450 ;
        RECT 211.940 -39.440 212.110 -28.460 ;
        RECT 212.560 -39.440 212.730 -28.460 ;
        RECT 214.510 -33.930 214.680 -33.760 ;
        RECT 214.850 -33.930 215.020 -33.760 ;
        RECT 215.190 -33.930 215.360 -33.760 ;
        RECT 215.530 -33.930 215.700 -33.760 ;
        RECT -149.930 -40.260 -148.010 -40.090 ;
        RECT -149.930 -40.270 -149.140 -40.260 ;
        RECT 213.690 -39.210 213.860 -39.200 ;
        RECT 211.590 -40.630 213.510 -40.450 ;
        RECT 211.600 -40.980 213.520 -40.810 ;
        RECT 212.730 -40.990 213.520 -40.980 ;
        RECT 213.690 -41.070 213.870 -39.210 ;
        RECT -150.040 -42.010 -149.110 -41.810 ;
        RECT -150.270 -45.580 -150.090 -42.420 ;
        RECT -147.170 -43.080 -143.870 -42.730 ;
        RECT -152.090 -55.120 -151.920 -54.950 ;
        RECT -151.750 -55.120 -151.580 -54.950 ;
        RECT -151.410 -55.120 -151.240 -54.950 ;
        RECT -151.070 -55.120 -150.900 -54.950 ;
        RECT -148.380 -53.580 -148.210 -44.130 ;
        RECT -147.630 -53.590 -147.460 -44.200 ;
        RECT -146.910 -53.560 -146.740 -44.160 ;
        RECT -146.250 -53.550 -146.080 -44.180 ;
        RECT -145.600 -53.560 -145.430 -44.110 ;
        RECT -144.960 -53.550 -144.790 -44.160 ;
        RECT -152.110 -61.800 -151.940 -61.630 ;
        RECT -151.770 -61.800 -151.600 -61.630 ;
        RECT -151.430 -61.800 -151.260 -61.630 ;
        RECT -151.090 -61.800 -150.920 -61.630 ;
        RECT -150.270 -67.080 -150.100 -67.070 ;
        RECT -150.280 -68.940 -150.100 -67.080 ;
        RECT -149.140 -67.310 -148.970 -56.330 ;
        RECT -148.520 -67.310 -148.350 -56.330 ;
        RECT -147.900 -67.300 -147.730 -56.320 ;
        RECT -147.320 -67.280 -147.150 -56.300 ;
        RECT -146.730 -67.270 -146.560 -56.290 ;
        RECT -146.130 -67.270 -145.960 -56.290 ;
        RECT -145.530 -67.320 -145.360 -56.340 ;
        RECT -144.920 -67.310 -144.750 -56.330 ;
        RECT -144.320 -67.320 -144.150 -56.340 ;
        RECT 212.700 -42.730 213.630 -42.530 ;
        RECT 207.460 -43.800 210.760 -43.450 ;
        RECT 208.380 -54.270 208.550 -44.880 ;
        RECT 209.020 -54.280 209.190 -44.830 ;
        RECT 209.670 -54.270 209.840 -44.900 ;
        RECT 210.330 -54.280 210.500 -44.880 ;
        RECT 211.050 -54.310 211.220 -44.920 ;
        RECT 211.800 -54.300 211.970 -44.850 ;
        RECT 213.680 -46.300 213.860 -43.140 ;
        RECT 214.490 -55.840 214.660 -55.670 ;
        RECT 214.830 -55.840 215.000 -55.670 ;
        RECT 215.170 -55.840 215.340 -55.670 ;
        RECT 215.510 -55.840 215.680 -55.670 ;
        RECT -149.920 -68.500 -148.000 -68.320 ;
        RECT 207.740 -68.040 207.910 -57.060 ;
        RECT 208.340 -68.030 208.510 -57.050 ;
        RECT 208.950 -68.040 209.120 -57.060 ;
        RECT 209.550 -67.990 209.720 -57.010 ;
        RECT 210.150 -67.990 210.320 -57.010 ;
        RECT 210.740 -68.000 210.910 -57.020 ;
        RECT 211.320 -68.020 211.490 -57.040 ;
        RECT 211.940 -68.030 212.110 -57.050 ;
        RECT 212.560 -68.030 212.730 -57.050 ;
        RECT 214.510 -62.520 214.680 -62.350 ;
        RECT 214.850 -62.520 215.020 -62.350 ;
        RECT 215.190 -62.520 215.360 -62.350 ;
        RECT 215.530 -62.520 215.700 -62.350 ;
        RECT -149.930 -68.850 -148.010 -68.680 ;
        RECT -149.930 -68.860 -149.140 -68.850 ;
        RECT 213.690 -67.800 213.860 -67.790 ;
        RECT 211.590 -69.220 213.510 -69.040 ;
        RECT 211.600 -69.570 213.520 -69.400 ;
        RECT 212.730 -69.580 213.520 -69.570 ;
        RECT 213.690 -69.660 213.870 -67.800 ;
        RECT -150.040 -70.600 -149.110 -70.400 ;
        RECT -150.270 -74.170 -150.090 -71.010 ;
        RECT -147.170 -71.670 -143.870 -71.320 ;
        RECT -152.090 -83.710 -151.920 -83.540 ;
        RECT -151.750 -83.710 -151.580 -83.540 ;
        RECT -151.410 -83.710 -151.240 -83.540 ;
        RECT -151.070 -83.710 -150.900 -83.540 ;
        RECT -148.380 -82.170 -148.210 -72.720 ;
        RECT -147.630 -82.180 -147.460 -72.790 ;
        RECT -146.910 -82.150 -146.740 -72.750 ;
        RECT -146.250 -82.140 -146.080 -72.770 ;
        RECT -145.600 -82.150 -145.430 -72.700 ;
        RECT -144.960 -82.140 -144.790 -72.750 ;
        RECT -152.110 -90.390 -151.940 -90.220 ;
        RECT -151.770 -90.390 -151.600 -90.220 ;
        RECT -151.430 -90.390 -151.260 -90.220 ;
        RECT -151.090 -90.390 -150.920 -90.220 ;
        RECT -150.270 -95.670 -150.100 -95.660 ;
        RECT -150.280 -97.530 -150.100 -95.670 ;
        RECT -149.140 -95.900 -148.970 -84.920 ;
        RECT -148.520 -95.900 -148.350 -84.920 ;
        RECT -147.900 -95.890 -147.730 -84.910 ;
        RECT -147.320 -95.870 -147.150 -84.890 ;
        RECT -146.730 -95.860 -146.560 -84.880 ;
        RECT -146.130 -95.860 -145.960 -84.880 ;
        RECT -145.530 -95.910 -145.360 -84.930 ;
        RECT -144.920 -95.900 -144.750 -84.920 ;
        RECT -144.320 -95.910 -144.150 -84.930 ;
        RECT -149.920 -97.090 -148.000 -96.910 ;
        RECT -149.930 -97.440 -148.010 -97.270 ;
        RECT -149.930 -97.450 -149.140 -97.440 ;
        RECT -150.040 -99.190 -149.110 -98.990 ;
        RECT -150.270 -102.760 -150.090 -99.600 ;
        RECT -147.170 -100.260 -143.870 -99.910 ;
        RECT -152.090 -112.300 -151.920 -112.130 ;
        RECT -151.750 -112.300 -151.580 -112.130 ;
        RECT -151.410 -112.300 -151.240 -112.130 ;
        RECT -151.070 -112.300 -150.900 -112.130 ;
        RECT -148.380 -110.760 -148.210 -101.310 ;
        RECT -147.630 -110.770 -147.460 -101.380 ;
        RECT -146.910 -110.740 -146.740 -101.340 ;
        RECT -146.250 -110.730 -146.080 -101.360 ;
        RECT -145.600 -110.740 -145.430 -101.290 ;
        RECT -144.960 -110.730 -144.790 -101.340 ;
        RECT -152.110 -118.980 -151.940 -118.810 ;
        RECT -151.770 -118.980 -151.600 -118.810 ;
        RECT -151.430 -118.980 -151.260 -118.810 ;
        RECT -151.090 -118.980 -150.920 -118.810 ;
        RECT -150.270 -124.260 -150.100 -124.250 ;
        RECT -150.280 -126.120 -150.100 -124.260 ;
        RECT -149.140 -124.490 -148.970 -113.510 ;
        RECT -148.520 -124.490 -148.350 -113.510 ;
        RECT -147.900 -124.480 -147.730 -113.500 ;
        RECT -147.320 -124.460 -147.150 -113.480 ;
        RECT -146.730 -124.450 -146.560 -113.470 ;
        RECT -146.130 -124.450 -145.960 -113.470 ;
        RECT -145.530 -124.500 -145.360 -113.520 ;
        RECT -144.920 -124.490 -144.750 -113.510 ;
        RECT -144.320 -124.500 -144.150 -113.520 ;
        RECT -149.920 -125.680 -148.000 -125.500 ;
        RECT -149.930 -126.030 -148.010 -125.860 ;
        RECT -149.930 -126.040 -149.140 -126.030 ;
        RECT -150.040 -127.780 -149.110 -127.580 ;
        RECT -150.270 -131.350 -150.090 -128.190 ;
        RECT -147.170 -128.850 -143.870 -128.500 ;
        RECT -152.090 -140.890 -151.920 -140.720 ;
        RECT -151.750 -140.890 -151.580 -140.720 ;
        RECT -151.410 -140.890 -151.240 -140.720 ;
        RECT -151.070 -140.890 -150.900 -140.720 ;
        RECT -148.380 -139.350 -148.210 -129.900 ;
        RECT -147.630 -139.360 -147.460 -129.970 ;
        RECT -146.910 -139.330 -146.740 -129.930 ;
        RECT -146.250 -139.320 -146.080 -129.950 ;
        RECT -145.600 -139.330 -145.430 -129.880 ;
        RECT -144.960 -139.320 -144.790 -129.930 ;
        RECT -152.110 -147.570 -151.940 -147.400 ;
        RECT -151.770 -147.570 -151.600 -147.400 ;
        RECT -151.430 -147.570 -151.260 -147.400 ;
        RECT -151.090 -147.570 -150.920 -147.400 ;
        RECT -150.270 -152.850 -150.100 -152.840 ;
        RECT -150.280 -154.710 -150.100 -152.850 ;
        RECT -149.140 -153.080 -148.970 -142.100 ;
        RECT -148.520 -153.080 -148.350 -142.100 ;
        RECT -147.900 -153.070 -147.730 -142.090 ;
        RECT -147.320 -153.050 -147.150 -142.070 ;
        RECT -146.730 -153.040 -146.560 -142.060 ;
        RECT -146.130 -153.040 -145.960 -142.060 ;
        RECT -145.530 -153.090 -145.360 -142.110 ;
        RECT -144.920 -153.080 -144.750 -142.100 ;
        RECT -144.320 -153.090 -144.150 -142.110 ;
        RECT -149.920 -154.270 -148.000 -154.090 ;
        RECT -149.930 -154.620 -148.010 -154.450 ;
        RECT -149.930 -154.630 -149.140 -154.620 ;
        RECT -150.040 -156.370 -149.110 -156.170 ;
        RECT -150.270 -159.940 -150.090 -156.780 ;
        RECT -147.170 -157.440 -143.870 -157.090 ;
        RECT -152.090 -169.480 -151.920 -169.310 ;
        RECT -151.750 -169.480 -151.580 -169.310 ;
        RECT -151.410 -169.480 -151.240 -169.310 ;
        RECT -151.070 -169.480 -150.900 -169.310 ;
        RECT -148.380 -167.940 -148.210 -158.490 ;
        RECT -147.630 -167.950 -147.460 -158.560 ;
        RECT -146.910 -167.920 -146.740 -158.520 ;
        RECT -146.250 -167.910 -146.080 -158.540 ;
        RECT -145.600 -167.920 -145.430 -158.470 ;
        RECT -144.960 -167.910 -144.790 -158.520 ;
        RECT -152.110 -176.160 -151.940 -175.990 ;
        RECT -151.770 -176.160 -151.600 -175.990 ;
        RECT -151.430 -176.160 -151.260 -175.990 ;
        RECT -151.090 -176.160 -150.920 -175.990 ;
        RECT -150.270 -181.440 -150.100 -181.430 ;
        RECT -150.280 -183.300 -150.100 -181.440 ;
        RECT -149.140 -181.670 -148.970 -170.690 ;
        RECT -148.520 -181.670 -148.350 -170.690 ;
        RECT -147.900 -181.660 -147.730 -170.680 ;
        RECT -147.320 -181.640 -147.150 -170.660 ;
        RECT -146.730 -181.630 -146.560 -170.650 ;
        RECT -146.130 -181.630 -145.960 -170.650 ;
        RECT -145.530 -181.680 -145.360 -170.700 ;
        RECT -144.920 -181.670 -144.750 -170.690 ;
        RECT -144.320 -181.680 -144.150 -170.700 ;
        RECT -149.920 -182.860 -148.000 -182.680 ;
        RECT -149.930 -183.210 -148.010 -183.040 ;
        RECT -149.930 -183.220 -149.140 -183.210 ;
        RECT -150.040 -184.960 -149.110 -184.760 ;
        RECT -150.270 -188.530 -150.090 -185.370 ;
        RECT -147.170 -186.030 -143.870 -185.680 ;
        RECT -152.090 -198.070 -151.920 -197.900 ;
        RECT -151.750 -198.070 -151.580 -197.900 ;
        RECT -151.410 -198.070 -151.240 -197.900 ;
        RECT -151.070 -198.070 -150.900 -197.900 ;
        RECT -148.380 -196.530 -148.210 -187.080 ;
        RECT -147.630 -196.540 -147.460 -187.150 ;
        RECT -146.910 -196.510 -146.740 -187.110 ;
        RECT -146.250 -196.500 -146.080 -187.130 ;
        RECT -145.600 -196.510 -145.430 -187.060 ;
        RECT -144.960 -196.500 -144.790 -187.110 ;
        RECT -152.110 -204.750 -151.940 -204.580 ;
        RECT -151.770 -204.750 -151.600 -204.580 ;
        RECT -151.430 -204.750 -151.260 -204.580 ;
        RECT -151.090 -204.750 -150.920 -204.580 ;
        RECT -150.270 -210.030 -150.100 -210.020 ;
        RECT -150.280 -211.890 -150.100 -210.030 ;
        RECT -149.140 -210.260 -148.970 -199.280 ;
        RECT -148.520 -210.260 -148.350 -199.280 ;
        RECT -147.900 -210.250 -147.730 -199.270 ;
        RECT -147.320 -210.230 -147.150 -199.250 ;
        RECT -146.730 -210.220 -146.560 -199.240 ;
        RECT -146.130 -210.220 -145.960 -199.240 ;
        RECT -145.530 -210.270 -145.360 -199.290 ;
        RECT -144.920 -210.260 -144.750 -199.280 ;
        RECT -144.320 -210.270 -144.150 -199.290 ;
        RECT -149.920 -211.450 -148.000 -211.270 ;
        RECT -149.930 -211.800 -148.010 -211.630 ;
        RECT -149.930 -211.810 -149.140 -211.800 ;
        RECT -150.040 -213.550 -149.110 -213.350 ;
        RECT -150.270 -217.120 -150.090 -213.960 ;
        RECT -147.170 -214.620 -143.870 -214.270 ;
        RECT -152.090 -226.660 -151.920 -226.490 ;
        RECT -151.750 -226.660 -151.580 -226.490 ;
        RECT -151.410 -226.660 -151.240 -226.490 ;
        RECT -151.070 -226.660 -150.900 -226.490 ;
        RECT -148.380 -225.120 -148.210 -215.670 ;
        RECT -147.630 -225.130 -147.460 -215.740 ;
        RECT -146.910 -225.100 -146.740 -215.700 ;
        RECT -146.250 -225.090 -146.080 -215.720 ;
        RECT -145.600 -225.100 -145.430 -215.650 ;
        RECT -144.960 -225.090 -144.790 -215.700 ;
        RECT -152.110 -233.340 -151.940 -233.170 ;
        RECT -151.770 -233.340 -151.600 -233.170 ;
        RECT -151.430 -233.340 -151.260 -233.170 ;
        RECT -151.090 -233.340 -150.920 -233.170 ;
        RECT -150.270 -238.620 -150.100 -238.610 ;
        RECT -150.280 -240.480 -150.100 -238.620 ;
        RECT -149.140 -238.850 -148.970 -227.870 ;
        RECT -148.520 -238.850 -148.350 -227.870 ;
        RECT -147.900 -238.840 -147.730 -227.860 ;
        RECT -147.320 -238.820 -147.150 -227.840 ;
        RECT -146.730 -238.810 -146.560 -227.830 ;
        RECT -146.130 -238.810 -145.960 -227.830 ;
        RECT -145.530 -238.860 -145.360 -227.880 ;
        RECT -144.920 -238.850 -144.750 -227.870 ;
        RECT -144.320 -238.860 -144.150 -227.880 ;
        RECT -149.920 -240.040 -148.000 -239.860 ;
        RECT -149.930 -240.390 -148.010 -240.220 ;
        RECT -149.930 -240.400 -149.140 -240.390 ;
      LAYER met1 ;
        RECT -4.490 143.690 -2.080 144.330 ;
        RECT -124.420 143.120 -124.070 143.270 ;
        RECT -95.830 143.120 -95.480 143.270 ;
        RECT -67.240 143.120 -66.890 143.270 ;
        RECT -124.430 142.170 -124.060 143.120 ;
        RECT -95.840 142.170 -95.470 143.120 ;
        RECT -67.250 142.170 -66.880 143.120 ;
        RECT -4.470 142.340 -4.060 143.690 ;
        RECT 2.260 142.760 2.670 143.800 ;
        RECT 10.140 143.740 14.030 145.710 ;
        RECT 10.140 143.150 14.040 143.740 ;
        RECT -126.210 141.800 -122.310 142.170 ;
        RECT -97.620 141.800 -93.720 142.170 ;
        RECT -69.030 141.800 -65.130 142.170 ;
        RECT -25.220 142.150 -0.850 142.170 ;
        RECT -138.330 141.000 -135.960 141.630 ;
        RECT -138.300 139.040 -137.350 141.000 ;
        RECT -136.600 140.980 -136.020 141.000 ;
        RECT -126.220 140.340 -122.310 141.800 ;
        RECT -114.990 141.150 -110.860 141.550 ;
        RECT -114.990 141.060 -110.850 141.150 ;
        RECT -135.930 140.330 -122.310 140.340 ;
        RECT -138.070 133.370 -137.350 139.040 ;
        RECT -136.600 139.770 -122.310 140.330 ;
        RECT -111.380 140.160 -110.850 141.060 ;
        RECT -109.740 141.000 -107.370 141.630 ;
        RECT -136.600 135.470 -113.250 139.770 ;
        RECT -109.710 139.040 -108.760 141.000 ;
        RECT -108.010 140.980 -107.430 141.000 ;
        RECT -97.630 140.340 -93.720 141.800 ;
        RECT -86.400 141.150 -82.270 141.550 ;
        RECT -86.400 141.060 -82.260 141.150 ;
        RECT -107.340 140.330 -93.720 140.340 ;
        RECT -112.480 138.350 -111.910 138.360 ;
        RECT -136.600 135.190 -122.310 135.470 ;
        RECT -126.220 133.640 -122.310 135.190 ;
        RECT -112.480 134.930 -111.860 138.350 ;
        RECT -112.480 134.920 -111.910 134.930 ;
        RECT -126.240 132.100 -122.290 133.640 ;
        RECT -113.310 133.290 -112.750 133.790 ;
        RECT -109.480 133.370 -108.760 139.040 ;
        RECT -108.010 139.770 -93.720 140.330 ;
        RECT -82.790 140.160 -82.260 141.060 ;
        RECT -81.150 141.000 -78.780 141.630 ;
        RECT -108.010 135.470 -84.660 139.770 ;
        RECT -81.120 139.040 -80.170 141.000 ;
        RECT -79.420 140.980 -78.840 141.000 ;
        RECT -69.040 140.340 -65.130 141.800 ;
        RECT -25.280 141.760 -0.850 142.150 ;
        RECT -57.810 141.150 -53.680 141.550 ;
        RECT -57.810 141.060 -53.670 141.150 ;
        RECT -78.750 140.330 -65.130 140.340 ;
        RECT -83.890 138.350 -83.320 138.360 ;
        RECT -108.010 135.190 -93.720 135.470 ;
        RECT -97.630 133.640 -93.720 135.190 ;
        RECT -83.890 134.930 -83.270 138.350 ;
        RECT -83.890 134.920 -83.320 134.930 ;
        RECT -113.300 133.070 -112.750 133.290 ;
        RECT -97.650 132.870 -93.700 133.640 ;
        RECT -84.720 133.290 -84.160 133.790 ;
        RECT -80.890 133.370 -80.170 139.040 ;
        RECT -79.420 139.770 -65.130 140.330 ;
        RECT -54.200 140.160 -53.670 141.060 ;
        RECT -79.420 135.470 -56.070 139.770 ;
        RECT -55.300 138.350 -54.730 138.360 ;
        RECT -79.420 135.190 -65.130 135.470 ;
        RECT -69.040 133.640 -65.130 135.190 ;
        RECT -55.300 134.930 -54.680 138.350 ;
        RECT -55.300 134.920 -54.730 134.930 ;
        RECT -84.710 133.070 -84.160 133.290 ;
        RECT -97.640 132.100 -93.690 132.870 ;
        RECT -69.060 132.100 -65.110 133.640 ;
        RECT -56.130 133.290 -55.570 133.790 ;
        RECT -25.280 133.510 -24.870 141.760 ;
        RECT 1.320 141.630 3.680 142.760 ;
        RECT 10.140 142.170 10.430 143.150 ;
        RECT 16.780 143.120 17.130 143.270 ;
        RECT 45.370 143.120 45.720 143.270 ;
        RECT 73.960 143.120 74.310 143.270 ;
        RECT 102.550 143.120 102.900 143.270 ;
        RECT 131.140 143.120 131.490 143.270 ;
        RECT 159.730 143.120 160.080 143.270 ;
        RECT 188.320 143.120 188.670 143.270 ;
        RECT 16.770 142.170 17.140 143.120 ;
        RECT 45.360 142.170 45.730 143.120 ;
        RECT 73.950 142.170 74.320 143.120 ;
        RECT 102.540 142.170 102.910 143.120 ;
        RECT 131.130 142.170 131.500 143.120 ;
        RECT 159.720 142.170 160.090 143.120 ;
        RECT 188.310 142.170 188.680 143.120 ;
        RECT 7.950 142.160 28.240 142.170 ;
        RECT 7.890 142.150 28.240 142.160 ;
        RECT 7.890 141.770 29.180 142.150 ;
        RECT 43.580 141.800 47.480 142.170 ;
        RECT 72.170 141.800 76.070 142.170 ;
        RECT 100.760 141.800 104.660 142.170 ;
        RECT 129.350 141.800 133.250 142.170 ;
        RECT 157.940 141.800 161.840 142.170 ;
        RECT 186.530 141.800 190.430 142.170 ;
        RECT 7.890 141.760 29.150 141.770 ;
        RECT 1.320 141.000 5.240 141.630 ;
        RECT 1.320 134.260 3.850 141.000 ;
        RECT 4.600 140.980 5.180 141.000 ;
        RECT 14.980 140.340 18.890 141.760 ;
        RECT 26.210 141.150 30.340 141.550 ;
        RECT 26.210 141.060 30.350 141.150 ;
        RECT 5.270 140.330 18.890 140.340 ;
        RECT 4.600 139.770 18.890 140.330 ;
        RECT 29.820 140.160 30.350 141.060 ;
        RECT 31.460 141.000 33.830 141.630 ;
        RECT 4.600 135.470 27.950 139.770 ;
        RECT 31.490 139.040 32.440 141.000 ;
        RECT 33.190 140.980 33.770 141.000 ;
        RECT 43.570 140.340 47.480 141.800 ;
        RECT 54.800 141.150 58.930 141.550 ;
        RECT 54.800 141.060 58.940 141.150 ;
        RECT 33.860 140.330 47.480 140.340 ;
        RECT 28.720 138.350 29.290 138.360 ;
        RECT 4.600 135.190 18.890 135.470 ;
        RECT 1.200 133.440 3.850 134.260 ;
        RECT 14.980 133.640 18.890 135.190 ;
        RECT 28.720 134.930 29.340 138.350 ;
        RECT 28.720 134.920 29.290 134.930 ;
        RECT 3.130 133.370 3.850 133.440 ;
        RECT -56.120 133.120 -55.570 133.290 ;
        RECT -56.170 133.070 -55.570 133.120 ;
        RECT -150.030 129.880 -149.040 129.890 ;
        RECT -150.430 129.360 -149.040 129.880 ;
        RECT -150.430 125.750 -149.940 129.360 ;
        RECT -147.230 128.830 -143.810 128.880 ;
        RECT -147.240 128.260 -143.800 128.830 ;
        RECT -148.650 118.430 -144.350 127.490 ;
        RECT -142.670 127.440 -141.950 127.990 ;
        RECT -142.670 127.430 -142.170 127.440 ;
        RECT -125.540 122.220 -122.310 132.100 ;
        RECT -96.950 125.630 -93.720 132.100 ;
        RECT -68.360 129.920 -65.130 132.100 ;
        RECT -68.790 127.180 -64.960 129.920 ;
        RECT -56.170 126.560 -55.650 133.070 ;
        RECT -56.230 126.050 -55.580 126.560 ;
        RECT -97.110 122.740 -93.610 125.630 ;
        RECT -127.710 118.600 -122.310 122.220 ;
        RECT -140.150 118.520 -136.760 118.590 ;
        RECT -142.520 118.440 -141.750 118.450 ;
        RECT -141.120 118.440 -136.760 118.520 ;
        RECT -142.520 118.430 -136.760 118.440 ;
        RECT -151.050 116.680 -136.760 118.430 ;
        RECT -127.710 118.420 -124.770 118.600 ;
        RECT -56.170 118.370 -55.650 126.050 ;
        RECT -52.770 122.140 -52.360 133.350 ;
        RECT -25.660 132.870 -24.500 133.260 ;
        RECT -26.290 132.100 -23.810 132.870 ;
        RECT 14.960 132.110 18.910 133.640 ;
        RECT 27.890 133.400 28.450 133.790 ;
        RECT 27.300 133.260 28.450 133.400 ;
        RECT -25.660 131.350 -24.500 132.100 ;
        RECT -25.660 130.220 1.700 131.350 ;
        RECT -25.660 130.020 1.890 130.220 ;
        RECT 0.370 129.630 1.700 130.020 ;
        RECT 0.360 129.180 1.700 129.630 ;
        RECT -25.740 128.340 -25.240 128.820 ;
        RECT 0.360 128.760 13.880 129.180 ;
        RECT 15.660 129.110 18.890 132.110 ;
        RECT 27.280 131.300 28.460 133.260 ;
        RECT 26.480 130.390 28.460 131.300 ;
        RECT 26.480 130.210 28.290 130.390 ;
        RECT 31.720 130.250 32.440 139.040 ;
        RECT 33.190 139.770 47.480 140.330 ;
        RECT 58.410 140.160 58.940 141.060 ;
        RECT 60.050 141.000 62.420 141.630 ;
        RECT 33.190 135.470 56.540 139.770 ;
        RECT 60.080 139.040 61.030 141.000 ;
        RECT 61.780 140.980 62.360 141.000 ;
        RECT 72.160 140.340 76.070 141.800 ;
        RECT 83.390 141.150 87.520 141.550 ;
        RECT 83.390 141.060 87.530 141.150 ;
        RECT 62.450 140.330 76.070 140.340 ;
        RECT 57.310 138.350 57.880 138.360 ;
        RECT 33.190 135.190 47.480 135.470 ;
        RECT 43.570 133.640 47.480 135.190 ;
        RECT 57.310 134.930 57.930 138.350 ;
        RECT 57.310 134.920 57.880 134.930 ;
        RECT 43.550 132.100 47.500 133.640 ;
        RECT 56.480 133.290 57.040 133.790 ;
        RECT 56.490 133.070 57.040 133.290 ;
        RECT 52.430 132.350 52.770 132.490 ;
        RECT 60.310 132.350 61.030 139.040 ;
        RECT 61.780 139.770 76.070 140.330 ;
        RECT 87.000 140.160 87.530 141.060 ;
        RECT 88.640 141.000 91.010 141.630 ;
        RECT 61.780 135.470 85.130 139.770 ;
        RECT 88.670 139.040 89.620 141.000 ;
        RECT 90.370 140.980 90.950 141.000 ;
        RECT 100.750 140.340 104.660 141.800 ;
        RECT 111.980 141.150 116.110 141.550 ;
        RECT 111.980 141.060 116.120 141.150 ;
        RECT 91.040 140.330 104.660 140.340 ;
        RECT 85.900 138.350 86.470 138.360 ;
        RECT 61.780 135.190 76.070 135.470 ;
        RECT 72.160 133.640 76.070 135.190 ;
        RECT 85.900 134.930 86.520 138.350 ;
        RECT 85.900 134.920 86.470 134.930 ;
        RECT 15.670 129.090 18.860 129.110 ;
        RECT 0.360 128.620 1.700 128.760 ;
        RECT -52.890 121.670 -52.360 122.140 ;
        RECT -56.370 117.640 -55.650 118.370 ;
        RECT -152.000 116.670 -136.760 116.680 ;
        RECT -152.150 116.320 -136.760 116.670 ;
        RECT -152.000 116.310 -136.760 116.320 ;
        RECT -151.050 114.530 -136.760 116.310 ;
        RECT -150.680 114.520 -136.760 114.530 ;
        RECT -149.220 104.810 -144.070 114.520 ;
        RECT -142.520 114.500 -141.120 114.520 ;
        RECT -150.510 104.720 -149.880 104.780 ;
        RECT -150.510 104.140 -149.860 104.720 ;
        RECT -149.210 104.140 -144.070 104.810 ;
        RECT -150.510 103.390 -149.880 104.140 ;
        RECT -150.510 102.670 -142.250 103.390 ;
        RECT -150.510 102.440 -147.920 102.670 ;
        RECT -150.510 102.410 -149.880 102.440 ;
        RECT -150.030 101.290 -149.040 101.300 ;
        RECT -150.430 100.770 -149.040 101.290 ;
        RECT -150.430 97.160 -149.940 100.770 ;
        RECT -147.230 100.240 -143.810 100.290 ;
        RECT -147.240 99.670 -143.800 100.240 ;
        RECT -148.650 89.840 -144.350 98.900 ;
        RECT -142.670 98.850 -141.950 99.400 ;
        RECT -142.670 98.840 -142.170 98.850 ;
        RECT -142.520 89.840 -141.120 89.860 ;
        RECT -130.980 89.840 -128.720 89.880 ;
        RECT -151.050 88.090 -128.720 89.840 ;
        RECT -152.000 88.080 -128.720 88.090 ;
        RECT -152.150 87.730 -128.720 88.080 ;
        RECT -152.000 87.720 -128.720 87.730 ;
        RECT -151.050 86.610 -128.720 87.720 ;
        RECT -151.050 85.940 -141.120 86.610 ;
        RECT -130.980 86.570 -128.720 86.610 ;
        RECT -150.680 85.930 -141.120 85.940 ;
        RECT -149.220 76.220 -144.070 85.930 ;
        RECT -142.520 85.920 -141.120 85.930 ;
        RECT -142.520 85.910 -141.750 85.920 ;
        RECT -56.170 82.290 -55.650 117.640 ;
        RECT -52.770 117.420 -52.360 121.670 ;
        RECT -25.640 125.380 -25.250 128.340 ;
        RECT -5.050 128.020 -2.280 128.260 ;
        RECT -23.270 127.560 -23.010 127.760 ;
        RECT -20.410 127.720 -20.150 127.810 ;
        RECT -23.330 127.250 -22.950 127.560 ;
        RECT -21.920 127.250 -20.890 127.560 ;
        RECT -20.420 127.490 -20.130 127.720 ;
        RECT -23.280 126.460 -23.020 126.730 ;
        RECT -22.590 126.460 -22.270 126.700 ;
        RECT -21.870 126.460 -21.610 126.740 ;
        RECT -23.320 125.800 -21.570 126.460 ;
        RECT -23.280 125.540 -23.020 125.800 ;
        RECT -22.590 125.540 -22.270 125.800 ;
        RECT -21.850 125.560 -21.590 125.800 ;
        RECT -25.640 124.890 -25.170 125.380 ;
        RECT -25.640 124.880 -25.190 124.890 ;
        RECT -52.910 116.830 -52.290 117.420 ;
        RECT -56.250 81.690 -55.620 82.290 ;
        RECT -52.770 81.270 -52.360 116.830 ;
        RECT -52.820 80.770 -52.340 81.270 ;
        RECT -150.510 76.130 -149.880 76.190 ;
        RECT -150.510 75.550 -149.860 76.130 ;
        RECT -149.210 75.550 -144.070 76.220 ;
        RECT -150.510 74.800 -149.880 75.550 ;
        RECT -150.510 74.080 -142.250 74.800 ;
        RECT -150.510 73.850 -147.920 74.080 ;
        RECT -150.510 73.820 -149.880 73.850 ;
        RECT -150.030 72.700 -149.040 72.710 ;
        RECT -150.430 72.180 -149.040 72.700 ;
        RECT -150.430 68.570 -149.940 72.180 ;
        RECT -147.230 71.650 -143.810 71.700 ;
        RECT -147.240 71.080 -143.800 71.650 ;
        RECT -148.650 61.250 -144.350 70.310 ;
        RECT -142.670 70.260 -141.950 70.810 ;
        RECT -142.670 70.250 -142.170 70.260 ;
        RECT -25.640 66.770 -25.250 124.880 ;
        RECT -23.260 124.510 -23.030 125.030 ;
        RECT -23.280 124.190 -23.020 124.510 ;
        RECT -24.230 123.740 -23.970 124.060 ;
        RECT -24.220 121.520 -23.980 123.740 ;
        RECT -23.260 123.620 -23.030 124.190 ;
        RECT -21.850 123.620 -21.620 125.030 ;
        RECT -21.130 124.480 -20.890 127.250 ;
        RECT -5.050 126.930 -4.810 128.020 ;
        RECT -20.470 126.800 -20.080 126.930 ;
        RECT -20.470 126.510 -20.050 126.800 ;
        RECT -5.050 126.670 -4.820 126.930 ;
        RECT -20.750 125.950 -20.430 126.270 ;
        RECT -20.700 125.720 -20.470 125.950 ;
        RECT -20.280 125.570 -20.050 126.510 ;
        RECT -5.060 126.450 -4.820 126.670 ;
        RECT -7.200 125.640 -6.880 125.960 ;
        RECT -5.840 125.720 -5.520 126.040 ;
        RECT -5.150 125.710 -4.830 126.030 ;
        RECT -20.410 125.500 -20.050 125.570 ;
        RECT -20.470 125.390 -20.050 125.500 ;
        RECT -20.470 125.270 -20.080 125.390 ;
        RECT -21.170 123.940 -20.850 124.260 ;
        RECT -20.410 124.100 -20.140 125.270 ;
        RECT -5.050 124.130 -4.810 124.770 ;
        RECT -20.410 123.870 -20.080 124.100 ;
        RECT -5.050 123.870 -4.820 124.130 ;
        RECT -5.060 123.220 -4.820 123.870 ;
        RECT -22.610 122.740 -22.290 123.060 ;
        RECT -21.180 122.760 -20.860 123.080 ;
        RECT -23.400 122.160 -23.080 122.480 ;
        RECT -22.470 122.160 -22.150 122.480 ;
        RECT -21.770 122.160 -21.450 122.480 ;
        RECT -21.030 122.160 -20.710 122.480 ;
        RECT -20.320 122.150 -20.000 122.470 ;
        RECT -24.310 121.040 -23.890 121.520 ;
        RECT -18.420 120.280 -18.130 122.970 ;
        RECT -5.060 122.580 -4.810 123.220 ;
        RECT -7.920 121.980 -7.600 122.300 ;
        RECT -18.440 119.610 -18.030 120.280 ;
        RECT -5.060 118.920 -4.820 122.580 ;
        RECT -5.110 118.580 -4.770 118.920 ;
        RECT -7.860 118.480 -7.370 118.490 ;
        RECT -11.790 109.790 -11.560 113.270 ;
        RECT -11.120 112.650 -10.900 113.270 ;
        RECT -10.010 112.740 -9.690 113.060 ;
        RECT -8.920 112.750 -8.600 113.070 ;
        RECT -11.150 112.330 -10.890 112.650 ;
        RECT -10.480 112.600 -10.160 112.650 ;
        RECT -10.480 112.370 -9.930 112.600 ;
        RECT -10.480 112.330 -10.160 112.370 ;
        RECT -11.120 111.730 -10.900 112.330 ;
        RECT -10.010 111.820 -9.690 112.140 ;
        RECT -8.920 111.830 -8.600 112.150 ;
        RECT -11.180 111.410 -10.900 111.730 ;
        RECT -10.480 111.680 -10.160 111.730 ;
        RECT -10.480 111.450 -9.930 111.680 ;
        RECT -10.480 111.410 -10.160 111.450 ;
        RECT -11.120 110.810 -10.900 111.410 ;
        RECT -10.010 110.900 -9.690 111.220 ;
        RECT -8.920 110.910 -8.600 111.230 ;
        RECT -11.170 110.490 -10.900 110.810 ;
        RECT -10.480 110.760 -10.160 110.810 ;
        RECT -10.480 110.530 -9.930 110.760 ;
        RECT -10.480 110.490 -10.160 110.530 ;
        RECT -11.820 109.470 -11.560 109.790 ;
        RECT -11.790 108.830 -11.560 109.470 ;
        RECT -11.860 108.510 -11.560 108.830 ;
        RECT -11.790 107.870 -11.560 108.510 ;
        RECT -11.820 107.550 -11.560 107.870 ;
        RECT -11.790 92.800 -11.560 107.550 ;
        RECT -11.120 92.800 -10.900 110.490 ;
        RECT -10.200 109.920 -9.880 110.240 ;
        RECT -8.900 109.820 -8.580 110.140 ;
        RECT -10.200 109.740 -9.880 109.780 ;
        RECT -10.430 109.510 -9.880 109.740 ;
        RECT -10.200 109.460 -9.880 109.510 ;
        RECT -10.200 108.960 -9.880 109.280 ;
        RECT -8.900 108.860 -8.580 109.180 ;
        RECT -10.200 108.780 -9.880 108.820 ;
        RECT -10.430 108.550 -9.880 108.780 ;
        RECT -10.200 108.500 -9.880 108.550 ;
        RECT -10.200 108.000 -9.880 108.320 ;
        RECT -8.900 107.900 -8.580 108.220 ;
        RECT -10.200 107.820 -9.880 107.860 ;
        RECT -10.430 107.590 -9.880 107.820 ;
        RECT -8.430 107.730 -8.210 117.540 ;
        RECT -7.870 117.330 -7.360 118.480 ;
        RECT -2.520 117.550 -2.280 128.020 ;
        RECT 0.790 127.690 3.820 127.960 ;
        RECT 0.790 126.710 1.060 127.690 ;
        RECT 0.800 124.500 1.060 124.520 ;
        RECT 0.760 118.520 1.070 124.500 ;
        RECT 1.940 122.000 2.260 122.320 ;
        RECT 0.680 118.150 1.070 118.520 ;
        RECT 3.550 118.010 3.820 127.690 ;
        RECT 5.500 126.670 5.760 128.760 ;
        RECT 13.460 125.510 13.880 128.760 ;
        RECT 17.270 126.270 17.690 129.090 ;
        RECT 17.270 125.790 17.740 126.270 ;
        RECT 13.420 125.030 13.900 125.510 ;
        RECT 4.730 123.960 4.960 124.130 ;
        RECT 4.720 122.090 4.970 123.960 ;
        RECT 18.970 123.420 19.410 123.920 ;
        RECT 24.690 123.420 25.130 123.920 ;
        RECT 14.550 122.400 14.990 122.900 ;
        RECT 4.720 121.910 4.980 122.090 ;
        RECT 4.720 119.010 4.970 121.910 ;
        RECT 11.760 119.660 12.080 119.710 ;
        RECT 11.670 119.370 12.080 119.660 ;
        RECT 4.680 118.650 5.010 119.010 ;
        RECT 3.510 117.700 3.850 118.010 ;
        RECT -7.920 117.230 -7.360 117.330 ;
        RECT -2.570 117.230 -2.230 117.550 ;
        RECT -8.030 116.830 -7.360 117.230 ;
        RECT 11.370 117.080 11.610 117.130 ;
        RECT -8.030 116.800 -7.370 116.830 ;
        RECT -8.030 112.580 -7.810 116.800 ;
        RECT 11.670 116.730 11.910 119.370 ;
        RECT 14.610 117.130 14.920 122.400 ;
        RECT 14.310 117.060 14.920 117.130 ;
        RECT 18.740 117.080 19.030 117.130 ;
        RECT 14.610 116.730 14.920 117.060 ;
        RECT 19.040 116.730 19.330 123.420 ;
        RECT 20.230 122.430 20.730 122.870 ;
        RECT 11.560 115.870 11.910 116.730 ;
        RECT 12.980 116.090 13.330 116.380 ;
        RECT 12.980 116.070 13.180 116.090 ;
        RECT 10.820 115.230 11.230 115.560 ;
        RECT -6.810 114.680 -6.460 115.140 ;
        RECT 9.620 114.700 9.990 115.010 ;
        RECT -7.410 114.320 -7.160 114.440 ;
        RECT -7.440 113.860 -7.120 114.320 ;
        RECT -8.040 112.290 -7.810 112.580 ;
        RECT -10.200 107.540 -9.880 107.590 ;
        RECT -8.490 107.500 -8.200 107.730 ;
        RECT -11.900 92.270 -11.560 92.800 ;
        RECT -11.240 92.270 -10.900 92.800 ;
        RECT -13.210 91.530 -12.980 91.600 ;
        RECT -13.250 91.270 -12.930 91.530 ;
        RECT -13.700 91.160 -13.470 91.200 ;
        RECT -13.740 90.840 -13.470 91.160 ;
        RECT -23.050 89.600 -22.330 90.300 ;
        RECT -23.040 84.450 -22.380 89.600 ;
        RECT -13.700 87.320 -13.470 90.840 ;
        RECT -13.210 88.800 -12.980 91.270 ;
        RECT -11.790 91.180 -11.560 92.270 ;
        RECT -11.120 91.540 -10.900 92.270 ;
        RECT -9.360 91.560 -9.090 91.600 ;
        RECT -11.140 91.220 -10.880 91.540 ;
        RECT -9.380 91.230 -9.090 91.560 ;
        RECT -11.800 90.860 -11.540 91.180 ;
        RECT -11.080 90.260 -10.760 90.580 ;
        RECT -10.430 90.260 -10.110 90.580 ;
        RECT -12.300 89.820 -11.980 90.140 ;
        RECT -11.600 89.820 -11.280 90.140 ;
        RECT -9.910 88.810 -9.620 89.720 ;
        RECT -13.210 88.790 -12.480 88.800 ;
        RECT -13.210 88.470 -12.460 88.790 ;
        RECT -13.210 88.430 -12.480 88.470 ;
        RECT -13.700 87.250 -13.440 87.320 ;
        RECT -13.720 87.240 -13.440 87.250 ;
        RECT -13.750 86.930 -13.430 87.240 ;
        RECT -17.850 85.070 -17.420 85.500 ;
        RECT -23.040 83.730 -22.300 84.450 ;
        RECT -17.800 79.260 -17.430 85.070 ;
        RECT -13.750 83.840 -13.430 84.160 ;
        RECT -13.210 83.490 -12.980 88.430 ;
        RECT -12.710 88.180 -12.480 88.430 ;
        RECT -10.000 88.240 -9.680 88.280 ;
        RECT -9.360 88.260 -9.090 91.230 ;
        RECT -9.480 88.240 -9.090 88.260 ;
        RECT -12.710 87.960 -12.490 88.180 ;
        RECT -10.000 88.010 -9.090 88.240 ;
        RECT -8.880 91.160 -8.640 91.200 ;
        RECT -8.880 90.840 -8.620 91.160 ;
        RECT -10.000 87.960 -9.680 88.010 ;
        RECT -12.690 87.530 -12.470 87.750 ;
        RECT -12.700 87.240 -12.470 87.530 ;
        RECT -9.990 87.700 -9.670 87.740 ;
        RECT -8.880 87.700 -8.640 90.840 ;
        RECT -9.990 87.470 -8.640 87.700 ;
        RECT -9.990 87.420 -9.670 87.470 ;
        RECT -12.720 86.920 -12.460 87.240 ;
        RECT -9.920 86.790 -9.650 86.970 ;
        RECT -9.940 86.470 -9.620 86.790 ;
        RECT -9.920 86.300 -9.650 86.470 ;
        RECT -12.270 85.940 -11.950 86.260 ;
        RECT -11.580 85.930 -11.260 86.250 ;
        RECT -11.100 85.160 -10.780 85.480 ;
        RECT -10.390 85.100 -10.070 85.420 ;
        RECT -10.440 84.280 -10.120 84.600 ;
        RECT -12.650 83.850 -12.330 84.170 ;
        RECT -11.560 83.850 -11.240 84.170 ;
        RECT -10.430 83.810 -10.110 84.130 ;
        RECT -13.210 83.170 -12.880 83.490 ;
        RECT -12.100 83.170 -11.780 83.490 ;
        RECT -11.000 83.170 -10.680 83.490 ;
        RECT -13.210 82.120 -12.980 83.170 ;
        RECT -10.290 83.000 -10.000 83.430 ;
        RECT -10.290 82.980 -9.820 83.000 ;
        RECT -10.280 82.680 -9.820 82.980 ;
        RECT -10.280 82.150 -10.000 82.680 ;
        RECT -13.210 81.800 -12.880 82.120 ;
        RECT -12.100 81.800 -11.780 82.120 ;
        RECT -11.000 81.800 -10.680 82.120 ;
        RECT -13.750 81.070 -13.430 81.390 ;
        RECT -13.210 80.930 -12.980 81.800 ;
        RECT -12.650 81.070 -12.330 81.390 ;
        RECT -11.560 81.070 -11.240 81.390 ;
        RECT -13.210 80.700 -10.760 80.930 ;
        RECT -11.080 80.370 -10.760 80.700 ;
        RECT -13.760 79.730 -13.440 80.050 ;
        RECT -12.650 79.720 -12.330 80.040 ;
        RECT -11.560 79.700 -11.240 80.020 ;
        RECT -17.840 78.830 -17.410 79.260 ;
        RECT -13.200 79.030 -12.880 79.350 ;
        RECT -12.100 79.020 -11.780 79.340 ;
        RECT -11.010 79.020 -10.690 79.340 ;
        RECT -10.320 78.800 -9.990 78.830 ;
        RECT -10.460 78.720 -9.990 78.800 ;
        RECT -10.700 78.480 -9.990 78.720 ;
        RECT -10.320 78.410 -9.990 78.480 ;
        RECT -14.830 73.170 -14.540 73.520 ;
        RECT -14.820 72.600 -14.560 73.170 ;
        RECT -14.180 72.070 -13.920 77.050 ;
        RECT -10.400 76.720 -10.080 77.040 ;
        RECT -13.710 76.280 -13.390 76.600 ;
        RECT -12.610 76.290 -12.290 76.610 ;
        RECT -11.520 76.290 -11.200 76.610 ;
        RECT -10.390 76.250 -10.070 76.570 ;
        RECT -13.160 75.610 -12.840 75.930 ;
        RECT -12.060 75.610 -11.740 75.930 ;
        RECT -10.960 75.610 -10.640 75.930 ;
        RECT -13.160 74.240 -12.840 74.560 ;
        RECT -12.060 74.240 -11.740 74.560 ;
        RECT -10.960 74.240 -10.640 74.560 ;
        RECT -13.710 73.510 -13.390 73.830 ;
        RECT -12.610 73.510 -12.290 73.830 ;
        RECT -11.520 73.510 -11.200 73.830 ;
        RECT -8.880 72.810 -8.640 87.470 ;
        RECT -8.430 86.800 -8.210 107.500 ;
        RECT -8.030 89.410 -7.810 112.290 ;
        RECT -7.410 113.070 -7.160 113.860 ;
        RECT -7.410 112.750 -7.120 113.070 ;
        RECT -7.410 112.150 -7.160 112.750 ;
        RECT -7.410 111.830 -7.120 112.150 ;
        RECT -7.410 111.230 -7.160 111.830 ;
        RECT -7.410 110.910 -7.150 111.230 ;
        RECT -7.410 90.560 -7.160 110.910 ;
        RECT -6.790 110.140 -6.530 114.680 ;
        RECT 8.980 112.980 9.370 113.350 ;
        RECT 8.400 111.490 8.790 111.880 ;
        RECT -6.790 109.820 -6.510 110.140 ;
        RECT 7.760 109.900 8.150 110.280 ;
        RECT 7.790 109.890 8.130 109.900 ;
        RECT -6.790 109.180 -6.530 109.820 ;
        RECT 7.150 109.700 7.490 109.710 ;
        RECT 7.140 109.310 7.500 109.700 ;
        RECT -6.790 108.860 -6.500 109.180 ;
        RECT -6.790 108.220 -6.530 108.860 ;
        RECT -6.790 107.900 -6.510 108.220 ;
        RECT -7.410 90.540 -7.150 90.560 ;
        RECT -7.420 90.260 -7.140 90.540 ;
        RECT -7.410 90.240 -7.150 90.260 ;
        RECT -8.070 89.090 -7.750 89.410 ;
        RECT -8.470 86.480 -8.190 86.800 ;
        RECT -8.430 73.510 -8.210 86.480 ;
        RECT -8.030 81.270 -7.810 89.090 ;
        RECT -8.030 80.790 -7.740 81.270 ;
        RECT -8.030 78.830 -7.810 80.790 ;
        RECT -8.050 78.410 -7.790 78.830 ;
        RECT -8.030 73.790 -7.810 78.410 ;
        RECT -7.410 75.170 -7.160 90.240 ;
        RECT -6.790 86.230 -6.530 107.900 ;
        RECT 6.530 107.750 6.890 108.140 ;
        RECT 5.880 106.210 6.290 106.610 ;
        RECT 5.350 104.650 5.710 105.040 ;
        RECT 4.770 99.590 5.100 99.610 ;
        RECT 4.710 99.170 5.100 99.590 ;
        RECT 4.140 97.980 4.470 98.000 ;
        RECT 4.090 97.590 4.480 97.980 ;
        RECT 3.520 96.430 3.850 96.440 ;
        RECT 3.490 96.040 3.850 96.430 ;
        RECT 2.870 94.560 3.260 94.960 ;
        RECT 2.200 89.390 2.630 89.790 ;
        RECT 1.540 87.820 1.950 88.220 ;
        RECT -6.800 85.910 -6.490 86.230 ;
        RECT 0.930 86.180 1.320 86.580 ;
        RECT -7.450 74.770 -7.150 75.170 ;
        RECT -8.030 73.650 -7.790 73.790 ;
        RECT -8.470 73.160 -8.160 73.510 ;
        RECT -8.020 73.020 -7.790 73.650 ;
        RECT -13.720 72.170 -13.400 72.490 ;
        RECT -12.610 72.160 -12.290 72.480 ;
        RECT -11.520 72.140 -11.200 72.460 ;
        RECT -9.670 72.250 -8.640 72.810 ;
        RECT -8.030 72.990 -7.790 73.020 ;
        RECT -9.670 72.140 -8.880 72.250 ;
        RECT -14.230 71.260 -13.920 72.070 ;
        RECT -13.160 71.470 -12.840 71.790 ;
        RECT -12.060 71.460 -11.740 71.780 ;
        RECT -10.970 71.460 -10.650 71.780 ;
        RECT -8.030 71.600 -7.810 72.990 ;
        RECT -14.180 71.060 -13.920 71.260 ;
        RECT -9.560 67.920 -7.140 71.600 ;
        RECT -6.790 67.630 -6.530 85.910 ;
        RECT 0.240 84.740 0.650 85.130 ;
        RECT -3.970 79.590 -3.040 81.240 ;
        RECT -3.880 79.110 -3.140 79.590 ;
        RECT -6.880 67.220 -6.530 67.630 ;
        RECT -25.810 66.250 -25.250 66.770 ;
        RECT 0.300 61.400 0.630 84.740 ;
        RECT 0.250 61.390 0.680 61.400 ;
        RECT -142.520 61.250 -141.750 61.270 ;
        RECT -127.070 61.250 -124.840 61.330 ;
        RECT -151.050 59.500 -124.840 61.250 ;
        RECT 0.220 60.930 0.710 61.390 ;
        RECT 0.250 60.910 0.680 60.930 ;
        RECT 0.950 60.610 1.280 86.180 ;
        RECT 0.860 60.120 1.350 60.610 ;
        RECT 1.600 59.900 1.930 87.820 ;
        RECT -152.000 59.490 -124.840 59.500 ;
        RECT -152.150 59.140 -124.840 59.490 ;
        RECT 1.570 59.440 1.970 59.900 ;
        RECT -152.000 59.130 -124.840 59.140 ;
        RECT -151.050 58.020 -124.840 59.130 ;
        RECT 1.360 58.950 1.940 59.060 ;
        RECT 2.270 58.950 2.600 89.390 ;
        RECT 2.910 63.530 3.240 94.560 ;
        RECT 2.910 59.070 3.230 63.530 ;
        RECT 3.520 59.680 3.850 96.040 ;
        RECT 4.140 59.930 4.470 97.590 ;
        RECT 4.770 60.960 5.100 99.170 ;
        RECT 5.370 61.260 5.700 104.650 ;
        RECT 5.950 61.830 6.280 106.210 ;
        RECT 6.560 62.860 6.890 107.750 ;
        RECT 7.150 63.470 7.480 109.310 ;
        RECT 7.790 64.140 8.120 109.890 ;
        RECT 8.410 64.790 8.740 111.490 ;
        RECT 9.010 65.420 9.340 112.980 ;
        RECT 9.640 66.030 9.970 114.700 ;
        RECT 10.820 113.680 11.230 114.010 ;
        RECT 10.820 112.130 11.230 112.460 ;
        RECT 11.560 110.940 11.800 115.870 ;
        RECT 14.500 115.800 14.920 116.730 ;
        RECT 17.860 116.190 18.180 116.490 ;
        RECT 18.930 115.820 19.330 116.730 ;
        RECT 12.980 114.540 13.330 114.830 ;
        RECT 12.980 114.520 13.180 114.540 ;
        RECT 12.980 112.990 13.330 113.280 ;
        RECT 12.980 112.970 13.180 112.990 ;
        RECT 12.980 111.440 13.330 111.730 ;
        RECT 12.980 111.420 13.180 111.440 ;
        RECT 14.500 110.950 14.810 115.800 ;
        RECT 15.060 115.340 15.340 115.670 ;
        RECT 17.860 114.640 18.180 114.940 ;
        RECT 15.060 113.790 15.340 114.120 ;
        RECT 17.860 113.090 18.180 113.390 ;
        RECT 15.060 112.240 15.340 112.570 ;
        RECT 17.860 111.540 18.180 111.840 ;
        RECT 10.820 110.580 11.230 110.910 ;
        RECT 11.370 110.890 11.800 110.940 ;
        RECT 14.310 110.890 14.810 110.950 ;
        RECT 11.560 110.490 11.800 110.890 ;
        RECT 14.500 110.490 14.810 110.890 ;
        RECT 15.060 110.690 15.340 111.020 ;
        RECT 18.930 110.940 19.220 115.820 ;
        RECT 18.740 110.890 19.220 110.940 ;
        RECT 18.930 110.490 19.220 110.890 ;
        RECT 14.910 109.870 14.920 109.880 ;
        RECT 11.670 109.790 11.910 109.870 ;
        RECT 14.610 109.790 14.920 109.870 ;
        RECT 19.040 109.790 19.330 109.870 ;
        RECT 20.500 109.430 20.690 122.430 ;
        RECT 22.570 110.190 22.850 110.840 ;
        RECT 22.570 109.590 22.960 110.190 ;
        RECT 10.820 108.750 11.230 109.080 ;
        RECT 11.560 108.770 11.800 109.170 ;
        RECT 14.500 108.770 14.810 109.170 ;
        RECT 11.370 108.720 11.800 108.770 ;
        RECT 10.820 107.200 11.230 107.530 ;
        RECT 10.820 105.650 11.230 105.980 ;
        RECT 10.820 104.100 11.230 104.430 ;
        RECT 11.560 103.790 11.800 108.720 ;
        RECT 14.310 108.710 14.810 108.770 ;
        RECT 12.980 108.220 13.180 108.240 ;
        RECT 12.980 107.930 13.330 108.220 ;
        RECT 12.980 106.670 13.180 106.690 ;
        RECT 12.980 106.380 13.330 106.670 ;
        RECT 12.980 105.120 13.180 105.140 ;
        RECT 12.980 104.830 13.330 105.120 ;
        RECT 14.500 103.860 14.810 108.710 ;
        RECT 15.060 108.640 15.340 108.970 ;
        RECT 18.930 108.770 19.220 109.170 ;
        RECT 18.740 108.720 19.220 108.770 ;
        RECT 17.860 107.820 18.180 108.120 ;
        RECT 15.060 107.090 15.340 107.420 ;
        RECT 17.860 106.270 18.180 106.570 ;
        RECT 15.060 105.540 15.340 105.870 ;
        RECT 17.860 104.720 18.180 105.020 ;
        RECT 15.060 103.990 15.340 104.320 ;
        RECT 11.560 102.930 11.910 103.790 ;
        RECT 12.980 103.570 13.180 103.590 ;
        RECT 12.980 103.280 13.330 103.570 ;
        RECT 14.500 102.930 14.920 103.860 ;
        RECT 18.930 103.840 19.220 108.720 ;
        RECT 22.570 106.040 22.850 109.590 ;
        RECT 23.100 109.380 23.290 110.840 ;
        RECT 24.780 110.460 25.030 123.420 ;
        RECT 26.480 123.380 27.210 130.210 ;
        RECT 31.630 130.100 32.610 130.250 ;
        RECT 26.640 112.990 26.810 123.380 ;
        RECT 31.640 122.850 32.610 130.100 ;
        RECT 44.250 129.110 47.480 132.100 ;
        RECT 52.430 131.630 61.030 132.350 ;
        RECT 72.140 132.100 76.090 133.640 ;
        RECT 85.070 133.290 85.630 133.790 ;
        RECT 85.080 133.070 85.630 133.290 ;
        RECT 81.770 132.720 81.960 132.730 ;
        RECT 88.900 132.720 89.620 139.040 ;
        RECT 90.370 139.770 104.660 140.330 ;
        RECT 115.590 140.160 116.120 141.060 ;
        RECT 117.230 141.000 119.600 141.630 ;
        RECT 90.370 135.470 113.720 139.770 ;
        RECT 117.260 139.040 118.210 141.000 ;
        RECT 118.960 140.980 119.540 141.000 ;
        RECT 129.340 140.340 133.250 141.800 ;
        RECT 140.570 141.150 144.700 141.550 ;
        RECT 140.570 141.060 144.710 141.150 ;
        RECT 119.630 140.330 133.250 140.340 ;
        RECT 114.490 138.350 115.060 138.360 ;
        RECT 90.370 135.190 104.660 135.470 ;
        RECT 100.750 133.640 104.660 135.190 ;
        RECT 114.490 134.930 115.110 138.350 ;
        RECT 114.490 134.920 115.060 134.930 ;
        RECT 81.770 132.370 89.620 132.720 ;
        RECT 44.260 129.080 47.450 129.110 ;
        RECT 37.030 125.010 38.500 125.540 ;
        RECT 31.620 122.380 32.630 122.850 ;
        RECT 34.660 122.400 35.100 122.900 ;
        RECT 28.860 118.650 29.200 118.940 ;
        RECT 28.910 118.620 29.170 118.650 ;
        RECT 27.030 115.090 27.290 115.410 ;
        RECT 27.060 112.860 27.250 115.090 ;
        RECT 28.930 112.840 29.140 118.620 ;
        RECT 32.500 118.020 32.760 118.030 ;
        RECT 32.480 117.720 32.780 118.020 ;
        RECT 32.500 117.710 32.760 117.720 ;
        RECT 29.330 116.690 29.670 117.010 ;
        RECT 29.400 112.860 29.590 116.690 ;
        RECT 29.770 114.600 30.060 114.920 ;
        RECT 29.810 112.840 30.020 114.600 ;
        RECT 30.810 114.120 31.150 114.440 ;
        RECT 30.890 112.870 31.070 114.120 ;
        RECT 24.500 110.020 25.030 110.460 ;
        RECT 24.780 109.390 25.030 110.020 ;
        RECT 29.580 109.630 29.810 110.840 ;
        RECT 30.800 109.870 31.030 110.840 ;
        RECT 23.070 109.350 23.290 109.380 ;
        RECT 23.060 109.080 23.310 109.350 ;
        RECT 23.060 109.070 23.300 109.080 ;
        RECT 23.070 108.830 23.300 109.070 ;
        RECT 24.340 109.060 24.660 109.380 ;
        RECT 29.550 108.840 29.810 109.630 ;
        RECT 30.790 109.690 31.030 109.870 ;
        RECT 30.790 109.620 31.190 109.690 ;
        RECT 30.800 109.470 31.190 109.620 ;
        RECT 31.600 109.470 31.920 109.790 ;
        RECT 32.530 109.690 32.730 117.710 ;
        RECT 34.760 112.820 34.990 122.400 ;
        RECT 35.660 118.630 35.940 118.950 ;
        RECT 35.220 117.720 35.500 118.040 ;
        RECT 30.720 108.980 31.190 109.470 ;
        RECT 31.580 109.330 31.950 109.350 ;
        RECT 31.530 109.070 31.950 109.330 ;
        RECT 31.580 109.060 31.950 109.070 ;
        RECT 23.100 106.800 23.260 108.830 ;
        RECT 23.450 108.270 23.690 108.400 ;
        RECT 23.430 107.950 23.690 108.270 ;
        RECT 23.430 107.350 23.690 107.670 ;
        RECT 23.450 107.230 23.690 107.350 ;
        RECT 26.540 106.970 26.820 107.020 ;
        RECT 23.070 106.560 23.300 106.800 ;
        RECT 26.540 106.690 26.860 106.970 ;
        RECT 27.070 106.960 27.260 107.020 ;
        RECT 29.580 106.690 29.810 108.840 ;
        RECT 30.800 108.820 31.190 108.980 ;
        RECT 30.540 108.720 31.190 108.820 ;
        RECT 30.540 108.540 31.230 108.720 ;
        RECT 30.800 108.430 31.230 108.540 ;
        RECT 30.800 107.830 31.190 108.430 ;
        RECT 30.800 107.720 31.230 107.830 ;
        RECT 30.540 107.540 31.230 107.720 ;
        RECT 30.540 107.440 31.190 107.540 ;
        RECT 30.800 107.280 31.190 107.440 ;
        RECT 30.720 106.790 31.190 107.280 ;
        RECT 32.310 107.350 32.730 109.690 ;
        RECT 31.580 107.190 31.950 107.200 ;
        RECT 31.530 106.930 31.950 107.190 ;
        RECT 31.580 106.910 31.950 106.930 ;
        RECT 32.310 107.020 32.790 107.350 ;
        RECT 23.060 106.550 23.300 106.560 ;
        RECT 23.060 106.280 23.310 106.550 ;
        RECT 24.340 106.300 24.660 106.620 ;
        RECT 23.070 106.250 23.290 106.280 ;
        RECT 22.570 105.440 22.960 106.040 ;
        RECT 22.570 104.790 22.850 105.440 ;
        RECT 23.100 104.790 23.290 106.250 ;
        RECT 29.550 105.900 29.810 106.690 ;
        RECT 30.800 106.540 31.190 106.790 ;
        RECT 30.720 106.050 31.190 106.540 ;
        RECT 31.580 106.400 31.950 106.420 ;
        RECT 31.530 106.140 31.950 106.400 ;
        RECT 31.580 106.130 31.950 106.140 ;
        RECT 24.500 105.170 24.810 105.610 ;
        RECT 29.580 104.790 29.810 105.900 ;
        RECT 30.800 105.890 31.190 106.050 ;
        RECT 30.540 105.790 31.190 105.890 ;
        RECT 30.540 105.610 31.230 105.790 ;
        RECT 31.630 105.780 31.950 106.100 ;
        RECT 30.800 105.500 31.230 105.610 ;
        RECT 30.800 104.900 31.190 105.500 ;
        RECT 30.800 104.790 31.230 104.900 ;
        RECT 30.540 104.510 30.860 104.790 ;
        RECT 31.000 104.610 31.230 104.790 ;
        RECT 31.000 104.350 31.190 104.610 ;
        RECT 30.720 103.860 31.190 104.350 ;
        RECT 31.580 104.260 31.950 104.270 ;
        RECT 31.530 104.000 31.950 104.260 ;
        RECT 31.580 103.980 31.950 104.000 ;
        RECT 17.860 103.170 18.180 103.470 ;
        RECT 18.930 102.930 19.330 103.840 ;
        RECT 11.370 102.530 11.610 102.580 ;
        RECT 11.670 99.420 11.910 102.930 ;
        RECT 14.610 102.600 14.920 102.930 ;
        RECT 14.310 102.530 14.920 102.600 ;
        RECT 18.740 102.530 19.030 102.580 ;
        RECT 14.610 99.350 14.920 102.530 ;
        RECT 19.040 99.370 19.330 102.930 ;
        RECT 20.500 99.380 20.690 103.780 ;
        RECT 21.810 99.570 22.040 103.820 ;
        RECT 24.780 99.570 25.030 103.840 ;
        RECT 31.000 103.640 31.190 103.860 ;
        RECT 32.310 103.640 32.540 107.020 ;
        RECT 33.090 104.800 33.510 110.840 ;
        RECT 35.250 109.690 35.470 117.720 ;
        RECT 35.250 109.470 35.530 109.690 ;
        RECT 35.680 109.470 35.910 118.630 ;
        RECT 37.050 112.630 37.470 125.010 ;
        RECT 38.080 112.630 38.500 125.010 ;
        RECT 40.460 122.360 40.900 122.860 ;
        RECT 40.560 115.380 40.790 122.360 ;
        RECT 44.980 117.110 46.260 129.080 ;
        RECT 48.740 123.890 49.020 124.010 ;
        RECT 48.740 123.390 49.070 123.890 ;
        RECT 44.980 117.030 46.280 117.110 ;
        RECT 44.970 116.730 46.280 117.030 ;
        RECT 41.750 116.080 42.050 116.400 ;
        RECT 40.430 115.370 40.790 115.380 ;
        RECT 40.400 114.520 40.790 115.370 ;
        RECT 40.430 114.510 40.790 114.520 ;
        RECT 40.560 112.820 40.790 114.510 ;
        RECT 41.780 112.820 42.010 116.080 ;
        RECT 48.060 115.530 48.490 115.870 ;
        RECT 48.300 112.860 48.490 115.530 ;
        RECT 48.740 112.770 49.020 123.390 ;
        RECT 50.440 118.630 50.700 118.950 ;
        RECT 49.550 117.760 49.810 118.080 ;
        RECT 49.580 114.040 49.770 117.760 ;
        RECT 50.460 114.040 50.680 118.630 ;
        RECT 52.430 115.410 52.770 131.630 ;
        RECT 72.840 130.230 76.070 132.100 ;
        RECT 81.770 130.430 81.960 132.370 ;
        RECT 100.730 132.180 104.680 133.640 ;
        RECT 113.660 133.290 114.220 133.790 ;
        RECT 117.490 133.370 118.210 139.040 ;
        RECT 118.960 139.770 133.250 140.330 ;
        RECT 144.180 140.160 144.710 141.060 ;
        RECT 145.820 141.000 148.190 141.630 ;
        RECT 118.960 135.470 142.310 139.770 ;
        RECT 145.850 139.040 146.800 141.000 ;
        RECT 147.550 140.980 148.130 141.000 ;
        RECT 157.930 140.340 161.840 141.800 ;
        RECT 169.160 141.150 173.290 141.550 ;
        RECT 169.160 141.060 173.300 141.150 ;
        RECT 148.220 140.330 161.840 140.340 ;
        RECT 143.080 138.350 143.650 138.360 ;
        RECT 118.960 135.190 133.250 135.470 ;
        RECT 129.340 133.640 133.250 135.190 ;
        RECT 143.080 134.930 143.700 138.350 ;
        RECT 143.080 134.920 143.650 134.930 ;
        RECT 113.670 133.070 114.220 133.290 ;
        RECT 129.320 132.870 133.270 133.640 ;
        RECT 142.250 133.290 142.810 133.790 ;
        RECT 146.080 133.370 146.800 139.040 ;
        RECT 147.550 139.770 161.840 140.330 ;
        RECT 172.770 140.160 173.300 141.060 ;
        RECT 174.410 141.000 176.780 141.630 ;
        RECT 147.550 135.470 170.900 139.770 ;
        RECT 174.440 139.040 175.390 141.000 ;
        RECT 176.140 140.980 176.720 141.000 ;
        RECT 186.520 140.340 190.430 141.800 ;
        RECT 197.750 141.150 201.880 141.550 ;
        RECT 197.750 141.060 201.890 141.150 ;
        RECT 176.810 140.330 190.430 140.340 ;
        RECT 171.670 138.350 172.240 138.360 ;
        RECT 147.550 135.190 161.840 135.470 ;
        RECT 157.930 133.640 161.840 135.190 ;
        RECT 171.670 134.930 172.290 138.350 ;
        RECT 171.670 134.920 172.240 134.930 ;
        RECT 142.260 133.070 142.810 133.290 ;
        RECT 100.670 132.100 104.680 132.180 ;
        RECT 129.330 132.100 133.280 132.870 ;
        RECT 157.910 132.100 161.860 133.640 ;
        RECT 170.840 133.290 171.400 133.790 ;
        RECT 174.670 133.370 175.390 139.040 ;
        RECT 176.140 139.770 190.430 140.330 ;
        RECT 201.360 140.160 201.890 141.060 ;
        RECT 176.140 135.470 199.490 139.770 ;
        RECT 200.260 138.350 200.830 138.360 ;
        RECT 176.140 135.190 190.430 135.470 ;
        RECT 186.520 133.640 190.430 135.190 ;
        RECT 200.260 134.930 200.880 138.350 ;
        RECT 200.260 134.920 200.830 134.930 ;
        RECT 170.850 133.070 171.400 133.290 ;
        RECT 186.500 132.100 190.450 133.640 ;
        RECT 199.430 133.290 199.990 133.790 ;
        RECT 199.440 133.070 199.990 133.290 ;
        RECT 100.670 131.900 104.660 132.100 ;
        RECT 100.650 131.700 104.660 131.900 ;
        RECT 81.770 130.240 81.980 130.430 ;
        RECT 72.830 129.110 76.070 130.230 ;
        RECT 56.930 128.170 57.300 128.180 ;
        RECT 56.880 127.720 57.380 128.170 ;
        RECT 53.080 119.310 53.400 119.680 ;
        RECT 53.100 115.470 53.370 119.310 ;
        RECT 52.380 115.330 52.770 115.410 ;
        RECT 52.370 114.560 52.770 115.330 ;
        RECT 52.380 114.490 52.770 114.560 ;
        RECT 49.410 113.350 50.090 114.040 ;
        RECT 50.450 113.350 51.130 114.040 ;
        RECT 52.430 112.710 52.770 114.490 ;
        RECT 52.820 114.820 52.980 115.470 ;
        RECT 52.820 114.270 53.090 114.820 ;
        RECT 52.810 114.220 53.090 114.270 ;
        RECT 52.810 114.130 52.980 114.220 ;
        RECT 52.820 110.840 52.980 114.130 ;
        RECT 53.100 113.980 53.420 115.470 ;
        RECT 55.100 115.100 55.310 115.470 ;
        RECT 54.630 114.650 54.940 115.090 ;
        RECT 55.090 114.810 55.320 115.100 ;
        RECT 53.100 113.930 53.440 113.980 ;
        RECT 53.100 113.430 53.780 113.930 ;
        RECT 53.100 112.780 53.390 113.430 ;
        RECT 54.230 113.120 54.550 113.440 ;
        RECT 55.100 113.110 55.310 114.810 ;
        RECT 55.570 114.540 55.760 115.470 ;
        RECT 55.560 114.250 55.790 114.540 ;
        RECT 53.230 111.430 53.390 112.780 ;
        RECT 53.580 112.610 53.820 113.030 ;
        RECT 55.090 112.820 55.320 113.110 ;
        RECT 55.100 112.680 55.310 112.820 ;
        RECT 53.550 112.290 53.820 112.610 ;
        RECT 53.580 111.860 53.820 112.290 ;
        RECT 55.570 112.220 55.760 114.250 ;
        RECT 55.980 112.750 56.190 115.470 ;
        RECT 55.950 112.240 56.190 112.750 ;
        RECT 55.120 112.040 55.310 112.170 ;
        RECT 55.100 111.750 55.330 112.040 ;
        RECT 55.560 111.930 55.790 112.220 ;
        RECT 54.220 111.430 54.540 111.750 ;
        RECT 53.200 111.190 53.430 111.430 ;
        RECT 53.190 111.180 53.430 111.190 ;
        RECT 53.190 110.910 53.440 111.180 ;
        RECT 53.200 110.880 53.420 110.910 ;
        RECT 34.040 109.310 34.380 109.360 ;
        RECT 34.040 109.290 34.600 109.310 ;
        RECT 33.920 109.120 34.600 109.290 ;
        RECT 34.040 109.080 34.600 109.120 ;
        RECT 34.040 109.040 34.380 109.080 ;
        RECT 35.250 108.400 35.920 109.470 ;
        RECT 35.250 107.860 35.530 108.400 ;
        RECT 35.680 107.860 35.910 108.400 ;
        RECT 34.040 107.180 34.380 107.220 ;
        RECT 34.040 107.140 34.600 107.180 ;
        RECT 33.550 106.930 33.780 107.010 ;
        RECT 33.920 106.970 34.600 107.140 ;
        RECT 34.040 106.950 34.600 106.970 ;
        RECT 34.040 106.900 34.380 106.950 ;
        RECT 34.770 106.930 35.000 107.010 ;
        RECT 35.250 106.790 35.920 107.860 ;
        RECT 37.060 106.860 38.500 107.020 ;
        RECT 40.560 106.930 40.790 107.020 ;
        RECT 41.780 106.940 42.010 107.020 ;
        RECT 35.250 106.540 35.530 106.790 ;
        RECT 35.680 106.540 35.910 106.790 ;
        RECT 34.040 106.380 34.380 106.430 ;
        RECT 34.040 106.360 34.600 106.380 ;
        RECT 33.920 106.190 34.600 106.360 ;
        RECT 34.040 106.150 34.600 106.190 ;
        RECT 35.250 106.180 35.920 106.540 ;
        RECT 34.040 106.110 34.380 106.150 ;
        RECT 35.240 106.110 35.920 106.180 ;
        RECT 35.230 105.510 35.920 106.110 ;
        RECT 35.240 105.480 35.920 105.510 ;
        RECT 35.250 105.470 35.920 105.480 ;
        RECT 35.250 104.930 35.530 105.470 ;
        RECT 34.040 104.250 34.380 104.290 ;
        RECT 34.040 104.210 34.600 104.250 ;
        RECT 33.920 104.040 34.600 104.210 ;
        RECT 34.800 104.200 34.970 104.370 ;
        RECT 34.040 104.020 34.600 104.040 ;
        RECT 34.040 103.970 34.380 104.020 ;
        RECT 34.780 103.610 35.100 103.910 ;
        RECT 35.250 103.860 35.920 104.930 ;
        RECT 42.040 104.790 42.460 110.840 ;
        RECT 44.520 104.790 44.750 110.840 ;
        RECT 45.740 109.630 45.970 110.840 ;
        RECT 50.740 110.020 51.050 110.460 ;
        RECT 45.740 108.840 46.000 109.630 ;
        RECT 52.260 109.380 52.450 110.840 ;
        RECT 52.700 110.670 52.980 110.840 ;
        RECT 52.700 110.190 53.090 110.670 ;
        RECT 52.590 110.070 53.090 110.190 ;
        RECT 52.590 109.590 52.980 110.070 ;
        RECT 50.890 109.060 51.210 109.380 ;
        RECT 52.260 109.350 52.480 109.380 ;
        RECT 52.240 109.080 52.490 109.350 ;
        RECT 52.250 109.070 52.490 109.080 ;
        RECT 45.740 106.690 45.970 108.840 ;
        RECT 52.250 108.830 52.480 109.070 ;
        RECT 51.860 108.270 52.100 108.400 ;
        RECT 51.860 107.950 52.120 108.270 ;
        RECT 51.860 107.350 52.120 107.670 ;
        RECT 51.860 107.230 52.100 107.350 ;
        RECT 52.290 107.020 52.450 108.830 ;
        RECT 52.700 107.990 52.980 109.590 ;
        RECT 53.230 109.420 53.420 110.880 ;
        RECT 54.630 109.800 54.940 110.240 ;
        RECT 55.120 110.130 55.310 111.750 ;
        RECT 55.570 110.640 55.760 111.930 ;
        RECT 55.550 110.350 55.780 110.640 ;
        RECT 55.120 109.920 55.350 110.130 ;
        RECT 55.110 109.840 55.350 109.920 ;
        RECT 55.110 109.420 55.340 109.840 ;
        RECT 55.570 109.420 55.760 110.350 ;
        RECT 55.980 109.420 56.190 112.240 ;
        RECT 56.930 111.650 57.300 127.720 ;
        RECT 57.720 124.270 58.180 124.700 ;
        RECT 56.770 111.630 57.370 111.650 ;
        RECT 56.610 111.590 57.370 111.630 ;
        RECT 56.610 111.330 57.300 111.590 ;
        RECT 52.700 107.670 53.060 107.990 ;
        RECT 52.700 107.020 52.980 107.670 ;
        RECT 48.300 106.940 48.490 107.020 ;
        RECT 48.740 106.970 49.020 107.020 ;
        RECT 45.740 105.900 46.000 106.690 ;
        RECT 48.740 106.670 49.060 106.970 ;
        RECT 50.490 106.680 50.810 107.000 ;
        RECT 52.290 106.800 52.980 107.020 ;
        RECT 53.090 106.870 53.370 107.020 ;
        RECT 50.890 106.300 51.210 106.620 ;
        RECT 51.470 106.400 51.790 106.720 ;
        RECT 52.250 106.550 52.980 106.800 ;
        RECT 52.240 106.280 52.980 106.550 ;
        RECT 45.740 104.790 45.970 105.900 ;
        RECT 50.640 105.850 50.960 106.170 ;
        RECT 51.420 105.750 51.740 106.070 ;
        RECT 49.530 105.320 49.850 105.640 ;
        RECT 50.740 105.170 51.050 105.610 ;
        RECT 50.750 105.160 50.960 105.170 ;
        RECT 50.730 104.840 50.990 105.160 ;
        RECT 51.420 104.920 51.740 105.240 ;
        RECT 40.590 104.200 40.760 104.370 ;
        RECT 50.260 104.040 50.580 104.360 ;
        RECT 35.250 103.640 35.530 103.860 ;
        RECT 34.810 103.510 34.980 103.610 ;
        RECT 35.250 102.280 35.470 103.640 ;
        RECT 40.480 103.540 40.800 103.860 ;
        RECT 50.750 103.550 50.960 104.840 ;
        RECT 52.260 104.790 52.980 106.280 ;
        RECT 53.100 105.440 53.370 106.870 ;
        RECT 53.720 106.450 54.040 106.770 ;
        RECT 53.100 105.150 53.380 105.440 ;
        RECT 51.470 104.270 51.790 104.590 ;
        RECT 38.140 102.880 38.300 103.530 ;
        RECT 38.140 102.330 38.410 102.880 ;
        RECT 38.130 102.280 38.410 102.330 ;
        RECT 38.550 102.540 38.740 103.530 ;
        RECT 38.950 102.850 39.110 103.530 ;
        RECT 40.590 103.520 40.760 103.540 ;
        RECT 38.910 102.830 39.110 102.850 ;
        RECT 39.930 102.840 40.250 103.160 ;
        RECT 38.900 102.590 39.130 102.830 ;
        RECT 38.550 102.420 38.720 102.540 ;
        RECT 35.250 102.190 35.600 102.280 ;
        RECT 38.130 102.190 38.300 102.280 ;
        RECT 35.250 101.970 35.760 102.190 ;
        RECT 38.140 101.830 38.300 102.190 ;
        RECT 38.130 101.740 38.300 101.830 ;
        RECT 38.130 101.690 38.410 101.740 ;
        RECT 38.140 101.390 38.410 101.690 ;
        RECT 38.550 101.600 38.710 102.420 ;
        RECT 38.910 102.370 39.110 102.590 ;
        RECT 38.950 101.650 39.110 102.370 ;
        RECT 39.930 102.290 40.250 102.610 ;
        RECT 40.890 102.370 41.130 103.530 ;
        RECT 38.550 101.480 38.720 101.600 ;
        RECT 26.540 100.140 26.820 101.250 ;
        RECT 27.070 100.560 27.260 101.160 ;
        RECT 29.070 100.720 29.460 100.740 ;
        RECT 29.060 100.630 29.460 100.720 ;
        RECT 27.070 100.370 28.700 100.560 ;
        RECT 26.540 99.860 28.260 100.140 ;
        RECT 27.980 99.630 28.260 99.860 ;
        RECT 28.510 99.590 28.700 100.370 ;
        RECT 28.910 100.380 29.460 100.630 ;
        RECT 28.910 100.360 29.450 100.380 ;
        RECT 28.910 99.510 29.070 100.360 ;
        RECT 33.030 100.290 33.410 100.310 ;
        RECT 33.550 100.290 33.780 101.200 ;
        RECT 33.030 100.060 33.780 100.290 ;
        RECT 34.770 100.200 35.000 101.200 ;
        RECT 38.080 100.210 38.500 101.390 ;
        RECT 38.550 100.620 38.740 101.480 ;
        RECT 38.910 101.430 39.110 101.650 ;
        RECT 38.900 101.190 39.130 101.430 ;
        RECT 39.930 101.410 40.250 101.730 ;
        RECT 40.880 101.710 41.150 102.370 ;
        RECT 38.910 101.170 39.110 101.190 ;
        RECT 38.520 100.390 38.760 100.620 ;
        RECT 31.000 99.400 31.190 99.620 ;
        RECT 10.820 98.620 11.230 98.950 ;
        RECT 11.560 98.640 11.800 99.040 ;
        RECT 14.500 98.640 14.810 99.040 ;
        RECT 11.370 98.590 11.800 98.640 ;
        RECT 10.820 97.070 11.230 97.400 ;
        RECT 10.820 95.520 11.230 95.850 ;
        RECT 10.820 93.970 11.230 94.300 ;
        RECT 11.560 93.660 11.800 98.590 ;
        RECT 14.310 98.580 14.810 98.640 ;
        RECT 12.980 98.090 13.180 98.110 ;
        RECT 12.980 97.800 13.330 98.090 ;
        RECT 12.980 96.540 13.180 96.560 ;
        RECT 12.980 96.250 13.330 96.540 ;
        RECT 12.980 94.990 13.180 95.010 ;
        RECT 12.980 94.700 13.330 94.990 ;
        RECT 14.500 93.730 14.810 98.580 ;
        RECT 15.060 98.510 15.340 98.840 ;
        RECT 18.930 98.640 19.220 99.040 ;
        RECT 30.720 98.910 31.190 99.400 ;
        RECT 31.580 99.260 31.950 99.280 ;
        RECT 31.530 99.000 31.950 99.260 ;
        RECT 31.580 98.990 31.950 99.000 ;
        RECT 18.740 98.590 19.220 98.640 ;
        RECT 17.860 97.690 18.180 97.990 ;
        RECT 15.060 96.960 15.340 97.290 ;
        RECT 17.860 96.140 18.180 96.440 ;
        RECT 15.060 95.410 15.340 95.740 ;
        RECT 17.860 94.590 18.180 94.890 ;
        RECT 15.060 93.860 15.340 94.190 ;
        RECT 11.560 92.800 11.910 93.660 ;
        RECT 12.980 93.440 13.180 93.460 ;
        RECT 12.980 93.150 13.330 93.440 ;
        RECT 14.500 92.800 14.920 93.730 ;
        RECT 18.930 93.710 19.220 98.590 ;
        RECT 30.540 98.470 30.860 98.750 ;
        RECT 31.000 98.650 31.190 98.910 ;
        RECT 31.000 98.360 31.230 98.650 ;
        RECT 31.000 97.760 31.190 98.360 ;
        RECT 30.540 97.370 30.860 97.650 ;
        RECT 31.000 97.470 31.230 97.760 ;
        RECT 31.000 97.210 31.190 97.470 ;
        RECT 30.720 96.720 31.190 97.210 ;
        RECT 31.580 97.120 31.950 97.130 ;
        RECT 31.530 96.860 31.950 97.120 ;
        RECT 31.580 96.840 31.950 96.860 ;
        RECT 31.000 96.470 31.190 96.720 ;
        RECT 30.720 95.980 31.190 96.470 ;
        RECT 31.580 96.330 31.950 96.350 ;
        RECT 31.530 96.070 31.950 96.330 ;
        RECT 31.580 96.060 31.950 96.070 ;
        RECT 30.540 95.540 30.860 95.820 ;
        RECT 31.000 95.720 31.190 95.980 ;
        RECT 31.000 95.430 31.230 95.720 ;
        RECT 31.000 94.830 31.190 95.430 ;
        RECT 30.540 94.440 30.860 94.720 ;
        RECT 31.000 94.540 31.230 94.830 ;
        RECT 31.000 94.280 31.190 94.540 ;
        RECT 30.720 93.790 31.190 94.280 ;
        RECT 31.580 94.190 31.950 94.200 ;
        RECT 31.530 93.930 31.950 94.190 ;
        RECT 31.580 93.910 31.950 93.930 ;
        RECT 17.860 93.040 18.180 93.340 ;
        RECT 18.930 92.800 19.330 93.710 ;
        RECT 11.370 92.400 11.610 92.450 ;
        RECT 11.670 89.890 11.910 92.800 ;
        RECT 14.610 92.470 14.920 92.800 ;
        RECT 14.310 92.400 14.920 92.470 ;
        RECT 18.740 92.400 19.030 92.450 ;
        RECT 14.610 89.890 14.920 92.400 ;
        RECT 19.040 89.890 19.330 92.800 ;
        RECT 20.500 89.620 20.690 93.710 ;
        RECT 21.810 92.670 22.040 93.750 ;
        RECT 21.720 92.190 22.050 92.670 ;
        RECT 21.810 89.580 22.040 92.190 ;
        RECT 24.780 89.790 25.030 93.770 ;
        RECT 25.440 93.060 25.600 93.710 ;
        RECT 25.440 92.510 25.710 93.060 ;
        RECT 25.430 92.460 25.710 92.510 ;
        RECT 25.850 92.720 26.040 93.710 ;
        RECT 26.250 93.030 26.410 93.710 ;
        RECT 26.210 93.010 26.410 93.030 ;
        RECT 27.230 93.020 27.550 93.340 ;
        RECT 26.200 92.770 26.430 93.010 ;
        RECT 25.850 92.600 26.020 92.720 ;
        RECT 25.430 92.370 25.600 92.460 ;
        RECT 25.440 92.010 25.600 92.370 ;
        RECT 25.430 91.920 25.600 92.010 ;
        RECT 25.430 91.870 25.710 91.920 ;
        RECT 25.440 91.320 25.710 91.870 ;
        RECT 25.850 91.780 26.010 92.600 ;
        RECT 26.210 92.550 26.410 92.770 ;
        RECT 26.250 91.830 26.410 92.550 ;
        RECT 27.230 92.470 27.550 92.790 ;
        RECT 25.850 91.660 26.020 91.780 ;
        RECT 25.440 90.050 25.600 91.320 ;
        RECT 25.850 90.800 26.040 91.660 ;
        RECT 26.210 91.610 26.410 91.830 ;
        RECT 26.200 91.370 26.430 91.610 ;
        RECT 27.230 91.590 27.550 91.910 ;
        RECT 26.210 91.350 26.410 91.370 ;
        RECT 25.820 90.570 26.060 90.800 ;
        RECT 25.440 89.500 25.710 90.050 ;
        RECT 25.430 89.450 25.710 89.500 ;
        RECT 25.850 89.710 26.040 90.570 ;
        RECT 26.250 90.020 26.410 91.350 ;
        RECT 27.230 91.040 27.550 91.360 ;
        RECT 26.210 90.000 26.410 90.020 ;
        RECT 27.230 90.010 27.550 90.330 ;
        RECT 26.200 89.760 26.430 90.000 ;
        RECT 25.850 89.590 26.020 89.710 ;
        RECT 25.430 89.360 25.600 89.450 ;
        RECT 10.820 88.850 11.230 89.180 ;
        RECT 11.560 88.870 11.800 89.270 ;
        RECT 14.500 88.870 14.810 89.270 ;
        RECT 11.370 88.820 11.800 88.870 ;
        RECT 10.820 87.300 11.230 87.630 ;
        RECT 10.820 85.750 11.230 86.080 ;
        RECT 10.820 84.200 11.230 84.530 ;
        RECT 11.560 83.890 11.800 88.820 ;
        RECT 14.310 88.810 14.810 88.870 ;
        RECT 12.980 88.320 13.180 88.340 ;
        RECT 12.980 88.030 13.330 88.320 ;
        RECT 12.980 86.770 13.180 86.790 ;
        RECT 12.980 86.480 13.330 86.770 ;
        RECT 12.980 85.220 13.180 85.240 ;
        RECT 12.980 84.930 13.330 85.220 ;
        RECT 14.500 83.960 14.810 88.810 ;
        RECT 15.060 88.740 15.340 89.070 ;
        RECT 18.930 88.870 19.220 89.270 ;
        RECT 25.440 89.010 25.600 89.360 ;
        RECT 25.430 88.920 25.600 89.010 ;
        RECT 25.430 88.870 25.710 88.920 ;
        RECT 18.740 88.820 19.220 88.870 ;
        RECT 17.860 87.920 18.180 88.220 ;
        RECT 15.060 87.190 15.340 87.520 ;
        RECT 17.860 86.370 18.180 86.670 ;
        RECT 15.060 85.640 15.340 85.970 ;
        RECT 17.860 84.820 18.180 85.120 ;
        RECT 15.060 84.090 15.340 84.420 ;
        RECT 11.560 83.030 11.910 83.890 ;
        RECT 12.980 83.670 13.180 83.690 ;
        RECT 12.980 83.380 13.330 83.670 ;
        RECT 14.500 83.030 14.920 83.960 ;
        RECT 18.930 83.940 19.220 88.820 ;
        RECT 25.440 88.320 25.710 88.870 ;
        RECT 25.850 88.780 26.010 89.590 ;
        RECT 26.210 89.540 26.410 89.760 ;
        RECT 26.250 88.830 26.410 89.540 ;
        RECT 27.230 89.460 27.550 89.780 ;
        RECT 28.100 89.730 28.260 93.780 ;
        RECT 28.310 89.890 28.560 93.710 ;
        RECT 30.370 91.790 30.750 93.710 ;
        RECT 30.850 93.570 31.190 93.790 ;
        RECT 32.310 93.710 32.540 99.620 ;
        RECT 33.030 99.290 33.410 100.060 ;
        RECT 34.770 99.900 35.020 100.200 ;
        RECT 34.780 99.430 35.020 99.900 ;
        RECT 38.080 99.820 38.540 100.210 ;
        RECT 35.280 99.400 35.530 99.620 ;
        RECT 34.040 99.240 34.380 99.290 ;
        RECT 34.040 99.220 34.600 99.240 ;
        RECT 33.920 99.050 34.600 99.220 ;
        RECT 34.040 99.010 34.600 99.050 ;
        RECT 34.040 98.970 34.380 99.010 ;
        RECT 35.280 98.330 35.920 99.400 ;
        RECT 38.140 99.320 38.540 99.820 ;
        RECT 38.130 99.270 38.540 99.320 ;
        RECT 38.550 99.530 38.740 100.390 ;
        RECT 38.950 99.840 39.110 101.170 ;
        RECT 39.930 100.860 40.250 101.180 ;
        RECT 40.480 101.030 40.800 101.330 ;
        RECT 40.560 100.220 40.790 101.030 ;
        RECT 38.910 99.820 39.110 99.840 ;
        RECT 39.930 99.830 40.250 100.150 ;
        RECT 40.560 99.870 40.820 100.220 ;
        RECT 38.900 99.580 39.130 99.820 ;
        RECT 40.580 99.710 40.820 99.870 ;
        RECT 40.890 99.710 41.130 101.710 ;
        RECT 43.070 101.610 43.450 103.530 ;
        RECT 44.820 102.350 45.060 103.530 ;
        RECT 44.810 101.690 45.070 102.350 ;
        RECT 41.780 100.310 42.010 101.200 ;
        RECT 41.760 99.930 42.570 100.310 ;
        RECT 38.550 99.410 38.720 99.530 ;
        RECT 38.130 99.180 38.300 99.270 ;
        RECT 38.140 98.830 38.300 99.180 ;
        RECT 38.130 98.740 38.300 98.830 ;
        RECT 38.130 98.690 38.410 98.740 ;
        RECT 35.280 97.790 35.530 98.330 ;
        RECT 38.140 98.140 38.410 98.690 ;
        RECT 38.550 98.600 38.710 99.410 ;
        RECT 38.910 99.360 39.110 99.580 ;
        RECT 38.950 98.650 39.110 99.360 ;
        RECT 39.930 99.280 40.250 99.600 ;
        RECT 40.580 99.430 41.130 99.710 ;
        RECT 41.190 99.660 41.380 99.710 ;
        RECT 41.590 99.660 41.750 99.710 ;
        RECT 40.620 99.370 41.130 99.430 ;
        RECT 40.890 99.120 41.130 99.370 ;
        RECT 42.190 99.290 42.570 99.930 ;
        RECT 43.070 99.750 43.460 101.610 ;
        RECT 40.880 98.800 41.140 99.120 ;
        RECT 38.550 98.480 38.720 98.600 ;
        RECT 34.040 97.110 34.380 97.150 ;
        RECT 34.040 97.070 34.600 97.110 ;
        RECT 33.920 96.900 34.600 97.070 ;
        RECT 34.040 96.880 34.600 96.900 ;
        RECT 34.040 96.830 34.380 96.880 ;
        RECT 35.280 96.720 35.920 97.790 ;
        RECT 38.140 97.490 38.300 98.140 ;
        RECT 38.550 97.490 38.740 98.480 ;
        RECT 38.910 98.430 39.110 98.650 ;
        RECT 38.900 98.190 39.130 98.430 ;
        RECT 39.930 98.410 40.250 98.730 ;
        RECT 38.910 98.170 39.110 98.190 ;
        RECT 38.950 97.490 39.110 98.170 ;
        RECT 39.930 97.860 40.250 98.180 ;
        RECT 40.890 97.480 41.130 98.800 ;
        RECT 43.070 97.480 43.450 99.750 ;
        RECT 43.530 99.620 43.770 99.710 ;
        RECT 44.820 99.080 45.060 101.690 ;
        RECT 47.100 100.180 47.500 103.530 ;
        RECT 50.730 103.260 50.960 103.550 ;
        RECT 51.470 103.440 51.790 103.760 ;
        RECT 51.420 102.790 51.740 103.110 ;
        RECT 51.420 101.960 51.740 102.280 ;
        RECT 48.300 100.180 48.490 101.160 ;
        RECT 46.470 99.810 46.750 100.130 ;
        RECT 46.900 99.990 48.490 100.180 ;
        RECT 45.710 99.610 46.090 99.710 ;
        RECT 46.530 99.510 46.690 99.810 ;
        RECT 46.900 99.640 47.090 99.990 ;
        RECT 47.100 99.800 47.500 99.990 ;
        RECT 48.740 99.800 49.020 101.250 ;
        RECT 50.920 101.170 51.250 101.460 ;
        RECT 51.470 101.310 51.790 101.630 ;
        RECT 52.430 101.170 52.770 104.790 ;
        RECT 50.910 101.030 52.770 101.170 ;
        RECT 52.430 100.970 52.770 101.030 ;
        RECT 53.100 102.850 53.370 105.150 ;
        RECT 53.770 104.230 54.090 104.550 ;
        RECT 53.760 103.530 54.080 103.830 ;
        RECT 53.460 103.510 54.080 103.530 ;
        RECT 53.100 102.560 53.380 102.850 ;
        RECT 53.100 100.970 53.370 102.560 ;
        RECT 53.460 101.580 53.860 103.510 ;
        RECT 55.900 102.350 56.140 103.530 ;
        RECT 55.890 101.690 56.150 102.350 ;
        RECT 53.460 101.260 54.000 101.580 ;
        RECT 47.100 99.520 49.020 99.800 ;
        RECT 53.460 99.710 53.860 101.260 ;
        RECT 49.740 99.580 50.140 99.710 ;
        RECT 50.820 99.610 51.220 99.710 ;
        RECT 53.260 99.660 53.860 99.710 ;
        RECT 44.810 98.760 45.070 99.080 ;
        RECT 44.820 97.480 45.060 98.760 ;
        RECT 47.100 97.480 47.500 99.520 ;
        RECT 50.140 99.350 50.820 99.570 ;
        RECT 53.460 97.480 53.860 99.660 ;
        RECT 54.870 99.610 55.250 99.710 ;
        RECT 55.900 99.080 56.140 101.690 ;
        RECT 56.930 100.810 57.300 111.330 ;
        RECT 57.740 103.530 58.110 124.270 ;
        RECT 58.490 119.560 58.940 119.990 ;
        RECT 57.510 101.610 58.110 103.530 ;
        RECT 56.900 100.350 57.350 100.810 ;
        RECT 56.930 100.310 57.300 100.350 ;
        RECT 57.500 100.220 58.110 101.610 ;
        RECT 57.500 99.760 58.150 100.220 ;
        RECT 57.500 99.750 58.110 99.760 ;
        RECT 57.510 99.710 58.110 99.750 ;
        RECT 57.190 99.640 57.430 99.710 ;
        RECT 55.890 98.760 56.150 99.080 ;
        RECT 55.900 97.480 56.140 98.760 ;
        RECT 57.510 97.480 57.890 99.710 ;
        RECT 58.510 97.870 58.880 119.560 ;
        RECT 65.060 118.510 65.640 119.070 ;
        RECT 61.850 116.940 62.410 117.590 ;
        RECT 62.800 117.430 63.360 118.010 ;
        RECT 63.880 117.890 64.440 118.480 ;
        RECT 59.380 114.480 59.810 114.920 ;
        RECT 59.050 111.540 59.260 111.650 ;
        RECT 59.060 105.610 59.290 105.730 ;
        RECT 59.390 99.710 59.760 114.480 ;
        RECT 60.930 111.650 61.160 115.470 ;
        RECT 59.930 111.590 60.140 111.650 ;
        RECT 60.930 111.580 61.190 111.650 ;
        RECT 60.930 109.420 61.160 111.580 ;
        RECT 61.870 103.530 62.370 116.940 ;
        RECT 62.800 115.470 63.300 117.430 ;
        RECT 62.800 109.420 63.640 115.470 ;
        RECT 62.800 103.530 63.300 109.420 ;
        RECT 59.830 102.370 60.070 103.530 ;
        RECT 60.710 102.840 61.030 103.160 ;
        RECT 61.850 102.830 62.410 103.530 ;
        RECT 62.660 102.880 63.300 103.530 ;
        RECT 59.810 101.710 60.080 102.370 ;
        RECT 60.710 102.290 61.030 102.610 ;
        RECT 61.830 102.590 62.410 102.830 ;
        RECT 59.830 99.710 60.070 101.710 ;
        RECT 60.710 101.410 61.030 101.730 ;
        RECT 61.850 101.430 62.410 102.590 ;
        RECT 62.550 102.280 63.300 102.880 ;
        RECT 62.660 101.740 63.300 102.280 ;
        RECT 61.830 101.190 62.410 101.430 ;
        RECT 60.710 100.860 61.030 101.180 ;
        RECT 61.850 100.620 62.410 101.190 ;
        RECT 62.550 101.140 63.300 101.740 ;
        RECT 61.850 100.390 62.440 100.620 ;
        RECT 60.710 99.830 61.030 100.150 ;
        RECT 61.850 99.820 62.410 100.390 ;
        RECT 62.660 99.870 63.300 101.140 ;
        RECT 59.210 99.660 59.370 99.710 ;
        RECT 59.390 99.660 59.770 99.710 ;
        RECT 59.830 99.670 60.180 99.710 ;
        RECT 58.480 97.860 58.880 97.870 ;
        RECT 58.470 97.440 58.890 97.860 ;
        RECT 58.510 97.430 58.880 97.440 ;
        RECT 35.280 96.470 35.530 96.720 ;
        RECT 34.040 96.310 34.380 96.360 ;
        RECT 34.040 96.290 34.600 96.310 ;
        RECT 33.920 96.120 34.600 96.290 ;
        RECT 34.040 96.080 34.600 96.120 ;
        RECT 34.040 96.040 34.380 96.080 ;
        RECT 35.280 95.400 35.920 96.470 ;
        RECT 35.280 94.860 35.530 95.400 ;
        RECT 34.040 94.180 34.380 94.220 ;
        RECT 34.040 94.140 34.600 94.180 ;
        RECT 32.310 93.570 32.590 93.710 ;
        RECT 30.370 89.930 30.760 91.790 ;
        RECT 30.850 90.140 31.090 93.570 ;
        RECT 28.310 89.820 28.700 89.890 ;
        RECT 28.910 89.820 29.070 89.890 ;
        RECT 28.310 89.270 28.560 89.820 ;
        RECT 30.370 89.640 30.750 89.930 ;
        RECT 30.830 89.890 31.220 90.140 ;
        RECT 30.970 89.640 31.220 89.890 ;
        RECT 32.320 89.860 32.590 93.570 ;
        RECT 28.290 89.240 28.570 89.270 ;
        RECT 28.280 88.960 28.580 89.240 ;
        RECT 30.370 89.150 31.190 89.640 ;
        RECT 31.580 89.500 31.950 89.520 ;
        RECT 31.530 89.240 31.950 89.500 ;
        RECT 32.310 89.240 32.590 89.860 ;
        RECT 33.030 89.510 33.410 94.000 ;
        RECT 33.920 93.970 34.600 94.140 ;
        RECT 34.040 93.950 34.600 93.970 ;
        RECT 34.040 93.900 34.380 93.950 ;
        RECT 34.780 93.710 35.020 93.860 ;
        RECT 34.400 90.120 35.020 93.710 ;
        RECT 35.280 93.790 35.920 94.860 ;
        RECT 35.280 93.570 35.530 93.790 ;
        RECT 34.400 89.850 35.250 90.120 ;
        RECT 34.040 89.480 34.380 89.530 ;
        RECT 34.400 89.480 34.800 89.850 ;
        RECT 34.980 89.620 35.250 89.850 ;
        RECT 35.280 89.640 35.530 89.860 ;
        RECT 34.040 89.460 34.800 89.480 ;
        RECT 33.920 89.290 34.800 89.460 ;
        RECT 34.040 89.250 34.800 89.290 ;
        RECT 31.580 89.230 31.950 89.240 ;
        RECT 30.370 88.990 30.750 89.150 ;
        RECT 28.290 88.940 28.570 88.960 ;
        RECT 26.210 88.800 26.410 88.830 ;
        RECT 25.850 88.660 26.020 88.780 ;
        RECT 25.440 87.670 25.600 88.320 ;
        RECT 25.850 87.670 26.040 88.660 ;
        RECT 26.130 88.460 26.450 88.800 ;
        RECT 27.230 88.590 27.550 88.910 ;
        RECT 26.200 88.370 26.430 88.460 ;
        RECT 17.860 83.270 18.180 83.570 ;
        RECT 18.930 83.320 19.330 83.940 ;
        RECT 19.540 83.340 19.880 83.660 ;
        RECT 18.930 83.030 19.360 83.320 ;
        RECT 11.370 82.630 11.610 82.680 ;
        RECT 11.670 71.260 11.910 83.030 ;
        RECT 14.610 82.810 14.920 83.030 ;
        RECT 19.010 82.970 19.360 83.030 ;
        RECT 14.570 82.700 14.940 82.810 ;
        RECT 14.310 82.630 14.940 82.700 ;
        RECT 18.740 82.630 19.030 82.680 ;
        RECT 14.570 82.480 14.940 82.630 ;
        RECT 19.040 82.510 19.330 82.970 ;
        RECT 19.540 82.730 19.790 83.340 ;
        RECT 20.500 82.750 20.690 83.950 ;
        RECT 24.780 83.280 25.030 84.010 ;
        RECT 26.210 83.700 26.420 88.370 ;
        RECT 27.230 88.040 27.550 88.360 ;
        RECT 27.240 87.960 27.500 88.040 ;
        RECT 27.230 87.760 27.500 87.960 ;
        RECT 27.230 87.070 27.440 87.760 ;
        RECT 28.310 87.660 28.560 88.940 ;
        RECT 30.370 88.710 30.860 88.990 ;
        RECT 31.000 88.890 31.190 89.150 ;
        RECT 32.300 88.930 32.610 89.240 ;
        RECT 34.040 89.210 34.380 89.250 ;
        RECT 30.370 88.580 30.750 88.710 ;
        RECT 31.000 88.600 31.230 88.890 ;
        RECT 30.370 88.260 30.770 88.580 ;
        RECT 30.370 87.890 30.750 88.260 ;
        RECT 31.000 88.000 31.190 88.600 ;
        RECT 30.370 87.660 30.860 87.890 ;
        RECT 30.540 87.610 30.860 87.660 ;
        RECT 31.000 87.710 31.230 88.000 ;
        RECT 31.000 87.450 31.190 87.710 ;
        RECT 27.220 87.020 27.480 87.070 ;
        RECT 27.220 86.770 27.860 87.020 ;
        RECT 30.720 86.960 31.190 87.450 ;
        RECT 32.310 87.660 32.590 88.930 ;
        RECT 34.400 87.660 34.800 89.250 ;
        RECT 35.280 88.570 35.920 89.640 ;
        RECT 37.060 89.490 37.460 94.020 ;
        RECT 40.580 93.720 40.820 93.860 ;
        RECT 40.580 93.660 40.940 93.720 ;
        RECT 41.190 93.670 41.380 93.730 ;
        RECT 41.590 93.670 41.750 93.730 ;
        RECT 43.530 93.660 43.770 93.740 ;
        RECT 45.710 93.660 46.090 93.750 ;
        RECT 47.460 93.660 47.700 93.730 ;
        RECT 49.740 93.660 50.140 93.780 ;
        RECT 50.820 93.660 51.220 93.780 ;
        RECT 53.260 93.660 53.500 93.730 ;
        RECT 54.870 93.660 55.250 93.810 ;
        RECT 59.390 93.730 59.760 99.660 ;
        RECT 59.830 99.370 60.340 99.670 ;
        RECT 59.830 99.120 60.070 99.370 ;
        RECT 60.710 99.280 61.030 99.600 ;
        RECT 61.830 99.580 62.410 99.820 ;
        RECT 59.820 98.800 60.080 99.120 ;
        RECT 59.830 97.480 60.070 98.800 ;
        RECT 60.710 98.410 61.030 98.730 ;
        RECT 61.850 98.430 62.410 99.580 ;
        RECT 62.550 99.270 63.300 99.870 ;
        RECT 62.660 98.740 63.300 99.270 ;
        RECT 61.830 98.190 62.410 98.430 ;
        RECT 60.710 97.860 61.030 98.180 ;
        RECT 61.850 97.490 62.410 98.190 ;
        RECT 62.550 98.140 63.300 98.740 ;
        RECT 62.660 97.490 63.300 98.140 ;
        RECT 57.190 93.660 57.430 93.720 ;
        RECT 59.210 93.670 59.370 93.730 ;
        RECT 59.390 93.670 59.770 93.730 ;
        RECT 60.020 93.670 60.180 93.730 ;
        RECT 40.580 91.350 40.820 93.660 ;
        RECT 59.390 92.690 59.760 93.670 ;
        RECT 59.350 92.180 59.840 92.690 ;
        RECT 59.390 92.150 59.760 92.180 ;
        RECT 40.580 91.110 41.160 91.350 ;
        RECT 38.580 89.110 38.900 89.430 ;
        RECT 35.280 88.030 35.530 88.570 ;
        RECT 38.730 88.430 39.050 88.750 ;
        RECT 31.580 87.360 31.950 87.370 ;
        RECT 31.530 87.100 31.950 87.360 ;
        RECT 31.580 87.080 31.950 87.100 ;
        RECT 27.220 86.750 27.480 86.770 ;
        RECT 26.750 85.670 27.090 86.010 ;
        RECT 26.790 85.650 27.010 85.670 ;
        RECT 26.180 83.380 26.460 83.700 ;
        RECT 26.790 83.370 26.990 85.650 ;
        RECT 27.140 84.710 27.460 85.030 ;
        RECT 27.250 84.180 27.440 84.190 ;
        RECT 27.190 83.860 27.510 84.180 ;
        RECT 27.250 83.690 27.440 83.860 ;
        RECT 24.750 82.990 25.090 83.280 ;
        RECT 26.750 83.050 27.030 83.370 ;
        RECT 27.210 83.360 27.490 83.690 ;
        RECT 14.610 81.270 14.920 82.480 ;
        RECT 18.470 82.230 19.330 82.510 ;
        RECT 18.390 82.220 19.330 82.230 ;
        RECT 19.490 82.620 19.790 82.730 ;
        RECT 18.390 81.750 18.850 82.220 ;
        RECT 14.560 80.790 14.980 81.270 ;
        RECT 19.490 81.110 19.680 82.620 ;
        RECT 20.440 82.430 20.760 82.750 ;
        RECT 23.120 82.220 23.870 82.410 ;
        RECT 23.370 81.380 23.870 82.220 ;
        RECT 27.680 82.140 27.860 86.770 ;
        RECT 31.000 86.710 31.190 86.960 ;
        RECT 30.720 86.700 31.190 86.710 ;
        RECT 30.510 86.380 31.190 86.700 ;
        RECT 31.580 86.570 31.950 86.590 ;
        RECT 30.510 86.060 30.670 86.380 ;
        RECT 30.720 86.220 31.190 86.380 ;
        RECT 31.530 86.310 31.950 86.570 ;
        RECT 31.580 86.300 31.950 86.310 ;
        RECT 30.510 85.780 30.860 86.060 ;
        RECT 31.000 85.960 31.190 86.220 ;
        RECT 30.510 85.520 30.670 85.780 ;
        RECT 30.350 85.200 30.670 85.520 ;
        RECT 31.000 85.670 31.230 85.960 ;
        RECT 31.000 85.070 31.190 85.670 ;
        RECT 30.540 84.680 30.860 84.960 ;
        RECT 31.000 84.780 31.230 85.070 ;
        RECT 31.000 84.520 31.190 84.780 ;
        RECT 30.720 84.090 31.190 84.520 ;
        RECT 31.580 84.430 31.950 84.440 ;
        RECT 31.530 84.170 31.950 84.430 ;
        RECT 31.580 84.150 31.950 84.170 ;
        RECT 30.720 84.030 31.220 84.090 ;
        RECT 29.000 83.300 29.260 83.330 ;
        RECT 28.980 83.000 29.280 83.300 ;
        RECT 29.000 82.990 29.260 83.000 ;
        RECT 27.680 81.840 28.160 82.140 ;
        RECT 29.010 82.070 29.230 82.990 ;
        RECT 30.970 82.860 31.220 84.030 ;
        RECT 32.310 83.810 32.540 87.660 ;
        RECT 34.040 87.350 34.380 87.390 ;
        RECT 34.040 87.310 34.600 87.350 ;
        RECT 33.920 87.140 34.600 87.310 ;
        RECT 34.040 87.120 34.600 87.140 ;
        RECT 34.040 87.070 34.380 87.120 ;
        RECT 35.280 86.960 35.920 88.030 ;
        RECT 38.730 87.540 39.050 87.860 ;
        RECT 35.280 86.710 35.530 86.960 ;
        RECT 38.580 86.860 38.900 87.180 ;
        RECT 34.040 86.550 34.380 86.600 ;
        RECT 34.040 86.530 34.600 86.550 ;
        RECT 33.920 86.360 34.600 86.530 ;
        RECT 34.040 86.320 34.600 86.360 ;
        RECT 34.040 86.280 34.380 86.320 ;
        RECT 35.280 85.640 35.920 86.710 ;
        RECT 38.580 86.340 38.900 86.660 ;
        RECT 38.730 85.660 39.050 85.980 ;
        RECT 35.280 85.100 35.530 85.640 ;
        RECT 34.040 84.420 34.380 84.460 ;
        RECT 34.040 84.380 34.600 84.420 ;
        RECT 33.920 84.210 34.600 84.380 ;
        RECT 34.040 84.190 34.600 84.210 ;
        RECT 34.040 84.140 34.380 84.190 ;
        RECT 33.030 83.840 33.410 83.940 ;
        RECT 34.980 82.880 35.250 84.110 ;
        RECT 35.280 84.030 35.920 85.100 ;
        RECT 38.730 84.770 39.050 85.090 ;
        RECT 38.580 84.090 38.900 84.410 ;
        RECT 35.280 83.810 35.530 84.030 ;
        RECT 39.660 83.840 39.890 89.890 ;
        RECT 40.920 89.770 41.160 91.110 ;
        RECT 40.920 85.540 41.150 89.770 ;
        RECT 46.040 88.710 46.300 88.770 ;
        RECT 46.030 88.450 46.300 88.710 ;
        RECT 45.520 87.520 45.780 87.840 ;
        RECT 45.050 85.680 45.310 86.000 ;
        RECT 40.880 85.530 41.160 85.540 ;
        RECT 40.880 85.210 41.180 85.530 ;
        RECT 37.800 83.310 38.230 83.710 ;
        RECT 30.960 82.600 31.280 82.860 ;
        RECT 34.980 82.570 35.330 82.880 ;
        RECT 27.760 81.730 28.160 81.840 ;
        RECT 28.950 81.670 29.290 82.070 ;
        RECT 29.010 81.590 29.230 81.670 ;
        RECT 32.960 81.400 33.900 82.330 ;
        RECT 37.840 81.520 38.190 83.310 ;
        RECT 39.660 82.750 39.880 83.840 ;
        RECT 40.920 83.350 41.150 85.210 ;
        RECT 44.550 84.750 44.810 85.070 ;
        RECT 40.920 83.120 44.130 83.350 ;
        RECT 40.920 83.110 41.150 83.120 ;
        RECT 39.370 82.510 39.880 82.750 ;
        RECT 19.050 80.790 19.680 81.110 ;
        RECT 22.880 81.060 23.120 81.380 ;
        RECT 24.120 81.060 24.360 81.380 ;
        RECT 32.690 81.080 32.930 81.400 ;
        RECT 33.930 81.080 34.170 81.400 ;
        RECT 39.370 81.260 39.600 82.510 ;
        RECT 43.900 82.150 44.130 83.120 ;
        RECT 43.850 81.750 44.160 82.150 ;
        RECT 39.260 80.820 39.720 81.260 ;
        RECT 19.050 80.690 19.490 80.790 ;
        RECT 22.880 79.720 23.120 80.040 ;
        RECT 24.120 79.710 24.360 80.030 ;
        RECT 32.690 79.740 32.930 80.060 ;
        RECT 33.930 79.730 34.170 80.050 ;
        RECT 43.900 78.580 44.130 81.750 ;
        RECT 43.770 78.360 44.130 78.580 ;
        RECT 22.480 78.090 22.740 78.290 ;
        RECT 24.500 78.090 24.760 78.290 ;
        RECT 19.210 77.570 19.530 77.890 ;
        RECT 20.300 77.570 20.620 77.890 ;
        RECT 21.400 77.560 21.720 77.880 ;
        RECT 22.480 77.280 22.790 78.090 ;
        RECT 24.450 77.280 24.760 78.090 ;
        RECT 32.290 78.120 32.550 78.320 ;
        RECT 34.310 78.120 34.570 78.320 ;
        RECT 43.570 78.130 44.130 78.360 ;
        RECT 43.570 78.120 44.110 78.130 ;
        RECT 25.520 77.560 25.840 77.880 ;
        RECT 26.620 77.570 26.940 77.890 ;
        RECT 27.710 77.570 28.030 77.890 ;
        RECT 29.020 77.600 29.340 77.920 ;
        RECT 30.110 77.600 30.430 77.920 ;
        RECT 31.210 77.590 31.530 77.910 ;
        RECT 32.290 77.310 32.600 78.120 ;
        RECT 34.260 77.310 34.570 78.120 ;
        RECT 35.330 77.590 35.650 77.910 ;
        RECT 36.430 77.600 36.750 77.920 ;
        RECT 37.520 77.600 37.840 77.920 ;
        RECT 41.070 77.570 41.390 77.890 ;
        RECT 42.170 77.580 42.490 77.900 ;
        RECT 43.260 77.580 43.580 77.900 ;
        RECT 19.260 75.510 19.580 77.260 ;
        RECT 19.760 76.890 20.080 77.210 ;
        RECT 20.850 76.870 21.170 77.190 ;
        RECT 21.960 76.860 22.280 77.180 ;
        RECT 19.760 75.520 20.080 75.840 ;
        RECT 20.850 75.520 21.170 75.840 ;
        RECT 21.950 75.520 22.270 75.840 ;
        RECT 19.140 74.910 19.680 75.510 ;
        RECT 19.200 74.790 19.520 74.910 ;
        RECT 20.300 74.790 20.620 75.110 ;
        RECT 21.400 74.790 21.720 75.110 ;
        RECT 19.200 73.420 19.520 73.740 ;
        RECT 20.300 73.420 20.620 73.740 ;
        RECT 21.400 73.420 21.720 73.740 ;
        RECT 18.630 72.780 18.950 73.100 ;
        RECT 19.760 72.740 20.080 73.060 ;
        RECT 20.850 72.740 21.170 73.060 ;
        RECT 21.950 72.750 22.270 73.070 ;
        RECT 18.640 72.310 18.960 72.630 ;
        RECT 22.480 72.300 22.740 77.280 ;
        RECT 22.880 76.950 23.120 77.270 ;
        RECT 24.120 76.940 24.360 77.260 ;
        RECT 23.120 76.290 23.380 76.750 ;
        RECT 23.860 76.310 24.120 76.750 ;
        RECT 23.110 75.950 23.390 76.290 ;
        RECT 23.850 75.970 24.130 76.310 ;
        RECT 23.120 74.540 23.380 75.950 ;
        RECT 23.860 74.540 24.120 75.970 ;
        RECT 11.270 69.940 11.920 71.260 ;
        RECT 23.120 71.110 24.120 74.540 ;
        RECT 24.500 72.300 24.760 77.280 ;
        RECT 24.960 76.860 25.280 77.180 ;
        RECT 26.070 76.870 26.390 77.190 ;
        RECT 27.160 76.890 27.480 77.210 ;
        RECT 24.970 75.520 25.290 75.840 ;
        RECT 26.070 75.520 26.390 75.840 ;
        RECT 27.160 75.520 27.480 75.840 ;
        RECT 27.630 75.110 27.970 77.280 ;
        RECT 29.060 75.140 29.400 77.270 ;
        RECT 29.570 76.920 29.890 77.240 ;
        RECT 30.660 76.900 30.980 77.220 ;
        RECT 31.770 76.890 32.090 77.210 ;
        RECT 29.570 75.550 29.890 75.870 ;
        RECT 30.660 75.550 30.980 75.870 ;
        RECT 31.760 75.550 32.080 75.870 ;
        RECT 25.520 74.790 25.840 75.110 ;
        RECT 26.620 74.790 26.940 75.110 ;
        RECT 27.630 74.790 28.040 75.110 ;
        RECT 29.010 74.820 29.400 75.140 ;
        RECT 30.110 74.820 30.430 75.140 ;
        RECT 31.210 74.820 31.530 75.140 ;
        RECT 27.630 74.490 27.970 74.790 ;
        RECT 27.570 73.970 28.030 74.490 ;
        RECT 29.060 73.770 29.400 74.820 ;
        RECT 25.520 73.420 25.840 73.740 ;
        RECT 26.620 73.420 26.940 73.740 ;
        RECT 27.720 73.420 28.040 73.740 ;
        RECT 29.010 73.600 29.400 73.770 ;
        RECT 28.440 73.100 28.760 73.130 ;
        RECT 24.970 72.750 25.290 73.070 ;
        RECT 26.070 72.740 26.390 73.060 ;
        RECT 27.160 72.740 27.480 73.060 ;
        RECT 28.290 72.810 28.760 73.100 ;
        RECT 28.970 73.080 29.490 73.600 ;
        RECT 30.110 73.450 30.430 73.770 ;
        RECT 31.210 73.450 31.530 73.770 ;
        RECT 28.290 72.780 28.610 72.810 ;
        RECT 29.570 72.770 29.890 73.090 ;
        RECT 30.660 72.770 30.980 73.090 ;
        RECT 31.760 72.780 32.080 73.100 ;
        RECT 28.450 72.630 28.770 72.660 ;
        RECT 28.280 72.340 28.770 72.630 ;
        RECT 28.280 72.310 28.600 72.340 ;
        RECT 32.290 72.330 32.550 77.310 ;
        RECT 32.690 76.970 32.930 77.290 ;
        RECT 33.930 76.970 34.170 77.290 ;
        RECT 32.930 76.290 33.190 76.780 ;
        RECT 32.920 75.950 33.200 76.290 ;
        RECT 32.930 74.770 33.190 75.950 ;
        RECT 33.670 74.770 33.930 76.780 ;
        RECT 32.930 71.130 33.930 74.770 ;
        RECT 34.310 72.330 34.570 77.310 ;
        RECT 34.770 76.890 35.090 77.210 ;
        RECT 35.880 76.900 36.200 77.220 ;
        RECT 36.970 76.920 37.290 77.240 ;
        RECT 34.780 75.550 35.100 75.870 ;
        RECT 35.880 75.550 36.200 75.870 ;
        RECT 36.970 75.550 37.290 75.870 ;
        RECT 37.480 75.140 37.750 77.310 ;
        RECT 40.510 76.870 40.830 77.190 ;
        RECT 41.620 76.880 41.940 77.200 ;
        RECT 42.710 76.900 43.030 77.220 ;
        RECT 44.550 76.910 44.800 84.750 ;
        RECT 45.050 77.810 45.300 85.680 ;
        RECT 45.530 78.720 45.780 87.520 ;
        RECT 46.030 79.610 46.280 88.450 ;
        RECT 61.870 81.110 62.370 97.490 ;
        RECT 62.800 86.390 63.300 97.490 ;
        RECT 63.930 91.620 64.430 117.890 ;
        RECT 65.060 105.950 65.560 118.510 ;
        RECT 73.920 116.910 75.200 129.110 ;
        RECT 73.910 115.570 75.200 116.910 ;
        RECT 67.170 111.500 67.590 111.650 ;
        RECT 68.200 111.500 68.620 111.650 ;
        RECT 71.900 111.570 72.130 111.650 ;
        RECT 67.170 111.360 68.620 111.500 ;
        RECT 72.160 109.420 72.580 115.470 ;
        RECT 73.920 115.080 75.200 115.570 ;
        RECT 74.640 112.610 74.870 115.080 ;
        RECT 74.370 112.130 74.870 112.610 ;
        RECT 74.470 109.420 74.870 112.130 ;
        RECT 75.860 114.260 76.090 115.470 ;
        RECT 80.860 114.650 81.170 115.090 ;
        RECT 75.860 113.470 76.120 114.260 ;
        RECT 78.280 113.900 78.480 113.930 ;
        RECT 75.860 111.320 76.090 113.470 ;
        RECT 78.190 113.400 78.500 113.900 ;
        RECT 81.010 113.690 81.330 114.010 ;
        RECT 78.280 111.650 78.480 113.400 ;
        RECT 81.790 113.030 81.980 130.240 ;
        RECT 100.470 128.000 104.820 131.700 ;
        RECT 130.020 127.520 133.250 132.100 ;
        RECT 129.720 123.470 133.270 127.520 ;
        RECT 158.610 121.890 161.840 132.100 ;
        RECT 85.130 121.580 85.950 121.670 ;
        RECT 85.070 120.890 85.950 121.580 ;
        RECT 82.380 114.010 82.570 115.470 ;
        RECT 82.820 114.820 83.100 115.470 ;
        RECT 82.710 114.220 83.100 114.820 ;
        RECT 82.380 113.980 82.600 114.010 ;
        RECT 82.360 113.710 82.610 113.980 ;
        RECT 82.370 113.700 82.610 113.710 ;
        RECT 82.370 113.460 82.600 113.700 ;
        RECT 81.790 112.900 82.220 113.030 ;
        RECT 81.790 112.580 82.240 112.900 ;
        RECT 81.790 112.300 81.980 112.580 ;
        RECT 81.790 111.980 82.240 112.300 ;
        RECT 81.790 111.860 82.220 111.980 ;
        RECT 78.280 111.570 78.610 111.650 ;
        RECT 78.860 111.630 79.140 111.650 ;
        RECT 78.860 111.570 79.200 111.630 ;
        RECT 75.860 110.530 76.120 111.320 ;
        RECT 75.860 109.420 76.090 110.530 ;
        RECT 78.280 109.480 78.480 111.570 ;
        RECT 78.880 111.330 79.200 111.570 ;
        RECT 80.610 111.310 80.930 111.630 ;
        RECT 81.790 111.350 81.980 111.860 ;
        RECT 82.410 111.650 82.570 113.460 ;
        RECT 82.820 112.620 83.100 114.220 ;
        RECT 82.820 112.300 83.180 112.620 ;
        RECT 82.820 111.650 83.100 112.300 ;
        RECT 82.410 111.430 83.100 111.650 ;
        RECT 83.210 111.500 83.490 111.650 ;
        RECT 81.010 110.930 81.330 111.250 ;
        RECT 81.590 111.030 81.980 111.350 ;
        RECT 82.370 111.180 83.100 111.430 ;
        RECT 80.760 110.480 81.080 110.800 ;
        RECT 81.790 110.700 81.980 111.030 ;
        RECT 82.360 110.910 83.100 111.180 ;
        RECT 81.540 110.380 81.980 110.700 ;
        RECT 79.180 109.920 79.500 110.240 ;
        RECT 79.650 109.950 79.970 110.270 ;
        RECT 80.180 109.800 80.410 110.090 ;
        RECT 80.750 109.920 81.170 110.240 ;
        RECT 80.860 109.800 81.170 109.920 ;
        RECT 81.310 109.870 81.540 110.100 ;
        RECT 81.790 109.870 81.980 110.380 ;
        RECT 81.310 109.810 81.980 109.870 ;
        RECT 70.380 108.930 70.850 109.420 ;
        RECT 64.830 105.650 65.560 105.950 ;
        RECT 65.060 96.790 65.560 105.650 ;
        RECT 65.010 96.230 65.560 96.790 ;
        RECT 63.920 91.060 64.440 91.620 ;
        RECT 62.790 85.870 63.310 86.390 ;
        RECT 61.710 80.540 62.370 81.110 ;
        RECT 45.980 79.030 46.350 79.610 ;
        RECT 45.450 78.140 45.820 78.720 ;
        RECT 44.960 77.230 45.330 77.810 ;
        RECT 40.520 75.530 40.840 75.850 ;
        RECT 41.620 75.530 41.940 75.850 ;
        RECT 42.710 75.530 43.030 75.850 ;
        RECT 35.330 74.820 35.650 75.140 ;
        RECT 36.430 74.820 36.750 75.140 ;
        RECT 37.480 74.820 37.850 75.140 ;
        RECT 43.220 75.120 43.550 76.690 ;
        RECT 44.490 76.340 44.840 76.910 ;
        RECT 37.480 73.770 37.750 74.820 ;
        RECT 41.070 74.800 41.390 75.120 ;
        RECT 42.170 74.800 42.490 75.120 ;
        RECT 43.220 74.800 43.590 75.120 ;
        RECT 35.330 73.450 35.650 73.770 ;
        RECT 36.430 73.450 36.750 73.770 ;
        RECT 37.480 73.450 37.850 73.770 ;
        RECT 43.220 73.750 43.550 74.800 ;
        RECT 43.990 74.240 44.270 74.770 ;
        RECT 43.990 73.940 44.450 74.240 ;
        RECT 43.980 73.920 44.450 73.940 ;
        RECT 34.780 72.780 35.100 73.100 ;
        RECT 35.880 72.770 36.200 73.090 ;
        RECT 36.970 72.770 37.290 73.090 ;
        RECT 37.480 72.720 37.750 73.450 ;
        RECT 41.070 73.430 41.390 73.750 ;
        RECT 42.170 73.430 42.490 73.750 ;
        RECT 43.220 73.430 43.590 73.750 ;
        RECT 43.980 73.490 44.270 73.920 ;
        RECT 38.100 72.810 38.420 73.130 ;
        RECT 40.520 72.760 40.840 73.080 ;
        RECT 41.620 72.750 41.940 73.070 ;
        RECT 42.710 72.750 43.030 73.070 ;
        RECT 37.370 72.160 37.860 72.720 ;
        RECT 38.090 72.340 38.410 72.660 ;
        RECT 34.060 71.130 34.950 71.170 ;
        RECT 22.640 71.070 24.570 71.110 ;
        RECT 22.100 69.880 24.570 71.070 ;
        RECT 9.620 65.650 9.990 66.030 ;
        RECT 8.970 65.030 9.360 65.420 ;
        RECT 8.370 64.400 8.750 64.790 ;
        RECT 7.780 63.770 8.130 64.140 ;
        RECT 7.140 63.090 7.500 63.470 ;
        RECT 6.550 62.850 6.890 62.860 ;
        RECT 6.530 62.480 6.910 62.850 ;
        RECT 6.550 62.470 6.880 62.480 ;
        RECT 4.770 60.630 5.120 60.960 ;
        RECT 4.790 60.570 5.120 60.630 ;
        RECT 3.500 59.350 3.850 59.680 ;
        RECT 3.500 59.280 3.830 59.350 ;
        RECT 1.360 58.620 2.600 58.950 ;
        RECT 2.890 58.650 3.330 59.070 ;
        RECT 1.360 58.510 1.940 58.620 ;
        RECT 22.100 58.390 23.040 69.880 ;
        RECT 32.450 69.850 34.950 71.130 ;
        RECT 34.060 59.850 34.950 69.850 ;
        RECT 43.220 66.700 43.550 73.430 ;
        RECT 43.840 72.790 44.160 73.110 ;
        RECT 43.830 72.320 44.150 72.640 ;
        RECT 61.870 72.230 62.370 80.540 ;
        RECT 62.800 73.140 63.300 85.870 ;
        RECT 63.930 74.010 64.430 91.060 ;
        RECT 65.060 75.520 65.560 96.230 ;
        RECT 70.430 105.950 70.830 108.930 ;
        RECT 71.350 108.320 71.770 108.680 ;
        RECT 70.430 105.650 70.950 105.950 ;
        RECT 67.950 83.080 68.530 83.640 ;
        RECT 67.980 83.070 68.490 83.080 ;
        RECT 65.060 74.960 65.620 75.520 ;
        RECT 65.060 74.830 65.560 74.960 ;
        RECT 67.980 71.200 68.480 83.070 ;
        RECT 67.350 69.920 68.480 71.200 ;
        RECT 69.230 70.440 69.460 72.510 ;
        RECT 69.220 70.210 69.510 70.440 ;
        RECT 69.230 68.830 69.460 70.210 ;
        RECT 69.220 68.600 69.510 68.830 ;
        RECT 69.230 67.230 69.460 68.600 ;
        RECT 69.220 67.000 69.510 67.230 ;
        RECT 43.160 66.310 43.590 66.700 ;
        RECT 69.230 65.610 69.460 67.000 ;
        RECT 70.430 66.140 70.830 105.650 ;
        RECT 70.430 66.120 70.960 66.140 ;
        RECT 71.360 66.120 71.750 108.320 ;
        RECT 72.270 105.930 72.720 106.360 ;
        RECT 72.290 66.120 72.680 105.930 ;
        RECT 73.130 105.670 73.510 105.680 ;
        RECT 73.110 105.370 73.530 105.670 ;
        RECT 70.430 65.920 72.950 66.120 ;
        RECT 69.220 65.380 69.510 65.610 ;
        RECT 70.430 65.580 70.830 65.920 ;
        RECT 69.230 64.010 69.460 65.380 ;
        RECT 70.420 65.120 70.890 65.580 ;
        RECT 71.360 64.780 71.750 65.920 ;
        RECT 69.950 64.400 70.270 64.480 ;
        RECT 71.330 64.400 71.790 64.780 ;
        RECT 69.950 64.220 72.040 64.400 ;
        RECT 71.530 64.180 72.040 64.220 ;
        RECT 71.750 64.170 72.040 64.180 ;
        RECT 69.220 63.780 69.510 64.010 ;
        RECT 72.290 63.960 72.680 65.920 ;
        RECT 69.230 62.390 69.460 63.780 ;
        RECT 72.270 63.500 72.740 63.960 ;
        RECT 72.780 62.890 72.950 65.920 ;
        RECT 73.130 63.160 73.510 105.370 ;
        RECT 74.470 82.140 74.700 109.420 ;
        RECT 77.770 109.260 78.000 109.450 ;
        RECT 77.770 109.160 78.120 109.260 ;
        RECT 78.270 109.190 78.500 109.480 ;
        RECT 80.200 109.330 80.390 109.800 ;
        RECT 80.870 109.790 81.080 109.800 ;
        RECT 80.850 109.470 81.110 109.790 ;
        RECT 77.780 108.940 78.120 109.160 ;
        RECT 77.780 108.510 78.120 108.730 ;
        RECT 77.770 108.410 78.120 108.510 ;
        RECT 78.280 108.480 78.480 109.190 ;
        RECT 80.130 109.010 80.390 109.330 ;
        RECT 80.380 108.670 80.700 108.990 ;
        RECT 77.770 108.220 78.000 108.410 ;
        RECT 78.270 108.190 78.500 108.480 ;
        RECT 80.130 108.340 80.390 108.660 ;
        RECT 78.280 106.460 78.480 108.190 ;
        RECT 80.200 107.870 80.390 108.340 ;
        RECT 80.870 108.180 81.080 109.470 ;
        RECT 81.310 109.320 81.500 109.810 ;
        RECT 81.540 109.550 81.980 109.810 ;
        RECT 81.790 109.480 81.980 109.550 ;
        RECT 81.140 109.070 81.500 109.320 ;
        RECT 81.770 109.220 82.000 109.480 ;
        RECT 82.380 109.420 83.100 110.910 ;
        RECT 83.220 110.070 83.490 111.500 ;
        RECT 83.840 111.080 84.160 111.400 ;
        RECT 83.220 109.780 83.500 110.070 ;
        RECT 81.590 109.190 82.000 109.220 ;
        RECT 81.140 109.000 81.400 109.070 ;
        RECT 81.590 108.900 81.980 109.190 ;
        RECT 81.140 108.600 81.400 108.670 ;
        RECT 81.140 108.350 81.500 108.600 ;
        RECT 81.790 108.480 81.980 108.900 ;
        RECT 81.770 108.390 82.000 108.480 ;
        RECT 80.850 107.890 81.080 108.180 ;
        RECT 79.180 107.430 79.500 107.750 ;
        RECT 80.180 107.580 80.410 107.870 ;
        RECT 81.310 107.860 81.500 108.350 ;
        RECT 81.590 108.190 82.000 108.390 ;
        RECT 81.590 108.070 81.980 108.190 ;
        RECT 80.750 107.430 81.070 107.750 ;
        RECT 81.310 107.740 81.540 107.860 ;
        RECT 81.790 107.740 81.980 108.070 ;
        RECT 81.310 107.570 81.980 107.740 ;
        RECT 81.540 107.420 81.980 107.570 ;
        RECT 79.180 106.900 79.500 107.220 ;
        RECT 80.180 106.780 80.410 107.070 ;
        RECT 80.750 106.900 81.070 107.220 ;
        RECT 81.310 106.910 81.540 107.080 ;
        RECT 81.790 106.910 81.980 107.420 ;
        RECT 81.310 106.790 81.980 106.910 ;
        RECT 77.770 106.240 78.000 106.430 ;
        RECT 77.770 106.140 78.120 106.240 ;
        RECT 78.270 106.170 78.500 106.460 ;
        RECT 80.200 106.310 80.390 106.780 ;
        RECT 77.780 105.920 78.120 106.140 ;
        RECT 77.780 105.490 78.120 105.710 ;
        RECT 77.770 105.390 78.120 105.490 ;
        RECT 78.280 105.650 78.480 106.170 ;
        RECT 80.130 105.990 80.390 106.310 ;
        RECT 81.310 106.300 81.500 106.790 ;
        RECT 81.540 106.590 81.980 106.790 ;
        RECT 81.790 106.460 81.980 106.590 ;
        RECT 81.140 106.100 81.500 106.300 ;
        RECT 81.770 106.260 82.000 106.460 ;
        RECT 81.020 106.050 81.500 106.100 ;
        RECT 81.590 106.170 82.000 106.260 ;
        RECT 81.020 105.980 81.400 106.050 ;
        RECT 81.020 105.800 81.340 105.980 ;
        RECT 81.590 105.940 81.980 106.170 ;
        RECT 81.790 105.800 81.980 105.940 ;
        RECT 82.550 105.800 82.890 109.420 ;
        RECT 81.020 105.740 82.890 105.800 ;
        RECT 81.070 105.660 82.890 105.740 ;
        RECT 78.280 105.600 78.610 105.650 ;
        RECT 78.860 105.600 79.140 105.650 ;
        RECT 78.280 105.460 78.480 105.600 ;
        RECT 77.770 105.200 78.000 105.390 ;
        RECT 78.270 105.170 78.500 105.460 ;
        RECT 80.130 105.320 80.390 105.640 ;
        RECT 81.140 105.580 81.400 105.650 ;
        RECT 81.140 105.330 81.500 105.580 ;
        RECT 81.790 105.460 81.980 105.660 ;
        RECT 82.550 105.600 82.890 105.660 ;
        RECT 83.220 107.480 83.490 109.780 ;
        RECT 83.890 108.860 84.210 109.180 ;
        RECT 83.880 108.140 84.200 108.460 ;
        RECT 83.220 107.190 83.500 107.480 ;
        RECT 83.220 105.600 83.490 107.190 ;
        RECT 83.800 105.890 84.120 106.210 ;
        RECT 78.280 104.300 78.480 105.170 ;
        RECT 80.200 104.850 80.390 105.320 ;
        RECT 79.180 104.410 79.500 104.730 ;
        RECT 80.180 104.560 80.410 104.850 ;
        RECT 81.310 104.840 81.500 105.330 ;
        RECT 81.770 105.170 82.000 105.460 ;
        RECT 80.750 104.410 81.070 104.730 ;
        RECT 81.310 104.550 81.540 104.840 ;
        RECT 81.790 104.300 81.980 105.170 ;
        RECT 85.070 101.890 85.780 120.890 ;
        RECT 158.410 119.360 162.000 121.890 ;
        RECT 187.200 118.400 190.430 132.100 ;
        RECT 212.630 129.160 213.620 129.170 ;
        RECT 212.630 128.640 214.020 129.160 ;
        RECT 207.400 128.110 210.820 128.160 ;
        RECT 207.390 127.540 210.830 128.110 ;
        RECT 205.540 126.720 206.260 127.270 ;
        RECT 205.760 126.710 206.260 126.720 ;
        RECT 186.890 114.780 190.650 118.400 ;
        RECT 201.240 117.750 204.650 118.030 ;
        RECT 201.240 117.730 205.360 117.750 ;
        RECT 201.240 117.710 206.110 117.730 ;
        RECT 207.940 117.710 212.240 126.770 ;
        RECT 213.530 125.030 214.020 128.640 ;
        RECT 201.240 115.960 214.640 117.710 ;
        RECT 201.240 115.950 215.590 115.960 ;
        RECT 201.240 115.600 215.740 115.950 ;
        RECT 201.240 115.590 215.590 115.600 ;
        RECT 84.940 101.100 85.780 101.890 ;
        RECT 109.560 84.320 113.980 114.430 ;
        RECT 201.240 113.990 214.640 115.590 ;
        RECT 204.650 113.810 214.640 113.990 ;
        RECT 204.650 113.800 214.270 113.810 ;
        RECT 204.650 113.790 206.110 113.800 ;
        RECT 205.340 113.780 206.110 113.790 ;
        RECT 207.660 104.090 212.810 113.800 ;
        RECT 207.660 103.420 212.800 104.090 ;
        RECT 213.470 104.000 214.100 104.060 ;
        RECT 213.450 103.420 214.100 104.000 ;
        RECT 213.470 102.670 214.100 103.420 ;
        RECT 205.840 101.950 214.100 102.670 ;
        RECT 211.510 101.720 214.100 101.950 ;
        RECT 213.470 101.690 214.100 101.720 ;
        RECT 212.630 100.570 213.620 100.580 ;
        RECT 212.630 100.050 214.020 100.570 ;
        RECT 207.400 99.520 210.820 99.570 ;
        RECT 207.390 98.950 210.830 99.520 ;
        RECT 205.540 98.130 206.260 98.680 ;
        RECT 205.760 98.120 206.260 98.130 ;
        RECT 192.830 89.120 195.150 89.200 ;
        RECT 204.640 89.140 205.340 89.150 ;
        RECT 204.640 89.120 206.110 89.140 ;
        RECT 207.940 89.120 212.240 98.180 ;
        RECT 213.530 96.440 214.020 100.050 ;
        RECT 192.830 87.370 214.640 89.120 ;
        RECT 192.830 87.360 215.590 87.370 ;
        RECT 192.830 87.010 215.740 87.360 ;
        RECT 192.830 87.000 215.590 87.010 ;
        RECT 192.830 85.890 214.640 87.000 ;
        RECT 192.830 85.830 195.150 85.890 ;
        RECT 204.640 85.220 214.640 85.890 ;
        RECT 204.640 85.210 214.270 85.220 ;
        RECT 204.640 85.190 206.110 85.210 ;
        RECT 80.660 83.060 81.380 83.630 ;
        RECT 74.470 81.910 74.710 82.140 ;
        RECT 74.470 76.100 74.700 81.910 ;
        RECT 80.720 76.050 81.230 83.060 ;
        RECT 109.530 83.000 114.000 84.320 ;
        RECT 80.580 76.000 81.230 76.050 ;
        RECT 80.570 75.820 81.230 76.000 ;
        RECT 80.540 75.810 81.230 75.820 ;
        RECT 80.540 75.440 81.140 75.810 ;
        RECT 80.540 73.570 81.120 75.440 ;
        RECT 80.190 72.580 81.120 73.570 ;
        RECT 80.540 71.800 81.120 72.580 ;
        RECT 80.550 71.190 81.120 71.800 ;
        RECT 80.540 70.190 81.120 71.190 ;
        RECT 74.730 69.430 75.050 69.750 ;
        RECT 80.550 69.590 81.120 70.190 ;
        RECT 74.730 68.760 75.050 69.080 ;
        RECT 74.850 67.790 75.170 67.840 ;
        RECT 74.620 67.560 75.170 67.790 ;
        RECT 74.850 67.520 75.170 67.560 ;
        RECT 74.850 66.180 75.170 66.230 ;
        RECT 74.620 65.950 75.170 66.180 ;
        RECT 74.850 65.910 75.170 65.950 ;
        RECT 74.840 64.570 75.160 64.620 ;
        RECT 74.610 64.340 75.160 64.570 ;
        RECT 74.840 64.300 75.160 64.340 ;
        RECT 72.360 62.670 72.950 62.890 ;
        RECT 73.100 62.700 73.540 63.160 ;
        RECT 74.840 62.950 75.160 63.000 ;
        RECT 74.610 62.720 75.160 62.950 ;
        RECT 74.840 62.680 75.160 62.720 ;
        RECT 72.360 62.660 72.650 62.670 ;
        RECT 69.220 62.160 69.510 62.390 ;
        RECT 69.230 60.790 69.460 62.160 ;
        RECT 80.540 62.150 81.120 69.590 ;
        RECT 80.550 61.550 81.120 62.150 ;
        RECT 74.840 61.340 75.160 61.390 ;
        RECT 74.610 61.110 75.160 61.340 ;
        RECT 74.840 61.070 75.160 61.110 ;
        RECT 69.220 60.560 69.510 60.790 ;
        RECT 80.540 60.730 81.120 61.550 ;
        RECT 80.540 60.720 81.080 60.730 ;
        RECT 34.060 59.120 34.980 59.850 ;
        RECT 69.230 59.170 69.460 60.560 ;
        RECT 74.470 59.470 74.790 59.790 ;
        RECT 74.520 59.240 74.750 59.470 ;
        RECT 34.030 58.390 34.950 59.120 ;
        RECT 69.220 58.940 69.510 59.170 ;
        RECT 74.850 58.140 75.170 58.190 ;
        RECT -151.050 57.350 -141.110 58.020 ;
        RECT -127.070 57.870 -124.840 58.020 ;
        RECT 74.620 57.910 75.170 58.140 ;
        RECT 74.850 57.870 75.170 57.910 ;
        RECT -150.680 57.340 -141.110 57.350 ;
        RECT -149.220 47.630 -144.070 57.340 ;
        RECT -142.520 57.320 -141.110 57.340 ;
        RECT -141.750 57.310 -141.110 57.320 ;
        RECT 74.840 56.550 75.160 56.600 ;
        RECT 71.640 56.470 71.960 56.520 ;
        RECT 72.580 56.470 72.900 56.520 ;
        RECT 71.410 56.240 71.960 56.470 ;
        RECT 72.350 56.240 72.900 56.470 ;
        RECT 73.530 56.410 73.850 56.460 ;
        RECT 71.640 56.200 71.960 56.240 ;
        RECT 72.580 56.200 72.900 56.240 ;
        RECT 73.300 56.180 73.850 56.410 ;
        RECT 74.610 56.320 75.160 56.550 ;
        RECT 74.840 56.280 75.160 56.320 ;
        RECT 73.530 56.140 73.850 56.180 ;
        RECT -150.510 47.540 -149.880 47.600 ;
        RECT -150.510 46.960 -149.860 47.540 ;
        RECT -149.210 46.960 -144.070 47.630 ;
        RECT -150.510 46.210 -149.880 46.960 ;
        RECT -150.510 45.490 -142.250 46.210 ;
        RECT -150.510 45.260 -147.920 45.490 ;
        RECT -150.510 45.230 -149.880 45.260 ;
        RECT -150.030 44.110 -149.040 44.120 ;
        RECT -150.430 43.590 -149.040 44.110 ;
        RECT -150.430 39.980 -149.940 43.590 ;
        RECT -147.230 43.060 -143.810 43.110 ;
        RECT -147.240 42.490 -143.800 43.060 ;
        RECT -148.650 32.660 -144.350 41.720 ;
        RECT -142.670 41.670 -141.950 42.220 ;
        RECT -142.670 41.660 -142.170 41.670 ;
        RECT -142.520 32.670 -141.750 32.680 ;
        RECT -142.520 32.660 -141.120 32.670 ;
        RECT -122.560 32.660 -120.150 32.760 ;
        RECT -151.050 30.910 -120.150 32.660 ;
        RECT -152.000 30.900 -120.150 30.910 ;
        RECT -152.150 30.550 -120.150 30.900 ;
        RECT -152.000 30.540 -120.150 30.550 ;
        RECT -151.050 29.430 -120.150 30.540 ;
        RECT -151.050 28.760 -141.120 29.430 ;
        RECT -122.560 29.330 -120.150 29.430 ;
        RECT -150.680 28.750 -141.120 28.760 ;
        RECT -149.220 19.040 -144.070 28.750 ;
        RECT -142.520 28.730 -141.120 28.750 ;
        RECT -150.510 18.950 -149.880 19.010 ;
        RECT -150.510 18.370 -149.860 18.950 ;
        RECT -149.210 18.370 -144.070 19.040 ;
        RECT -150.510 17.620 -149.880 18.370 ;
        RECT -150.510 16.900 -142.250 17.620 ;
        RECT -150.510 16.670 -147.920 16.900 ;
        RECT -150.510 16.640 -149.880 16.670 ;
        RECT -150.030 15.520 -149.040 15.530 ;
        RECT -150.430 15.000 -149.040 15.520 ;
        RECT -150.430 11.390 -149.940 15.000 ;
        RECT -147.230 14.470 -143.810 14.520 ;
        RECT -147.240 13.900 -143.800 14.470 ;
        RECT -148.650 4.070 -144.350 13.130 ;
        RECT -142.670 13.080 -141.950 13.630 ;
        RECT -142.670 13.070 -142.170 13.080 ;
        RECT -142.520 4.070 -141.110 4.090 ;
        RECT -118.000 4.070 -115.730 4.140 ;
        RECT -151.050 2.320 -115.730 4.070 ;
        RECT -152.000 2.310 -115.730 2.320 ;
        RECT -152.150 1.960 -115.730 2.310 ;
        RECT -152.000 1.950 -115.730 1.960 ;
        RECT -151.050 0.840 -115.730 1.950 ;
        RECT -151.050 0.170 -141.110 0.840 ;
        RECT -118.000 0.740 -115.730 0.840 ;
        RECT -150.680 0.160 -141.110 0.170 ;
        RECT -149.220 -9.550 -144.070 0.160 ;
        RECT -142.520 0.150 -141.110 0.160 ;
        RECT -142.520 0.140 -141.750 0.150 ;
        RECT -150.510 -9.640 -149.880 -9.580 ;
        RECT -150.510 -10.220 -149.860 -9.640 ;
        RECT -149.210 -10.220 -144.070 -9.550 ;
        RECT -150.510 -10.970 -149.880 -10.220 ;
        RECT -150.510 -11.690 -142.250 -10.970 ;
        RECT -150.510 -11.920 -147.920 -11.690 ;
        RECT -150.510 -11.950 -149.880 -11.920 ;
        RECT -150.030 -13.070 -149.040 -13.060 ;
        RECT -150.430 -13.590 -149.040 -13.070 ;
        RECT -150.430 -17.200 -149.940 -13.590 ;
        RECT -147.230 -14.120 -143.810 -14.070 ;
        RECT -147.240 -14.690 -143.800 -14.120 ;
        RECT -148.650 -24.520 -144.350 -15.460 ;
        RECT -142.670 -15.510 -141.950 -14.960 ;
        RECT -142.670 -15.520 -142.170 -15.510 ;
        RECT -142.520 -24.520 -141.120 -24.500 ;
        RECT -113.640 -24.520 -111.390 -24.460 ;
        RECT -151.050 -26.270 -111.390 -24.520 ;
        RECT -152.000 -26.280 -111.390 -26.270 ;
        RECT -152.150 -26.630 -111.390 -26.280 ;
        RECT -152.000 -26.640 -111.390 -26.630 ;
        RECT -151.050 -27.750 -111.390 -26.640 ;
        RECT -151.050 -28.420 -141.120 -27.750 ;
        RECT -113.640 -27.830 -111.390 -27.750 ;
        RECT -150.680 -28.430 -141.120 -28.420 ;
        RECT -149.220 -38.140 -144.070 -28.430 ;
        RECT -142.520 -28.440 -141.120 -28.430 ;
        RECT -142.520 -28.450 -141.750 -28.440 ;
        RECT -150.510 -38.230 -149.880 -38.170 ;
        RECT -150.510 -38.810 -149.860 -38.230 ;
        RECT -149.210 -38.810 -144.070 -38.140 ;
        RECT -150.510 -39.560 -149.880 -38.810 ;
        RECT -150.510 -40.280 -142.250 -39.560 ;
        RECT -150.510 -40.510 -147.920 -40.280 ;
        RECT -150.510 -40.540 -149.880 -40.510 ;
        RECT -150.030 -41.660 -149.040 -41.650 ;
        RECT -150.430 -42.180 -149.040 -41.660 ;
        RECT -150.430 -45.790 -149.940 -42.180 ;
        RECT -147.230 -42.710 -143.810 -42.660 ;
        RECT -147.240 -43.280 -143.800 -42.710 ;
        RECT -148.650 -53.110 -144.350 -44.050 ;
        RECT -142.670 -44.100 -141.950 -43.550 ;
        RECT -142.670 -44.110 -142.170 -44.100 ;
        RECT -142.520 -53.110 -141.120 -53.090 ;
        RECT -109.320 -53.110 -107.070 -53.000 ;
        RECT -151.050 -54.860 -106.920 -53.110 ;
        RECT -152.000 -54.870 -106.920 -54.860 ;
        RECT -152.150 -55.220 -106.920 -54.870 ;
        RECT -152.000 -55.230 -106.920 -55.220 ;
        RECT -151.050 -56.340 -106.920 -55.230 ;
        RECT -151.050 -57.010 -141.120 -56.340 ;
        RECT -109.320 -56.450 -107.070 -56.340 ;
        RECT -150.680 -57.020 -141.120 -57.010 ;
        RECT -149.220 -66.730 -144.070 -57.020 ;
        RECT -142.520 -57.030 -141.120 -57.020 ;
        RECT -142.520 -57.040 -141.750 -57.030 ;
        RECT -150.510 -66.820 -149.880 -66.760 ;
        RECT -150.510 -67.400 -149.860 -66.820 ;
        RECT -149.210 -67.400 -144.070 -66.730 ;
        RECT -150.510 -68.150 -149.880 -67.400 ;
        RECT -150.510 -68.870 -142.250 -68.150 ;
        RECT -150.510 -69.100 -147.920 -68.870 ;
        RECT -150.510 -69.130 -149.880 -69.100 ;
        RECT -150.030 -70.250 -149.040 -70.240 ;
        RECT -150.430 -70.770 -149.040 -70.250 ;
        RECT -150.430 -74.380 -149.940 -70.770 ;
        RECT -147.230 -71.300 -143.810 -71.250 ;
        RECT -147.240 -71.870 -143.800 -71.300 ;
        RECT -148.650 -81.700 -144.350 -72.640 ;
        RECT -142.670 -72.690 -141.950 -72.140 ;
        RECT -142.670 -72.700 -142.170 -72.690 ;
        RECT 109.560 -78.300 113.980 83.000 ;
        RECT 207.660 75.500 212.810 85.210 ;
        RECT 207.660 74.830 212.800 75.500 ;
        RECT 213.470 75.410 214.100 75.470 ;
        RECT 213.450 74.830 214.100 75.410 ;
        RECT 213.470 74.080 214.100 74.830 ;
        RECT 205.840 73.360 214.100 74.080 ;
        RECT 211.510 73.130 214.100 73.360 ;
        RECT 213.470 73.100 214.100 73.130 ;
        RECT 212.630 71.980 213.620 71.990 ;
        RECT 212.630 71.460 214.020 71.980 ;
        RECT 207.400 70.930 210.820 70.980 ;
        RECT 207.390 70.360 210.830 70.930 ;
        RECT 205.540 69.540 206.260 70.090 ;
        RECT 205.760 69.530 206.260 69.540 ;
        RECT 188.660 60.530 191.020 60.660 ;
        RECT 204.660 60.550 205.360 60.560 ;
        RECT 204.660 60.530 206.110 60.550 ;
        RECT 207.940 60.530 212.240 69.590 ;
        RECT 213.530 67.850 214.020 71.460 ;
        RECT 188.660 58.780 214.640 60.530 ;
        RECT 188.660 58.770 215.590 58.780 ;
        RECT 188.660 58.420 215.740 58.770 ;
        RECT 188.660 58.410 215.590 58.420 ;
        RECT 188.660 57.300 214.640 58.410 ;
        RECT 188.660 57.200 191.020 57.300 ;
        RECT 204.660 56.630 214.640 57.300 ;
        RECT 204.660 56.620 214.270 56.630 ;
        RECT 204.660 56.600 206.110 56.620 ;
        RECT 207.660 46.910 212.810 56.620 ;
        RECT 207.660 46.240 212.800 46.910 ;
        RECT 213.470 46.820 214.100 46.880 ;
        RECT 213.450 46.240 214.100 46.820 ;
        RECT 213.470 45.490 214.100 46.240 ;
        RECT 205.840 44.770 214.100 45.490 ;
        RECT 211.510 44.540 214.100 44.770 ;
        RECT 213.470 44.510 214.100 44.540 ;
        RECT 212.630 43.390 213.620 43.400 ;
        RECT 212.630 42.870 214.020 43.390 ;
        RECT 207.400 42.340 210.820 42.390 ;
        RECT 207.390 41.770 210.830 42.340 ;
        RECT 205.540 40.950 206.260 41.500 ;
        RECT 205.760 40.940 206.260 40.950 ;
        RECT 184.650 31.940 186.930 32.100 ;
        RECT 204.640 31.960 205.340 31.970 ;
        RECT 204.640 31.940 206.110 31.960 ;
        RECT 207.940 31.940 212.240 41.000 ;
        RECT 213.530 39.260 214.020 42.870 ;
        RECT 184.650 30.190 214.640 31.940 ;
        RECT 184.650 30.180 215.590 30.190 ;
        RECT 184.650 29.830 215.740 30.180 ;
        RECT 184.650 29.820 215.590 29.830 ;
        RECT 184.650 28.710 214.640 29.820 ;
        RECT 184.650 28.600 186.930 28.710 ;
        RECT 204.640 28.040 214.640 28.710 ;
        RECT 204.640 28.030 214.270 28.040 ;
        RECT 204.640 28.010 206.110 28.030 ;
        RECT 207.660 18.320 212.810 28.030 ;
        RECT 207.660 17.650 212.800 18.320 ;
        RECT 213.470 18.230 214.100 18.290 ;
        RECT 213.450 17.650 214.100 18.230 ;
        RECT 213.470 16.900 214.100 17.650 ;
        RECT 205.840 16.180 214.100 16.900 ;
        RECT 211.510 15.950 214.100 16.180 ;
        RECT 213.470 15.920 214.100 15.950 ;
        RECT 212.630 14.800 213.620 14.810 ;
        RECT 212.630 14.280 214.020 14.800 ;
        RECT 207.400 13.750 210.820 13.800 ;
        RECT 207.390 13.180 210.830 13.750 ;
        RECT 205.540 12.360 206.260 12.910 ;
        RECT 205.760 12.350 206.260 12.360 ;
        RECT 180.350 3.350 182.770 3.470 ;
        RECT 204.640 3.350 206.110 3.370 ;
        RECT 207.940 3.350 212.240 12.410 ;
        RECT 213.530 10.670 214.020 14.280 ;
        RECT 180.350 1.600 214.640 3.350 ;
        RECT 180.350 1.590 215.590 1.600 ;
        RECT 180.350 1.240 215.740 1.590 ;
        RECT 180.350 1.230 215.590 1.240 ;
        RECT 180.350 0.120 214.640 1.230 ;
        RECT 180.350 -0.040 182.770 0.120 ;
        RECT 204.640 -0.550 214.640 0.120 ;
        RECT 204.640 -0.560 214.270 -0.550 ;
        RECT 204.640 -0.580 206.110 -0.560 ;
        RECT 204.640 -0.590 205.340 -0.580 ;
        RECT 207.660 -10.270 212.810 -0.560 ;
        RECT 207.660 -10.940 212.800 -10.270 ;
        RECT 213.470 -10.360 214.100 -10.300 ;
        RECT 213.450 -10.940 214.100 -10.360 ;
        RECT 213.470 -11.690 214.100 -10.940 ;
        RECT 205.840 -12.410 214.100 -11.690 ;
        RECT 211.510 -12.640 214.100 -12.410 ;
        RECT 213.470 -12.670 214.100 -12.640 ;
        RECT 212.630 -13.790 213.620 -13.780 ;
        RECT 212.630 -14.310 214.020 -13.790 ;
        RECT 207.400 -14.840 210.820 -14.790 ;
        RECT 207.390 -15.410 210.830 -14.840 ;
        RECT 205.540 -16.230 206.260 -15.680 ;
        RECT 205.760 -16.240 206.260 -16.230 ;
        RECT 176.460 -25.240 178.730 -25.130 ;
        RECT 204.650 -25.220 205.350 -25.210 ;
        RECT 204.650 -25.240 206.110 -25.220 ;
        RECT 207.940 -25.240 212.240 -16.180 ;
        RECT 213.530 -17.920 214.020 -14.310 ;
        RECT 176.460 -26.990 214.640 -25.240 ;
        RECT 176.460 -27.000 215.590 -26.990 ;
        RECT 176.460 -27.350 215.740 -27.000 ;
        RECT 176.460 -27.360 215.590 -27.350 ;
        RECT 176.460 -28.470 214.640 -27.360 ;
        RECT 176.460 -28.600 178.730 -28.470 ;
        RECT 204.650 -29.140 214.640 -28.470 ;
        RECT 204.650 -29.150 214.270 -29.140 ;
        RECT 204.650 -29.170 206.110 -29.150 ;
        RECT 207.660 -38.860 212.810 -29.150 ;
        RECT 207.660 -39.530 212.800 -38.860 ;
        RECT 213.470 -38.950 214.100 -38.890 ;
        RECT 213.450 -39.530 214.100 -38.950 ;
        RECT 213.470 -40.280 214.100 -39.530 ;
        RECT 205.840 -41.000 214.100 -40.280 ;
        RECT 211.510 -41.230 214.100 -41.000 ;
        RECT 213.470 -41.260 214.100 -41.230 ;
        RECT 212.630 -42.380 213.620 -42.370 ;
        RECT 212.630 -42.900 214.020 -42.380 ;
        RECT 207.400 -43.430 210.820 -43.380 ;
        RECT 207.390 -44.000 210.830 -43.430 ;
        RECT 205.540 -44.820 206.260 -44.270 ;
        RECT 205.760 -44.830 206.260 -44.820 ;
        RECT 172.060 -53.830 174.360 -53.750 ;
        RECT 204.650 -53.830 206.110 -53.810 ;
        RECT 207.940 -53.830 212.240 -44.770 ;
        RECT 213.530 -46.510 214.020 -42.900 ;
        RECT 172.060 -55.580 214.640 -53.830 ;
        RECT 172.060 -55.590 215.590 -55.580 ;
        RECT 172.060 -55.940 215.740 -55.590 ;
        RECT 172.060 -55.950 215.590 -55.940 ;
        RECT 172.060 -57.060 214.640 -55.950 ;
        RECT 172.060 -57.160 174.360 -57.060 ;
        RECT 204.650 -57.730 214.640 -57.060 ;
        RECT 204.650 -57.740 214.270 -57.730 ;
        RECT 204.650 -57.760 206.110 -57.740 ;
        RECT 204.650 -57.770 205.350 -57.760 ;
        RECT 207.660 -67.450 212.810 -57.740 ;
        RECT 207.660 -68.120 212.800 -67.450 ;
        RECT 213.470 -67.540 214.100 -67.480 ;
        RECT 213.450 -68.120 214.100 -67.540 ;
        RECT 213.470 -68.870 214.100 -68.120 ;
        RECT 205.840 -69.590 214.100 -68.870 ;
        RECT 211.510 -69.820 214.100 -69.590 ;
        RECT 213.470 -69.850 214.100 -69.820 ;
        RECT -142.520 -81.690 -141.750 -81.680 ;
        RECT -142.520 -81.700 -141.120 -81.690 ;
        RECT -105.260 -81.700 -102.850 -81.600 ;
        RECT -151.050 -83.450 -102.850 -81.700 ;
        RECT 108.640 -82.040 113.980 -78.300 ;
        RECT 108.640 -83.000 113.400 -82.040 ;
        RECT -152.000 -83.460 -102.850 -83.450 ;
        RECT -152.150 -83.810 -102.850 -83.460 ;
        RECT -152.000 -83.820 -102.850 -83.810 ;
        RECT -151.050 -84.930 -102.850 -83.820 ;
        RECT -151.050 -85.600 -141.120 -84.930 ;
        RECT -105.260 -85.110 -102.850 -84.930 ;
        RECT -150.680 -85.610 -141.120 -85.600 ;
        RECT -149.220 -95.320 -144.070 -85.610 ;
        RECT -142.520 -85.630 -141.120 -85.610 ;
        RECT -150.510 -95.410 -149.880 -95.350 ;
        RECT -150.510 -95.990 -149.860 -95.410 ;
        RECT -149.210 -95.990 -144.070 -95.320 ;
        RECT -150.510 -96.740 -149.880 -95.990 ;
        RECT -150.510 -97.460 -142.250 -96.740 ;
        RECT -150.510 -97.690 -147.920 -97.460 ;
        RECT -150.510 -97.720 -149.880 -97.690 ;
        RECT -150.030 -98.840 -149.040 -98.830 ;
        RECT -150.430 -99.360 -149.040 -98.840 ;
        RECT -150.430 -102.970 -149.940 -99.360 ;
        RECT -147.230 -99.890 -143.810 -99.840 ;
        RECT -147.240 -100.460 -143.800 -99.890 ;
        RECT -148.650 -110.290 -144.350 -101.230 ;
        RECT -142.670 -101.280 -141.950 -100.730 ;
        RECT -142.670 -101.290 -142.170 -101.280 ;
        RECT -142.520 -110.280 -141.750 -110.270 ;
        RECT -142.520 -110.290 -141.120 -110.280 ;
        RECT -100.980 -110.290 -98.520 -110.220 ;
        RECT -151.050 -112.040 -98.520 -110.290 ;
        RECT -152.000 -112.050 -98.520 -112.040 ;
        RECT -152.150 -112.400 -98.520 -112.050 ;
        RECT -152.000 -112.410 -98.520 -112.400 ;
        RECT -151.050 -113.520 -98.520 -112.410 ;
        RECT -151.050 -114.190 -141.120 -113.520 ;
        RECT -100.980 -113.570 -98.520 -113.520 ;
        RECT -150.680 -114.200 -141.120 -114.190 ;
        RECT -149.220 -123.910 -144.070 -114.200 ;
        RECT -142.520 -114.220 -141.120 -114.200 ;
        RECT -150.510 -124.000 -149.880 -123.940 ;
        RECT -150.510 -124.580 -149.860 -124.000 ;
        RECT -149.210 -124.580 -144.070 -123.910 ;
        RECT -150.510 -125.330 -149.880 -124.580 ;
        RECT -150.510 -126.050 -142.250 -125.330 ;
        RECT -150.510 -126.280 -147.920 -126.050 ;
        RECT -150.510 -126.310 -149.880 -126.280 ;
        RECT -150.030 -127.430 -149.040 -127.420 ;
        RECT -150.430 -127.950 -149.040 -127.430 ;
        RECT -150.430 -131.560 -149.940 -127.950 ;
        RECT -147.230 -128.480 -143.810 -128.430 ;
        RECT -147.240 -129.050 -143.800 -128.480 ;
        RECT -148.650 -138.880 -144.350 -129.820 ;
        RECT -142.670 -129.870 -141.950 -129.320 ;
        RECT -142.670 -129.880 -142.170 -129.870 ;
        RECT -141.770 -138.860 -141.130 -138.850 ;
        RECT -142.520 -138.880 -141.130 -138.860 ;
        RECT -96.610 -138.880 -94.210 -138.740 ;
        RECT -151.050 -140.630 -94.210 -138.880 ;
        RECT -152.000 -140.640 -94.210 -140.630 ;
        RECT -152.150 -140.990 -94.210 -140.640 ;
        RECT -152.000 -141.000 -94.210 -140.990 ;
        RECT -151.050 -142.110 -94.210 -141.000 ;
        RECT -151.050 -142.780 -141.130 -142.110 ;
        RECT -96.610 -142.210 -94.210 -142.110 ;
        RECT -150.680 -142.790 -141.130 -142.780 ;
        RECT -149.220 -152.500 -144.070 -142.790 ;
        RECT -142.520 -142.810 -141.750 -142.790 ;
        RECT -150.510 -152.590 -149.880 -152.530 ;
        RECT -150.510 -153.170 -149.860 -152.590 ;
        RECT -149.210 -153.170 -144.070 -152.500 ;
        RECT -150.510 -153.920 -149.880 -153.170 ;
        RECT -150.510 -154.640 -142.250 -153.920 ;
        RECT -150.510 -154.870 -147.920 -154.640 ;
        RECT -150.510 -154.900 -149.880 -154.870 ;
        RECT -150.030 -156.020 -149.040 -156.010 ;
        RECT -150.430 -156.540 -149.040 -156.020 ;
        RECT -150.430 -160.150 -149.940 -156.540 ;
        RECT -147.230 -157.070 -143.810 -157.020 ;
        RECT -147.240 -157.640 -143.800 -157.070 ;
        RECT -148.650 -167.470 -144.350 -158.410 ;
        RECT -142.670 -158.460 -141.950 -157.910 ;
        RECT -142.670 -158.470 -142.170 -158.460 ;
        RECT -142.520 -167.470 -141.130 -167.450 ;
        RECT -92.670 -167.470 -90.180 -167.390 ;
        RECT -151.050 -169.220 -90.180 -167.470 ;
        RECT -152.000 -169.230 -90.180 -169.220 ;
        RECT -152.150 -169.580 -90.180 -169.230 ;
        RECT -152.000 -169.590 -90.180 -169.580 ;
        RECT -151.050 -170.700 -90.180 -169.590 ;
        RECT -151.050 -171.370 -141.130 -170.700 ;
        RECT -92.670 -170.890 -90.180 -170.700 ;
        RECT -150.680 -171.380 -141.130 -171.370 ;
        RECT -149.220 -181.090 -144.070 -171.380 ;
        RECT -142.520 -171.390 -141.130 -171.380 ;
        RECT -142.520 -171.400 -141.750 -171.390 ;
        RECT -150.510 -181.180 -149.880 -181.120 ;
        RECT -150.510 -181.760 -149.860 -181.180 ;
        RECT -149.210 -181.760 -144.070 -181.090 ;
        RECT -150.510 -182.510 -149.880 -181.760 ;
        RECT -150.510 -183.230 -142.250 -182.510 ;
        RECT -150.510 -183.460 -147.920 -183.230 ;
        RECT -150.510 -183.490 -149.880 -183.460 ;
        RECT -150.030 -184.610 -149.040 -184.600 ;
        RECT -150.430 -185.130 -149.040 -184.610 ;
        RECT -150.430 -188.740 -149.940 -185.130 ;
        RECT -147.230 -185.660 -143.810 -185.610 ;
        RECT -147.240 -186.230 -143.800 -185.660 ;
        RECT -148.650 -196.060 -144.350 -187.000 ;
        RECT -142.670 -187.050 -141.950 -186.500 ;
        RECT -142.670 -187.060 -142.170 -187.050 ;
        RECT -142.520 -196.050 -141.750 -196.040 ;
        RECT -142.520 -196.060 -141.110 -196.050 ;
        RECT -88.200 -196.060 -85.850 -195.960 ;
        RECT -151.050 -197.810 -85.850 -196.060 ;
        RECT -152.000 -197.820 -85.850 -197.810 ;
        RECT -152.150 -198.170 -85.850 -197.820 ;
        RECT -152.000 -198.180 -85.850 -198.170 ;
        RECT -151.050 -199.290 -85.850 -198.180 ;
        RECT -151.050 -199.960 -141.110 -199.290 ;
        RECT -88.200 -199.420 -85.850 -199.290 ;
        RECT -150.680 -199.970 -141.110 -199.960 ;
        RECT -149.220 -209.680 -144.070 -199.970 ;
        RECT -142.520 -199.990 -141.110 -199.970 ;
        RECT -150.510 -209.770 -149.880 -209.710 ;
        RECT -150.510 -210.350 -149.860 -209.770 ;
        RECT -149.210 -210.350 -144.070 -209.680 ;
        RECT -150.510 -211.100 -149.880 -210.350 ;
        RECT -150.510 -211.820 -142.250 -211.100 ;
        RECT -150.510 -212.050 -147.920 -211.820 ;
        RECT -150.510 -212.080 -149.880 -212.050 ;
        RECT -150.030 -213.200 -149.040 -213.190 ;
        RECT -150.430 -213.720 -149.040 -213.200 ;
        RECT -150.430 -217.330 -149.940 -213.720 ;
        RECT -147.230 -214.250 -143.810 -214.200 ;
        RECT -147.240 -214.820 -143.800 -214.250 ;
        RECT -148.650 -224.650 -144.350 -215.590 ;
        RECT -142.670 -215.640 -141.950 -215.090 ;
        RECT -142.670 -215.650 -142.170 -215.640 ;
        RECT -141.750 -224.630 -141.110 -224.620 ;
        RECT -142.520 -224.650 -141.110 -224.630 ;
        RECT -84.200 -224.650 -81.490 -224.590 ;
        RECT -151.050 -226.400 -81.490 -224.650 ;
        RECT -152.000 -226.410 -81.490 -226.400 ;
        RECT -152.150 -226.760 -81.490 -226.410 ;
        RECT -152.000 -226.770 -81.490 -226.760 ;
        RECT -151.050 -227.880 -81.490 -226.770 ;
        RECT -151.050 -228.550 -141.110 -227.880 ;
        RECT -84.200 -228.000 -81.490 -227.880 ;
        RECT -150.680 -228.560 -141.110 -228.550 ;
        RECT -149.220 -238.270 -144.070 -228.560 ;
        RECT -142.520 -228.580 -141.750 -228.560 ;
        RECT -150.510 -238.360 -149.880 -238.300 ;
        RECT -150.510 -238.940 -149.860 -238.360 ;
        RECT -149.210 -238.940 -144.070 -238.270 ;
        RECT -150.510 -239.690 -149.880 -238.940 ;
        RECT -150.510 -240.410 -142.250 -239.690 ;
        RECT -150.510 -240.640 -147.920 -240.410 ;
        RECT -150.510 -240.670 -149.880 -240.640 ;
      LAYER via ;
        RECT -138.110 141.150 -136.080 141.480 ;
        RECT -138.170 140.290 -137.470 140.910 ;
        RECT -114.720 141.150 -111.730 141.500 ;
        RECT -109.520 141.150 -107.490 141.480 ;
        RECT -111.290 140.350 -110.940 141.110 ;
        RECT -109.580 140.290 -108.880 140.910 ;
        RECT -86.130 141.150 -83.140 141.500 ;
        RECT -80.930 141.150 -78.900 141.480 ;
        RECT -112.320 135.060 -111.900 138.230 ;
        RECT -113.290 133.240 -112.770 133.760 ;
        RECT -82.700 140.350 -82.350 141.110 ;
        RECT -80.990 140.290 -80.290 140.910 ;
        RECT -24.730 141.850 -0.930 142.110 ;
        RECT -57.540 141.150 -54.550 141.500 ;
        RECT -83.730 135.060 -83.310 138.230 ;
        RECT -84.700 133.240 -84.180 133.760 ;
        RECT -54.110 140.350 -53.760 141.110 ;
        RECT -55.140 135.060 -54.720 138.230 ;
        RECT -56.110 133.240 -55.590 133.760 ;
        RECT 7.950 141.850 28.810 142.110 ;
        RECT 3.090 141.150 5.120 141.480 ;
        RECT 3.030 140.290 3.730 140.910 ;
        RECT 26.480 141.150 29.470 141.500 ;
        RECT 31.680 141.150 33.710 141.480 ;
        RECT 29.910 140.350 30.260 141.110 ;
        RECT 31.620 140.290 32.320 140.910 ;
        RECT 55.070 141.150 58.060 141.500 ;
        RECT 60.270 141.150 62.300 141.480 ;
        RECT 28.880 135.060 29.300 138.230 ;
        RECT -149.990 129.450 -149.230 129.800 ;
        RECT -150.380 126.020 -150.030 129.010 ;
        RECT -147.110 128.420 -143.940 128.840 ;
        RECT -142.640 127.450 -142.120 127.970 ;
        RECT -68.360 127.360 -65.130 129.610 ;
        RECT -56.170 126.080 -55.650 126.450 ;
        RECT -96.950 122.870 -93.720 125.120 ;
        RECT -127.370 118.600 -125.120 121.830 ;
        RECT -138.900 115.200 -137.040 118.430 ;
        RECT 27.910 133.240 28.430 133.760 ;
        RECT -25.690 128.390 -25.300 128.780 ;
        RECT 58.500 140.350 58.850 141.110 ;
        RECT 60.210 140.290 60.910 140.910 ;
        RECT 83.660 141.150 86.650 141.500 ;
        RECT 88.860 141.150 90.890 141.480 ;
        RECT 57.470 135.060 57.890 138.230 ;
        RECT 56.500 133.240 57.020 133.760 ;
        RECT 87.090 140.350 87.440 141.110 ;
        RECT 88.800 140.290 89.500 140.910 ;
        RECT 112.250 141.150 115.240 141.500 ;
        RECT 117.450 141.150 119.480 141.480 ;
        RECT 86.060 135.060 86.480 138.230 ;
        RECT -52.830 121.700 -52.420 122.110 ;
        RECT -56.310 117.760 -55.790 118.280 ;
        RECT -150.360 102.630 -150.030 104.660 ;
        RECT -149.790 102.570 -149.170 103.270 ;
        RECT -149.990 100.860 -149.230 101.210 ;
        RECT -150.380 97.430 -150.030 100.420 ;
        RECT -147.110 99.830 -143.940 100.250 ;
        RECT -142.640 98.860 -142.120 99.380 ;
        RECT -130.850 86.610 -128.770 89.840 ;
        RECT -23.270 127.470 -23.010 127.730 ;
        RECT -20.410 127.520 -20.150 127.780 ;
        RECT -23.280 126.440 -23.020 126.700 ;
        RECT -22.560 126.410 -22.300 126.670 ;
        RECT -21.870 126.450 -21.610 126.710 ;
        RECT -23.280 125.990 -23.020 126.250 ;
        RECT -21.870 126.010 -21.610 126.270 ;
        RECT -23.280 125.570 -23.020 125.830 ;
        RECT -22.560 125.570 -22.300 125.830 ;
        RECT -21.850 125.590 -21.590 125.850 ;
        RECT -25.610 124.940 -25.220 125.330 ;
        RECT -52.780 116.910 -52.370 117.320 ;
        RECT -56.210 81.740 -55.690 82.260 ;
        RECT -52.780 80.800 -52.370 81.240 ;
        RECT -150.360 74.040 -150.030 76.070 ;
        RECT -149.790 73.980 -149.170 74.680 ;
        RECT -149.990 72.270 -149.230 72.620 ;
        RECT -150.380 68.840 -150.030 71.830 ;
        RECT -147.110 71.240 -143.940 71.660 ;
        RECT -142.640 70.270 -142.120 70.790 ;
        RECT -23.280 124.220 -23.020 124.480 ;
        RECT -24.230 123.770 -23.970 124.030 ;
        RECT -20.720 125.980 -20.460 126.240 ;
        RECT -7.170 125.670 -6.910 125.930 ;
        RECT -5.810 125.750 -5.550 126.010 ;
        RECT -5.120 125.740 -4.860 126.000 ;
        RECT -21.140 123.970 -20.880 124.230 ;
        RECT -22.580 122.770 -22.320 123.030 ;
        RECT -21.150 122.790 -20.890 123.050 ;
        RECT -23.370 122.190 -23.110 122.450 ;
        RECT -22.440 122.190 -22.180 122.450 ;
        RECT -21.740 122.190 -21.480 122.450 ;
        RECT -21.000 122.190 -20.740 122.450 ;
        RECT -20.290 122.180 -20.030 122.440 ;
        RECT -24.310 121.070 -23.890 121.490 ;
        RECT -7.890 122.010 -7.630 122.270 ;
        RECT -18.360 119.670 -18.070 120.250 ;
        RECT -5.070 118.610 -4.810 118.870 ;
        RECT -9.980 112.770 -9.720 113.030 ;
        RECT -8.890 112.780 -8.630 113.040 ;
        RECT -11.150 112.360 -10.890 112.620 ;
        RECT -10.450 112.360 -10.190 112.620 ;
        RECT -9.980 111.850 -9.720 112.110 ;
        RECT -8.890 111.860 -8.630 112.120 ;
        RECT -11.180 111.440 -10.920 111.700 ;
        RECT -10.450 111.440 -10.190 111.700 ;
        RECT -9.980 110.930 -9.720 111.190 ;
        RECT -8.890 110.940 -8.630 111.200 ;
        RECT -11.170 110.520 -10.910 110.780 ;
        RECT -10.450 110.520 -10.190 110.780 ;
        RECT -11.820 109.500 -11.560 109.760 ;
        RECT -11.860 108.540 -11.600 108.800 ;
        RECT -11.820 107.580 -11.560 107.840 ;
        RECT -10.170 109.950 -9.910 110.210 ;
        RECT -8.870 109.850 -8.610 110.110 ;
        RECT -10.170 109.490 -9.910 109.750 ;
        RECT -10.170 108.990 -9.910 109.250 ;
        RECT -8.870 108.890 -8.610 109.150 ;
        RECT -10.170 108.530 -9.910 108.790 ;
        RECT -10.170 108.030 -9.910 108.290 ;
        RECT -8.870 107.930 -8.610 108.190 ;
        RECT -10.170 107.570 -9.910 107.830 ;
        RECT 1.970 122.030 2.230 122.290 ;
        RECT 0.720 118.180 1.030 118.490 ;
        RECT 17.300 125.820 17.720 126.240 ;
        RECT 13.450 125.060 13.870 125.480 ;
        RECT 18.970 123.450 19.410 123.890 ;
        RECT 24.690 123.450 25.130 123.890 ;
        RECT 26.510 123.420 26.950 123.860 ;
        RECT 14.550 122.430 14.990 122.870 ;
        RECT 11.790 119.410 12.050 119.670 ;
        RECT 4.720 118.720 4.980 118.980 ;
        RECT 3.550 117.730 3.820 117.990 ;
        RECT -7.780 116.950 -7.430 117.300 ;
        RECT -2.530 117.260 -2.270 117.520 ;
        RECT 20.260 122.430 20.700 122.870 ;
        RECT 13.030 116.100 13.290 116.360 ;
        RECT 10.930 115.260 11.190 115.520 ;
        RECT -6.760 114.710 -6.500 115.100 ;
        RECT 9.640 114.720 9.970 114.980 ;
        RECT -7.400 113.890 -7.140 114.290 ;
        RECT -11.860 92.300 -11.600 92.770 ;
        RECT -11.220 92.300 -10.960 92.770 ;
        RECT -13.220 91.270 -12.960 91.530 ;
        RECT -13.740 90.870 -13.480 91.130 ;
        RECT -23.020 89.620 -22.360 90.280 ;
        RECT -11.140 91.250 -10.880 91.510 ;
        RECT -9.380 91.260 -9.110 91.530 ;
        RECT -11.800 90.890 -11.540 91.150 ;
        RECT -11.050 90.290 -10.790 90.550 ;
        RECT -10.400 90.290 -10.140 90.550 ;
        RECT -12.270 89.850 -12.010 90.110 ;
        RECT -11.570 89.850 -11.310 90.110 ;
        RECT -9.890 89.120 -9.630 89.380 ;
        RECT -12.720 88.500 -12.460 88.760 ;
        RECT -13.720 86.960 -13.460 87.220 ;
        RECT -17.810 85.100 -17.440 85.470 ;
        RECT -22.980 83.760 -22.320 84.420 ;
        RECT -13.720 83.870 -13.460 84.130 ;
        RECT -9.970 87.990 -9.710 88.250 ;
        RECT -8.880 90.870 -8.620 91.130 ;
        RECT -9.960 87.450 -9.700 87.710 ;
        RECT -12.720 86.950 -12.460 87.210 ;
        RECT -9.910 86.500 -9.650 86.760 ;
        RECT -12.240 85.970 -11.980 86.230 ;
        RECT -11.550 85.960 -11.290 86.220 ;
        RECT -11.070 85.190 -10.810 85.450 ;
        RECT -10.360 85.130 -10.100 85.390 ;
        RECT -10.410 84.310 -10.150 84.570 ;
        RECT -12.620 83.880 -12.360 84.140 ;
        RECT -11.530 83.880 -11.270 84.140 ;
        RECT -10.400 83.840 -10.140 84.100 ;
        RECT -13.170 83.200 -12.910 83.460 ;
        RECT -12.070 83.200 -11.810 83.460 ;
        RECT -10.970 83.200 -10.710 83.460 ;
        RECT -13.170 81.830 -12.910 82.090 ;
        RECT -12.070 81.830 -11.810 82.090 ;
        RECT -10.970 81.830 -10.710 82.090 ;
        RECT -13.720 81.100 -13.460 81.360 ;
        RECT -12.620 81.100 -12.360 81.360 ;
        RECT -11.530 81.100 -11.270 81.360 ;
        RECT -13.730 79.760 -13.470 80.020 ;
        RECT -12.620 79.750 -12.360 80.010 ;
        RECT -11.530 79.730 -11.270 79.990 ;
        RECT -17.820 78.860 -17.450 79.230 ;
        RECT -13.170 79.060 -12.910 79.320 ;
        RECT -12.070 79.050 -11.810 79.310 ;
        RECT -10.980 79.050 -10.720 79.310 ;
        RECT -10.280 78.440 -10.020 78.800 ;
        RECT -14.830 73.200 -14.540 73.490 ;
        RECT -10.370 76.750 -10.110 77.010 ;
        RECT -13.680 76.310 -13.420 76.570 ;
        RECT -12.580 76.320 -12.320 76.580 ;
        RECT -11.490 76.320 -11.230 76.580 ;
        RECT -10.360 76.280 -10.100 76.540 ;
        RECT -13.130 75.640 -12.870 75.900 ;
        RECT -12.030 75.640 -11.770 75.900 ;
        RECT -10.930 75.640 -10.670 75.900 ;
        RECT -13.130 74.270 -12.870 74.530 ;
        RECT -12.030 74.270 -11.770 74.530 ;
        RECT -10.930 74.270 -10.670 74.530 ;
        RECT -13.680 73.540 -13.420 73.800 ;
        RECT -12.580 73.540 -12.320 73.800 ;
        RECT -11.490 73.540 -11.230 73.800 ;
        RECT -7.380 112.780 -7.120 113.040 ;
        RECT -7.380 111.860 -7.120 112.120 ;
        RECT -7.410 110.940 -7.150 111.200 ;
        RECT 9.010 113.000 9.340 113.330 ;
        RECT 8.440 111.520 8.770 111.850 ;
        RECT -6.770 109.850 -6.510 110.110 ;
        RECT 7.800 109.920 8.130 110.250 ;
        RECT 7.160 109.350 7.490 109.680 ;
        RECT -6.760 108.890 -6.500 109.150 ;
        RECT -6.770 107.930 -6.510 108.190 ;
        RECT -7.410 90.270 -7.150 90.530 ;
        RECT -8.030 89.120 -7.770 89.380 ;
        RECT -8.450 86.510 -8.190 86.770 ;
        RECT -8.010 80.820 -7.750 81.240 ;
        RECT -8.050 78.440 -7.790 78.800 ;
        RECT 6.550 107.780 6.880 108.110 ;
        RECT 5.920 106.250 6.250 106.580 ;
        RECT 5.360 104.680 5.690 105.010 ;
        RECT 4.740 99.210 5.070 99.540 ;
        RECT 4.110 97.620 4.440 97.950 ;
        RECT 3.490 96.070 3.820 96.400 ;
        RECT 2.890 94.590 3.220 94.920 ;
        RECT 2.250 89.420 2.580 89.750 ;
        RECT 1.580 87.850 1.910 88.180 ;
        RECT -6.770 85.940 -6.510 86.200 ;
        RECT 0.960 86.210 1.290 86.540 ;
        RECT -7.430 74.810 -7.170 75.140 ;
        RECT -8.460 73.190 -8.170 73.480 ;
        RECT -13.690 72.200 -13.430 72.460 ;
        RECT -12.580 72.190 -12.320 72.450 ;
        RECT -11.490 72.170 -11.230 72.430 ;
        RECT -9.620 72.180 -9.020 72.780 ;
        RECT -13.130 71.500 -12.870 71.760 ;
        RECT -12.030 71.490 -11.770 71.750 ;
        RECT -10.940 71.490 -10.680 71.750 ;
        RECT 0.280 84.770 0.610 85.100 ;
        RECT -3.760 80.410 -3.180 81.120 ;
        RECT -6.840 67.250 -6.580 67.590 ;
        RECT -25.750 66.310 -25.360 66.700 ;
        RECT -126.950 58.020 -124.870 61.250 ;
        RECT 0.250 60.940 0.680 61.370 ;
        RECT 0.900 60.150 1.330 60.580 ;
        RECT 1.570 59.470 1.970 59.870 ;
        RECT 1.400 58.530 1.910 59.040 ;
        RECT 10.930 113.710 11.190 113.970 ;
        RECT 10.930 112.160 11.190 112.420 ;
        RECT 17.890 116.200 18.150 116.460 ;
        RECT 13.030 114.550 13.290 114.810 ;
        RECT 13.030 113.000 13.290 113.260 ;
        RECT 13.030 111.450 13.290 111.710 ;
        RECT 15.070 115.380 15.330 115.640 ;
        RECT 17.890 114.650 18.150 114.910 ;
        RECT 15.070 113.830 15.330 114.090 ;
        RECT 17.890 113.100 18.150 113.360 ;
        RECT 15.070 112.280 15.330 112.540 ;
        RECT 17.890 111.550 18.150 111.810 ;
        RECT 10.930 110.610 11.190 110.870 ;
        RECT 15.070 110.730 15.330 110.990 ;
        RECT 10.930 108.790 11.190 109.050 ;
        RECT 10.930 107.240 11.190 107.500 ;
        RECT 10.930 105.690 11.190 105.950 ;
        RECT 10.930 104.140 11.190 104.400 ;
        RECT 13.030 107.950 13.290 108.210 ;
        RECT 13.030 106.400 13.290 106.660 ;
        RECT 13.030 104.850 13.290 105.110 ;
        RECT 15.070 108.670 15.330 108.930 ;
        RECT 17.890 107.850 18.150 108.110 ;
        RECT 15.070 107.120 15.330 107.380 ;
        RECT 17.890 106.300 18.150 106.560 ;
        RECT 15.070 105.570 15.330 105.830 ;
        RECT 17.890 104.750 18.150 105.010 ;
        RECT 15.070 104.020 15.330 104.280 ;
        RECT 13.030 103.300 13.290 103.560 ;
        RECT 85.090 133.240 85.610 133.760 ;
        RECT 115.680 140.350 116.030 141.110 ;
        RECT 117.390 140.290 118.090 140.910 ;
        RECT 140.840 141.150 143.830 141.500 ;
        RECT 146.040 141.150 148.070 141.480 ;
        RECT 114.650 135.060 115.070 138.230 ;
        RECT 37.070 125.060 38.420 125.480 ;
        RECT 31.650 122.420 32.600 122.830 ;
        RECT 34.660 122.430 35.100 122.870 ;
        RECT 28.910 118.650 29.170 118.910 ;
        RECT 27.030 115.120 27.290 115.380 ;
        RECT 32.500 117.740 32.760 118.000 ;
        RECT 29.370 116.720 29.630 116.980 ;
        RECT 29.790 114.630 30.050 114.890 ;
        RECT 30.850 114.150 31.110 114.410 ;
        RECT 24.520 110.050 24.780 110.310 ;
        RECT 24.370 109.090 24.630 109.350 ;
        RECT 31.630 109.500 31.890 109.760 ;
        RECT 35.670 118.660 35.930 118.920 ;
        RECT 35.230 117.750 35.490 118.010 ;
        RECT 31.660 109.070 31.920 109.330 ;
        RECT 23.430 107.980 23.690 108.240 ;
        RECT 23.430 107.380 23.690 107.640 ;
        RECT 26.570 106.700 26.830 106.960 ;
        RECT 30.570 108.550 30.830 108.810 ;
        RECT 30.570 107.450 30.830 107.710 ;
        RECT 31.660 106.930 31.920 107.190 ;
        RECT 32.490 107.050 32.760 107.320 ;
        RECT 24.370 106.330 24.630 106.590 ;
        RECT 31.660 106.140 31.920 106.400 ;
        RECT 24.520 105.320 24.780 105.580 ;
        RECT 30.570 105.620 30.830 105.880 ;
        RECT 31.660 105.810 31.920 106.070 ;
        RECT 30.570 104.520 30.830 104.780 ;
        RECT 31.660 104.000 31.920 104.260 ;
        RECT 17.890 103.200 18.150 103.460 ;
        RECT 40.460 122.390 40.900 122.830 ;
        RECT 48.790 123.420 49.070 123.860 ;
        RECT 45.010 116.760 46.230 117.020 ;
        RECT 41.770 116.110 42.030 116.370 ;
        RECT 48.100 115.570 48.360 115.830 ;
        RECT 50.440 118.660 50.700 118.920 ;
        RECT 49.550 117.790 49.810 118.050 ;
        RECT 113.680 133.240 114.200 133.760 ;
        RECT 144.270 140.350 144.620 141.110 ;
        RECT 145.980 140.290 146.680 140.910 ;
        RECT 169.430 141.150 172.420 141.500 ;
        RECT 174.630 141.150 176.660 141.480 ;
        RECT 143.240 135.060 143.660 138.230 ;
        RECT 142.270 133.240 142.790 133.760 ;
        RECT 172.860 140.350 173.210 141.110 ;
        RECT 174.570 140.290 175.270 140.910 ;
        RECT 198.020 141.150 201.010 141.500 ;
        RECT 171.830 135.060 172.250 138.230 ;
        RECT 170.860 133.240 171.380 133.760 ;
        RECT 201.450 140.350 201.800 141.110 ;
        RECT 200.420 135.060 200.840 138.230 ;
        RECT 199.450 133.240 199.970 133.760 ;
        RECT 56.960 127.760 57.330 128.130 ;
        RECT 53.110 119.370 53.370 119.640 ;
        RECT 49.550 113.580 49.810 113.840 ;
        RECT 50.570 113.590 50.830 113.850 ;
        RECT 54.650 114.680 54.910 114.940 ;
        RECT 53.320 113.470 53.750 113.900 ;
        RECT 54.260 113.150 54.520 113.410 ;
        RECT 53.550 112.320 53.810 112.580 ;
        RECT 54.250 111.460 54.510 111.720 ;
        RECT 34.070 109.070 34.330 109.330 ;
        RECT 34.070 106.930 34.330 107.190 ;
        RECT 34.070 106.140 34.330 106.400 ;
        RECT 34.070 104.000 34.330 104.260 ;
        RECT 34.810 103.630 35.070 103.890 ;
        RECT 50.770 110.050 51.030 110.310 ;
        RECT 50.920 109.090 51.180 109.350 ;
        RECT 51.860 107.980 52.120 108.240 ;
        RECT 51.860 107.380 52.120 107.640 ;
        RECT 54.650 109.950 54.910 110.210 ;
        RECT 57.780 124.300 58.150 124.670 ;
        RECT 56.640 111.350 56.900 111.610 ;
        RECT 52.800 107.700 53.060 107.960 ;
        RECT 48.770 106.690 49.030 106.950 ;
        RECT 50.520 106.710 50.780 106.970 ;
        RECT 50.920 106.330 51.180 106.590 ;
        RECT 51.500 106.430 51.760 106.690 ;
        RECT 50.670 105.880 50.930 106.140 ;
        RECT 51.450 105.780 51.710 106.040 ;
        RECT 49.560 105.350 49.820 105.610 ;
        RECT 50.770 105.320 51.030 105.580 ;
        RECT 50.730 104.870 50.990 105.130 ;
        RECT 51.450 104.950 51.710 105.210 ;
        RECT 50.290 104.070 50.550 104.330 ;
        RECT 40.510 103.570 40.770 103.830 ;
        RECT 53.750 106.480 54.010 106.740 ;
        RECT 51.500 104.300 51.760 104.560 ;
        RECT 39.960 102.870 40.220 103.130 ;
        RECT 39.960 102.320 40.220 102.580 ;
        RECT 29.130 100.410 29.410 100.690 ;
        RECT 39.960 101.440 40.220 101.700 ;
        RECT 10.930 98.660 11.190 98.920 ;
        RECT 10.930 97.110 11.190 97.370 ;
        RECT 10.930 95.560 11.190 95.820 ;
        RECT 10.930 94.010 11.190 94.270 ;
        RECT 13.030 97.820 13.290 98.080 ;
        RECT 13.030 96.270 13.290 96.530 ;
        RECT 13.030 94.720 13.290 94.980 ;
        RECT 15.070 98.540 15.330 98.800 ;
        RECT 31.660 99.000 31.920 99.260 ;
        RECT 17.890 97.720 18.150 97.980 ;
        RECT 15.070 96.990 15.330 97.250 ;
        RECT 17.890 96.170 18.150 96.430 ;
        RECT 15.070 95.440 15.330 95.700 ;
        RECT 17.890 94.620 18.150 94.880 ;
        RECT 15.070 93.890 15.330 94.150 ;
        RECT 13.030 93.170 13.290 93.430 ;
        RECT 30.570 98.480 30.830 98.740 ;
        RECT 30.570 97.380 30.830 97.640 ;
        RECT 31.660 96.860 31.920 97.120 ;
        RECT 31.660 96.070 31.920 96.330 ;
        RECT 30.570 95.550 30.830 95.810 ;
        RECT 30.570 94.450 30.830 94.710 ;
        RECT 31.660 93.930 31.920 94.190 ;
        RECT 17.890 93.070 18.150 93.330 ;
        RECT 21.760 92.220 22.020 92.630 ;
        RECT 27.260 93.050 27.520 93.310 ;
        RECT 27.260 92.500 27.520 92.760 ;
        RECT 27.260 91.620 27.520 91.880 ;
        RECT 27.260 91.070 27.520 91.330 ;
        RECT 27.260 90.040 27.520 90.300 ;
        RECT 10.930 88.890 11.190 89.150 ;
        RECT 10.930 87.340 11.190 87.600 ;
        RECT 10.930 85.790 11.190 86.050 ;
        RECT 10.930 84.240 11.190 84.500 ;
        RECT 13.030 88.050 13.290 88.310 ;
        RECT 13.030 86.500 13.290 86.760 ;
        RECT 13.030 84.950 13.290 85.210 ;
        RECT 15.070 88.770 15.330 89.030 ;
        RECT 17.890 87.950 18.150 88.210 ;
        RECT 15.070 87.220 15.330 87.480 ;
        RECT 17.890 86.400 18.150 86.660 ;
        RECT 15.070 85.670 15.330 85.930 ;
        RECT 17.890 84.850 18.150 85.110 ;
        RECT 15.070 84.120 15.330 84.380 ;
        RECT 13.030 83.400 13.290 83.660 ;
        RECT 27.260 89.490 27.520 89.750 ;
        RECT 34.070 99.000 34.330 99.260 ;
        RECT 39.960 100.890 40.220 101.150 ;
        RECT 40.510 101.050 40.770 101.310 ;
        RECT 39.960 99.860 40.220 100.120 ;
        RECT 39.960 99.310 40.220 99.570 ;
        RECT 40.650 99.390 40.910 99.650 ;
        RECT 40.880 98.830 41.140 99.090 ;
        RECT 34.070 96.860 34.330 97.120 ;
        RECT 39.960 98.440 40.220 98.700 ;
        RECT 39.960 97.890 40.220 98.150 ;
        RECT 51.500 103.470 51.760 103.730 ;
        RECT 51.450 102.820 51.710 103.080 ;
        RECT 51.450 101.990 51.710 102.250 ;
        RECT 46.480 99.840 46.740 100.100 ;
        RECT 50.950 101.180 51.220 101.440 ;
        RECT 51.500 101.340 51.760 101.600 ;
        RECT 53.800 104.260 54.060 104.520 ;
        RECT 53.790 103.540 54.050 103.800 ;
        RECT 53.710 101.290 53.970 101.550 ;
        RECT 44.810 98.790 45.070 99.050 ;
        RECT 58.550 119.590 58.920 119.960 ;
        RECT 56.970 100.390 57.340 100.760 ;
        RECT 57.740 99.800 58.110 100.170 ;
        RECT 55.890 98.790 56.150 99.050 ;
        RECT 65.100 118.540 65.600 119.040 ;
        RECT 61.880 116.980 62.380 117.480 ;
        RECT 62.830 117.470 63.330 117.970 ;
        RECT 63.910 117.940 64.410 118.440 ;
        RECT 59.430 114.520 59.800 114.890 ;
        RECT 60.740 102.870 61.000 103.130 ;
        RECT 60.740 102.320 61.000 102.580 ;
        RECT 60.740 101.440 61.000 101.700 ;
        RECT 60.740 100.890 61.000 101.150 ;
        RECT 60.740 99.860 61.000 100.120 ;
        RECT 58.480 97.470 58.850 97.840 ;
        RECT 34.070 96.070 34.330 96.330 ;
        RECT 30.530 89.340 30.790 89.600 ;
        RECT 28.300 88.970 28.560 89.230 ;
        RECT 31.660 89.240 31.920 89.500 ;
        RECT 34.070 93.930 34.330 94.190 ;
        RECT 34.070 89.240 34.330 89.500 ;
        RECT 26.160 88.500 26.420 88.760 ;
        RECT 27.260 88.620 27.520 88.880 ;
        RECT 17.890 83.300 18.150 83.560 ;
        RECT 19.580 83.370 19.840 83.630 ;
        RECT 19.040 83.000 19.330 83.290 ;
        RECT 14.600 82.490 14.910 82.800 ;
        RECT 27.260 88.070 27.520 88.330 ;
        RECT 27.240 87.790 27.500 88.050 ;
        RECT 30.570 88.720 30.830 88.980 ;
        RECT 32.320 88.950 32.590 89.210 ;
        RECT 30.510 88.290 30.770 88.550 ;
        RECT 30.570 87.620 30.830 87.880 ;
        RECT 27.220 86.780 27.480 87.040 ;
        RECT 60.050 99.390 60.310 99.650 ;
        RECT 60.740 99.310 61.000 99.570 ;
        RECT 59.820 98.830 60.080 99.090 ;
        RECT 60.740 98.440 61.000 98.700 ;
        RECT 60.740 97.890 61.000 98.150 ;
        RECT 59.410 92.220 59.780 92.630 ;
        RECT 38.610 89.140 38.870 89.400 ;
        RECT 38.760 88.460 39.020 88.720 ;
        RECT 31.660 87.100 31.920 87.360 ;
        RECT 26.790 85.720 27.050 85.980 ;
        RECT 26.190 83.410 26.450 83.670 ;
        RECT 27.170 84.740 27.430 85.000 ;
        RECT 27.220 83.890 27.480 84.150 ;
        RECT 27.220 83.400 27.480 83.660 ;
        RECT 24.790 83.000 25.050 83.260 ;
        RECT 26.760 83.080 27.020 83.340 ;
        RECT 18.410 81.780 18.830 82.200 ;
        RECT 14.560 80.820 14.980 81.240 ;
        RECT 20.470 82.460 20.730 82.720 ;
        RECT 30.510 86.410 30.770 86.670 ;
        RECT 31.660 86.310 31.920 86.570 ;
        RECT 30.570 85.790 30.830 86.050 ;
        RECT 30.350 85.230 30.610 85.490 ;
        RECT 30.570 84.690 30.830 84.950 ;
        RECT 31.660 84.170 31.920 84.430 ;
        RECT 29.000 83.020 29.260 83.280 ;
        RECT 27.800 81.770 28.130 82.100 ;
        RECT 34.070 87.100 34.330 87.360 ;
        RECT 38.760 87.570 39.020 87.830 ;
        RECT 38.610 86.890 38.870 87.150 ;
        RECT 34.070 86.310 34.330 86.570 ;
        RECT 38.610 86.370 38.870 86.630 ;
        RECT 38.760 85.690 39.020 85.950 ;
        RECT 34.070 84.170 34.330 84.430 ;
        RECT 38.760 84.800 39.020 85.060 ;
        RECT 38.610 84.120 38.870 84.380 ;
        RECT 46.040 88.480 46.300 88.740 ;
        RECT 45.520 87.550 45.780 87.810 ;
        RECT 45.050 85.710 45.310 85.970 ;
        RECT 40.890 85.240 41.160 85.510 ;
        RECT 37.840 83.330 38.190 83.680 ;
        RECT 30.990 82.600 31.250 82.860 ;
        RECT 35.030 82.570 35.300 82.840 ;
        RECT 28.950 81.700 29.290 82.040 ;
        RECT 44.550 84.780 44.810 85.040 ;
        RECT 37.880 81.560 38.140 81.880 ;
        RECT 43.870 81.780 44.130 82.120 ;
        RECT 19.090 80.730 19.410 81.050 ;
        RECT 39.300 80.850 39.680 81.230 ;
        RECT 19.240 77.600 19.500 77.860 ;
        RECT 20.330 77.600 20.590 77.860 ;
        RECT 21.430 77.590 21.690 77.850 ;
        RECT 25.550 77.590 25.810 77.850 ;
        RECT 26.650 77.600 26.910 77.860 ;
        RECT 27.740 77.600 28.000 77.860 ;
        RECT 29.050 77.630 29.310 77.890 ;
        RECT 30.140 77.630 30.400 77.890 ;
        RECT 31.240 77.620 31.500 77.880 ;
        RECT 35.360 77.620 35.620 77.880 ;
        RECT 36.460 77.630 36.720 77.890 ;
        RECT 37.550 77.630 37.810 77.890 ;
        RECT 41.100 77.600 41.360 77.860 ;
        RECT 42.200 77.610 42.460 77.870 ;
        RECT 43.290 77.610 43.550 77.870 ;
        RECT 19.790 76.920 20.050 77.180 ;
        RECT 20.880 76.900 21.140 77.160 ;
        RECT 21.990 76.890 22.250 77.150 ;
        RECT 19.790 75.550 20.050 75.810 ;
        RECT 20.880 75.550 21.140 75.810 ;
        RECT 21.980 75.550 22.240 75.810 ;
        RECT 19.190 74.950 19.650 75.410 ;
        RECT 19.230 74.820 19.490 74.950 ;
        RECT 20.330 74.820 20.590 75.080 ;
        RECT 21.430 74.820 21.690 75.080 ;
        RECT 19.230 73.450 19.490 73.710 ;
        RECT 20.330 73.450 20.590 73.710 ;
        RECT 21.430 73.450 21.690 73.710 ;
        RECT 18.660 72.810 18.920 73.070 ;
        RECT 19.790 72.770 20.050 73.030 ;
        RECT 20.880 72.770 21.140 73.030 ;
        RECT 21.980 72.780 22.240 73.040 ;
        RECT 18.670 72.340 18.930 72.600 ;
        RECT 23.110 75.980 23.390 76.260 ;
        RECT 23.850 76.000 24.130 76.280 ;
        RECT 24.990 76.890 25.250 77.150 ;
        RECT 26.100 76.900 26.360 77.160 ;
        RECT 27.190 76.920 27.450 77.180 ;
        RECT 25.000 75.550 25.260 75.810 ;
        RECT 26.100 75.550 26.360 75.810 ;
        RECT 27.190 75.550 27.450 75.810 ;
        RECT 29.600 76.950 29.860 77.210 ;
        RECT 30.690 76.930 30.950 77.190 ;
        RECT 31.800 76.920 32.060 77.180 ;
        RECT 29.600 75.580 29.860 75.840 ;
        RECT 30.690 75.580 30.950 75.840 ;
        RECT 31.790 75.580 32.050 75.840 ;
        RECT 25.550 74.820 25.810 75.080 ;
        RECT 26.650 74.820 26.910 75.080 ;
        RECT 27.750 74.820 28.010 75.080 ;
        RECT 29.040 74.850 29.300 75.110 ;
        RECT 30.140 74.850 30.400 75.110 ;
        RECT 31.240 74.850 31.500 75.110 ;
        RECT 27.570 74.000 28.030 74.460 ;
        RECT 25.550 73.450 25.810 73.710 ;
        RECT 26.650 73.450 26.910 73.710 ;
        RECT 27.750 73.450 28.010 73.710 ;
        RECT 29.040 73.570 29.300 73.740 ;
        RECT 28.470 73.070 28.730 73.100 ;
        RECT 25.000 72.780 25.260 73.040 ;
        RECT 26.100 72.770 26.360 73.030 ;
        RECT 27.190 72.770 27.450 73.030 ;
        RECT 28.320 72.840 28.730 73.070 ;
        RECT 29.000 73.110 29.460 73.570 ;
        RECT 30.140 73.480 30.400 73.740 ;
        RECT 31.240 73.480 31.500 73.740 ;
        RECT 28.320 72.810 28.580 72.840 ;
        RECT 29.600 72.800 29.860 73.060 ;
        RECT 30.690 72.800 30.950 73.060 ;
        RECT 31.790 72.810 32.050 73.070 ;
        RECT 28.480 72.600 28.740 72.630 ;
        RECT 28.310 72.370 28.740 72.600 ;
        RECT 28.310 72.340 28.570 72.370 ;
        RECT 32.920 75.980 33.200 76.260 ;
        RECT 34.800 76.920 35.060 77.180 ;
        RECT 35.910 76.930 36.170 77.190 ;
        RECT 37.000 76.950 37.260 77.210 ;
        RECT 34.810 75.580 35.070 75.840 ;
        RECT 35.910 75.580 36.170 75.840 ;
        RECT 37.000 75.580 37.260 75.840 ;
        RECT 40.540 76.900 40.800 77.160 ;
        RECT 41.650 76.910 41.910 77.170 ;
        RECT 42.740 76.930 43.000 77.190 ;
        RECT 73.910 115.600 75.190 116.880 ;
        RECT 74.400 112.160 74.660 112.580 ;
        RECT 80.890 114.680 81.150 114.940 ;
        RECT 78.230 113.440 78.490 113.870 ;
        RECT 81.040 113.720 81.300 113.980 ;
        RECT 101.430 128.670 104.660 130.730 ;
        RECT 130.020 123.780 132.080 127.080 ;
        RECT 85.180 120.930 85.890 121.640 ;
        RECT 81.980 112.610 82.240 112.870 ;
        RECT 81.980 112.010 82.240 112.270 ;
        RECT 78.910 111.350 79.170 111.610 ;
        RECT 80.640 111.340 80.900 111.600 ;
        RECT 82.920 112.330 83.180 112.590 ;
        RECT 81.040 110.960 81.300 111.220 ;
        RECT 81.620 111.060 81.880 111.320 ;
        RECT 80.790 110.510 81.050 110.770 ;
        RECT 81.570 110.410 81.830 110.670 ;
        RECT 79.210 109.950 79.470 110.210 ;
        RECT 79.680 109.980 79.940 110.240 ;
        RECT 80.780 109.950 81.150 110.210 ;
        RECT 70.400 108.960 70.800 109.360 ;
        RECT 64.860 105.670 65.120 105.930 ;
        RECT 65.010 96.260 65.510 96.760 ;
        RECT 63.930 91.070 64.430 91.540 ;
        RECT 62.800 85.880 63.300 86.380 ;
        RECT 61.750 80.580 62.250 81.080 ;
        RECT 46.020 79.070 46.280 79.570 ;
        RECT 45.480 78.170 45.740 78.670 ;
        RECT 45.010 77.270 45.270 77.770 ;
        RECT 40.550 75.560 40.810 75.820 ;
        RECT 41.650 75.560 41.910 75.820 ;
        RECT 42.740 75.560 43.000 75.820 ;
        RECT 35.360 74.850 35.620 75.110 ;
        RECT 36.460 74.850 36.720 75.110 ;
        RECT 44.530 76.370 44.790 76.870 ;
        RECT 37.560 74.850 37.820 75.110 ;
        RECT 41.100 74.830 41.360 75.090 ;
        RECT 42.200 74.830 42.460 75.090 ;
        RECT 43.300 74.830 43.560 75.090 ;
        RECT 35.360 73.480 35.620 73.740 ;
        RECT 36.460 73.480 36.720 73.740 ;
        RECT 37.560 73.480 37.820 73.740 ;
        RECT 41.100 73.460 41.360 73.720 ;
        RECT 34.810 72.810 35.070 73.070 ;
        RECT 35.910 72.800 36.170 73.060 ;
        RECT 37.000 72.800 37.260 73.060 ;
        RECT 42.200 73.460 42.460 73.720 ;
        RECT 43.300 73.460 43.560 73.720 ;
        RECT 38.130 72.840 38.390 73.100 ;
        RECT 40.550 72.790 40.810 73.050 ;
        RECT 41.650 72.780 41.910 73.040 ;
        RECT 42.740 72.780 43.000 73.040 ;
        RECT 37.390 72.200 37.850 72.660 ;
        RECT 38.120 72.370 38.380 72.630 ;
        RECT 11.320 69.970 11.580 71.090 ;
        RECT 23.430 71.030 24.550 71.050 ;
        RECT 22.690 69.930 24.550 71.030 ;
        RECT 22.690 69.910 23.810 69.930 ;
        RECT 32.500 69.880 34.360 71.070 ;
        RECT 9.640 65.680 9.970 66.010 ;
        RECT 9.020 65.060 9.350 65.390 ;
        RECT 8.390 64.430 8.720 64.760 ;
        RECT 7.790 63.800 8.120 64.130 ;
        RECT 7.150 63.120 7.480 63.450 ;
        RECT 6.550 62.500 6.880 62.830 ;
        RECT 5.950 61.860 6.280 62.190 ;
        RECT 5.370 61.290 5.700 61.620 ;
        RECT 4.790 60.600 5.120 60.930 ;
        RECT 4.140 59.960 4.470 60.290 ;
        RECT 3.500 59.310 3.830 59.650 ;
        RECT 2.920 58.670 3.290 59.040 ;
        RECT 43.870 72.820 44.130 73.080 ;
        RECT 71.380 108.320 71.740 108.680 ;
        RECT 70.660 105.670 70.920 105.930 ;
        RECT 67.990 83.100 68.490 83.600 ;
        RECT 65.120 74.990 65.620 75.490 ;
        RECT 63.930 74.040 64.430 74.500 ;
        RECT 62.800 73.170 63.300 73.630 ;
        RECT 43.860 72.350 44.120 72.610 ;
        RECT 61.870 72.260 62.370 72.720 ;
        RECT 67.410 69.970 68.350 71.090 ;
        RECT 43.200 66.340 43.530 66.670 ;
        RECT 72.300 105.950 72.690 106.340 ;
        RECT 73.130 105.390 73.510 105.650 ;
        RECT 70.460 65.150 70.860 65.550 ;
        RECT 69.980 64.220 70.240 64.480 ;
        RECT 71.370 64.350 71.760 64.740 ;
        RECT 72.300 63.530 72.690 63.920 ;
        RECT 77.860 108.970 78.120 109.230 ;
        RECT 80.850 109.500 81.110 109.760 ;
        RECT 77.860 108.440 78.120 108.700 ;
        RECT 80.130 109.040 80.390 109.300 ;
        RECT 80.410 108.700 80.670 108.960 ;
        RECT 80.130 108.370 80.390 108.630 ;
        RECT 81.570 109.580 81.830 109.840 ;
        RECT 81.140 109.030 81.400 109.290 ;
        RECT 83.870 111.110 84.130 111.370 ;
        RECT 81.620 108.930 81.880 109.190 ;
        RECT 81.140 108.380 81.400 108.640 ;
        RECT 79.210 107.460 79.470 107.720 ;
        RECT 81.620 108.100 81.880 108.360 ;
        RECT 80.780 107.460 81.040 107.720 ;
        RECT 81.570 107.450 81.830 107.710 ;
        RECT 79.210 106.930 79.470 107.190 ;
        RECT 80.780 106.930 81.040 107.190 ;
        RECT 77.860 105.950 78.120 106.210 ;
        RECT 81.570 106.620 81.830 106.880 ;
        RECT 77.860 105.420 78.120 105.680 ;
        RECT 80.130 106.020 80.390 106.280 ;
        RECT 81.140 106.080 81.400 106.270 ;
        RECT 81.050 106.010 81.400 106.080 ;
        RECT 81.050 105.820 81.310 106.010 ;
        RECT 81.620 105.970 81.880 106.230 ;
        RECT 80.130 105.350 80.390 105.610 ;
        RECT 81.140 105.360 81.400 105.620 ;
        RECT 83.920 108.890 84.180 109.150 ;
        RECT 83.910 108.170 84.170 108.430 ;
        RECT 83.830 105.920 84.090 106.180 ;
        RECT 79.210 104.440 79.470 104.700 ;
        RECT 80.780 104.440 81.040 104.700 ;
        RECT 158.610 119.530 161.840 121.590 ;
        RECT 212.820 128.730 213.580 129.080 ;
        RECT 207.530 127.700 210.700 128.120 ;
        RECT 205.710 126.730 206.230 127.250 ;
        RECT 187.200 115.120 190.430 117.170 ;
        RECT 213.620 125.300 213.970 128.290 ;
        RECT 201.540 114.480 203.530 117.710 ;
        RECT 84.990 101.140 85.700 101.850 ;
        RECT 109.800 113.500 112.020 113.820 ;
        RECT 212.760 101.850 213.380 102.550 ;
        RECT 213.620 101.910 213.950 103.940 ;
        RECT 212.820 100.140 213.580 100.490 ;
        RECT 207.530 99.110 210.700 99.530 ;
        RECT 205.710 98.140 206.230 98.660 ;
        RECT 213.620 96.710 213.970 99.700 ;
        RECT 192.990 85.890 195.080 89.120 ;
        RECT 80.790 83.090 81.300 83.600 ;
        RECT 109.640 83.110 113.920 84.200 ;
        RECT 74.760 69.460 75.020 69.720 ;
        RECT 74.760 68.790 75.020 69.050 ;
        RECT 74.880 67.550 75.140 67.810 ;
        RECT 74.880 65.940 75.140 66.200 ;
        RECT 74.870 64.330 75.130 64.590 ;
        RECT 73.120 62.740 73.500 63.120 ;
        RECT 74.870 62.710 75.130 62.970 ;
        RECT 74.870 61.100 75.130 61.360 ;
        RECT 74.500 59.500 74.760 59.760 ;
        RECT 74.880 57.900 75.140 58.160 ;
        RECT 71.670 56.230 71.930 56.490 ;
        RECT 72.610 56.230 72.870 56.490 ;
        RECT 73.560 56.170 73.820 56.430 ;
        RECT 74.870 56.310 75.130 56.570 ;
        RECT -150.360 45.450 -150.030 47.480 ;
        RECT -149.790 45.390 -149.170 46.090 ;
        RECT -149.990 43.680 -149.230 44.030 ;
        RECT -150.380 40.250 -150.030 43.240 ;
        RECT -147.110 42.650 -143.940 43.070 ;
        RECT -142.640 41.680 -142.120 42.200 ;
        RECT -122.320 29.430 -120.240 32.660 ;
        RECT -150.360 16.860 -150.030 18.890 ;
        RECT -149.790 16.800 -149.170 17.500 ;
        RECT -149.990 15.090 -149.230 15.440 ;
        RECT -150.380 11.660 -150.030 14.650 ;
        RECT -147.110 14.060 -143.940 14.480 ;
        RECT -142.640 13.090 -142.120 13.610 ;
        RECT -117.910 0.840 -115.830 4.070 ;
        RECT -150.360 -11.730 -150.030 -9.700 ;
        RECT -149.790 -11.790 -149.170 -11.090 ;
        RECT -149.990 -13.500 -149.230 -13.150 ;
        RECT -150.380 -16.930 -150.030 -13.940 ;
        RECT -147.110 -14.530 -143.940 -14.110 ;
        RECT -142.640 -15.500 -142.120 -14.980 ;
        RECT -113.570 -27.750 -111.490 -24.520 ;
        RECT -150.360 -40.320 -150.030 -38.290 ;
        RECT -149.790 -40.380 -149.170 -39.680 ;
        RECT -149.990 -42.090 -149.230 -41.740 ;
        RECT -150.380 -45.520 -150.030 -42.530 ;
        RECT -147.110 -43.120 -143.940 -42.700 ;
        RECT -142.640 -44.090 -142.120 -43.570 ;
        RECT -150.360 -68.910 -150.030 -66.880 ;
        RECT -149.790 -68.970 -149.170 -68.270 ;
        RECT -149.990 -70.680 -149.230 -70.330 ;
        RECT -150.380 -74.110 -150.030 -71.120 ;
        RECT -147.110 -71.710 -143.940 -71.290 ;
        RECT -142.640 -72.680 -142.120 -72.160 ;
        RECT 212.760 73.260 213.380 73.960 ;
        RECT 213.620 73.320 213.950 75.350 ;
        RECT 212.820 71.550 213.580 71.900 ;
        RECT 207.530 70.520 210.700 70.940 ;
        RECT 205.710 69.550 206.230 70.070 ;
        RECT 213.620 68.120 213.970 71.110 ;
        RECT 188.740 57.300 190.830 60.530 ;
        RECT 212.760 44.670 213.380 45.370 ;
        RECT 213.620 44.730 213.950 46.760 ;
        RECT 212.820 42.960 213.580 43.310 ;
        RECT 207.530 41.930 210.700 42.350 ;
        RECT 205.710 40.960 206.230 41.480 ;
        RECT 213.620 39.530 213.970 42.520 ;
        RECT 184.760 28.710 186.850 31.940 ;
        RECT 212.760 16.080 213.380 16.780 ;
        RECT 213.620 16.140 213.950 18.170 ;
        RECT 212.820 14.370 213.580 14.720 ;
        RECT 207.530 13.340 210.700 13.760 ;
        RECT 205.710 12.370 206.230 12.890 ;
        RECT 213.620 10.940 213.970 13.930 ;
        RECT 180.510 0.120 182.600 3.350 ;
        RECT 212.760 -12.510 213.380 -11.810 ;
        RECT 213.620 -12.450 213.950 -10.420 ;
        RECT 212.820 -14.220 213.580 -13.870 ;
        RECT 207.530 -15.250 210.700 -14.830 ;
        RECT 205.710 -16.220 206.230 -15.700 ;
        RECT 213.620 -17.650 213.970 -14.660 ;
        RECT 176.570 -28.470 178.660 -25.240 ;
        RECT 212.760 -41.100 213.380 -40.400 ;
        RECT 213.620 -41.040 213.950 -39.010 ;
        RECT 212.820 -42.810 213.580 -42.460 ;
        RECT 207.530 -43.840 210.700 -43.420 ;
        RECT 205.710 -44.810 206.230 -44.290 ;
        RECT 213.620 -46.240 213.970 -43.250 ;
        RECT 212.760 -69.690 213.380 -68.990 ;
        RECT 213.620 -69.630 213.950 -67.600 ;
        RECT -105.030 -84.930 -102.950 -81.700 ;
        RECT 108.820 -82.830 113.240 -78.410 ;
        RECT -150.360 -97.500 -150.030 -95.470 ;
        RECT -149.790 -97.560 -149.170 -96.860 ;
        RECT -149.990 -99.270 -149.230 -98.920 ;
        RECT -150.380 -102.700 -150.030 -99.710 ;
        RECT -147.110 -100.300 -143.940 -99.880 ;
        RECT -142.640 -101.270 -142.120 -100.750 ;
        RECT -150.360 -126.090 -150.030 -124.060 ;
        RECT -149.790 -126.150 -149.170 -125.450 ;
        RECT -149.990 -127.860 -149.230 -127.510 ;
        RECT -150.380 -131.290 -150.030 -128.300 ;
        RECT -147.110 -128.890 -143.940 -128.470 ;
        RECT -142.640 -129.860 -142.120 -129.340 ;
        RECT -96.410 -142.110 -94.330 -138.880 ;
        RECT -150.360 -154.680 -150.030 -152.650 ;
        RECT -149.790 -154.740 -149.170 -154.040 ;
        RECT -149.990 -156.450 -149.230 -156.100 ;
        RECT -150.380 -159.880 -150.030 -156.890 ;
        RECT -147.110 -157.480 -143.940 -157.060 ;
        RECT -142.640 -158.450 -142.120 -157.930 ;
        RECT -92.440 -170.700 -90.360 -167.470 ;
        RECT -150.360 -183.270 -150.030 -181.240 ;
        RECT -149.790 -183.330 -149.170 -182.630 ;
        RECT -149.990 -185.040 -149.230 -184.690 ;
        RECT -150.380 -188.470 -150.030 -185.480 ;
        RECT -147.110 -186.070 -143.940 -185.650 ;
        RECT -142.640 -187.040 -142.120 -186.520 ;
        RECT -88.000 -199.290 -85.920 -196.060 ;
        RECT -150.360 -211.860 -150.030 -209.830 ;
        RECT -149.790 -211.920 -149.170 -211.220 ;
        RECT -149.990 -213.630 -149.230 -213.280 ;
        RECT -150.380 -217.060 -150.030 -214.070 ;
        RECT -147.110 -214.660 -143.940 -214.240 ;
        RECT -142.640 -215.630 -142.120 -215.110 ;
        RECT -83.700 -227.880 -81.620 -224.650 ;
        RECT -150.360 -240.450 -150.030 -238.420 ;
        RECT -149.790 -240.510 -149.170 -239.810 ;
      LAYER met2 ;
        RECT 87.770 129.440 88.630 129.480 ;
        RECT 100.280 129.440 105.080 131.530 ;
        RECT 56.900 128.130 57.360 128.150 ;
        RECT 87.770 128.130 105.130 129.440 ;
        RECT -20.440 127.730 -20.120 127.780 ;
        RECT 56.900 127.760 105.130 128.130 ;
        RECT 56.900 127.740 57.360 127.760 ;
        RECT -23.300 127.490 -20.120 127.730 ;
        RECT -23.300 127.470 -22.980 127.490 ;
        RECT 87.770 127.380 105.130 127.760 ;
        RECT -97.040 125.380 -93.660 125.490 ;
        RECT 13.430 125.480 13.880 125.500 ;
        RECT 13.420 125.470 13.900 125.480 ;
        RECT 37.040 125.470 38.460 125.510 ;
        RECT -26.950 125.380 -26.270 125.390 ;
        RECT -97.450 124.510 -26.270 125.380 ;
        RECT 13.420 125.070 38.510 125.470 ;
        RECT 87.770 125.310 88.630 125.350 ;
        RECT 129.870 125.310 133.180 127.370 ;
        RECT 13.420 125.060 13.900 125.070 ;
        RECT 13.430 125.040 13.880 125.060 ;
        RECT 37.040 125.030 38.460 125.070 ;
        RECT 57.730 124.670 58.170 124.690 ;
        RECT 87.770 124.670 133.500 125.310 ;
        RECT -97.450 124.480 -23.290 124.510 ;
        RECT -97.450 124.220 -22.990 124.480 ;
        RECT 57.730 124.300 133.500 124.670 ;
        RECT 57.730 124.280 58.170 124.300 ;
        RECT -97.450 124.190 -23.290 124.220 ;
        RECT -97.450 123.130 -26.270 124.190 ;
        RECT -21.170 124.030 -20.860 124.260 ;
        RECT -24.260 123.930 -20.860 124.030 ;
        RECT -24.260 123.800 -20.880 123.930 ;
        RECT -24.260 123.770 -23.940 123.800 ;
        RECT 87.770 123.250 133.500 124.300 ;
        RECT -97.040 122.810 -93.660 123.130 ;
        RECT -26.950 123.070 -26.270 123.130 ;
        RECT -127.580 120.890 -124.940 122.070 ;
        RECT 85.150 121.490 85.920 121.640 ;
        RECT -24.340 121.070 85.920 121.490 ;
        RECT 85.150 120.930 85.920 121.070 ;
        RECT 87.740 121.230 88.600 121.260 ;
        RECT 158.260 121.230 162.190 121.680 ;
        RECT -27.400 120.890 -26.720 120.920 ;
        RECT -127.660 120.250 -26.720 120.890 ;
        RECT -18.480 120.250 -18.010 120.270 ;
        RECT -127.660 119.670 -18.010 120.250 ;
        RECT -127.660 119.430 -26.680 119.670 ;
        RECT -18.480 119.650 -18.010 119.670 ;
        RECT 58.510 119.960 58.930 119.980 ;
        RECT 87.740 119.960 162.190 121.230 ;
        RECT 58.510 119.590 162.190 119.960 ;
        RECT 58.510 119.570 58.930 119.590 ;
        RECT -127.660 118.640 -26.720 119.430 ;
        RECT 87.740 119.170 162.190 119.590 ;
        RECT 87.740 119.160 88.600 119.170 ;
        RECT 158.260 119.160 162.190 119.170 ;
        RECT -139.810 116.550 -136.920 118.510 ;
        RECT -127.580 118.470 -124.940 118.640 ;
        RECT -27.400 118.600 -26.720 118.640 ;
        RECT 29.340 116.950 29.660 116.990 ;
        RECT 44.990 116.950 46.270 117.050 ;
        RECT 19.260 116.610 19.370 116.810 ;
        RECT 29.340 116.740 46.270 116.950 ;
        RECT 29.340 116.710 29.660 116.740 ;
        RECT -27.720 116.550 -26.450 116.560 ;
        RECT -139.840 115.100 -26.450 116.550 ;
        RECT 17.860 116.410 18.180 116.460 ;
        RECT 10.570 115.630 10.660 115.950 ;
        RECT 13.030 115.590 13.290 116.390 ;
        RECT 17.860 116.210 19.490 116.410 ;
        RECT 17.860 116.200 18.180 116.210 ;
        RECT 48.070 115.800 48.380 115.860 ;
        RECT 19.770 115.790 48.380 115.800 ;
        RECT 15.030 115.590 15.370 115.650 ;
        RECT 19.440 115.600 48.380 115.790 ;
        RECT 19.440 115.590 20.020 115.600 ;
        RECT 10.760 115.230 11.220 115.550 ;
        RECT 12.930 115.370 15.370 115.590 ;
        RECT 48.070 115.540 48.380 115.600 ;
        RECT 27.000 115.330 27.320 115.380 ;
        RECT -16.370 115.100 -16.070 115.110 ;
        RECT -6.780 115.100 -6.490 115.120 ;
        RECT -139.840 114.710 -6.460 115.100 ;
        RECT 19.260 115.060 19.370 115.260 ;
        RECT 22.000 115.130 27.370 115.330 ;
        RECT 17.860 114.860 18.180 114.910 ;
        RECT -139.840 114.690 -26.450 114.710 ;
        RECT -6.780 114.690 -6.490 114.710 ;
        RECT -27.720 114.680 -26.450 114.690 ;
        RECT 10.570 114.080 10.660 114.400 ;
        RECT 13.030 114.040 13.290 114.840 ;
        RECT 17.860 114.660 19.490 114.860 ;
        RECT 17.860 114.650 18.180 114.660 ;
        RECT 22.000 114.250 22.200 115.130 ;
        RECT 27.000 115.120 27.320 115.130 ;
        RECT 29.760 114.890 30.070 114.900 ;
        RECT 29.760 114.860 30.080 114.890 ;
        RECT 19.760 114.240 22.200 114.250 ;
        RECT 15.030 114.040 15.370 114.100 ;
        RECT 19.470 114.050 22.200 114.240 ;
        RECT 22.510 114.660 30.080 114.860 ;
        RECT 19.470 114.040 19.960 114.050 ;
        RECT 10.760 113.680 11.220 114.000 ;
        RECT 12.930 113.820 15.370 114.040 ;
        RECT 19.260 113.510 19.370 113.710 ;
        RECT 17.860 113.310 18.180 113.360 ;
        RECT -16.070 113.210 -15.700 113.220 ;
        RECT -17.860 112.980 -15.700 113.210 ;
        RECT -10.010 112.980 -9.700 113.070 ;
        RECT -17.860 112.850 -9.700 112.980 ;
        RECT -17.860 112.150 -17.240 112.850 ;
        RECT -16.070 112.810 -9.700 112.850 ;
        RECT -10.010 112.740 -9.700 112.810 ;
        RECT 10.570 112.530 10.660 112.850 ;
        RECT 13.030 112.490 13.290 113.290 ;
        RECT 17.860 113.110 19.490 113.310 ;
        RECT 17.860 113.100 18.180 113.110 ;
        RECT 22.510 112.700 22.710 114.660 ;
        RECT 29.760 114.630 30.080 114.660 ;
        RECT 29.760 114.620 30.070 114.630 ;
        RECT 30.820 114.380 31.140 114.420 ;
        RECT 19.760 112.690 22.710 112.700 ;
        RECT 15.030 112.490 15.370 112.550 ;
        RECT 19.470 112.500 22.710 112.690 ;
        RECT 23.060 114.180 31.220 114.380 ;
        RECT 19.470 112.490 19.970 112.500 ;
        RECT -16.070 112.150 -15.700 112.190 ;
        RECT -18.390 112.060 -15.700 112.150 ;
        RECT -10.010 112.060 -9.700 112.150 ;
        RECT 10.760 112.130 11.220 112.450 ;
        RECT 12.930 112.270 15.370 112.490 ;
        RECT -18.390 111.890 -9.700 112.060 ;
        RECT 19.260 111.960 19.370 112.160 ;
        RECT -18.390 111.780 -15.700 111.890 ;
        RECT -10.010 111.820 -9.700 111.890 ;
        RECT -18.390 111.670 -17.240 111.780 ;
        RECT 17.860 111.760 18.180 111.810 ;
        RECT -18.390 111.220 -17.280 111.670 ;
        RECT -16.070 111.220 -15.700 111.260 ;
        RECT -18.390 111.140 -15.700 111.220 ;
        RECT -10.010 111.140 -9.700 111.230 ;
        RECT -18.390 110.970 -9.700 111.140 ;
        RECT 10.570 110.980 10.660 111.300 ;
        RECT -18.390 110.850 -15.700 110.970 ;
        RECT -10.010 110.900 -9.700 110.970 ;
        RECT 13.030 110.940 13.290 111.740 ;
        RECT 17.860 111.560 19.490 111.760 ;
        RECT 17.860 111.550 18.180 111.560 ;
        RECT 23.060 111.150 23.260 114.180 ;
        RECT 30.820 114.140 31.140 114.180 ;
        RECT 54.230 111.570 54.540 111.760 ;
        RECT 56.610 111.570 56.930 111.630 ;
        RECT 54.230 111.510 63.980 111.570 ;
        RECT 78.880 111.510 79.200 111.630 ;
        RECT 54.230 111.430 79.200 111.510 ;
        RECT 54.260 111.380 79.200 111.430 ;
        RECT 56.610 111.330 79.200 111.380 ;
        RECT 19.770 111.140 23.260 111.150 ;
        RECT 15.030 110.940 15.370 111.000 ;
        RECT 19.470 110.950 23.260 111.140 ;
        RECT 56.410 110.970 56.490 111.150 ;
        RECT 19.470 110.940 19.930 110.950 ;
        RECT -18.390 110.810 -17.490 110.850 ;
        RECT -126.790 107.140 -26.950 107.230 ;
        RECT -126.790 106.260 -25.730 107.140 ;
        RECT -18.390 106.260 -18.020 110.810 ;
        RECT 10.760 110.580 11.220 110.900 ;
        RECT 12.930 110.720 15.370 110.940 ;
        RECT 50.560 110.340 51.160 110.510 ;
        RECT 54.160 110.340 59.390 110.570 ;
        RECT -10.200 110.140 -9.890 110.250 ;
        RECT 41.690 110.160 53.220 110.340 ;
        RECT -16.910 110.120 -9.890 110.140 ;
        RECT -126.790 105.890 -18.020 106.260 ;
        RECT -17.200 109.950 -9.890 110.120 ;
        RECT -17.200 109.770 -15.700 109.950 ;
        RECT -10.200 109.920 -9.890 109.950 ;
        RECT -8.900 110.080 -8.590 110.150 ;
        RECT -6.800 110.080 -6.480 110.110 ;
        RECT -8.900 109.880 -6.380 110.080 ;
        RECT 50.560 109.950 51.160 110.160 ;
        RECT 54.630 110.100 54.940 110.240 ;
        RECT 52.460 110.090 54.940 110.100 ;
        RECT 52.460 109.940 63.980 110.090 ;
        RECT 52.460 109.920 54.940 109.940 ;
        RECT 54.630 109.910 54.940 109.920 ;
        RECT -8.900 109.820 -8.590 109.880 ;
        RECT -6.800 109.850 -6.480 109.880 ;
        RECT -17.200 109.180 -16.540 109.770 ;
        RECT -16.070 109.730 -15.700 109.770 ;
        RECT 31.610 109.750 31.920 109.800 ;
        RECT 31.610 109.740 32.070 109.750 ;
        RECT 31.610 109.560 33.860 109.740 ;
        RECT 31.610 109.470 31.920 109.560 ;
        RECT 54.170 109.520 59.390 109.740 ;
        RECT 50.890 109.320 51.200 109.390 ;
        RECT -10.200 109.180 -9.890 109.290 ;
        RECT -17.200 108.990 -9.890 109.180 ;
        RECT -17.200 108.810 -15.700 108.990 ;
        RECT -10.200 108.960 -9.890 108.990 ;
        RECT -8.900 109.120 -8.590 109.190 ;
        RECT -6.790 109.120 -6.470 109.150 ;
        RECT -8.900 108.920 -6.380 109.120 ;
        RECT 50.890 109.100 53.220 109.320 ;
        RECT -8.900 108.860 -8.590 108.920 ;
        RECT -6.790 108.890 -6.470 108.920 ;
        RECT -17.200 108.800 -16.530 108.810 ;
        RECT -17.200 108.760 -16.540 108.800 ;
        RECT -16.070 108.770 -15.700 108.810 ;
        RECT 10.760 108.760 11.220 109.080 ;
        RECT 50.890 109.060 51.200 109.100 ;
        RECT -126.790 105.260 -25.730 105.890 ;
        RECT -126.790 105.150 -26.950 105.260 ;
        RECT -126.790 61.320 -124.710 105.150 ;
        RECT -127.010 57.910 -124.710 61.320 ;
        RECT -126.790 57.580 -124.710 57.910 ;
        RECT -122.450 102.390 -26.950 102.410 ;
        RECT -122.450 101.500 -25.790 102.390 ;
        RECT -17.200 101.500 -16.830 108.760 ;
        RECT 12.930 108.720 15.370 108.940 ;
        RECT 19.770 108.730 20.070 108.760 ;
        RECT 19.770 108.720 20.160 108.730 ;
        RECT 10.570 108.360 10.660 108.680 ;
        RECT -10.200 108.220 -9.890 108.330 ;
        RECT -122.450 101.130 -16.830 101.500 ;
        RECT -16.070 108.030 -9.890 108.220 ;
        RECT -122.450 100.510 -25.790 101.130 ;
        RECT -122.450 100.330 -26.950 100.510 ;
        RECT -122.450 32.840 -120.370 100.330 ;
        RECT -117.910 97.570 -26.950 97.710 ;
        RECT -117.910 96.660 -25.730 97.570 ;
        RECT -16.070 96.660 -15.700 108.030 ;
        RECT -10.200 108.000 -9.890 108.030 ;
        RECT -8.900 108.160 -8.590 108.230 ;
        RECT -6.800 108.160 -6.480 108.190 ;
        RECT -8.900 107.960 -6.380 108.160 ;
        RECT -8.900 107.900 -8.590 107.960 ;
        RECT -6.800 107.930 -6.480 107.960 ;
        RECT 13.030 107.920 13.290 108.720 ;
        RECT 15.030 108.660 15.370 108.720 ;
        RECT 19.470 108.520 20.160 108.720 ;
        RECT 30.390 108.600 30.870 108.830 ;
        RECT 30.530 108.530 30.870 108.600 ;
        RECT 23.400 108.120 33.860 108.340 ;
        RECT 17.860 108.100 18.180 108.110 ;
        RECT 17.860 107.900 19.490 108.100 ;
        RECT 23.400 107.980 23.720 108.120 ;
        RECT 17.860 107.850 18.180 107.900 ;
        RECT 10.760 107.210 11.220 107.530 ;
        RECT 19.260 107.500 19.370 107.700 ;
        RECT 23.420 107.640 23.680 107.980 ;
        RECT 19.740 107.410 20.070 107.610 ;
        RECT 12.930 107.170 15.370 107.390 ;
        RECT 19.740 107.190 19.920 107.410 ;
        RECT 23.400 107.380 23.720 107.640 ;
        RECT 25.770 107.490 26.500 107.670 ;
        RECT 30.530 107.660 30.870 107.730 ;
        RECT 25.770 107.280 25.950 107.490 ;
        RECT 30.390 107.430 30.870 107.660 ;
        RECT 19.720 107.170 19.920 107.190 ;
        RECT 10.570 106.810 10.660 107.130 ;
        RECT 13.030 106.370 13.290 107.170 ;
        RECT 15.030 107.110 15.370 107.170 ;
        RECT 19.470 106.970 19.920 107.170 ;
        RECT 25.380 107.100 25.950 107.280 ;
        RECT 54.940 107.060 59.390 107.220 ;
        RECT 54.910 107.020 59.390 107.060 ;
        RECT 26.540 106.850 26.860 106.970 ;
        RECT 48.740 106.850 49.060 106.970 ;
        RECT 26.540 106.670 49.060 106.850 ;
        RECT 24.350 106.560 24.660 106.630 ;
        RECT 17.860 106.550 18.180 106.560 ;
        RECT 17.860 106.350 19.490 106.550 ;
        RECT 22.330 106.380 33.860 106.560 ;
        RECT 34.040 106.380 34.360 106.400 ;
        RECT 22.330 106.350 34.360 106.380 ;
        RECT 17.860 106.300 18.180 106.350 ;
        RECT 23.640 106.340 34.360 106.350 ;
        RECT 24.350 106.300 24.660 106.340 ;
        RECT 10.760 105.660 11.220 105.980 ;
        RECT 19.260 105.950 19.370 106.150 ;
        RECT 25.870 106.130 26.050 106.340 ;
        RECT 25.380 105.950 26.050 106.130 ;
        RECT 31.630 106.190 34.360 106.340 ;
        RECT 31.630 106.110 31.950 106.190 ;
        RECT 34.040 106.180 34.360 106.190 ;
        RECT 34.040 106.140 36.060 106.180 ;
        RECT 31.640 106.030 31.950 106.110 ;
        RECT 12.930 105.620 15.370 105.840 ;
        RECT 19.720 105.780 20.070 105.850 ;
        RECT 19.720 105.620 20.110 105.780 ;
        RECT 30.390 105.670 30.870 105.900 ;
        RECT 31.640 105.820 33.860 106.030 ;
        RECT 34.150 106.020 36.060 106.140 ;
        RECT 34.870 106.000 36.060 106.020 ;
        RECT 31.640 105.780 31.950 105.820 ;
        RECT 35.200 105.740 36.040 105.940 ;
        RECT 10.570 105.260 10.660 105.580 ;
        RECT 13.030 104.820 13.290 105.620 ;
        RECT 15.030 105.560 15.370 105.620 ;
        RECT 19.530 105.550 20.110 105.620 ;
        RECT 19.530 105.420 19.920 105.550 ;
        RECT 24.500 105.470 24.810 105.610 ;
        RECT 30.530 105.600 30.870 105.670 ;
        RECT 22.330 105.460 24.810 105.470 ;
        RECT 22.330 105.310 33.860 105.460 ;
        RECT 22.330 105.290 24.810 105.310 ;
        RECT 24.500 105.280 24.810 105.290 ;
        RECT 17.860 105.000 18.180 105.010 ;
        RECT 17.860 104.800 19.490 105.000 ;
        RECT 17.860 104.750 18.180 104.800 ;
        RECT 30.530 104.730 30.870 104.800 ;
        RECT 10.760 104.110 11.220 104.430 ;
        RECT 19.260 104.400 19.370 104.600 ;
        RECT 19.810 104.470 20.070 104.680 ;
        RECT 30.390 104.500 30.870 104.730 ;
        RECT 51.470 104.540 51.780 104.590 ;
        RECT 53.770 104.540 54.080 104.560 ;
        RECT 54.910 104.540 55.140 107.020 ;
        RECT 56.410 106.100 56.490 106.280 ;
        RECT 79.180 104.620 79.490 104.740 ;
        RECT 78.410 104.610 79.530 104.620 ;
        RECT 80.750 104.610 81.060 104.740 ;
        RECT 12.930 104.070 15.370 104.290 ;
        RECT 19.810 104.070 20.010 104.470 ;
        RECT 35.600 104.320 44.610 104.520 ;
        RECT 50.540 104.360 51.160 104.460 ;
        RECT 50.260 104.320 51.160 104.360 ;
        RECT 34.810 104.310 44.610 104.320 ;
        RECT 34.120 104.300 44.610 104.310 ;
        RECT 25.380 104.090 26.150 104.270 ;
        RECT 10.570 103.710 10.660 104.030 ;
        RECT 13.030 103.270 13.290 104.070 ;
        RECT 15.030 104.010 15.370 104.070 ;
        RECT 19.670 103.870 20.010 104.070 ;
        RECT 19.810 103.860 20.010 103.870 ;
        RECT 17.860 103.450 18.180 103.460 ;
        RECT 17.860 103.250 19.490 103.450 ;
        RECT 17.860 103.200 18.180 103.250 ;
        RECT 19.260 102.850 19.370 103.050 ;
        RECT 25.970 101.650 26.150 104.090 ;
        RECT 31.630 104.210 31.950 104.290 ;
        RECT 34.120 104.260 36.060 104.300 ;
        RECT 34.040 104.210 36.060 104.260 ;
        RECT 31.630 104.150 36.060 104.210 ;
        RECT 31.630 104.020 34.360 104.150 ;
        RECT 34.810 104.140 36.060 104.150 ;
        RECT 31.630 103.970 31.950 104.020 ;
        RECT 34.040 104.000 34.360 104.020 ;
        RECT 34.780 103.860 35.100 103.910 ;
        RECT 34.780 103.610 40.800 103.860 ;
        RECT 40.480 103.540 40.800 103.610 ;
        RECT 39.940 103.030 40.250 103.170 ;
        RECT 44.390 103.030 44.610 104.300 ;
        RECT 49.940 104.080 51.160 104.320 ;
        RECT 51.470 104.310 55.140 104.540 ;
        RECT 55.750 104.410 59.390 104.610 ;
        RECT 59.760 104.410 81.060 104.610 ;
        RECT 51.470 104.260 51.780 104.310 ;
        RECT 53.770 104.230 54.080 104.310 ;
        RECT 50.260 104.030 51.160 104.080 ;
        RECT 50.540 103.930 51.160 104.030 ;
        RECT 51.470 103.710 51.780 103.770 ;
        RECT 53.760 103.710 54.070 103.840 ;
        RECT 55.750 103.710 55.950 104.410 ;
        RECT 78.410 104.400 79.530 104.410 ;
        RECT 51.470 103.560 55.950 103.710 ;
        RECT 51.470 103.490 55.920 103.560 ;
        RECT 51.470 103.440 51.780 103.490 ;
        RECT 60.710 103.030 61.020 103.170 ;
        RECT 37.780 102.850 47.850 103.030 ;
        RECT 53.110 102.850 63.180 103.030 ;
        RECT 39.940 102.840 40.250 102.850 ;
        RECT 35.650 102.600 41.310 102.740 ;
        RECT 44.390 102.690 44.610 102.850 ;
        RECT 60.710 102.840 61.020 102.850 ;
        RECT 44.390 102.600 47.240 102.690 ;
        RECT 87.700 102.640 88.600 102.650 ;
        RECT 60.710 102.600 61.020 102.620 ;
        RECT 35.650 102.520 47.850 102.600 ;
        RECT 37.780 102.420 47.850 102.520 ;
        RECT 53.110 102.420 63.180 102.600 ;
        RECT 39.940 102.290 40.250 102.420 ;
        RECT 35.150 102.220 35.630 102.230 ;
        RECT 35.150 101.980 36.040 102.220 ;
        RECT 41.090 102.190 41.310 102.420 ;
        RECT 60.710 102.290 61.020 102.420 ;
        RECT 51.420 102.240 51.730 102.280 ;
        RECT 45.460 102.190 51.730 102.240 ;
        RECT 41.090 102.030 51.730 102.190 ;
        RECT 41.090 101.970 45.850 102.030 ;
        RECT 51.420 101.950 51.730 102.030 ;
        RECT 84.960 101.730 85.740 101.880 ;
        RECT 87.700 101.730 190.930 102.640 ;
        RECT 25.970 101.470 26.510 101.650 ;
        RECT 39.940 101.600 40.250 101.730 ;
        RECT 37.780 101.420 47.860 101.600 ;
        RECT 51.470 101.550 51.780 101.630 ;
        RECT 60.710 101.600 61.020 101.730 ;
        RECT 53.100 101.550 63.180 101.600 ;
        RECT 51.470 101.420 63.180 101.550 ;
        RECT 39.940 101.400 40.250 101.420 ;
        RECT 51.470 101.320 54.180 101.420 ;
        RECT 60.710 101.400 61.020 101.420 ;
        RECT 51.470 101.300 51.780 101.320 ;
        RECT 53.680 101.260 53.990 101.320 ;
        RECT 84.960 101.260 190.930 101.730 ;
        RECT 60.710 101.170 61.020 101.180 ;
        RECT 53.100 100.990 63.180 101.170 ;
        RECT 84.960 101.110 85.740 101.260 ;
        RECT 60.710 100.850 61.020 100.990 ;
        RECT 29.110 100.710 29.430 100.720 ;
        RECT 56.920 100.710 57.380 100.780 ;
        RECT 29.110 100.430 57.380 100.710 ;
        RECT 87.700 100.560 190.930 101.260 ;
        RECT 88.580 100.550 190.930 100.560 ;
        RECT 29.110 100.380 29.430 100.430 ;
        RECT 56.920 100.370 57.380 100.430 ;
        RECT 39.940 100.020 40.250 100.160 ;
        RECT 57.710 100.110 58.140 100.190 ;
        RECT 37.780 100.010 40.250 100.020 ;
        RECT 46.450 100.010 58.140 100.110 ;
        RECT 60.710 100.020 61.020 100.160 ;
        RECT 60.710 100.010 63.180 100.020 ;
        RECT 37.780 99.850 63.180 100.010 ;
        RECT 37.780 99.840 47.840 99.850 ;
        RECT 53.120 99.840 63.180 99.850 ;
        RECT 39.940 99.830 40.250 99.840 ;
        RECT 57.710 99.780 58.140 99.840 ;
        RECT 60.710 99.830 61.020 99.840 ;
        RECT 31.630 99.240 31.950 99.290 ;
        RECT 34.040 99.240 34.360 99.260 ;
        RECT 26.140 99.050 27.920 99.170 ;
        RECT 25.550 98.990 27.920 99.050 ;
        RECT 31.630 99.100 34.360 99.240 ;
        RECT 31.630 99.050 36.060 99.100 ;
        RECT 10.760 98.630 11.220 98.950 ;
        RECT 25.550 98.870 26.390 98.990 ;
        RECT 31.630 98.970 31.950 99.050 ;
        RECT 34.040 99.000 36.060 99.050 ;
        RECT 40.420 99.030 40.560 99.220 ;
        RECT 60.450 99.030 60.540 99.210 ;
        RECT 34.080 98.930 36.060 99.000 ;
        RECT 35.540 98.920 36.060 98.930 ;
        RECT 12.930 98.590 15.370 98.810 ;
        RECT 19.810 98.690 20.060 98.710 ;
        RECT 19.810 98.590 20.070 98.690 ;
        RECT 10.570 98.230 10.660 98.550 ;
        RECT 13.030 97.790 13.290 98.590 ;
        RECT 15.030 98.530 15.370 98.590 ;
        RECT 19.470 98.390 20.070 98.590 ;
        RECT 30.390 98.530 30.870 98.760 ;
        RECT 39.940 98.610 40.250 98.730 ;
        RECT 40.420 98.610 40.560 98.790 ;
        RECT 47.680 98.610 48.240 98.740 ;
        RECT 60.450 98.610 60.540 98.780 ;
        RECT 60.710 98.610 61.020 98.730 ;
        RECT 39.940 98.600 48.240 98.610 ;
        RECT 30.530 98.460 30.870 98.530 ;
        RECT 37.780 98.560 48.240 98.600 ;
        RECT 53.120 98.600 61.020 98.610 ;
        RECT 37.780 98.440 47.840 98.560 ;
        RECT 53.120 98.440 63.180 98.600 ;
        RECT 37.780 98.420 40.340 98.440 ;
        RECT 39.940 98.400 40.250 98.420 ;
        RECT 45.520 98.350 47.060 98.440 ;
        RECT 53.900 98.350 55.440 98.440 ;
        RECT 60.620 98.420 63.180 98.440 ;
        RECT 60.710 98.400 61.020 98.420 ;
        RECT 39.940 98.170 40.250 98.180 ;
        RECT 60.710 98.170 61.020 98.180 ;
        RECT 37.780 98.000 47.840 98.170 ;
        RECT 53.120 98.000 63.180 98.170 ;
        RECT 37.780 97.990 40.250 98.000 ;
        RECT 17.860 97.970 18.180 97.980 ;
        RECT 17.860 97.770 19.490 97.970 ;
        RECT 39.940 97.850 40.250 97.990 ;
        RECT 60.710 97.990 63.180 98.000 ;
        RECT 17.860 97.720 18.180 97.770 ;
        RECT 30.530 97.590 30.870 97.660 ;
        RECT 40.420 97.600 40.570 97.790 ;
        RECT 58.450 97.740 58.890 97.860 ;
        RECT 60.710 97.850 61.020 97.990 ;
        RECT 10.760 97.080 11.220 97.400 ;
        RECT 19.260 97.370 19.370 97.570 ;
        RECT 19.660 97.340 20.040 97.540 ;
        RECT 30.390 97.360 30.870 97.590 ;
        RECT 47.690 97.560 58.890 97.740 ;
        RECT 60.420 97.600 60.550 97.780 ;
        RECT 58.450 97.460 58.890 97.560 ;
        RECT 19.660 97.310 20.030 97.340 ;
        RECT 12.930 97.040 15.370 97.260 ;
        RECT 19.660 97.040 19.860 97.310 ;
        RECT 26.160 97.210 27.920 97.310 ;
        RECT 10.570 96.680 10.660 97.000 ;
        RECT -117.910 96.290 -15.700 96.660 ;
        RECT -117.910 95.690 -25.730 96.290 ;
        RECT 13.030 96.240 13.290 97.040 ;
        RECT 15.030 96.980 15.370 97.040 ;
        RECT 19.470 96.840 19.860 97.040 ;
        RECT 25.560 97.130 27.920 97.210 ;
        RECT 25.560 97.030 26.440 97.130 ;
        RECT 31.630 97.070 31.950 97.150 ;
        RECT 34.110 97.120 36.060 97.260 ;
        RECT 40.420 97.170 40.550 97.350 ;
        RECT 60.410 97.170 60.550 97.350 ;
        RECT 34.040 97.100 36.060 97.120 ;
        RECT 34.040 97.070 34.360 97.100 ;
        RECT 34.840 97.090 36.060 97.100 ;
        RECT 35.540 97.080 36.060 97.090 ;
        RECT 31.630 96.880 34.360 97.070 ;
        RECT 31.630 96.830 31.950 96.880 ;
        RECT 34.040 96.860 34.360 96.880 ;
        RECT 17.860 96.420 18.180 96.430 ;
        RECT 17.860 96.220 19.490 96.420 ;
        RECT 31.630 96.310 31.950 96.360 ;
        RECT 34.040 96.310 34.360 96.330 ;
        RECT 17.860 96.170 18.180 96.220 ;
        RECT 26.170 96.060 27.920 96.160 ;
        RECT -117.910 95.630 -26.950 95.690 ;
        RECT -122.660 29.240 -120.090 32.840 ;
        RECT -122.450 29.200 -120.370 29.240 ;
        RECT -117.910 4.220 -115.830 95.630 ;
        RECT 10.760 95.530 11.220 95.850 ;
        RECT 19.260 95.820 19.370 96.020 ;
        RECT 25.560 95.980 27.920 96.060 ;
        RECT 31.630 96.120 34.360 96.310 ;
        RECT 31.630 96.040 31.950 96.120 ;
        RECT 34.040 96.110 34.360 96.120 ;
        RECT 34.040 96.070 36.060 96.110 ;
        RECT 25.560 95.880 26.440 95.980 ;
        RECT 34.150 95.950 36.060 96.070 ;
        RECT 40.420 96.020 40.490 96.200 ;
        RECT 60.460 96.020 60.550 96.200 ;
        RECT 34.870 95.930 36.060 95.950 ;
        RECT 12.930 95.490 15.370 95.710 ;
        RECT 19.870 95.490 20.070 95.770 ;
        RECT 30.390 95.600 30.870 95.830 ;
        RECT 30.530 95.530 30.870 95.600 ;
        RECT 40.420 95.590 40.490 95.770 ;
        RECT 60.460 95.590 60.550 95.770 ;
        RECT 10.570 95.130 10.660 95.450 ;
        RECT 13.030 94.690 13.290 95.490 ;
        RECT 15.030 95.430 15.370 95.490 ;
        RECT 19.470 95.290 20.070 95.490 ;
        RECT 47.120 95.040 53.880 95.220 ;
        RECT 17.860 94.870 18.180 94.880 ;
        RECT 17.860 94.670 19.490 94.870 ;
        RECT 17.860 94.620 18.180 94.670 ;
        RECT 30.530 94.660 30.870 94.730 ;
        RECT 10.760 93.980 11.220 94.300 ;
        RECT 19.260 94.270 19.370 94.470 ;
        RECT 12.930 93.940 15.370 94.160 ;
        RECT 19.870 93.940 20.070 94.610 ;
        RECT 30.390 94.430 30.870 94.660 ;
        RECT 40.420 94.600 40.490 94.780 ;
        RECT 60.460 94.600 60.550 94.780 ;
        RECT 26.140 94.200 27.920 94.310 ;
        RECT 34.810 94.240 36.060 94.250 ;
        RECT 25.560 94.130 27.920 94.200 ;
        RECT 31.630 94.140 31.950 94.220 ;
        RECT 34.120 94.190 36.060 94.240 ;
        RECT 34.040 94.140 36.060 94.190 ;
        RECT 40.420 94.170 40.490 94.350 ;
        RECT 60.460 94.170 60.550 94.350 ;
        RECT 25.560 94.020 26.440 94.130 ;
        RECT 31.630 94.080 36.060 94.140 ;
        RECT 10.570 93.580 10.660 93.900 ;
        RECT -113.560 93.350 -26.950 93.450 ;
        RECT -113.560 92.510 -25.790 93.350 ;
        RECT 13.030 93.140 13.290 93.940 ;
        RECT 15.030 93.880 15.370 93.940 ;
        RECT 19.470 93.740 20.070 93.940 ;
        RECT 31.630 93.950 34.360 94.080 ;
        RECT 34.810 94.070 36.060 94.080 ;
        RECT 31.630 93.900 31.950 93.950 ;
        RECT 34.040 93.930 34.360 93.950 ;
        RECT 17.860 93.320 18.180 93.330 ;
        RECT 17.860 93.120 19.490 93.320 ;
        RECT 27.240 93.210 27.550 93.350 ;
        RECT 17.860 93.070 18.180 93.120 ;
        RECT 25.080 93.030 27.650 93.210 ;
        RECT 27.240 93.020 27.550 93.030 ;
        RECT 19.260 92.720 19.370 92.920 ;
        RECT -113.560 92.140 -17.360 92.510 ;
        RECT -113.560 91.470 -25.790 92.140 ;
        RECT -113.560 91.370 -26.950 91.470 ;
        RECT -118.070 0.650 -115.680 4.220 ;
        RECT -117.910 0.120 -115.830 0.650 ;
        RECT -113.560 -24.390 -111.480 91.370 ;
        RECT -17.730 90.790 -17.360 92.140 ;
        RECT -17.730 90.780 -15.700 90.790 ;
        RECT -17.730 90.600 -15.480 90.780 ;
        RECT -17.730 90.540 -14.080 90.600 ;
        RECT -11.080 90.540 -10.770 90.580 ;
        RECT -17.730 90.420 -10.770 90.540 ;
        RECT -16.070 90.380 -10.770 90.420 ;
        RECT -15.700 90.320 -10.770 90.380 ;
        RECT -23.070 90.130 -22.300 90.320 ;
        RECT -11.080 90.250 -10.770 90.320 ;
        RECT 27.240 90.200 27.550 90.340 ;
        RECT 25.070 90.190 27.550 90.200 ;
        RECT -16.070 90.130 -15.680 90.150 ;
        RECT -23.070 90.090 -15.680 90.130 ;
        RECT -12.300 90.090 -11.990 90.140 ;
        RECT -23.070 89.880 -11.990 90.090 ;
        RECT 25.070 90.020 27.670 90.190 ;
        RECT 27.240 90.010 27.550 90.020 ;
        RECT -23.070 89.760 -15.690 89.880 ;
        RECT -12.300 89.810 -11.990 89.880 ;
        RECT -23.070 89.580 -22.300 89.760 ;
        RECT -16.070 89.740 -15.700 89.760 ;
        RECT -109.220 89.250 -26.950 89.380 ;
        RECT -109.220 88.480 -25.730 89.250 ;
        RECT 25.410 89.210 27.740 89.390 ;
        RECT 28.270 89.180 28.590 89.240 ;
        RECT 32.290 89.180 32.620 89.210 ;
        RECT 10.760 88.860 11.220 89.180 ;
        RECT 12.930 88.820 15.370 89.040 ;
        RECT 28.270 89.010 32.620 89.180 ;
        RECT 28.270 88.960 28.590 89.010 ;
        RECT 32.290 88.950 32.620 89.010 ;
        RECT -109.220 88.110 -21.010 88.480 ;
        RECT 10.570 88.460 10.660 88.780 ;
        RECT -109.220 87.370 -25.730 88.110 ;
        RECT -109.220 87.300 -26.950 87.370 ;
        RECT -113.740 -27.910 -111.290 -24.390 ;
        RECT -113.560 -28.030 -111.480 -27.910 ;
        RECT -109.220 -52.900 -107.140 87.300 ;
        RECT -21.380 86.450 -21.010 88.110 ;
        RECT 13.030 88.020 13.290 88.820 ;
        RECT 15.030 88.760 15.370 88.820 ;
        RECT 19.450 88.620 20.100 88.820 ;
        RECT 17.860 88.200 18.180 88.210 ;
        RECT 17.860 88.000 19.490 88.200 ;
        RECT 17.860 87.950 18.180 88.000 ;
        RECT 10.760 87.310 11.220 87.630 ;
        RECT 19.260 87.600 19.370 87.800 ;
        RECT 19.830 87.570 20.080 87.800 ;
        RECT 12.930 87.270 15.370 87.490 ;
        RECT 19.830 87.270 20.030 87.570 ;
        RECT 10.570 86.910 10.660 87.230 ;
        RECT 13.030 86.470 13.290 87.270 ;
        RECT 15.030 87.210 15.370 87.270 ;
        RECT 19.470 87.070 20.030 87.270 ;
        RECT 25.410 87.350 27.750 87.530 ;
        RECT 25.410 87.250 25.590 87.350 ;
        RECT 17.860 86.650 18.180 86.660 ;
        RECT 17.860 86.450 19.490 86.650 ;
        RECT -21.380 86.270 -15.430 86.450 ;
        RECT 17.860 86.400 18.180 86.450 ;
        RECT -21.380 86.200 -15.360 86.270 ;
        RECT -13.970 86.200 -12.700 86.210 ;
        RECT -12.270 86.200 -11.960 86.260 ;
        RECT -21.380 86.080 -11.960 86.200 ;
        RECT -16.070 86.040 -11.960 86.080 ;
        RECT -15.710 85.990 -11.960 86.040 ;
        RECT -12.270 85.930 -11.960 85.990 ;
        RECT -11.580 86.180 -11.270 86.250 ;
        RECT -6.790 86.200 -6.500 86.220 ;
        RECT -11.580 86.170 -9.440 86.180 ;
        RECT -6.800 86.170 -6.480 86.200 ;
        RECT -11.580 85.970 -6.480 86.170 ;
        RECT -11.580 85.920 -11.270 85.970 ;
        RECT -9.650 85.960 -6.480 85.970 ;
        RECT -17.840 85.470 -17.430 85.490 ;
        RECT -16.070 85.470 -14.080 85.490 ;
        RECT -17.840 85.430 -14.080 85.470 ;
        RECT -11.100 85.430 -10.790 85.480 ;
        RECT -105.060 85.160 -26.950 85.230 ;
        RECT -17.840 85.210 -10.790 85.430 ;
        RECT -105.060 84.340 -25.730 85.160 ;
        RECT -17.840 85.100 -15.690 85.210 ;
        RECT -11.100 85.150 -10.790 85.210 ;
        RECT -10.390 85.350 -10.080 85.420 ;
        RECT -9.650 85.350 -9.440 85.960 ;
        RECT -6.800 85.940 -6.480 85.960 ;
        RECT -6.790 85.920 -6.500 85.940 ;
        RECT 10.760 85.760 11.220 86.080 ;
        RECT 19.260 86.050 19.370 86.250 ;
        RECT 25.420 86.200 27.740 86.380 ;
        RECT 27.190 86.190 27.350 86.200 ;
        RECT 19.840 86.010 20.040 86.020 ;
        RECT 12.930 85.720 15.370 85.940 ;
        RECT 19.840 85.740 20.130 86.010 ;
        RECT 19.840 85.720 20.040 85.740 ;
        RECT 10.570 85.360 10.660 85.680 ;
        RECT -10.390 85.140 -9.440 85.350 ;
        RECT -17.840 85.080 -17.430 85.100 ;
        RECT -16.070 85.080 -15.700 85.100 ;
        RECT -10.390 85.090 -10.080 85.140 ;
        RECT 13.030 84.920 13.290 85.720 ;
        RECT 15.030 85.660 15.370 85.720 ;
        RECT 19.430 85.520 20.040 85.720 ;
        RECT 40.860 85.430 41.190 85.520 ;
        RECT 34.510 85.260 41.190 85.430 ;
        RECT 40.860 85.230 41.190 85.260 ;
        RECT 17.860 85.100 18.180 85.110 ;
        RECT 17.860 84.900 19.490 85.100 ;
        RECT 17.860 84.850 18.180 84.900 ;
        RECT 19.820 84.860 20.120 84.900 ;
        RECT -23.070 84.340 -22.270 84.480 ;
        RECT -105.060 83.840 -22.270 84.340 ;
        RECT -10.430 84.270 -9.820 84.600 ;
        RECT -105.060 83.280 -25.730 83.840 ;
        RECT -23.070 83.710 -22.270 83.840 ;
        RECT -10.420 83.780 -9.820 84.270 ;
        RECT 10.760 84.210 11.220 84.530 ;
        RECT 19.260 84.500 19.370 84.700 ;
        RECT 19.810 84.620 20.120 84.860 ;
        RECT 27.140 84.710 27.450 85.040 ;
        RECT 30.530 84.900 30.870 84.970 ;
        RECT 30.390 84.670 30.870 84.900 ;
        RECT 12.930 84.170 15.370 84.390 ;
        RECT 19.810 84.170 20.010 84.620 ;
        RECT 27.210 84.530 27.370 84.540 ;
        RECT 25.420 84.350 27.740 84.530 ;
        RECT 34.810 84.480 36.060 84.490 ;
        RECT 31.630 84.380 31.950 84.460 ;
        RECT 34.120 84.430 36.060 84.480 ;
        RECT 34.040 84.380 36.060 84.430 ;
        RECT 31.630 84.350 36.060 84.380 ;
        RECT 38.580 84.360 38.890 84.420 ;
        RECT 38.030 84.350 38.890 84.360 ;
        RECT 10.570 83.810 10.660 84.130 ;
        RECT 13.030 83.370 13.290 84.170 ;
        RECT 15.030 84.110 15.370 84.170 ;
        RECT 19.460 83.970 20.010 84.170 ;
        RECT 27.190 84.070 27.500 84.190 ;
        RECT 30.450 84.130 38.890 84.350 ;
        RECT 30.450 84.120 38.040 84.130 ;
        RECT 30.450 84.110 31.220 84.120 ;
        RECT 30.450 84.070 30.690 84.110 ;
        RECT 38.580 84.090 38.890 84.130 ;
        RECT 27.190 83.870 30.690 84.070 ;
        RECT 27.190 83.860 29.880 83.870 ;
        RECT 27.190 83.580 27.510 83.670 ;
        RECT 37.810 83.580 38.220 83.690 ;
        RECT 17.860 83.550 18.180 83.560 ;
        RECT 17.860 83.350 19.490 83.550 ;
        RECT 27.190 83.420 38.220 83.580 ;
        RECT 27.190 83.390 27.510 83.420 ;
        RECT 17.860 83.300 18.180 83.350 ;
        RECT 37.810 83.320 38.220 83.420 ;
        RECT -105.060 83.150 -26.950 83.280 ;
        RECT -109.470 -56.630 -106.870 -52.900 ;
        RECT -109.220 -56.960 -107.140 -56.630 ;
        RECT -105.060 -81.530 -102.980 83.150 ;
        RECT 43.850 82.120 44.150 82.140 ;
        RECT 37.510 81.540 38.170 81.900 ;
        RECT 43.140 81.780 44.160 82.120 ;
        RECT 43.850 81.760 44.160 81.780 ;
        RECT 39.260 80.820 39.710 81.250 ;
        RECT -100.810 80.010 -26.950 80.080 ;
        RECT -100.810 79.230 -25.790 80.010 ;
        RECT -17.830 79.230 -17.420 79.250 ;
        RECT -100.810 78.860 -17.420 79.230 ;
        RECT -100.810 78.130 -25.790 78.860 ;
        RECT -17.830 78.840 -17.420 78.860 ;
        RECT -100.810 78.000 -26.950 78.130 ;
        RECT -105.480 -85.200 -102.770 -81.530 ;
        RECT -105.060 -85.920 -102.980 -85.200 ;
        RECT -100.810 -110.150 -98.730 78.000 ;
        RECT 88.010 77.040 88.020 77.050 ;
        RECT -10.390 76.710 -9.780 77.040 ;
        RECT -10.380 76.220 -9.780 76.710 ;
        RECT -16.110 75.840 -15.740 75.850 ;
        RECT -96.550 75.720 -26.950 75.820 ;
        RECT -96.550 75.020 -25.730 75.720 ;
        RECT -17.430 75.460 -14.900 75.840 ;
        RECT -17.430 75.020 -17.050 75.460 ;
        RECT -16.110 75.440 -15.740 75.460 ;
        RECT -96.550 74.640 -17.050 75.020 ;
        RECT -96.550 73.840 -25.730 74.640 ;
        RECT -96.550 73.740 -26.950 73.840 ;
        RECT -101.140 -113.630 -98.400 -110.150 ;
        RECT -100.810 -114.440 -98.730 -113.630 ;
        RECT -96.550 -138.440 -94.470 73.740 ;
        RECT 18.340 72.640 18.940 73.130 ;
        RECT 18.340 72.310 18.950 72.640 ;
        RECT -92.400 70.700 -26.950 70.780 ;
        RECT -92.400 69.790 -25.730 70.700 ;
        RECT -92.400 69.410 -17.030 69.790 ;
        RECT 74.900 69.740 75.190 69.800 ;
        RECT 74.730 69.430 75.190 69.740 ;
        RECT -92.400 68.820 -25.730 69.410 ;
        RECT -92.400 68.700 -26.950 68.820 ;
        RECT -96.770 -142.490 -93.980 -138.440 ;
        RECT -96.550 -142.770 -94.470 -142.490 ;
        RECT -92.400 -167.220 -90.320 68.700 ;
        RECT -17.410 68.560 -17.030 69.410 ;
        RECT 74.900 69.390 75.190 69.430 ;
        RECT 74.910 69.070 75.190 69.390 ;
        RECT 74.730 68.760 75.190 69.070 ;
        RECT 74.910 68.640 75.190 68.760 ;
        RECT -16.110 68.560 -15.740 68.570 ;
        RECT -17.410 68.180 -14.690 68.560 ;
        RECT -16.110 68.160 -15.740 68.180 ;
        RECT -6.860 67.590 -6.550 67.610 ;
        RECT -11.090 67.250 -6.550 67.590 ;
        RECT -6.860 67.230 -6.550 67.250 ;
        RECT -88.050 65.160 -26.950 65.170 ;
        RECT -88.050 63.280 -25.860 65.160 ;
        RECT -88.050 63.090 -26.950 63.280 ;
        RECT -92.890 -171.000 -90.060 -167.220 ;
        RECT -92.400 -171.560 -90.320 -171.000 ;
        RECT -88.050 -195.800 -85.970 63.090 ;
        RECT 188.840 60.710 190.930 100.550 ;
        RECT -83.890 60.410 -26.950 60.470 ;
        RECT -83.890 58.530 -25.790 60.410 ;
        RECT -83.890 58.390 -26.950 58.530 ;
        RECT -88.400 -199.520 -85.750 -195.800 ;
        RECT -88.050 -199.530 -85.970 -199.520 ;
        RECT -83.890 -224.500 -81.810 58.390 ;
        RECT -84.080 -228.030 -81.410 -224.500 ;
        RECT -22.350 -233.860 -19.010 58.530 ;
        RECT 188.600 57.140 191.110 60.710 ;
        RECT 71.640 56.200 71.960 56.520 ;
      LAYER via2 ;
        RECT 50.690 110.060 51.030 110.400 ;
        RECT 50.710 104.010 51.050 104.370 ;
  END
END sky130_hilas_TopProtectStructure

MACRO sky130_hilas_nFETLarge
  CLASS CORE ;
  FOREIGN sky130_hilas_nFETLarge ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.370 BY 5.830 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    USE ANALOG ;
    ANTENNAGATEAREA 6.396000 ;
    PORT
      LAYER met2 ;
        RECT 0.000 0.330 0.600 0.820 ;
        RECT 0.000 0.000 0.610 0.330 ;
    END
  END GATE
  PIN SOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 4.231200 ;
    PORT
      LAYER met2 ;
        RECT 0.330 5.590 3.390 5.600 ;
        RECT 0.240 5.260 3.390 5.590 ;
        RECT 0.240 2.810 0.560 5.260 ;
        RECT 3.060 5.250 3.370 5.260 ;
        RECT 0.240 2.480 3.400 2.810 ;
        RECT 0.240 1.440 0.560 2.480 ;
        RECT 0.240 1.120 3.400 1.440 ;
        RECT 0.860 1.110 1.170 1.120 ;
        RECT 1.960 1.110 2.270 1.120 ;
        RECT 3.060 1.110 3.370 1.120 ;
    END
  END SOURCE
  PIN DRAIN
    USE ANALOG ;
    ANTENNADIFFAREA 4.231200 ;
    PORT
      LAYER met2 ;
        RECT 1.420 4.880 1.730 4.910 ;
        RECT 2.510 4.880 2.820 4.890 ;
        RECT 1.420 4.580 4.370 4.880 ;
        RECT 2.510 4.560 2.820 4.580 ;
        RECT 3.620 4.540 4.370 4.580 ;
        RECT 3.990 4.410 4.370 4.540 ;
        RECT 4.020 3.540 4.370 4.410 ;
        RECT 1.420 3.210 4.370 3.540 ;
        RECT 4.020 0.770 4.370 3.210 ;
        RECT 1.430 0.760 4.370 0.770 ;
        RECT 1.420 0.450 4.370 0.760 ;
        RECT 1.420 0.440 4.140 0.450 ;
        RECT 1.420 0.430 1.730 0.440 ;
        RECT 2.510 0.430 2.820 0.440 ;
    END
  END DRAIN
  PIN VGND
    ANTENNADIFFAREA 1.444000 ;
    PORT
      LAYER met1 ;
        RECT 0.180 1.920 0.460 2.450 ;
        RECT 0.000 1.620 0.460 1.920 ;
        RECT 0.000 1.600 0.470 1.620 ;
        RECT 0.180 1.170 0.470 1.600 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.950 5.550 1.120 5.580 ;
        RECT 0.880 5.510 1.200 5.550 ;
        RECT 0.880 5.320 1.210 5.510 ;
        RECT 0.880 5.290 1.200 5.320 ;
        RECT 0.950 2.770 1.120 5.290 ;
        RECT 1.500 4.870 1.670 5.580 ;
        RECT 2.050 5.550 2.220 5.580 ;
        RECT 1.970 5.510 2.290 5.550 ;
        RECT 1.970 5.320 2.300 5.510 ;
        RECT 1.970 5.290 2.290 5.320 ;
        RECT 1.430 4.830 1.750 4.870 ;
        RECT 1.430 4.640 1.760 4.830 ;
        RECT 1.430 4.610 1.750 4.640 ;
        RECT 1.500 3.500 1.670 4.610 ;
        RECT 1.430 3.460 1.750 3.500 ;
        RECT 1.430 3.270 1.760 3.460 ;
        RECT 1.430 3.240 1.750 3.270 ;
        RECT 0.870 2.730 1.190 2.770 ;
        RECT 0.870 2.540 1.200 2.730 ;
        RECT 0.870 2.510 1.190 2.540 ;
        RECT 0.240 1.200 0.410 2.390 ;
        RECT 0.950 1.400 1.120 2.510 ;
        RECT 0.870 1.360 1.190 1.400 ;
        RECT 0.870 1.170 1.200 1.360 ;
        RECT 0.870 1.140 1.190 1.170 ;
        RECT 0.190 0.750 0.700 1.010 ;
        RECT 0.190 0.680 0.710 0.750 ;
        RECT 0.200 0.000 0.710 0.680 ;
        RECT 0.950 0.400 1.120 1.140 ;
        RECT 1.500 0.720 1.670 3.240 ;
        RECT 2.050 2.770 2.220 5.290 ;
        RECT 2.600 4.850 2.770 5.580 ;
        RECT 3.150 5.540 3.320 5.580 ;
        RECT 3.070 5.500 3.390 5.540 ;
        RECT 3.070 5.310 3.400 5.500 ;
        RECT 3.070 5.280 3.390 5.310 ;
        RECT 2.520 4.810 2.840 4.850 ;
        RECT 2.520 4.620 2.850 4.810 ;
        RECT 2.520 4.590 2.840 4.620 ;
        RECT 2.600 3.500 2.770 4.590 ;
        RECT 2.520 3.460 2.840 3.500 ;
        RECT 2.520 3.270 2.850 3.460 ;
        RECT 2.520 3.240 2.840 3.270 ;
        RECT 1.970 2.730 2.290 2.770 ;
        RECT 1.970 2.540 2.300 2.730 ;
        RECT 1.970 2.510 2.290 2.540 ;
        RECT 2.050 1.400 2.220 2.510 ;
        RECT 1.970 1.360 2.290 1.400 ;
        RECT 1.970 1.170 2.300 1.360 ;
        RECT 1.970 1.140 2.290 1.170 ;
        RECT 1.430 0.680 1.750 0.720 ;
        RECT 1.430 0.490 1.760 0.680 ;
        RECT 1.430 0.460 1.750 0.490 ;
        RECT 1.500 0.400 1.670 0.460 ;
        RECT 2.050 0.400 2.220 1.140 ;
        RECT 2.600 0.720 2.770 3.240 ;
        RECT 3.150 2.770 3.320 5.280 ;
        RECT 3.700 4.840 3.870 5.580 ;
        RECT 3.630 4.800 3.950 4.840 ;
        RECT 3.630 4.610 3.960 4.800 ;
        RECT 3.630 4.580 3.950 4.610 ;
        RECT 3.700 3.500 3.870 4.580 ;
        RECT 3.620 3.460 3.940 3.500 ;
        RECT 3.620 3.270 3.950 3.460 ;
        RECT 3.620 3.240 3.940 3.270 ;
        RECT 3.070 2.730 3.390 2.770 ;
        RECT 3.070 2.540 3.400 2.730 ;
        RECT 3.070 2.510 3.390 2.540 ;
        RECT 3.150 1.400 3.320 2.510 ;
        RECT 3.070 1.360 3.390 1.400 ;
        RECT 3.070 1.170 3.400 1.360 ;
        RECT 3.070 1.140 3.390 1.170 ;
        RECT 2.520 0.680 2.840 0.720 ;
        RECT 2.520 0.490 2.850 0.680 ;
        RECT 2.520 0.460 2.840 0.490 ;
        RECT 2.600 0.400 2.770 0.460 ;
        RECT 3.150 0.400 3.320 1.140 ;
        RECT 3.700 0.730 3.870 3.240 ;
        RECT 3.620 0.690 3.940 0.730 ;
        RECT 3.620 0.500 3.950 0.690 ;
        RECT 3.620 0.470 3.940 0.500 ;
        RECT 3.700 0.400 3.870 0.470 ;
      LAYER mcon ;
        RECT 0.940 5.330 1.110 5.500 ;
        RECT 2.030 5.330 2.200 5.500 ;
        RECT 1.490 4.650 1.660 4.820 ;
        RECT 1.490 3.280 1.660 3.450 ;
        RECT 0.930 2.550 1.100 2.720 ;
        RECT 0.240 2.220 0.410 2.390 ;
        RECT 0.240 1.880 0.410 2.050 ;
        RECT 0.240 1.540 0.410 1.710 ;
        RECT 0.930 1.180 1.100 1.350 ;
        RECT 0.360 0.540 0.530 0.710 ;
        RECT 3.130 5.320 3.300 5.490 ;
        RECT 2.580 4.630 2.750 4.800 ;
        RECT 2.580 3.280 2.750 3.450 ;
        RECT 2.030 2.550 2.200 2.720 ;
        RECT 2.030 1.180 2.200 1.350 ;
        RECT 1.490 0.500 1.660 0.670 ;
        RECT 3.690 4.620 3.860 4.790 ;
        RECT 3.680 3.280 3.850 3.450 ;
        RECT 3.130 2.550 3.300 2.720 ;
        RECT 3.130 1.180 3.300 1.350 ;
        RECT 2.580 0.500 2.750 0.670 ;
        RECT 3.680 0.510 3.850 0.680 ;
        RECT 0.370 0.070 0.540 0.240 ;
      LAYER met1 ;
        RECT 0.870 5.260 1.190 5.580 ;
        RECT 1.960 5.260 2.280 5.580 ;
        RECT 3.060 5.250 3.380 5.570 ;
        RECT 1.420 4.580 1.740 4.900 ;
        RECT 2.510 4.560 2.830 4.880 ;
        RECT 3.620 4.550 3.940 4.870 ;
        RECT 1.420 3.210 1.740 3.530 ;
        RECT 2.510 3.210 2.830 3.530 ;
        RECT 3.610 3.210 3.930 3.530 ;
        RECT 0.860 2.480 1.180 2.800 ;
        RECT 1.960 2.480 2.280 2.800 ;
        RECT 3.060 2.480 3.380 2.800 ;
        RECT 0.860 1.110 1.180 1.430 ;
        RECT 1.960 1.110 2.280 1.430 ;
        RECT 3.060 1.110 3.380 1.430 ;
        RECT 0.290 0.470 0.610 0.790 ;
        RECT 1.420 0.430 1.740 0.750 ;
        RECT 2.510 0.430 2.830 0.750 ;
        RECT 3.610 0.440 3.930 0.760 ;
        RECT 0.300 0.000 0.620 0.320 ;
      LAYER via ;
        RECT 0.900 5.290 1.160 5.550 ;
        RECT 1.990 5.290 2.250 5.550 ;
        RECT 3.090 5.280 3.350 5.540 ;
        RECT 1.450 4.610 1.710 4.870 ;
        RECT 2.540 4.590 2.800 4.850 ;
        RECT 3.650 4.580 3.910 4.840 ;
        RECT 1.450 3.240 1.710 3.500 ;
        RECT 2.540 3.240 2.800 3.500 ;
        RECT 3.640 3.240 3.900 3.500 ;
        RECT 0.890 2.510 1.150 2.770 ;
        RECT 1.990 2.510 2.250 2.770 ;
        RECT 3.090 2.510 3.350 2.770 ;
        RECT 0.890 1.140 1.150 1.400 ;
        RECT 1.990 1.140 2.250 1.400 ;
        RECT 3.090 1.140 3.350 1.400 ;
        RECT 0.320 0.500 0.580 0.760 ;
        RECT 1.450 0.460 1.710 0.720 ;
        RECT 2.540 0.460 2.800 0.720 ;
        RECT 3.640 0.470 3.900 0.730 ;
        RECT 0.330 0.030 0.590 0.290 ;
  END
END sky130_hilas_nFETLarge

END LIBRARY