magic
tech sky130A
timestamp 1629137261
<< checkpaint >>
rect -587 1861 1397 2123
rect -587 -145 1756 1861
rect -587 -200 1553 -145
rect -256 -630 1553 -200
<< error_s >>
rect 783 832 784 833
<< nwell >>
rect 0 1048 191 1049
rect 0 488 560 1048
rect 760 1031 888 1049
rect 0 470 43 488
rect 0 447 71 470
rect 0 445 43 447
rect 760 444 888 463
<< nsubdiff >>
rect 19 965 50 1002
rect 19 948 25 965
rect 42 948 50 965
rect 19 931 50 948
rect 19 914 25 931
rect 42 914 50 931
rect 19 897 50 914
rect 19 880 25 897
rect 42 880 50 897
rect 19 863 50 880
rect 19 846 25 863
rect 42 846 50 863
rect 19 829 50 846
rect 19 812 25 829
rect 42 812 50 829
rect 19 797 50 812
rect 18 662 50 695
rect 18 645 26 662
rect 43 645 50 662
rect 18 628 50 645
rect 18 611 26 628
rect 43 611 50 628
rect 18 594 50 611
rect 18 577 26 594
rect 43 577 50 594
rect 18 560 50 577
rect 18 543 26 560
rect 43 543 50 560
rect 18 526 50 543
rect 18 509 26 526
rect 43 509 50 526
rect 18 494 50 509
<< nsubdiffcont >>
rect 25 948 42 965
rect 25 914 42 931
rect 25 880 42 897
rect 25 846 42 863
rect 25 812 42 829
rect 26 645 43 662
rect 26 611 43 628
rect 26 577 43 594
rect 26 543 43 560
rect 26 509 43 526
<< locali >>
rect 67 1001 101 1002
rect 42 977 101 1001
rect 42 928 84 977
rect 765 902 767 919
rect 784 902 790 919
rect 765 865 790 902
rect 765 849 786 865
rect 765 832 767 849
rect 784 832 786 849
rect 765 830 786 832
rect 25 795 42 812
rect 26 501 43 509
<< viali >>
rect 25 965 42 982
rect 25 931 42 948
rect 84 960 101 977
rect 84 926 101 943
rect 25 897 42 914
rect 25 863 42 880
rect 25 829 42 846
rect 767 902 784 919
rect 767 832 784 849
rect 26 662 43 679
rect 26 628 43 645
rect 26 594 43 611
rect 26 560 43 577
rect 26 526 43 543
<< metal1 >>
rect 692 1035 726 1049
rect 759 1034 786 1049
rect 22 1002 75 1003
rect 22 1001 101 1002
rect 22 995 104 1001
rect 22 982 34 995
rect 22 965 25 982
rect 93 977 104 995
rect 22 948 34 965
rect 101 971 104 977
rect 101 960 107 971
rect 22 931 25 948
rect 93 943 107 960
rect 22 923 34 931
rect 101 942 107 943
rect 101 926 104 942
rect 93 923 104 926
rect 22 917 104 923
rect 762 919 794 923
rect 22 914 86 917
rect 22 897 25 914
rect 42 897 86 914
rect 22 880 86 897
rect 22 863 25 880
rect 42 863 86 880
rect 22 846 86 863
rect 22 829 25 846
rect 42 829 86 846
rect 762 833 763 919
rect 789 833 794 919
rect 762 832 767 833
rect 784 832 794 833
rect 762 831 794 832
rect 765 830 794 831
rect 22 679 86 829
rect 22 662 26 679
rect 43 662 86 679
rect 22 645 86 662
rect 22 628 26 645
rect 43 628 86 645
rect 22 611 86 628
rect 22 594 26 611
rect 43 594 86 611
rect 22 577 86 594
rect 22 560 26 577
rect 43 560 86 577
rect 22 543 86 560
rect 22 526 26 543
rect 43 526 86 543
rect 22 499 86 526
rect 44 498 86 499
rect 692 444 726 463
rect 759 444 786 465
<< via1 >>
rect 34 982 93 995
rect 34 965 42 982
rect 42 977 93 982
rect 42 965 84 977
rect 34 960 84 965
rect 84 960 93 977
rect 34 948 93 960
rect 34 931 42 948
rect 42 943 93 948
rect 42 931 84 943
rect 34 926 84 931
rect 84 926 93 943
rect 34 923 93 926
rect 763 902 767 919
rect 767 902 784 919
rect 784 902 789 919
rect 763 849 789 902
rect 763 833 767 849
rect 767 833 784 849
rect 784 833 789 849
<< metal2 >>
rect 79 1002 103 1049
rect 439 1022 464 1048
rect 27 995 103 1002
rect 27 923 34 995
rect 93 967 103 995
rect 93 944 481 967
rect 93 923 103 944
rect 27 920 103 923
rect 27 919 72 920
rect 458 908 481 944
rect 545 924 570 961
rect 760 919 793 923
rect 760 908 763 919
rect 188 875 407 897
rect 458 888 763 908
rect 484 887 763 888
rect 548 839 569 868
rect 760 833 763 887
rect 789 833 793 919
rect 760 830 793 833
rect 873 778 888 800
rect 443 755 468 778
rect 1 714 147 738
rect 287 714 315 738
rect 1 713 65 714
rect 873 696 888 718
rect 392 631 569 651
rect 235 596 251 614
rect 233 595 251 596
rect 211 582 251 595
rect 211 533 247 582
rect 363 550 569 571
rect 5 447 170 470
rect 283 446 309 471
<< rmetal2 >>
rect 72 919 103 920
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1629137248
transform 1 0 733 0 1 485
box 0 0 393 746
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1629137146
transform 1 0 89 0 1 1013
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1629137146
transform 1 0 173 0 1 885
box 0 0 34 33
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_2
timestamp 1628285143
transform 1 0 -90 0 1 884
box 133 -454 682 609
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1628285143
transform 1 0 241 0 -1 609
box 133 -454 682 609
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_0
timestamp 1628285143
transform 1 0 85 0 1 884
box 133 -454 682 609
<< labels >>
rlabel metal1 692 444 726 450 0 VGND
port 3 nsew ground default
rlabel metal1 759 444 786 450 0 VPWR
port 4 nsew power default
rlabel metal1 692 1044 726 1049 0 VGND
port 3 nsew ground default
rlabel metal1 759 1044 786 1049 0 VPWR
port 4 nsew power default
rlabel metal2 287 714 310 738 0 VIN11
port 7 nsew analog default
rlabel metal2 443 755 468 778 0 VIN21
port 6 nsew analog default
rlabel metal2 283 446 306 471 0 VIN12
port 8 nsew analog default
rlabel metal2 439 1022 464 1048 0 VIN22
port 5 nsew analog default
rlabel metal2 873 696 888 718 0 VOUT_AMP1
port 2 nsew analog default
rlabel metal2 873 778 888 800 0 VOUT_AMP2
port 1 nsew analog default
rlabel metal2 79 1041 103 1049 0 VPWR
port 4 nsew power default
rlabel metal2 43 714 50 738 0 VBIAS1
port 10 nsew analog default
rlabel metal2 43 447 50 470 0 VBIAS2
port 9 nsew analog default
<< end >>
