* NGSPICE file created from /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_TA2Cell_1FG_Strong.ext - technology: sky130A

.subckt sky130_hilas_nFET03 a_n62_n12# a_54_n12# $SUB a_0_n38#
X0 a_54_n12# a_0_n38# a_n62_n12# $SUB sky130_fd_pr__nfet_01v8 w=350000u l=270000u
.ends

.subckt sky130_hilas_nMirror03 sky130_hilas_nFET03_1/a_n62_n12# a_n92_86# $SUB a_168_16#
Xsky130_hilas_nFET03_0 a_n92_86# $SUB $SUB a_n92_86# sky130_hilas_nFET03
Xsky130_hilas_nFET03_1 sky130_hilas_nFET03_1/a_n62_n12# $SUB $SUB a_n92_86# sky130_hilas_nFET03
.ends

.subckt sky130_hilas_pFETmirror02 w_n122_178# a_n80_650# $SUB a_n80_262#
X0 a_n80_650# a_n80_262# w_n122_178# w_n122_178# sky130_fd_pr__pfet_01v8 w=680000u l=300000u
X1 w_n122_178# a_n80_262# a_n80_262# w_n122_178# sky130_fd_pr__pfet_01v8 w=680000u l=300000u
.ends

.subckt sky130_hilas_DualTACore01 sky130_hilas_nMirror03_3/a_n92_86# sky130_hilas_nMirror03_2/a_n92_86#
+ sky130_hilas_nMirror03_1/a_n92_86# sky130_hilas_nMirror03_0/a_n92_86# m1_n82_n44#
+ $SUB m2_n272_422# m1_52_n42# output1
Xsky130_hilas_nMirror03_3 output1 sky130_hilas_nMirror03_3/a_n92_86# $SUB m1_n82_n44#
+ sky130_hilas_nMirror03
Xsky130_hilas_pFETmirror02_0 m1_52_n42# m2_n272_422# $SUB m2_n274_n12# sky130_hilas_pFETmirror02
Xsky130_hilas_pFETmirror02_1 m1_52_n42# output1 $SUB m2_n272_1014# sky130_hilas_pFETmirror02
Xsky130_hilas_nMirror03_0 m2_n274_n12# sky130_hilas_nMirror03_0/a_n92_86# $SUB m1_n82_n44#
+ sky130_hilas_nMirror03
Xsky130_hilas_nMirror03_2 m2_n272_1014# sky130_hilas_nMirror03_2/a_n92_86# $SUB m1_n82_n44#
+ sky130_hilas_nMirror03
Xsky130_hilas_nMirror03_1 m2_n272_422# sky130_hilas_nMirror03_1/a_n92_86# $SUB m1_n82_n44#
+ sky130_hilas_nMirror03
.ends

.subckt sky130_hilas_TunCap01 $SUB a_n2872_n666# w_n2902_n800#
X0 a_n2872_n666# w_n2902_n800# w_n2902_n800# sky130_fd_pr__cap_var w=590000u l=500000u
.ends

.subckt sky130_hilas_horizTransCell01 a_n512_284# a_n952_238# a_n346_284# a_n654_284#
+ a_n926_284# $SUB a_n952_338# a_n952_496# a_n654_438# a_n926_438# a_n300_130# a_n512_162#
+ w_n728_96# a_n654_596# a_n926_596#
X0 a_n654_438# a_n952_338# a_n654_284# w_n728_96# sky130_fd_pr__pfet_g5v0d10v5 w=390000u l=500000u
X1 w_n728_96# a_n300_130# a_n344_162# w_n728_96# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
X2 a_n346_284# a_n952_238# a_n512_284# w_n728_96# sky130_fd_pr__pfet_g5v0d10v5 w=1.84e+06u l=510000u
X3 a_n344_162# a_n952_238# a_n512_162# w_n728_96# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
X4 a_n926_596# a_n952_496# a_n926_438# $SUB sky130_fd_pr__nfet_g5v0d10v5 w=400000u l=500000u
X5 a_n926_438# a_n952_338# a_n926_284# $SUB sky130_fd_pr__nfet_g5v0d10v5 w=400000u l=500000u
X6 a_n654_596# a_n952_496# a_n654_438# w_n728_96# sky130_fd_pr__pfet_g5v0d10v5 w=390000u l=500000u
.ends

.subckt sky130_hilas_FGVaractorCapacitor02 a_n1882_n644# $SUB w_n2010_n760#
X0 a_n1882_n644# w_n2010_n760# w_n2010_n760# sky130_fd_pr__cap_var w=1.11e+06u l=500000u
.ends

.subckt sky130_hilas_FGBias2x1cell Vtun GND gate_control drain1 drain4 Vinj output1
+ output2 GateColSelect
Xsky130_hilas_TunCap01_1 GND a_n560_n620# Vtun sky130_hilas_TunCap01
Xsky130_hilas_horizTransCell01_0 output2 a_n560_n620# Vinj sky130_hilas_horizTransCell01_0/a_n654_284#
+ sky130_hilas_horizTransCell01_0/a_n926_284# GND sky130_hilas_horizTransCell01_0/a_n952_338#
+ sky130_hilas_horizTransCell01_0/a_n952_496# li_934_n408# sky130_hilas_horizTransCell01_0/a_n926_438#
+ GateColSelect drain4 Vinj li_948_n216# sky130_hilas_horizTransCell01_0/a_n926_596#
+ sky130_hilas_horizTransCell01
Xsky130_hilas_TunCap01_3 GND a_n474_252# Vtun sky130_hilas_TunCap01
Xsky130_hilas_horizTransCell01_1 output1 a_n474_252# Vinj sky130_hilas_horizTransCell01_1/a_n654_284#
+ sky130_hilas_horizTransCell01_1/a_n926_284# GND sky130_hilas_horizTransCell01_1/a_n952_338#
+ sky130_hilas_horizTransCell01_1/a_n952_496# li_934_56# sky130_hilas_horizTransCell01_1/a_n926_438#
+ GateColSelect drain1 Vinj li_948_n216# sky130_hilas_horizTransCell01_1/a_n926_596#
+ sky130_hilas_horizTransCell01
Xsky130_hilas_FGVaractorCapacitor02_0 a_n560_n620# GND gate_control sky130_hilas_FGVaractorCapacitor02
Xsky130_hilas_FGVaractorCapacitor02_2 a_n474_252# GND gate_control sky130_hilas_FGVaractorCapacitor02
.ends

.subckt sky130_hilas_pTransistorVert01 a_n658_n792# a_n596_n822# a_n496_n792# $SUB
+ w_n726_n888#
X0 a_n496_n792# a_n596_n822# a_n658_n792# w_n726_n888# sky130_fd_pr__pfet_g5v0d10v5 w=2.03e+06u l=500000u
.ends

.subckt sky130_hilas_pTransistorPair m2_510_n704# w_534_n338# li_348_n384# a_454_n814#
+ $SUB a_450_n208# m2_546_n498#
Xsky130_hilas_pTransistorVert01_0 li_348_n384# a_450_n208# m2_546_n498# $SUB w_534_n338#
+ sky130_hilas_pTransistorVert01
Xsky130_hilas_pTransistorVert01_1 li_348_n384# a_454_n814# m2_510_n704# $SUB w_534_n338#
+ sky130_hilas_pTransistorVert01
.ends

.subckt sky130_hilas_FGtrans2x1cell GateSelect Vinj drain1 drain4 prog run Gate1 Gate2
+ ProgGate GND Vtun drain Vs
Xsky130_hilas_TunCap01_1 GND a_n560_n620# Vtun sky130_hilas_TunCap01
Xsky130_hilas_horizTransCell01_0 drain a_n560_n620# Vs ProgGate Gate1 GND run prog
+ li_724_n408# li_724_n408# GateSelect drain4 Vinj Gate1 ProgGate sky130_hilas_horizTransCell01
Xsky130_hilas_TunCap01_3 GND a_n474_252# Vtun sky130_hilas_TunCap01
Xsky130_hilas_horizTransCell01_1 drain1 a_n474_252# Vs ProgGate Gate2 GND run prog
+ li_724_56# li_724_56# GateSelect drain1 Vinj Gate2 ProgGate sky130_hilas_horizTransCell01
Xsky130_hilas_FGVaractorCapacitor02_0 a_n560_n620# GND li_724_n408# sky130_hilas_FGVaractorCapacitor02
Xsky130_hilas_FGVaractorCapacitor02_2 a_n474_252# GND li_724_56# sky130_hilas_FGVaractorCapacitor02
.ends

.subckt home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_TA2Cell_1FG_Strong
+ Vin+_Amp2 Vin-_Amp2 Vdd GateColSelect Vin+_Amp1 GND output2 output1 Vinj
Xsky130_hilas_DualTACore01_0 m2_n294_1062# m2_n308_1242# sky130_hilas_FGBias2x1cell_0/drain1
+ sky130_hilas_FGtrans2x1cell_0/drain GND $SUB output2 Vdd output1 sky130_hilas_DualTACore01
Xsky130_hilas_FGBias2x1cell_0 sky130_hilas_FGBias2x1cell_0/Vtun $SUB sky130_hilas_FGBias2x1cell_0/gate_control
+ sky130_hilas_FGBias2x1cell_0/drain1 sky130_hilas_FGBias2x1cell_0/drain4 Vinj sky130_hilas_FGBias2x1cell_0/output1
+ sky130_hilas_FGtrans2x1cell_0/Vs GateColSelect sky130_hilas_FGBias2x1cell
Xsky130_hilas_pTransistorPair_1 m2_n308_1242# Vinj sky130_hilas_FGBias2x1cell_0/output1
+ Vin-_Amp2 $SUB Vin+_Amp2 m2_n294_1062# sky130_hilas_pTransistorPair
Xsky130_hilas_FGtrans2x1cell_0 sky130_hilas_FGtrans2x1cell_0/GateSelect sky130_hilas_FGtrans2x1cell_0/Vinj
+ sky130_hilas_FGBias2x1cell_0/drain1 sky130_hilas_FGtrans2x1cell_0/drain4 sky130_hilas_FGtrans2x1cell_0/prog
+ sky130_hilas_FGtrans2x1cell_0/run Vin-_Amp1 Vin+_Amp1 sky130_hilas_FGtrans2x1cell_0/ProgGate
+ $SUB sky130_hilas_FGBias2x1cell_0/Vtun sky130_hilas_FGtrans2x1cell_0/drain sky130_hilas_FGtrans2x1cell_0/Vs
+ sky130_hilas_FGtrans2x1cell
.ends

