magic
tech sky130A
timestamp 1627737364
<< error_s >>
rect 309 425 336 432
rect 309 383 336 390
rect 309 333 336 340
rect 309 291 336 298
rect 309 241 336 248
rect 309 199 336 206
rect 301 135 340 138
rect 273 96 276 112
rect 301 93 340 96
rect 301 39 340 42
rect 273 0 276 16
rect 301 -3 340 0
rect 301 -57 340 -54
rect 273 -96 276 -80
rect 301 -99 340 -96
<< nwell >>
rect 401 -87 455 159
rect 383 -132 455 -87
rect 198 -150 455 -132
<< psubdiff >>
rect 397 368 439 375
rect 397 351 410 368
rect 427 351 439 368
rect 397 344 439 351
<< nsubdiff >>
rect 396 -110 437 -105
rect 396 -127 408 -110
rect 425 -127 437 -110
rect 396 -132 437 -127
<< psubdiffcont >>
rect 410 351 427 368
<< nsubdiffcont >>
rect 408 -127 425 -110
<< locali >>
rect 411 376 428 381
rect 410 373 428 376
rect 410 368 453 373
rect 427 351 453 368
rect 410 348 453 351
rect 410 342 427 348
rect 396 -127 408 -110
rect 425 -127 438 -110
<< metal1 >>
rect 409 -150 431 438
rect 449 -150 471 438
<< metal2 >>
rect 191 398 198 415
rect 389 399 471 416
rect 191 357 198 374
rect 191 306 198 323
rect 389 307 471 324
rect 191 265 198 282
rect 191 214 198 231
rect 389 215 471 232
rect 191 173 198 190
rect 191 112 198 131
rect 391 105 471 125
rect 191 70 198 89
rect 191 16 198 35
rect 391 9 471 29
rect 191 -26 198 -7
rect 191 -80 198 -61
rect 390 -87 471 -67
rect 191 -122 198 -103
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1627737364
transform 1 0 458 0 1 354
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1627737364
transform 0 1 411 -1 0 -120
box -10 -8 13 21
use sky130_hilas_nFET03a  sky130_hilas_nFET03a_3
timestamp 1627737364
transform 1 0 309 0 1 396
box -111 -47 97 42
use sky130_hilas_nFET03a  sky130_hilas_nFET03a_1
timestamp 1627737364
transform 1 0 309 0 1 304
box -111 -47 97 42
use sky130_hilas_nFET03a  sky130_hilas_nFET03a_0
timestamp 1627737364
transform 1 0 309 0 1 212
box -111 -47 97 42
use sky130_hilas_pFETdevice01e  sky130_hilas_pFETdevice01e_2
timestamp 1627737364
transform 1 0 319 0 1 -77
box -121 -55 82 44
use sky130_hilas_pFETdevice01e  sky130_hilas_pFETdevice01e_1
timestamp 1627737364
transform 1 0 319 0 1 19
box -121 -55 82 44
use sky130_hilas_pFETdevice01e  sky130_hilas_pFETdevice01e_0
timestamp 1627737364
transform 1 0 319 0 1 115
box -121 -55 82 44
<< labels >>
rlabel metal1 409 -150 431 -141 0 WELL
port 13 nsew power default
rlabel metal1 449 -150 471 -141 0 VGND
port 14 nsew ground default
rlabel metal1 409 429 431 438 0 WELL
port 13 nsew ground default
rlabel metal1 449 429 471 438 0 VGND
port 14 nsew power default
rlabel metal2 191 398 198 415 0 NFET_SOURCE1
port 1 nsew analog default
rlabel metal2 191 357 198 374 0 NFET_GATE1
port 2 nsew analog default
rlabel metal2 191 306 198 323 0 NFET_SOURCE2
port 3 nsew analog default
rlabel metal2 191 265 198 282 0 NFET_GATE2
port 4 nsew analog default
rlabel metal2 191 214 198 231 0 NFET_SOURCE3
port 5 nsew analog default
rlabel metal2 191 173 198 190 0 NFET_GATE3
port 6 nsew analog default
rlabel metal2 191 70 198 89 0 PFET_GATE1
port 8 nsew analog default
rlabel metal2 191 112 198 131 0 PFET_SOURCE1
port 7 nsew analog default
rlabel metal2 191 16 198 35 0 PFET_SOURCE2
port 9 nsew analog default
rlabel metal2 191 -26 198 -7 0 PFET_GATE2
port 10 nsew analog default
rlabel metal2 191 -80 198 -61 0 PFET_SOURCE3
port 11 nsew analog default
rlabel metal2 191 -122 198 -103 0 PFET_GATE3
port 12 nsew analog default
rlabel metal2 465 105 471 125 0 PFET_DRAIN1
port 17 nsew analog default
rlabel metal2 465 9 471 29 0 PFET_DRAIN2
port 16 nsew analog default
rlabel metal2 465 -87 471 -67 0 PFET_DRAIN3
port 15 nsew analog default
rlabel metal2 466 399 471 416 0 NFET_DRAIN1
port 20 nsew analog default
rlabel metal2 466 307 471 324 0 NFET_DRAIN2
port 19 nsew analog default
rlabel metal2 466 215 471 232 0 NFET_DRAIN3
port 18 nsew analog default
<< end >>
