magic
tech sky130A
timestamp 1624927090
<< error_p >>
rect -550 -62 -538 -50
rect -411 -57 -399 -50
rect -407 -62 -399 -57
rect -562 -69 -550 -62
rect -562 -79 -528 -69
rect -399 -70 -387 -62
rect -393 -71 -387 -70
rect -399 -74 -387 -71
rect -399 -79 -391 -74
rect -550 -84 -538 -79
rect -554 -91 -538 -84
rect -407 -87 -399 -79
rect -554 -96 -542 -91
rect -408 -96 -400 -88
rect -566 -113 -554 -96
rect -400 -101 -392 -96
rect -400 -104 -388 -101
rect -393 -105 -388 -104
rect -400 -113 -388 -105
rect -554 -125 -542 -113
rect -412 -125 -400 -113
<< mvndiff >>
rect -558 543 599 548
rect -558 526 -552 543
rect 593 526 599 543
rect -558 517 599 526
rect -558 486 -527 517
rect -558 479 599 486
rect -558 462 -552 479
rect 593 462 599 479
rect -558 455 599 462
rect -558 424 -527 455
rect -558 417 599 424
rect -558 400 -552 417
rect 592 400 599 417
rect -558 394 599 400
rect -558 364 -527 394
rect -558 357 599 364
rect -558 340 -552 357
rect 593 340 599 357
rect -558 334 599 340
rect -558 304 -527 334
rect -558 298 599 304
rect -558 281 -552 298
rect 593 281 599 298
rect -558 275 599 281
rect -558 245 -527 275
rect -558 239 599 245
rect -558 222 -552 239
rect 593 222 599 239
rect -558 216 599 222
rect -558 186 -527 216
rect -558 180 599 186
rect -558 163 -552 180
rect 592 163 599 180
rect -558 156 599 163
rect -558 125 -527 156
rect 568 155 599 156
rect -558 119 599 125
rect -558 102 -552 119
rect 593 102 599 119
rect -558 95 599 102
rect -558 64 -527 95
rect -558 57 599 64
rect -558 40 -551 57
rect 593 40 599 57
rect -558 34 599 40
rect -558 4 -527 34
rect -559 -4 599 4
rect -559 -21 -552 -4
rect 592 -21 599 -4
rect -559 -26 599 -21
<< mvndiffc >>
rect -552 526 593 543
rect -552 462 593 479
rect -552 400 592 417
rect -552 340 593 357
rect -552 281 593 298
rect -552 222 593 239
rect -552 163 592 180
rect -552 102 593 119
rect -551 40 593 57
rect -552 -21 592 -4
<< psubdiff >>
rect -528 -62 -393 -57
rect -399 -79 -393 -62
rect -528 -96 -393 -79
rect -400 -109 -393 -96
<< psubdiffcont >>
rect -550 -79 -399 -62
rect -554 -113 -400 -96
<< locali >>
rect -552 544 -535 552
rect 572 544 595 553
rect -552 543 595 544
rect -553 526 -552 543
rect 593 526 595 543
rect -553 510 595 526
rect -553 493 -519 510
rect 579 493 595 510
rect -553 479 595 493
rect -553 462 -552 479
rect 593 462 595 479
rect -553 448 595 462
rect -553 431 -519 448
rect 579 431 595 448
rect -553 417 595 431
rect -553 400 -552 417
rect 592 400 595 417
rect -553 386 595 400
rect -553 369 -518 386
rect 580 369 595 386
rect -553 357 595 369
rect -553 340 -552 357
rect 593 340 595 357
rect -553 328 595 340
rect -553 311 -516 328
rect 582 311 595 328
rect -553 298 595 311
rect -553 281 -552 298
rect 593 281 595 298
rect -553 269 595 281
rect -553 252 -515 269
rect 583 252 595 269
rect -553 239 595 252
rect -553 222 -552 239
rect 593 222 595 239
rect -553 209 595 222
rect -553 192 -515 209
rect 583 192 595 209
rect -553 180 595 192
rect -553 163 -552 180
rect 592 163 595 180
rect -553 149 595 163
rect -553 132 -520 149
rect 578 132 595 149
rect -553 119 595 132
rect -553 102 -552 119
rect 593 102 595 119
rect -553 88 595 102
rect -553 71 -519 88
rect 579 71 595 88
rect -553 57 595 71
rect -553 40 -551 57
rect 593 40 595 57
rect -553 28 595 40
rect -553 11 -520 28
rect 578 11 595 28
rect -553 -4 595 11
rect -560 -21 -552 -4
rect 592 -21 595 -4
rect -553 -27 -534 -21
rect 572 -45 595 -21
rect -523 -96 -506 -79
<< viali >>
rect -519 493 579 510
rect -519 431 579 448
rect -518 369 580 386
rect -516 311 582 328
rect -515 252 583 269
rect -515 192 583 209
rect -520 132 578 149
rect -519 71 579 88
rect -520 11 578 28
<< metal1 >>
rect -528 510 589 518
rect -528 493 -519 510
rect 579 493 589 510
rect -528 448 589 493
rect -528 431 -519 448
rect 579 431 589 448
rect -528 386 589 431
rect -528 369 -518 386
rect 580 369 589 386
rect -528 328 589 369
rect -528 311 -516 328
rect 582 311 589 328
rect -528 269 589 311
rect -528 252 -515 269
rect 583 252 589 269
rect -528 209 589 252
rect -528 192 -515 209
rect 583 192 589 209
rect -528 149 589 192
rect -528 132 -520 149
rect 578 132 589 149
rect -528 88 589 132
rect -528 71 -519 88
rect 579 71 589 88
rect -528 28 589 71
rect -528 11 -520 28
rect 578 11 589 28
rect -528 3 589 11
<< end >>
