magic
tech sky130A
timestamp 1634057737
<< nmos >>
rect 28 13 54 259
<< ndiff >>
rect 0 250 28 259
rect 0 233 5 250
rect 22 233 28 250
rect 0 216 28 233
rect 0 199 5 216
rect 22 199 28 216
rect 0 182 28 199
rect 0 165 5 182
rect 22 165 28 182
rect 0 148 28 165
rect 0 131 5 148
rect 22 131 28 148
rect 0 114 28 131
rect 0 97 5 114
rect 22 97 28 114
rect 0 80 28 97
rect 0 63 5 80
rect 22 63 28 80
rect 0 46 28 63
rect 0 29 5 46
rect 22 29 28 46
rect 0 13 28 29
rect 54 250 82 259
rect 54 233 60 250
rect 77 233 82 250
rect 54 216 82 233
rect 54 199 60 216
rect 77 199 82 216
rect 54 182 82 199
rect 54 165 60 182
rect 77 165 82 182
rect 54 148 82 165
rect 54 131 60 148
rect 77 131 82 148
rect 54 114 82 131
rect 54 97 60 114
rect 77 97 82 114
rect 54 80 82 97
rect 54 63 60 80
rect 77 63 82 80
rect 54 46 82 63
rect 54 29 60 46
rect 77 29 82 46
rect 54 13 82 29
<< ndiffc >>
rect 5 233 22 250
rect 5 199 22 216
rect 5 165 22 182
rect 5 131 22 148
rect 5 97 22 114
rect 5 63 22 80
rect 5 29 22 46
rect 60 233 77 250
rect 60 199 77 216
rect 60 165 77 182
rect 60 131 77 148
rect 60 97 77 114
rect 60 63 77 80
rect 60 29 77 46
<< poly >>
rect 28 259 54 272
rect 28 0 54 13
<< locali >>
rect 5 250 22 258
rect 5 216 22 233
rect 5 182 22 199
rect 5 148 22 165
rect 5 114 22 131
rect 5 80 22 97
rect 5 46 22 63
rect 5 18 22 29
rect 60 250 77 258
rect 60 216 77 233
rect 60 182 77 199
rect 60 148 77 165
rect 60 114 77 131
rect 60 80 77 97
rect 60 46 77 63
rect 60 18 77 29
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
