magic
tech sky130A
timestamp 1627400425
<< metal1 >>
rect 74 601 94 605
rect 657 601 676 605
rect 74 0 94 4
rect 657 0 676 4
<< metal2 >>
rect 0 574 5 594
rect 0 526 5 546
rect 0 476 6 496
rect 701 476 708 496
rect 0 411 6 431
rect 702 411 708 431
rect 0 361 5 381
rect 0 313 5 333
rect 0 272 5 292
rect 0 224 5 244
rect 0 174 6 194
rect 702 174 708 194
rect 0 109 6 129
rect 702 109 708 129
rect 0 59 5 79
rect 0 11 5 31
use sky130_hilas_TgateDouble01  sky130_hilas_TgateDouble01_2
timestamp 1608225149
transform 1 0 263 0 -1 122
box -263 -181 445 -29
use sky130_hilas_TgateDouble01  sky130_hilas_TgateDouble01_3
timestamp 1608225149
transform 1 0 263 0 1 483
box -263 -181 445 -29
use sky130_hilas_TgateDouble01  sky130_hilas_TgateDouble01_0
timestamp 1608225149
transform 1 0 263 0 -1 424
box -263 -181 445 -29
use sky130_hilas_TgateDouble01  sky130_hilas_TgateDouble01_1
timestamp 1608225149
transform 1 0 263 0 1 181
box -263 -181 445 -29
<< labels >>
rlabel metal1 657 601 676 605 0 VPWR
port 13 nsew
rlabel metal1 74 601 94 605 0 VGND
port 1 nsew ground default
rlabel metal2 701 476 708 496 0 OUTPUT1
port 17 nsew
rlabel metal2 702 174 708 194 0 OUTPUT3
port 15 nsew
rlabel metal2 702 411 708 431 0 OUTPUT2
port 16 nsew
rlabel metal2 702 109 708 129 0 OUTPUT4
port 14 nsew
rlabel metal2 0 476 6 496 0 SELECT1
port 4 nsew
rlabel metal2 0 411 6 431 0 SELECT2
port 5 nsew
rlabel metal2 0 174 6 194 0 SELECT3
port 8 nsew
rlabel metal2 0 109 6 129 0 SELECT4
port 10 nsew
rlabel metal1 657 0 676 4 0 VGND
port 1 nsew
rlabel metal1 74 0 94 4 0 VPWR
port 13 nsew
rlabel metal2 0 574 5 594 0 INPUT1_1
port 2 nsew
rlabel metal2 0 313 5 333 0 INPUT1_2
port 7 nsew
rlabel metal2 0 361 5 381 0 INPUT2_2
port 6 nsew
rlabel metal2 0 272 5 292 0 INPUT1_3
port 19 nsew
rlabel metal2 0 224 5 244 0 INPUT2_3
port 9 nsew
rlabel metal2 0 59 5 79 0 INPUT2_4
port 11 nsew
rlabel metal2 0 11 5 31 0 INPUT1_4
port 12 nsew
rlabel metal2 0 526 5 546 0 INPUT2_1
port 18 nsew
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
