magic
tech sky130A
timestamp 1608384750
<< nwell >>
rect 192 727 319 745
rect -381 571 -162 593
rect -526 410 -434 434
rect -282 410 -254 434
rect 191 140 319 159
<< metal1 >>
rect 123 731 157 745
rect 190 730 217 745
rect 123 140 157 159
rect 190 140 217 161
<< metal2 >>
rect -490 695 -466 745
rect -130 718 -105 744
rect -24 620 1 657
rect -381 571 -162 593
rect -21 535 0 564
rect 304 474 319 496
rect -126 451 -101 474
rect -526 410 -422 434
rect -282 410 -254 434
rect 304 392 319 414
rect -177 327 0 347
rect -334 292 -318 310
rect -336 291 -318 292
rect -358 278 -318 291
rect -358 229 -322 278
rect -206 246 0 267
rect -526 143 -399 166
rect -286 142 -260 167
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_0
timestamp 1608384750
transform 1 0 -484 0 1 580
box 133 -440 320 165
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1608384750
transform 1 0 -328 0 -1 305
box 133 -440 320 165
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_2
timestamp 1608384750
transform 1 0 -659 0 1 580
box 133 -440 320 165
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1607089160
transform 1 0 -396 0 1 581
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1607089160
transform 1 0 -480 0 1 682
box -14 -15 20 18
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1608069483
transform 1 0 164 0 1 181
box -172 -22 155 550
<< labels >>
rlabel metal1 123 140 157 146 0 VGND
port 3 nsew ground default
rlabel metal1 190 140 217 146 0 VPWR
port 4 nsew power default
rlabel metal1 123 740 157 745 0 VGND
port 3 nsew ground default
rlabel metal1 190 740 217 745 0 VPWR
port 4 nsew power default
rlabel metal2 -282 410 -259 434 0 VINP_AMP1
port 7 nsew analog default
rlabel metal2 -126 451 -101 474 0 VINP_AMP2
port 6 nsew analog default
rlabel metal2 -286 142 -263 167 0 VINN_AMP1
port 8 nsew analog default
rlabel metal2 -130 718 -105 744 0 VINN_AMP2
port 5 nsew analog default
rlabel metal2 304 392 319 414 0 VOUT_AMP1
port 2 nsew analog default
rlabel metal2 304 474 319 496 0 VOUT_AMP2
port 1 nsew analog default
rlabel metal2 -490 737 -466 745 0 VPWR
port 4 nsew power default
rlabel metal2 -526 410 -519 434 0 VBIAS1
port 10 nsew analog default
rlabel metal2 -526 143 -519 166 0 VBIAS2
port 9 nsew analog default
<< end >>
