magic
tech sky130A
timestamp 1628707312
<< checkpaint >>
rect 822 1649 2255 1682
rect 820 1329 2255 1649
rect 556 1290 2259 1329
rect 556 1287 2284 1290
rect 80 1208 2284 1287
rect -628 -411 2284 1208
rect -253 -519 2284 -411
rect 80 -588 2284 -519
rect 556 -601 2284 -588
rect 556 -630 2259 -601
<< error_s >>
rect 964 624 1014 630
rect 1036 624 1086 630
rect 964 582 1014 588
rect 1036 582 1086 588
rect 964 111 1014 117
rect 1036 111 1086 117
rect 964 69 1014 75
rect 1036 69 1086 75
<< nwell >>
rect 822 651 1153 652
rect 1057 648 1076 651
rect 59 187 115 429
<< psubdiff >>
rect 301 387 326 550
rect 301 370 304 387
rect 323 370 326 387
rect 301 357 326 370
rect 301 354 663 357
rect 301 353 542 354
rect 301 336 325 353
rect 344 336 368 353
rect 387 336 412 353
rect 431 336 452 353
rect 471 336 496 353
rect 515 337 542 353
rect 561 353 663 354
rect 561 337 586 353
rect 515 336 586 337
rect 605 336 632 353
rect 651 336 663 353
rect 301 332 663 336
rect 301 319 326 332
rect 301 302 304 319
rect 323 302 326 319
rect 301 148 326 302
<< mvnsubdiff >>
rect 59 187 115 429
<< psubdiffcont >>
rect 304 370 323 387
rect 325 336 344 353
rect 368 336 387 353
rect 412 336 431 353
rect 452 336 471 353
rect 496 336 515 353
rect 542 337 561 354
rect 586 336 605 353
rect 632 336 651 353
rect 304 302 323 319
<< poly >>
rect 159 563 728 580
rect 159 555 211 563
rect 441 520 460 563
rect 616 519 633 563
rect 442 136 459 169
rect 616 136 633 169
rect 116 119 727 136
<< locali >>
rect 304 387 323 395
rect 304 354 323 370
rect 304 353 542 354
rect 304 336 325 353
rect 344 336 368 353
rect 387 336 412 353
rect 431 336 452 353
rect 471 336 496 353
rect 515 337 542 353
rect 561 353 659 354
rect 561 337 586 353
rect 515 336 586 337
rect 605 336 632 353
rect 651 336 659 353
rect 304 319 323 336
rect 304 294 323 302
rect 407 232 430 236
<< metal1 >>
rect 35 47 77 652
rect 283 47 306 652
rect 405 47 428 652
rect 1057 648 1076 652
rect 1057 47 1076 52
rect 1101 47 1129 652
<< metal2 >>
rect 0 584 912 602
rect 950 478 1153 500
rect 1018 331 1136 366
rect 949 203 1153 224
rect 906 114 922 116
rect 0 109 922 114
rect 0 99 910 109
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1628707287
transform 1 0 293 0 1 337
box 0 0 23 29
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628707307
transform 1 0 934 0 1 213
box 0 0 34 33
use sky130_hilas_m12m2  sky130_hilas_m12m2_2
timestamp 1628705688
transform 1 0 1117 0 1 345
box 0 0 32 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1628705688
transform 1 0 1023 0 1 313
box 0 0 32 32
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_2
timestamp 1628705756
transform 1 0 1382 0 -1 198
box 0 0 272 169
use sky130_hilas_horizTransCell01  sky130_hilas_horizTransCell01_0
timestamp 1628705693
transform 1 0 1186 0 1 0
box 0 0 443 317
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628707307
transform 1 0 934 0 1 489
box 0 0 34 33
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1628705688
transform 1 0 1023 0 1 373
box 0 0 32 32
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_1
timestamp 1628707260
transform 1 0 1452 0 1 448
box 0 0 173 190
use sky130_hilas_wellContact  sky130_hilas_wellContact_0
timestamp 1628707306
transform 1 0 1450 0 1 660
box 0 0 173 186
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_0
timestamp 1628705756
transform 1 0 1382 0 1 491
box 0 0 272 169
use sky130_hilas_horizTransCell01  sky130_hilas_horizTransCell01_1
timestamp 1628705693
transform 1 0 1186 0 -1 699
box 0 0 443 317
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_3
timestamp 1628707260
transform 1 0 1452 0 1 862
box 0 0 173 190
use sky130_hilas_wellContact  sky130_hilas_wellContact_1
timestamp 1628707306
transform 1 0 1450 0 1 833
box 0 0 173 186
<< labels >>
rlabel metal1 35 645 77 652 0 VTUN
port 1 nsew analog default
rlabel metal1 283 645 306 652 0 VGND
port 2 nsew ground default
rlabel metal1 405 644 428 652 0 GATE_CONTROL
port 3 nsew analog default
rlabel metal1 1101 645 1129 652 0 VINJ
port 7 nsew power default
rlabel metal2 1145 478 1153 500 0 OUTPUT1
port 8 nsew analog default
rlabel metal2 1146 203 1153 224 0 OUTPUT2
port 9 nsew analog default
rlabel metal1 35 47 77 59 0 VTUN
port 1 nsew analog default
rlabel metal1 405 47 428 53 0 GATE_CONTROL
port 4 nsew analog default
rlabel metal1 283 47 306 53 0 VGND
port 2 nsew ground default
rlabel metal2 0 584 7 602 0 DRAIN1
port 5 nsew analog default
rlabel metal2 0 99 6 114 0 DRAIN4
port 6 nsew analog default
rlabel metal1 1057 648 1076 652 0 GATECOL
port 10 nsew
rlabel metal1 1057 47 1076 52 0 GATECOL
port 10 nsew
rlabel metal1 1101 47 1129 52 0 VINJ
port 11 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
