VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_capacitorSize04
  CLASS BLOCK ;
  FOREIGN sky130_hilas_capacitorSize04 ;
  ORIGIN -14.150 0.180 ;
  SIZE 5.780 BY 5.290 ;
  PIN Cap1Term02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 19.570 3.850 19.920 4.130 ;
    END
  END Cap1Term02
  PIN Cap2Term02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 19.570 0.850 19.930 1.130 ;
    END
  END Cap2Term02
  PIN Cap2Term01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 14.170 0.850 14.450 1.130 ;
    END
  END Cap2Term01
  PIN Cap1Term01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 14.170 3.850 14.420 4.130 ;
    END
  END Cap1Term01
  OBS
      LAYER met2 ;
        RECT 14.170 4.410 19.920 4.980 ;
        RECT 14.700 3.570 19.290 4.410 ;
        RECT 14.170 1.410 19.920 3.570 ;
        RECT 14.730 0.570 19.290 1.410 ;
        RECT 14.170 -0.050 19.920 0.570 ;
      LAYER met3 ;
        RECT 14.150 -0.180 19.810 5.110 ;
      LAYER met4 ;
        RECT 14.240 0.560 19.770 4.310 ;
  END
END sky130_hilas_capacitorSize04
END LIBRARY

