magic
tech sky130A
timestamp 1628617013
<< error_p >>
rect 307 88 308 91
<< nwell >>
rect 0 0 198 164
<< mvnmos >>
rect 263 33 315 65
<< mvpmos >>
rect 84 33 137 66
<< mvndiff >>
rect 235 58 263 65
rect 235 41 240 58
rect 257 41 263 58
rect 235 33 263 41
rect 315 57 343 65
rect 315 40 321 57
rect 338 40 343 57
rect 315 33 343 40
<< mvpdiff >>
rect 57 58 84 66
rect 57 41 61 58
rect 78 41 84 58
rect 57 33 84 41
rect 137 58 165 66
rect 137 41 143 58
rect 160 41 165 58
rect 137 33 165 41
<< mvndiffc >>
rect 240 41 257 58
rect 321 40 338 57
<< mvpdiffc >>
rect 61 41 78 58
rect 143 41 160 58
<< psubdiff >>
rect 307 112 351 120
rect 307 95 321 112
rect 338 95 351 112
rect 307 88 351 95
<< mvnsubdiff >>
rect 50 123 91 131
rect 50 106 62 123
rect 79 106 91 123
rect 50 97 91 106
<< psubdiffcont >>
rect 321 95 338 112
<< mvnsubdiffcont >>
rect 62 106 79 123
<< poly >>
rect 14 80 300 83
rect 14 68 315 80
rect 14 58 41 68
rect 84 66 137 68
rect 14 41 19 58
rect 36 41 41 58
rect 14 33 41 41
rect 263 65 315 68
rect 84 20 137 33
rect 263 20 315 33
<< polycont >>
rect 19 41 36 58
<< locali >>
rect 62 123 79 135
rect 62 104 64 106
rect 321 112 338 120
rect 62 94 79 104
rect 321 85 338 95
rect 19 58 36 66
rect 34 39 36 41
rect 19 33 36 39
rect 61 60 78 66
rect 61 58 86 60
rect 78 53 86 58
rect 61 36 65 41
rect 82 36 86 53
rect 135 58 160 66
rect 135 41 143 58
rect 160 41 199 58
rect 216 41 240 58
rect 257 41 265 58
rect 321 57 338 68
rect 61 33 86 36
rect 62 31 86 33
rect 143 32 160 41
rect 313 40 321 57
rect 338 40 346 57
<< viali >>
rect 64 106 79 121
rect 79 106 81 121
rect 64 104 81 106
rect 321 68 338 85
rect 17 41 19 56
rect 19 41 34 56
rect 17 39 34 41
rect 65 41 78 53
rect 78 41 82 53
rect 65 36 82 41
rect 199 41 216 58
<< metal1 >>
rect 61 126 83 160
rect 61 121 84 126
rect 61 104 64 121
rect 81 104 84 121
rect 61 100 84 104
rect 8 61 39 67
rect 8 35 11 61
rect 37 35 39 61
rect 8 32 39 35
rect 61 60 83 100
rect 318 85 341 160
rect 318 68 321 85
rect 338 68 341 85
rect 61 53 86 60
rect 61 36 65 53
rect 82 36 86 53
rect 191 36 194 62
rect 220 36 223 62
rect 61 29 86 36
rect 61 9 83 29
rect 318 9 341 68
<< via1 >>
rect 11 56 37 61
rect 11 39 17 56
rect 17 39 34 56
rect 34 39 37 56
rect 11 35 37 39
rect 194 58 220 62
rect 194 41 199 58
rect 199 41 216 58
rect 216 41 220 58
rect 194 36 220 41
<< metal2 >>
rect 0 103 361 121
rect 8 51 11 61
rect 7 35 11 51
rect 37 35 40 61
rect 191 36 194 62
rect 220 54 223 62
rect 220 36 361 54
<< labels >>
rlabel metal1 61 9 83 15 0 Vinj
rlabel metal1 61 153 83 160 0 Vinj
rlabel metal1 318 151 341 160 0 GND
rlabel metal1 318 9 341 15 0 GND
rlabel metal2 0 103 10 121 0 Input
rlabel metal2 352 103 361 121 0 Input
rlabel metal2 352 36 361 54 0 Output
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
