magic
tech sky130A
timestamp 1628704229
<< checkpaint >>
rect 821 1203 2254 1640
rect 236 1147 2254 1203
rect 189 946 2254 1147
rect -348 -224 2254 946
rect -348 -285 1519 -224
rect -348 -343 1518 -285
rect 189 -374 1518 -343
rect 190 -392 1518 -374
rect 190 -532 1516 -392
rect 233 -583 1516 -532
<< error_s >>
rect 963 582 1013 588
rect 1035 582 1085 588
rect 963 540 1013 546
rect 1035 540 1085 546
rect 720 438 722 488
rect 762 438 764 488
rect 855 438 858 488
rect 897 438 900 488
rect 720 359 722 409
rect 762 359 764 409
rect 855 359 858 409
rect 897 359 900 409
rect 720 206 722 256
rect 762 206 764 256
rect 855 206 858 256
rect 897 206 900 256
rect 720 127 722 177
rect 762 127 764 177
rect 855 127 858 177
rect 897 127 900 177
rect 963 69 1013 75
rect 1035 69 1085 75
rect 963 27 1013 33
rect 1035 27 1085 33
<< nwell >>
rect 58 145 114 387
rect 34 6 76 13
<< psubdiff >>
rect 300 345 325 508
rect 300 328 303 345
rect 322 328 325 345
rect 300 315 325 328
rect 300 312 663 315
rect 300 311 541 312
rect 300 294 324 311
rect 343 294 367 311
rect 386 294 411 311
rect 430 294 451 311
rect 470 294 495 311
rect 514 295 541 311
rect 560 311 663 312
rect 560 295 585 311
rect 514 294 585 295
rect 604 294 631 311
rect 650 294 663 311
rect 300 290 663 294
rect 300 277 325 290
rect 300 260 303 277
rect 322 260 325 277
rect 300 106 325 260
<< mvnsubdiff >>
rect 58 145 114 387
<< psubdiffcont >>
rect 303 328 322 345
rect 324 294 343 311
rect 367 294 386 311
rect 411 294 430 311
rect 451 294 470 311
rect 495 294 514 311
rect 541 295 560 312
rect 585 294 604 311
rect 631 294 650 311
rect 303 260 322 277
<< poly >>
rect 158 523 726 538
rect 158 521 714 523
rect 158 513 210 521
rect 393 478 415 521
rect 561 478 583 521
rect 671 438 709 488
rect 671 177 686 438
rect 779 359 793 360
rect 779 256 801 359
rect 671 154 711 177
rect 667 149 711 154
rect 667 132 675 149
rect 692 132 711 149
rect 667 127 711 132
rect 392 94 412 127
rect 564 94 584 127
rect 667 124 695 127
rect 115 92 712 94
rect 115 77 726 92
<< polycont >>
rect 675 132 692 149
<< locali >>
rect 781 550 869 567
rect 781 511 798 550
rect 759 494 798 511
rect 839 494 861 511
rect 616 415 724 432
rect 757 415 865 432
rect 303 345 322 353
rect 859 336 867 353
rect 303 312 322 328
rect 303 311 541 312
rect 303 294 324 311
rect 343 294 367 311
rect 386 294 411 311
rect 430 294 451 311
rect 470 294 495 311
rect 514 295 541 311
rect 560 311 658 312
rect 560 295 585 311
rect 514 294 585 295
rect 604 294 631 311
rect 650 294 658 311
rect 303 277 322 294
rect 733 279 750 336
rect 751 276 759 277
rect 817 276 822 277
rect 751 272 822 276
rect 749 268 822 272
rect 303 252 322 260
rect 742 256 826 268
rect 859 262 864 279
rect 601 183 725 200
rect 757 183 865 200
rect 675 151 692 157
rect 675 123 692 130
rect 759 120 805 121
rect 758 105 805 120
rect 759 104 805 105
rect 840 104 861 121
rect 786 70 805 104
rect 786 52 882 70
<< viali >>
rect 673 149 694 151
rect 673 132 675 149
rect 675 132 692 149
rect 692 132 694 149
rect 673 130 694 132
<< metal1 >>
rect 34 5 76 610
rect 282 5 305 610
rect 674 157 692 610
rect 669 151 698 157
rect 669 130 673 151
rect 694 130 698 151
rect 669 123 698 130
rect 674 5 692 123
rect 779 5 800 610
rect 822 5 841 610
rect 867 331 888 610
rect 1056 604 1075 610
rect 1100 605 1116 610
rect 1016 286 1040 328
rect 867 55 886 280
rect 917 55 918 56
rect 864 5 887 55
rect 1056 5 1075 10
rect 1100 5 1116 10
<< metal2 >>
rect 879 560 911 562
rect 0 542 911 560
rect 1144 542 1152 560
rect 0 387 971 406
rect 0 314 1016 318
rect 0 295 1017 314
rect 0 201 972 220
rect 905 72 921 74
rect 0 67 921 72
rect 0 57 909 67
rect 1144 55 1152 73
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_0
timestamp 1628285143
transform -1 0 -357 0 1 449
box -1005 -380 -733 -211
use sky130_hilas_wellContact  sky130_hilas_wellContact_0
timestamp 1628285143
transform 1 0 1449 0 1 618
box -1448 -441 -1275 -255
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1628285143
transform 1 0 292 0 1 295
box -10 -8 13 21
use sky130_hilas_poly2m1  sky130_hilas_poly2m1_0
timestamp 1628285143
transform 1 0 784 0 1 313
box -9 -26 24 25
use sky130_hilas_horizTransCell01a  sky130_hilas_horizTransCell01a_1
timestamp 1628285143
transform 1 0 1185 0 -1 657
box -476 42 -33 359
use sky130_hilas_horizTransCell01a  sky130_hilas_horizTransCell01a_0
timestamp 1628285143
transform 1 0 1185 0 1 -42
box -476 42 -33 359
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1628285143
transform 1 0 829 0 1 264
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_3
timestamp 1628285143
transform 1 0 875 0 1 246
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_2
timestamp 1628285143
transform 1 0 830 0 1 106
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_5
timestamp 1628285143
transform 1 0 873 0 1 55
box -10 -8 13 21
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1628285143
transform 1 0 1023 0 1 302
box -9 -10 23 22
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628285143
transform 1 0 958 0 1 221
box -14 -15 20 18
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_2
timestamp 1628285143
transform -1 0 -357 0 -1 156
box -1005 -380 -733 -211
use sky130_hilas_wellContact  sky130_hilas_wellContact_1
timestamp 1628285143
transform 1 0 1449 0 1 791
box -1448 -441 -1275 -255
use sky130_hilas_li2m1  sky130_hilas_li2m1_6
timestamp 1628285143
transform 1 0 876 0 1 552
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_4
timestamp 1628285143
transform 1 0 829 0 1 496
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_7
timestamp 1628285143
transform 1 0 876 0 1 353
box -10 -8 13 21
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628285143
transform 1 0 957 0 1 390
box -14 -15 20 18
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_1
timestamp 1628704213
transform 1 0 1451 0 1 406
box 0 0 173 190
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_3
timestamp 1628704213
transform 1 0 1451 0 1 820
box 0 0 173 190
<< labels >>
rlabel metal1 34 603 76 610 0 VTUN
port 11 nsew analog default
rlabel metal1 282 603 305 610 0 VGND
port 10 nsew ground default
rlabel space 1100 604 1116 609 0 VINJ
port 2 nsew analog default
rlabel metal2 0 57 4 72 3 DRAIN2
port 12 e analog default
rlabel metal2 0 542 6 560 0 DRAIN1
port 15 nsew analog default
rlabel metal1 822 604 841 610 0 GATE1
port 9 nsew analog default
rlabel metal1 864 6 887 30 0 VIN2
port 7 nsew analog default
rlabel metal1 674 5 692 12 0 RUN
port 6 nsew analog default
rlabel metal1 779 5 800 12 0 PROG
port 5 nsew analog default
rlabel metal1 674 603 692 610 0 RUN
port 6 nsew analog default
rlabel metal1 779 604 800 610 0 PROG
port 5 nsew analog default
rlabel metal1 867 578 888 609 0 VIN1
port 8 nsew analog default
rlabel metal1 1056 604 1075 610 0 COLSEL1
port 1 nsew analog default
rlabel metal1 1056 5 1075 10 0 COLSEL1
port 1 nsew analog default
rlabel metal1 1100 5 1116 10 0 VINJ
port 2 nsew analog default
rlabel metal2 1144 542 1152 560 0 DRAIN1
port 3 nsew analog default
rlabel metal2 1144 55 1152 73 0 DRAIN2
port 4 nsew analog default
rlabel metal1 822 6 841 11 0 GATE1
port 9 nsew analog default
rlabel metal1 282 5 305 12 0 VGND
port 10 nsew ground default
rlabel metal1 34 6 76 13 0 VTUN
port 11 nsew analog default
rlabel metal2 0 295 6 318 0 COL1
port 16 nsew
rlabel metal2 0 387 6 406 0 ROW1
port 17 nsew
rlabel metal2 0 201 6 220 0 ROW2
port 18 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
