magic
tech sky130A
magscale 1 2
timestamp 1632256366
<< checkpaint >>
rect -1260 11418 7284 16772
rect 7476 12012 11774 13848
rect 7476 11670 15122 12012
rect 15872 11670 27780 15858
rect 2876 9320 6090 11418
rect 7476 8674 27780 11670
rect 7476 7990 26572 8674
rect 3546 5484 7002 7944
rect 2408 4238 7002 5484
rect 7468 7468 26572 7990
rect 7468 6206 24594 7468
rect 7468 4410 21166 6206
rect 2408 1750 5944 4238
rect 7468 3896 15642 4410
rect 9048 2020 15642 3896
rect 9048 2014 13680 2020
<< error_s >>
rect 2522 13918 2562 13950
rect 2644 13946 2655 13957
rect 2866 13946 2964 13972
rect 2997 13950 3008 13957
rect 2997 13946 3054 13950
rect 2644 13938 3054 13946
rect 2644 13924 2866 13938
rect 2964 13918 3054 13938
rect 34 13830 72 13864
rect 22 13816 72 13830
rect 76 13794 110 13822
rect 186 13810 202 13862
rect 214 13794 230 13842
rect 318 13832 352 13864
rect 2522 13850 2523 13851
rect 2644 13850 2866 13918
rect 2964 13850 3008 13918
rect 3053 13850 3054 13851
rect 298 13822 352 13832
rect 298 13816 390 13822
rect 54 13788 106 13794
rect 352 13792 390 13816
rect 2422 13792 2456 13850
rect 2521 13849 2580 13850
rect 2522 13834 2580 13849
rect 2522 13806 2540 13834
rect 2562 13824 2580 13834
rect 2644 13824 2896 13850
rect 2964 13849 3055 13850
rect 2964 13834 3054 13849
rect 2644 13806 2866 13824
rect 2964 13806 3008 13834
rect 3034 13806 3054 13834
rect 2522 13793 2580 13806
rect 2644 13793 2896 13806
rect 2964 13794 3054 13806
rect 3008 13793 3054 13794
rect 2521 13792 2581 13793
rect 2644 13792 2897 13793
rect 2995 13792 2996 13793
rect 3008 13792 3055 13793
rect 3118 13792 3154 13850
rect 334 13790 390 13792
rect 2522 13791 2523 13792
rect 2579 13791 2580 13792
rect 54 13782 96 13788
rect 334 13782 376 13790
rect 2644 13774 2866 13792
rect 2895 13791 2896 13792
rect 2996 13791 2997 13792
rect 3053 13791 3054 13792
rect 2644 13736 3008 13774
rect 578 13662 602 13730
rect 2644 13722 2866 13736
rect 2964 13722 3008 13736
rect 2522 13692 2580 13722
rect 2866 13692 2896 13722
rect 2964 13694 3054 13722
rect 3176 13712 3188 13966
rect 2964 13683 2975 13694
rect 2996 13692 3054 13694
rect 2997 13683 3008 13692
rect 646 13662 698 13664
rect 646 13630 670 13662
rect 772 13638 824 13662
rect 2388 13656 3188 13678
rect 3430 13656 3442 13712
rect 136 13604 200 13624
rect 272 13616 334 13624
rect 142 13598 164 13604
rect 270 13602 334 13616
rect 418 13606 482 13624
rect 424 13600 446 13606
rect 108 13576 228 13596
rect 244 13588 362 13596
rect 152 13572 164 13576
rect 242 13574 362 13588
rect 390 13578 510 13596
rect 396 13572 446 13578
rect 142 13570 164 13572
rect 142 13508 152 13516
rect 234 13506 366 13526
rect 620 13510 638 13630
rect 646 13628 740 13630
rect 642 13616 740 13628
rect 646 13606 740 13616
rect 648 13582 712 13602
rect 722 13598 740 13606
rect 648 13562 666 13582
rect 694 13570 712 13582
rect 648 13538 712 13562
rect 142 13480 152 13488
rect 268 13484 332 13492
rect 266 13472 332 13484
rect 630 13464 638 13510
rect 658 13492 666 13538
rect 670 13510 724 13534
rect 2530 13506 3074 13656
rect 3410 13588 3470 13608
rect 3516 13588 3552 13590
rect 3598 13588 3752 13712
rect 3502 13568 3552 13582
rect 3430 13554 3752 13568
rect 3852 13554 4192 13588
rect 3400 13460 3410 13512
rect 698 13376 726 13394
rect 760 13376 824 13394
rect 646 13361 685 13376
rect 646 13344 670 13361
rect 772 13354 824 13376
rect 2522 13358 2580 13390
rect 2680 13358 2738 13390
rect 2838 13358 2896 13390
rect 2996 13358 3054 13390
rect 672 13344 698 13346
rect 646 13330 703 13344
rect 726 13330 771 13344
rect 646 13320 698 13330
rect 2522 13290 2523 13291
rect 2579 13290 2580 13291
rect 2680 13290 2681 13291
rect 2737 13290 2738 13291
rect 2838 13290 2839 13291
rect 2895 13290 2896 13291
rect 2996 13290 2997 13291
rect 3053 13290 3054 13291
rect 108 13230 228 13240
rect 614 13232 636 13248
rect 2422 13232 2456 13290
rect 2521 13289 2581 13290
rect 2679 13289 2739 13290
rect 2837 13289 2897 13290
rect 2995 13289 3055 13290
rect 2522 13274 2580 13289
rect 2680 13274 2738 13289
rect 2838 13274 2896 13289
rect 2996 13274 3054 13289
rect 2522 13246 2540 13274
rect 3034 13246 3054 13274
rect 2522 13233 2580 13246
rect 2680 13233 2738 13246
rect 2838 13233 2896 13246
rect 2996 13233 3054 13246
rect 2521 13232 2581 13233
rect 2679 13232 2739 13233
rect 2837 13232 2897 13233
rect 2995 13232 3055 13233
rect 3118 13232 3154 13290
rect 2522 13231 2523 13232
rect 2579 13231 2580 13232
rect 2680 13231 2681 13232
rect 2737 13231 2738 13232
rect 2838 13231 2839 13232
rect 2895 13231 2896 13232
rect 2996 13231 2997 13232
rect 3053 13231 3054 13232
rect 136 13202 200 13212
rect 2522 13132 2580 13162
rect 2680 13132 2738 13162
rect 2838 13132 2896 13162
rect 2996 13132 3054 13162
rect 662 13106 676 13112
rect 326 13062 348 13100
rect 662 13068 678 13106
rect 696 13076 712 13110
rect 304 13040 358 13062
rect 360 13032 382 13066
rect 590 13054 608 13062
rect 662 13060 676 13068
rect 2522 13048 2580 13080
rect 2680 13048 2738 13080
rect 2838 13048 2896 13080
rect 2996 13048 3054 13080
rect 2522 12980 2523 12981
rect 2579 12980 2580 12981
rect 2680 12980 2681 12981
rect 2737 12980 2738 12981
rect 2838 12980 2839 12981
rect 2895 12980 2896 12981
rect 2996 12980 2997 12981
rect 3053 12980 3054 12981
rect 2422 12922 2456 12980
rect 2521 12979 2581 12980
rect 2679 12979 2739 12980
rect 2837 12979 2897 12980
rect 2995 12979 3055 12980
rect 2522 12964 2580 12979
rect 2680 12964 2738 12979
rect 2838 12964 2896 12979
rect 2996 12964 3054 12979
rect 2522 12936 2540 12964
rect 3034 12936 3054 12964
rect 2522 12923 2580 12936
rect 2680 12923 2738 12936
rect 2838 12923 2896 12936
rect 2996 12923 3054 12936
rect 2521 12922 2581 12923
rect 2679 12922 2739 12923
rect 2837 12922 2897 12923
rect 2995 12922 3055 12923
rect 3118 12922 3154 12980
rect 2522 12921 2523 12922
rect 2579 12921 2580 12922
rect 2680 12921 2681 12922
rect 2737 12921 2738 12922
rect 2838 12921 2839 12922
rect 2895 12921 2896 12922
rect 2996 12921 2997 12922
rect 3053 12921 3054 12922
rect 268 12874 330 12896
rect 554 12878 616 12896
rect 240 12846 358 12868
rect 526 12850 644 12868
rect 3226 12852 3270 13432
rect 3430 13424 3896 13554
rect 3420 13318 3896 13424
rect 3430 13314 3644 13318
rect 3786 13316 3896 13318
rect 3430 13282 3588 13314
rect 3642 13278 3756 13314
rect 3852 13278 3896 13316
rect 3954 13278 4192 13316
rect 3954 13276 4020 13278
rect 4974 13102 5018 13182
rect 5632 13172 5690 13208
rect 5632 13108 5633 13109
rect 5689 13108 5690 13109
rect 4908 13036 5084 13102
rect 5532 13050 5568 13108
rect 5631 13107 5691 13108
rect 5632 13088 5690 13107
rect 5632 13070 5652 13088
rect 5670 13070 5690 13088
rect 5632 13051 5690 13070
rect 5631 13050 5691 13051
rect 5754 13050 5790 13108
rect 5632 13049 5633 13050
rect 5689 13049 5690 13050
rect 4908 13014 5142 13036
rect 4908 12948 5084 13014
rect 5632 12950 5690 12986
rect 2522 12822 2580 12852
rect 2680 12822 2738 12852
rect 2838 12822 2896 12852
rect 2996 12822 3054 12852
rect 810 12802 812 12812
rect 290 12770 292 12798
rect 430 12770 432 12798
rect 578 12770 580 12798
rect 256 12736 292 12764
rect 396 12736 432 12764
rect 544 12736 580 12764
rect 588 12758 646 12762
rect 762 12756 788 12762
rect 1304 12748 3038 12762
rect 2944 12744 3038 12748
rect 616 12730 674 12734
rect 762 12728 816 12734
rect 1304 12720 3066 12734
rect 2916 12716 3066 12720
rect 8924 12502 9278 12656
rect 9480 12490 9532 12586
rect 9678 12522 9734 12534
rect 9798 12502 9834 12586
rect 9962 12520 10018 12534
rect 10232 12522 10332 12534
rect 10170 12520 10388 12522
rect 9984 12502 10388 12520
rect 16574 12502 16584 12510
rect 8934 12414 8974 12432
rect 9480 12378 9834 12490
rect 10052 12482 10196 12502
rect 10388 12483 10456 12502
rect 10373 12482 10456 12483
rect 16456 12482 16584 12502
rect 10052 12468 10456 12482
rect 16573 12471 16584 12482
rect 24164 12502 24174 12510
rect 24164 12482 24292 12502
rect 24164 12471 24175 12482
rect 10052 12450 10388 12468
rect 9962 12436 10018 12450
rect 10052 12446 10088 12450
rect 10122 12446 10158 12450
rect 10018 12420 10030 12432
rect 10000 12386 10008 12402
rect 10052 12386 10158 12446
rect 10182 12438 10382 12450
rect 10182 12418 10232 12438
rect 10254 12407 10322 12422
rect 10332 12418 10382 12438
rect 10388 12414 10426 12424
rect 10422 12396 10476 12406
rect 10484 12396 10552 12446
rect 10172 12386 10178 12396
rect 10206 12386 10312 12396
rect 9340 12366 9834 12378
rect 9874 12378 10312 12386
rect 10422 12378 10552 12396
rect 9874 12366 10484 12378
rect 9368 12338 9460 12350
rect 8924 12170 9278 12306
rect 9480 12268 9834 12366
rect 9966 12360 10088 12366
rect 10116 12363 10178 12366
rect 10122 12360 10178 12363
rect 10254 12362 10484 12366
rect 10236 12360 10518 12362
rect 9966 12358 10017 12360
rect 10036 12358 10088 12360
rect 10159 12358 10518 12360
rect 9874 12350 10518 12358
rect 9874 12338 10278 12350
rect 9976 12336 10116 12338
rect 9978 12332 10116 12336
rect 10128 12334 10278 12338
rect 10036 12321 10116 12332
rect 10021 12307 10116 12321
rect 10126 12332 10278 12334
rect 10126 12312 10274 12332
rect 10126 12307 10242 12312
rect 10312 12310 10313 12350
rect 10322 12320 10374 12350
rect 10021 12306 10242 12307
rect 10280 12307 10313 12310
rect 10438 12307 10470 12350
rect 10472 12344 10518 12350
rect 10472 12328 10526 12344
rect 10476 12307 10536 12328
rect 10540 12307 10552 12378
rect 10280 12306 10552 12307
rect 10052 12294 10116 12306
rect 10244 12302 10278 12306
rect 10280 12302 10330 12306
rect 9528 12250 9562 12264
rect 10020 12254 10022 12264
rect 10052 12258 10088 12294
rect 10180 12290 10330 12302
rect 10438 12294 10470 12306
rect 10118 12266 10482 12290
rect 10036 12244 10088 12258
rect 10116 12260 10482 12266
rect 10116 12250 10322 12260
rect 10342 12252 10482 12260
rect 10052 12238 10088 12244
rect 10118 12240 10322 12250
rect 10102 12238 10456 12240
rect 9480 12222 9562 12236
rect 8774 12100 8802 12164
rect 8972 12152 8974 12166
rect 9480 12140 9532 12222
rect 9678 12172 9734 12184
rect 9962 12170 10018 12184
rect 10052 12172 10456 12238
rect 10052 12157 10232 12172
rect 10342 12164 10456 12172
rect 4690 11780 4698 11830
rect 4724 11802 4732 11854
rect 8924 11820 9278 11956
rect 9480 11918 9834 12140
rect 10052 12132 10196 12157
rect 10388 12133 10456 12164
rect 10373 12132 10456 12133
rect 10052 12118 10456 12132
rect 10052 12100 10388 12118
rect 9962 12086 10018 12100
rect 10052 12096 10088 12100
rect 10122 12096 10158 12100
rect 10018 12070 10030 12082
rect 10000 12036 10008 12052
rect 10052 12036 10158 12096
rect 10182 12088 10382 12100
rect 10182 12068 10232 12088
rect 10254 12057 10322 12072
rect 10332 12068 10382 12088
rect 10484 12092 10552 12096
rect 10484 12074 10566 12092
rect 10172 12036 10178 12046
rect 10194 12036 10318 12048
rect 10000 12028 10318 12036
rect 10422 12046 10476 12056
rect 10484 12046 10552 12074
rect 10422 12028 10552 12046
rect 10000 12026 10484 12028
rect 10002 12024 10484 12026
rect 10002 12018 10088 12024
rect 9966 12010 10088 12018
rect 10116 12013 10178 12024
rect 10206 12016 10484 12024
rect 10122 12010 10178 12013
rect 10222 12012 10484 12016
rect 10222 12010 10518 12012
rect 9966 12008 10017 12010
rect 10036 12008 10088 12010
rect 10159 12008 10518 12010
rect 9966 12000 10518 12008
rect 9966 11996 10290 12000
rect 9966 11994 10098 11996
rect 10159 11995 10290 11996
rect 10172 11994 10290 11995
rect 9966 11992 10116 11994
rect 9976 11986 10116 11992
rect 9978 11982 10116 11986
rect 10128 11984 10278 11994
rect 10036 11971 10116 11982
rect 10021 11957 10116 11971
rect 10126 11982 10278 11984
rect 10126 11962 10274 11982
rect 10126 11957 10242 11962
rect 10312 11960 10313 12000
rect 10322 11970 10374 12000
rect 10021 11956 10242 11957
rect 10280 11957 10313 11960
rect 10438 11957 10470 12000
rect 10472 11994 10518 12000
rect 10472 11978 10526 11994
rect 10476 11957 10536 11978
rect 10540 11957 10552 12028
rect 10280 11956 10552 11957
rect 10052 11944 10116 11956
rect 10244 11952 10278 11956
rect 10280 11952 10330 11956
rect 9528 11900 9576 11914
rect 10020 11904 10022 11914
rect 10052 11908 10088 11944
rect 10180 11940 10330 11952
rect 10438 11944 10470 11956
rect 10480 11940 10514 11956
rect 10118 11936 10514 11940
rect 10118 11916 10482 11936
rect 16306 11922 16316 11940
rect 10036 11894 10088 11908
rect 10116 11910 10482 11916
rect 10116 11900 10322 11910
rect 10342 11902 10482 11910
rect 10052 11888 10088 11894
rect 10118 11890 10322 11900
rect 16334 11894 16400 11920
rect 16514 11916 16526 12010
rect 16542 11944 16554 12038
rect 16780 11894 16996 11920
rect 17358 11918 17390 11946
rect 17440 11916 17478 11944
rect 22800 11928 23462 12094
rect 24194 11968 24206 12038
rect 24222 11968 24234 12010
rect 24036 11956 24136 11968
rect 24180 11956 24280 11968
rect 24194 11944 24206 11956
rect 23270 11926 23308 11928
rect 23270 11920 23438 11926
rect 10102 11888 10456 11890
rect 9480 11872 9576 11886
rect 8972 11788 9020 11816
rect 9480 11790 9532 11872
rect 9678 11822 9734 11834
rect 9962 11820 10018 11834
rect 10052 11822 10456 11888
rect 16400 11884 16780 11894
rect 16468 11856 16568 11884
rect 16612 11868 16712 11884
rect 16996 11868 17022 11894
rect 23968 11884 24036 11928
rect 24136 11884 24180 11928
rect 24222 11916 24234 11956
rect 24280 11884 24348 11928
rect 23980 11874 24004 11876
rect 24036 11874 24136 11884
rect 24180 11874 24280 11884
rect 16468 11852 16526 11856
rect 9576 11802 9622 11818
rect 10052 11807 10232 11822
rect 10342 11814 10456 11822
rect 4108 11756 4178 11758
rect 8794 11750 8802 11786
rect 4136 11676 4164 11730
rect 4532 11678 4696 11700
rect 4572 11672 4598 11678
rect 4108 11648 4192 11672
rect 4504 11662 4724 11672
rect 4504 11656 4744 11662
rect 4504 11654 4746 11656
rect 4512 11650 4746 11654
rect 4542 11642 4598 11650
rect 4724 11646 4746 11650
rect 4542 11632 4608 11642
rect 4696 11640 4716 11646
rect 4544 11630 4570 11632
rect 4572 11630 4598 11632
rect 4544 11596 4636 11630
rect 4548 11568 4636 11596
rect 4692 11588 4716 11640
rect 4724 11612 4748 11646
rect 4724 11604 4746 11612
rect 4724 11598 4744 11604
rect 4692 11582 4700 11588
rect 4136 11492 4164 11526
rect 4164 11410 4170 11444
rect 4192 11438 4198 11472
rect 4254 11438 4256 11486
rect 4192 11428 4256 11438
rect 4282 11410 4284 11468
rect 4478 11410 4492 11416
rect 4506 11410 4520 11444
rect 4164 11400 4284 11410
rect 4544 11398 4570 11462
rect 4572 11378 4598 11490
rect 8924 11470 9278 11606
rect 9480 11568 9834 11790
rect 10052 11782 10196 11807
rect 10388 11783 10456 11814
rect 10373 11782 10456 11783
rect 10052 11768 10456 11782
rect 16400 11826 16468 11828
rect 16480 11826 16526 11852
rect 16612 11838 17220 11868
rect 17796 11858 17834 11864
rect 23980 11858 24350 11874
rect 16400 11822 16574 11826
rect 16614 11822 16716 11838
rect 16952 11834 17084 11838
rect 10052 11750 10388 11768
rect 16400 11754 16780 11822
rect 16844 11768 16922 11822
rect 16996 11768 17022 11834
rect 17114 11768 17194 11822
rect 17286 11792 17314 11828
rect 17796 11824 17798 11858
rect 17818 11824 17834 11858
rect 17796 11818 17834 11824
rect 17852 11808 17868 11842
rect 23986 11836 24350 11858
rect 23986 11822 24030 11836
rect 24128 11830 24350 11836
rect 24128 11822 24134 11830
rect 24222 11822 24268 11830
rect 23986 11782 24032 11822
rect 9962 11736 10018 11750
rect 10052 11746 10088 11750
rect 10122 11746 10158 11750
rect 10018 11720 10030 11732
rect 10000 11686 10008 11702
rect 10052 11686 10158 11746
rect 10182 11738 10382 11750
rect 10182 11718 10232 11738
rect 10254 11707 10322 11722
rect 10332 11718 10382 11738
rect 10484 11742 10552 11746
rect 10484 11724 10566 11742
rect 10172 11686 10178 11696
rect 10194 11686 10318 11698
rect 10000 11678 10318 11686
rect 10422 11696 10476 11706
rect 10484 11696 10552 11724
rect 16372 11723 16780 11754
rect 16818 11723 17220 11768
rect 17878 11730 17890 11740
rect 16361 11713 16780 11723
rect 16807 11713 17231 11723
rect 16334 11712 17231 11713
rect 10422 11678 10552 11696
rect 10000 11676 10484 11678
rect 10002 11674 10484 11676
rect 10002 11668 10088 11674
rect 9966 11660 10088 11668
rect 10116 11663 10178 11674
rect 10206 11666 10484 11674
rect 10122 11660 10178 11663
rect 10222 11662 10484 11666
rect 10222 11660 10518 11662
rect 9966 11658 10017 11660
rect 10036 11658 10088 11660
rect 10159 11658 10518 11660
rect 9966 11650 10518 11658
rect 9966 11646 10290 11650
rect 9966 11644 10098 11646
rect 10159 11645 10290 11646
rect 10172 11644 10290 11645
rect 9966 11642 10116 11644
rect 9976 11636 10116 11642
rect 9978 11632 10116 11636
rect 10128 11634 10278 11644
rect 10036 11621 10116 11632
rect 10021 11607 10116 11621
rect 10126 11632 10278 11634
rect 10126 11612 10274 11632
rect 10126 11607 10242 11612
rect 10312 11610 10313 11650
rect 10322 11620 10374 11650
rect 10021 11606 10242 11607
rect 10280 11607 10313 11610
rect 10438 11607 10470 11650
rect 10472 11644 10518 11650
rect 10472 11628 10526 11644
rect 10476 11607 10536 11628
rect 10540 11607 10552 11678
rect 16528 11660 16530 11712
rect 16556 11654 16656 11712
rect 16838 11668 16844 11712
rect 16922 11668 16928 11712
rect 17110 11668 17114 11712
rect 17194 11668 17198 11712
rect 23986 11692 24030 11782
rect 24128 11672 24190 11822
rect 24244 11804 24350 11822
rect 24294 11768 24350 11804
rect 24222 11720 24268 11722
rect 24214 11672 24268 11720
rect 24292 11672 24350 11722
rect 10280 11606 10552 11607
rect 16456 11638 16548 11654
rect 16456 11622 16550 11638
rect 16556 11632 16574 11654
rect 10052 11594 10116 11606
rect 10244 11602 10278 11606
rect 10280 11602 10330 11606
rect 9528 11550 9576 11564
rect 10020 11554 10022 11564
rect 10052 11558 10088 11594
rect 10180 11590 10330 11602
rect 10438 11594 10470 11606
rect 10476 11590 10514 11606
rect 10118 11586 10514 11590
rect 16456 11594 16548 11622
rect 16558 11594 16574 11632
rect 23000 11624 23024 11630
rect 23030 11626 23034 11636
rect 16456 11586 16574 11594
rect 10118 11566 10482 11586
rect 10036 11544 10088 11558
rect 10116 11560 10482 11566
rect 10116 11550 10322 11560
rect 10342 11552 10482 11560
rect 10052 11538 10088 11544
rect 10118 11540 10322 11550
rect 10102 11538 10456 11540
rect 9480 11522 9576 11536
rect 4692 11384 4700 11434
rect 4726 11406 4734 11458
rect 8794 11400 8802 11456
rect 8972 11438 9020 11466
rect 9480 11438 9532 11522
rect 9678 11472 9734 11484
rect 9962 11470 10018 11484
rect 10052 11472 10456 11538
rect 9576 11452 9622 11468
rect 10052 11457 10232 11472
rect 10342 11464 10456 11472
rect 10052 11432 10196 11457
rect 10388 11433 10456 11464
rect 10373 11432 10456 11433
rect 10052 11418 10456 11432
rect 10052 11400 10388 11418
rect 9678 11388 9734 11400
rect 9962 11386 10018 11400
rect 10052 11396 10088 11400
rect 10122 11396 10158 11400
rect 4532 11366 4710 11378
rect 4136 11336 4164 11342
rect 4136 11308 4178 11336
rect 4456 11306 4498 11332
rect 4524 11328 4532 11338
rect 4556 11320 4648 11336
rect 4188 11280 4206 11296
rect 4460 11294 4462 11306
rect 4488 11298 4490 11304
rect 4460 11286 4468 11294
rect 4460 11280 4462 11286
rect 4160 11226 4168 11260
rect 4188 11254 4196 11280
rect 4488 11272 4532 11298
rect 4488 11258 4496 11272
rect 4488 11254 4494 11258
rect 4544 11254 4552 11304
rect 4556 11256 4558 11278
rect 4188 11230 4250 11254
rect 4460 11226 4466 11254
rect 4488 11240 4552 11254
rect 4520 11226 4524 11240
rect 4160 11202 4278 11226
rect 4460 11212 4552 11226
rect 4572 11212 4580 11320
rect 4716 11206 4722 11256
rect 4750 11226 4756 11278
rect 4364 11192 4496 11198
rect 4542 11192 4593 11197
rect 4542 11184 4598 11192
rect 4392 11164 4468 11170
rect 4136 11104 4164 11142
rect 4460 11134 4506 11136
rect 4544 11134 4570 11164
rect 4460 11112 4570 11134
rect 4460 11110 4506 11112
rect 4460 11102 4462 11110
rect 4488 11100 4506 11108
rect 4512 11106 4570 11112
rect 4544 11100 4570 11106
rect 4488 11092 4554 11100
rect 4488 11080 4556 11092
rect 4488 11078 4558 11080
rect 4488 11056 4494 11078
rect 4460 11042 4466 11056
rect 4488 11048 4524 11056
rect 4488 11042 4494 11048
rect 4520 11018 4524 11048
rect 4544 11042 4552 11078
rect 4556 11058 4558 11078
rect 4572 11072 4598 11184
rect 8746 11134 8782 11142
rect 8924 11120 9278 11270
rect 9480 11218 9532 11374
rect 10018 11370 10030 11382
rect 9580 11328 9636 11340
rect 10000 11336 10008 11352
rect 10052 11336 10158 11396
rect 10182 11388 10382 11400
rect 10182 11368 10232 11388
rect 10254 11357 10322 11372
rect 10332 11368 10382 11388
rect 10484 11392 10552 11396
rect 10484 11374 10566 11392
rect 16334 11388 16340 11512
rect 16494 11456 16520 11586
rect 16522 11484 16548 11586
rect 16838 11512 16844 11610
rect 16922 11512 16928 11610
rect 16558 11498 16600 11502
rect 16614 11498 16626 11502
rect 16512 11448 16520 11456
rect 16540 11448 16548 11456
rect 16558 11454 16626 11498
rect 16504 11400 16572 11448
rect 16540 11378 16548 11400
rect 16690 11388 16996 11512
rect 17110 11510 17114 11610
rect 17194 11510 17198 11610
rect 23028 11602 23056 11626
rect 23068 11614 23092 11616
rect 23068 11608 23090 11614
rect 22934 11584 23014 11598
rect 23028 11574 23056 11598
rect 23102 11580 23126 11582
rect 23102 11576 23124 11580
rect 17796 11460 17834 11466
rect 17796 11426 17798 11460
rect 17822 11426 17834 11448
rect 17796 11420 17834 11426
rect 17856 11380 17890 11414
rect 10172 11336 10178 11346
rect 10194 11336 10318 11348
rect 10000 11328 10318 11336
rect 10422 11346 10476 11356
rect 10484 11346 10552 11374
rect 17530 11364 17544 11370
rect 10422 11328 10552 11346
rect 10000 11326 10484 11328
rect 10002 11324 10484 11326
rect 10002 11318 10088 11324
rect 9966 11310 10088 11318
rect 10116 11313 10178 11324
rect 10206 11316 10484 11324
rect 10122 11310 10178 11313
rect 10222 11312 10484 11316
rect 10222 11310 10518 11312
rect 9966 11308 10017 11310
rect 10036 11308 10088 11310
rect 10159 11308 10518 11310
rect 9966 11300 10518 11308
rect 9966 11296 10290 11300
rect 9966 11294 10098 11296
rect 10159 11295 10290 11296
rect 10172 11294 10290 11295
rect 9966 11292 10116 11294
rect 9976 11286 10116 11292
rect 9978 11282 10116 11286
rect 10128 11284 10278 11294
rect 10036 11271 10116 11282
rect 10021 11257 10116 11271
rect 10126 11282 10278 11284
rect 10126 11262 10274 11282
rect 10126 11257 10242 11262
rect 10312 11260 10313 11300
rect 10322 11270 10374 11300
rect 10021 11256 10242 11257
rect 10280 11257 10313 11260
rect 10438 11257 10470 11300
rect 10472 11294 10518 11300
rect 10472 11278 10526 11294
rect 10476 11257 10536 11278
rect 10540 11257 10552 11328
rect 17528 11318 17544 11364
rect 17558 11336 17572 11344
rect 16572 11296 16582 11304
rect 17556 11298 17572 11336
rect 17938 11306 17946 11464
rect 17966 11334 17974 11436
rect 16454 11276 16582 11296
rect 10280 11256 10552 11257
rect 9580 11244 9636 11256
rect 10052 11244 10116 11256
rect 10244 11252 10278 11256
rect 10280 11252 10330 11256
rect 10052 11218 10088 11244
rect 10180 11240 10330 11252
rect 10438 11244 10470 11256
rect 10482 11240 10514 11256
rect 10020 11204 10022 11214
rect 10118 11195 10131 11240
rect 10280 11236 10514 11240
rect 10280 11222 10482 11236
rect 10278 11212 10482 11222
rect 10280 11210 10482 11212
rect 10342 11202 10482 11210
rect 10180 11156 10280 11168
rect 4572 11014 4580 11072
rect 4716 11008 4722 11058
rect 4750 11028 4756 11080
rect 8774 11050 8802 11114
rect 8934 11014 8982 11042
rect 9522 11014 9584 11042
rect 10388 11014 10446 11042
rect 16512 11036 16520 11240
rect 16540 11064 16548 11268
rect 16571 11265 16582 11276
rect 17890 11282 17928 11288
rect 17890 11278 17906 11282
rect 17912 11278 17928 11282
rect 17890 11266 17928 11278
rect 17798 11246 17836 11252
rect 16560 11224 16582 11246
rect 16552 11192 16606 11224
rect 17798 11212 17800 11246
rect 17828 11212 17836 11246
rect 17862 11242 17928 11266
rect 18076 11262 18738 11320
rect 17946 11260 17980 11262
rect 18072 11260 18738 11262
rect 17946 11254 17962 11260
rect 17862 11232 17896 11242
rect 17938 11220 17962 11254
rect 18056 11232 18738 11260
rect 17798 11206 17836 11212
rect 16558 11186 16582 11192
rect 16558 11156 16600 11186
rect 16564 11154 16600 11156
rect 17618 11150 17674 11176
rect 18076 11154 18738 11232
rect 18076 11152 18434 11154
rect 4542 10994 4593 10999
rect 4542 10986 4598 10994
rect 4122 10946 4164 10974
rect 4544 10960 4570 10966
rect 4136 10912 4164 10946
rect 4392 10902 4570 10960
rect 4122 10866 4164 10890
rect 4122 10862 4136 10866
rect 4150 10842 4164 10866
rect 4392 10882 4556 10902
rect 4392 10860 4558 10882
rect 4572 10874 4598 10986
rect 16512 10986 16528 11036
rect 16540 11014 16556 11064
rect 16838 11036 16844 11136
rect 16922 11036 16928 11136
rect 17110 11036 17114 11136
rect 17194 11036 17198 11136
rect 17646 11122 17702 11148
rect 18088 11062 18100 11152
rect 18116 11150 18180 11152
rect 18188 11150 18208 11152
rect 18116 11090 18128 11150
rect 18160 11090 18284 11150
rect 18576 11104 18592 11154
rect 18604 11132 18646 11154
rect 18698 11138 18736 11154
rect 18780 11142 18822 11170
rect 18188 11062 18208 11090
rect 18076 11018 18104 11054
rect 16512 10958 16530 10986
rect 16540 10958 16558 11014
rect 4392 10844 4556 10860
rect 4572 10844 4580 10874
rect 4150 10834 4192 10842
rect 4392 10820 4628 10844
rect 4392 10790 4636 10820
rect 4392 10788 4598 10790
rect 4122 10748 4164 10776
rect 4392 10768 4556 10788
rect 4392 10748 4570 10768
rect 4136 10720 4570 10748
rect 4150 10706 4570 10720
rect 4150 10616 4520 10706
rect 4544 10704 4570 10706
rect 4572 10676 4598 10788
rect 4624 10774 4636 10790
rect 4652 10746 4664 10848
rect 4716 10810 4722 10860
rect 4750 10830 4756 10882
rect 8946 10802 9300 10948
rect 8994 10780 9042 10802
rect 9582 10780 9644 10808
rect 10074 10802 10574 10948
rect 16469 10947 16582 10958
rect 16480 10926 16534 10947
rect 16540 10934 16582 10947
rect 16480 10916 16526 10926
rect 16540 10916 16586 10934
rect 11730 10810 11904 10916
rect 16480 10910 16586 10916
rect 16480 10900 16582 10910
rect 16480 10892 16554 10900
rect 11730 10808 12066 10810
rect 10448 10772 10506 10802
rect 11730 10748 11762 10808
rect 11898 10740 11930 10808
rect 16412 10770 16414 10774
rect 16458 10764 16460 10832
rect 16480 10821 16526 10892
rect 16532 10876 16554 10892
rect 16469 10816 16537 10821
rect 16540 10816 16554 10876
rect 16558 10876 16582 10900
rect 16838 10878 16844 10978
rect 16922 10878 16928 10978
rect 17110 10878 17114 10978
rect 17194 10878 17198 10978
rect 17876 10950 17888 10960
rect 18038 10950 18074 10952
rect 18072 10948 18074 10950
rect 19296 10932 19540 11548
rect 21208 11166 21452 11548
rect 23062 11528 23082 11562
rect 23102 11536 23116 11576
rect 23388 11568 23414 11656
rect 24092 11654 24190 11672
rect 23416 11568 23442 11628
rect 23140 11560 23152 11562
rect 23062 11514 23076 11528
rect 22934 11500 23014 11514
rect 23228 11508 23456 11544
rect 22986 11462 22994 11484
rect 22934 11450 23014 11462
rect 22872 11402 22888 11418
rect 22894 11402 22902 11420
rect 22958 11418 22966 11450
rect 22986 11446 22994 11450
rect 23010 11402 23020 11412
rect 22888 11386 22904 11392
rect 23026 11386 23042 11402
rect 22934 11366 23014 11378
rect 23130 11340 23456 11508
rect 23752 11388 24054 11602
rect 24174 11586 24190 11654
rect 24202 11644 24292 11654
rect 24214 11610 24292 11644
rect 24214 11594 24284 11610
rect 24118 11498 24134 11502
rect 24148 11498 24190 11502
rect 24118 11454 24190 11498
rect 24200 11448 24204 11456
rect 24228 11448 24232 11484
rect 24172 11400 24244 11448
rect 24172 11376 24194 11392
rect 24200 11378 24204 11400
rect 24404 11388 24414 11512
rect 23192 11334 23390 11340
rect 23192 11332 23202 11334
rect 22670 11290 22938 11320
rect 23000 11290 23322 11304
rect 22244 11206 22246 11222
rect 22220 11166 22248 11206
rect 22368 11204 22408 11232
rect 22570 11166 22634 11258
rect 21174 11138 21452 11166
rect 21208 10932 21452 11138
rect 22244 11130 22246 11166
rect 22478 11138 22516 11166
rect 22566 11154 22634 11166
rect 22570 11150 22634 11154
rect 22670 11152 22888 11290
rect 22894 11198 22908 11290
rect 23186 11240 23322 11290
rect 23596 11286 23634 11310
rect 23654 11286 23662 11318
rect 22894 11188 22916 11198
rect 22900 11174 22916 11188
rect 21970 11088 22016 11122
rect 22246 11054 22412 11130
rect 22634 11090 22738 11150
rect 22770 11122 22888 11152
rect 22974 11136 23322 11240
rect 23440 11264 23696 11286
rect 23440 11246 23726 11264
rect 23906 11258 23950 11348
rect 24106 11336 24118 11354
rect 24072 11302 24084 11336
rect 24106 11320 24122 11336
rect 24072 11286 24090 11302
rect 24162 11296 24172 11304
rect 24162 11276 24290 11296
rect 24162 11265 24173 11276
rect 23440 11236 23696 11246
rect 23440 11206 23712 11236
rect 23752 11220 23950 11258
rect 23724 11214 23950 11220
rect 24062 11218 24084 11246
rect 24162 11224 24188 11246
rect 24032 11214 24084 11218
rect 23724 11212 24084 11214
rect 23724 11206 23950 11212
rect 22974 11122 23396 11136
rect 22770 11016 23396 11122
rect 23408 11096 23414 11182
rect 23440 11180 23950 11206
rect 24032 11198 24084 11212
rect 24062 11192 24084 11198
rect 24138 11192 24192 11224
rect 23968 11180 24084 11192
rect 24162 11186 24190 11192
rect 23440 11178 24084 11180
rect 23440 11158 23950 11178
rect 23968 11158 24084 11178
rect 23440 11154 24084 11158
rect 24148 11156 24190 11186
rect 24148 11154 24184 11156
rect 23436 11136 24084 11154
rect 23436 11124 23696 11136
rect 23440 11118 23696 11124
rect 23724 11128 24084 11136
rect 23724 11124 23950 11128
rect 23968 11124 24084 11128
rect 23724 11118 24084 11124
rect 23736 11110 23920 11118
rect 23752 11102 23920 11110
rect 23740 11100 23920 11102
rect 23458 11092 23490 11100
rect 23564 11092 23682 11094
rect 23736 11074 23920 11100
rect 23948 11094 24084 11118
rect 23964 11090 24084 11094
rect 23968 11078 24084 11090
rect 23430 11064 23462 11072
rect 23592 11064 23654 11066
rect 23560 11048 23592 11064
rect 23674 11062 23736 11074
rect 23594 11048 23626 11058
rect 23560 11016 23626 11048
rect 23650 11050 23658 11058
rect 23650 11016 23660 11050
rect 23674 11037 23694 11062
rect 23684 11020 23694 11037
rect 23706 11020 23724 11062
rect 23728 11059 23736 11062
rect 23740 11034 23758 11074
rect 23790 11073 23920 11074
rect 23802 11036 23842 11052
rect 23852 11036 23920 11073
rect 23948 11054 24084 11078
rect 24200 11064 24204 11268
rect 23948 11048 23964 11054
rect 23968 11048 24084 11054
rect 23790 11034 23852 11036
rect 23752 11026 23858 11034
rect 23736 11020 23858 11026
rect 23674 11016 23858 11020
rect 22220 10970 22248 11010
rect 22770 10986 23414 11016
rect 23560 11000 23858 11016
rect 23560 10998 23592 11000
rect 23416 10986 23442 10988
rect 22770 10978 23442 10986
rect 23564 10978 23570 10998
rect 23624 10996 23858 11000
rect 22770 10968 23228 10978
rect 22950 10958 22962 10968
rect 22934 10944 23014 10958
rect 22950 10940 22962 10944
rect 23130 10942 23184 10958
rect 23388 10952 23414 10978
rect 23416 10952 23442 10978
rect 23596 10968 23858 10996
rect 23612 10966 23858 10968
rect 23648 10964 23662 10966
rect 23674 10965 23858 10966
rect 23872 10965 23898 11036
rect 23948 10996 24084 11048
rect 24192 11014 24204 11064
rect 24228 11036 24232 11240
rect 23968 10980 24084 10996
rect 23674 10964 23898 10965
rect 22876 10922 23076 10934
rect 22876 10888 23082 10922
rect 23102 10896 23116 10942
rect 23140 10920 23152 10922
rect 23228 10888 23456 10952
rect 23624 10914 23778 10964
rect 23964 10948 24084 10980
rect 24190 10958 24204 11014
rect 24220 10986 24232 11036
rect 24218 10958 24232 10986
rect 24162 10954 24279 10958
rect 23674 10896 23728 10900
rect 23752 10896 23858 10914
rect 17720 10882 17808 10884
rect 16558 10846 16586 10876
rect 17748 10854 17800 10870
rect 16558 10824 16582 10846
rect 16464 10810 16466 10816
rect 16468 10810 16582 10816
rect 16410 10756 16480 10762
rect 16451 10750 16468 10756
rect 16414 10747 16466 10750
rect 16414 10740 16454 10747
rect 4664 10706 4724 10716
rect 4664 10616 4688 10706
rect 8774 10468 8802 10532
rect 8924 10480 9278 10630
rect 9522 10556 9584 10584
rect 10388 10544 10446 10572
rect 9226 10462 9278 10480
rect 10052 10412 10088 10480
rect 10180 10414 10280 10426
rect 10020 10402 10088 10412
rect 10052 10394 10088 10402
rect 10052 10367 10242 10394
rect 10244 10367 10552 10394
rect 8774 10118 8802 10182
rect 8924 10144 9278 10280
rect 8972 10130 9020 10144
rect 8746 10090 8798 10114
rect 9226 10112 9278 10144
rect 9480 10268 9532 10364
rect 9580 10326 9636 10338
rect 10052 10330 10552 10367
rect 10052 10326 10242 10330
rect 10244 10326 10552 10330
rect 10021 10311 10088 10326
rect 10036 10300 10088 10311
rect 10165 10300 10242 10326
rect 10280 10322 10313 10326
rect 9978 10296 10098 10300
rect 10165 10299 10278 10300
rect 10174 10298 10278 10299
rect 9976 10290 10098 10296
rect 10172 10290 10278 10298
rect 9966 10288 10278 10290
rect 9966 10282 10290 10288
rect 10312 10282 10313 10322
rect 10322 10282 10374 10312
rect 10438 10282 10470 10326
rect 10476 10304 10536 10326
rect 10472 10288 10526 10304
rect 10472 10282 10518 10288
rect 9966 10274 10299 10282
rect 9480 10046 9834 10268
rect 9966 10264 10088 10274
rect 10002 10258 10088 10264
rect 10094 10272 10299 10274
rect 10094 10258 10178 10272
rect 10222 10267 10299 10272
rect 10312 10270 10518 10282
rect 10222 10266 10290 10267
rect 10312 10266 10484 10270
rect 10206 10258 10484 10266
rect 10002 10256 10484 10258
rect 10000 10255 10484 10256
rect 10540 10255 10552 10326
rect 10000 10254 10552 10255
rect 10000 10250 10318 10254
rect 10000 10246 10332 10250
rect 10000 10242 10008 10246
rect 9988 10230 10008 10242
rect 10052 10218 10158 10246
rect 10172 10236 10178 10246
rect 10194 10234 10332 10246
rect 9962 10182 10018 10196
rect 10052 10182 10154 10218
rect 10232 10214 10332 10234
rect 10422 10236 10484 10254
rect 10422 10226 10476 10236
rect 10492 10218 10538 10236
rect 10182 10182 10382 10214
rect 10520 10190 10566 10208
rect 10052 10164 10232 10182
rect 10332 10164 10388 10182
rect 10052 10125 10196 10164
rect 10373 10149 10456 10164
rect 10052 10124 10232 10125
rect 10388 10124 10456 10149
rect 10052 10112 10456 10124
rect 9962 10098 10018 10112
rect 10052 10080 10088 10112
rect 10170 10110 10456 10112
rect 10232 10098 10332 10110
rect 9994 10066 10088 10080
rect 10052 10062 10088 10066
rect 10124 10064 10142 10066
rect 10180 10064 10280 10076
rect 10020 10052 10088 10062
rect 10118 10060 10180 10064
rect 10052 10044 10088 10052
rect 10116 10049 10180 10060
rect 10280 10056 10442 10064
rect 10280 10055 10343 10056
rect 10280 10051 10342 10055
rect 10116 10044 10178 10049
rect 9528 10018 9576 10032
rect 10052 10017 10242 10044
rect 10244 10017 10552 10044
rect 8794 9800 8802 9832
rect 8924 9794 9278 9930
rect 8972 9780 9020 9794
rect 8780 9768 8794 9772
rect 9226 9762 9278 9794
rect 9480 9918 9532 10014
rect 9580 9976 9636 9988
rect 10052 9980 10552 10017
rect 10052 9976 10242 9980
rect 10244 9976 10552 9980
rect 10021 9961 10088 9976
rect 10036 9950 10088 9961
rect 10165 9950 10242 9976
rect 10280 9972 10313 9976
rect 9978 9946 10098 9950
rect 10165 9949 10278 9950
rect 10174 9948 10278 9949
rect 9976 9940 10098 9946
rect 10172 9940 10278 9948
rect 9966 9938 10278 9940
rect 9966 9932 10290 9938
rect 10312 9932 10313 9972
rect 10322 9932 10374 9962
rect 10438 9932 10470 9976
rect 10476 9954 10536 9976
rect 10472 9938 10526 9954
rect 10472 9932 10518 9938
rect 9966 9924 10299 9932
rect 8780 9740 8782 9744
rect 9480 9696 9834 9918
rect 9966 9914 10088 9924
rect 10002 9908 10088 9914
rect 10094 9922 10299 9924
rect 10094 9908 10178 9922
rect 10222 9917 10299 9922
rect 10312 9920 10518 9932
rect 10222 9916 10290 9917
rect 10312 9916 10484 9920
rect 10206 9908 10484 9916
rect 10002 9906 10484 9908
rect 10000 9905 10484 9906
rect 10540 9905 10552 9976
rect 10000 9904 10552 9905
rect 10000 9900 10318 9904
rect 10000 9896 10332 9900
rect 10000 9892 10008 9896
rect 9988 9880 10008 9892
rect 10052 9868 10158 9896
rect 10172 9886 10178 9896
rect 10194 9884 10332 9896
rect 9962 9832 10018 9846
rect 10052 9832 10154 9868
rect 10232 9864 10332 9884
rect 10422 9886 10484 9904
rect 10422 9876 10476 9886
rect 10492 9868 10538 9886
rect 10182 9832 10382 9864
rect 10520 9840 10566 9858
rect 10052 9814 10232 9832
rect 10332 9814 10388 9832
rect 10052 9775 10196 9814
rect 10373 9799 10456 9814
rect 10052 9774 10232 9775
rect 10388 9774 10456 9799
rect 10052 9762 10456 9774
rect 9962 9748 10018 9762
rect 10052 9730 10088 9762
rect 10170 9760 10456 9762
rect 10232 9748 10332 9760
rect 9994 9716 10088 9730
rect 10052 9712 10088 9716
rect 10124 9714 10142 9716
rect 10180 9714 10280 9726
rect 10020 9702 10088 9712
rect 10118 9710 10180 9714
rect 10052 9694 10088 9702
rect 10116 9699 10180 9710
rect 10280 9706 10442 9714
rect 10280 9705 10343 9706
rect 10280 9701 10342 9705
rect 10116 9694 10178 9699
rect 11900 9698 11928 10740
rect 16412 10736 16454 10740
rect 16486 10736 16488 10804
rect 16512 10762 16526 10810
rect 16540 10762 16554 10810
rect 16752 10804 16858 10826
rect 17286 10818 17314 10854
rect 17780 10852 17800 10854
rect 17840 10848 17860 10858
rect 17754 10820 17756 10846
rect 17754 10818 17782 10820
rect 16768 10776 16830 10798
rect 16512 10756 16612 10762
rect 16414 10724 16454 10736
rect 16412 10722 16454 10724
rect 12840 10672 12878 10700
rect 13102 10686 13146 10698
rect 16398 10678 16466 10722
rect 16512 10710 16526 10756
rect 16540 10738 16554 10756
rect 16595 10750 16612 10756
rect 16595 10747 16610 10750
rect 16726 10736 16762 10750
rect 16780 10736 16816 10750
rect 16726 10734 16830 10736
rect 16726 10724 16762 10734
rect 16768 10732 16830 10734
rect 16780 10724 16816 10732
rect 17360 10728 17390 10746
rect 17448 10738 17478 10746
rect 16724 10722 16762 10724
rect 16778 10722 16816 10724
rect 16568 10690 16610 10722
rect 16712 10716 16816 10722
rect 17438 10718 17478 10738
rect 19438 10734 19522 10888
rect 22876 10874 23076 10888
rect 22934 10866 23014 10874
rect 23228 10868 23460 10888
rect 23624 10884 23858 10896
rect 22232 10852 22248 10864
rect 22882 10844 23142 10866
rect 23168 10864 23460 10868
rect 23158 10844 23460 10864
rect 23596 10872 23858 10884
rect 23596 10856 23898 10872
rect 23612 10846 23898 10856
rect 23648 10844 23662 10846
rect 23674 10844 23898 10846
rect 22718 10806 22724 10822
rect 22746 10794 22752 10822
rect 22882 10818 23460 10844
rect 22882 10810 23144 10818
rect 22854 10754 22866 10810
rect 22876 10778 22882 10810
rect 22888 10788 22900 10810
rect 22888 10780 22908 10788
rect 22888 10778 22912 10780
rect 22958 10778 22966 10810
rect 22986 10806 22994 10810
rect 23074 10796 23144 10810
rect 22872 10776 22912 10778
rect 22872 10772 22916 10776
rect 22872 10764 22922 10772
rect 22872 10762 22934 10764
rect 23010 10762 23020 10772
rect 22854 10746 22874 10754
rect 22876 10746 22882 10762
rect 22888 10758 22964 10762
rect 22888 10752 22922 10758
rect 22888 10746 22904 10752
rect 23026 10746 23042 10762
rect 22854 10742 22882 10746
rect 23074 10745 23142 10796
rect 22854 10740 22884 10742
rect 23014 10741 23142 10745
rect 23168 10741 23460 10818
rect 23564 10812 23570 10832
rect 23624 10812 23898 10844
rect 23968 10834 24084 10948
rect 23948 10818 24084 10834
rect 24128 10947 24279 10954
rect 24128 10916 24204 10947
rect 24214 10926 24268 10947
rect 24222 10916 24268 10926
rect 24128 10904 24268 10916
rect 24128 10900 24350 10904
rect 24128 10824 24190 10900
rect 24192 10878 24350 10900
rect 24192 10846 24248 10878
rect 24194 10832 24204 10846
rect 23528 10778 23548 10812
rect 23560 10810 23592 10812
rect 23560 10804 23598 10810
rect 23624 10804 23872 10812
rect 23560 10784 23872 10804
rect 23986 10790 24030 10818
rect 24086 10790 24136 10804
rect 24192 10790 24204 10832
rect 24222 10804 24232 10846
rect 24294 10842 24350 10878
rect 24220 10794 24268 10804
rect 24220 10790 24280 10794
rect 23986 10784 24136 10790
rect 23560 10778 23736 10784
rect 23790 10778 23872 10784
rect 23980 10778 24136 10784
rect 23560 10762 23626 10778
rect 23560 10746 23592 10762
rect 23594 10752 23626 10762
rect 23650 10760 23660 10778
rect 23650 10752 23658 10760
rect 23674 10758 23694 10778
rect 23706 10758 23724 10778
rect 23740 10766 23758 10776
rect 23790 10774 23898 10778
rect 23852 10766 23920 10774
rect 23986 10770 24136 10778
rect 24180 10776 24280 10790
rect 23980 10768 24136 10770
rect 23674 10751 23728 10758
rect 23736 10751 23920 10766
rect 23986 10762 24136 10768
rect 24178 10762 24280 10776
rect 23014 10740 23460 10741
rect 22854 10738 23460 10740
rect 19522 10720 19606 10734
rect 22854 10728 22900 10738
rect 22934 10736 23014 10738
rect 23128 10736 23460 10738
rect 23674 10738 23920 10751
rect 23968 10752 24348 10762
rect 23968 10750 24024 10752
rect 24034 10750 24036 10752
rect 24178 10750 24180 10752
rect 23932 10744 24038 10750
rect 23932 10738 24024 10744
rect 24192 10738 24204 10752
rect 23674 10736 24068 10738
rect 22934 10730 23026 10736
rect 16712 10708 16814 10716
rect 17438 10710 17476 10718
rect 20686 10708 20834 10720
rect 22854 10718 22930 10728
rect 22934 10726 23014 10730
rect 23168 10720 23460 10736
rect 23694 10728 23728 10736
rect 16712 10704 16828 10708
rect 22840 10704 22888 10706
rect 16712 10690 16814 10704
rect 22866 10694 22888 10704
rect 23168 10700 23456 10720
rect 23736 10711 23898 10736
rect 23918 10734 24068 10736
rect 23918 10732 24024 10734
rect 23932 10724 24024 10732
rect 23736 10710 23801 10711
rect 23814 10710 23898 10711
rect 23922 10722 24024 10724
rect 23922 10710 24034 10722
rect 23740 10708 23812 10710
rect 16566 10678 16610 10690
rect 16710 10678 16778 10690
rect 20714 10680 20806 10692
rect 22812 10670 22854 10672
rect 22934 10670 22950 10694
rect 22996 10686 23076 10696
rect 16742 10668 16766 10670
rect 16396 10660 16766 10668
rect 16396 10624 16566 10660
rect 16568 10652 16766 10660
rect 16568 10630 16760 10652
rect 16568 10624 16618 10630
rect 16478 10616 16524 10624
rect 16612 10616 16618 10624
rect 16716 10616 16760 10630
rect 21126 10626 21932 10650
rect 21976 10642 22188 10650
rect 21976 10626 22030 10642
rect 22220 10628 22248 10668
rect 22832 10660 22854 10670
rect 22866 10638 22880 10640
rect 22800 10628 22880 10638
rect 22894 10628 22908 10666
rect 22938 10628 22953 10643
rect 22996 10628 23076 10636
rect 23117 10628 23132 10643
rect 23168 10628 23322 10698
rect 23646 10678 23724 10686
rect 23750 10678 23812 10708
rect 23814 10706 24040 10710
rect 23814 10704 24034 10706
rect 23814 10678 23898 10704
rect 23646 10674 23736 10678
rect 23750 10674 23898 10678
rect 23596 10650 23602 10670
rect 23646 10666 23724 10674
rect 23646 10664 23726 10666
rect 23646 10642 23670 10664
rect 23674 10662 23704 10664
rect 23790 10662 23898 10674
rect 23922 10678 24034 10704
rect 24136 10690 24178 10722
rect 24220 10710 24232 10752
rect 24294 10724 24334 10750
rect 24292 10722 24334 10724
rect 24134 10678 24178 10690
rect 23674 10642 23736 10662
rect 23790 10642 23872 10662
rect 23922 10648 23974 10678
rect 23978 10668 24002 10670
rect 24258 10668 24260 10704
rect 24280 10690 24348 10722
rect 24278 10678 24346 10690
rect 24286 10668 24288 10676
rect 24332 10668 24334 10670
rect 23978 10664 24348 10668
rect 23978 10650 24134 10664
rect 23612 10640 23724 10642
rect 23728 10640 23872 10642
rect 12488 10596 12588 10606
rect 12848 10596 12948 10608
rect 13128 10596 13228 10606
rect 16396 10598 16524 10616
rect 13398 10560 14022 10580
rect 16412 10562 16524 10598
rect 12736 10524 12746 10538
rect 12488 10512 12588 10522
rect 12848 10512 12948 10524
rect 13128 10512 13228 10522
rect 12342 10468 12348 10470
rect 12324 10446 12348 10468
rect 12438 10462 12488 10502
rect 12432 10452 12488 10462
rect 12588 10462 12638 10502
rect 13078 10462 13128 10502
rect 12588 10452 12644 10462
rect 12432 10448 12447 10452
rect 12312 10434 12348 10446
rect 12418 10446 12447 10448
rect 12629 10446 12644 10452
rect 13068 10452 13128 10462
rect 13068 10446 13083 10452
rect 12356 10436 12376 10442
rect 12282 10420 12350 10434
rect 12356 10430 12398 10436
rect 12312 10406 12346 10420
rect 12282 10392 12350 10406
rect 12356 10396 12380 10430
rect 12384 10396 12398 10430
rect 12418 10414 12492 10446
rect 12584 10414 13134 10446
rect 13240 10416 13274 10444
rect 13320 10418 13354 10446
rect 13398 10416 13854 10560
rect 13410 10412 13854 10416
rect 12312 10380 12348 10392
rect 12356 10390 12398 10396
rect 12356 10384 12376 10390
rect 12324 10358 12348 10380
rect 12418 10380 12492 10412
rect 12584 10380 13134 10412
rect 13320 10380 13354 10408
rect 12418 10378 12447 10380
rect 12432 10374 12447 10378
rect 12629 10374 12644 10380
rect 12432 10364 12488 10374
rect 12342 10356 12348 10358
rect 12438 10324 12488 10364
rect 12588 10364 12644 10374
rect 13068 10374 13083 10380
rect 13068 10364 13128 10374
rect 13856 10372 14022 10560
rect 16478 10548 16524 10562
rect 16398 10534 16454 10548
rect 16396 10466 16454 10516
rect 16556 10466 16618 10616
rect 16714 10576 16760 10616
rect 21154 10598 21932 10622
rect 21976 10614 22258 10622
rect 21976 10598 22058 10614
rect 22192 10600 22258 10614
rect 22800 10606 23322 10628
rect 23646 10630 23670 10640
rect 23646 10624 23668 10630
rect 23602 10622 23668 10624
rect 23674 10628 23736 10640
rect 23790 10628 23852 10640
rect 23984 10630 24134 10650
rect 23602 10620 23664 10622
rect 23674 10620 23724 10628
rect 23602 10616 23724 10620
rect 23602 10614 23728 10616
rect 22804 10602 23322 10606
rect 22804 10598 22996 10602
rect 21154 10586 21774 10598
rect 21898 10586 21932 10592
rect 22192 10586 22258 10594
rect 22816 10578 22880 10598
rect 16716 10486 16760 10576
rect 21696 10572 21740 10574
rect 19102 10484 19106 10504
rect 16556 10448 16654 10466
rect 19136 10454 19140 10484
rect 19172 10478 19174 10542
rect 19200 10450 19202 10570
rect 21126 10558 21746 10572
rect 21926 10558 21932 10564
rect 22220 10526 22248 10566
rect 22828 10560 22880 10578
rect 22866 10554 22880 10560
rect 22894 10558 22908 10598
rect 22946 10592 22996 10598
rect 23076 10598 23322 10602
rect 23624 10612 23724 10614
rect 23802 10613 23920 10628
rect 23984 10616 24028 10630
rect 24126 10624 24134 10630
rect 24136 10624 24278 10664
rect 24280 10624 24348 10664
rect 24126 10616 24132 10624
rect 24220 10616 24266 10624
rect 24286 10616 24288 10624
rect 23624 10598 23674 10612
rect 23684 10606 23724 10612
rect 23684 10604 23712 10606
rect 23684 10598 23724 10604
rect 23076 10592 23126 10598
rect 22946 10588 23126 10592
rect 23168 10588 23322 10598
rect 23612 10596 23728 10598
rect 22946 10586 23322 10588
rect 23602 10586 23728 10596
rect 22934 10582 23322 10586
rect 22934 10580 22996 10582
rect 22938 10566 22996 10580
rect 23076 10566 23322 10582
rect 23612 10572 23728 10586
rect 22894 10534 22916 10558
rect 22938 10551 22953 10566
rect 23117 10551 23132 10566
rect 22832 10524 22854 10534
rect 22894 10528 22908 10534
rect 22812 10522 22854 10524
rect 22882 10502 23142 10524
rect 23168 10502 23322 10566
rect 23596 10552 23602 10572
rect 23612 10570 23712 10572
rect 23724 10570 23728 10572
rect 23650 10568 23670 10570
rect 23684 10568 23724 10570
rect 23736 10568 23770 10612
rect 23802 10606 23842 10613
rect 23802 10570 23842 10604
rect 23852 10570 23920 10613
rect 23966 10582 24030 10616
rect 23956 10576 24030 10582
rect 23624 10544 23674 10568
rect 23684 10556 23712 10568
rect 23684 10544 23704 10556
rect 23624 10536 23726 10544
rect 23790 10542 23852 10570
rect 23872 10542 23898 10570
rect 23956 10548 24028 10576
rect 23736 10536 23920 10542
rect 23624 10528 23920 10536
rect 23624 10520 23684 10528
rect 23724 10520 23920 10528
rect 23624 10518 23920 10520
rect 22882 10500 23322 10502
rect 23646 10500 23724 10518
rect 23736 10510 23920 10518
rect 23750 10502 23920 10510
rect 23740 10500 23920 10502
rect 22866 10496 23362 10500
rect 22866 10490 23142 10496
rect 22840 10488 23142 10490
rect 22882 10484 23142 10488
rect 22882 10480 23200 10484
rect 22770 10472 23228 10480
rect 23674 10474 23702 10492
rect 23736 10474 23920 10500
rect 22770 10468 23362 10472
rect 16454 10404 16544 10448
rect 16454 10388 16532 10404
rect 16556 10388 16572 10448
rect 22770 10446 23228 10468
rect 23282 10456 23362 10468
rect 23560 10448 23592 10464
rect 23646 10458 23654 10466
rect 23674 10462 23736 10474
rect 23594 10448 23626 10458
rect 23236 10446 23252 10448
rect 22770 10442 23252 10446
rect 22770 10404 23236 10442
rect 23298 10432 23362 10446
rect 23402 10432 23456 10446
rect 23434 10420 23466 10430
rect 23298 10404 23362 10418
rect 23402 10404 23460 10418
rect 23560 10416 23626 10448
rect 23646 10450 23658 10458
rect 23646 10420 23660 10450
rect 23674 10448 23702 10462
rect 23674 10437 23694 10448
rect 23684 10420 23694 10437
rect 23706 10420 23724 10462
rect 23728 10459 23736 10462
rect 23740 10434 23758 10474
rect 23790 10473 23920 10474
rect 23802 10436 23842 10452
rect 23852 10436 23920 10473
rect 23966 10486 24028 10548
rect 23790 10434 23852 10436
rect 23750 10426 23858 10434
rect 23736 10420 23858 10426
rect 23650 10416 23660 10420
rect 23674 10416 23858 10420
rect 23560 10406 23858 10416
rect 16454 10380 16572 10388
rect 22192 10386 22260 10398
rect 22770 10386 23228 10404
rect 23560 10400 23598 10406
rect 23560 10398 23592 10400
rect 12588 10324 12638 10364
rect 13078 10324 13128 10364
rect 21018 10342 21208 10372
rect 12488 10304 12588 10314
rect 12848 10302 12948 10314
rect 13128 10304 13228 10314
rect 12734 10288 12746 10302
rect 13034 10278 13048 10296
rect 12488 10220 12588 10230
rect 12714 10164 13398 10278
rect 13860 10238 13896 10298
rect 13914 10238 13950 10294
rect 13638 10196 13666 10228
rect 13832 10226 13896 10238
rect 13914 10126 13956 10226
rect 16332 10182 16994 10306
rect 13832 10110 13896 10126
rect 16540 10110 16708 10182
rect 17480 10170 17544 10178
rect 17502 10142 17554 10150
rect 13860 10090 13896 10110
rect 13778 10058 13896 10090
rect 13914 10068 13950 10110
rect 13914 10060 14136 10068
rect 13778 10004 13896 10036
rect 12488 9956 12588 9966
rect 12848 9956 12948 9968
rect 13032 9936 13052 9946
rect 13060 9936 13080 9974
rect 13128 9956 13228 9966
rect 13860 9964 13896 10004
rect 13914 10006 14136 10014
rect 13914 9964 13950 10006
rect 13914 9958 13980 9964
rect 12930 9884 13008 9928
rect 13068 9890 13156 9928
rect 12488 9872 12588 9882
rect 12848 9872 12948 9884
rect 13032 9882 13052 9890
rect 13060 9882 13156 9890
rect 13060 9874 13080 9882
rect 12984 9862 13102 9874
rect 13128 9872 13228 9882
rect 12342 9828 12348 9830
rect 12324 9806 12348 9828
rect 12438 9822 12488 9862
rect 12432 9812 12488 9822
rect 12588 9822 12638 9862
rect 12588 9812 12644 9822
rect 12432 9808 12447 9812
rect 12312 9794 12348 9806
rect 12418 9806 12447 9808
rect 12629 9806 12644 9812
rect 12984 9812 13128 9862
rect 12984 9806 13036 9812
rect 13048 9808 13102 9812
rect 13068 9806 13106 9808
rect 12356 9796 12376 9802
rect 12282 9780 12350 9794
rect 12356 9790 12398 9796
rect 12312 9766 12346 9780
rect 12282 9752 12350 9766
rect 12356 9756 12380 9790
rect 12384 9756 12398 9790
rect 12418 9774 12492 9806
rect 12584 9790 13036 9806
rect 12584 9782 13016 9790
rect 13048 9782 13116 9806
rect 12584 9774 13116 9782
rect 13126 9774 13134 9806
rect 13240 9776 13274 9804
rect 13320 9778 13354 9806
rect 13398 9774 13664 9940
rect 13914 9888 13956 9958
rect 18076 9948 18472 10114
rect 18076 9946 18344 9948
rect 13832 9880 13908 9888
rect 13778 9864 13908 9880
rect 13832 9830 13908 9864
rect 13734 9774 13746 9800
rect 12984 9772 13102 9774
rect 12312 9740 12348 9752
rect 12356 9750 12398 9756
rect 12356 9744 12376 9750
rect 12324 9718 12348 9740
rect 12418 9740 12492 9772
rect 12584 9740 13058 9772
rect 12418 9738 12447 9740
rect 12432 9734 12447 9738
rect 12629 9734 12644 9740
rect 12432 9724 12488 9734
rect 12342 9716 12348 9718
rect 9528 9668 9576 9682
rect 10052 9667 10242 9694
rect 10244 9667 10552 9694
rect 8774 9418 8802 9482
rect 8924 9444 9278 9580
rect 9226 9412 9278 9444
rect 9480 9568 9532 9664
rect 9580 9626 9636 9638
rect 10052 9630 10552 9667
rect 10052 9626 10242 9630
rect 10244 9626 10552 9630
rect 10021 9611 10088 9626
rect 10036 9600 10088 9611
rect 10165 9600 10242 9626
rect 10280 9622 10313 9626
rect 9978 9596 10098 9600
rect 10165 9599 10278 9600
rect 10174 9598 10278 9599
rect 9976 9590 10098 9596
rect 10172 9590 10278 9598
rect 9966 9588 10278 9590
rect 9966 9582 10290 9588
rect 10312 9582 10313 9622
rect 10322 9582 10374 9612
rect 10438 9582 10470 9626
rect 10476 9604 10536 9626
rect 10472 9588 10526 9604
rect 10472 9582 10518 9588
rect 9966 9574 10299 9582
rect 9480 9346 9834 9568
rect 9966 9564 10088 9574
rect 10002 9558 10088 9564
rect 10094 9572 10299 9574
rect 10094 9558 10178 9572
rect 10222 9567 10299 9572
rect 10312 9570 10518 9582
rect 10222 9566 10290 9567
rect 10312 9566 10484 9570
rect 10206 9558 10484 9566
rect 10002 9556 10484 9558
rect 10000 9555 10484 9556
rect 10540 9555 10552 9626
rect 10000 9554 10552 9555
rect 10000 9550 10318 9554
rect 10000 9546 10332 9550
rect 10000 9542 10008 9546
rect 9988 9530 10008 9542
rect 10052 9518 10158 9546
rect 10172 9536 10178 9546
rect 10194 9534 10332 9546
rect 9962 9482 10018 9496
rect 10052 9482 10154 9518
rect 10232 9514 10332 9534
rect 10422 9536 10484 9554
rect 10422 9526 10476 9536
rect 10492 9518 10538 9536
rect 10182 9482 10382 9514
rect 10520 9490 10566 9508
rect 11900 9490 11930 9698
rect 12438 9684 12488 9724
rect 12588 9724 12644 9734
rect 12984 9734 13058 9740
rect 13068 9762 13106 9772
rect 13068 9734 13102 9762
rect 13126 9740 13134 9772
rect 13320 9740 13354 9768
rect 13860 9740 13908 9830
rect 13914 9830 13928 9880
rect 13914 9780 13962 9830
rect 12984 9726 13128 9734
rect 13068 9724 13128 9726
rect 12588 9684 12638 9724
rect 13078 9692 13128 9724
rect 13060 9684 13128 9692
rect 12488 9664 12588 9674
rect 12848 9662 12948 9674
rect 12734 9648 12746 9662
rect 13032 9656 13052 9664
rect 13060 9656 13080 9684
rect 13128 9664 13228 9674
rect 12488 9580 12588 9590
rect 12848 9578 12948 9590
rect 13128 9580 13228 9590
rect 13860 9588 13896 9658
rect 14066 9656 14248 9910
rect 18076 9848 18090 9946
rect 18096 9866 18100 9946
rect 18124 9894 18128 9946
rect 18160 9938 18180 9946
rect 18188 9938 18208 9946
rect 18578 9918 18592 9998
rect 18606 9946 18652 9974
rect 19294 9958 19538 10342
rect 20922 10238 20958 10294
rect 20976 10238 21012 10298
rect 21018 10276 21450 10342
rect 22220 10330 22248 10370
rect 22752 10360 23228 10386
rect 23282 10372 23362 10384
rect 23564 10378 23570 10398
rect 23624 10396 23858 10406
rect 23872 10396 23898 10436
rect 23624 10394 23906 10396
rect 23612 10366 23906 10394
rect 23648 10364 23662 10366
rect 23674 10364 23906 10366
rect 22770 10358 23228 10360
rect 22752 10346 23228 10358
rect 23624 10356 23906 10364
rect 23966 10386 24024 10486
rect 24126 10466 24188 10616
rect 24242 10598 24348 10616
rect 24292 10562 24348 10598
rect 24220 10514 24266 10516
rect 24212 10466 24266 10514
rect 24290 10466 24348 10516
rect 24090 10448 24188 10466
rect 23966 10358 24084 10386
rect 24172 10380 24188 10448
rect 24200 10438 24290 10448
rect 24212 10404 24290 10438
rect 24212 10388 24282 10404
rect 22752 10332 23422 10346
rect 22770 10328 23422 10332
rect 23596 10328 23906 10356
rect 23962 10340 24084 10358
rect 22934 10320 23422 10328
rect 21746 10300 22188 10316
rect 22998 10312 23422 10320
rect 23624 10314 23906 10328
rect 22998 10294 23456 10312
rect 23648 10300 23662 10314
rect 23674 10296 23728 10300
rect 23750 10296 23906 10314
rect 20976 10226 21040 10238
rect 20976 10126 21018 10226
rect 20976 10110 21040 10126
rect 20922 10068 20958 10110
rect 20736 10060 20958 10068
rect 20976 10090 21012 10110
rect 20976 10058 21094 10090
rect 21208 10042 21450 10276
rect 21746 10272 22216 10288
rect 22030 10252 22216 10266
rect 22030 10244 22260 10252
rect 21882 10218 21970 10226
rect 22030 10216 22188 10238
rect 22220 10216 22248 10224
rect 22232 10198 22248 10216
rect 21910 10190 21970 10198
rect 22590 10180 22608 10208
rect 22618 10186 22620 10252
rect 22876 10250 23456 10294
rect 23624 10274 23906 10296
rect 22934 10236 23456 10250
rect 23612 10246 23906 10274
rect 23966 10262 24084 10340
rect 24132 10263 24134 10328
rect 24132 10262 24149 10263
rect 23966 10256 24149 10262
rect 23620 10244 23906 10246
rect 22922 10196 22934 10226
rect 22950 10224 22962 10236
rect 22998 10226 23456 10236
rect 22964 10210 23028 10226
rect 23166 10224 23456 10226
rect 23158 10216 23456 10224
rect 23596 10236 23906 10244
rect 23948 10248 24149 10256
rect 23948 10240 24084 10248
rect 23596 10216 23950 10236
rect 24030 10222 24084 10240
rect 22936 10182 23056 10198
rect 23130 10156 23144 10196
rect 23158 10184 23186 10216
rect 23200 10208 23212 10216
rect 23228 10208 23456 10216
rect 23560 10210 23592 10212
rect 23624 10210 23950 10216
rect 23388 10178 23412 10208
rect 23416 10206 23440 10208
rect 23560 10206 23950 10210
rect 24069 10208 24084 10222
rect 23560 10194 23674 10206
rect 23560 10188 23662 10194
rect 23200 10170 23264 10178
rect 23560 10162 23626 10188
rect 23190 10142 23292 10150
rect 23560 10146 23592 10162
rect 23594 10152 23626 10162
rect 23650 10160 23660 10188
rect 23684 10173 23694 10204
rect 23650 10152 23658 10160
rect 23674 10158 23694 10173
rect 23706 10158 23724 10204
rect 23736 10184 23950 10206
rect 23750 10182 23950 10184
rect 24082 10182 24084 10184
rect 24162 10182 24412 10306
rect 23740 10166 23758 10176
rect 23790 10174 23852 10182
rect 23836 10166 23852 10174
rect 23674 10151 23728 10158
rect 23736 10151 23852 10166
rect 23428 10114 23452 10140
rect 23674 10136 23852 10151
rect 23906 10142 23920 10174
rect 23694 10128 23728 10136
rect 21756 10042 21806 10050
rect 22668 10042 22770 10114
rect 23736 10112 23790 10136
rect 19294 9946 19572 9958
rect 18730 9894 18776 9916
rect 19294 9894 19538 9946
rect 19732 9926 19752 10042
rect 19760 9974 19780 10014
rect 20736 10006 20958 10014
rect 19760 9954 19824 9974
rect 20922 9964 20958 10006
rect 20976 10004 21094 10036
rect 21180 10022 21984 10042
rect 21208 10014 21450 10022
rect 21756 10014 21757 10022
rect 21806 10014 21832 10022
rect 22230 10014 22248 10028
rect 20976 9964 21012 10004
rect 21180 9994 21984 10014
rect 22368 10002 22408 10030
rect 22646 10020 22770 10042
rect 22668 10014 22770 10020
rect 22876 10092 23166 10108
rect 22876 10072 23168 10092
rect 23190 10080 23200 10090
rect 23264 10080 23362 10090
rect 23456 10086 23480 10112
rect 23526 10080 23696 10112
rect 23736 10111 23852 10112
rect 23736 10110 23801 10111
rect 23740 10108 23778 10110
rect 23438 10074 23696 10080
rect 23724 10088 23778 10092
rect 23780 10090 23812 10110
rect 23780 10088 23848 10090
rect 23724 10078 23848 10088
rect 23724 10074 23872 10078
rect 22876 10062 23322 10072
rect 22876 10052 23362 10062
rect 23438 10052 23872 10074
rect 23904 10052 23950 10142
rect 24070 10080 24088 10182
rect 24104 10114 24131 10148
rect 24083 10066 24084 10080
rect 20892 9958 20958 9964
rect 21208 9960 21450 9994
rect 19770 9930 19816 9954
rect 19742 9902 19752 9926
rect 18124 9878 19618 9894
rect 19294 9866 19538 9878
rect 18096 9850 19590 9866
rect 18090 9812 18244 9848
rect 19090 9832 19208 9834
rect 19088 9822 19208 9832
rect 16467 9737 16543 9748
rect 16478 9720 16532 9737
rect 16478 9698 16524 9720
rect 16396 9672 16502 9698
rect 13914 9588 13950 9644
rect 14320 9600 14502 9656
rect 16412 9636 16502 9672
rect 16556 9618 16618 9748
rect 19088 9736 19114 9822
rect 19118 9804 19180 9806
rect 19116 9794 19180 9804
rect 19116 9764 19142 9794
rect 19172 9764 19180 9794
rect 19116 9740 19180 9764
rect 19142 9736 19172 9740
rect 19200 9736 19208 9822
rect 16716 9620 16760 9728
rect 19088 9712 19208 9736
rect 19294 9726 19538 9850
rect 17790 9664 17806 9678
rect 17746 9650 17806 9664
rect 17762 9646 17806 9650
rect 16716 9616 16850 9620
rect 16716 9600 16856 9616
rect 14320 9588 14554 9600
rect 14598 9588 14698 9600
rect 16478 9588 16524 9598
rect 13832 9586 13896 9588
rect 10052 9464 10232 9482
rect 10332 9464 10388 9482
rect 12840 9476 12878 9504
rect 13102 9476 13148 9504
rect 13734 9490 13746 9504
rect 13914 9486 13956 9586
rect 14320 9516 14502 9588
rect 16466 9584 16524 9588
rect 16610 9596 16660 9598
rect 16716 9596 16760 9600
rect 16466 9556 16566 9584
rect 16610 9556 16994 9596
rect 14696 9516 14756 9520
rect 14970 9518 15002 9546
rect 15052 9518 15090 9546
rect 15132 9520 15164 9548
rect 16398 9546 16994 9556
rect 14320 9504 14554 9516
rect 14598 9508 14756 9516
rect 16644 9512 16994 9546
rect 17438 9512 17476 9540
rect 14598 9504 14698 9508
rect 10052 9425 10196 9464
rect 10373 9449 10456 9464
rect 13832 9460 13896 9486
rect 14320 9474 14502 9504
rect 14724 9484 14784 9492
rect 14724 9480 14780 9484
rect 10052 9424 10232 9425
rect 10388 9424 10456 9449
rect 13860 9434 13896 9460
rect 10052 9412 10456 9424
rect 13778 9418 13896 9434
rect 13914 9420 13950 9460
rect 14066 9420 14248 9474
rect 9962 9398 10018 9412
rect 10052 9380 10088 9412
rect 10170 9410 10456 9412
rect 13914 9410 14248 9420
rect 10232 9398 10332 9410
rect 9994 9366 10088 9380
rect 10052 9362 10088 9366
rect 10124 9364 10142 9366
rect 10180 9364 10280 9376
rect 13778 9364 13896 9380
rect 14066 9366 14248 9410
rect 10020 9352 10088 9362
rect 10118 9360 10180 9364
rect 10052 9344 10088 9352
rect 10116 9349 10180 9360
rect 10280 9356 10442 9364
rect 10280 9355 10343 9356
rect 10280 9351 10342 9355
rect 10116 9344 10178 9349
rect 9528 9318 9562 9332
rect 10052 9317 10242 9344
rect 10244 9317 10552 9344
rect 8924 9094 9278 9248
rect 9480 9080 9532 9314
rect 9580 9276 9636 9288
rect 10052 9280 10552 9317
rect 13860 9310 13896 9364
rect 13914 9356 14248 9366
rect 13914 9310 13950 9356
rect 13832 9308 13896 9310
rect 10052 9276 10242 9280
rect 10244 9276 10552 9280
rect 10021 9261 10088 9276
rect 10036 9250 10088 9261
rect 10165 9250 10242 9276
rect 10280 9272 10313 9276
rect 9978 9246 10098 9250
rect 10165 9249 10278 9250
rect 10174 9248 10278 9249
rect 9976 9240 10098 9246
rect 10172 9240 10278 9248
rect 9966 9238 10278 9240
rect 9966 9232 10290 9238
rect 10312 9232 10313 9272
rect 10322 9232 10374 9262
rect 10438 9232 10470 9276
rect 10476 9254 10536 9276
rect 10472 9238 10526 9254
rect 10472 9232 10518 9238
rect 9966 9224 10299 9232
rect 9966 9214 10088 9224
rect 10002 9208 10088 9214
rect 10094 9222 10299 9224
rect 10094 9208 10178 9222
rect 10222 9217 10299 9222
rect 10312 9220 10518 9232
rect 10222 9216 10290 9217
rect 10312 9216 10484 9220
rect 10206 9208 10484 9216
rect 10002 9206 10484 9208
rect 10000 9205 10484 9206
rect 10540 9205 10552 9276
rect 13914 9208 13956 9308
rect 14066 9220 14248 9356
rect 14320 9458 14832 9474
rect 14320 9422 14842 9458
rect 14320 9274 14832 9422
rect 16426 9418 16994 9512
rect 15828 9336 16050 9392
rect 10000 9204 10552 9205
rect 9580 9192 9636 9204
rect 10000 9200 10318 9204
rect 10000 9196 10332 9200
rect 10422 9196 10484 9204
rect 10000 9192 10008 9196
rect 9988 9180 10008 9192
rect 10052 9168 10158 9196
rect 10172 9186 10178 9196
rect 10194 9184 10332 9196
rect 10388 9186 10484 9196
rect 9678 9132 9734 9144
rect 9962 9132 10018 9146
rect 10052 9132 10154 9168
rect 10232 9164 10332 9184
rect 10422 9176 10476 9186
rect 13832 9182 13896 9208
rect 10182 9132 10382 9164
rect 13860 9140 13896 9182
rect 13914 9132 13950 9182
rect 10052 9114 10232 9132
rect 10332 9114 10388 9132
rect 10052 9080 10154 9114
rect 10170 9080 10196 9114
rect 10373 9099 10456 9114
rect 10388 9080 10456 9099
rect 14320 9064 14502 9220
rect 14598 9116 14698 9128
rect 14798 9072 14832 9194
rect 15762 9158 16116 9336
rect 16680 9324 16798 9404
rect 16898 9342 16912 9418
rect 17960 9342 17974 9474
rect 18074 9342 18192 9404
rect 16614 9170 16864 9324
rect 16898 9306 17066 9342
rect 17960 9324 18192 9342
rect 18822 9336 19044 9392
rect 17960 9306 18258 9324
rect 18008 9170 18258 9306
rect 18756 9158 19110 9336
rect 19276 9296 19300 9602
rect 20174 9588 20274 9600
rect 20318 9588 20418 9600
rect 19304 9296 19328 9574
rect 19782 9518 19820 9546
rect 19870 9518 19902 9546
rect 20116 9516 20176 9520
rect 20116 9508 20274 9516
rect 20174 9504 20274 9508
rect 20318 9504 20418 9516
rect 20088 9484 20148 9492
rect 20092 9480 20148 9484
rect 19748 9420 19752 9448
rect 19798 9426 19810 9432
rect 19770 9420 19816 9426
rect 19764 9414 19822 9420
rect 19764 9408 19782 9414
rect 19776 9398 19782 9408
rect 19764 9390 19782 9398
rect 19804 9408 19822 9414
rect 19804 9398 19816 9408
rect 19804 9390 19822 9398
rect 19764 9386 19822 9390
rect 19748 9356 19752 9386
rect 19776 9384 19810 9386
rect 19798 9374 19810 9384
rect 19744 9216 19752 9354
rect 19772 9250 19780 9326
rect 20040 9274 20552 9474
rect 20624 9420 20806 9910
rect 20976 9888 21018 9958
rect 21176 9948 21450 9960
rect 21196 9932 21450 9948
rect 20964 9880 21040 9888
rect 20944 9830 20958 9880
rect 20910 9780 20958 9830
rect 20964 9864 21094 9880
rect 20964 9830 21040 9864
rect 20964 9740 21012 9830
rect 21208 9726 21450 9932
rect 21756 9715 21757 9994
rect 21806 9874 21832 9994
rect 22618 9992 22784 10014
rect 22876 10000 23322 10052
rect 23438 10034 23950 10052
rect 23998 10040 24009 10051
rect 24023 10040 24081 10051
rect 23962 10034 24009 10040
rect 23438 10026 24030 10034
rect 24034 10026 24081 10040
rect 22486 9960 22516 9972
rect 22476 9954 22516 9960
rect 22592 9954 22622 9972
rect 22476 9948 22478 9954
rect 22514 9944 22516 9954
rect 22566 9948 22578 9954
rect 22514 9916 22550 9940
rect 21968 9882 22014 9916
rect 22536 9876 22550 9916
rect 22564 9878 22578 9948
rect 22620 9944 22622 9954
rect 22668 9970 22770 9992
rect 22868 9984 23322 10000
rect 22876 9978 23322 9984
rect 22668 9958 22822 9970
rect 22866 9958 23322 9978
rect 23410 9972 23412 10014
rect 22668 9946 23322 9958
rect 22620 9916 22628 9938
rect 22770 9904 23322 9946
rect 21770 9726 21806 9874
rect 23086 9854 23110 9872
rect 23400 9868 23402 9894
rect 23406 9890 23412 9972
rect 23438 10006 24088 10026
rect 23438 9992 23961 10006
rect 24030 9992 24084 10006
rect 23438 9972 24090 9992
rect 23438 9952 23950 9972
rect 23964 9958 24084 9972
rect 23966 9952 24084 9958
rect 23438 9950 24084 9952
rect 24132 9971 24149 9986
rect 23438 9948 24082 9950
rect 23434 9930 24082 9948
rect 23434 9918 23694 9930
rect 23438 9912 23694 9918
rect 23722 9922 24082 9930
rect 23722 9918 23948 9922
rect 23966 9918 24082 9922
rect 23722 9912 24090 9918
rect 23596 9904 23634 9912
rect 23456 9886 23488 9894
rect 23646 9888 23662 9912
rect 23734 9904 23918 9912
rect 23750 9896 23918 9904
rect 23738 9894 23918 9896
rect 23562 9886 23680 9888
rect 23646 9876 23662 9886
rect 23734 9868 23918 9894
rect 23946 9902 24090 9912
rect 24132 9902 24134 9971
rect 23946 9888 24086 9902
rect 24146 9894 24188 9931
rect 23962 9884 24086 9888
rect 24132 9884 24188 9894
rect 23966 9872 24086 9884
rect 23400 9858 23460 9866
rect 23590 9858 23652 9860
rect 23130 9844 23142 9854
rect 22670 9800 22760 9826
rect 22888 9802 22904 9808
rect 22922 9802 22930 9820
rect 22934 9816 23014 9828
rect 23130 9818 23200 9844
rect 23400 9840 23430 9858
rect 23558 9842 23590 9858
rect 23672 9856 23734 9868
rect 23592 9842 23624 9852
rect 21806 9715 21832 9726
rect 21756 9714 21832 9715
rect 22402 9704 22774 9800
rect 23026 9792 23042 9808
rect 22872 9776 22888 9792
rect 23010 9782 23020 9792
rect 22958 9744 22966 9776
rect 22996 9748 23006 9758
rect 23130 9748 23142 9818
rect 23170 9816 23200 9818
rect 23282 9816 23362 9828
rect 22986 9744 22994 9748
rect 22934 9732 23014 9744
rect 23130 9737 23144 9748
rect 23174 9737 23200 9816
rect 23224 9792 23228 9816
rect 23558 9810 23624 9842
rect 23648 9844 23656 9852
rect 23648 9810 23658 9844
rect 23672 9831 23692 9856
rect 23682 9814 23692 9831
rect 23704 9814 23722 9856
rect 23726 9853 23734 9856
rect 23738 9828 23756 9868
rect 23788 9867 23918 9868
rect 23800 9830 23840 9846
rect 23850 9830 23918 9867
rect 23946 9848 24086 9872
rect 24106 9874 24188 9884
rect 24106 9868 24172 9874
rect 24106 9850 24120 9868
rect 24122 9850 24172 9868
rect 23946 9842 23962 9848
rect 23966 9842 24086 9848
rect 23788 9828 23850 9830
rect 23750 9820 23856 9828
rect 23734 9814 23856 9820
rect 23672 9810 23856 9814
rect 23236 9802 23252 9808
rect 23558 9800 23856 9810
rect 23558 9794 23596 9800
rect 23558 9792 23590 9794
rect 23220 9776 23236 9792
rect 23434 9780 23466 9790
rect 23224 9744 23228 9776
rect 23562 9772 23568 9792
rect 23622 9788 23856 9800
rect 23610 9760 23856 9788
rect 23672 9759 23856 9760
rect 23870 9759 23896 9830
rect 23946 9816 24086 9842
rect 24132 9840 24172 9850
rect 23946 9790 24082 9816
rect 23966 9774 24082 9790
rect 23672 9758 23896 9759
rect 23130 9736 23200 9737
rect 22986 9710 22994 9732
rect 21978 9660 22188 9674
rect 22402 9658 22838 9704
rect 22934 9680 23014 9694
rect 23130 9686 23144 9736
rect 23282 9732 23362 9744
rect 23622 9708 23776 9758
rect 23962 9742 24082 9774
rect 23672 9690 23726 9694
rect 23750 9690 23856 9708
rect 23622 9668 23856 9690
rect 23610 9666 23856 9668
rect 20922 9588 20958 9644
rect 20976 9588 21012 9658
rect 22402 9646 22774 9658
rect 21950 9632 22216 9646
rect 22558 9630 22632 9646
rect 22640 9630 22788 9646
rect 23068 9632 23082 9666
rect 23106 9658 23118 9666
rect 22606 9626 22630 9630
rect 22640 9626 22696 9630
rect 22640 9612 22664 9626
rect 22674 9620 22696 9626
rect 22614 9598 22630 9612
rect 20976 9586 21040 9588
rect 20976 9486 21018 9586
rect 22586 9574 22604 9596
rect 22640 9592 22648 9612
rect 22702 9592 22724 9630
rect 23028 9614 23082 9616
rect 22934 9596 23014 9610
rect 23028 9596 23086 9614
rect 23102 9612 23116 9658
rect 23610 9640 23896 9666
rect 23672 9638 23896 9640
rect 23622 9636 23813 9638
rect 23814 9636 23896 9638
rect 23388 9610 23412 9626
rect 23416 9610 23440 9626
rect 23028 9588 23042 9596
rect 23028 9586 23054 9588
rect 23028 9568 23058 9586
rect 23228 9568 23456 9610
rect 23562 9606 23568 9626
rect 23622 9606 23896 9636
rect 23966 9628 24082 9742
rect 23946 9612 24082 9628
rect 24126 9618 24188 9748
rect 24201 9737 24277 9748
rect 24212 9720 24266 9737
rect 24220 9698 24266 9720
rect 24242 9672 24348 9698
rect 24292 9636 24348 9672
rect 23526 9572 23546 9606
rect 23558 9604 23590 9606
rect 23558 9598 23596 9604
rect 23622 9598 23870 9606
rect 23558 9578 23870 9598
rect 23984 9584 24028 9612
rect 24084 9584 24134 9598
rect 24220 9588 24266 9598
rect 24220 9584 24278 9588
rect 23984 9578 24134 9584
rect 23558 9572 23734 9578
rect 23788 9572 23870 9578
rect 23978 9572 24134 9578
rect 22702 9542 22744 9564
rect 22718 9522 22764 9536
rect 22694 9514 22764 9522
rect 22694 9506 22744 9514
rect 23268 9512 23306 9540
rect 23388 9538 23412 9568
rect 23416 9566 23440 9568
rect 23558 9556 23624 9572
rect 23558 9540 23590 9556
rect 23592 9546 23624 9556
rect 23648 9554 23658 9572
rect 23648 9546 23656 9554
rect 23672 9552 23692 9572
rect 23704 9552 23722 9572
rect 23738 9560 23756 9570
rect 23788 9568 23896 9572
rect 23850 9560 23918 9568
rect 23984 9564 24134 9572
rect 23978 9562 24134 9564
rect 23672 9545 23726 9552
rect 23734 9545 23918 9560
rect 23984 9556 24134 9562
rect 24178 9556 24278 9584
rect 23672 9532 23918 9545
rect 23966 9546 24346 9556
rect 23966 9544 24022 9546
rect 23930 9538 24036 9544
rect 23930 9532 24022 9538
rect 23672 9530 24066 9532
rect 23692 9522 23726 9530
rect 23734 9506 23896 9530
rect 23916 9528 24066 9530
rect 23916 9526 24022 9528
rect 23930 9510 24022 9526
rect 22718 9490 22724 9506
rect 23734 9505 23850 9506
rect 23734 9504 23799 9505
rect 23870 9504 23896 9506
rect 23956 9504 24022 9510
rect 23738 9502 23810 9504
rect 20976 9460 21040 9486
rect 22718 9478 22764 9490
rect 23750 9486 23810 9502
rect 23622 9480 23682 9486
rect 23722 9484 23810 9486
rect 23870 9498 23942 9504
rect 23956 9500 24038 9504
rect 23722 9480 23846 9484
rect 23622 9472 23846 9480
rect 23870 9472 23896 9498
rect 23956 9486 24022 9500
rect 23966 9484 24022 9486
rect 23622 9468 24412 9472
rect 23622 9464 23722 9468
rect 20922 9420 20958 9460
rect 20624 9410 20958 9420
rect 20976 9434 21012 9460
rect 23610 9458 23726 9464
rect 23610 9436 23702 9458
rect 23722 9436 23726 9458
rect 23644 9434 23668 9436
rect 23672 9434 23722 9436
rect 23734 9434 24412 9468
rect 20976 9418 21094 9434
rect 23622 9432 23702 9434
rect 23622 9418 23722 9432
rect 23750 9418 24412 9434
rect 23600 9410 23722 9418
rect 20624 9366 20806 9410
rect 23600 9408 23726 9410
rect 23622 9406 23722 9408
rect 23622 9392 23672 9406
rect 23682 9400 23722 9406
rect 23682 9392 23722 9398
rect 23610 9390 23726 9392
rect 23600 9380 23726 9390
rect 20624 9356 20958 9366
rect 19772 9248 19784 9250
rect 19806 9248 19812 9250
rect 19772 9244 19812 9248
rect 19820 9244 19844 9266
rect 19778 9242 19844 9244
rect 19778 9232 19790 9242
rect 19800 9236 19844 9242
rect 19800 9230 19812 9236
rect 19816 9232 19844 9236
rect 9678 9048 9734 9060
rect 9962 9048 10018 9062
rect 10232 9048 10332 9060
rect 14598 9032 14698 9044
rect 14798 9036 14842 9072
rect 14724 9010 14780 9014
rect 14724 9002 14784 9010
rect 14696 8974 14756 8986
rect 14728 8948 14780 8952
rect 14400 8932 14440 8948
rect 14696 8932 14780 8948
rect 14798 8940 14832 9036
rect 14886 8940 15256 9106
rect 14886 8938 15086 8940
rect 15088 8938 15256 8940
rect 14292 8900 14724 8924
rect 14696 8898 14718 8900
rect 14320 8872 14724 8896
rect 14728 8894 14780 8932
rect 15018 8928 15256 8938
rect 15018 8876 15042 8928
rect 15046 8906 15256 8928
rect 15046 8904 15070 8906
rect 15046 8900 15094 8904
rect 15052 8892 15080 8900
rect 15106 8896 15132 8906
rect 18076 8902 18092 9006
rect 15106 8890 15122 8896
rect 18048 8888 18116 8902
rect 15018 8872 15122 8876
rect 18076 8874 18092 8888
rect 14696 8860 14756 8872
rect 15024 8864 15102 8872
rect 14724 8836 14784 8844
rect 18076 8838 18244 8874
rect 14724 8832 14780 8836
rect 14320 8810 14832 8828
rect 18048 8810 18120 8836
rect 14320 8774 14842 8810
rect 14320 8626 14832 8774
rect 18182 8770 18268 8774
rect 15550 8682 15568 8748
rect 15578 8710 15616 8738
rect 15658 8710 15690 8738
rect 15828 8696 16050 8744
rect 16052 8730 16058 8748
rect 16052 8702 16094 8730
rect 16102 8696 16122 8748
rect 16482 8700 16558 8728
rect 15762 8680 16122 8696
rect 16680 8684 16798 8748
rect 18074 8746 18192 8748
rect 18074 8742 18296 8746
rect 16842 8720 16880 8736
rect 17288 8694 17368 8722
rect 17504 8700 17584 8728
rect 17992 8720 18030 8738
rect 15424 8618 15452 8654
rect 15496 8652 15520 8674
rect 15518 8624 15520 8646
rect 8774 8442 8802 8506
rect 8924 8454 9278 8604
rect 12836 8578 12874 8606
rect 13098 8576 13144 8604
rect 14320 8558 14382 8574
rect 9522 8530 9584 8558
rect 10388 8518 10446 8546
rect 15424 8532 15452 8568
rect 12484 8502 12584 8512
rect 12844 8502 12944 8514
rect 13124 8502 13224 8512
rect 15762 8510 16116 8680
rect 16614 8514 16864 8684
rect 17368 8666 17396 8692
rect 17476 8672 17504 8692
rect 18074 8684 18192 8742
rect 18822 8734 19044 8744
rect 18314 8720 18342 8728
rect 18778 8706 19044 8734
rect 19182 8720 19200 8738
rect 18822 8696 19044 8706
rect 18008 8514 18258 8684
rect 18756 8510 19110 8696
rect 19276 8674 19300 9164
rect 19274 8554 19300 8674
rect 19304 8646 19328 9164
rect 19616 8940 19986 9106
rect 19616 8938 19784 8940
rect 19820 8938 19986 8940
rect 19734 8930 19986 8938
rect 19734 8924 19760 8930
rect 19750 8916 19760 8924
rect 19774 8916 19986 8930
rect 19750 8906 19986 8916
rect 20040 8906 20074 9194
rect 20174 9116 20274 9128
rect 20624 9064 20806 9356
rect 20922 9310 20958 9356
rect 20976 9364 21094 9380
rect 23610 9366 23726 9380
rect 23610 9364 23702 9366
rect 23722 9364 23726 9366
rect 20976 9310 21012 9364
rect 23648 9362 23668 9364
rect 23682 9362 23722 9364
rect 23734 9362 23768 9406
rect 23800 9400 23840 9418
rect 23800 9364 23840 9398
rect 23622 9330 23672 9362
rect 23682 9332 23702 9362
rect 23788 9336 23850 9364
rect 23734 9330 23850 9336
rect 23622 9314 23682 9330
rect 23722 9322 23838 9330
rect 23722 9314 23870 9322
rect 23622 9312 23870 9314
rect 20976 9308 21040 9310
rect 20976 9208 21018 9308
rect 23644 9294 23722 9312
rect 23734 9304 23870 9312
rect 23738 9294 23776 9296
rect 23778 9294 23870 9304
rect 23672 9268 23700 9286
rect 23734 9282 23768 9294
rect 23788 9292 23870 9294
rect 23734 9268 23788 9282
rect 23558 9242 23590 9258
rect 23644 9252 23652 9260
rect 23672 9256 23734 9268
rect 23592 9242 23624 9252
rect 23558 9220 23624 9242
rect 23644 9244 23656 9252
rect 23644 9220 23658 9244
rect 23672 9242 23700 9256
rect 23672 9231 23692 9242
rect 23558 9210 23658 9220
rect 23682 9214 23692 9231
rect 23704 9214 23722 9256
rect 23726 9253 23734 9256
rect 23738 9228 23756 9268
rect 23788 9267 23850 9268
rect 23836 9246 23850 9267
rect 23800 9230 23850 9246
rect 23788 9220 23850 9230
rect 23734 9214 23850 9220
rect 23672 9210 23850 9214
rect 20976 9182 21040 9208
rect 23558 9200 23850 9210
rect 23558 9194 23596 9200
rect 23600 9198 23850 9200
rect 23600 9194 23838 9198
rect 23558 9192 23590 9194
rect 20922 9132 20958 9182
rect 20976 9140 21012 9182
rect 23562 9172 23568 9192
rect 23622 9188 23838 9194
rect 23610 9180 23838 9188
rect 23610 9178 23812 9180
rect 23610 9160 23813 9178
rect 23672 9158 23788 9160
rect 23622 9108 23776 9158
rect 23672 9090 23726 9094
rect 23622 9068 23776 9090
rect 20174 9032 20274 9044
rect 20092 9010 20148 9014
rect 20088 9002 20148 9010
rect 20116 8974 20176 8986
rect 22588 8974 22606 9002
rect 22616 8980 22618 9046
rect 23610 9040 23818 9068
rect 23618 9038 23788 9040
rect 23562 9006 23568 9026
rect 23622 9014 23776 9038
rect 23788 9020 23813 9038
rect 23788 9018 23812 9020
rect 23788 9016 23838 9018
rect 23788 9014 23846 9016
rect 23558 9004 23590 9006
rect 20092 8948 20144 8952
rect 20092 8932 20176 8948
rect 20432 8932 20472 8948
rect 19750 8872 19752 8904
rect 19768 8896 19794 8906
rect 19768 8890 19784 8896
rect 19820 8892 19826 8900
rect 20092 8894 20144 8932
rect 20154 8898 20176 8914
rect 20116 8860 20176 8872
rect 19392 8744 19410 8852
rect 20088 8836 20148 8844
rect 20092 8832 20148 8836
rect 19426 8744 19438 8770
rect 19410 8742 19560 8744
rect 19398 8686 19560 8742
rect 19410 8684 19560 8686
rect 19352 8652 19376 8674
rect 19426 8658 19438 8684
rect 19302 8582 19328 8646
rect 19352 8624 19354 8646
rect 19430 8618 19458 8654
rect 20040 8626 20552 8828
rect 22644 8814 22754 8836
rect 22616 8786 22782 8808
rect 23128 8780 23438 9000
rect 23558 8998 23596 9004
rect 23622 9000 23846 9014
rect 23622 8998 23672 9000
rect 23558 8988 23672 8998
rect 23558 8956 23624 8988
rect 23558 8940 23590 8956
rect 23592 8946 23624 8956
rect 23648 8954 23658 8988
rect 23682 8967 23692 8998
rect 23648 8946 23656 8954
rect 23672 8952 23692 8967
rect 23704 8952 23722 8998
rect 23734 8978 23850 9000
rect 23738 8960 23756 8970
rect 23788 8968 23850 8978
rect 23672 8945 23726 8952
rect 23734 8945 23850 8960
rect 23672 8930 23850 8945
rect 23500 8906 23606 8926
rect 23692 8922 23726 8930
rect 23734 8906 23788 8930
rect 23500 8866 23694 8906
rect 23734 8905 23850 8906
rect 23734 8904 23799 8905
rect 23738 8902 23776 8904
rect 23722 8882 23776 8886
rect 23778 8884 23810 8904
rect 23778 8882 23846 8884
rect 23722 8868 23846 8882
rect 23500 8844 23702 8866
rect 23722 8844 23726 8864
rect 23734 8844 23768 8868
rect 23500 8834 23768 8844
rect 23788 8834 23850 8868
rect 23500 8798 23762 8834
rect 22476 8738 22514 8766
rect 22564 8738 22620 8766
rect 23128 8758 23490 8780
rect 23500 8776 23694 8798
rect 23722 8784 23788 8798
rect 23332 8746 23490 8758
rect 23436 8738 23490 8746
rect 23904 8738 23948 9030
rect 22484 8710 22548 8734
rect 24070 8696 24088 8712
rect 24098 8696 24132 8730
rect 24070 8662 24082 8696
rect 24104 8662 24120 8678
rect 24104 8644 24116 8662
rect 22668 8594 22758 8620
rect 15396 8504 15466 8508
rect 9226 8436 9278 8454
rect 10052 8386 10088 8454
rect 12732 8430 12742 8444
rect 12484 8418 12584 8428
rect 12844 8418 12944 8430
rect 13124 8418 13224 8428
rect 10180 8388 10280 8400
rect 10020 8376 10088 8386
rect 10052 8368 10088 8376
rect 12338 8374 12344 8376
rect 10052 8341 10242 8368
rect 10244 8341 10552 8368
rect 12320 8352 12344 8374
rect 12434 8368 12484 8408
rect 12428 8358 12484 8368
rect 12584 8368 12634 8408
rect 13074 8368 13124 8408
rect 12584 8358 12640 8368
rect 12428 8354 12443 8358
rect 8774 8092 8802 8156
rect 8924 8118 9278 8254
rect 8972 8104 9020 8118
rect 9226 8086 9278 8118
rect 9480 8242 9532 8338
rect 9580 8300 9636 8312
rect 10052 8304 10552 8341
rect 12308 8340 12344 8352
rect 12414 8352 12443 8354
rect 12625 8352 12640 8358
rect 13064 8358 13124 8368
rect 13064 8352 13079 8358
rect 12352 8342 12372 8348
rect 12278 8326 12346 8340
rect 12352 8336 12394 8342
rect 12308 8312 12342 8326
rect 10052 8300 10242 8304
rect 10244 8300 10552 8304
rect 10021 8285 10088 8300
rect 10036 8274 10088 8285
rect 10165 8274 10242 8300
rect 10280 8296 10313 8300
rect 9978 8270 10098 8274
rect 10165 8273 10278 8274
rect 10174 8272 10278 8273
rect 9976 8264 10098 8270
rect 10172 8264 10278 8272
rect 9966 8262 10278 8264
rect 9966 8256 10290 8262
rect 10312 8256 10313 8296
rect 10322 8256 10374 8286
rect 10438 8256 10470 8300
rect 10476 8278 10536 8300
rect 10472 8262 10526 8278
rect 10472 8256 10518 8262
rect 9966 8248 10299 8256
rect 8746 8064 8768 8078
rect 9480 8020 9834 8242
rect 9966 8238 10088 8248
rect 10002 8232 10088 8238
rect 10094 8246 10299 8248
rect 10094 8232 10178 8246
rect 10222 8241 10299 8246
rect 10312 8244 10518 8256
rect 10222 8240 10290 8241
rect 10312 8240 10484 8244
rect 10206 8232 10484 8240
rect 10002 8230 10484 8232
rect 10000 8229 10484 8230
rect 10540 8229 10552 8300
rect 12278 8298 12346 8312
rect 12352 8302 12376 8336
rect 12380 8302 12394 8336
rect 12414 8320 12488 8352
rect 12580 8320 13130 8352
rect 13236 8322 13270 8350
rect 13316 8324 13350 8352
rect 13394 8322 13782 8486
rect 13978 8434 14014 8496
rect 14032 8434 14068 8490
rect 14598 8470 14698 8482
rect 13950 8424 14014 8434
rect 14032 8324 14074 8424
rect 14598 8386 14698 8398
rect 14814 8390 14842 8426
rect 14724 8364 14780 8368
rect 14724 8356 14784 8364
rect 15270 8346 15450 8416
rect 18302 8390 18446 8414
rect 18276 8388 18446 8390
rect 18330 8362 18418 8386
rect 18304 8360 18418 8362
rect 14454 8332 14554 8344
rect 14598 8340 14698 8344
rect 14598 8332 14756 8340
rect 14696 8328 14756 8332
rect 13692 8318 13742 8322
rect 12308 8286 12344 8298
rect 12352 8296 12394 8302
rect 12352 8290 12372 8296
rect 12320 8264 12344 8286
rect 12414 8286 12488 8318
rect 12580 8286 13130 8318
rect 13316 8286 13350 8314
rect 13950 8306 14014 8324
rect 15270 8310 15452 8346
rect 12414 8284 12443 8286
rect 12428 8280 12443 8284
rect 12625 8280 12640 8286
rect 12428 8270 12484 8280
rect 12338 8262 12344 8264
rect 12434 8230 12484 8270
rect 12584 8270 12640 8280
rect 13064 8280 13079 8286
rect 13064 8270 13124 8280
rect 13978 8278 14014 8306
rect 12584 8230 12634 8270
rect 13074 8230 13124 8270
rect 13896 8256 14014 8278
rect 14032 8256 14068 8306
rect 15270 8260 15450 8310
rect 14454 8248 14554 8260
rect 14598 8248 14698 8260
rect 15270 8248 15592 8260
rect 10000 8228 10552 8229
rect 10000 8224 10318 8228
rect 10000 8220 10332 8224
rect 10000 8216 10008 8220
rect 9988 8204 10008 8216
rect 10052 8192 10158 8220
rect 10172 8210 10178 8220
rect 10194 8208 10332 8220
rect 9962 8156 10018 8170
rect 10052 8156 10154 8192
rect 10232 8188 10332 8208
rect 10422 8210 10484 8228
rect 15424 8224 15592 8248
rect 19276 8246 19300 8554
rect 19304 8274 19328 8582
rect 19430 8532 19458 8568
rect 19402 8504 19476 8508
rect 22400 8498 22772 8594
rect 20174 8470 20274 8482
rect 22400 8452 22836 8498
rect 22400 8440 22772 8452
rect 20040 8390 20068 8426
rect 22604 8420 22628 8440
rect 22638 8420 22694 8440
rect 22638 8406 22662 8420
rect 22672 8414 22694 8420
rect 20174 8386 20274 8398
rect 22612 8392 22628 8406
rect 22584 8368 22602 8390
rect 22638 8386 22646 8406
rect 22700 8386 22722 8440
rect 20092 8364 20148 8368
rect 20088 8356 20148 8364
rect 19436 8310 19464 8346
rect 20174 8340 20274 8344
rect 20116 8332 20274 8340
rect 20318 8332 20418 8344
rect 22700 8336 22742 8358
rect 20116 8328 20176 8332
rect 22716 8316 22762 8330
rect 22692 8308 22762 8316
rect 22692 8300 22742 8308
rect 22716 8284 22722 8300
rect 22716 8272 22762 8284
rect 19436 8224 19464 8260
rect 20174 8248 20274 8260
rect 20318 8248 20418 8260
rect 12484 8210 12584 8220
rect 10422 8200 10476 8210
rect 10492 8192 10538 8210
rect 12844 8208 12944 8220
rect 13124 8210 13224 8220
rect 12730 8194 12742 8208
rect 13896 8202 14014 8224
rect 10182 8156 10382 8188
rect 10520 8164 10566 8182
rect 10052 8138 10232 8156
rect 10332 8138 10388 8156
rect 10052 8099 10196 8138
rect 10373 8123 10456 8138
rect 12484 8126 12584 8136
rect 10052 8098 10232 8099
rect 10388 8098 10456 8123
rect 10052 8086 10456 8098
rect 9962 8072 10018 8086
rect 10052 8054 10088 8086
rect 10170 8084 10456 8086
rect 10232 8072 10332 8084
rect 12710 8070 12982 8182
rect 13124 8126 13224 8136
rect 13328 8070 13394 8182
rect 13978 8152 14014 8202
rect 14032 8152 14068 8202
rect 14032 8146 14098 8152
rect 14032 8076 14074 8146
rect 14014 8068 14026 8076
rect 9994 8040 10088 8054
rect 13896 8052 14026 8068
rect 10052 8036 10088 8040
rect 10124 8038 10142 8040
rect 10180 8038 10280 8050
rect 10020 8026 10088 8036
rect 10118 8034 10180 8038
rect 10052 8018 10088 8026
rect 10116 8023 10180 8034
rect 10280 8030 10442 8038
rect 10280 8029 10343 8030
rect 10280 8025 10342 8029
rect 10116 8018 10178 8023
rect 13950 8018 14026 8052
rect 9528 7992 9576 8006
rect 10052 7991 10242 8018
rect 10244 7991 10552 8018
rect 8746 7714 8772 7782
rect 8774 7742 8802 7806
rect 8924 7768 9278 7904
rect 8972 7754 9020 7768
rect 9226 7736 9278 7768
rect 9480 7892 9532 7988
rect 9580 7950 9636 7962
rect 10052 7954 10552 7991
rect 10052 7950 10242 7954
rect 10244 7950 10552 7954
rect 10021 7935 10088 7950
rect 10036 7924 10088 7935
rect 10165 7924 10242 7950
rect 10280 7946 10313 7950
rect 9978 7920 10098 7924
rect 10165 7923 10278 7924
rect 10174 7922 10278 7923
rect 9976 7914 10098 7920
rect 10172 7914 10278 7922
rect 9966 7912 10278 7914
rect 9966 7906 10290 7912
rect 10312 7906 10313 7946
rect 10322 7906 10374 7936
rect 10438 7906 10470 7950
rect 10476 7928 10536 7950
rect 10472 7912 10526 7928
rect 10472 7906 10518 7912
rect 9966 7898 10299 7906
rect 9480 7670 9834 7892
rect 9966 7888 10088 7898
rect 10002 7882 10088 7888
rect 10094 7896 10299 7898
rect 10094 7882 10178 7896
rect 10222 7891 10299 7896
rect 10312 7894 10518 7906
rect 10222 7890 10290 7891
rect 10312 7890 10484 7894
rect 10206 7882 10484 7890
rect 10002 7880 10484 7882
rect 10000 7879 10484 7880
rect 10532 7879 10538 7882
rect 10540 7879 10552 7950
rect 13978 7928 14026 8018
rect 14032 8018 14046 8068
rect 14032 7968 14080 8018
rect 13102 7914 13220 7916
rect 10000 7878 10552 7879
rect 10000 7874 10318 7878
rect 10000 7870 10332 7874
rect 10000 7866 10008 7870
rect 9988 7854 10008 7866
rect 10052 7842 10158 7870
rect 10172 7860 10178 7870
rect 10194 7858 10332 7870
rect 9962 7806 10018 7820
rect 10052 7806 10154 7842
rect 10232 7838 10332 7858
rect 10422 7860 10484 7878
rect 10532 7860 10538 7878
rect 10422 7850 10476 7860
rect 10492 7842 10538 7860
rect 10182 7806 10382 7838
rect 10560 7832 10566 7888
rect 12484 7862 12584 7872
rect 12844 7862 12944 7874
rect 13124 7862 13224 7872
rect 13064 7860 13274 7862
rect 14184 7852 14366 8106
rect 15424 7970 15452 8006
rect 19430 7970 19458 8006
rect 15424 7884 15452 7920
rect 19430 7884 19458 7920
rect 10520 7814 10566 7832
rect 10052 7788 10232 7806
rect 10332 7788 10388 7806
rect 10052 7749 10196 7788
rect 10373 7773 10456 7788
rect 12484 7778 12584 7788
rect 12844 7778 12944 7790
rect 13124 7778 13224 7788
rect 10052 7748 10232 7749
rect 10388 7748 10456 7773
rect 10052 7736 10456 7748
rect 9962 7722 10018 7736
rect 10052 7704 10088 7736
rect 10170 7734 10456 7736
rect 12338 7734 12344 7736
rect 10232 7722 10332 7734
rect 12320 7712 12344 7734
rect 12434 7728 12484 7768
rect 12428 7718 12484 7728
rect 12584 7728 12634 7768
rect 13074 7728 13124 7768
rect 12584 7718 12640 7728
rect 12428 7714 12443 7718
rect 9994 7690 10088 7704
rect 12308 7700 12344 7712
rect 12414 7712 12443 7714
rect 12625 7712 12640 7718
rect 13064 7718 13124 7728
rect 13064 7712 13079 7718
rect 12352 7702 12372 7708
rect 10052 7686 10088 7690
rect 10124 7688 10142 7690
rect 10180 7688 10280 7700
rect 10020 7676 10088 7686
rect 10118 7684 10180 7688
rect 10052 7668 10088 7676
rect 10116 7673 10180 7684
rect 10280 7680 10442 7688
rect 12278 7686 12346 7700
rect 12352 7696 12394 7702
rect 10280 7679 10343 7680
rect 10280 7675 10342 7679
rect 10116 7668 10178 7673
rect 12308 7672 12342 7686
rect 9528 7642 9576 7656
rect 10052 7641 10242 7668
rect 10244 7641 10552 7668
rect 12278 7658 12346 7672
rect 12352 7662 12376 7696
rect 12380 7662 12394 7696
rect 12414 7680 12488 7712
rect 12580 7680 13130 7712
rect 13236 7682 13270 7710
rect 13316 7684 13350 7712
rect 13394 7680 13782 7846
rect 13978 7776 14014 7846
rect 14032 7776 14068 7832
rect 14438 7796 14620 7852
rect 14438 7784 14672 7796
rect 14716 7784 14816 7796
rect 13950 7774 14014 7776
rect 13692 7678 13742 7680
rect 12308 7646 12344 7658
rect 12352 7656 12394 7662
rect 12352 7650 12372 7656
rect 8774 7392 8802 7456
rect 8924 7418 9278 7554
rect 9226 7386 9278 7418
rect 9480 7542 9532 7638
rect 9580 7600 9636 7612
rect 10052 7604 10552 7641
rect 12320 7624 12344 7646
rect 12414 7646 12488 7678
rect 12580 7646 13130 7678
rect 14032 7674 14074 7774
rect 14438 7712 14620 7784
rect 14814 7712 14874 7716
rect 14438 7700 14672 7712
rect 14716 7704 14874 7712
rect 14716 7700 14816 7704
rect 15088 7702 15120 7730
rect 15170 7702 15208 7730
rect 15250 7702 15282 7730
rect 14438 7674 14620 7700
rect 14842 7680 14902 7688
rect 14842 7676 14898 7680
rect 13316 7646 13350 7674
rect 13950 7648 14014 7674
rect 12414 7644 12443 7646
rect 12428 7640 12443 7644
rect 12625 7640 12640 7646
rect 12428 7630 12484 7640
rect 12338 7622 12344 7624
rect 10052 7600 10242 7604
rect 10244 7600 10552 7604
rect 10021 7585 10088 7600
rect 10036 7574 10088 7585
rect 10165 7574 10242 7600
rect 10280 7596 10313 7600
rect 9978 7570 10098 7574
rect 10165 7573 10278 7574
rect 10174 7572 10278 7573
rect 9976 7564 10098 7570
rect 10172 7564 10278 7572
rect 9966 7562 10278 7564
rect 9966 7556 10290 7562
rect 10312 7556 10313 7596
rect 10322 7556 10374 7586
rect 10438 7556 10470 7600
rect 10476 7578 10536 7600
rect 10472 7562 10526 7578
rect 10472 7556 10518 7562
rect 9966 7548 10299 7556
rect 9480 7320 9834 7542
rect 9966 7538 10088 7548
rect 10002 7532 10088 7538
rect 10094 7546 10299 7548
rect 10094 7532 10178 7546
rect 10222 7541 10299 7546
rect 10312 7544 10518 7556
rect 10222 7540 10290 7541
rect 10312 7540 10484 7544
rect 10206 7532 10484 7540
rect 10002 7530 10484 7532
rect 10000 7529 10484 7530
rect 10540 7529 10552 7600
rect 12434 7590 12484 7630
rect 12584 7630 12640 7640
rect 13064 7640 13079 7646
rect 13064 7630 13124 7640
rect 13978 7630 14014 7648
rect 12584 7590 12634 7630
rect 13074 7590 13124 7630
rect 13896 7606 14014 7630
rect 14032 7616 14068 7648
rect 14184 7616 14366 7674
rect 14032 7598 14366 7616
rect 10000 7528 10552 7529
rect 10000 7524 10318 7528
rect 10000 7520 10332 7524
rect 10000 7516 10008 7520
rect 9988 7504 10008 7516
rect 10052 7492 10158 7520
rect 10172 7510 10178 7520
rect 10194 7508 10332 7520
rect 9962 7456 10018 7470
rect 10052 7456 10154 7492
rect 10232 7488 10332 7508
rect 10422 7510 10484 7528
rect 10422 7500 10476 7510
rect 10492 7492 10538 7510
rect 10182 7456 10382 7488
rect 10520 7464 10566 7482
rect 12288 7456 12292 7570
rect 12316 7484 12320 7582
rect 12484 7570 12584 7580
rect 12844 7568 12944 7580
rect 13124 7570 13224 7580
rect 12730 7554 12742 7568
rect 13896 7552 14014 7576
rect 14184 7562 14366 7598
rect 13978 7506 14014 7552
rect 14032 7544 14366 7562
rect 14032 7506 14068 7544
rect 13950 7504 14014 7506
rect 12484 7486 12584 7496
rect 12844 7484 12944 7496
rect 13124 7486 13224 7496
rect 10052 7438 10232 7456
rect 10332 7438 10388 7456
rect 10052 7399 10196 7438
rect 10373 7423 10456 7438
rect 10052 7398 10232 7399
rect 10388 7398 10456 7423
rect 10052 7386 10456 7398
rect 12858 7392 12874 7410
rect 9962 7372 10018 7386
rect 10052 7354 10088 7386
rect 10170 7384 10456 7386
rect 10232 7372 10332 7384
rect 13098 7382 13144 7410
rect 13692 7382 13742 7410
rect 14032 7404 14074 7504
rect 14184 7420 14366 7544
rect 14438 7654 14950 7674
rect 15424 7664 15452 7700
rect 19430 7664 19458 7700
rect 14438 7618 14960 7654
rect 15016 7622 15044 7658
rect 14438 7470 14950 7618
rect 15424 7578 15452 7614
rect 15016 7536 15044 7572
rect 15496 7510 15528 7538
rect 15578 7512 15616 7540
rect 15658 7524 15662 7540
rect 15946 7532 16168 7580
rect 13950 7378 14014 7404
rect 9994 7340 10088 7354
rect 10052 7336 10088 7340
rect 10124 7338 10142 7340
rect 10180 7338 10280 7350
rect 10020 7326 10088 7336
rect 10118 7334 10180 7338
rect 10052 7318 10088 7326
rect 10116 7323 10180 7334
rect 10280 7330 10442 7338
rect 13978 7336 14014 7378
rect 10280 7329 10343 7330
rect 10280 7325 10342 7329
rect 14032 7328 14068 7378
rect 10116 7318 10178 7323
rect 9528 7292 9562 7306
rect 10052 7291 10242 7318
rect 10244 7291 10552 7318
rect 8924 7068 9278 7222
rect 9480 7054 9532 7288
rect 9580 7250 9636 7262
rect 10052 7254 10552 7291
rect 14438 7260 14620 7420
rect 14716 7316 14816 7328
rect 10052 7250 10242 7254
rect 10244 7250 10552 7254
rect 10021 7235 10088 7250
rect 10036 7224 10088 7235
rect 10165 7224 10242 7250
rect 10280 7246 10313 7250
rect 9978 7220 10098 7224
rect 10165 7223 10278 7224
rect 10174 7222 10278 7223
rect 9976 7214 10098 7220
rect 10172 7214 10278 7222
rect 9966 7212 10278 7214
rect 9966 7206 10290 7212
rect 10312 7206 10313 7246
rect 10322 7206 10374 7236
rect 10438 7206 10470 7250
rect 10476 7228 10536 7250
rect 10472 7212 10526 7228
rect 10472 7206 10518 7212
rect 9966 7198 10299 7206
rect 9966 7188 10088 7198
rect 10002 7182 10088 7188
rect 10094 7196 10299 7198
rect 10094 7182 10178 7196
rect 10222 7191 10299 7196
rect 10312 7194 10518 7206
rect 10222 7190 10290 7191
rect 10312 7190 10484 7194
rect 10206 7182 10484 7190
rect 10002 7180 10484 7182
rect 10000 7179 10484 7180
rect 10540 7179 10552 7250
rect 14916 7258 14950 7382
rect 15034 7340 15044 7354
rect 14716 7232 14816 7244
rect 14916 7236 14960 7258
rect 14842 7210 14898 7214
rect 14842 7202 14902 7210
rect 10000 7178 10552 7179
rect 9580 7166 9636 7178
rect 10000 7174 10318 7178
rect 10000 7170 10332 7174
rect 10422 7170 10484 7178
rect 14814 7174 14874 7186
rect 10000 7166 10008 7170
rect 9988 7154 10008 7166
rect 10052 7166 10158 7170
rect 10172 7166 10178 7170
rect 10194 7166 10332 7170
rect 10388 7166 10484 7170
rect 10052 7158 10538 7166
rect 10004 7140 10006 7154
rect 10052 7142 10212 7158
rect 10232 7142 10538 7158
rect 14438 7150 14842 7166
rect 14846 7144 14898 7152
rect 10052 7138 10154 7142
rect 10232 7138 10332 7142
rect 14518 7138 14558 7144
rect 14814 7138 14898 7144
rect 9976 7120 10006 7138
rect 9678 7106 9734 7118
rect 9962 7106 10018 7120
rect 10052 7114 10566 7138
rect 14410 7132 14898 7138
rect 14410 7122 14842 7132
rect 10052 7106 10154 7114
rect 10182 7106 10382 7114
rect 10052 7088 10232 7106
rect 10332 7088 10388 7106
rect 14814 7098 14836 7110
rect 14846 7090 14898 7132
rect 14916 7128 14950 7236
rect 15004 7130 15374 7294
rect 15510 7264 15528 7396
rect 15880 7346 16234 7532
rect 16518 7528 16558 7538
rect 16798 7522 16916 7592
rect 19430 7578 19458 7614
rect 23126 7552 23498 7794
rect 16732 7358 16982 7522
rect 17288 7510 17368 7538
rect 17504 7510 17584 7538
rect 17992 7510 18040 7538
rect 18314 7510 18390 7540
rect 18778 7510 18826 7538
rect 19182 7524 19200 7540
rect 19344 7512 19376 7540
rect 15482 7258 15556 7264
rect 15510 7244 15528 7258
rect 15528 7236 15678 7244
rect 15504 7228 15678 7236
rect 15504 7208 15532 7228
rect 15004 7126 15216 7130
rect 15230 7126 15374 7130
rect 15088 7120 15120 7126
rect 15144 7122 15374 7126
rect 15144 7120 15150 7122
rect 15170 7106 15374 7122
rect 10052 7054 10154 7088
rect 10170 7054 10196 7088
rect 10373 7073 10456 7088
rect 15192 7080 15198 7100
rect 15224 7096 15250 7106
rect 15224 7090 15240 7096
rect 10388 7054 10456 7073
rect 14814 7044 14932 7068
rect 9678 7022 9734 7034
rect 9962 7022 10018 7036
rect 10232 7022 10332 7034
rect 14842 7024 14904 7040
rect 14438 7006 14950 7024
rect 14438 6970 14960 7006
rect 15016 6974 15044 7010
rect 14438 6822 14950 6970
rect 15378 6940 16056 7082
rect 15016 6888 15044 6924
rect 15378 6916 16168 6940
rect 15378 6882 15464 6916
rect 15546 6914 16168 6916
rect 15546 6902 15648 6914
rect 15546 6884 15632 6902
rect 15582 6882 15632 6884
rect 4658 6752 4716 6780
rect 8738 6714 8814 6722
rect 8776 6712 8810 6714
rect 4778 6644 5030 6664
rect 5028 6638 5030 6644
rect 5088 6638 5092 6664
rect 4806 6616 5030 6636
rect 5000 6610 5030 6616
rect 5088 6610 5120 6636
rect 4940 6504 4948 6546
rect 4968 6476 4976 6526
rect 5006 6462 5032 6526
rect 5034 6434 5060 6554
rect 5184 6542 5208 6642
rect 5212 6570 5236 6614
rect 5254 6570 5276 6614
rect 5212 6550 5276 6570
rect 5212 6548 5274 6550
rect 5282 6542 5304 6642
rect 5184 6522 5304 6542
rect 5314 6542 5334 6642
rect 8766 6630 8794 6694
rect 8916 6642 9270 6792
rect 9514 6718 9576 6746
rect 9582 6738 9604 6758
rect 12834 6742 12884 6766
rect 10380 6706 10438 6734
rect 12842 6724 12880 6742
rect 13104 6722 13150 6750
rect 13246 6716 13312 6732
rect 13234 6688 13284 6704
rect 14716 6666 14816 6678
rect 15016 6668 15044 6704
rect 15546 6660 15632 6882
rect 15662 6874 15676 6914
rect 15778 6902 15810 6914
rect 15946 6906 16168 6914
rect 16602 6916 16678 7064
rect 15946 6890 16206 6906
rect 16602 6896 16770 6916
rect 15946 6878 16168 6890
rect 15946 6876 16178 6878
rect 15880 6838 16234 6876
rect 16798 6872 16916 6944
rect 17408 6916 17488 7056
rect 17488 6888 17576 6916
rect 15880 6812 16458 6838
rect 15880 6810 16234 6812
rect 15880 6784 16458 6810
rect 15880 6706 16234 6784
rect 16732 6710 16982 6872
rect 18070 6668 18152 6684
rect 12490 6648 12590 6658
rect 12850 6648 12950 6660
rect 13130 6648 13230 6658
rect 9218 6624 9270 6642
rect 5342 6570 5362 6614
rect 10044 6574 10080 6642
rect 10172 6576 10272 6588
rect 12738 6576 12748 6590
rect 5342 6548 5404 6570
rect 10012 6564 10080 6574
rect 12490 6564 12590 6574
rect 12850 6564 12950 6576
rect 13130 6564 13230 6574
rect 10044 6556 10080 6564
rect 5184 6520 5302 6522
rect 5314 6520 5432 6542
rect 10044 6529 10234 6556
rect 10236 6529 10544 6556
rect 5364 6458 5388 6504
rect 4806 6232 4856 6276
rect 5418 6272 5442 6458
rect 8766 6280 8794 6344
rect 8916 6306 9270 6442
rect 8964 6292 9012 6306
rect 9218 6274 9270 6306
rect 9472 6430 9524 6526
rect 9572 6488 9628 6500
rect 10044 6492 10544 6529
rect 12344 6520 12350 6522
rect 12326 6498 12350 6520
rect 12440 6514 12490 6554
rect 12434 6504 12490 6514
rect 12590 6514 12640 6554
rect 13080 6514 13130 6554
rect 12590 6504 12646 6514
rect 12434 6500 12449 6504
rect 10044 6488 10234 6492
rect 10236 6488 10544 6492
rect 10013 6473 10080 6488
rect 10028 6462 10080 6473
rect 10157 6462 10234 6488
rect 10272 6484 10305 6488
rect 9970 6458 10090 6462
rect 10157 6461 10270 6462
rect 10166 6460 10270 6461
rect 9968 6452 10090 6458
rect 10164 6452 10270 6460
rect 9958 6450 10270 6452
rect 9958 6444 10282 6450
rect 10304 6444 10305 6484
rect 10314 6444 10366 6474
rect 10430 6444 10462 6488
rect 10468 6466 10528 6488
rect 10464 6450 10518 6466
rect 10464 6444 10510 6450
rect 9958 6436 10291 6444
rect 4868 6208 4884 6260
rect 9472 6208 9826 6430
rect 9958 6426 10080 6436
rect 9994 6420 10080 6426
rect 10086 6434 10291 6436
rect 10086 6420 10170 6434
rect 10214 6429 10291 6434
rect 10304 6432 10510 6444
rect 10214 6428 10282 6429
rect 10304 6428 10476 6432
rect 10198 6420 10476 6428
rect 9994 6418 10476 6420
rect 9992 6417 10476 6418
rect 10532 6417 10544 6488
rect 12314 6486 12350 6498
rect 12420 6498 12449 6500
rect 12631 6498 12646 6504
rect 13070 6504 13130 6514
rect 13070 6498 13085 6504
rect 12358 6488 12378 6494
rect 12284 6472 12352 6486
rect 12358 6482 12400 6488
rect 12314 6458 12348 6472
rect 12284 6444 12352 6458
rect 12358 6448 12382 6482
rect 12386 6448 12400 6482
rect 12420 6466 12494 6498
rect 12586 6466 13136 6498
rect 13242 6468 13276 6496
rect 13322 6470 13356 6498
rect 13400 6468 13864 6632
rect 14716 6582 14816 6594
rect 14932 6586 14960 6622
rect 15016 6582 15044 6618
rect 14842 6560 14898 6564
rect 14842 6552 14902 6560
rect 14904 6552 14914 6574
rect 14572 6528 14672 6540
rect 14716 6536 14816 6540
rect 14886 6536 14902 6552
rect 14716 6528 14874 6536
rect 14814 6524 14874 6528
rect 14858 6508 14874 6524
rect 14886 6520 14932 6536
rect 15088 6508 15120 6536
rect 15170 6508 15208 6536
rect 15250 6508 15282 6536
rect 15376 6530 15464 6614
rect 15544 6530 15632 6660
rect 16082 6628 16096 6646
rect 16110 6644 16124 6668
rect 16100 6628 16124 6644
rect 18036 6662 18152 6668
rect 18156 6662 18258 6668
rect 18036 6644 18258 6662
rect 18036 6620 18044 6644
rect 18070 6640 18196 6644
rect 18064 6632 18286 6640
rect 18064 6616 18122 6632
rect 18064 6592 18068 6616
rect 18070 6590 18122 6616
rect 18138 6616 18286 6632
rect 18138 6604 18196 6616
rect 18138 6590 18153 6604
rect 18070 6584 18130 6590
rect 18064 6582 18130 6584
rect 18132 6586 18164 6590
rect 18064 6576 18128 6582
rect 18064 6574 18126 6576
rect 18064 6554 18126 6556
rect 18064 6548 18128 6554
rect 18132 6548 18184 6586
rect 18064 6546 18184 6548
rect 17556 6534 17558 6546
rect 18070 6544 18184 6546
rect 18250 6544 18284 6586
rect 18362 6544 18396 6586
rect 18476 6544 18510 6586
rect 18544 6544 18578 6586
rect 18070 6540 18164 6544
rect 14858 6492 14904 6508
rect 13698 6464 13748 6468
rect 12314 6432 12350 6444
rect 12358 6442 12400 6448
rect 12358 6436 12378 6442
rect 9992 6416 10544 6417
rect 9992 6412 10310 6416
rect 9992 6408 10324 6412
rect 9992 6404 10000 6408
rect 9980 6392 10000 6404
rect 10044 6380 10150 6408
rect 10164 6398 10170 6408
rect 10186 6396 10324 6408
rect 9954 6344 10010 6358
rect 10044 6344 10146 6380
rect 10224 6376 10324 6396
rect 10414 6398 10476 6416
rect 12326 6410 12350 6432
rect 12420 6432 12494 6464
rect 12586 6432 13136 6464
rect 13322 6432 13356 6460
rect 14572 6444 14672 6456
rect 14716 6444 14816 6456
rect 15376 6446 15442 6530
rect 15544 6468 15610 6530
rect 17720 6494 17742 6518
rect 17748 6490 17770 6494
rect 18036 6490 18044 6510
rect 18064 6490 18068 6538
rect 18070 6526 18153 6540
rect 18070 6496 18196 6526
rect 18100 6468 18196 6496
rect 12420 6430 12449 6432
rect 12434 6426 12449 6430
rect 12631 6426 12646 6432
rect 12434 6416 12490 6426
rect 12344 6408 12350 6410
rect 10414 6388 10468 6398
rect 10484 6380 10530 6398
rect 12440 6376 12490 6416
rect 12590 6416 12646 6426
rect 13070 6426 13085 6432
rect 13070 6416 13130 6426
rect 12590 6376 12640 6416
rect 13080 6376 13130 6416
rect 15544 6406 15632 6468
rect 18100 6446 18152 6468
rect 10174 6344 10374 6376
rect 10512 6352 10558 6370
rect 12490 6356 12590 6366
rect 12850 6354 12950 6366
rect 13130 6356 13230 6366
rect 10044 6326 10224 6344
rect 10324 6326 10380 6344
rect 12736 6340 12748 6354
rect 10044 6287 10188 6326
rect 10365 6311 10448 6326
rect 10044 6286 10224 6287
rect 10380 6286 10448 6311
rect 10044 6274 10448 6286
rect 9954 6260 10010 6274
rect 10044 6242 10080 6274
rect 10162 6272 10448 6274
rect 12490 6272 12590 6282
rect 10224 6260 10324 6272
rect 9986 6228 10080 6242
rect 10044 6224 10080 6228
rect 10116 6226 10134 6228
rect 10172 6226 10272 6238
rect 10012 6214 10080 6224
rect 10110 6222 10172 6226
rect 10044 6206 10080 6214
rect 10108 6211 10172 6222
rect 10272 6218 10434 6226
rect 10272 6217 10335 6218
rect 10272 6213 10334 6217
rect 12716 6216 13400 6328
rect 10108 6206 10170 6211
rect 5320 6190 5334 6194
rect 4986 6164 4996 6165
rect 4904 6130 4938 6150
rect 4850 6114 4880 6118
rect 4884 6084 4914 6114
rect 4918 6082 4924 6130
rect 4946 6110 4952 6158
rect 4986 6150 5001 6164
rect 5320 6152 5388 6190
rect 9520 6180 9568 6194
rect 10044 6179 10234 6206
rect 10236 6179 10544 6206
rect 5320 6150 5334 6152
rect 5348 6150 5388 6152
rect 4986 6120 5042 6150
rect 5256 6120 5280 6150
rect 5320 6120 5388 6150
rect 5510 6130 5538 6176
rect 4986 6105 5001 6120
rect 5320 6096 5334 6120
rect 5348 6102 5422 6120
rect 5373 6096 5388 6102
rect 4934 6078 4944 6094
rect 4986 6092 5042 6093
rect 4986 6078 5150 6092
rect 5241 6078 5280 6093
rect 5320 6080 5388 6096
rect 5320 6074 5402 6080
rect 5322 6060 5334 6074
rect 4920 6048 5056 6056
rect 5322 6038 5342 6060
rect 5350 6048 5370 6058
rect 5350 6046 5412 6048
rect 5350 6038 5370 6046
rect 5322 6002 5344 6038
rect 5322 5996 5342 6002
rect 4806 5924 4856 5968
rect 5322 5966 5334 5996
rect 5350 5994 5372 6038
rect 4868 5898 4884 5950
rect 4942 5768 4950 5772
rect 4668 5738 4680 5765
rect 4668 5684 4683 5738
rect 4942 5726 4956 5768
rect 4668 5670 4680 5684
rect 4942 5670 4950 5726
rect 4974 5698 4984 5750
rect 5384 5742 5400 5998
rect 5420 5778 5436 5962
rect 4976 5692 4984 5698
rect 4668 5629 4683 5670
rect 5512 5634 5568 6028
rect 8766 5930 8794 5994
rect 8916 5956 9270 6092
rect 8964 5942 9012 5956
rect 9218 5924 9270 5956
rect 9472 6080 9524 6176
rect 9572 6138 9628 6150
rect 10044 6142 10544 6179
rect 10044 6138 10234 6142
rect 10236 6138 10544 6142
rect 10013 6123 10080 6138
rect 10028 6112 10080 6123
rect 10157 6112 10234 6138
rect 10272 6134 10305 6138
rect 9970 6108 10090 6112
rect 10157 6111 10270 6112
rect 10166 6110 10270 6111
rect 9968 6102 10090 6108
rect 10164 6102 10270 6110
rect 9958 6100 10270 6102
rect 9958 6094 10282 6100
rect 10304 6094 10305 6134
rect 10314 6094 10366 6124
rect 10430 6094 10462 6138
rect 10468 6116 10528 6138
rect 10464 6100 10518 6116
rect 10464 6094 10510 6100
rect 9958 6086 10291 6094
rect 9472 5858 9826 6080
rect 9958 6076 10080 6086
rect 9994 6070 10080 6076
rect 10086 6084 10291 6086
rect 10086 6070 10170 6084
rect 10214 6079 10291 6084
rect 10304 6082 10510 6094
rect 10214 6078 10282 6079
rect 10304 6078 10476 6082
rect 10198 6070 10476 6078
rect 9994 6068 10476 6070
rect 9992 6067 10476 6068
rect 10532 6067 10544 6138
rect 9992 6066 10544 6067
rect 9992 6062 10310 6066
rect 9992 6058 10324 6062
rect 9992 6054 10000 6058
rect 9980 6042 10000 6054
rect 10044 6030 10150 6058
rect 10164 6048 10170 6058
rect 10186 6046 10324 6058
rect 9954 5994 10010 6008
rect 10044 5994 10146 6030
rect 10224 6026 10324 6046
rect 10414 6048 10476 6066
rect 10414 6038 10468 6048
rect 10484 6030 10530 6048
rect 10174 5994 10374 6026
rect 10512 6002 10558 6020
rect 12490 6008 12590 6018
rect 12850 6008 12950 6020
rect 13130 6008 13230 6018
rect 10044 5976 10224 5994
rect 10324 5976 10380 5994
rect 10044 5937 10188 5976
rect 10365 5961 10448 5976
rect 10044 5936 10224 5937
rect 10380 5936 10448 5961
rect 10044 5924 10448 5936
rect 12490 5924 12590 5934
rect 12850 5924 12950 5936
rect 13130 5924 13230 5934
rect 9954 5910 10010 5924
rect 10044 5892 10080 5924
rect 10162 5922 10448 5924
rect 10224 5910 10324 5922
rect 9986 5878 10080 5892
rect 10044 5874 10080 5878
rect 10116 5876 10134 5878
rect 10172 5876 10272 5888
rect 12344 5880 12350 5882
rect 10012 5864 10080 5874
rect 10110 5872 10172 5876
rect 10044 5856 10080 5864
rect 10108 5861 10172 5872
rect 10272 5868 10434 5876
rect 10272 5867 10335 5868
rect 10272 5863 10334 5867
rect 10108 5856 10170 5861
rect 12326 5858 12350 5880
rect 12440 5874 12490 5914
rect 12434 5864 12490 5874
rect 12590 5874 12640 5914
rect 13080 5874 13130 5914
rect 12590 5864 12646 5874
rect 12434 5860 12449 5864
rect 9520 5830 9568 5844
rect 10044 5829 10234 5856
rect 10236 5829 10544 5856
rect 12314 5846 12350 5858
rect 12420 5858 12449 5860
rect 12631 5858 12646 5864
rect 13070 5864 13130 5874
rect 13070 5858 13085 5864
rect 12358 5848 12378 5854
rect 12284 5832 12352 5846
rect 12358 5842 12400 5848
rect 4668 5554 4685 5629
rect 5180 5570 5198 5614
rect 4668 5526 4704 5554
rect 5208 5542 5226 5594
rect 5254 5530 5272 5594
rect 4632 5500 4704 5526
rect 5282 5502 5300 5622
rect 4650 5486 4704 5500
rect 5322 5490 5334 5610
rect 5350 5518 5362 5582
rect 8766 5580 8794 5644
rect 8916 5606 9270 5742
rect 9218 5574 9270 5606
rect 9472 5730 9524 5826
rect 9572 5788 9628 5800
rect 10044 5792 10544 5829
rect 12314 5818 12348 5832
rect 12284 5804 12352 5818
rect 12358 5808 12382 5842
rect 12386 5808 12400 5842
rect 12420 5826 12494 5858
rect 12586 5826 13136 5858
rect 13242 5828 13276 5856
rect 13322 5830 13356 5858
rect 13400 5826 13864 5992
rect 15400 5966 15452 5968
rect 15438 5940 15454 5950
rect 15428 5938 15454 5940
rect 15438 5926 15454 5938
rect 13698 5824 13748 5826
rect 12314 5792 12350 5804
rect 12358 5802 12400 5808
rect 12358 5796 12378 5802
rect 10044 5788 10234 5792
rect 10236 5788 10544 5792
rect 10013 5773 10080 5788
rect 10028 5762 10080 5773
rect 10157 5762 10234 5788
rect 10272 5784 10305 5788
rect 9970 5758 10090 5762
rect 10157 5761 10270 5762
rect 10166 5760 10270 5761
rect 9968 5752 10090 5758
rect 10164 5752 10270 5760
rect 9958 5750 10270 5752
rect 9958 5744 10282 5750
rect 10304 5744 10305 5784
rect 10314 5744 10366 5774
rect 10430 5744 10462 5788
rect 10468 5766 10528 5788
rect 10464 5750 10518 5766
rect 10464 5744 10510 5750
rect 9958 5736 10291 5744
rect 9472 5508 9826 5730
rect 9958 5726 10080 5736
rect 9994 5720 10080 5726
rect 10086 5734 10291 5736
rect 10086 5720 10170 5734
rect 10214 5729 10291 5734
rect 10304 5732 10510 5744
rect 10214 5728 10282 5729
rect 10304 5728 10476 5732
rect 10198 5720 10476 5728
rect 9994 5718 10476 5720
rect 9992 5717 10476 5718
rect 10532 5717 10544 5788
rect 12326 5770 12350 5792
rect 12420 5792 12494 5824
rect 12586 5792 13136 5824
rect 13322 5792 13356 5820
rect 12420 5790 12449 5792
rect 12434 5786 12449 5790
rect 12631 5786 12646 5792
rect 12434 5776 12490 5786
rect 12344 5768 12350 5770
rect 9992 5716 10544 5717
rect 12110 5716 12356 5748
rect 12440 5736 12490 5776
rect 12590 5776 12646 5786
rect 13070 5786 13085 5792
rect 13070 5776 13130 5786
rect 15522 5780 15526 5782
rect 15546 5780 15632 6406
rect 16082 6304 16132 6320
rect 16082 6300 16116 6304
rect 16110 6276 16160 6292
rect 16110 6272 16144 6276
rect 18036 6268 18082 6308
rect 18288 6268 18334 6310
rect 18070 6114 18152 6130
rect 18036 6108 18152 6114
rect 18156 6108 18258 6114
rect 18036 6090 18258 6108
rect 18036 6066 18044 6090
rect 18070 6086 18196 6090
rect 18064 6078 18286 6086
rect 18064 6062 18122 6078
rect 18064 6038 18068 6062
rect 18070 6036 18122 6062
rect 18138 6062 18286 6078
rect 18138 6054 18262 6062
rect 18138 6050 18196 6054
rect 18138 6036 18153 6050
rect 18180 6046 18186 6050
rect 18224 6046 18226 6054
rect 18224 6044 18228 6046
rect 18224 6042 18232 6044
rect 18070 6028 18130 6036
rect 18132 6032 18164 6036
rect 18168 6032 18234 6042
rect 18252 6032 18260 6054
rect 18064 6022 18128 6028
rect 18132 6026 18234 6032
rect 18064 5996 18128 6000
rect 18132 5996 18184 6026
rect 18224 5996 18232 6026
rect 18064 5994 18234 5996
rect 18070 5990 18234 5994
rect 18250 5990 18284 6032
rect 18362 5990 18396 6032
rect 18476 5990 18510 6032
rect 18544 5990 18578 6032
rect 18070 5986 18164 5990
rect 18036 5936 18044 5956
rect 18064 5936 18068 5984
rect 18070 5972 18153 5986
rect 18168 5984 18234 5990
rect 18224 5980 18232 5984
rect 18070 5968 18196 5972
rect 18252 5968 18260 5990
rect 18070 5956 18262 5968
rect 18070 5942 18196 5956
rect 18252 5952 18260 5956
rect 18100 5914 18196 5942
rect 18100 5892 18152 5914
rect 12590 5736 12640 5776
rect 13080 5736 13130 5776
rect 15516 5742 15526 5780
rect 15544 5770 15632 5780
rect 12490 5716 12590 5726
rect 9992 5712 10310 5716
rect 9992 5708 10324 5712
rect 9992 5704 10000 5708
rect 9980 5692 10000 5704
rect 10044 5680 10150 5708
rect 10164 5698 10170 5708
rect 10186 5696 10324 5708
rect 9954 5644 10010 5658
rect 10044 5644 10146 5680
rect 10224 5676 10324 5696
rect 10414 5698 10476 5716
rect 10414 5688 10468 5698
rect 10484 5680 10530 5698
rect 10174 5644 10374 5676
rect 10512 5652 10558 5670
rect 10044 5626 10224 5644
rect 10324 5626 10380 5644
rect 10044 5587 10188 5626
rect 10365 5611 10448 5626
rect 10044 5586 10224 5587
rect 10380 5586 10448 5611
rect 12110 5586 12364 5716
rect 12850 5714 12950 5726
rect 13130 5716 13230 5726
rect 15522 5718 15526 5742
rect 12736 5700 12748 5714
rect 15546 5708 15632 5770
rect 15550 5690 15554 5708
rect 16602 5706 16678 5734
rect 17928 5706 17974 5756
rect 18180 5706 18226 5756
rect 12490 5632 12590 5642
rect 12850 5630 12950 5642
rect 13130 5632 13230 5642
rect 10044 5574 10448 5586
rect 9954 5560 10010 5574
rect 10044 5542 10080 5574
rect 10162 5572 10448 5574
rect 10224 5560 10324 5572
rect 9986 5528 10080 5542
rect 10044 5524 10080 5528
rect 10116 5526 10134 5528
rect 10172 5526 10272 5538
rect 13104 5528 13150 5556
rect 10012 5514 10080 5524
rect 10110 5522 10172 5526
rect 10044 5506 10080 5514
rect 10108 5511 10172 5522
rect 10272 5518 10434 5526
rect 10272 5517 10335 5518
rect 10272 5513 10334 5517
rect 10108 5506 10170 5511
rect 4650 5450 4676 5486
rect 9520 5480 9562 5494
rect 10044 5479 10234 5506
rect 10236 5479 10544 5506
rect 13670 5500 13690 5570
rect 13698 5528 13748 5556
rect 8916 5256 9270 5410
rect 9472 5242 9524 5476
rect 9572 5438 9628 5450
rect 10044 5442 10544 5479
rect 10044 5438 10234 5442
rect 10236 5438 10544 5442
rect 10013 5423 10080 5438
rect 10028 5412 10080 5423
rect 10157 5412 10234 5438
rect 10272 5434 10305 5438
rect 9970 5408 10090 5412
rect 10157 5411 10270 5412
rect 10166 5410 10270 5411
rect 9968 5402 10090 5408
rect 10164 5402 10270 5410
rect 9958 5400 10270 5402
rect 9958 5394 10282 5400
rect 10304 5394 10305 5434
rect 10314 5394 10366 5424
rect 10430 5394 10462 5438
rect 10468 5416 10528 5438
rect 10464 5400 10518 5416
rect 10464 5394 10510 5400
rect 9958 5386 10291 5394
rect 9958 5376 10080 5386
rect 9994 5370 10080 5376
rect 10086 5384 10291 5386
rect 10086 5370 10170 5384
rect 10214 5379 10291 5384
rect 10304 5382 10510 5394
rect 10214 5378 10282 5379
rect 10304 5378 10476 5382
rect 10198 5370 10476 5378
rect 9994 5368 10476 5370
rect 9992 5367 10476 5368
rect 10532 5367 10544 5438
rect 9992 5366 10544 5367
rect 9572 5354 9628 5366
rect 9992 5362 10310 5366
rect 9992 5358 10324 5362
rect 10414 5358 10476 5366
rect 9992 5354 10000 5358
rect 9980 5342 10000 5354
rect 10044 5330 10150 5358
rect 10164 5348 10170 5358
rect 10186 5346 10324 5358
rect 10380 5348 10476 5358
rect 9670 5294 9726 5306
rect 9954 5294 10010 5308
rect 10044 5294 10146 5330
rect 10224 5326 10324 5346
rect 10414 5344 10468 5348
rect 10380 5338 10468 5344
rect 10380 5330 10418 5338
rect 10174 5316 10374 5326
rect 10174 5302 10418 5316
rect 10174 5294 10374 5302
rect 10044 5276 10224 5294
rect 10324 5276 10380 5294
rect 10044 5242 10146 5276
rect 10162 5242 10188 5276
rect 10365 5261 10448 5276
rect 10380 5242 10448 5261
rect 9670 5210 9726 5222
rect 9954 5210 10010 5224
rect 10224 5210 10324 5222
rect 10390 5214 10410 5242
rect 3934 5142 3936 5174
rect 3968 5158 3970 5196
rect 4127 5154 4142 5169
rect 3976 5124 4034 5154
rect 4086 5124 4142 5154
rect 4154 5142 4156 5174
rect 4188 5158 4190 5194
rect 4254 5174 4266 5184
rect 4374 5124 4376 5174
rect 4408 5158 4410 5194
rect 4474 5174 4486 5184
rect 4127 5109 4142 5124
rect 13232 5094 13254 5122
rect 13398 5094 13420 5122
rect 11216 5026 11264 5090
rect 11464 5026 11512 5090
rect 13178 5030 13226 5094
rect 13426 5030 13474 5094
rect 3594 4996 3646 5026
rect 3704 4996 3756 5026
rect 3814 4996 3866 5026
rect 3924 4996 3976 5026
rect 4034 4996 4086 5026
rect 11216 4758 11264 4822
rect 11464 4756 11512 4820
rect 13178 4762 13226 4826
rect 13426 4760 13474 4824
rect 4127 4598 4142 4613
rect 3976 4568 4034 4598
rect 4086 4568 4142 4598
rect 4127 4553 4142 4568
rect 14392 4518 14588 4546
rect 14392 4508 14407 4518
rect 12260 4502 12278 4508
rect 12370 4502 12388 4508
rect 14392 4506 14426 4508
rect 10434 4476 10484 4488
rect 10536 4476 10594 4488
rect 10646 4476 10704 4488
rect 10756 4476 10806 4488
rect 11922 4476 11972 4488
rect 12024 4476 12082 4488
rect 12134 4482 12184 4488
rect 12302 4482 12320 4502
rect 12412 4482 12430 4502
rect 12498 4482 12556 4494
rect 12608 4482 12666 4494
rect 12718 4482 12768 4494
rect 13884 4482 13934 4494
rect 13986 4482 14044 4494
rect 14096 4482 14154 4494
rect 14206 4482 14256 4494
rect 14392 4482 14436 4506
rect 12134 4476 12168 4482
rect 12177 4476 12226 4482
rect 12287 4476 12336 4482
rect 12397 4478 12446 4482
rect 12759 4478 12774 4482
rect 10797 4472 10812 4476
rect 10432 4438 10484 4472
rect 10536 4438 10594 4472
rect 10646 4438 10704 4472
rect 10756 4438 10812 4472
rect 11916 4472 11931 4476
rect 12177 4472 12192 4476
rect 12287 4472 12320 4476
rect 3842 4012 3856 4132
rect 3880 4104 3924 4188
rect 3870 4040 3924 4104
rect 4520 4090 4550 4158
rect 4610 4104 4618 4137
rect 4634 4116 4656 4158
rect 4676 4090 4698 4116
rect 4508 4075 4671 4090
rect 3880 3866 3924 4040
rect 4520 4070 4656 4075
rect 4520 4016 4566 4070
rect 4612 4044 4656 4070
rect 4612 4036 4693 4044
rect 4618 4016 4656 4036
rect 3756 3612 3924 3866
rect 3942 3660 3944 3662
rect 3842 3458 3856 3578
rect 3880 3550 3924 3612
rect 3942 3586 3944 3624
rect 3954 3612 3956 3772
rect 4042 3662 4052 3672
rect 4144 3638 4210 3866
rect 4262 3662 4272 3672
rect 4144 3634 4224 3638
rect 4052 3612 4054 3628
rect 3954 3604 4122 3612
rect 4144 3604 4236 3634
rect 4052 3586 4054 3604
rect 4156 3586 4164 3604
rect 4180 3598 4196 3604
rect 4204 3598 4224 3604
rect 4180 3589 4195 3598
rect 4238 3592 4258 3638
rect 4266 3592 4272 3662
rect 4300 3634 4306 3696
rect 4316 3694 4334 3696
rect 4314 3634 4334 3694
rect 4350 3660 4368 3662
rect 4288 3604 4346 3634
rect 4300 3598 4306 3604
rect 4314 3598 4334 3604
rect 4348 3594 4368 3660
rect 4350 3592 4368 3594
rect 4376 3660 4384 3662
rect 4376 3628 4382 3660
rect 4410 3634 4416 3682
rect 4482 3662 4492 3672
rect 4424 3634 4444 3638
rect 4376 3592 4384 3628
rect 4398 3604 4456 3634
rect 4410 3598 4416 3604
rect 4424 3598 4444 3604
rect 4458 3592 4478 3638
rect 4486 3626 4492 3662
rect 4520 3634 4560 4016
rect 10432 3989 10470 4438
rect 10797 4423 10812 4438
rect 11108 4274 11124 4280
rect 11108 4266 11126 4274
rect 11108 4230 11128 4266
rect 11108 4216 11124 4230
rect 11136 4188 11152 4308
rect 11158 4300 11160 4304
rect 11158 4258 11162 4300
rect 11188 4270 11198 4296
rect 11236 4268 11280 4450
rect 11568 4300 11570 4304
rect 11530 4270 11540 4294
rect 11216 4204 11280 4268
rect 11236 4148 11280 4204
rect 11464 4202 11512 4266
rect 11566 4258 11570 4300
rect 11576 4188 11592 4308
rect 11616 4280 11660 4450
rect 11916 4438 11972 4472
rect 12024 4438 12082 4472
rect 12134 4438 12226 4472
rect 12278 4467 12302 4472
rect 12278 4439 12296 4467
rect 11916 4423 11931 4438
rect 12192 4434 12214 4438
rect 12146 4416 12214 4434
rect 12245 4434 12296 4439
rect 12302 4434 12324 4445
rect 12394 4444 12446 4478
rect 12498 4444 12556 4478
rect 12608 4444 12666 4478
rect 12718 4444 12774 4478
rect 13878 4478 13893 4482
rect 12245 4428 12324 4434
rect 12355 4434 12388 4439
rect 12394 4434 12434 4444
rect 12355 4428 12434 4434
rect 12465 4434 12498 4439
rect 12465 4428 12544 4434
rect 12759 4429 12774 4444
rect 12146 4400 12225 4416
rect 12256 4400 12324 4428
rect 12366 4400 12434 4428
rect 12476 4400 12544 4428
rect 12146 4394 12180 4400
rect 12256 4394 12296 4400
rect 12366 4394 12432 4400
rect 12476 4394 12510 4400
rect 12192 4366 12225 4377
rect 12278 4371 12296 4394
rect 12394 4377 12432 4394
rect 12146 4364 12225 4366
rect 12245 4366 12296 4371
rect 12302 4366 12324 4377
rect 12146 4332 12214 4364
rect 12245 4360 12324 4366
rect 12355 4366 12388 4371
rect 12394 4366 12434 4377
rect 12355 4360 12434 4366
rect 12465 4366 12498 4371
rect 12465 4360 12544 4366
rect 12256 4332 12324 4360
rect 12366 4332 12434 4360
rect 12476 4332 12544 4360
rect 12146 4326 12180 4332
rect 12256 4326 12296 4332
rect 12366 4326 12432 4332
rect 12476 4326 12510 4332
rect 12192 4298 12214 4309
rect 12278 4303 12296 4326
rect 12394 4309 12432 4326
rect 11604 4274 11660 4280
rect 11602 4266 11660 4274
rect 11600 4230 11660 4266
rect 12146 4264 12214 4298
rect 12245 4298 12296 4303
rect 12302 4298 12324 4309
rect 12245 4292 12324 4298
rect 12355 4298 12388 4303
rect 12394 4298 12434 4309
rect 12355 4292 12434 4298
rect 12465 4298 12498 4303
rect 12465 4292 12544 4298
rect 12256 4264 12324 4292
rect 12366 4264 12434 4292
rect 12476 4264 12544 4292
rect 13070 4280 13086 4286
rect 13070 4272 13088 4280
rect 12146 4258 12180 4264
rect 12256 4258 12296 4264
rect 12366 4258 12432 4264
rect 12476 4258 12510 4264
rect 12192 4230 12214 4241
rect 12278 4235 12296 4258
rect 12394 4241 12432 4258
rect 11604 4216 11660 4230
rect 11616 4148 11660 4216
rect 12146 4196 12214 4230
rect 12245 4230 12296 4235
rect 12302 4230 12324 4241
rect 12245 4224 12324 4230
rect 12355 4230 12388 4235
rect 12394 4230 12434 4241
rect 13070 4236 13090 4272
rect 12355 4224 12434 4230
rect 12465 4230 12498 4235
rect 12465 4224 12544 4230
rect 12256 4196 12324 4224
rect 12366 4196 12434 4224
rect 12476 4196 12544 4224
rect 13070 4222 13086 4236
rect 12146 4190 12180 4196
rect 12256 4190 12296 4196
rect 12366 4190 12432 4196
rect 12476 4190 12510 4196
rect 13098 4194 13114 4314
rect 13120 4306 13122 4310
rect 13120 4264 13124 4306
rect 13150 4276 13160 4300
rect 13198 4272 13242 4456
rect 13530 4306 13532 4310
rect 13492 4276 13502 4300
rect 13178 4208 13242 4272
rect 13426 4208 13474 4272
rect 13528 4264 13532 4306
rect 12192 4162 12214 4173
rect 12278 4167 12296 4190
rect 12394 4173 12432 4190
rect 10426 3978 10484 3989
rect 10264 3948 10316 3978
rect 10374 3974 10536 3978
rect 10374 3948 10426 3974
rect 10432 3936 10470 3974
rect 10484 3948 10536 3974
rect 10594 3948 10646 3978
rect 10704 3948 10756 3978
rect 10592 3936 10600 3938
rect 10782 3936 10848 4148
rect 11036 3936 11038 4054
rect 11112 4012 11280 4148
rect 11108 3948 11280 4012
rect 11112 3936 11280 3948
rect 10432 3914 10468 3936
rect 10484 3914 10512 3936
rect 10592 3918 11280 3936
rect 10432 3910 10512 3914
rect 10426 3896 10484 3910
rect 10500 3896 10506 3910
rect 10514 3896 10534 3912
rect 10536 3910 10594 3914
rect 10564 3908 10572 3910
rect 10610 3908 10616 3912
rect 10624 3908 10644 3912
rect 10646 3910 10704 3914
rect 10720 3908 10726 3918
rect 10734 3908 10754 3918
rect 10782 3914 10848 3918
rect 10756 3910 10848 3914
rect 10782 3908 10848 3910
rect 10862 3908 10864 3912
rect 10972 3908 10974 3912
rect 11036 3908 11038 3918
rect 11082 3908 11084 3912
rect 11112 3908 11280 3918
rect 10564 3900 11280 3908
rect 10548 3896 11280 3900
rect 10426 3895 11280 3896
rect 4486 3592 4494 3626
rect 4508 3604 4560 3634
rect 4520 3603 4560 3604
rect 10432 3894 10472 3895
rect 10478 3894 11280 3895
rect 11492 4042 11660 4148
rect 11690 4042 11692 4054
rect 11880 4042 11946 4148
rect 12146 4128 12214 4162
rect 12245 4162 12296 4167
rect 12302 4162 12324 4173
rect 12245 4156 12324 4162
rect 12355 4162 12388 4167
rect 12394 4162 12434 4173
rect 12355 4156 12434 4162
rect 12465 4162 12498 4167
rect 12465 4156 12544 4162
rect 12256 4128 12324 4156
rect 12366 4128 12434 4156
rect 12476 4128 12544 4156
rect 13198 4154 13242 4208
rect 13538 4194 13554 4314
rect 13578 4286 13622 4456
rect 13878 4444 13934 4478
rect 13986 4444 14044 4478
rect 14096 4444 14154 4478
rect 14206 4444 14258 4478
rect 14392 4471 14484 4482
rect 14391 4460 14484 4471
rect 13878 4429 13893 4444
rect 13566 4280 13622 4286
rect 13564 4272 13622 4280
rect 13562 4236 13622 4272
rect 13566 4222 13622 4236
rect 13578 4154 13622 4222
rect 12146 4122 12180 4128
rect 12256 4122 12296 4128
rect 12366 4122 12432 4128
rect 12476 4122 12510 4128
rect 12192 4094 12214 4105
rect 12278 4099 12296 4122
rect 12394 4105 12432 4122
rect 12146 4060 12214 4094
rect 12245 4094 12296 4099
rect 12302 4094 12324 4105
rect 12245 4088 12324 4094
rect 12355 4094 12388 4099
rect 12394 4094 12434 4105
rect 12355 4088 12434 4094
rect 12465 4094 12498 4099
rect 12465 4088 12544 4094
rect 12256 4060 12324 4088
rect 12366 4060 12434 4088
rect 12476 4060 12544 4088
rect 12146 4054 12180 4060
rect 12256 4054 12296 4060
rect 12366 4054 12432 4060
rect 12476 4054 12510 4060
rect 11492 4016 11698 4042
rect 11800 4016 11946 4042
rect 12018 4016 12136 4042
rect 12192 4026 12214 4037
rect 12278 4031 12296 4054
rect 12394 4037 12432 4054
rect 11492 4014 11660 4016
rect 11492 3988 11670 4014
rect 11492 3936 11660 3988
rect 11690 3936 11692 4016
rect 11880 4014 11946 4016
rect 11828 3988 11946 4014
rect 12046 3988 12108 4014
rect 12146 3992 12214 4026
rect 12245 4026 12296 4031
rect 12302 4026 12324 4037
rect 12245 4020 12324 4026
rect 12355 4026 12388 4031
rect 12394 4026 12434 4037
rect 12355 4020 12434 4026
rect 12465 4026 12498 4031
rect 12465 4020 12544 4026
rect 12256 3992 12324 4020
rect 12366 3992 12434 4020
rect 12476 4018 12544 4020
rect 12744 4018 12810 4154
rect 12998 4018 13000 4060
rect 13074 4018 13242 4154
rect 12476 4016 12582 4018
rect 12644 4016 12810 4018
rect 12862 4016 13020 4018
rect 12476 3992 12544 4016
rect 11880 3936 11946 3988
rect 12146 3986 12180 3992
rect 12256 3989 12296 3992
rect 12256 3986 12302 3989
rect 12366 3986 12432 3992
rect 12476 3986 12510 3992
rect 12744 3990 12810 4016
rect 12998 3990 13000 4016
rect 12554 3988 12582 3990
rect 12644 3988 12810 3990
rect 12862 3988 13020 3990
rect 12278 3984 12302 3986
rect 12388 3984 12432 3986
rect 12498 3984 12513 3986
rect 12192 3980 12258 3984
rect 12278 3980 12513 3984
rect 11972 3948 12024 3978
rect 12082 3948 12134 3978
rect 12192 3974 12513 3980
rect 12192 3954 12258 3974
rect 12260 3954 12296 3974
rect 12192 3948 12244 3954
rect 12258 3948 12296 3954
rect 12302 3954 12388 3974
rect 12394 3954 12498 3974
rect 12556 3954 12608 3984
rect 12666 3954 12718 3984
rect 12302 3948 12354 3954
rect 12394 3948 12464 3954
rect 12260 3936 12296 3948
rect 12394 3942 12432 3948
rect 12336 3936 12338 3942
rect 11492 3918 12136 3936
rect 11492 3908 11660 3918
rect 11678 3908 11680 3912
rect 11690 3908 11692 3918
rect 11880 3914 11946 3918
rect 11788 3908 11790 3912
rect 11880 3910 11972 3914
rect 11880 3908 11946 3910
rect 11974 3908 11994 3918
rect 12002 3908 12008 3918
rect 12302 3916 12338 3936
rect 12394 3916 12430 3942
rect 12446 3936 12474 3942
rect 12744 3936 12810 3988
rect 12998 3936 13000 3988
rect 13070 3954 13242 4018
rect 13074 3936 13242 3954
rect 12554 3924 13242 3936
rect 12024 3910 12082 3914
rect 12086 3908 12104 3912
rect 12112 3908 12120 3912
rect 12134 3910 12168 3914
rect 12177 3912 12226 3916
rect 12177 3910 12230 3912
rect 11492 3894 12164 3908
rect 12177 3901 12192 3910
rect 12222 3906 12230 3910
rect 12278 3910 12336 3916
rect 12388 3910 12446 3916
rect 12222 3894 12228 3906
rect 12278 3901 12302 3910
rect 12388 3906 12432 3910
rect 12388 3901 12434 3906
rect 10432 3890 11280 3894
rect 10432 3864 10594 3890
rect 10610 3872 10616 3890
rect 4508 3592 4566 3603
rect 4236 3588 4288 3592
rect 4346 3588 4398 3592
rect 4456 3588 4618 3592
rect 4186 3584 4560 3588
rect 4236 3562 4288 3584
rect 4346 3562 4398 3584
rect 4456 3562 4508 3584
rect 3870 3486 3924 3550
rect 4522 3550 4560 3584
rect 4566 3562 4618 3588
rect 4676 3562 4728 3592
rect 3934 3514 4092 3534
rect 4154 3514 4310 3534
rect 4372 3514 4400 3534
rect 4522 3524 4550 3550
rect 4566 3524 4602 3550
rect 4508 3509 4566 3524
rect 3934 3486 4092 3506
rect 4154 3486 4310 3506
rect 4372 3486 4428 3506
rect 3830 3198 3834 3240
rect 3832 3194 3834 3198
rect 3840 3190 3856 3310
rect 3880 3282 3924 3486
rect 3868 3268 3924 3282
rect 3864 3232 3924 3268
rect 3866 3224 3924 3232
rect 3868 3218 3924 3224
rect 3880 3048 3924 3218
rect 4180 3060 4195 3075
rect 4522 3060 4560 3509
rect 10299 3482 10426 3509
rect 10432 3482 10472 3864
rect 10478 3804 10570 3864
rect 10576 3816 10582 3864
rect 10608 3838 10616 3872
rect 10610 3836 10616 3838
rect 10624 3836 10644 3890
rect 10646 3864 10704 3890
rect 10658 3804 10678 3864
rect 10658 3802 10676 3804
rect 10686 3802 10692 3864
rect 10720 3836 10726 3890
rect 10734 3870 10754 3890
rect 10756 3870 10812 3890
rect 10830 3872 10836 3890
rect 11036 3886 11280 3890
rect 10734 3864 10812 3870
rect 10734 3860 10764 3864
rect 10768 3860 10788 3864
rect 10796 3849 10812 3864
rect 10796 3816 10802 3849
rect 10828 3838 10836 3872
rect 10974 3860 10984 3870
rect 11048 3838 11050 3852
rect 10830 3836 10836 3838
rect 10862 3836 10864 3838
rect 11082 3836 11084 3838
rect 10299 3462 10472 3482
rect 10336 3441 10472 3462
rect 10301 3423 10472 3441
rect 10301 3408 10484 3423
rect 10336 3382 10358 3408
rect 10484 3382 10514 3408
rect 11108 3394 11122 3458
rect 11136 3366 11150 3486
rect 11236 3310 11280 3886
rect 11616 3890 12228 3894
rect 11578 3366 11592 3486
rect 11616 3458 11660 3890
rect 11690 3886 11858 3890
rect 11880 3886 11972 3890
rect 11892 3872 11898 3886
rect 11744 3860 11754 3870
rect 11678 3836 11680 3852
rect 11892 3836 11900 3872
rect 11916 3870 11972 3886
rect 11974 3870 11994 3890
rect 11916 3864 11994 3870
rect 11916 3849 11932 3864
rect 11940 3860 11960 3864
rect 11964 3860 11994 3864
rect 11926 3816 11932 3849
rect 12002 3836 12008 3890
rect 12024 3864 12082 3890
rect 12036 3802 12042 3864
rect 12050 3804 12070 3864
rect 12084 3838 12104 3890
rect 12086 3836 12104 3838
rect 12112 3872 12118 3890
rect 12112 3836 12120 3872
rect 12134 3864 12228 3890
rect 12256 3873 12262 3900
rect 12278 3873 12296 3901
rect 12394 3900 12434 3901
rect 12146 3836 12228 3864
rect 12245 3868 12296 3873
rect 12302 3868 12324 3879
rect 12245 3862 12324 3868
rect 12355 3868 12388 3873
rect 12394 3870 12446 3900
rect 12462 3873 12468 3918
rect 12476 3900 12496 3918
rect 12498 3916 12556 3920
rect 12572 3908 12578 3918
rect 12586 3908 12606 3918
rect 12608 3916 12666 3920
rect 12682 3908 12688 3924
rect 12696 3908 12716 3924
rect 12744 3920 12810 3924
rect 12718 3916 12810 3920
rect 12744 3908 12810 3916
rect 12824 3910 12826 3918
rect 12934 3910 12936 3918
rect 12998 3908 13000 3924
rect 13044 3914 13046 3918
rect 13074 3908 13242 3924
rect 12526 3906 13242 3908
rect 12510 3900 13242 3906
rect 13454 3936 13622 4154
rect 13652 3936 13654 4060
rect 13842 3936 13908 4154
rect 14220 3995 14258 4444
rect 14392 4403 14484 4460
rect 14391 4392 14484 4403
rect 14392 4335 14484 4392
rect 14391 4324 14484 4335
rect 14392 4267 14484 4324
rect 14391 4256 14484 4267
rect 14392 4199 14484 4256
rect 14391 4188 14484 4199
rect 14392 4131 14484 4188
rect 14391 4120 14484 4131
rect 14392 4058 14484 4120
rect 14520 4058 14588 4518
rect 14981 4444 14996 4459
rect 14830 4414 14888 4444
rect 14940 4414 14996 4444
rect 14981 4399 14996 4414
rect 14392 4054 14610 4058
rect 14438 4030 14520 4054
rect 14448 4028 14520 4030
rect 14558 4028 14610 4054
rect 14668 4028 14720 4058
rect 14778 4028 14830 4058
rect 14888 4028 14940 4058
rect 14469 4022 14520 4028
rect 14206 3984 14264 3995
rect 14438 3990 14520 4022
rect 14392 3984 14484 3990
rect 13934 3954 13986 3984
rect 14044 3954 14096 3984
rect 14154 3980 14316 3984
rect 14154 3954 14206 3980
rect 14220 3942 14258 3980
rect 14264 3954 14316 3980
rect 14374 3980 14484 3984
rect 14374 3954 14436 3980
rect 14438 3974 14470 3980
rect 13454 3924 14098 3936
rect 13454 3908 13622 3924
rect 13640 3914 13642 3918
rect 13652 3908 13654 3924
rect 13842 3920 13908 3924
rect 13750 3910 13752 3918
rect 13842 3916 13934 3920
rect 13842 3908 13908 3916
rect 13936 3908 13956 3924
rect 13964 3908 13970 3924
rect 14220 3920 14248 3942
rect 13986 3916 14044 3920
rect 14048 3910 14066 3918
rect 14046 3908 14066 3910
rect 14074 3910 14082 3918
rect 14096 3916 14154 3920
rect 14158 3912 14176 3918
rect 14074 3908 14080 3910
rect 13454 3906 14126 3908
rect 13454 3900 14142 3906
rect 12498 3896 13242 3900
rect 12498 3873 12556 3896
rect 12572 3878 12578 3896
rect 12462 3870 12556 3873
rect 12394 3868 12434 3870
rect 12355 3862 12434 3868
rect 12146 3834 12225 3836
rect 12256 3834 12324 3862
rect 12146 3828 12180 3834
rect 12256 3828 12296 3834
rect 12366 3828 12434 3862
rect 12462 3868 12498 3870
rect 12538 3868 12544 3870
rect 12462 3862 12544 3868
rect 12462 3842 12468 3862
rect 12476 3834 12544 3862
rect 12570 3844 12578 3878
rect 12572 3842 12578 3844
rect 12586 3842 12606 3896
rect 12608 3870 12666 3896
rect 12476 3828 12510 3834
rect 12146 3816 12152 3828
rect 12052 3802 12070 3804
rect 12192 3800 12214 3811
rect 12256 3805 12262 3828
rect 12278 3805 12296 3828
rect 12146 3766 12214 3800
rect 12245 3800 12296 3805
rect 12302 3800 12324 3811
rect 12245 3794 12324 3800
rect 12355 3800 12388 3805
rect 12394 3800 12434 3828
rect 12538 3822 12544 3834
rect 12620 3810 12640 3870
rect 12620 3808 12638 3810
rect 12648 3808 12654 3870
rect 12682 3842 12688 3896
rect 12696 3876 12716 3896
rect 12718 3876 12774 3896
rect 12792 3878 12798 3896
rect 12998 3892 13242 3896
rect 12696 3870 12774 3876
rect 12696 3866 12726 3870
rect 12730 3866 12750 3870
rect 12758 3855 12774 3870
rect 12758 3822 12764 3855
rect 12790 3844 12798 3878
rect 12936 3866 12946 3876
rect 13010 3844 13012 3858
rect 12792 3842 12798 3844
rect 12824 3842 12826 3844
rect 13044 3842 13046 3844
rect 12355 3794 12434 3800
rect 12465 3800 12498 3805
rect 12465 3794 12544 3800
rect 12256 3766 12324 3794
rect 12146 3760 12180 3766
rect 12256 3760 12296 3766
rect 12366 3760 12434 3794
rect 12476 3766 12544 3794
rect 12476 3760 12510 3766
rect 12192 3732 12214 3743
rect 12278 3737 12296 3760
rect 12146 3698 12214 3732
rect 12245 3732 12296 3737
rect 12302 3732 12324 3743
rect 12245 3726 12324 3732
rect 12355 3732 12388 3737
rect 12394 3732 12434 3760
rect 12355 3726 12434 3732
rect 12465 3732 12498 3737
rect 12465 3726 12544 3732
rect 12256 3698 12324 3726
rect 12146 3692 12180 3698
rect 12256 3692 12296 3698
rect 12366 3692 12434 3726
rect 12476 3698 12544 3726
rect 12476 3692 12510 3698
rect 12192 3664 12214 3675
rect 12278 3669 12296 3692
rect 12146 3630 12214 3664
rect 12245 3664 12296 3669
rect 12302 3664 12324 3675
rect 12245 3658 12324 3664
rect 12355 3664 12388 3669
rect 12394 3664 12434 3692
rect 12355 3658 12434 3664
rect 12465 3664 12498 3669
rect 12465 3658 12544 3664
rect 12256 3630 12324 3658
rect 12146 3624 12180 3630
rect 12256 3624 12296 3630
rect 12366 3624 12434 3658
rect 12476 3630 12544 3658
rect 12476 3624 12510 3630
rect 12148 3614 12246 3622
rect 12154 3608 12246 3614
rect 12192 3596 12214 3607
rect 12278 3601 12296 3624
rect 12146 3594 12214 3596
rect 12245 3596 12296 3601
rect 12302 3596 12324 3607
rect 12146 3586 12220 3594
rect 12245 3590 12324 3596
rect 12355 3596 12388 3601
rect 12394 3596 12434 3624
rect 12355 3590 12434 3596
rect 12465 3596 12498 3601
rect 12465 3590 12544 3596
rect 12146 3562 12225 3586
rect 12256 3562 12324 3590
rect 12146 3556 12180 3562
rect 12256 3556 12296 3562
rect 12366 3556 12434 3590
rect 12476 3562 12544 3590
rect 12476 3556 12510 3562
rect 12192 3528 12214 3539
rect 12278 3533 12296 3556
rect 12146 3494 12214 3528
rect 12245 3528 12296 3533
rect 12302 3528 12324 3539
rect 12245 3522 12324 3528
rect 12355 3528 12388 3533
rect 12394 3528 12434 3556
rect 12355 3522 12434 3528
rect 12465 3528 12498 3533
rect 12465 3522 12544 3528
rect 12256 3515 12324 3522
rect 12366 3515 12434 3522
rect 12256 3500 12434 3515
rect 12256 3498 12446 3500
rect 12146 3488 12180 3494
rect 12256 3488 12448 3498
rect 12476 3494 12544 3522
rect 12476 3488 12510 3494
rect 12192 3460 12214 3471
rect 12261 3468 12448 3488
rect 12278 3465 12448 3468
rect 11606 3394 11660 3458
rect 12146 3426 12214 3460
rect 12245 3454 12448 3465
rect 12465 3460 12498 3465
rect 12528 3460 12582 3464
rect 12465 3454 12582 3460
rect 12256 3430 12448 3454
rect 12476 3452 12582 3454
rect 12644 3452 12800 3464
rect 12862 3452 13020 3464
rect 12146 3420 12180 3426
rect 12256 3420 12434 3430
rect 12476 3426 12550 3452
rect 12476 3420 12510 3426
rect 12556 3424 12582 3436
rect 12644 3424 12800 3436
rect 12862 3424 13020 3436
rect 12263 3414 12434 3420
rect 12498 3414 12513 3420
rect 12244 3408 12427 3414
rect 12464 3408 12513 3414
rect 12328 3400 12334 3408
rect 12356 3406 12362 3408
rect 12406 3406 12420 3408
rect 12310 3398 12344 3400
rect 12556 3398 12578 3424
rect 13070 3400 13084 3464
rect 12312 3394 12344 3398
rect 11616 3310 11660 3394
rect 12256 3382 12286 3388
rect 12330 3332 12332 3370
rect 12346 3360 12378 3394
rect 13098 3372 13112 3492
rect 12312 3326 12344 3332
rect 12358 3326 12360 3360
rect 12330 3306 12332 3326
rect 12346 3298 12378 3326
rect 13198 3316 13242 3892
rect 13578 3896 14154 3900
rect 13540 3372 13554 3492
rect 13578 3464 13622 3896
rect 13652 3892 13820 3896
rect 13842 3892 13934 3896
rect 13854 3878 13860 3892
rect 13706 3866 13716 3876
rect 13640 3842 13642 3858
rect 13854 3842 13862 3878
rect 13878 3876 13934 3892
rect 13936 3876 13956 3896
rect 13878 3870 13956 3876
rect 13878 3855 13894 3870
rect 13902 3866 13922 3870
rect 13926 3866 13956 3870
rect 13888 3822 13894 3855
rect 13964 3842 13970 3896
rect 13986 3870 14044 3896
rect 13998 3808 14004 3870
rect 14012 3810 14032 3870
rect 14046 3844 14066 3896
rect 14048 3842 14066 3844
rect 14074 3878 14080 3896
rect 14074 3842 14082 3878
rect 14096 3876 14154 3896
rect 14156 3876 14176 3912
rect 14096 3870 14176 3876
rect 14108 3822 14114 3870
rect 14122 3866 14142 3870
rect 14146 3866 14176 3870
rect 14184 3912 14192 3918
rect 14206 3916 14256 3920
rect 14264 3916 14300 3942
rect 14392 3916 14436 3954
rect 14184 3842 14190 3912
rect 14206 3901 14264 3916
rect 14392 3915 14484 3916
rect 14391 3904 14484 3915
rect 14218 3900 14258 3901
rect 14206 3870 14258 3900
rect 14014 3808 14032 3810
rect 14218 3488 14258 3870
rect 14392 3847 14484 3904
rect 14391 3836 14484 3847
rect 14392 3779 14484 3836
rect 14391 3768 14484 3779
rect 14392 3711 14484 3768
rect 14391 3700 14484 3711
rect 14392 3643 14484 3700
rect 14391 3632 14484 3643
rect 14392 3575 14484 3632
rect 14391 3564 14484 3575
rect 14264 3488 14391 3515
rect 14392 3499 14484 3564
rect 14520 3499 14588 3990
rect 14726 3920 15246 3936
rect 14726 3892 15274 3908
rect 14981 3888 14996 3892
rect 14788 3838 14790 3870
rect 14830 3858 14888 3888
rect 14940 3858 14996 3888
rect 14822 3816 14824 3854
rect 14981 3843 14996 3858
rect 15008 3838 15010 3870
rect 15074 3862 15086 3872
rect 15042 3818 15044 3854
rect 15228 3838 15230 3888
rect 15294 3862 15306 3872
rect 15262 3818 15264 3854
rect 14392 3498 14588 3499
rect 14218 3474 14391 3488
rect 14438 3474 14484 3498
rect 14218 3468 14410 3474
rect 14448 3472 14484 3474
rect 13568 3400 13622 3464
rect 13632 3452 13790 3464
rect 13852 3452 14008 3464
rect 14070 3452 14124 3464
rect 14218 3447 14264 3468
rect 14296 3452 14410 3468
rect 14469 3460 14484 3472
rect 14472 3457 14484 3460
rect 14780 3452 14938 3460
rect 15000 3452 15156 3460
rect 15218 3452 15272 3460
rect 15444 3452 15558 3470
rect 14310 3447 14354 3452
rect 13632 3424 13790 3436
rect 13852 3424 14008 3436
rect 14070 3424 14096 3436
rect 14218 3429 14389 3447
rect 14206 3414 14389 3429
rect 14780 3424 14938 3432
rect 15000 3424 15156 3432
rect 15218 3424 15244 3432
rect 15444 3424 15530 3442
rect 13578 3316 13622 3400
rect 14218 3388 14248 3414
rect 14374 3388 14396 3414
rect 14082 3370 14096 3388
rect 14232 3376 14242 3378
rect 14110 3346 14124 3360
rect 14204 3358 14214 3360
rect 14202 3356 14214 3358
rect 14230 3356 14242 3376
rect 14656 3368 15244 3384
rect 14702 3366 15244 3368
rect 14110 3342 14118 3346
rect 14202 3284 14212 3356
rect 14230 3312 14240 3356
rect 14628 3340 15272 3356
rect 14674 3338 15272 3340
rect 21112 3328 21344 3398
rect 4744 3138 4774 3154
rect 4786 3138 4822 3164
rect 4180 3026 4236 3060
rect 4288 3026 4346 3060
rect 4398 3026 4456 3060
rect 4508 3026 4560 3060
rect 4722 3120 4786 3138
rect 4722 3070 4808 3120
rect 4722 3036 4786 3070
rect 4180 3022 4195 3026
rect 4724 3022 4786 3036
rect 4186 3010 4236 3022
rect 4288 3010 4346 3022
rect 4398 3010 4456 3022
rect 4508 3010 4558 3022
rect 4724 2996 4728 3022
rect 4724 2985 4735 2996
rect 4822 2986 4848 3138
rect 20920 3074 21090 3328
rect 21112 3076 21880 3328
rect 21884 3200 21890 3278
rect 21992 3200 21998 3278
rect 22076 3200 22082 3278
rect 20960 2878 20966 2956
rect 21044 2878 21050 2956
rect 20960 2556 20966 2634
rect 21044 2556 21050 2634
rect 20960 2234 20966 2312
rect 21044 2234 21050 2312
rect 20798 1970 20806 2066
rect 20826 1998 20834 2038
rect 20960 1912 20966 1990
rect 21044 1912 21050 1990
rect 20920 1810 20992 1822
rect 20882 1790 20904 1794
rect 20880 1760 20904 1790
rect 20910 1762 20932 1766
rect 20908 1760 20932 1762
rect 20920 1684 21090 1720
rect 20882 1652 20904 1684
rect 20910 1680 21090 1684
rect 20920 1478 21090 1680
rect 21112 1718 21344 3074
rect 21416 2896 21422 2952
rect 21394 2874 21422 2896
rect 21500 2874 21506 2952
rect 21608 2874 21614 2952
rect 21692 2874 21698 2952
rect 21800 2874 21806 2952
rect 21884 2874 21890 2952
rect 21992 2878 21998 2956
rect 22076 2878 22082 2956
rect 21394 2862 21416 2874
rect 21428 2828 21450 2862
rect 21620 2828 21686 2830
rect 21626 2794 21664 2796
rect 21590 2758 21620 2764
rect 21488 2642 21494 2666
rect 21416 2552 21422 2630
rect 21488 2608 21528 2632
rect 21500 2552 21506 2608
rect 21608 2552 21614 2630
rect 21692 2552 21698 2630
rect 21800 2552 21806 2630
rect 21884 2552 21890 2630
rect 21992 2556 21998 2634
rect 22076 2556 22082 2634
rect 21640 2362 21652 2372
rect 21668 2362 21680 2400
rect 21598 2328 21606 2350
rect 21614 2313 21621 2362
rect 21640 2350 21692 2362
rect 21640 2347 21724 2350
rect 21640 2342 21652 2347
rect 21658 2334 21724 2347
rect 21760 2334 21766 2378
rect 21677 2319 21692 2334
rect 21416 2230 21422 2308
rect 21500 2230 21506 2308
rect 21608 2230 21614 2308
rect 21692 2230 21698 2308
rect 21800 2230 21806 2308
rect 21884 2230 21890 2308
rect 21992 2234 21998 2312
rect 22076 2234 22082 2312
rect 21422 2176 21441 2184
rect 21408 2128 21410 2150
rect 21358 2096 21410 2128
rect 21442 2116 21444 2184
rect 21440 1908 21446 1986
rect 21524 1908 21530 1986
rect 21568 1908 21592 2028
rect 21598 2006 21608 2028
rect 21614 1991 21623 2040
rect 21643 2028 21692 2040
rect 21643 2025 21724 2028
rect 21658 2012 21724 2025
rect 21760 2012 21766 2056
rect 21677 1997 21692 2012
rect 21608 1908 21614 1986
rect 21692 1908 21698 1986
rect 21800 1908 21806 1986
rect 21884 1908 21890 1986
rect 21992 1912 21998 1990
rect 22076 1912 22082 1990
rect 21465 1880 21524 1889
rect 21462 1854 21524 1880
rect 21462 1770 21488 1854
rect 21496 1804 21522 1846
rect 21568 1838 21598 1900
rect 21568 1834 21604 1838
rect 21568 1832 21676 1834
rect 21546 1808 21562 1816
rect 21568 1808 21688 1832
rect 21760 1808 21832 1818
rect 21952 1810 22024 1822
rect 21542 1792 21562 1808
rect 21584 1790 21612 1792
rect 21614 1790 21642 1792
rect 21584 1786 21600 1790
rect 21614 1786 21668 1790
rect 21584 1762 21800 1786
rect 21596 1730 21800 1762
rect 21596 1720 21846 1730
rect 21112 1506 21474 1718
rect 21488 1644 21546 1718
rect 21596 1644 22122 1720
rect 21488 1506 22122 1644
rect 21112 1498 22122 1506
rect 21112 1476 21474 1498
rect 21488 1488 22122 1498
rect 20920 1464 21090 1466
rect 21488 1464 21642 1488
rect 21688 1478 22122 1488
rect 21688 1476 21930 1478
rect 20960 1268 20966 1346
rect 21044 1268 21050 1346
rect 20960 946 20966 1024
rect 21044 946 21050 1024
rect 20960 624 20966 702
rect 21044 624 21050 702
rect 20960 302 20966 380
rect 21044 302 21050 380
rect 21112 178 21344 1464
rect 21598 1362 21606 1384
rect 21614 1347 21621 1396
rect 21643 1384 21692 1396
rect 21643 1381 21724 1384
rect 21658 1366 21724 1381
rect 21760 1366 21766 1412
rect 21677 1351 21692 1366
rect 21416 1264 21422 1342
rect 21500 1264 21506 1342
rect 21608 1264 21614 1342
rect 21692 1264 21698 1342
rect 21800 1264 21806 1342
rect 21884 1264 21890 1342
rect 21992 1268 21998 1346
rect 22076 1268 22082 1346
rect 21598 1040 21604 1062
rect 21614 1025 21619 1074
rect 21641 1062 21692 1074
rect 21641 1059 21722 1062
rect 21656 1044 21722 1059
rect 21760 1044 21764 1090
rect 21677 1029 21692 1044
rect 21416 942 21422 1020
rect 21500 942 21506 1020
rect 21608 942 21614 1020
rect 21692 942 21698 1020
rect 21800 942 21806 1020
rect 21884 942 21890 1020
rect 21992 946 21998 1024
rect 22076 946 22082 1024
rect 22666 930 22668 1004
rect 21568 842 21622 848
rect 21530 768 21547 790
rect 21474 764 21594 768
rect 21492 740 21494 744
rect 21499 740 21500 752
rect 21514 750 21578 764
rect 21526 740 21528 750
rect 21474 736 21566 740
rect 21486 722 21566 736
rect 21492 710 21494 722
rect 21526 720 21528 722
rect 21416 620 21422 698
rect 21500 620 21506 698
rect 21608 620 21614 698
rect 21692 620 21698 698
rect 21800 620 21806 698
rect 21884 620 21890 698
rect 21992 624 21998 702
rect 22076 624 22082 702
rect 21376 520 21448 522
rect 21568 520 21640 522
rect 21760 520 21832 522
rect 21598 396 21604 422
rect 21614 381 21619 432
rect 21641 422 21692 432
rect 21641 417 21722 422
rect 21656 404 21722 417
rect 21760 404 21764 450
rect 21677 389 21692 404
rect 21416 302 21422 380
rect 21500 302 21506 380
rect 21608 302 21614 380
rect 21692 302 21698 380
rect 21800 302 21806 380
rect 21884 302 21890 380
rect 21992 302 21998 380
rect 22076 302 22082 380
<< nwell >>
rect 11898 10808 11904 10810
rect 8946 10780 9300 10802
rect 10074 10780 10574 10802
rect 11762 10748 11904 10808
rect 11762 10740 11898 10748
rect 11760 9530 11900 10740
rect 13854 10322 13856 10560
rect 13854 10312 13864 10322
rect 13854 10292 13866 10312
rect 13856 10068 13866 10292
rect 16540 10110 16652 10218
rect 11762 9490 11900 9530
rect 11760 5586 12110 6780
rect 11760 5580 12364 5586
rect 12188 5548 12364 5580
rect 12140 4154 12544 5292
rect 22668 930 22938 4024
rect 22666 836 22938 930
<< psubdiff >>
rect 2432 12494 6036 12520
rect 2432 12352 5176 12494
rect 5354 12352 6036 12494
rect 2432 12338 6036 12352
rect 5854 4878 6036 12338
rect 14644 11884 17866 11894
rect 14644 11720 14670 11884
rect 14722 11882 17866 11884
rect 14722 11726 17336 11882
rect 17514 11726 17866 11882
rect 14722 11720 17866 11726
rect 14644 11712 17866 11720
rect 17684 8074 17866 11712
rect 5854 4810 5876 4878
rect 5910 4844 5944 4878
rect 5978 4844 6036 4878
rect 6012 4810 6036 4844
rect 5854 4774 6036 4810
rect 5854 4652 5882 4774
rect 5988 4652 6036 4774
rect 4722 3120 5224 3138
rect 4722 3036 4778 3120
rect 4724 2416 4778 3036
rect 4812 2416 4850 3120
rect 4884 2416 4920 3120
rect 4954 2416 4990 3120
rect 5024 2416 5062 3120
rect 5096 2416 5132 3120
rect 5166 2416 5224 3120
rect 4724 2390 5224 2416
rect 5854 2552 6036 4652
rect 17186 7892 17866 8074
rect 17186 2552 17368 7892
rect 4724 2388 4794 2390
rect 5854 2370 20170 2552
rect 5854 1576 6036 2370
<< nsubdiff >>
rect 22750 3962 22864 3978
rect 22750 3174 22776 3962
rect 22758 3054 22776 3174
rect 22750 2852 22776 3054
rect 22758 2732 22776 2852
rect 22750 2530 22776 2732
rect 22756 2410 22776 2530
rect 22750 2206 22776 2410
rect 22758 2086 22776 2206
rect 22750 1884 22776 2086
rect 22756 1764 22776 1884
rect 22750 1390 22776 1764
rect 22756 972 22776 1390
rect 22810 972 22864 3962
rect 22756 948 22864 972
<< psubdiffcont >>
rect 5176 12352 5354 12494
rect 14670 11720 14722 11884
rect 17336 11726 17514 11882
rect 5876 4844 5910 4878
rect 5944 4844 5978 4878
rect 5876 4810 6012 4844
rect 5882 4652 5988 4774
rect 4778 2416 4812 3120
rect 4850 2416 4884 3120
rect 4920 2416 4954 3120
rect 4990 2416 5024 3120
rect 5062 2416 5096 3120
rect 5132 2416 5166 3120
<< nsubdiffcont >>
rect 22776 972 22810 3962
<< locali >>
rect 5060 12504 5364 12506
rect 5060 12500 5370 12504
rect 5060 12352 5074 12500
rect 5160 12494 5370 12500
rect 5160 12352 5176 12494
rect 5354 12352 5370 12494
rect 5060 12346 5370 12352
rect 14654 11884 14788 11888
rect 14654 11720 14670 11884
rect 14722 11720 14732 11884
rect 14784 11720 14788 11884
rect 14654 11714 14788 11720
rect 17110 11884 17530 11888
rect 17110 11726 17122 11884
rect 17186 11882 17530 11884
rect 17186 11726 17336 11882
rect 17514 11726 17530 11882
rect 17110 11718 17530 11726
rect 5860 4810 5876 4878
rect 5938 4844 5944 4878
rect 5860 4794 6012 4810
rect 5864 4774 6012 4794
rect 5864 4652 5882 4774
rect 5988 4652 6012 4774
rect 5864 4636 6012 4652
rect 22776 3964 22850 3978
rect 22776 3962 22816 3964
rect 4730 3120 5208 3130
rect 4730 3056 4742 3120
rect 4740 2416 4742 3056
rect 4776 2416 4778 3120
rect 4812 2416 4814 3120
rect 4848 2416 4850 3120
rect 4884 2416 4886 3120
rect 4954 2416 4990 3120
rect 5058 2416 5062 3120
rect 5130 2416 5132 3120
rect 5166 2416 5168 3120
rect 5202 2416 5208 3120
rect 4740 2404 5208 2416
rect 4740 2402 5206 2404
rect 22810 974 22816 3962
rect 22850 974 22852 1004
rect 22810 972 22852 974
rect 22776 954 22852 972
<< viali >>
rect 5074 12352 5160 12500
rect 14732 11720 14784 11884
rect 17122 11726 17186 11884
rect 5904 4844 5910 4878
rect 5910 4844 5938 4878
rect 5978 4844 6012 4878
rect 5904 4810 5938 4844
rect 5978 4810 6012 4844
rect 4742 2416 4776 3120
rect 4814 2416 4848 3120
rect 4886 2416 4920 3120
rect 5024 2416 5058 3120
rect 5096 2416 5130 3120
rect 5168 2416 5202 3120
rect 22816 974 22850 3964
<< metal1 >>
rect 17126 15284 17194 15312
rect 18702 15284 18846 15632
rect 17126 15140 18846 15284
rect 6712 14650 6980 14740
rect 1492 14570 1592 14578
rect 1492 14492 1502 14570
rect 1580 14492 1592 14570
rect 6712 14566 9416 14650
rect 9774 14632 10412 14856
rect 6712 14538 6980 14566
rect 1492 14482 1592 14492
rect 1512 13890 1590 14482
rect 5630 14418 6184 14466
rect 5630 14336 5678 14418
rect 1512 13880 1606 13890
rect 1512 13802 1518 13880
rect 1596 13802 1606 13880
rect 1512 13792 1606 13802
rect 1512 13790 1602 13792
rect 1512 2168 1590 13790
rect 1794 13620 1846 13626
rect 1794 13562 1846 13568
rect 1796 13118 1844 13562
rect 1778 13112 1862 13118
rect 1778 13022 1862 13028
rect 2956 12870 3014 13254
rect 2952 12864 3034 12870
rect 2952 12748 2968 12864
rect 3026 12748 3034 12864
rect 2952 12736 3034 12748
rect 5628 12598 5676 13244
rect 5618 12588 5686 12598
rect 5618 12536 5626 12588
rect 5678 12536 5686 12588
rect 5618 12530 5686 12536
rect 5068 12510 5166 12512
rect 5066 12500 5168 12510
rect 5066 12352 5074 12500
rect 5160 12352 5168 12500
rect 4282 10772 4328 11468
rect 4416 11344 4460 11468
rect 4954 11412 4998 12322
rect 5066 12280 5168 12352
rect 6136 12324 6184 14418
rect 6798 14352 7404 14406
rect 7740 14354 7792 14566
rect 6792 12518 6854 13258
rect 6776 12512 6854 12518
rect 6776 12450 6784 12512
rect 6846 12450 6854 12512
rect 6776 12444 6854 12450
rect 7350 12416 7404 14352
rect 9332 13916 9416 14566
rect 10094 14068 10178 14632
rect 10094 14062 10188 14068
rect 10094 13978 10100 14062
rect 10184 13978 10188 14062
rect 10094 13972 10188 13978
rect 9324 13910 9420 13916
rect 9324 13826 9330 13910
rect 9414 13826 9420 13910
rect 9324 13820 9420 13826
rect 10434 13592 10522 13598
rect 10434 13498 10522 13504
rect 11578 13592 11666 13598
rect 11578 13498 11666 13504
rect 11936 13586 12082 14864
rect 12966 14834 13162 14864
rect 11936 13498 11942 13586
rect 12030 13498 12082 13586
rect 9550 13388 9638 13394
rect 9550 13294 9638 13300
rect 7584 12616 7634 13246
rect 8992 12748 9056 12756
rect 8992 12746 8998 12748
rect 8974 12696 8998 12746
rect 9050 12696 9056 12748
rect 8974 12688 9056 12696
rect 7576 12610 7642 12616
rect 7576 12558 7584 12610
rect 7636 12558 7642 12610
rect 7576 12544 7642 12558
rect 7342 12412 7410 12416
rect 7342 12360 7350 12412
rect 7404 12360 7410 12412
rect 7342 12354 7410 12360
rect 5056 12274 5168 12280
rect 5056 12260 5084 12274
rect 5034 12204 5084 12260
rect 5154 12204 5168 12274
rect 6126 12318 6194 12324
rect 6126 12266 6134 12318
rect 6186 12266 6194 12318
rect 6126 12260 6194 12266
rect 5034 12180 5168 12204
rect 5034 12174 5166 12180
rect 5034 11412 5078 12174
rect 8974 11988 9022 12688
rect 9562 11974 9624 13294
rect 10448 11978 10506 13498
rect 10686 13300 10692 13388
rect 10780 13300 10786 13388
rect 5278 11834 5348 11842
rect 5278 11756 5288 11834
rect 5340 11756 5348 11834
rect 5278 11750 5348 11756
rect 8564 11810 8638 11816
rect 8564 11758 8568 11810
rect 8634 11758 8638 11810
rect 8564 11754 8638 11758
rect 5158 11678 5208 11702
rect 5152 11672 5216 11678
rect 5152 11592 5160 11672
rect 5212 11592 5216 11672
rect 5152 11586 5216 11592
rect 5158 11428 5208 11586
rect 5158 11422 5216 11428
rect 5158 11370 5164 11422
rect 5158 11364 5216 11370
rect 4410 11338 4462 11344
rect 4410 11280 4462 11286
rect 4416 11160 4460 11280
rect 4404 11154 4460 11160
rect 4456 11102 4460 11154
rect 4404 11096 4460 11102
rect 4416 10976 4460 11096
rect 4406 10970 4460 10976
rect 4458 10918 4460 10970
rect 4406 10912 4460 10918
rect 4276 10766 4328 10772
rect 4276 10708 4328 10714
rect 4282 10580 4328 10708
rect 4268 10574 4328 10580
rect 4320 10522 4328 10574
rect 4268 10516 4328 10522
rect 4282 10388 4328 10516
rect 4276 10382 4328 10388
rect 4276 10324 4328 10330
rect 4282 7374 4328 10324
rect 4416 7374 4460 10912
rect 5158 11244 5208 11364
rect 5158 11238 5216 11244
rect 5158 11186 5164 11238
rect 5158 11180 5216 11186
rect 5158 11060 5208 11180
rect 5158 11054 5210 11060
rect 5158 10996 5210 11002
rect 4260 7368 4328 7374
rect 4260 7274 4268 7368
rect 4320 7274 4328 7368
rect 4260 7268 4328 7274
rect 4392 7368 4460 7374
rect 4392 7274 4396 7368
rect 4448 7274 4460 7368
rect 4392 7268 4460 7274
rect 3998 7120 4044 7134
rect 3990 7068 3996 7120
rect 4048 7068 4054 7120
rect 3900 7046 3946 7054
rect 3892 7040 3946 7046
rect 3944 6988 3946 7040
rect 3892 6982 3946 6988
rect 2030 6870 2174 6874
rect 2030 6738 2036 6870
rect 2168 6738 2174 6870
rect 2030 6734 2174 6738
rect 2032 5704 2164 6734
rect 3900 6278 3946 6982
rect 3998 6574 4044 7068
rect 4282 7050 4328 7268
rect 4416 7122 4460 7268
rect 4768 7126 4822 7134
rect 4412 7116 4464 7122
rect 4412 7058 4464 7064
rect 4764 7120 4822 7126
rect 4818 7066 4822 7120
rect 4764 7060 4822 7066
rect 4280 7044 4332 7050
rect 4280 6986 4332 6992
rect 4658 6752 4716 6758
rect 3998 6500 4144 6574
rect 3900 6264 3952 6278
rect 3896 6262 3952 6264
rect 3890 6258 3954 6262
rect 3890 6206 3896 6258
rect 3948 6206 3954 6258
rect 3890 6200 3954 6206
rect 3070 5908 3156 5914
rect 3070 5834 3078 5908
rect 3152 5834 3156 5908
rect 3070 5828 3156 5834
rect 2032 5698 2180 5704
rect 2032 5566 2044 5698
rect 2176 5566 2180 5698
rect 2032 5560 2180 5566
rect 3080 4666 3154 5828
rect 3998 5000 4044 6500
rect 4768 6466 4822 7060
rect 4744 6416 4822 6466
rect 4864 7046 4912 7054
rect 4864 7040 4916 7046
rect 4864 6982 4916 6988
rect 4864 6354 4912 6982
rect 4744 6308 4912 6354
rect 3998 4954 4488 5000
rect 4424 4888 4488 4954
rect 3072 4660 3158 4666
rect 3072 4586 3076 4660
rect 3150 4586 3158 4660
rect 3072 4580 3158 4586
rect 4576 4574 4642 4580
rect 4548 4558 4584 4574
rect 4500 4510 4584 4558
rect 4576 4502 4584 4510
rect 4636 4502 4642 4574
rect 4576 4496 4642 4502
rect 3674 3512 3732 3518
rect 3674 3448 3732 3454
rect 3676 3334 3728 3448
rect 4864 3376 4912 6308
rect 4954 6174 4998 10324
rect 5034 6696 5078 10324
rect 5158 6926 5208 10996
rect 5282 10842 5334 11750
rect 8436 11480 8514 11484
rect 8436 11414 8442 11480
rect 8508 11414 8514 11480
rect 8436 11410 8514 11414
rect 8320 11184 8398 11190
rect 8320 11118 8328 11184
rect 8394 11118 8398 11184
rect 8320 11112 8398 11118
rect 8192 10864 8270 10870
rect 5282 10836 5338 10842
rect 5282 10784 5286 10836
rect 8192 10798 8200 10864
rect 8266 10798 8270 10864
rect 8192 10794 8270 10798
rect 5282 10778 5338 10784
rect 8198 10792 8266 10794
rect 5282 10650 5334 10778
rect 8070 10754 8138 10756
rect 8068 10750 8140 10754
rect 8068 10684 8072 10750
rect 8138 10684 8140 10750
rect 8068 10676 8140 10684
rect 5282 10644 5340 10650
rect 5282 10592 5288 10644
rect 5282 10586 5340 10592
rect 5282 10458 5334 10586
rect 5282 10452 5338 10458
rect 5282 10400 5286 10452
rect 5282 10394 5338 10400
rect 7946 10436 8018 10442
rect 5158 6922 5210 6926
rect 5156 6920 5212 6922
rect 5156 6868 5158 6920
rect 5210 6868 5212 6920
rect 5156 6866 5212 6868
rect 5158 6862 5210 6866
rect 5026 6690 5090 6696
rect 5026 6638 5034 6690
rect 5086 6638 5090 6690
rect 5026 6632 5090 6638
rect 4946 6168 5002 6174
rect 4946 6116 4950 6168
rect 4946 6110 5002 6116
rect 4954 3516 4998 6110
rect 5034 5068 5078 6632
rect 5034 5062 5092 5068
rect 5034 4978 5038 5062
rect 5090 4978 5092 5062
rect 5034 4972 5092 4978
rect 5034 4580 5078 4972
rect 5030 4574 5082 4580
rect 5030 4496 5082 4502
rect 5034 3572 5078 4496
rect 5158 3848 5208 6862
rect 5282 6060 5334 10394
rect 7946 10370 7950 10436
rect 8016 10370 8018 10436
rect 7946 10364 8018 10370
rect 7816 10130 7898 10136
rect 7816 10064 7824 10130
rect 7890 10064 7898 10130
rect 7816 10056 7898 10064
rect 7710 9816 7782 9822
rect 7710 9750 7712 9816
rect 7778 9750 7782 9816
rect 7710 9744 7782 9750
rect 7594 8732 7660 8736
rect 7582 8722 7660 8732
rect 7582 8656 7588 8722
rect 7654 8656 7660 8722
rect 7582 8648 7660 8656
rect 7468 8410 7534 8414
rect 7458 8404 7536 8410
rect 7458 8338 7462 8404
rect 7528 8338 7536 8404
rect 7458 8332 7536 8338
rect 7344 8100 7410 8102
rect 7338 8094 7410 8100
rect 7404 8028 7410 8094
rect 7338 8022 7410 8028
rect 7214 7798 7292 7806
rect 7214 7732 7218 7798
rect 7284 7732 7292 7798
rect 7214 7726 7292 7732
rect 7080 6764 7166 6772
rect 7080 6698 7090 6764
rect 7156 6698 7166 6764
rect 7080 6692 7166 6698
rect 6948 6450 7030 6458
rect 6948 6384 6956 6450
rect 7022 6384 7030 6450
rect 6948 6378 7030 6384
rect 6826 6122 6904 6130
rect 5280 6054 5342 6060
rect 5280 6002 5286 6054
rect 5338 6002 5342 6054
rect 6826 6056 6832 6122
rect 6898 6056 6904 6122
rect 6826 6050 6904 6056
rect 5280 5996 5342 6002
rect 5150 3842 5210 3848
rect 5150 3776 5154 3842
rect 5206 3776 5210 3842
rect 5150 3768 5210 3776
rect 5034 3544 5082 3572
rect 4946 3510 5008 3516
rect 4946 3452 4948 3510
rect 5006 3452 5008 3510
rect 4946 3446 5008 3452
rect 5036 3418 5082 3544
rect 4706 3370 4912 3376
rect 4706 3250 4716 3370
rect 4836 3264 4912 3370
rect 5034 3412 5082 3418
rect 4836 3250 4864 3264
rect 4706 3242 4864 3250
rect 5034 3134 5078 3412
rect 4728 3120 5212 3134
rect 4728 2416 4742 3120
rect 4776 2416 4814 3120
rect 4848 2416 4886 3120
rect 4920 2416 5024 3120
rect 5058 2416 5096 3120
rect 5130 2416 5168 3120
rect 5202 2416 5212 3120
rect 4728 2398 5212 2416
rect 5282 2340 5334 5996
rect 6688 5834 6770 5840
rect 6688 5768 6696 5834
rect 6762 5768 6770 5834
rect 6688 5762 6770 5768
rect 5846 5038 6032 5062
rect 5846 4896 5888 5038
rect 6004 4896 6032 5038
rect 5846 4878 6032 4896
rect 5846 4810 5904 4878
rect 5938 4810 5978 4878
rect 6012 4810 6032 4878
rect 5846 4732 6032 4810
rect 5864 4636 6012 4732
rect 5264 2332 5334 2340
rect 5264 2264 5272 2332
rect 5324 2264 5334 2332
rect 5264 2258 5334 2264
rect 1478 2154 1590 2168
rect 1478 2076 1490 2154
rect 1568 2076 1590 2154
rect 1478 2064 1590 2076
rect 6700 1094 6766 5762
rect 6690 1092 6776 1094
rect 6684 1088 6782 1092
rect 6684 1002 6690 1088
rect 6776 1002 6782 1088
rect 6684 1000 6782 1002
rect 6690 996 6776 1000
rect 6830 936 6896 6050
rect 6812 930 6910 936
rect 6812 844 6820 930
rect 6906 844 6910 930
rect 6812 838 6910 844
rect 6960 794 7026 6378
rect 6954 788 7034 794
rect 6954 702 7034 708
rect 6912 622 7028 626
rect 6912 520 6920 622
rect 7022 604 7028 622
rect 7094 604 7160 6692
rect 7222 1520 7288 7726
rect 7222 628 7286 1520
rect 7344 750 7410 8022
rect 7468 872 7534 8332
rect 7594 1006 7660 8648
rect 7714 1138 7780 9744
rect 7830 1252 7896 10056
rect 7952 1386 8018 10364
rect 8070 1508 8136 10676
rect 8198 1642 8264 10792
rect 8322 1772 8388 11112
rect 8442 1898 8508 11410
rect 8568 2020 8634 11754
rect 8994 10780 9042 10802
rect 9582 10780 9644 10802
rect 10448 10772 10506 10804
rect 10740 10700 10778 13300
rect 11596 10692 11646 13498
rect 11936 13490 12082 13498
rect 11968 11412 12002 13490
rect 12968 13384 13162 14834
rect 15492 14630 16130 14854
rect 14046 13910 14340 13922
rect 14046 13826 14054 13910
rect 14324 13826 14340 13910
rect 14046 13816 14340 13826
rect 13572 13388 13660 13394
rect 12964 13380 13166 13384
rect 12964 13298 12970 13380
rect 13160 13298 13166 13380
rect 12964 13290 13166 13298
rect 13572 13294 13660 13300
rect 12412 12596 12480 12602
rect 12412 12544 12422 12596
rect 12474 12544 12480 12596
rect 12422 12538 12474 12544
rect 12046 11890 12098 11896
rect 12046 11832 12098 11838
rect 12052 11386 12090 11832
rect 12426 11382 12468 12538
rect 13140 12418 13192 12420
rect 13136 12414 13196 12418
rect 13136 12362 13140 12414
rect 13192 12362 13196 12414
rect 13136 12358 13196 12362
rect 13140 12356 13192 12358
rect 12506 12210 12574 12216
rect 12506 12158 12514 12210
rect 12566 12158 12574 12210
rect 12506 12152 12574 12158
rect 12520 11386 12558 12152
rect 12594 11792 12652 11798
rect 12594 11740 12598 11792
rect 12650 11740 12652 11792
rect 12594 11734 12652 11740
rect 12602 11382 12644 11734
rect 12802 11696 12870 11702
rect 12802 11644 12810 11696
rect 12862 11644 12870 11696
rect 12802 11638 12870 11644
rect 12818 11388 12854 11638
rect 13146 10310 13186 12356
rect 13592 11378 13638 13294
rect 13772 12598 13828 12604
rect 13772 12546 13774 12598
rect 13826 12546 13828 12598
rect 13772 12540 13828 12546
rect 13684 12416 13740 12422
rect 13684 12364 13686 12416
rect 13738 12364 13740 12416
rect 13684 12358 13740 12364
rect 13142 10284 13186 10310
rect 13132 10278 13198 10284
rect 13132 10224 13138 10278
rect 13192 10224 13198 10278
rect 13132 10218 13198 10224
rect 13638 10196 13640 10228
rect 13690 10050 13734 12358
rect 13688 10036 13734 10050
rect 13686 9916 13726 10036
rect 13776 9946 13822 12540
rect 14050 11340 14134 13816
rect 14256 11340 14340 13816
rect 14732 13380 14820 13386
rect 14732 13286 14820 13292
rect 14752 11890 14798 13286
rect 15636 12236 15892 14630
rect 16388 13592 16444 13616
rect 16388 13586 16454 13592
rect 16388 13498 16398 13586
rect 16388 13492 16454 13498
rect 15636 12220 15896 12236
rect 15634 12218 15896 12220
rect 15634 12166 15642 12218
rect 15886 12166 15896 12218
rect 15634 12160 15896 12166
rect 14990 12088 15050 12094
rect 14990 12036 14994 12088
rect 15046 12036 15050 12088
rect 14990 12030 15050 12036
rect 14726 11888 14798 11890
rect 14720 11884 14798 11888
rect 14720 11720 14732 11884
rect 14784 11720 14798 11884
rect 14720 11710 14798 11720
rect 14752 11378 14798 11710
rect 14996 11378 15042 12030
rect 16252 11980 16338 11988
rect 16252 11928 16260 11980
rect 16312 11928 16338 11980
rect 16252 11920 16338 11928
rect 16300 11386 16338 11920
rect 16388 11368 16444 13492
rect 16728 12598 16780 12604
rect 16728 12540 16780 12546
rect 16550 12424 16602 12430
rect 16550 12366 16602 12372
rect 16556 11622 16594 12366
rect 16732 11622 16776 12540
rect 17126 11896 17194 15140
rect 21206 14636 21844 14860
rect 18026 14448 18100 14450
rect 18016 14440 18116 14448
rect 18016 14366 18032 14440
rect 18106 14366 18116 14440
rect 18016 14358 18116 14366
rect 17256 12742 17320 12750
rect 17256 12688 17262 12742
rect 17314 12688 17320 12742
rect 17256 12676 17320 12688
rect 17116 11884 17194 11896
rect 17116 11880 17122 11884
rect 17114 11726 17122 11880
rect 17186 11726 17194 11884
rect 17116 11712 17194 11726
rect 16522 11582 16658 11622
rect 16522 11530 16550 11582
rect 16602 11530 16658 11582
rect 16522 11484 16658 11530
rect 16730 11584 16866 11622
rect 16730 11532 16754 11584
rect 16806 11532 16866 11584
rect 16730 11484 16866 11532
rect 17126 11356 17194 11712
rect 17260 11600 17314 12676
rect 17260 11594 17396 11600
rect 17260 11508 17304 11594
rect 17390 11508 17396 11594
rect 17260 11500 17396 11508
rect 17260 11370 17314 11500
rect 13688 9910 13734 9916
rect 8974 8698 9022 9572
rect 9562 8684 9624 9586
rect 10448 8688 10506 9582
rect 10740 8790 10778 9570
rect 11002 8810 11048 9578
rect 11596 8812 11646 9582
rect 13690 9270 13734 9910
rect 13690 9252 13760 9270
rect 13690 9208 13792 9252
rect 10736 8690 10778 8790
rect 10998 8728 11048 8810
rect 11592 8728 11646 8812
rect 11948 8842 12004 9064
rect 12054 8926 12092 9046
rect 12454 8958 12532 8962
rect 12452 8952 12532 8958
rect 12452 8940 12466 8952
rect 12422 8938 12466 8940
rect 12054 8888 12374 8926
rect 11948 8786 12292 8842
rect 12252 8740 12292 8786
rect 10736 8664 10774 8690
rect 10998 8642 11044 8728
rect 11592 8654 11642 8728
rect 12254 8680 12286 8740
rect 12336 8664 12374 8888
rect 12416 8896 12466 8938
rect 12522 8896 12532 8952
rect 12416 8890 12532 8896
rect 12416 8886 12530 8890
rect 12416 8884 12454 8886
rect 12416 8716 12450 8884
rect 13350 8872 13396 9054
rect 13594 8878 13640 9054
rect 13246 8858 13396 8872
rect 13240 8826 13396 8858
rect 13590 8866 13640 8878
rect 14256 8892 14340 9092
rect 13240 8736 13322 8826
rect 12416 8662 12448 8716
rect 13240 8638 13316 8736
rect 13590 8666 13638 8866
rect 14256 8856 14342 8892
rect 14256 8778 14344 8856
rect 14752 8814 14798 9054
rect 14262 8736 14344 8778
rect 14262 8634 14342 8736
rect 14750 8666 14798 8814
rect 14996 8876 15042 9054
rect 14996 8800 15148 8876
rect 16300 8850 16338 9046
rect 15072 8708 15148 8800
rect 15934 8834 15990 8840
rect 15934 8782 15936 8834
rect 15988 8782 15990 8834
rect 15934 8776 15990 8782
rect 16020 8812 16338 8850
rect 15940 8680 15972 8776
rect 16020 8746 16058 8812
rect 16388 8774 16444 9064
rect 18026 8976 18100 14358
rect 18184 13748 18276 13754
rect 18184 13674 18196 13748
rect 18270 13674 18276 13748
rect 18184 13668 18276 13674
rect 18020 8966 18110 8976
rect 18020 8892 18034 8966
rect 18108 8892 18110 8966
rect 18020 8884 18110 8892
rect 18026 8876 18100 8884
rect 18188 8858 18262 13668
rect 18338 12806 18428 12812
rect 18338 12732 18350 12806
rect 18424 12732 18428 12806
rect 18338 12726 18428 12732
rect 16110 8772 16444 8774
rect 16014 8724 16058 8746
rect 16014 8664 16052 8724
rect 16102 8718 16444 8772
rect 18182 8848 18270 8858
rect 18182 8774 18188 8848
rect 18262 8774 18270 8848
rect 18182 8766 18270 8774
rect 18188 8756 18262 8766
rect 16102 8680 16134 8718
rect 18342 8388 18416 12726
rect 19652 12622 19768 12628
rect 19652 12522 19660 12622
rect 19760 12522 19768 12622
rect 19652 12516 19768 12522
rect 19416 12502 19528 12510
rect 19200 12408 19312 12416
rect 19010 12310 19122 12332
rect 19010 12210 19016 12310
rect 19116 12210 19122 12310
rect 19010 12202 19122 12210
rect 19200 12308 19206 12408
rect 19306 12308 19312 12408
rect 19416 12402 19422 12502
rect 19522 12402 19528 12502
rect 19416 12392 19528 12402
rect 19200 12300 19312 12308
rect 18516 11792 18602 11798
rect 18516 11718 18526 11792
rect 18600 11718 18602 11792
rect 18516 11710 18602 11718
rect 18336 8386 18416 8388
rect 18334 8382 18418 8386
rect 18334 8308 18336 8382
rect 18410 8308 18418 8382
rect 18334 8302 18418 8308
rect 18342 8300 18416 8302
rect 8974 7374 9022 7546
rect 9562 7374 9624 7560
rect 8974 6792 9042 7374
rect 9562 6792 9644 7374
rect 10448 6792 10506 7556
rect 8994 6744 9042 6792
rect 9582 6738 9644 6792
rect 10740 6738 10778 7556
rect 11002 7348 11048 7564
rect 10984 7340 11050 7348
rect 10984 7258 10992 7340
rect 11044 7258 11050 7340
rect 10984 7252 11050 7258
rect 11002 6730 11048 7252
rect 11596 6772 11646 7568
rect 12260 6760 12292 7570
rect 12810 6842 12858 7586
rect 12806 6792 12884 6842
rect 12834 6742 12884 6792
rect 13246 6716 13322 7614
rect 13596 6838 13644 7586
rect 13596 6784 13690 6838
rect 13636 6738 13690 6784
rect 14052 6712 14132 7618
rect 14756 7084 14804 7586
rect 18518 7352 18592 11710
rect 18510 7340 18608 7352
rect 18510 7258 18522 7340
rect 18596 7258 18608 7340
rect 18510 7250 18608 7258
rect 18518 7244 18592 7250
rect 14756 7036 14872 7084
rect 14824 6768 14872 7036
rect 11866 6566 11930 6574
rect 11866 6514 11872 6566
rect 11924 6514 11930 6566
rect 15848 6562 15900 6568
rect 11866 6506 11930 6514
rect 15846 6510 15848 6556
rect 8974 3066 9022 5592
rect 9562 5376 9624 5606
rect 10448 5478 10506 5602
rect 10548 5540 10616 5546
rect 10548 5488 10556 5540
rect 10608 5488 10616 5540
rect 10548 5482 10616 5488
rect 10442 5472 10512 5478
rect 10442 5414 10448 5472
rect 10506 5414 10512 5472
rect 10442 5408 10512 5414
rect 9554 5374 9628 5376
rect 9554 5312 9560 5374
rect 9622 5312 9628 5374
rect 10448 5316 10506 5408
rect 10548 5360 10598 5482
rect 10740 5364 10778 5604
rect 11596 5470 11646 5616
rect 11882 5554 11924 6506
rect 15846 6504 15900 6510
rect 15744 6376 15796 6382
rect 15744 6318 15796 6324
rect 12134 6168 12212 6218
rect 11990 6010 12058 6016
rect 11990 5958 11998 6010
rect 12050 5958 12058 6010
rect 11990 5948 12058 5958
rect 11998 5944 12042 5948
rect 11876 5548 11932 5554
rect 11876 5496 11878 5548
rect 11930 5496 11932 5548
rect 11876 5490 11932 5496
rect 11998 5488 12038 5944
rect 12090 5580 12128 5652
rect 12082 5546 12138 5580
rect 12082 5494 12084 5546
rect 12136 5494 12138 5546
rect 11990 5482 12046 5488
rect 12082 5486 12138 5494
rect 11590 5466 11658 5470
rect 11590 5414 11598 5466
rect 11650 5414 11658 5466
rect 11990 5430 11992 5482
rect 12044 5430 12046 5482
rect 11990 5424 12046 5430
rect 11590 5412 11658 5414
rect 9554 5310 9628 5312
rect 9562 5068 9624 5310
rect 10334 5260 10506 5316
rect 10318 5258 10506 5260
rect 10538 5338 10598 5360
rect 10728 5358 10792 5364
rect 10318 5254 10410 5258
rect 10318 5170 10322 5254
rect 10406 5170 10410 5254
rect 10318 5164 10410 5170
rect 9552 5062 9636 5068
rect 10538 5036 10576 5338
rect 10728 5306 10734 5358
rect 10786 5306 10792 5358
rect 10728 5300 10792 5306
rect 11264 5258 11414 5296
rect 11314 5090 11414 5258
rect 12176 5242 12212 6168
rect 15650 6008 15702 6014
rect 15650 5950 15702 5956
rect 15550 5822 15602 5828
rect 15550 5764 15602 5770
rect 12440 5474 12492 5480
rect 12436 5470 12496 5474
rect 12436 5418 12440 5470
rect 12492 5418 12496 5470
rect 12436 5414 12496 5418
rect 12440 5412 12492 5414
rect 12176 5234 12272 5242
rect 12176 5182 12200 5234
rect 12192 5168 12200 5182
rect 12266 5168 12272 5234
rect 12442 5228 12486 5412
rect 12834 5386 12884 5632
rect 13636 5390 13690 5636
rect 14200 5550 14286 5556
rect 14200 5480 14208 5550
rect 14278 5480 14286 5550
rect 14200 5476 14286 5480
rect 12832 5334 12838 5386
rect 12890 5334 12896 5386
rect 13636 5382 13706 5390
rect 13636 5328 13646 5382
rect 13700 5328 13706 5382
rect 12192 5160 12272 5168
rect 12430 5222 12498 5228
rect 12430 5148 12498 5154
rect 12442 5132 12486 5148
rect 13232 5094 13420 5280
rect 14208 5190 14278 5476
rect 14572 5364 14616 5628
rect 14824 5484 14870 5628
rect 14824 5438 15466 5484
rect 14824 5436 14870 5438
rect 14208 5126 14216 5190
rect 14268 5126 14278 5190
rect 14208 5118 14278 5126
rect 14514 5316 14616 5364
rect 9552 4972 9636 4978
rect 10450 5024 10576 5036
rect 11216 5026 11264 5090
rect 11464 5026 11512 5090
rect 13178 5030 13226 5094
rect 13426 5030 13474 5094
rect 14514 5066 14560 5316
rect 15420 5244 15466 5438
rect 15410 5238 15472 5244
rect 15410 5170 15414 5238
rect 15466 5170 15472 5238
rect 15410 5164 15472 5170
rect 14492 5060 14584 5066
rect 10450 4960 10458 5024
rect 10522 4972 10576 5024
rect 14492 4984 14500 5060
rect 14576 4984 14584 5060
rect 14492 4978 14584 4984
rect 10522 4960 10538 4972
rect 10450 4952 10538 4960
rect 11216 4758 11264 4822
rect 11464 4756 11512 4820
rect 13178 4762 13226 4826
rect 13426 4760 13474 4824
rect 15420 4530 15466 5164
rect 15394 4486 15466 4530
rect 15354 4440 15466 4486
rect 15354 4438 15462 4440
rect 10492 3916 10556 4266
rect 11216 4204 11264 4268
rect 11464 4202 11512 4266
rect 11264 4072 11316 4164
rect 11412 4076 11464 4164
rect 11262 4066 11318 4072
rect 11262 4004 11318 4010
rect 11410 4070 11466 4076
rect 11410 4008 11466 4014
rect 10468 3896 10576 3916
rect 10468 3804 10478 3896
rect 10570 3804 10576 3896
rect 10468 3796 10576 3804
rect 11264 3722 11316 4004
rect 11412 3722 11464 4008
rect 8894 3032 9024 3066
rect 11264 3036 11464 3722
rect 12166 3712 12234 4270
rect 12154 3706 12246 3712
rect 12154 3608 12246 3614
rect 12452 3534 12520 4268
rect 13178 4208 13226 4272
rect 13426 4208 13474 4272
rect 13226 4072 13278 4170
rect 13224 4066 13280 4072
rect 13224 4004 13280 4010
rect 13226 3768 13278 4004
rect 13374 3768 13426 4170
rect 12434 3528 12538 3534
rect 12434 3436 12440 3528
rect 12532 3436 12538 3528
rect 12434 3430 12538 3436
rect 13226 3048 13426 3768
rect 14136 3358 14190 4276
rect 15550 4196 15600 5764
rect 15650 4376 15700 5950
rect 15746 4558 15796 6318
rect 15846 4736 15896 6504
rect 19014 5036 19114 12202
rect 19200 6092 19300 12300
rect 19426 7138 19526 12392
rect 19652 8172 19752 12516
rect 21424 12196 21680 14636
rect 21422 12190 21680 12196
rect 21678 11934 21680 12190
rect 21422 11928 21680 11934
rect 21424 11830 21680 11928
rect 22296 11594 22336 11600
rect 22278 11588 22340 11594
rect 22278 11502 22286 11588
rect 22338 11502 22340 11588
rect 22278 11494 22340 11502
rect 21514 11330 21584 11336
rect 21514 11246 21520 11330
rect 21572 11246 21584 11330
rect 21514 11240 21584 11246
rect 20716 10686 20810 10698
rect 20716 10606 20720 10686
rect 20800 10606 20810 10686
rect 20716 10600 20810 10606
rect 19642 8166 19752 8172
rect 19742 8066 19752 8166
rect 19642 8060 19752 8066
rect 19424 7122 19528 7138
rect 19424 7028 19426 7122
rect 19526 7028 19528 7122
rect 19424 7026 19528 7028
rect 19198 6090 19302 6092
rect 19198 5990 19200 6090
rect 19300 5990 19302 6090
rect 19198 5988 19302 5990
rect 18982 5030 19114 5036
rect 18982 4930 18990 5030
rect 19090 4930 19114 5030
rect 18982 4922 19114 4930
rect 15836 4728 15910 4736
rect 15836 4628 15844 4728
rect 15896 4628 15910 4728
rect 15836 4620 15910 4628
rect 15730 4548 15804 4558
rect 15730 4448 15736 4548
rect 15788 4448 15804 4548
rect 15730 4442 15804 4448
rect 15632 4368 15706 4376
rect 15632 4268 15642 4368
rect 15694 4268 15706 4368
rect 15632 4260 15706 4268
rect 15538 4188 15608 4196
rect 14114 3346 14212 3358
rect 14114 3254 14118 3346
rect 14210 3254 14212 3346
rect 14114 3246 14212 3254
rect 13226 3040 13630 3048
rect 8894 2808 8904 3032
rect 8956 2808 9024 3032
rect 11168 3028 11554 3036
rect 8894 2802 9024 2808
rect 11060 3024 11554 3028
rect 11060 3020 11326 3024
rect 11060 2796 11178 3020
rect 11550 2800 11554 3024
rect 11402 2796 11554 2800
rect 11060 2790 11554 2796
rect 13130 3028 13630 3040
rect 13130 2790 13140 3028
rect 13512 2790 13630 3028
rect 8564 2016 8638 2020
rect 8564 1950 8568 2016
rect 8634 1950 8638 2016
rect 8564 1944 8638 1950
rect 8434 1892 8512 1898
rect 8434 1826 8444 1892
rect 8510 1826 8512 1892
rect 8434 1820 8512 1826
rect 8314 1766 8390 1772
rect 8314 1700 8318 1766
rect 8384 1700 8390 1766
rect 8314 1694 8390 1700
rect 8196 1640 8266 1642
rect 8196 1574 8198 1640
rect 8264 1574 8266 1640
rect 8196 1568 8266 1574
rect 8068 1504 8140 1508
rect 8068 1438 8070 1504
rect 8136 1438 8140 1504
rect 8068 1432 8140 1438
rect 7950 1384 8018 1386
rect 7946 1380 8022 1384
rect 7946 1314 7950 1380
rect 8016 1314 8022 1380
rect 7946 1310 8022 1314
rect 7950 1308 8016 1310
rect 7830 1180 7896 1186
rect 7714 1066 7780 1072
rect 7594 1000 7664 1006
rect 7594 940 7598 1000
rect 7598 928 7664 934
rect 7468 800 7534 806
rect 7340 744 7410 750
rect 7406 684 7410 744
rect 7340 670 7406 676
rect 7022 538 7160 604
rect 7218 622 7306 628
rect 7218 548 7224 622
rect 7298 548 7306 622
rect 7218 544 7306 548
rect 7022 520 7028 538
rect 6912 516 7028 520
rect 11060 492 11248 2790
rect 13130 2784 13630 2790
rect 13452 784 13630 2784
rect 15284 2154 15350 4152
rect 15538 4088 15546 4188
rect 15598 4088 15608 4188
rect 15538 4082 15608 4088
rect 19014 3358 19114 4922
rect 19200 3540 19300 5988
rect 19426 3714 19526 7026
rect 19652 3918 19752 8060
rect 20230 5534 20346 5542
rect 20230 5434 20238 5534
rect 20338 5434 20346 5534
rect 20230 5430 20346 5434
rect 20236 5428 20338 5430
rect 19652 3912 19764 3918
rect 19652 3812 19664 3912
rect 19652 3806 19764 3812
rect 19652 3780 19752 3806
rect 19426 3616 19526 3622
rect 19200 3442 19300 3448
rect 19014 3260 19114 3266
rect 20236 3054 20336 5428
rect 20110 3032 20336 3054
rect 20110 2808 20122 3032
rect 20310 2808 20336 3032
rect 20110 2798 20336 2808
rect 15272 2148 15358 2154
rect 15272 2082 15280 2148
rect 15346 2082 15358 2148
rect 15272 2076 15358 2082
rect 20726 1930 20806 10600
rect 20910 10478 20916 10550
rect 20988 10478 20994 10550
rect 20724 1924 20818 1930
rect 20724 1844 20732 1924
rect 20812 1844 20818 1924
rect 20724 1838 20818 1844
rect 20912 1770 20990 10478
rect 21094 10082 21184 10086
rect 21094 10004 21100 10082
rect 21178 10004 21184 10082
rect 21094 10000 21184 10004
rect 20906 1762 20998 1770
rect 20906 1684 20914 1762
rect 20992 1684 20998 1762
rect 20906 1676 20998 1684
rect 21098 1606 21176 10000
rect 21266 9948 21342 9950
rect 21262 9944 21346 9948
rect 21262 9892 21266 9944
rect 21342 9892 21346 9944
rect 21262 9888 21346 9892
rect 21094 1598 21188 1606
rect 21094 1520 21100 1598
rect 21178 1520 21188 1598
rect 21094 1514 21188 1520
rect 21266 1446 21342 9888
rect 21534 5242 21580 11240
rect 22296 10844 22336 11494
rect 22998 10846 23036 14900
rect 23666 13142 23830 13148
rect 23666 13130 23676 13142
rect 23654 13000 23676 13130
rect 23818 13000 23830 13142
rect 23654 12992 23830 13000
rect 23654 9192 23796 12992
rect 23628 9184 23796 9192
rect 23628 9042 23638 9184
rect 23780 9042 23796 9184
rect 23628 9034 23796 9042
rect 22772 5534 22916 5540
rect 22772 5432 22798 5534
rect 22900 5432 22916 5534
rect 22772 5426 22916 5432
rect 21534 5196 21582 5242
rect 21534 4034 21580 5196
rect 22784 4024 22886 5426
rect 22756 4014 22886 4024
rect 22754 3978 22886 4014
rect 22748 3976 22886 3978
rect 22748 3964 22868 3976
rect 22748 3528 22816 3964
rect 22678 3330 22816 3528
rect 22748 3174 22816 3330
rect 22758 3054 22816 3174
rect 22750 3052 22816 3054
rect 22748 2852 22816 3052
rect 22758 2732 22816 2852
rect 22748 2530 22816 2732
rect 22756 2410 22816 2530
rect 22748 2206 22816 2410
rect 22758 2086 22816 2206
rect 22748 1884 22816 2086
rect 22756 1764 22816 1884
rect 21260 1438 21348 1446
rect 21260 1362 21264 1438
rect 21340 1362 21348 1438
rect 22748 1390 22816 1764
rect 21260 1354 21348 1362
rect 22756 974 22816 1390
rect 22850 3902 22868 3964
rect 22850 974 22864 3902
rect 22756 948 22864 974
rect 13452 638 13636 784
rect 13446 492 13630 638
<< via1 >>
rect 1502 14492 1580 14570
rect 1518 13802 1596 13880
rect 1794 13568 1846 13620
rect 1778 13028 1862 13112
rect 2968 12748 3026 12864
rect 5626 12536 5678 12588
rect 6784 12450 6846 12512
rect 10100 13978 10184 14062
rect 9330 13826 9414 13910
rect 10434 13504 10522 13592
rect 11578 13504 11666 13592
rect 11942 13498 12030 13586
rect 9550 13300 9638 13388
rect 8998 12696 9050 12748
rect 7584 12558 7636 12610
rect 7350 12360 7404 12412
rect 5084 12204 5154 12274
rect 6134 12266 6186 12318
rect 10692 13300 10780 13388
rect 5288 11756 5340 11834
rect 8568 11758 8634 11810
rect 5160 11592 5212 11672
rect 5164 11370 5216 11422
rect 4410 11286 4462 11338
rect 4404 11102 4456 11154
rect 4406 10918 4458 10970
rect 4276 10714 4328 10766
rect 4268 10522 4320 10574
rect 4276 10330 4328 10382
rect 5164 11186 5216 11238
rect 5158 11002 5210 11054
rect 4268 7274 4320 7368
rect 4396 7274 4448 7368
rect 3996 7068 4048 7120
rect 3892 6988 3944 7040
rect 2036 6738 2168 6870
rect 4412 7064 4464 7116
rect 4764 7066 4818 7120
rect 4280 6992 4332 7044
rect 3896 6206 3948 6258
rect 3078 5834 3152 5908
rect 2044 5566 2176 5698
rect 4864 6988 4916 7040
rect 3076 4586 3150 4660
rect 4584 4502 4636 4574
rect 3674 3454 3732 3512
rect 8442 11414 8508 11480
rect 8328 11118 8394 11184
rect 5286 10784 5338 10836
rect 8200 10798 8266 10864
rect 8072 10684 8138 10750
rect 5288 10592 5340 10644
rect 5286 10400 5338 10452
rect 5158 6868 5210 6920
rect 5034 6638 5086 6690
rect 4950 6116 5002 6168
rect 5038 4978 5090 5062
rect 5030 4502 5082 4574
rect 7950 10370 8016 10436
rect 7824 10064 7890 10130
rect 7712 9750 7778 9816
rect 7588 8656 7654 8722
rect 7462 8338 7528 8404
rect 7338 8028 7404 8094
rect 7218 7732 7284 7798
rect 7090 6698 7156 6764
rect 6956 6384 7022 6450
rect 5286 6002 5338 6054
rect 6832 6056 6898 6122
rect 5154 3776 5206 3842
rect 4948 3452 5006 3510
rect 4716 3250 4836 3370
rect 6696 5768 6762 5834
rect 5888 4896 6004 5038
rect 5272 2264 5324 2332
rect 1490 2076 1568 2154
rect 6690 1002 6776 1088
rect 6820 844 6906 930
rect 6954 708 7034 788
rect 6920 520 7022 622
rect 14054 13826 14324 13910
rect 12970 13298 13160 13380
rect 13572 13300 13660 13388
rect 12422 12544 12474 12596
rect 12046 11838 12098 11890
rect 13140 12362 13192 12414
rect 12514 12158 12566 12210
rect 12598 11740 12650 11792
rect 12810 11644 12862 11696
rect 13774 12546 13826 12598
rect 13686 12364 13738 12416
rect 13138 10224 13192 10278
rect 14732 13292 14820 13380
rect 16398 13498 16454 13586
rect 15642 12166 15886 12218
rect 14994 12036 15046 12088
rect 16260 11928 16312 11980
rect 16728 12546 16780 12598
rect 16550 12372 16602 12424
rect 18032 14366 18106 14440
rect 17262 12688 17314 12742
rect 16550 11530 16602 11582
rect 16754 11532 16806 11584
rect 17304 11508 17390 11594
rect 12466 8896 12522 8952
rect 15936 8782 15988 8834
rect 18196 13674 18270 13748
rect 18034 8892 18108 8966
rect 18350 12732 18424 12806
rect 18188 8774 18262 8848
rect 19660 12522 19760 12622
rect 19016 12210 19116 12310
rect 19206 12308 19306 12408
rect 19422 12402 19522 12502
rect 18526 11718 18600 11792
rect 18336 8308 18410 8382
rect 10992 7258 11044 7340
rect 18522 7258 18596 7340
rect 11872 6514 11924 6566
rect 15848 6510 15900 6562
rect 10556 5488 10608 5540
rect 10448 5414 10506 5472
rect 9560 5312 9622 5374
rect 15744 6324 15796 6376
rect 11998 5958 12050 6010
rect 11878 5496 11930 5548
rect 12084 5494 12136 5546
rect 11598 5414 11650 5466
rect 11992 5430 12044 5482
rect 10322 5170 10406 5254
rect 9552 4978 9636 5062
rect 10734 5306 10786 5358
rect 15650 5956 15702 6008
rect 15550 5770 15602 5822
rect 12440 5418 12492 5470
rect 12200 5168 12266 5234
rect 14208 5480 14278 5550
rect 12838 5334 12890 5386
rect 13646 5328 13700 5382
rect 12430 5154 12498 5222
rect 14216 5126 14268 5190
rect 15414 5170 15466 5238
rect 10458 4960 10522 5024
rect 14500 4984 14576 5060
rect 11262 4010 11318 4066
rect 11410 4014 11466 4070
rect 10478 3804 10570 3896
rect 12154 3614 12246 3706
rect 13224 4010 13280 4066
rect 12440 3436 12532 3528
rect 21422 11934 21678 12190
rect 22286 11502 22338 11588
rect 21520 11246 21572 11330
rect 20720 10606 20800 10686
rect 19642 8066 19742 8166
rect 19426 7028 19526 7122
rect 19200 5990 19300 6090
rect 18990 4930 19090 5030
rect 15844 4628 15896 4728
rect 15736 4448 15788 4548
rect 15642 4268 15694 4368
rect 14118 3254 14210 3346
rect 8904 2808 8956 3032
rect 11326 3020 11550 3024
rect 11178 2800 11550 3020
rect 11178 2796 11402 2800
rect 13140 2790 13512 3028
rect 8568 1950 8634 2016
rect 8444 1826 8510 1892
rect 8318 1700 8384 1766
rect 8198 1574 8264 1640
rect 8070 1438 8136 1504
rect 7950 1314 8016 1380
rect 7830 1186 7896 1252
rect 7714 1072 7780 1138
rect 7598 934 7664 1000
rect 7468 806 7534 872
rect 7340 676 7406 744
rect 7224 548 7298 622
rect 15546 4088 15598 4188
rect 20238 5434 20338 5534
rect 19664 3812 19764 3912
rect 19426 3622 19526 3714
rect 19200 3448 19300 3540
rect 19014 3266 19114 3358
rect 20122 2808 20310 3032
rect 15280 2082 15346 2148
rect 20916 10478 20988 10550
rect 20732 1844 20812 1924
rect 21100 10004 21178 10082
rect 20914 1684 20992 1762
rect 21266 9892 21342 9944
rect 21100 1520 21178 1598
rect 23676 13000 23818 13142
rect 23638 9042 23780 9184
rect 22798 5432 22900 5534
rect 21264 1362 21340 1438
<< metal2 >>
rect 1250 14554 1386 14798
rect 1496 14570 1586 14574
rect 1496 14554 1502 14570
rect 1250 14508 1502 14554
rect 1250 14334 1386 14508
rect 1496 14492 1502 14508
rect 1580 14492 1586 14570
rect 1496 14488 1586 14492
rect 18020 14440 18112 14444
rect 24194 14440 24366 14710
rect 18020 14366 18032 14440
rect 18106 14366 24366 14440
rect 18020 14362 18112 14366
rect 24194 14290 24366 14366
rect 1220 14114 1716 14116
rect 1220 14036 2010 14114
rect 1674 13962 2010 14036
rect 5206 14096 5356 14098
rect 5206 14036 5530 14096
rect 10096 14062 10186 14066
rect 10094 14050 10100 14062
rect 5206 14002 5254 14036
rect 5470 13992 5530 14036
rect 5616 13990 10100 14050
rect 10094 13978 10100 13990
rect 10184 13978 10190 14062
rect 10096 13974 10186 13978
rect 9326 13910 9416 13914
rect 14048 13910 14332 13916
rect 1250 13716 1386 13892
rect 1516 13880 1602 13888
rect 1516 13802 1518 13880
rect 1596 13802 1602 13880
rect 9324 13826 9330 13910
rect 9414 13908 9420 13910
rect 14048 13908 14054 13910
rect 9414 13828 14054 13908
rect 9414 13826 9420 13828
rect 14048 13826 14054 13828
rect 14324 13908 14332 13910
rect 14324 13828 14342 13908
rect 14324 13826 14332 13828
rect 9326 13822 9416 13826
rect 14048 13820 14332 13826
rect 1516 13794 1602 13802
rect 1516 13792 1904 13794
rect 1534 13748 1904 13792
rect 18186 13748 18274 13752
rect 24194 13748 24366 13884
rect 1250 13652 1922 13716
rect 18186 13674 18196 13748
rect 18270 13674 24366 13748
rect 18186 13670 18274 13674
rect 1250 13428 1386 13652
rect 1788 13568 1794 13620
rect 1846 13574 1904 13620
rect 1846 13568 1852 13574
rect 10428 13504 10434 13592
rect 10522 13586 10528 13592
rect 11572 13586 11578 13592
rect 10522 13504 11578 13586
rect 11666 13586 11672 13592
rect 11666 13504 11942 13586
rect 10458 13498 11942 13504
rect 12030 13498 16398 13586
rect 16454 13498 16460 13586
rect 24194 13464 24366 13674
rect 10692 13388 10780 13394
rect 1650 13354 1956 13386
rect 1288 13288 1956 13354
rect 9544 13300 9550 13388
rect 9638 13384 9644 13388
rect 9638 13300 10692 13384
rect 13566 13384 13572 13388
rect 10780 13380 13572 13384
rect 10780 13300 12970 13380
rect 9574 13298 12970 13300
rect 13160 13300 13572 13380
rect 13660 13384 13666 13388
rect 13660 13380 14846 13384
rect 13660 13300 14732 13380
rect 13160 13298 14732 13300
rect 9574 13296 14732 13298
rect 10692 13294 10780 13296
rect 14726 13292 14732 13296
rect 14820 13296 14846 13380
rect 14820 13292 14826 13296
rect 1288 13274 1742 13288
rect 1288 13234 1368 13274
rect 1218 13154 1368 13234
rect 23670 13112 23676 13142
rect 1772 13028 1778 13112
rect 1862 13028 23676 13112
rect 23670 13000 23676 13028
rect 23818 13000 23824 13142
rect 1160 12864 1296 12998
rect 2944 12864 3038 12868
rect 1160 12748 2968 12864
rect 3026 12748 3038 12864
rect 18342 12806 18426 12810
rect 24188 12806 24360 13066
rect 1160 12700 1304 12748
rect 2944 12744 3038 12748
rect 8994 12748 9054 12754
rect 1160 12534 1296 12700
rect 8994 12696 8998 12748
rect 9050 12742 9054 12748
rect 17258 12742 17318 12748
rect 9050 12696 17262 12742
rect 8994 12690 9054 12696
rect 17258 12688 17262 12696
rect 17314 12696 17332 12742
rect 18342 12732 18350 12806
rect 18424 12732 24360 12806
rect 18342 12728 18426 12732
rect 17314 12688 17318 12696
rect 17258 12680 17318 12688
rect 24188 12646 24360 12732
rect 7578 12610 7640 12614
rect 5620 12594 5684 12596
rect 7578 12594 7584 12610
rect 5620 12588 7584 12594
rect 5620 12536 5626 12588
rect 5678 12558 7584 12588
rect 7636 12594 7642 12610
rect 12414 12596 12478 12600
rect 13768 12598 13832 12600
rect 12414 12594 12422 12596
rect 7636 12558 12422 12594
rect 5678 12548 12422 12558
rect 5678 12536 5684 12548
rect 7578 12546 7640 12548
rect 12414 12544 12422 12548
rect 12474 12594 12480 12596
rect 13768 12594 13774 12598
rect 12474 12548 13774 12594
rect 12474 12544 12480 12548
rect 13768 12546 13774 12548
rect 13826 12594 13832 12598
rect 16722 12594 16728 12598
rect 13826 12548 16728 12594
rect 13826 12546 13832 12548
rect 16722 12546 16728 12548
rect 16780 12594 16786 12598
rect 19654 12594 19660 12622
rect 16780 12548 19660 12594
rect 16780 12546 16786 12548
rect 13768 12544 13832 12546
rect 5620 12532 5684 12536
rect 19654 12522 19660 12548
rect 19760 12522 19766 12622
rect 19654 12520 19766 12522
rect 6778 12512 6852 12516
rect 1160 12434 1262 12458
rect 6778 12450 6784 12512
rect 6846 12504 6852 12512
rect 19418 12504 19526 12508
rect 6846 12502 19526 12504
rect 6846 12458 19422 12502
rect 6846 12450 6852 12458
rect 6778 12446 6852 12450
rect 1160 12376 1780 12434
rect 13680 12416 13744 12418
rect 13138 12414 13194 12416
rect 1262 12374 1780 12376
rect 7344 12412 7406 12414
rect 13134 12412 13140 12414
rect 7344 12360 7350 12412
rect 7404 12366 13140 12412
rect 7404 12360 7410 12366
rect 13134 12362 13140 12366
rect 13192 12412 13198 12414
rect 13680 12412 13686 12416
rect 13192 12366 13686 12412
rect 13192 12362 13198 12366
rect 13680 12364 13686 12366
rect 13738 12412 13744 12416
rect 16544 12412 16550 12424
rect 13738 12372 16550 12412
rect 16602 12412 16608 12424
rect 19202 12412 19310 12414
rect 16602 12408 19310 12412
rect 16602 12372 19206 12408
rect 13738 12366 19206 12372
rect 13738 12364 13744 12366
rect 13680 12362 13744 12364
rect 13138 12360 13194 12362
rect 7344 12356 7406 12360
rect 6128 12320 6192 12322
rect 19014 12320 19120 12326
rect 6128 12318 19120 12320
rect 1152 12274 1254 12278
rect 5080 12274 5160 12276
rect 1152 12204 5084 12274
rect 5154 12204 5160 12274
rect 6128 12266 6134 12318
rect 6186 12310 19120 12318
rect 6186 12274 19016 12310
rect 6186 12266 6192 12274
rect 6128 12262 6192 12266
rect 15638 12218 15894 12224
rect 1152 12196 1254 12204
rect 5080 12198 5160 12204
rect 12508 12210 12572 12212
rect 12508 12158 12514 12210
rect 12566 12204 12572 12210
rect 15638 12204 15642 12218
rect 12566 12166 15642 12204
rect 15886 12166 15894 12218
rect 19014 12210 19016 12274
rect 19116 12210 19120 12310
rect 19202 12308 19206 12366
rect 19306 12308 19310 12408
rect 19418 12402 19422 12458
rect 19522 12402 19526 12502
rect 19418 12396 19526 12402
rect 19202 12302 19310 12308
rect 19014 12204 19120 12210
rect 12566 12162 15894 12166
rect 12566 12158 12572 12162
rect 12508 12156 12572 12158
rect 1096 11834 1350 12126
rect 10520 12074 11090 12114
rect 14992 12088 15048 12092
rect 11050 11974 11090 12074
rect 14988 12036 14994 12088
rect 15046 12082 15052 12088
rect 21416 12082 21422 12190
rect 15046 12040 21422 12082
rect 15046 12036 15052 12040
rect 14992 12032 15048 12036
rect 16254 11980 16316 11986
rect 16254 11974 16260 11980
rect 8756 11904 8868 11938
rect 11050 11934 16260 11974
rect 16254 11928 16260 11934
rect 16312 11928 16316 11980
rect 21416 11934 21422 12040
rect 21678 11934 21684 12190
rect 16254 11922 16316 11928
rect 3366 11834 3426 11836
rect 5284 11834 5342 11838
rect 1096 11756 5288 11834
rect 5340 11756 5348 11834
rect 8562 11758 8568 11810
rect 8634 11792 8640 11810
rect 8756 11792 8790 11904
rect 12040 11880 12046 11890
rect 11040 11840 12046 11880
rect 8634 11758 8792 11792
rect 11040 11764 11080 11840
rect 12040 11838 12046 11840
rect 12098 11880 12104 11890
rect 12098 11840 12114 11880
rect 12098 11838 12104 11840
rect 12592 11792 12654 11794
rect 18518 11792 18604 11796
rect 24188 11792 24360 12188
rect 12592 11786 12598 11792
rect 1096 11750 1350 11756
rect 5284 11752 5342 11756
rect 10520 11724 11080 11764
rect 11142 11746 12598 11786
rect 5156 11672 5214 11676
rect 2666 11592 5160 11672
rect 5212 11592 5218 11672
rect 1154 11054 1408 11228
rect 2666 11054 2746 11592
rect 5156 11590 5214 11592
rect 8756 11538 8868 11572
rect 8442 11484 8508 11486
rect 8438 11480 8512 11484
rect 3426 11456 3500 11458
rect 3068 11410 3500 11456
rect 5158 11412 5164 11422
rect 3068 11384 4552 11410
rect 3068 11244 3192 11384
rect 3426 11376 4552 11384
rect 5044 11378 5164 11412
rect 5158 11370 5164 11378
rect 5216 11412 5222 11422
rect 8438 11414 8442 11480
rect 8508 11464 8512 11480
rect 8756 11464 8790 11538
rect 8508 11430 8790 11464
rect 8508 11414 8512 11430
rect 8756 11428 8790 11430
rect 11142 11414 11182 11746
rect 12592 11740 12598 11746
rect 12650 11740 12656 11792
rect 12592 11738 12654 11740
rect 18518 11718 18526 11792
rect 18600 11768 24360 11792
rect 18600 11718 24338 11768
rect 18518 11712 18600 11718
rect 12804 11696 12868 11698
rect 12804 11690 12810 11696
rect 5216 11378 5234 11412
rect 8438 11408 8512 11414
rect 5216 11370 5222 11378
rect 10520 11374 11182 11414
rect 11252 11650 12810 11690
rect 4404 11286 4410 11338
rect 4462 11328 4468 11338
rect 4462 11294 4552 11328
rect 4462 11286 4468 11294
rect 3426 11244 3500 11252
rect 1154 10974 2746 11054
rect 2962 11226 3500 11244
rect 5158 11228 5164 11238
rect 2962 11192 4552 11226
rect 5044 11194 5164 11228
rect 2962 11170 3500 11192
rect 5158 11186 5164 11194
rect 5216 11228 5222 11238
rect 5216 11194 5234 11228
rect 5216 11186 5222 11194
rect 8748 11192 8868 11226
rect 8322 11184 8400 11188
rect 2962 11148 3192 11170
rect 2962 11058 3184 11148
rect 4398 11102 4404 11154
rect 4456 11144 4462 11154
rect 4456 11110 4552 11144
rect 8322 11118 8328 11184
rect 8394 11168 8400 11184
rect 8748 11168 8782 11192
rect 8394 11134 8782 11168
rect 8394 11118 8400 11134
rect 8322 11114 8400 11118
rect 4456 11102 4462 11110
rect 3426 11058 3500 11066
rect 11252 11064 11292 11650
rect 12804 11644 12810 11650
rect 12862 11690 12868 11696
rect 12862 11650 12884 11690
rect 12862 11644 12868 11650
rect 12804 11642 12868 11644
rect 16532 11588 16648 11618
rect 16532 11582 16556 11588
rect 16532 11530 16550 11582
rect 16620 11530 16648 11588
rect 16736 11586 16852 11616
rect 16736 11584 16762 11586
rect 16736 11532 16754 11584
rect 16532 11524 16556 11530
rect 16620 11524 16660 11530
rect 16532 11492 16660 11524
rect 16612 11370 16660 11492
rect 16736 11522 16762 11532
rect 16826 11522 16852 11586
rect 16736 11490 16852 11522
rect 17300 11594 17394 11600
rect 17300 11508 17304 11594
rect 17390 11588 17394 11594
rect 22280 11590 22338 11592
rect 22280 11588 22340 11590
rect 24386 11588 24476 11592
rect 17390 11508 22286 11588
rect 17300 11502 22286 11508
rect 22338 11502 24478 11588
rect 22280 11500 22340 11502
rect 22280 11496 22338 11500
rect 24286 11366 24358 11368
rect 21516 11330 21576 11334
rect 24174 11330 24358 11366
rect 2962 11042 3500 11058
rect 5152 11044 5158 11054
rect 2962 11008 4552 11042
rect 5044 11010 5158 11044
rect 2962 10984 3500 11008
rect 5152 11002 5158 11010
rect 5210 11044 5216 11054
rect 5210 11010 5234 11044
rect 10512 11024 11292 11064
rect 11882 11290 11940 11326
rect 5210 11002 5216 11010
rect 2962 10976 3142 10984
rect 1154 10852 1408 10974
rect 1240 10066 1494 10242
rect 2962 10066 3036 10976
rect 4400 10918 4406 10970
rect 4458 10960 4464 10970
rect 4458 10926 4552 10960
rect 4458 10918 4464 10926
rect 8194 10864 8272 10866
rect 3258 10838 4556 10842
rect 1240 9992 3036 10066
rect 3200 10804 4556 10838
rect 5280 10830 5286 10836
rect 3200 10768 3500 10804
rect 5038 10790 5286 10830
rect 5280 10784 5286 10790
rect 5338 10830 5344 10836
rect 5338 10790 5364 10830
rect 8194 10798 8200 10864
rect 8266 10848 8272 10864
rect 8782 10848 8868 10882
rect 8266 10814 8908 10848
rect 8266 10798 8272 10814
rect 8782 10810 8816 10814
rect 8194 10796 8272 10798
rect 5338 10784 5344 10790
rect 3200 10650 3332 10768
rect 3426 10760 3500 10768
rect 4270 10714 4276 10766
rect 4328 10758 4334 10766
rect 4328 10720 4556 10758
rect 8066 10750 8144 10756
rect 4328 10714 4334 10720
rect 8066 10684 8072 10750
rect 8138 10734 8144 10750
rect 8138 10700 8908 10734
rect 11882 10722 11918 11290
rect 21514 11246 21520 11330
rect 21572 11310 24358 11330
rect 21572 11246 24366 11310
rect 21516 11242 21576 11246
rect 24174 11178 24366 11246
rect 16752 10894 16872 10916
rect 16752 10826 16778 10894
rect 16846 10826 16872 10894
rect 17472 10882 18518 10928
rect 18592 10882 20422 10928
rect 24186 10892 24366 11178
rect 16752 10804 16872 10826
rect 20364 10862 20422 10882
rect 21960 10862 22188 10878
rect 20364 10838 22188 10862
rect 20364 10822 22030 10838
rect 20364 10820 20422 10822
rect 8138 10684 8144 10700
rect 11728 10688 11918 10722
rect 17474 10718 18518 10762
rect 18592 10718 20234 10762
rect 8066 10680 8144 10684
rect 3200 10612 4556 10650
rect 5282 10638 5288 10644
rect 3200 10576 3500 10612
rect 5038 10598 5288 10638
rect 5282 10592 5288 10598
rect 5340 10638 5346 10644
rect 5340 10598 5364 10638
rect 10596 10602 10636 10626
rect 5340 10592 5346 10598
rect 3200 10574 3334 10576
rect 3200 10566 3332 10574
rect 3426 10568 3500 10576
rect 1240 9866 1494 9992
rect 1228 9114 1482 9292
rect 3200 9114 3274 10566
rect 4262 10522 4268 10574
rect 4320 10566 4326 10574
rect 4320 10528 4556 10566
rect 10596 10562 10666 10602
rect 10596 10558 10636 10562
rect 4320 10522 4326 10528
rect 10520 10518 10636 10558
rect 1228 9040 3274 9114
rect 3426 10420 4556 10458
rect 5280 10446 5286 10452
rect 1228 8916 1482 9040
rect 1240 8146 1494 8328
rect 3426 8146 3500 10420
rect 5038 10406 5286 10446
rect 5280 10400 5286 10406
rect 5338 10446 5344 10452
rect 5338 10406 5364 10446
rect 7944 10436 8022 10440
rect 5338 10400 5344 10406
rect 4270 10330 4276 10382
rect 4328 10374 4334 10382
rect 4328 10336 4556 10374
rect 7944 10370 7950 10436
rect 8016 10420 8022 10436
rect 8016 10386 8908 10420
rect 8016 10370 8022 10386
rect 7944 10366 8022 10370
rect 8798 10354 8868 10386
rect 4328 10330 4334 10336
rect 10586 10318 10660 10358
rect 10586 10208 10626 10318
rect 11794 10312 11940 10348
rect 20190 10342 20234 10718
rect 20714 10686 20806 10692
rect 20714 10606 20720 10686
rect 20800 10666 20806 10686
rect 21976 10666 22188 10682
rect 20800 10642 22188 10666
rect 23060 10642 23404 10682
rect 20800 10626 22030 10642
rect 23060 10626 23402 10642
rect 20800 10606 20806 10626
rect 20714 10602 20806 10606
rect 20916 10550 20988 10556
rect 23362 10536 23402 10626
rect 20988 10496 22188 10536
rect 23060 10496 23402 10536
rect 20916 10472 20988 10478
rect 20190 10340 20510 10342
rect 11794 10270 11830 10312
rect 20190 10300 22188 10340
rect 20190 10298 20510 10300
rect 23362 10286 23402 10496
rect 24180 10286 24360 10420
rect 13134 10280 13196 10282
rect 11716 10234 11830 10270
rect 13132 10278 13198 10280
rect 13132 10268 13138 10278
rect 13062 10258 13138 10268
rect 12416 10224 13138 10258
rect 13192 10224 13198 10278
rect 17628 10226 18518 10258
rect 12416 10214 13196 10224
rect 17622 10218 18518 10226
rect 18592 10238 22030 10258
rect 18592 10218 22188 10238
rect 10520 10168 10626 10208
rect 16540 10200 16652 10218
rect 7818 10130 7902 10132
rect 7818 10064 7824 10130
rect 7890 10114 7902 10130
rect 16540 10130 16564 10200
rect 16630 10130 16652 10200
rect 7890 10080 8798 10114
rect 7890 10064 7902 10080
rect 7818 10062 7902 10064
rect 8764 10044 8798 10080
rect 11814 10082 11924 10118
rect 16540 10110 16652 10130
rect 11814 10078 11850 10082
rect 11730 10046 11850 10078
rect 8764 10010 8868 10044
rect 10592 9896 10656 9984
rect 10592 9858 10632 9896
rect 10520 9818 10632 9858
rect 7706 9816 7784 9818
rect 7706 9750 7712 9816
rect 7778 9800 7784 9816
rect 7778 9766 8780 9800
rect 7778 9750 7784 9766
rect 7706 9748 7784 9750
rect 8748 9744 8780 9766
rect 8748 9684 8782 9744
rect 17622 9722 17668 10218
rect 21970 10198 22188 10218
rect 23362 10200 24360 10286
rect 21100 10084 21178 10088
rect 21098 10082 21180 10084
rect 21098 10004 21100 10082
rect 21178 10062 21180 10082
rect 23362 10062 23402 10200
rect 21178 10042 22030 10062
rect 21178 10022 22188 10042
rect 21178 10004 21180 10022
rect 21098 10002 21180 10004
rect 21984 10002 22188 10022
rect 23060 10002 23402 10062
rect 24180 10002 24360 10200
rect 21100 9998 21178 10002
rect 21264 9944 21344 9946
rect 21260 9892 21266 9944
rect 21342 9932 21348 9944
rect 23362 9932 23402 10002
rect 21342 9896 22030 9932
rect 23060 9896 23402 9932
rect 21342 9892 22188 9896
rect 21264 9890 21344 9892
rect 21960 9856 22188 9892
rect 23048 9868 23402 9896
rect 23048 9856 23400 9868
rect 8748 9650 8868 9684
rect 10578 9672 10654 9708
rect 16748 9688 16872 9706
rect 10578 9508 10614 9672
rect 11726 9582 11870 9618
rect 16748 9616 16782 9688
rect 16850 9616 16872 9688
rect 17472 9676 17668 9722
rect 17790 9696 18518 9736
rect 18592 9700 22030 9736
rect 18592 9696 22188 9700
rect 16748 9600 16872 9616
rect 10520 9468 10616 9508
rect 11834 9144 11870 9582
rect 17790 9556 17830 9696
rect 21978 9660 22188 9696
rect 17474 9526 17830 9556
rect 17474 9512 17824 9526
rect 23632 9184 23788 9190
rect 11834 9108 11942 9144
rect 23632 9042 23638 9184
rect 23780 9160 23788 9184
rect 24180 9160 24360 9344
rect 23780 9066 24360 9160
rect 23780 9042 23788 9066
rect 23632 9036 23788 9042
rect 18024 8966 18116 8970
rect 12462 8956 12526 8958
rect 18024 8956 18034 8966
rect 12462 8952 18034 8956
rect 12462 8896 12466 8952
rect 12522 8900 18034 8952
rect 12522 8896 12526 8900
rect 12462 8890 12526 8896
rect 18024 8892 18034 8900
rect 18108 8892 18116 8966
rect 24180 8926 24360 9066
rect 18024 8888 18116 8892
rect 18182 8848 18268 8852
rect 18182 8836 18188 8848
rect 15930 8834 18188 8836
rect 15930 8782 15936 8834
rect 15988 8784 18188 8834
rect 15988 8782 15994 8784
rect 18182 8774 18188 8784
rect 18262 8774 18268 8848
rect 18182 8770 18268 8774
rect 7584 8722 7658 8730
rect 7584 8656 7588 8722
rect 7654 8706 7658 8722
rect 7654 8672 8848 8706
rect 7654 8656 7658 8672
rect 7584 8650 7658 8656
rect 11818 8624 11854 8626
rect 11750 8602 11854 8624
rect 11750 8588 12220 8602
rect 11818 8566 12220 8588
rect 10534 8492 10654 8532
rect 7456 8404 7534 8406
rect 7456 8338 7462 8404
rect 7528 8388 7534 8404
rect 7528 8364 8848 8388
rect 18330 8382 18418 8386
rect 7528 8354 8868 8364
rect 18330 8362 18336 8382
rect 7528 8338 7534 8354
rect 7456 8336 7534 8338
rect 8790 8330 8868 8354
rect 18304 8326 18336 8362
rect 18328 8308 18336 8326
rect 18410 8308 18418 8382
rect 18328 8306 18418 8308
rect 18328 8294 18408 8306
rect 16162 8258 18408 8294
rect 10574 8252 10650 8254
rect 10570 8218 10650 8252
rect 10570 8182 10610 8218
rect 1240 8072 3500 8146
rect 10520 8142 10610 8182
rect 11766 8176 12232 8208
rect 11722 8172 12232 8176
rect 11722 8140 11802 8172
rect 19636 8166 19756 8174
rect 1240 7952 1494 8072
rect 7332 8028 7338 8094
rect 7404 8078 7410 8094
rect 7404 8044 8768 8078
rect 19636 8066 19642 8166
rect 19742 8162 19756 8166
rect 24180 8162 24360 8368
rect 19742 8068 24360 8162
rect 19742 8066 19756 8068
rect 19636 8058 19756 8066
rect 7404 8028 7410 8044
rect 8738 8030 8768 8044
rect 8738 8008 8772 8030
rect 8738 7974 8868 8008
rect 11726 7982 11806 7984
rect 11726 7954 11808 7982
rect 11726 7952 12228 7954
rect 11772 7918 12228 7952
rect 24180 7950 24360 8068
rect 10560 7862 10650 7888
rect 10560 7832 10658 7862
rect 10520 7822 10658 7832
rect 7210 7798 7294 7800
rect 7210 7732 7218 7798
rect 7284 7782 7294 7798
rect 10520 7792 10630 7822
rect 7284 7748 8772 7782
rect 7284 7732 7294 7748
rect 7210 7728 7294 7732
rect 8738 7650 8772 7748
rect 8738 7616 8868 7650
rect 10568 7578 10654 7624
rect 1228 7316 1482 7484
rect 10568 7482 10608 7578
rect 11764 7526 12224 7562
rect 11764 7524 11804 7526
rect 11722 7488 11804 7524
rect 10520 7442 10608 7482
rect 4262 7368 4324 7372
rect 4394 7368 4456 7372
rect 1228 7242 3168 7316
rect 4262 7274 4268 7368
rect 4320 7274 4396 7368
rect 4448 7274 5726 7368
rect 4262 7270 4324 7274
rect 4394 7270 4456 7274
rect 1228 7108 1482 7242
rect 3094 6972 3168 7242
rect 5632 7138 5726 7274
rect 10986 7340 11048 7344
rect 18514 7340 18604 7346
rect 10986 7258 10992 7340
rect 11044 7258 18522 7340
rect 18596 7258 18604 7340
rect 10986 7254 11048 7258
rect 18514 7254 18604 7258
rect 24186 7138 24366 7332
rect 3996 7120 4048 7126
rect 5632 7122 24366 7138
rect 4406 7112 4412 7116
rect 4048 7074 4412 7112
rect 3996 7062 4048 7068
rect 4406 7064 4412 7074
rect 4464 7112 4470 7116
rect 4758 7112 4764 7120
rect 4464 7074 4764 7112
rect 4464 7064 4470 7074
rect 4758 7066 4764 7074
rect 4818 7066 4824 7120
rect 5632 7044 19426 7122
rect 3886 6988 3892 7040
rect 3944 7032 3950 7040
rect 4274 7032 4280 7044
rect 3944 6994 4280 7032
rect 3944 6988 3950 6994
rect 4274 6992 4280 6994
rect 4332 7032 4338 7044
rect 4858 7032 4864 7040
rect 4332 6994 4864 7032
rect 4332 6992 4338 6994
rect 4858 6988 4864 6994
rect 4916 6988 4922 7040
rect 19418 7028 19426 7044
rect 19526 7044 24366 7122
rect 19526 7028 19532 7044
rect 19418 7020 19532 7028
rect 3094 6970 3500 6972
rect 3094 6934 3544 6970
rect 3094 6922 3824 6934
rect 3094 6898 4090 6922
rect 5154 6920 5214 6924
rect 5152 6916 5158 6920
rect 3426 6890 4090 6898
rect 3500 6878 4090 6890
rect 2026 6870 2180 6878
rect 2026 6738 2036 6870
rect 2168 6840 2180 6870
rect 4708 6872 5158 6916
rect 3426 6840 3504 6844
rect 2168 6832 3504 6840
rect 2168 6790 4088 6832
rect 2168 6766 3502 6790
rect 4708 6784 4752 6872
rect 5152 6868 5158 6872
rect 5210 6868 5216 6920
rect 24186 6914 24366 7044
rect 5154 6864 5214 6868
rect 8776 6856 8860 6890
rect 8776 6836 8852 6856
rect 8776 6792 8832 6836
rect 2168 6738 2180 6766
rect 3426 6762 3500 6766
rect 7082 6764 7164 6768
rect 2026 6730 2180 6738
rect 7082 6698 7090 6764
rect 7156 6748 7164 6764
rect 8776 6748 8830 6792
rect 7156 6714 8830 6748
rect 11728 6736 11790 6772
rect 7156 6698 7164 6714
rect 8776 6712 8810 6714
rect 7082 6696 7164 6698
rect 5030 6690 5088 6694
rect 5028 6682 5034 6690
rect 1240 6510 1494 6664
rect 4714 6644 5034 6682
rect 5028 6638 5034 6644
rect 5086 6638 5092 6690
rect 10512 6680 10634 6720
rect 11754 6700 12224 6736
rect 10594 6672 10634 6680
rect 5030 6634 5088 6638
rect 10594 6632 10678 6672
rect 11882 6574 12116 6604
rect 11870 6566 11926 6574
rect 1240 6436 2438 6510
rect 8764 6504 8860 6538
rect 11870 6514 11872 6566
rect 11924 6514 11926 6566
rect 15842 6552 15848 6562
rect 14886 6520 15848 6552
rect 11870 6508 11926 6514
rect 15842 6510 15848 6520
rect 15900 6510 15906 6562
rect 1240 6288 1494 6436
rect 2364 6104 2438 6436
rect 6950 6450 7028 6456
rect 6950 6384 6956 6450
rect 7022 6434 7028 6450
rect 8764 6446 8798 6504
rect 8764 6434 8796 6446
rect 7022 6402 8796 6434
rect 7022 6400 8726 6402
rect 7022 6384 7028 6400
rect 6950 6380 7028 6384
rect 10592 6370 10656 6402
rect 10512 6330 10656 6370
rect 15738 6366 15744 6376
rect 11750 6320 12108 6346
rect 14886 6334 15744 6366
rect 15738 6324 15744 6334
rect 15796 6324 15802 6376
rect 11722 6310 12108 6320
rect 11722 6280 11786 6310
rect 11722 6264 11758 6280
rect 3892 6258 3950 6260
rect 3890 6206 3896 6258
rect 3948 6254 3954 6258
rect 3948 6210 4090 6254
rect 3948 6206 3954 6210
rect 3892 6202 3950 6206
rect 4944 6168 5008 6172
rect 4944 6162 4950 6168
rect 4710 6120 4950 6162
rect 4944 6116 4950 6120
rect 5002 6116 5008 6168
rect 8748 6142 8860 6176
rect 8748 6134 8782 6142
rect 4944 6112 5008 6116
rect 6828 6126 6902 6128
rect 8748 6126 8780 6134
rect 6828 6122 8780 6126
rect 2364 6068 3554 6104
rect 2364 6054 3568 6068
rect 3846 6054 4090 6056
rect 5282 6054 5340 6058
rect 6828 6056 6832 6122
rect 6898 6092 8780 6122
rect 11732 6098 11772 6130
rect 6898 6056 6902 6092
rect 2364 6030 4090 6054
rect 5280 6048 5286 6054
rect 3426 6022 4090 6030
rect 3498 6012 4090 6022
rect 4710 6006 5286 6048
rect 3072 5908 3154 5912
rect 3426 5908 3824 5912
rect 1240 5682 1494 5846
rect 3072 5834 3078 5908
rect 3152 5900 3824 5908
rect 3152 5856 4090 5900
rect 3152 5834 3502 5856
rect 4710 5842 4752 6006
rect 5280 6002 5286 6006
rect 5338 6002 5344 6054
rect 6828 6050 6902 6056
rect 11736 6088 11772 6098
rect 19194 6090 19304 6092
rect 11736 6052 12114 6088
rect 10512 6016 10650 6020
rect 5282 5998 5340 6002
rect 10512 5980 10666 6016
rect 10608 5962 10666 5980
rect 11992 6010 12056 6014
rect 11992 5958 11998 6010
rect 12050 6006 12056 6010
rect 12050 5964 12114 6006
rect 15644 5998 15650 6008
rect 14886 5966 15650 5998
rect 12050 5958 12084 5964
rect 11992 5950 12084 5958
rect 15644 5956 15650 5966
rect 15702 5956 15708 6008
rect 19194 5990 19200 6090
rect 19300 6086 19306 6090
rect 24180 6086 24360 6316
rect 19300 5992 24360 6086
rect 19300 5990 19306 5992
rect 19194 5986 19304 5990
rect 24180 5898 24360 5992
rect 6690 5834 6768 5838
rect 3072 5830 3154 5834
rect 3426 5830 3500 5834
rect 6690 5768 6696 5834
rect 6762 5818 6768 5834
rect 8730 5818 8860 5832
rect 6762 5798 8860 5818
rect 15544 5812 15550 5822
rect 6762 5784 8788 5798
rect 10604 5786 10664 5794
rect 6762 5768 6768 5784
rect 8754 5780 8788 5784
rect 6690 5764 6768 5768
rect 10602 5738 10664 5786
rect 14886 5780 15550 5812
rect 15544 5770 15550 5780
rect 15602 5770 15608 5822
rect 2026 5698 2186 5710
rect 2026 5682 2044 5698
rect 1240 5582 2044 5682
rect 1240 5470 1494 5582
rect 2026 5566 2044 5582
rect 2176 5566 2186 5698
rect 10602 5670 10642 5738
rect 11784 5670 12110 5696
rect 10512 5630 10642 5670
rect 11722 5660 12110 5670
rect 11722 5634 11820 5660
rect 2026 5556 2186 5566
rect 11872 5548 11936 5550
rect 10550 5488 10556 5540
rect 10608 5530 10614 5540
rect 11872 5530 11878 5548
rect 10608 5498 11878 5530
rect 10608 5488 10614 5498
rect 11872 5496 11878 5498
rect 11930 5496 11936 5548
rect 11872 5494 11936 5496
rect 12078 5546 12142 5588
rect 12078 5494 12084 5546
rect 12136 5526 12142 5546
rect 14202 5550 14284 5552
rect 14202 5530 14208 5550
rect 12808 5526 14208 5530
rect 12136 5498 14208 5526
rect 12136 5494 12142 5498
rect 12078 5492 12142 5494
rect 12792 5484 14208 5498
rect 11990 5482 12046 5484
rect 10444 5472 10510 5476
rect 10442 5414 10448 5472
rect 10506 5456 10512 5472
rect 11592 5466 11656 5468
rect 11592 5456 11598 5466
rect 10506 5424 11598 5456
rect 10506 5414 10512 5424
rect 11592 5414 11598 5424
rect 11650 5414 11656 5466
rect 11986 5464 11992 5482
rect 11980 5432 11992 5464
rect 11986 5430 11992 5432
rect 12044 5464 12050 5482
rect 14202 5480 14208 5484
rect 14278 5480 14284 5550
rect 14202 5478 14284 5480
rect 20232 5534 20344 5538
rect 12434 5464 12440 5470
rect 12044 5432 12440 5464
rect 12044 5430 12050 5432
rect 11990 5428 12046 5430
rect 12434 5418 12440 5432
rect 12492 5418 12498 5470
rect 20232 5434 20238 5534
rect 20338 5524 20344 5534
rect 22776 5534 22912 5536
rect 22776 5524 22798 5534
rect 20338 5442 22798 5524
rect 20338 5434 20344 5442
rect 20232 5432 20344 5434
rect 22776 5432 22798 5442
rect 22900 5524 22912 5534
rect 24282 5524 24414 5652
rect 22900 5442 24414 5524
rect 22900 5432 22912 5442
rect 22776 5430 22912 5432
rect 24282 5422 24414 5442
rect 12438 5416 12494 5418
rect 10442 5410 10512 5414
rect 12836 5386 12892 5392
rect 9558 5374 9624 5380
rect 9558 5312 9560 5374
rect 9622 5332 9624 5374
rect 10730 5358 10790 5360
rect 10728 5332 10734 5358
rect 9622 5312 10734 5332
rect 9558 5306 10734 5312
rect 10786 5332 10792 5358
rect 12836 5334 12838 5386
rect 12890 5334 12892 5386
rect 12836 5332 12892 5334
rect 13642 5382 13702 5388
rect 13642 5332 13646 5382
rect 10786 5328 13646 5332
rect 13700 5328 13702 5382
rect 10786 5322 13700 5328
rect 10786 5306 13688 5322
rect 9558 5300 13688 5306
rect 10320 5256 10408 5258
rect 1256 5254 10408 5256
rect 1256 5172 10322 5254
rect 8950 5170 9046 5172
rect 10316 5170 10322 5172
rect 10406 5170 10412 5254
rect 12194 5234 12270 5240
rect 15410 5238 15470 5242
rect 10320 5168 10408 5170
rect 12194 5168 12200 5234
rect 12266 5168 12270 5234
rect 12194 5162 12270 5168
rect 12424 5154 12430 5222
rect 12498 5154 12504 5222
rect 14142 5190 14274 5194
rect 14142 5126 14216 5190
rect 14268 5126 14274 5190
rect 15268 5170 15414 5238
rect 15466 5170 15472 5238
rect 15410 5166 15472 5170
rect 14142 5122 14274 5126
rect 1252 4978 5038 5062
rect 5090 5038 9552 5062
rect 5090 4978 5888 5038
rect 5862 4896 5888 4978
rect 6004 4978 9552 5038
rect 9636 4978 9648 5062
rect 14492 5060 14582 5064
rect 10454 5024 10530 5030
rect 6004 4896 6028 4978
rect 10454 4960 10458 5024
rect 10522 4960 10530 5024
rect 14492 4984 14500 5060
rect 14576 4984 14582 5060
rect 14492 4978 14582 4984
rect 18984 5030 19104 5036
rect 10454 4954 10530 4960
rect 18984 4930 18990 5030
rect 19090 5026 19104 5030
rect 24266 5026 24686 5214
rect 19090 4932 24686 5026
rect 19090 4930 19104 4932
rect 18984 4924 19104 4930
rect 5862 4878 6028 4896
rect 1228 4660 1482 4816
rect 24266 4798 24686 4932
rect 24270 4796 24424 4798
rect 3074 4660 3156 4664
rect 1228 4586 3076 4660
rect 3150 4586 3156 4660
rect 15838 4628 15844 4728
rect 15896 4628 27146 4728
rect 1228 4440 1482 4586
rect 3074 4582 3156 4586
rect 4580 4574 4638 4578
rect 5026 4574 5088 4578
rect 4578 4502 4584 4574
rect 4636 4502 5030 4574
rect 5082 4502 5088 4574
rect 25926 4548 26328 4552
rect 4580 4498 4638 4502
rect 5026 4498 5088 4502
rect 15730 4448 15736 4548
rect 15788 4448 26328 4548
rect 15636 4268 15642 4368
rect 15694 4364 25490 4368
rect 15694 4268 25512 4364
rect 15540 4088 15546 4188
rect 15598 4186 24698 4188
rect 15598 4088 24740 4186
rect 11258 4070 13438 4072
rect 11258 4066 11410 4070
rect 11256 4010 11262 4066
rect 11318 4016 11410 4066
rect 11318 4010 11324 4016
rect 11404 4014 11410 4016
rect 11466 4066 13438 4070
rect 11466 4016 13224 4066
rect 11466 4014 11472 4016
rect 13218 4010 13224 4016
rect 13280 4016 13438 4066
rect 13280 4010 13286 4016
rect 3418 3982 3492 3984
rect 1240 3818 1494 3958
rect 3154 3906 3676 3982
rect 10472 3908 10572 3910
rect 19658 3908 19664 3912
rect 3154 3818 3230 3906
rect 3418 3902 3492 3906
rect 10472 3896 19664 3908
rect 5152 3842 5208 3844
rect 1240 3742 3230 3818
rect 4434 3776 5154 3842
rect 5206 3776 5212 3842
rect 10472 3804 10478 3896
rect 10570 3816 19664 3896
rect 10570 3804 10576 3816
rect 19658 3812 19664 3816
rect 19764 3812 19770 3912
rect 10472 3800 10572 3804
rect 5152 3772 5208 3776
rect 1240 3582 1494 3742
rect 12134 3714 19550 3726
rect 12134 3706 19426 3714
rect 12134 3634 12154 3706
rect 12148 3614 12154 3634
rect 12246 3634 19426 3706
rect 12246 3614 12252 3634
rect 19420 3622 19426 3634
rect 19526 3634 19550 3714
rect 19526 3622 19532 3634
rect 12422 3540 19332 3544
rect 12422 3530 19200 3540
rect 12420 3528 19200 3530
rect 3668 3454 3674 3512
rect 3732 3506 3738 3512
rect 4944 3510 5010 3518
rect 4942 3506 4948 3510
rect 3732 3454 4948 3506
rect 3676 3452 4948 3454
rect 5006 3506 5012 3510
rect 5006 3452 5674 3506
rect 3676 3448 5674 3452
rect 4944 3444 5010 3448
rect 4436 3370 4904 3380
rect 4436 3260 4716 3370
rect 4710 3250 4716 3260
rect 4836 3312 4904 3370
rect 4836 3264 4912 3312
rect 4836 3260 4904 3264
rect 4836 3250 4842 3260
rect 4710 3246 4842 3250
rect 4716 3244 4836 3246
rect 5614 3032 5672 3448
rect 12420 3436 12440 3528
rect 12532 3452 19200 3528
rect 12532 3436 12550 3452
rect 19194 3448 19200 3452
rect 19300 3452 19332 3540
rect 19300 3448 19306 3452
rect 12420 3426 12550 3436
rect 14110 3356 14214 3360
rect 19008 3356 19014 3358
rect 14110 3346 19014 3356
rect 14110 3254 14118 3346
rect 14210 3266 19014 3346
rect 19114 3356 19120 3358
rect 19114 3266 19138 3356
rect 14210 3264 19138 3266
rect 14210 3254 14216 3264
rect 14110 3244 14214 3254
rect 8898 3032 8962 3036
rect 20098 3032 20330 3038
rect 1240 2772 1494 2954
rect 5576 2808 8904 3032
rect 8956 3028 20122 3032
rect 8956 3024 13140 3028
rect 8956 3020 11326 3024
rect 8956 2808 11178 3020
rect 8898 2804 8962 2808
rect 11172 2796 11178 2808
rect 11550 2808 13140 3024
rect 11550 2800 11556 2808
rect 11402 2796 11556 2800
rect 11172 2792 11556 2796
rect 13134 2790 13140 2808
rect 13512 2808 20122 3028
rect 20310 2808 20330 3032
rect 13512 2790 13520 2808
rect 20098 2802 20330 2808
rect 13134 2786 13520 2790
rect 1240 2696 3234 2772
rect 1240 2578 1494 2696
rect 3158 2526 3234 2696
rect 3418 2526 3492 2528
rect 3158 2450 3702 2526
rect 3418 2446 3492 2450
rect 5268 2332 5330 2336
rect 4422 2264 5272 2332
rect 5324 2264 5330 2332
rect 5268 2260 5330 2264
rect 1482 2154 1582 2164
rect 1482 2076 1490 2154
rect 1568 2142 1582 2154
rect 15276 2148 15354 2150
rect 15274 2142 15280 2148
rect 1568 2086 15280 2142
rect 1568 2076 1582 2086
rect 15274 2082 15280 2086
rect 15346 2082 15354 2148
rect 15276 2080 15354 2082
rect 1482 2070 1582 2076
rect 8558 2016 8642 2018
rect 8558 1950 8568 2016
rect 8634 1966 16612 2016
rect 8634 1950 16614 1966
rect 8558 1948 8642 1950
rect 15406 1946 16614 1950
rect 8438 1892 8514 1894
rect 1214 1470 1468 1846
rect 8438 1826 8444 1892
rect 8510 1826 15798 1892
rect 8438 1824 8514 1826
rect 14584 1824 15798 1826
rect 8310 1766 8394 1768
rect 8310 1700 8318 1766
rect 8384 1700 14982 1766
rect 8310 1698 8394 1700
rect 8192 1640 8272 1642
rect 8192 1574 8198 1640
rect 8264 1638 8272 1640
rect 8264 1574 14180 1638
rect 8192 1572 14180 1574
rect 8192 1570 8272 1572
rect 8060 1504 8142 1506
rect 8058 1438 8070 1504
rect 8136 1438 13362 1504
rect 8060 1434 8142 1438
rect 7944 1380 8026 1382
rect 7944 1314 7950 1380
rect 8016 1376 12558 1380
rect 8016 1314 12560 1376
rect 7944 1312 8026 1314
rect 7824 1186 7830 1252
rect 7896 1250 7902 1252
rect 7896 1186 11762 1250
rect 7844 1184 11762 1186
rect 6680 1088 6788 1094
rect 6680 1086 6690 1088
rect 4114 1078 6690 1086
rect 4104 1002 6690 1078
rect 6776 1002 6788 1088
rect 7708 1072 7714 1138
rect 7780 1128 7786 1138
rect 7780 1072 10980 1128
rect 7760 1062 10980 1072
rect 4104 1000 6788 1002
rect 1228 520 1482 896
rect 4104 624 4506 1000
rect 6680 994 6788 1000
rect 7592 934 7598 1000
rect 7664 934 10140 1000
rect 6810 930 6918 932
rect 6810 918 6820 930
rect 4924 844 6820 918
rect 6906 844 6918 930
rect 8914 874 9318 878
rect 7482 872 9324 874
rect 4924 832 6918 844
rect 4924 630 5320 832
rect 7462 806 7468 872
rect 7534 808 9324 872
rect 7534 806 7540 808
rect 6946 788 7044 796
rect 6946 756 6954 788
rect 5824 752 6954 756
rect 5710 708 6954 752
rect 7034 708 7044 788
rect 5710 696 7044 708
rect 5710 676 7026 696
rect 7334 676 7340 744
rect 7406 676 8530 744
rect 5710 630 6106 676
rect 6912 630 7042 632
rect 4100 492 4506 624
rect 4914 498 5320 630
rect 5706 498 6112 630
rect 6506 622 7042 630
rect 6506 520 6920 622
rect 7022 520 7042 622
rect 7212 626 7322 630
rect 7212 622 7722 626
rect 8124 624 8532 676
rect 7212 548 7224 622
rect 7298 548 7722 622
rect 7212 540 7722 548
rect 6506 504 7042 520
rect 6506 498 6912 504
rect 7316 494 7722 540
rect 8122 492 8532 624
rect 8908 498 9324 808
rect 9730 674 10136 934
rect 9730 616 10138 674
rect 9732 494 10138 616
rect 10566 498 10972 1062
rect 11364 642 11762 1184
rect 11362 492 11768 642
rect 12160 638 12560 1314
rect 12154 498 12560 638
rect 12980 624 13362 1438
rect 13788 628 14178 1572
rect 14584 628 14982 1700
rect 15406 1760 15798 1824
rect 16226 1846 16614 1946
rect 20730 1924 20816 1928
rect 17030 1918 17422 1924
rect 20726 1918 20732 1924
rect 17030 1848 20732 1918
rect 15406 628 15796 1760
rect 16226 632 16612 1846
rect 12964 494 13370 624
rect 13778 498 14184 628
rect 14584 498 14990 628
rect 15394 498 15800 628
rect 16208 476 16614 632
rect 17030 628 17422 1848
rect 20726 1844 20732 1848
rect 20812 1844 20818 1924
rect 20730 1842 20816 1844
rect 20910 1762 20996 1766
rect 20908 1760 20914 1762
rect 17816 1684 20914 1760
rect 20992 1684 20998 1762
rect 17024 498 17430 628
rect 17816 624 18208 1684
rect 20910 1680 20996 1684
rect 21094 1596 21100 1598
rect 18646 1520 21100 1596
rect 21178 1520 21184 1598
rect 18646 628 19042 1520
rect 21262 1438 21346 1444
rect 19468 1362 21264 1438
rect 21340 1362 21346 1438
rect 17814 494 18220 624
rect 18638 498 19044 628
rect 19468 622 19864 1362
rect 21262 1356 21346 1362
rect 20482 764 21730 804
rect 20482 628 20522 764
rect 21914 722 21954 804
rect 21468 682 21954 722
rect 21468 628 21508 682
rect 22108 628 22150 806
rect 19466 492 19872 622
rect 20264 498 20670 628
rect 21068 568 21508 628
rect 21068 498 21474 568
rect 21884 498 22290 628
rect 22494 610 22536 806
rect 22688 768 22726 802
rect 22688 730 23688 768
rect 23650 638 23688 730
rect 22720 610 23126 628
rect 23650 624 23856 638
rect 24338 628 24740 4088
rect 22494 568 23126 610
rect 22720 498 23126 568
rect 23516 494 23922 624
rect 24326 524 24740 628
rect 25110 628 25512 4268
rect 24326 498 24732 524
rect 25110 498 25524 628
rect 25926 624 26328 4448
rect 26744 628 27146 4628
rect 25110 490 25512 498
rect 25926 494 26334 624
rect 26738 512 27146 628
rect 26738 498 27144 512
rect 25926 478 26328 494
<< via2 >>
rect 16556 11582 16620 11588
rect 16556 11530 16602 11582
rect 16602 11530 16620 11582
rect 16762 11584 16826 11586
rect 16762 11532 16806 11584
rect 16806 11532 16826 11584
rect 16556 11524 16620 11530
rect 16762 11522 16826 11532
rect 16778 10826 16846 10894
rect 16564 10130 16630 10200
rect 16782 9616 16850 9688
<< metal3 >>
rect 16542 11588 16632 11600
rect 16542 11524 16556 11588
rect 16620 11524 16632 11588
rect 16542 11450 16632 11524
rect 16750 11586 16840 11598
rect 16750 11522 16762 11586
rect 16826 11522 16840 11586
rect 16542 10218 16616 11450
rect 16750 11448 16840 11522
rect 16766 10920 16840 11448
rect 16766 10894 16854 10920
rect 16766 10826 16778 10894
rect 16846 10826 16854 10894
rect 16766 10800 16854 10826
rect 16542 10200 16640 10218
rect 16542 10152 16564 10200
rect 16552 10130 16564 10152
rect 16630 10130 16640 10200
rect 16552 10120 16640 10130
rect 16766 9778 16840 10800
rect 16764 9688 16858 9778
rect 16764 9616 16782 9688
rect 16850 9616 16858 9688
rect 16764 9604 16858 9616
use sky130_hilas_nFETLarge  sky130_hilas_nFETLarge_0
timestamp 1632255311
transform -1 0 4676 0 -1 5734
box 0 0 1114 1206
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_0
timestamp 1632256357
transform -1 0 4684 0 -1 4224
box 0 0 1016 1214
use sky130_hilas_nFETLarge  sky130_hilas_nFETLarge_1
timestamp 1632255311
transform -1 0 15530 0 1 3278
box 0 0 1114 1206
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_4
timestamp 1632256357
transform -1 0 14382 0 1 3280
box 0 0 1016 1214
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_1
timestamp 1632256357
transform 1 0 10308 0 1 3274
box 0 0 1016 1214
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_2
timestamp 1632256357
transform -1 0 12420 0 1 3274
box 0 0 1016 1214
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_3
timestamp 1632256357
transform 1 0 12270 0 1 3280
box 0 0 1016 1214
use sky130_hilas_DAC5bit01  sky130_hilas_DAC5bit01_0
timestamp 1632255311
transform 0 1 20484 1 0 0
box 0 0 3398 1638
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_1
timestamp 1632256361
transform -1 0 10514 0 -1 10568
box 0 0 1778 1574
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_2
timestamp 1632256361
transform -1 0 10514 0 -1 8542
box 0 0 1778 1574
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_3
timestamp 1632256361
transform -1 0 10506 0 -1 6730
box 0 0 1778 1574
use sky130_hilas_Trans2med  sky130_hilas_Trans2med_0
timestamp 1632256353
transform 1 0 4806 0 -1 6684
box 0 0 936 1186
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_2
timestamp 1632256352
transform -1 0 13858 0 -1 8658
box 0 0 1600 1228
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_3
timestamp 1632256352
transform -1 0 13864 0 -1 6804
box 0 0 1600 1228
use sky130_hilas_TA2Cell_1FG  sky130_hilas_TA2Cell_1FG_0
timestamp 1632256356
transform 1 0 17132 0 1 8728
box 0 0 8180 4664
use sky130_hilas_swc4x2cell  sky130_hilas_swc4x2cell_0
timestamp 1632256358
transform 1 0 14190 0 1 7466
box 0 0 9144 2944
use sky130_hilas_WTA4Stage01  sky130_hilas_WTA4Stage01_0
timestamp 1632256350
transform 1 0 14310 0 1 5670
box 0 0 5596 2974
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_0
timestamp 1632256361
transform -1 0 10514 0 1 11014
box 0 0 1778 1574
use sky130_hilas_FGcharacterization01  sky130_hilas_FGcharacterization01_0
timestamp 1632256360
transform -1 0 6024 0 1 12678
box 0 0 6024 2834
use sky130_hilas_Trans4small  sky130_hilas_Trans4small_0
timestamp 1632256349
transform 1 0 4136 0 1 10580
box 0 0 694 1292
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_1
timestamp 1632256352
transform -1 0 13862 0 -1 10752
box 0 0 1600 1228
use sky130_hilas_TA2Cell_1FG_Strong  sky130_hilas_TA2Cell_1FG_Strong_0
timestamp 1632256354
transform 1 0 17132 0 1 9934
box 0 0 9388 4664
use sky130_hilas_Tgate4Single01  sky130_hilas_Tgate4Single01_0
timestamp 1632256348
transform 1 0 22220 0 1 9956
box 0 0 1492 2094
<< labels >>
rlabel metal2 26738 498 27144 628 1 DIG24 
port 1 n
rlabel metal2 25928 494 26334 624 0 DIG23
port 2 nsew
rlabel metal2 25118 498 25524 628 0 DIG22
port 3 nsew
rlabel metal2 24326 498 24732 628 0 DIG21
port 4 nsew
rlabel metal2 23516 494 23922 624 0 DIG29
port 5 nsew
rlabel metal2 22720 498 23126 628 0 DIG28
port 6 nsew
rlabel metal2 21884 498 22290 628 0 DIG27
port 7 nsew
rlabel metal2 21068 498 21474 628 0 DIG26
port 8 nsew
rlabel metal2 20264 498 20670 628 0 DIG25
port 9 nsew
rlabel metal2 19466 492 19872 622 0 DIG20
port 10 nsew
rlabel metal2 18638 498 19044 628 0 DIG19
port 11 nsew
rlabel metal2 17814 494 18220 624 0 DIG18
port 12 nsew
rlabel metal2 17024 498 17430 628 0 DIG17
port 13 nsew
rlabel metal2 16208 502 16614 632 0 DIG16
port 14 nsew
rlabel metal2 15394 498 15800 628 0 DIG15
port 15 nsew
rlabel metal2 14584 498 14990 628 0 DIG14
port 16 nsew
rlabel metal2 13778 498 14184 628 0 DIG13
port 17 nsew
rlabel metal2 12964 494 13370 624 0 DIG12
port 18 nsew
rlabel metal2 12154 506 12560 638 0 DIG11
port 19 nsew
rlabel metal2 11362 510 11768 642 0 DIG10
port 20 nsew
rlabel metal2 10566 498 10972 630 0 DIG09
port 21 nsew
rlabel metal2 9732 494 10138 626 0 DIG08
port 22 nsew
rlabel metal2 8914 498 9320 630 0 DIG07
port 23 nsew
rlabel metal2 8122 492 8528 624 0 DIG06
port 24 nsew
rlabel metal2 7316 494 7722 626 0 DIG05
port 25 nsew
rlabel metal2 6506 498 6912 630 0 DIG04
port 26 nsew
rlabel metal2 5706 498 6112 630 0 DIG03
port 27 nsew
rlabel metal2 4914 498 5320 630 0 DIG02
port 28 nsew
rlabel metal2 4100 492 4506 624 0 DIG01
port 29 nsew
rlabel metal2 24270 4796 24424 5214 0 CAP2    
port 30 nsew
rlabel metal2 24180 5898 24360 6316 0 GENERALGATE01   
port 31 nsew
rlabel metal2 24186 6914 24366 7332 0 GATEANDCAP1    
port 32 nsew
rlabel metal2 24180 7950 24360 8368 0 GENERALGATE02
port 33 nsew
rlabel metal2 24180 8926 24360 9344 0 OUTPUTTA1    
port 34 nsew
rlabel metal2 24180 10002 24360 10420 0 GATENFET1   
port 35 nsew
rlabel metal2 24186 10892 24366 11310 0 DACOUTPUT  
port 36 nsew
rlabel metal2 24188 11768 24360 12188 0 DRAINOUT
port 37 nsew
rlabel metal2 24188 12646 24360 13066 0 ROWTERM2
port 38 nsew
rlabel metal2 24194 13464 24366 13884 0 COLUMN2
port 39 nsew
rlabel metal2 24194 14290 24366 14710 0 COLUMN1
port 40 nsew
rlabel metal1 21206 14636 21844 14860 0 GATE2
port 41 nsew
rlabel metal1 15492 14630 16130 14854 0 GATE1
port 61 nsew
rlabel metal1 9774 14632 10412 14856 0 DRAININJECT
port 42 nsew
rlabel metal1 6712 14538 6980 14740 0 VTUN
port 43 nsew
rlabel metal2 1250 14334 1386 14798 0 VREFCHAR
port 44 nsew
rlabel metal2 1250 13428 1386 13892 0 CHAROUTPUT
port 45 nsew
rlabel metal2 1160 12534 1296 12998 0 LARGECAPACITOR
port 46 nsew
rlabel metal2 3418 3902 3492 3984 0 DRAIN6N
port 47 nsew
rlabel metal2 3418 2446 3492 2528 0 DRAIN6P
port 48 nsew
rlabel metal2 3426 5830 3500 5912 0 DRAIN5P
port 49 nsew
rlabel metal2 3426 6022 3500 6104 0 DARIN4P
port 50 nsew
rlabel metal2 3426 6762 3500 6844 0 DRAIN5N
port 51 nsew
rlabel metal2 3426 6890 3500 6972 0 DRAIN4N
port 52 nsew
rlabel metal2 3426 10376 3500 10458 0 DRAIN3P
port 53 nsew
rlabel metal2 3426 10568 3500 10650 0 DRAIN2P
port 54 nsew
rlabel metal2 3426 10760 3500 10842 0 DRAIN1P
port 55 nsew
rlabel metal2 3426 10984 3500 11066 0 DRAIN3N
port 56 nsew
rlabel metal2 3426 11170 3500 11252 0 DRAIN2N
port 57 nsew
rlabel metal2 3426 11376 3500 11458 0 DRAIN1N
port 58 nsew
rlabel metal2 3366 11592 3426 11672 0 SOURCEN
port 59 nsew
rlabel metal2 3366 11756 3426 11836 0 SOURCEP
port 60 nsew
rlabel metal2 1218 13154 1308 13234 0 VGND
port 63 nsew
rlabel metal2 1226 14036 1316 14116 0 VINJ
port 62 nsew
rlabel metal2 1160 12376 1262 12458 0 VINJ
port 62 nsew
rlabel metal2 1152 12196 1254 12278 0 VGND
port 63 nsew
rlabel metal2 1256 5172 1382 5256 0 VINJ
port 62 nsew
rlabel metal2 1252 4978 1378 5062 0 VGND
port 63 nsew
rlabel metal2 24386 11502 24476 11592 0 VPWR
port 64 nsew
rlabel metal1 11936 14804 12082 14864 0 VINJ
port 62 nsew
rlabel metal1 12968 14822 13162 14864 0 VGND
port 63 nsew
rlabel metal2 24282 5422 24414 5652 0 VPWR
port 64 nsew
rlabel metal1 11060 492 11244 638 0 VPWR
port 64 nsew
rlabel metal1 13446 492 13630 638 0 VPWR
port 64 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
