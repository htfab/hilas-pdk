magic
tech sky130A
timestamp 1628707289
<< checkpaint >>
rect -331 19898 2016 20643
rect -560 -630 2016 19898
rect -560 -1375 1787 -630
<< metal1 >>
rect 1 17663 72 18059
rect 1156 17181 1228 17570
rect 0 14803 70 15199
rect 1156 14322 1228 14711
rect 2 11944 72 12340
rect 1156 11462 1228 11851
rect 0 9085 70 9481
rect 1156 8605 1228 8994
rect 0 6225 70 6621
rect 1155 5745 1227 6134
rect 1 3367 71 3763
rect 1156 2886 1228 3275
rect 1 507 71 903
rect 1156 26 1228 415
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_12
timestamp 1628705751
transform 0 1 299 1 0 17154
box 0 0 2859 1087
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_11
timestamp 1628705751
transform 0 1 299 1 0 14295
box 0 0 2859 1087
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_10
timestamp 1628705751
transform 0 1 299 1 0 11436
box 0 0 2859 1087
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_5
timestamp 1628705751
transform 0 1 299 1 0 8577
box 0 0 2859 1087
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_8
timestamp 1628705751
transform 0 1 299 1 0 5718
box 0 0 2859 1087
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_7
timestamp 1628705751
transform 0 1 299 1 0 2859
box 0 0 2859 1087
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_9
timestamp 1628705751
transform 0 1 299 1 0 0
box 0 0 2859 1087
<< labels >>
rlabel metal1 1156 26 1228 415 0 IO7
port 1 nsew
rlabel metal1 1156 2886 1228 3275 0 IO8
port 2 nsew
rlabel metal1 1155 5745 1227 6134 0 IO9
port 3 nsew
rlabel metal1 1156 8605 1228 8994 0 IO10
port 4 nsew
rlabel metal1 1156 11462 1228 11851 0 IO11
port 5 nsew
rlabel metal1 1156 14322 1228 14711 0 IO12
port 7 nsew
rlabel metal1 1156 17181 1228 17570 0 IO13
port 6 nsew
rlabel metal1 1 507 71 903 0 PIN1
port 8 nsew
rlabel metal1 1 3367 71 3763 0 PIN2
port 9 nsew
rlabel metal1 0 6225 70 6621 0 PIN3
port 10 nsew
rlabel metal1 0 9085 70 9481 0 PIN4
port 11 nsew
rlabel metal1 2 11944 72 12340 0 PIN5
port 12 nsew
rlabel metal1 0 14803 70 15199 0 PIN6
port 13 nsew
rlabel metal1 1 17663 71 18059 0 PIN7
port 14 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
