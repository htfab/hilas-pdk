VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_wtasinglestage01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_wtasinglestage01 ;
  ORIGIN 1.080 0.760 ;
  SIZE 2.830 BY 1.430 ;
  OBS
      LAYER li1 ;
        RECT 0.110 0.610 0.320 0.630 ;
        RECT 0.090 0.440 0.760 0.610 ;
        RECT 0.090 0.210 0.340 0.440 ;
        RECT -0.500 -0.300 -0.160 0.210 ;
        RECT 0.010 0.040 0.340 0.210 ;
        RECT 0.560 0.040 0.900 0.210 ;
        RECT 0.090 -0.130 0.260 0.040 ;
        RECT 0.650 -0.130 0.820 0.040 ;
        RECT 0.010 -0.300 0.340 -0.130 ;
        RECT 0.560 -0.300 0.900 -0.130 ;
        RECT 0.650 -0.530 0.820 -0.300 ;
        RECT 1.220 -0.380 1.730 0.290 ;
        RECT -0.640 -0.700 0.820 -0.530 ;
      LAYER mcon ;
        RECT 0.130 0.440 0.300 0.610 ;
        RECT 1.390 -0.130 1.560 0.040 ;
      LAYER met1 ;
        RECT 0.100 -0.760 0.330 0.670 ;
        RECT 1.360 -0.760 1.590 0.530 ;
      LAYER met2 ;
        RECT -0.540 -0.020 1.750 0.140 ;
        RECT -1.080 -0.720 -0.960 -0.510 ;
  END
END sky130_hilas_wtasinglestage01
END LIBRARY

