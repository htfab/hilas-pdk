VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_fgbias2x1cell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_fgbias2x1cell ;
  ORIGIN 3.960 3.820 ;
  SIZE 11.530 BY 6.050 ;
  OBS
      LAYER nwell ;
        RECT 4.260 2.220 7.570 2.230 ;
        RECT -3.370 -2.420 -2.810 0.000 ;
      LAYER li1 ;
        RECT 4.670 0.280 4.700 0.450 ;
        RECT -0.920 -0.750 -0.730 -0.340 ;
        RECT 4.670 -0.510 4.720 -0.340 ;
        RECT -0.920 -0.930 2.630 -0.750 ;
        RECT -0.920 -1.350 -0.730 -0.930 ;
        RECT 4.740 -1.080 4.910 -0.510 ;
        RECT 4.670 -1.250 4.690 -1.080 ;
        RECT 0.110 -1.970 0.340 -1.930 ;
        RECT 4.670 -2.040 4.700 -1.870 ;
      LAYER met1 ;
        RECT -3.610 -3.810 -3.190 2.230 ;
        RECT -1.130 -3.820 -0.900 2.230 ;
        RECT 0.090 -3.820 0.320 2.230 ;
        RECT 6.610 2.220 6.800 2.230 ;
        RECT 7.050 -3.820 7.330 2.230 ;
      LAYER met2 ;
        RECT 4.840 1.730 5.160 1.750 ;
        RECT -3.960 1.550 5.160 1.730 ;
        RECT 5.540 0.490 7.570 0.710 ;
        RECT 6.220 -0.980 7.400 -0.630 ;
        RECT 5.530 -2.260 7.570 -2.050 ;
        RECT 5.100 -3.150 5.260 -3.130 ;
        RECT -3.940 -3.200 5.260 -3.150 ;
        RECT -3.940 -3.300 5.140 -3.200 ;
  END
END sky130_hilas_fgbias2x1cell
END LIBRARY

