magic
tech sky130A
timestamp 1625669215
<< error_s >>
rect 6280 4601 6286 4607
rect 6333 4601 6339 4607
rect 6446 4601 6452 4607
rect 6499 4601 6505 4607
rect 6274 4551 6280 4557
rect 6339 4551 6345 4557
rect 6440 4551 6446 4557
rect 6505 4551 6511 4557
rect 5852 4542 5858 4548
rect 5957 4542 5963 4548
rect 6869 4542 6875 4548
rect 6974 4542 6980 4548
rect 5846 4492 5852 4498
rect 5963 4492 5969 4498
rect 6863 4492 6869 4498
rect 6980 4492 6986 4498
rect 5852 4241 5858 4247
rect 5957 4241 5963 4247
rect 6869 4241 6875 4247
rect 6974 4241 6980 4247
rect 5846 4191 5852 4197
rect 5963 4191 5969 4197
rect 6280 4187 6286 4193
rect 6333 4187 6339 4193
rect 6446 4187 6452 4193
rect 6499 4187 6505 4193
rect 6863 4191 6869 4197
rect 6980 4191 6986 4197
rect 6274 4137 6280 4143
rect 6339 4137 6345 4143
rect 6440 4137 6446 4143
rect 6505 4137 6511 4143
rect 3309 4086 3560 4099
rect 3956 4086 4133 4099
rect 6285 3856 6291 3862
rect 6338 3856 6344 3862
rect 6450 3856 6456 3862
rect 6503 3856 6509 3862
rect 6279 3806 6285 3812
rect 6344 3806 6350 3812
rect 6444 3806 6450 3812
rect 6509 3806 6515 3812
rect 5810 3797 5816 3803
rect 5915 3797 5921 3803
rect 6873 3797 6879 3803
rect 6978 3797 6984 3803
rect 5804 3747 5810 3753
rect 5921 3747 5927 3753
rect 6867 3747 6873 3753
rect 6984 3747 6990 3753
rect 6678 3612 6695 3613
rect 6678 3595 6695 3596
rect 6116 3578 6117 3591
rect 5810 3496 5816 3502
rect 5915 3496 5921 3502
rect 6873 3496 6879 3502
rect 6978 3496 6984 3502
rect 5804 3446 5810 3452
rect 5921 3446 5927 3452
rect 6285 3442 6291 3448
rect 6338 3442 6344 3448
rect 6450 3442 6456 3448
rect 6503 3442 6509 3448
rect 6867 3446 6873 3452
rect 6984 3446 6990 3452
rect 1649 3422 1666 3425
rect 6279 3392 6285 3398
rect 6344 3392 6350 3398
rect 6444 3392 6450 3398
rect 6509 3392 6515 3398
rect 5720 3092 5726 3098
rect 5825 3092 5831 3098
rect 6691 3092 6697 3098
rect 6796 3092 6802 3098
rect 6146 3082 6152 3088
rect 6199 3082 6205 3088
rect 6317 3082 6323 3088
rect 6370 3082 6376 3088
rect 5714 3028 5720 3034
rect 5831 3028 5837 3034
rect 6140 3032 6146 3038
rect 6205 3032 6211 3038
rect 6311 3032 6317 3038
rect 6376 3032 6382 3038
rect 6685 3028 6691 3034
rect 6802 3028 6808 3034
rect 5720 2975 5726 2981
rect 5825 2975 5831 2981
rect 6146 2973 6152 2979
rect 6199 2973 6205 2979
rect 6317 2973 6323 2979
rect 6370 2973 6376 2979
rect 6691 2975 6697 2981
rect 6796 2975 6802 2981
rect 6140 2923 6146 2929
rect 6205 2923 6211 2929
rect 6311 2923 6317 2929
rect 6376 2923 6382 2929
rect 5714 2911 5720 2917
rect 5831 2911 5837 2917
rect 6685 2911 6691 2917
rect 6802 2911 6808 2917
rect 5720 2790 5726 2796
rect 5825 2790 5831 2796
rect 6691 2790 6697 2796
rect 6796 2790 6802 2796
rect 6146 2784 6152 2790
rect 6199 2784 6205 2790
rect 6317 2784 6323 2790
rect 6370 2784 6376 2790
rect 6140 2734 6146 2740
rect 6205 2734 6211 2740
rect 6311 2734 6317 2740
rect 6376 2734 6382 2740
rect 5714 2726 5720 2732
rect 5831 2726 5837 2732
rect 6685 2726 6691 2732
rect 6802 2726 6808 2732
rect 5720 2674 5726 2680
rect 5825 2674 5831 2680
rect 6691 2674 6697 2680
rect 6796 2674 6802 2680
rect 6146 2667 6152 2673
rect 6199 2667 6205 2673
rect 6317 2667 6323 2673
rect 6370 2667 6376 2673
rect 6140 2617 6146 2623
rect 6205 2617 6211 2623
rect 6311 2617 6317 2623
rect 6376 2617 6382 2623
rect 5714 2610 5720 2616
rect 5831 2610 5837 2616
rect 6685 2610 6691 2616
rect 6802 2610 6808 2616
rect 5780 2289 5786 2295
rect 5885 2289 5891 2295
rect 6206 2279 6212 2285
rect 6259 2279 6265 2285
rect 5774 2225 5780 2231
rect 5891 2225 5897 2231
rect 6200 2229 6206 2235
rect 6265 2229 6271 2235
rect 5780 2172 5786 2178
rect 5885 2172 5891 2178
rect 6206 2170 6212 2176
rect 6259 2170 6265 2176
rect 6200 2120 6206 2126
rect 6265 2120 6271 2126
rect 5774 2108 5780 2114
rect 5891 2108 5897 2114
rect 5780 1987 5786 1993
rect 5885 1987 5891 1993
rect 6043 1982 6060 1986
rect 6206 1981 6212 1987
rect 6259 1981 6265 1987
rect 6200 1931 6206 1937
rect 6265 1931 6271 1937
rect 5774 1923 5780 1929
rect 5891 1923 5897 1929
rect 5780 1871 5786 1877
rect 5885 1871 5891 1877
rect 6206 1864 6212 1870
rect 6259 1864 6265 1870
rect 6200 1814 6206 1820
rect 6265 1814 6271 1820
rect 5774 1807 5780 1813
rect 5891 1807 5897 1813
rect 6181 1350 6210 1366
rect 6260 1350 6289 1366
rect 6339 1350 6368 1366
rect 6418 1350 6447 1366
rect 5321 1321 5327 1327
rect 5376 1321 5382 1327
rect 5791 1326 5797 1332
rect 5896 1326 5902 1332
rect 6728 1326 6734 1332
rect 7578 1326 7585 1332
rect 6181 1316 6182 1317
rect 6209 1316 6210 1317
rect 6260 1316 6261 1317
rect 6288 1316 6289 1317
rect 6339 1316 6340 1317
rect 6367 1316 6368 1317
rect 6418 1316 6419 1317
rect 6446 1316 6447 1317
rect 6131 1287 6149 1316
rect 6180 1315 6211 1316
rect 6259 1315 6290 1316
rect 6338 1315 6369 1316
rect 6417 1315 6448 1316
rect 6181 1308 6210 1315
rect 6260 1308 6289 1315
rect 6339 1308 6368 1315
rect 6418 1308 6447 1315
rect 6181 1294 6191 1308
rect 6438 1294 6447 1308
rect 6181 1288 6210 1294
rect 6260 1288 6289 1294
rect 6339 1288 6368 1294
rect 6418 1288 6447 1294
rect 6180 1287 6211 1288
rect 6259 1287 6290 1288
rect 6338 1287 6369 1288
rect 6417 1287 6448 1288
rect 6480 1287 6497 1316
rect 6181 1286 6182 1287
rect 6209 1286 6210 1287
rect 6260 1286 6261 1287
rect 6288 1286 6289 1287
rect 6339 1286 6340 1287
rect 6367 1286 6368 1287
rect 6418 1286 6419 1287
rect 6446 1286 6447 1287
rect 5315 1271 5321 1277
rect 5382 1271 5388 1277
rect 5785 1276 5791 1282
rect 5902 1276 5908 1282
rect 6181 1237 6210 1252
rect 6260 1237 6289 1252
rect 6339 1237 6368 1252
rect 6418 1237 6447 1252
rect 2006 1141 2008 1142
rect 6181 1070 6210 1086
rect 6260 1070 6289 1086
rect 6339 1070 6368 1086
rect 6418 1070 6447 1086
rect 7888 1067 7893 1068
rect 6181 1036 6182 1037
rect 6209 1036 6210 1037
rect 6260 1036 6261 1037
rect 6288 1036 6289 1037
rect 6339 1036 6340 1037
rect 6367 1036 6368 1037
rect 6418 1036 6419 1037
rect 6446 1036 6447 1037
rect 5791 1027 5797 1033
rect 5896 1027 5902 1033
rect 6131 1007 6149 1036
rect 6180 1035 6211 1036
rect 6259 1035 6290 1036
rect 6338 1035 6369 1036
rect 6417 1035 6448 1036
rect 6181 1028 6210 1035
rect 6260 1028 6289 1035
rect 6339 1028 6368 1035
rect 6418 1028 6447 1035
rect 6181 1014 6191 1028
rect 6438 1014 6447 1028
rect 6181 1008 6210 1014
rect 6260 1008 6289 1014
rect 6339 1008 6368 1014
rect 6418 1008 6447 1014
rect 6180 1007 6211 1008
rect 6259 1007 6290 1008
rect 6338 1007 6369 1008
rect 6417 1007 6448 1008
rect 6480 1007 6497 1036
rect 6181 1006 6182 1007
rect 6209 1006 6210 1007
rect 6260 1006 6261 1007
rect 6288 1006 6289 1007
rect 6339 1006 6340 1007
rect 6367 1006 6368 1007
rect 6418 1006 6419 1007
rect 6446 1006 6447 1007
rect 5322 988 5351 1006
rect 5785 977 5791 983
rect 5902 977 5908 983
rect 6181 957 6210 972
rect 6260 957 6289 972
rect 6339 957 6368 972
rect 6418 957 6447 972
rect 5322 956 5323 957
rect 5350 956 5351 957
rect 5272 927 5290 956
rect 5321 955 5352 956
rect 5322 946 5351 955
rect 5322 937 5332 946
rect 5341 937 5351 946
rect 5322 928 5351 937
rect 5321 927 5352 928
rect 5383 927 5401 956
rect 5322 926 5323 927
rect 5350 926 5351 927
rect 5791 926 5797 932
rect 5896 926 5902 932
rect 6181 915 6210 931
rect 6260 915 6289 931
rect 6339 915 6368 931
rect 6418 915 6447 931
rect 8180 900 8181 955
rect 5322 877 5351 895
rect 5785 876 5791 882
rect 5902 876 5908 882
rect 6181 881 6182 882
rect 6209 881 6210 882
rect 6260 881 6261 882
rect 6288 881 6289 882
rect 6339 881 6340 882
rect 6367 881 6368 882
rect 6418 881 6419 882
rect 6446 881 6447 882
rect 6131 852 6149 881
rect 6180 880 6211 881
rect 6259 880 6290 881
rect 6338 880 6369 881
rect 6417 880 6448 881
rect 6181 873 6210 880
rect 6260 873 6289 880
rect 6339 873 6368 880
rect 6418 873 6447 880
rect 6181 859 6191 873
rect 6438 859 6447 873
rect 6181 853 6210 859
rect 6260 853 6289 859
rect 6339 853 6368 859
rect 6418 853 6447 859
rect 6180 852 6211 853
rect 6259 852 6290 853
rect 6338 852 6369 853
rect 6417 852 6448 853
rect 6480 852 6497 881
rect 6722 860 6728 866
rect 7584 860 7590 866
rect 6181 851 6182 852
rect 6209 851 6210 852
rect 6260 851 6261 852
rect 6288 851 6289 852
rect 6339 851 6340 852
rect 6367 851 6368 852
rect 6418 851 6419 852
rect 6446 851 6447 852
rect 6181 802 6210 817
rect 6260 802 6289 817
rect 6339 802 6368 817
rect 6418 802 6447 817
use sky130_hilas_DAC5bit01  sky130_hilas_DAC5bit01_0
timestamp 1625056879
transform 1 0 943 0 1 252
box 382 524 2040 1121
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_0
timestamp 1608245216
transform 1 0 1261 0 1 1187
box 64 419 528 1018
use sky130_hilas_nFETLarge  sky130_hilas_nFETLarge_0
timestamp 1625426387
transform 1 0 1227 0 1 2063
box 64 420 501 1003
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_3
timestamp 1625405207
transform 1 0 3493 0 1 1717
box 1050 5 1614 610
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_3
timestamp 1624113741
transform 1 0 3478 0 1 1812
box -30 -102 850 522
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_2
timestamp 1625405207
transform 1 0 3436 0 1 2605
box 1050 5 1614 610
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_2
timestamp 1624113741
transform 1 0 3432 0 1 2608
box -30 -102 850 522
use sky130_hilas_swc4x2cell  sky130_hilas_swc4x2cell_0
timestamp 1625491916
transform 1 0 6259 0 1 2554
box -1004 -4 1009 601
use sky130_hilas_WTA4Stage01  sky130_hilas_WTA4Stage01_0
timestamp 1625404155
transform 1 0 6376 0 1 1790
box -1121 -43 296 562
use sky130_hilas_FGcharacterization01  sky130_hilas_FGcharacterization01_0
timestamp 1625074044
transform 1 0 6129 0 1 525
box -912 259 2083 864
use sky130_hilas_Trans2med  sky130_hilas_Trans2med_0
timestamp 1625425852
transform 1 0 1717 0 1 3456
box -380 -143 -27 452
use sky130_hilas_Trans4small  sky130_hilas_Trans4small_0
timestamp 1608234847
transform 1 0 1146 0 1 4305
box 191 -150 471 438
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_1
timestamp 1625405207
transform 1 0 3447 0 1 3343
box 1050 5 1614 610
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_1
timestamp 1624113741
transform 1 0 3409 0 1 3450
box -30 -102 850 522
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_0
timestamp 1625405207
transform 1 0 3424 0 1 4104
box 1050 5 1614 610
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_0
timestamp 1624113741
transform 1 0 3339 0 1 4188
box -30 -102 850 522
use sky130_hilas_TA2Cell_1FG_Strong  sky130_hilas_TA2Cell_1FG_Strong_0
timestamp 1625491312
transform 1 0 7861 0 1 3929
box -2617 140 193 745
use sky130_hilas_TA2Cell_1FG  sky130_hilas_TA2Cell_1FG_0
timestamp 1625491133
transform 1 0 7865 0 1 3184
box -2616 140 193 745
use sky130_hilas_Tgate4Single01  sky130_hilas_Tgate4Single01_0
timestamp 1608226321
transform 1 0 8789 0 1 3847
box -36 -141 440 464
<< end >>
