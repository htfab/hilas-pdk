magic
tech sky130A
timestamp 1634057804
<< nwell >>
rect 64 465 309 634
rect 64 464 175 465
<< nmos >>
rect 88 85 293 105
<< pmos >>
rect 90 531 291 551
<< ndiff >>
rect 88 128 293 132
rect 88 111 104 128
rect 278 111 293 128
rect 88 105 293 111
rect 88 79 293 85
rect 88 62 104 79
rect 278 62 293 79
rect 88 53 293 62
<< pdiff >>
rect 90 575 291 586
rect 90 558 102 575
rect 279 558 291 575
rect 90 551 291 558
rect 90 525 291 531
rect 90 508 102 525
rect 279 508 291 525
rect 90 503 291 508
<< ndiffc >>
rect 104 111 278 128
rect 104 62 278 79
<< pdiffc >>
rect 102 558 279 575
rect 102 508 279 525
<< psubdiff >>
rect 88 42 293 53
rect 88 40 142 42
rect 159 40 179 42
rect 196 40 214 42
rect 231 40 250 42
rect 267 40 293 42
rect 88 23 103 40
rect 279 23 293 40
rect 88 17 293 23
<< nsubdiff >>
rect 90 609 291 616
rect 90 592 102 609
rect 279 592 291 609
rect 90 586 291 592
<< psubdiffcont >>
rect 142 40 159 42
rect 179 40 196 42
rect 214 40 231 42
rect 250 40 267 42
rect 103 23 279 40
<< nsubdiffcont >>
rect 102 592 279 609
<< poly >>
rect 76 531 90 551
rect 291 531 320 551
rect 305 486 320 531
rect 76 478 320 486
rect 76 461 103 478
rect 276 461 320 478
rect 76 456 320 461
rect 75 168 316 173
rect 75 151 105 168
rect 279 151 316 168
rect 75 144 316 151
rect 301 105 316 144
rect 75 85 88 105
rect 293 85 316 105
<< polycont >>
rect 103 461 276 478
rect 105 151 279 168
<< locali >>
rect 94 609 291 611
rect 94 592 102 609
rect 279 592 291 609
rect 94 591 118 592
rect 135 591 183 592
rect 200 591 248 592
rect 265 591 291 592
rect 94 575 291 591
rect 94 558 102 575
rect 279 558 291 575
rect 94 555 150 558
rect 167 555 217 558
rect 234 555 291 558
rect 94 553 291 555
rect 245 525 289 528
rect 94 508 102 525
rect 279 508 289 525
rect 245 507 259 508
rect 276 507 289 508
rect 245 504 289 507
rect 95 478 135 481
rect 95 461 103 478
rect 276 461 284 478
rect 95 458 135 461
rect 97 151 105 168
rect 279 151 288 168
rect 248 149 288 151
rect 96 128 143 131
rect 96 111 104 128
rect 278 111 286 128
rect 96 110 107 111
rect 124 110 143 111
rect 96 108 143 110
rect 95 79 286 81
rect 95 62 104 79
rect 278 62 286 79
rect 95 61 125 62
rect 142 61 161 62
rect 178 61 197 62
rect 214 61 233 62
rect 250 61 286 62
rect 95 42 286 61
rect 95 40 106 42
rect 123 40 142 42
rect 95 23 103 40
rect 159 40 179 42
rect 196 40 214 42
rect 231 40 250 42
rect 267 40 286 42
rect 279 23 287 40
rect 95 20 279 23
<< viali >>
rect 118 592 135 608
rect 183 592 200 608
rect 248 592 265 608
rect 118 591 135 592
rect 183 591 200 592
rect 248 591 265 592
rect 150 558 167 572
rect 217 558 234 572
rect 150 555 167 558
rect 217 555 234 558
rect 259 508 276 524
rect 259 507 276 508
rect 108 461 125 478
rect 259 151 276 168
rect 107 111 124 128
rect 107 110 124 111
rect 125 62 142 78
rect 161 62 178 78
rect 197 62 214 78
rect 233 62 250 78
rect 125 61 142 62
rect 161 61 178 62
rect 197 61 214 62
rect 233 61 250 62
rect 106 40 123 42
rect 106 25 123 40
rect 142 25 159 42
rect 214 25 231 42
rect 250 25 267 42
<< metal1 >>
rect 111 644 272 646
rect 111 618 115 644
rect 141 618 179 644
rect 205 618 243 644
rect 269 618 272 644
rect 111 608 272 618
rect 111 591 118 608
rect 135 591 183 608
rect 200 591 248 608
rect 265 591 272 608
rect 111 588 272 591
rect 114 587 272 588
rect 114 572 288 587
rect 114 555 150 572
rect 167 555 217 572
rect 234 555 288 572
rect 114 552 288 555
rect 248 524 288 552
rect 248 507 259 524
rect 276 507 288 524
rect 98 478 138 482
rect 98 461 108 478
rect 125 461 138 478
rect 98 128 138 461
rect 248 168 288 507
rect 248 151 259 168
rect 276 151 288 168
rect 248 148 288 151
rect 98 110 107 128
rect 124 110 138 128
rect 98 81 138 110
rect 98 79 273 81
rect 101 78 273 79
rect 101 61 125 78
rect 142 61 161 78
rect 178 61 197 78
rect 214 61 233 78
rect 250 61 273 78
rect 101 47 273 61
rect 100 42 273 47
rect 100 40 106 42
rect 88 25 106 40
rect 123 34 142 42
rect 159 34 214 42
rect 231 34 250 42
rect 159 25 169 34
rect 88 23 117 25
rect 100 8 117 23
rect 143 8 169 25
rect 195 25 214 34
rect 247 25 250 34
rect 267 25 273 42
rect 195 8 221 25
rect 247 8 273 25
rect 100 4 273 8
<< via1 >>
rect 115 618 141 644
rect 179 618 205 644
rect 243 618 269 644
rect 117 25 123 34
rect 123 25 142 34
rect 142 25 143 34
rect 117 8 143 25
rect 169 8 195 34
rect 221 25 231 34
rect 231 25 247 34
rect 221 8 247 25
<< metal2 >>
rect 0 644 373 650
rect 0 618 115 644
rect 141 618 179 644
rect 205 618 243 644
rect 269 618 373 644
rect 0 612 373 618
rect 0 558 373 584
rect 0 494 373 520
rect 0 434 373 460
rect 0 380 373 406
rect 0 326 373 352
rect 0 274 373 300
rect 0 222 373 248
rect 0 170 373 196
rect 0 118 373 144
rect 0 66 373 92
rect 0 34 373 40
rect 0 8 117 34
rect 143 8 169 34
rect 195 8 221 34
rect 247 8 373 34
rect 0 0 373 8
<< labels >>
rlabel metal2 362 612 373 650 0 VPWR
port 1 nsew
rlabel metal2 0 612 10 650 0 VPWR
port 1 nsew
rlabel metal2 362 0 373 40 0 VGND
port 2 nsew
rlabel metal2 0 0 11 40 0 VGND
port 2 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
