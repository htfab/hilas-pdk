magic
tech sky130A
timestamp 1632256358
<< checkpaint >>
rect -630 -248 5202 2102
<< error_s >>
rect 484 1358 516 1364
rect 4056 1358 4088 1364
rect 484 1300 516 1308
rect 4056 1300 4088 1308
rect 525 1224 558 1227
rect 4014 1224 4047 1227
rect 484 1160 522 1189
rect 650 1073 692 1200
rect 728 1045 819 1073
rect 728 1039 845 1045
rect 867 1039 917 1045
rect 3655 1039 3705 1045
rect 3727 1039 3777 1045
rect 484 1038 516 1039
rect 728 1003 819 1039
rect 916 1003 946 1005
rect 1053 1004 1069 1018
rect 1094 1004 1113 1018
rect 1134 1005 1150 1019
rect 3422 1005 3438 1019
rect 3459 1004 3478 1018
rect 3503 1004 3519 1018
rect 728 997 845 1003
rect 867 999 946 1003
rect 3626 1003 3656 1005
rect 3626 999 3705 1003
rect 867 997 917 999
rect 3655 997 3705 999
rect 3727 997 3777 1003
rect 484 975 516 988
rect 728 982 819 997
rect 930 987 960 991
rect 3612 987 3642 991
rect 930 985 958 987
rect 3614 985 3642 987
rect 484 899 516 900
rect 650 855 692 982
rect 728 974 984 982
rect 728 956 989 974
rect 728 882 984 956
rect 1482 913 1593 941
rect 484 836 516 849
rect 728 777 819 855
rect 867 803 917 809
rect 967 781 984 842
rect 1449 824 1626 913
rect 1908 907 1967 947
rect 2017 916 2024 982
rect 2548 916 2555 982
rect 2605 916 2664 947
rect 1875 830 2000 907
rect 2017 898 2101 916
rect 2548 907 2664 916
rect 2979 913 3090 941
rect 2548 898 2697 907
rect 2572 830 2697 898
rect 2946 824 3123 913
rect 3588 882 3844 982
rect 867 761 917 767
rect 967 763 989 781
rect 930 750 958 752
rect 930 746 960 750
rect 916 732 946 738
rect 932 719 958 721
rect 768 711 788 719
rect 916 711 958 719
rect 967 715 984 763
rect 1011 715 1196 798
rect 1011 714 1111 715
rect 1112 714 1196 715
rect 3376 715 3561 798
rect 3376 714 3460 715
rect 3478 714 3561 715
rect 916 694 927 702
rect 932 692 958 711
rect 1088 709 1091 714
rect 1094 698 1196 714
rect 3435 710 3561 714
rect 3435 707 3448 710
rect 3443 703 3448 707
rect 3455 703 3561 710
rect 3443 698 3561 703
rect 3588 698 3605 842
rect 3655 803 3705 809
rect 3880 777 3922 1200
rect 4050 1160 4088 1189
rect 4056 1038 4088 1039
rect 4056 975 4088 988
rect 4056 899 4088 900
rect 4056 836 4088 849
rect 3655 761 3705 767
rect 3614 750 3642 752
rect 3612 746 3642 750
rect 3626 732 3656 738
rect 3614 719 3640 721
rect 3614 711 3656 719
rect 3784 711 3804 719
rect 1105 691 1108 695
rect 1121 693 1134 698
rect 3452 693 3465 698
rect 1121 690 1129 693
rect 3452 690 3460 693
rect 3478 691 3481 695
rect 3614 692 3640 711
rect 3645 694 3656 702
rect 916 675 946 681
rect 3626 675 3656 681
rect 930 663 960 667
rect 930 661 958 663
rect 728 650 984 659
rect 728 632 989 650
rect 728 558 984 632
rect 1343 586 1352 619
rect 1357 600 1376 614
rect 1397 600 1413 614
rect 1482 610 1593 617
rect 1482 596 1615 610
rect 1482 593 1593 596
rect 1809 595 1847 609
rect 1280 554 1294 572
rect 1316 571 1328 582
rect 1327 557 1328 568
rect 1280 511 1294 529
rect 1449 500 1626 593
rect 1908 587 1967 619
rect 1989 605 2008 613
rect 2212 592 2252 606
rect 2320 595 2360 609
rect 2564 605 2583 614
rect 1875 502 2000 587
rect 2252 578 2266 591
rect 2306 581 2320 591
rect 2605 587 2664 619
rect 2979 612 3090 617
rect 2725 595 2763 609
rect 2957 598 3090 612
rect 3159 600 3175 614
rect 3196 600 3215 614
rect 2979 593 3090 598
rect 2572 502 2697 587
rect 2946 500 3123 593
rect 3220 586 3229 619
rect 3264 617 3273 671
rect 3612 663 3642 667
rect 3614 661 3642 663
rect 3273 587 3348 617
rect 3244 571 3256 582
rect 3244 557 3245 568
rect 3283 554 3297 572
rect 3588 558 3844 659
rect 3283 511 3297 529
rect 1266 497 1301 499
rect 3269 497 3306 499
rect 867 480 917 486
rect 3655 480 3705 486
rect 867 438 917 444
rect 975 440 989 458
rect 930 427 958 429
rect 930 423 960 427
rect 1203 418 1293 453
rect 3588 440 3602 458
rect 3655 438 3705 444
rect 3614 427 3642 429
rect 3612 423 3642 427
rect 795 411 845 417
rect 867 415 917 417
rect 867 411 946 415
rect 916 409 946 411
rect 1203 400 1294 418
rect 3286 400 3300 418
rect 3655 415 3705 417
rect 3626 411 3705 415
rect 3727 411 3777 417
rect 3626 409 3656 411
rect 1203 375 1293 400
rect 795 369 845 375
rect 867 369 917 375
rect 1203 369 1364 375
rect 1280 357 1364 369
rect 3286 357 3300 375
rect 3655 369 3705 375
rect 3727 369 3777 375
rect 1280 230 1294 248
rect 3283 230 3297 248
rect 1280 187 1294 205
rect 3283 187 3297 205
rect 1280 77 1294 95
rect 3283 77 3297 95
rect 1280 34 1294 52
rect 3283 34 3297 52
rect 1316 0 1332 14
rect 1357 1 1376 15
rect 1397 1 1413 15
rect 1591 0 1615 14
rect 1809 0 1847 14
rect 1984 0 2008 14
rect 2212 0 2252 14
rect 2320 0 2360 14
rect 2564 0 2588 14
rect 2725 0 2763 15
rect 2957 0 2981 14
rect 3159 1 3175 15
rect 3196 1 3215 15
rect 3240 1 3256 15
<< nwell >>
rect 3264 587 3273 617
rect 1280 369 1293 375
rect 1280 357 1287 369
<< metal1 >>
rect 3241 615 3273 616
rect 1301 614 1332 615
rect 1301 601 1304 614
rect 1300 588 1304 601
rect 1330 588 1332 614
rect 3241 605 3244 615
rect 1357 600 1376 605
rect 1397 600 1413 605
rect 1591 596 1615 605
rect 1809 595 1847 605
rect 1984 599 2008 605
rect 2212 592 2252 605
rect 2320 595 2360 605
rect 2564 600 2588 605
rect 2725 595 2763 605
rect 2957 598 2981 605
rect 3159 600 3175 605
rect 3196 600 3215 605
rect 1300 586 1332 588
rect 1316 571 1332 586
rect 2252 569 2320 591
rect 3240 589 3244 605
rect 3270 589 3273 615
rect 3240 588 3273 589
rect 3240 571 3256 588
rect 1316 0 1332 6
rect 1357 1 1376 7
rect 1397 1 1413 7
rect 1591 0 1615 8
rect 1809 0 1847 9
rect 1984 0 2008 7
rect 2212 0 2252 12
rect 2320 0 2360 12
rect 2564 0 2588 7
rect 2725 0 2763 15
rect 2957 0 2981 6
rect 3159 1 3175 7
rect 3196 1 3215 7
rect 3240 1 3256 7
<< via1 >>
rect 1304 588 1330 614
rect 3244 589 3270 615
<< metal2 >>
rect 1300 615 3274 618
rect 1300 614 3244 615
rect 1300 588 1304 614
rect 1330 600 3244 614
rect 1330 588 1342 600
rect 1300 586 1342 588
rect 3240 589 3244 600
rect 3270 589 3274 615
rect 3240 587 3274 589
rect 1280 554 1286 572
rect 3283 554 3292 572
rect 1280 511 1287 529
rect 3283 511 3292 529
rect 1280 400 1286 418
rect 3286 400 3292 418
rect 1280 357 1293 375
rect 3286 357 3292 375
rect 1280 230 1287 248
rect 3283 230 3292 248
rect 1280 187 1287 205
rect 3283 187 3292 205
rect 1950 138 2626 156
rect 1280 77 1287 95
rect 3283 77 3292 95
rect 1280 34 1287 52
rect 3283 34 3292 52
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_1
timestamp 1632256337
transform -1 0 2024 0 1 382
box 0 0 2024 1090
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_0
timestamp 1632256337
transform 1 0 2548 0 1 382
box 0 0 2024 1090
<< labels >>
rlabel metal1 2725 595 2763 605 0 GATE2
port 1 nsew analog default
rlabel metal1 2212 0 2252 12 0 VTUN
port 2 nsew power default
rlabel metal1 2320 0 2360 12 0 VTUN
port 2 nsew power default
rlabel metal1 2320 595 2360 605 0 VTUN
port 2 nsew power default
rlabel metal1 2212 592 2252 605 0 VTUN
port 2 nsew power default
rlabel metal1 1809 595 1847 605 0 GATE1
port 3 nsew analog default
rlabel metal1 1809 0 1847 9 0 GATE1
port 3 nsew analog default
rlabel metal1 3240 1 3256 7 0 VINJ
port 4 nsew power default
rlabel metal1 2725 0 2763 15 0 GATE2
port 1 nsew analog default
rlabel metal1 3196 600 3215 605 0 SelectGate2
rlabel metal1 3240 600 3256 605 0 VINJ
port 6 nsew power default
rlabel metal1 1316 600 1332 605 0 VINJ
port 6 nsew power default
rlabel metal1 1357 600 1376 605 0 GATESELECT1
port 10 nsew analog default
rlabel metal1 1316 0 1332 6 0 VINJ
port 6 nsew power default
rlabel metal1 1357 1 1376 7 0 GATESELECT1
port 10 nsew analog default
rlabel metal1 1397 600 1413 605 0 COL1
port 12 nsew analog default
rlabel metal1 1397 1 1413 7 0 COL1
port 12 nsew analog default
rlabel metal1 3196 1 3215 7 0 GATESELECT2
port 11 nsew analog default
rlabel metal1 3159 1 3175 7 0 COL2
port 13 nsew analog default
rlabel metal1 3159 600 3175 605 0 COL2
port 13 nsew analog default
rlabel metal1 1591 599 1615 605 0 VGND
port 22 nsew
rlabel metal1 1591 0 1615 8 0 VGND
port 22 nsew
rlabel metal1 1984 0 2008 7 0 VGND
port 22 nsew
rlabel metal1 1984 599 2008 605 0 VGND
port 22 nsew
rlabel metal1 2564 0 2588 7 0 VGND
port 22 nsew
rlabel metal1 2957 0 2981 6 0 VGND
port 22 nsew
rlabel metal1 2564 600 2588 605 0 VGND
port 22 nsew
rlabel metal1 2957 598 2981 605 0 VGND
port 22 nsew
rlabel metal2 1280 34 1287 52 0 DRAIN4
port 21 nsew
rlabel metal2 1280 77 1287 95 0 ROW4
port 20 nsew
rlabel metal2 1280 187 1287 205 0 ROW3
port 19 nsew
rlabel metal2 1280 230 1287 248 0 DRAIN3
port 18 nsew
rlabel metal2 1280 357 1287 375 0 DRAIN2
port 17 nsew
rlabel metal2 1280 400 1286 418 0 ROW2
port 15 nsew
rlabel metal2 1280 511 1287 529 0 ROW1
port 14 nsew
rlabel metal2 1280 554 1286 572 0 DRAIN1
port 16 nsew
rlabel metal2 3283 511 3292 529 0 ROW1
port 14 nsew
rlabel metal2 3286 400 3292 418 0 ROW2
port 15 nsew
rlabel metal2 3286 357 3292 375 0 DRAIN2
port 17 nsew
rlabel metal2 3283 230 3292 248 0 DRAIN3
port 18 nsew
rlabel metal2 3283 187 3292 205 0 ROW3
port 19 nsew
rlabel metal2 3283 77 3292 95 0 ROW4
port 20 nsew
rlabel metal2 3283 34 3292 52 0 DRAIN4
port 21 nsew
rlabel metal2 3283 554 3292 572 0 DRAIN1
port 16 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
