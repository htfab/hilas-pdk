magic
tech sky130A
timestamp 1628707260
<< nwell >>
rect 0 0 173 190
<< mvvaractor >>
rect 57 67 116 117
<< mvnsubdiff >>
rect 57 117 116 153
rect 57 33 116 67
<< poly >>
rect 15 67 57 117
rect 116 67 158 117
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
