magic
tech sky130A
timestamp 1628285143
<< error_s >>
rect 35 554 85 560
rect 358 555 408 561
rect 515 554 543 561
rect 657 555 685 561
rect 35 512 85 518
rect 358 513 408 519
rect 515 512 543 519
rect 657 513 685 519
rect 106 488 156 494
rect 286 483 337 489
rect 466 483 494 489
rect 706 483 734 489
rect 106 446 156 452
rect 286 441 337 447
rect 466 441 494 447
rect 706 441 734 447
rect 35 379 85 385
rect 358 380 408 386
rect 515 379 543 386
rect 657 380 685 386
rect 35 337 85 343
rect 358 338 408 344
rect 515 337 543 344
rect 657 338 685 344
rect 106 313 156 319
rect 286 308 337 314
rect 466 308 494 314
rect 706 308 734 314
rect 106 271 156 277
rect 286 266 337 272
rect 466 266 494 272
rect 706 266 734 272
rect 35 204 85 210
rect 358 205 408 211
rect 515 204 543 211
rect 657 205 685 211
rect 35 162 85 168
rect 358 163 408 169
rect 515 162 543 169
rect 657 163 685 169
rect 106 138 156 144
rect 286 133 337 139
rect 466 133 494 139
rect 706 133 734 139
rect 106 96 156 102
rect 286 91 337 97
rect 466 91 494 97
rect 706 91 734 97
rect 35 29 85 35
rect 358 30 408 36
rect 515 29 543 36
rect 657 30 685 36
rect 35 -13 85 -7
rect 358 -12 408 -6
rect 515 -13 543 -6
rect 657 -12 685 -6
rect 106 -37 156 -31
rect 286 -42 337 -36
rect 466 -42 494 -36
rect 706 -42 734 -36
rect 106 -79 156 -73
rect 286 -84 337 -78
rect 466 -84 494 -78
rect 706 -84 734 -78
use sky130_hilas_StepUpDigital  StepUpDigital_2
timestamp 1628285143
transform 1 0 -49 0 1 463
box 19 -44 889 131
use sky130_hilas_StepUpDigital  StepUpDigital_1
timestamp 1628285143
transform 1 0 -49 0 1 288
box 19 -44 889 131
use sky130_hilas_StepUpDigital  StepUpDigital_3
timestamp 1628285143
transform 1 0 -49 0 1 -62
box 19 -44 889 131
use sky130_hilas_StepUpDigital  StepUpDigital_0
timestamp 1628285143
transform 1 0 -49 0 1 113
box 19 -44 889 131
<< labels >>
rlabel space 746 517 770 522 0 VPWR
port 5 nsew
rlabel metal1 746 -102 770 -97 0 VPWR
port 5 nsew
rlabel space 4 517 33 522 0 VINJ
port 6 nsew
rlabel metal1 4 -102 33 -97 0 VINJ
port 6 nsew
rlabel space -30 470 -19 490 0 OUTPUT1
port 7 nsew
rlabel space -30 315 -19 335 0 OUTPUT2
port 8 nsew
rlabel space -30 160 -19 180 0 OUTPUT3
port 9 nsew
rlabel metal2 -30 5 -19 25 0 OUTPUT4
port 10 nsew
rlabel space 445 515 476 522 0 VGND
port 11 nsew
rlabel metal1 445 -102 476 -96 0 VGND
port 11 nsew
<< end >>
