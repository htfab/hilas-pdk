magic
tech sky130A
timestamp 1627742263
<< nwell >>
rect -1451 -400 -1278 -210
<< mvvaractor >>
rect -1394 -333 -1335 -283
<< mvnsubdiff >>
rect -1394 -283 -1335 -247
rect -1394 -367 -1335 -333
<< poly >>
rect -1436 -333 -1394 -283
rect -1335 -333 -1293 -283
<< end >>
