magic
tech sky130A
timestamp 1637952898
<< error_p >>
rect -252 211 -199 218
rect -73 210 -21 218
rect -252 169 -199 176
rect -73 168 -21 176
<< nwell >>
rect -336 143 -138 308
<< mvnmos >>
rect -73 176 -21 210
<< mvpmos >>
rect -252 176 -199 211
<< mvndiff >>
rect -101 202 -73 210
rect -101 185 -96 202
rect -79 185 -73 202
rect -101 176 -73 185
rect -21 201 7 210
rect -21 184 -15 201
rect 2 184 7 201
rect -21 176 7 184
<< mvpdiff >>
rect -279 202 -252 211
rect -279 185 -275 202
rect -258 185 -252 202
rect -279 176 -252 185
rect -199 202 -171 211
rect -199 185 -193 202
rect -176 185 -171 202
rect -199 176 -171 185
<< mvndiffc >>
rect -96 185 -79 202
rect -15 184 2 201
<< mvpdiffc >>
rect -275 185 -258 202
rect -193 185 -176 202
<< psubdiff >>
rect -29 261 15 269
rect -29 244 -15 261
rect 2 244 15 261
rect -29 237 15 244
<< mvnsubdiff >>
rect -286 267 -245 275
rect -286 250 -274 267
rect -257 250 -245 267
rect -286 241 -245 250
<< psubdiffcont >>
rect -15 244 2 261
<< mvnsubdiffcont >>
rect -274 250 -257 267
<< poly >>
rect -325 224 -36 235
rect -325 219 -21 224
rect -325 203 -296 219
rect -252 211 -199 219
rect -325 186 -320 203
rect -303 186 -296 203
rect -325 174 -296 186
rect -73 210 -21 219
rect -252 163 -199 176
rect -73 163 -21 176
<< polycont >>
rect -320 186 -303 203
<< locali >>
rect -274 267 -257 279
rect -274 248 -272 250
rect -15 261 2 269
rect -274 238 -257 248
rect -15 229 2 244
rect -323 203 -300 218
rect -323 202 -320 203
rect -323 184 -321 202
rect -303 186 -300 203
rect -304 184 -300 186
rect -323 176 -300 184
rect -275 204 -258 210
rect -275 202 -250 204
rect -258 197 -250 202
rect -275 180 -271 185
rect -254 180 -250 197
rect -201 202 -176 210
rect -201 185 -193 202
rect -176 185 -137 202
rect -120 185 -96 202
rect -79 185 -71 202
rect -15 201 2 212
rect -275 177 -250 180
rect -274 175 -250 177
rect -193 176 -176 185
rect -23 184 -15 201
rect 2 184 10 201
<< viali >>
rect -272 250 -257 265
rect -257 250 -255 265
rect -272 248 -255 250
rect -15 212 2 229
rect -321 186 -320 202
rect -320 186 -304 202
rect -321 184 -304 186
rect -271 185 -258 197
rect -258 185 -254 197
rect -271 180 -254 185
rect -137 185 -120 202
<< metal1 >>
rect -275 270 -253 304
rect -275 265 -252 270
rect -275 248 -272 265
rect -255 248 -252 265
rect -275 244 -252 248
rect -325 208 -299 210
rect -326 207 -298 208
rect -326 181 -325 207
rect -299 181 -298 207
rect -326 177 -298 181
rect -275 204 -253 244
rect -18 229 5 304
rect -18 212 -15 229
rect 2 212 5 229
rect -275 197 -250 204
rect -275 180 -271 197
rect -254 180 -250 197
rect -145 180 -142 206
rect -116 180 -113 206
rect -275 173 -250 180
rect -275 153 -253 173
rect -18 153 5 212
<< via1 >>
rect -325 202 -299 207
rect -325 184 -321 202
rect -321 184 -304 202
rect -304 184 -299 202
rect -325 181 -299 184
rect -142 202 -116 206
rect -142 185 -137 202
rect -137 185 -120 202
rect -120 185 -116 202
rect -142 180 -116 185
<< metal2 >>
rect -336 247 25 265
rect -320 210 -299 247
rect -325 207 -299 210
rect -325 178 -299 181
rect -145 180 -142 206
rect -116 198 -113 206
rect -116 180 25 198
<< labels >>
rlabel metal1 -275 153 -253 159 0 Vinj
rlabel metal1 -275 297 -253 304 0 Vinj
rlabel metal1 -18 295 5 304 0 GND
rlabel metal1 -18 153 5 159 0 GND
rlabel metal2 -336 247 -326 265 0 Input
rlabel metal2 16 247 25 265 0 Input
rlabel metal2 16 180 25 198 0 Output
<< end >>
