magic
tech sky130A
timestamp 1632251375
<< error_p >>
rect 132 136 182 142
rect 289 135 317 142
rect 431 136 459 142
rect 132 94 182 100
rect 289 93 317 100
rect 431 94 459 100
rect 60 64 111 70
rect 240 64 268 70
rect 480 64 508 70
rect 60 22 111 28
rect 240 22 268 28
rect 480 22 508 28
<< nwell >>
rect 381 9 558 168
<< nmos >>
rect 289 100 317 135
rect 240 28 268 64
<< pmos >>
rect 431 100 459 136
rect 480 28 508 64
<< mvnmos >>
rect 132 100 182 136
rect 60 28 111 64
<< ndiff >>
rect 255 121 289 135
rect 255 104 266 121
rect 283 104 289 121
rect 255 100 289 104
rect 317 121 346 135
rect 317 104 323 121
rect 340 104 346 121
rect 317 100 346 104
rect 211 59 240 64
rect 211 42 217 59
rect 234 42 240 59
rect 211 28 240 42
rect 268 59 297 64
rect 268 42 274 59
rect 291 42 297 59
rect 268 28 297 42
<< pdiff >>
rect 400 121 431 136
rect 400 104 406 121
rect 424 104 431 121
rect 400 100 431 104
rect 459 121 495 136
rect 459 104 465 121
rect 482 104 495 121
rect 459 100 495 104
rect 451 59 480 64
rect 451 42 457 59
rect 474 42 480 59
rect 451 28 480 42
rect 508 59 539 64
rect 508 42 515 59
rect 532 42 539 59
rect 508 28 539 42
<< mvndiff >>
rect 104 124 132 136
rect 104 107 108 124
rect 126 107 132 124
rect 104 100 132 107
rect 182 124 213 136
rect 182 107 188 124
rect 206 107 213 124
rect 182 100 213 107
rect 28 56 60 64
rect 28 39 35 56
rect 53 39 60 56
rect 28 28 60 39
rect 111 54 142 64
rect 111 37 117 54
rect 135 37 142 54
rect 111 28 142 37
<< ndiffc >>
rect 266 104 283 121
rect 323 104 340 121
rect 217 42 234 59
rect 274 42 291 59
<< pdiffc >>
rect 406 104 424 121
rect 465 104 482 121
rect 457 42 474 59
rect 515 42 532 59
<< mvndiffc >>
rect 108 107 126 124
rect 188 107 206 124
rect 35 39 53 56
rect 117 37 135 54
<< psubdiff >>
rect 213 121 255 135
rect 213 104 225 121
rect 242 104 255 121
rect 213 100 255 104
<< nsubdiff >>
rect 495 121 540 136
rect 495 104 507 121
rect 524 104 540 121
rect 495 100 540 104
<< psubdiffcont >>
rect 225 104 242 121
<< nsubdiffcont >>
rect 507 104 524 121
<< poly >>
rect 167 158 236 159
rect 132 144 317 158
rect 132 136 182 144
rect 221 143 317 144
rect 289 135 317 143
rect 431 136 459 149
rect 132 86 182 100
rect 289 91 317 100
rect 431 91 459 100
rect 60 64 111 78
rect 240 64 268 82
rect 289 76 459 91
rect 156 48 183 63
rect 156 31 161 48
rect 178 31 183 48
rect 60 20 111 28
rect 156 20 183 31
rect 356 59 364 76
rect 381 59 389 76
rect 480 64 508 80
rect 356 58 389 59
rect 359 54 386 58
rect 565 43 603 53
rect 60 5 183 20
rect 240 20 268 28
rect 480 20 508 28
rect 565 26 575 43
rect 592 26 603 43
rect 565 20 603 26
rect 240 15 603 20
rect 240 5 593 15
<< polycont >>
rect 161 31 178 48
rect 364 59 381 76
rect 575 26 592 43
<< locali >>
rect 16 126 33 130
rect 357 129 392 131
rect 16 124 131 126
rect 16 107 108 124
rect 126 107 135 124
rect 180 107 188 124
rect 206 121 226 124
rect 357 121 363 129
rect 206 107 225 121
rect 209 104 225 107
rect 242 104 266 121
rect 283 104 291 121
rect 315 104 323 121
rect 340 108 363 121
rect 384 121 392 129
rect 384 108 406 121
rect 340 104 406 108
rect 424 104 432 121
rect 457 104 465 121
rect 482 104 507 121
rect 524 104 533 121
rect 209 90 235 104
rect 117 73 235 90
rect 510 103 533 104
rect 510 88 537 103
rect 0 39 35 56
rect 53 39 62 56
rect 117 54 135 73
rect 209 59 235 73
rect 356 76 389 85
rect 356 59 364 76
rect 381 59 389 76
rect 510 71 514 88
rect 531 71 537 88
rect 510 59 537 71
rect 117 29 135 37
rect 159 48 180 56
rect 159 31 161 48
rect 178 31 180 48
rect 209 42 217 59
rect 234 42 242 59
rect 266 42 274 59
rect 291 42 457 59
rect 474 42 482 59
rect 507 42 515 59
rect 532 42 540 59
rect 575 45 592 51
rect 209 37 226 42
rect 507 41 540 42
rect 159 23 180 31
rect 575 18 592 23
<< viali >>
rect 363 108 384 129
rect 514 71 531 88
rect 573 43 595 45
rect 573 26 575 43
rect 575 26 592 43
rect 592 26 595 43
rect 573 23 595 26
<< metal1 >>
rect 156 59 184 62
rect 156 33 157 59
rect 183 33 184 59
rect 156 29 184 33
rect 209 0 240 169
rect 357 131 392 133
rect 357 105 361 131
rect 387 105 392 131
rect 357 104 392 105
rect 372 102 392 104
rect 510 88 534 168
rect 510 71 514 88
rect 531 71 534 88
rect 510 0 534 71
rect 567 47 608 51
rect 567 21 571 47
rect 597 21 608 47
rect 567 18 608 21
<< via1 >>
rect 157 33 183 59
rect 361 129 387 131
rect 361 108 363 129
rect 363 108 384 129
rect 384 108 387 129
rect 361 105 387 108
rect 571 45 597 47
rect 571 23 573 45
rect 573 23 595 45
rect 595 23 597 45
rect 571 21 597 23
<< metal2 >>
rect 361 131 387 134
rect 153 59 187 60
rect 153 33 157 59
rect 183 54 187 59
rect 361 54 387 105
rect 183 33 397 54
rect 153 32 397 33
rect 568 47 614 50
rect 568 21 571 47
rect 597 21 614 47
rect 568 18 614 21
<< labels >>
rlabel metal2 607 18 614 50 0 Input
rlabel metal1 510 164 534 168 0 Vdd
rlabel metal1 510 9 534 13 0 Vdd
rlabel metal1 209 164 240 168 0 GND
rlabel metal1 209 9 240 14 0 GND
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
