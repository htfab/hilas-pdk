magic
tech sky130A
timestamp 1629421669
<< error_s >>
rect -626 12757 -597 12773
rect -547 12757 -518 12773
rect -468 12757 -439 12773
rect -389 12757 -360 12773
rect -626 12723 -625 12724
rect -598 12723 -597 12724
rect -547 12723 -546 12724
rect -519 12723 -518 12724
rect -468 12723 -467 12724
rect -440 12723 -439 12724
rect -389 12723 -388 12724
rect -361 12723 -360 12724
rect -676 12694 -659 12723
rect -627 12722 -596 12723
rect -548 12722 -517 12723
rect -469 12722 -438 12723
rect -390 12722 -359 12723
rect -626 12715 -597 12722
rect -547 12715 -518 12722
rect -468 12715 -439 12722
rect -389 12715 -360 12722
rect -626 12701 -617 12715
rect -370 12701 -360 12715
rect -626 12695 -597 12701
rect -547 12695 -518 12701
rect -468 12695 -439 12701
rect -389 12695 -360 12701
rect -627 12694 -596 12695
rect -548 12694 -517 12695
rect -469 12694 -438 12695
rect -390 12694 -359 12695
rect -328 12694 -310 12723
rect -626 12693 -625 12694
rect -598 12693 -597 12694
rect -547 12693 -546 12694
rect -519 12693 -518 12694
rect -468 12693 -467 12694
rect -440 12693 -439 12694
rect -389 12693 -388 12694
rect -361 12693 -360 12694
rect -626 12644 -597 12659
rect -547 12644 -518 12659
rect -468 12644 -439 12659
rect -389 12644 -360 12659
rect -626 12477 -597 12493
rect -547 12477 -518 12493
rect -468 12477 -439 12493
rect -389 12477 -360 12493
rect -626 12443 -625 12444
rect -598 12443 -597 12444
rect -547 12443 -546 12444
rect -519 12443 -518 12444
rect -468 12443 -467 12444
rect -440 12443 -439 12444
rect -389 12443 -388 12444
rect -361 12443 -360 12444
rect -676 12414 -659 12443
rect -627 12442 -596 12443
rect -548 12442 -517 12443
rect -469 12442 -438 12443
rect -390 12442 -359 12443
rect -626 12435 -597 12442
rect -547 12435 -518 12442
rect -468 12435 -439 12442
rect -389 12435 -360 12442
rect -626 12421 -617 12435
rect -370 12421 -360 12435
rect -626 12415 -597 12421
rect -547 12415 -518 12421
rect -468 12415 -439 12421
rect -389 12415 -360 12421
rect -627 12414 -596 12415
rect -548 12414 -517 12415
rect -469 12414 -438 12415
rect -390 12414 -359 12415
rect -328 12414 -310 12443
rect -626 12413 -625 12414
rect -598 12413 -597 12414
rect -547 12413 -546 12414
rect -519 12413 -518 12414
rect -468 12413 -467 12414
rect -440 12413 -439 12414
rect -389 12413 -388 12414
rect -361 12413 -360 12414
rect 470 12395 499 12413
rect -626 12364 -597 12379
rect -547 12364 -518 12379
rect -468 12364 -439 12379
rect -389 12364 -360 12379
rect 470 12363 471 12364
rect 498 12363 499 12364
rect -626 12322 -597 12338
rect -547 12322 -518 12338
rect -468 12322 -439 12338
rect -389 12322 -360 12338
rect 420 12334 438 12363
rect 469 12362 500 12363
rect 470 12353 499 12362
rect 470 12344 480 12353
rect 489 12344 499 12353
rect 470 12335 499 12344
rect 469 12334 500 12335
rect 531 12334 549 12363
rect 470 12333 471 12334
rect 498 12333 499 12334
rect -626 12288 -625 12289
rect -598 12288 -597 12289
rect -547 12288 -546 12289
rect -519 12288 -518 12289
rect -468 12288 -467 12289
rect -440 12288 -439 12289
rect -389 12288 -388 12289
rect -361 12288 -360 12289
rect -676 12259 -659 12288
rect -627 12287 -596 12288
rect -548 12287 -517 12288
rect -469 12287 -438 12288
rect -390 12287 -359 12288
rect -626 12280 -597 12287
rect -547 12280 -518 12287
rect -468 12280 -439 12287
rect -389 12280 -360 12287
rect -626 12266 -617 12280
rect -370 12266 -360 12280
rect -626 12260 -597 12266
rect -547 12260 -518 12266
rect -468 12260 -439 12266
rect -389 12260 -360 12266
rect -627 12259 -596 12260
rect -548 12259 -517 12260
rect -469 12259 -438 12260
rect -390 12259 -359 12260
rect -328 12259 -310 12288
rect 470 12284 499 12302
rect -626 12258 -625 12259
rect -598 12258 -597 12259
rect -547 12258 -546 12259
rect -519 12258 -518 12259
rect -468 12258 -467 12259
rect -440 12258 -439 12259
rect -389 12258 -388 12259
rect -361 12258 -360 12259
rect -626 12209 -597 12224
rect -547 12209 -518 12224
rect -468 12209 -439 12224
rect -389 12209 -360 12224
rect 1252 11655 1280 11661
rect 1394 11654 1422 11661
rect 1529 11655 1579 11661
rect 1852 11654 1902 11660
rect 1252 11613 1280 11619
rect 1394 11612 1422 11619
rect 1529 11613 1579 11619
rect 1852 11612 1902 11618
rect 1203 11583 1231 11589
rect 1443 11583 1471 11589
rect 1600 11583 1651 11589
rect 1781 11588 1831 11594
rect 1203 11541 1231 11547
rect 1443 11541 1471 11547
rect 1600 11541 1651 11547
rect 1781 11546 1831 11552
rect 1252 11480 1280 11486
rect 1394 11479 1422 11486
rect 1529 11480 1579 11486
rect 1852 11479 1902 11485
rect 1252 11438 1280 11444
rect 1394 11437 1422 11444
rect 1529 11438 1579 11444
rect 1852 11437 1902 11443
rect 1203 11408 1231 11414
rect 1443 11408 1471 11414
rect 1600 11408 1651 11414
rect 1781 11413 1831 11419
rect 1203 11366 1231 11372
rect 1443 11366 1471 11372
rect 1600 11366 1651 11372
rect 1781 11371 1831 11377
rect 1252 11305 1280 11311
rect 1394 11304 1422 11311
rect 1529 11305 1579 11311
rect 4595 11310 4680 11388
rect 1852 11304 1902 11310
rect 4595 11305 4596 11310
rect 2696 11277 2746 11283
rect 2768 11277 2818 11283
rect 4737 11277 4787 11283
rect 4809 11277 4859 11283
rect 5197 11281 5224 11287
rect 1252 11263 1280 11269
rect 1394 11262 1422 11269
rect 1529 11263 1579 11269
rect 1852 11262 1902 11268
rect 1203 11233 1231 11239
rect 1443 11233 1471 11239
rect 1600 11233 1651 11239
rect 1781 11238 1831 11244
rect 2696 11235 2746 11241
rect 2768 11235 2818 11241
rect 4737 11235 4787 11241
rect 4809 11235 4859 11241
rect 5197 11239 5224 11245
rect 5197 11214 5224 11220
rect 1203 11191 1231 11197
rect 1443 11191 1471 11197
rect 1600 11191 1651 11197
rect 1781 11196 1831 11202
rect 1252 11130 1280 11136
rect 1394 11129 1422 11136
rect 1529 11130 1579 11136
rect 1852 11129 1902 11135
rect 2881 11133 2884 11183
rect 2923 11133 2926 11183
rect 3017 11133 3019 11183
rect 3059 11133 3061 11183
rect 5197 11172 5224 11178
rect 5197 11131 5224 11137
rect 1252 11088 1280 11094
rect 1394 11087 1422 11094
rect 1529 11088 1579 11094
rect 1852 11087 1902 11093
rect 1203 11058 1231 11064
rect 1443 11058 1471 11064
rect 1600 11058 1651 11064
rect 1781 11063 1831 11069
rect 2881 11054 2884 11104
rect 2923 11054 2926 11104
rect 3017 11054 3019 11104
rect 3059 11054 3061 11104
rect 5197 11089 5224 11095
rect 5197 11064 5224 11070
rect 1203 11016 1231 11022
rect 1443 11016 1471 11022
rect 1600 11016 1651 11022
rect 1781 11021 1831 11027
rect 5197 11022 5224 11028
rect 7955 11024 7995 11030
rect 8105 11024 8145 11030
rect 5197 10981 5224 10987
rect 7955 10982 7995 10988
rect 8105 10982 8145 10988
rect 2106 10964 2156 10969
rect 2286 10964 2336 10970
rect 2426 10964 2476 10969
rect 1203 10955 1231 10961
rect 1443 10955 1471 10961
rect 1600 10955 1651 10961
rect 7879 10958 7919 10963
rect 8105 10956 8145 10963
rect 1781 10950 1831 10956
rect 2106 10922 2156 10927
rect 2286 10922 2336 10928
rect 2426 10922 2476 10927
rect 1203 10913 1231 10919
rect 1443 10913 1471 10919
rect 1600 10913 1651 10919
rect 1781 10908 1831 10914
rect 2106 10897 2156 10903
rect 2426 10897 2476 10903
rect 2881 10901 2884 10951
rect 2923 10901 2926 10951
rect 3017 10901 3019 10951
rect 3059 10901 3061 10951
rect 5197 10939 5224 10945
rect 5197 10914 5224 10920
rect 7879 10916 7919 10921
rect 8105 10914 8145 10921
rect 1252 10883 1280 10889
rect 1394 10883 1422 10890
rect 1529 10883 1579 10889
rect 1852 10884 1902 10890
rect 5197 10872 5224 10878
rect 2106 10855 2156 10861
rect 2426 10855 2476 10861
rect 1252 10841 1280 10847
rect 1394 10841 1422 10848
rect 1529 10841 1579 10847
rect 1852 10842 1902 10848
rect 2881 10822 2884 10872
rect 2923 10822 2926 10872
rect 3017 10822 3019 10872
rect 3059 10822 3061 10872
rect 7879 10854 7919 10859
rect 8105 10854 8145 10861
rect 5197 10831 5224 10837
rect 7879 10812 7919 10817
rect 8105 10812 8145 10819
rect 2106 10794 2156 10800
rect 2426 10794 2476 10800
rect 5197 10789 5224 10795
rect 7955 10787 7995 10793
rect 8105 10787 8145 10793
rect 1203 10780 1231 10786
rect 1443 10780 1471 10786
rect 1600 10780 1651 10786
rect 1781 10775 1831 10781
rect 2696 10764 2746 10770
rect 2768 10764 2818 10770
rect 2106 10752 2156 10758
rect 2426 10752 2476 10758
rect 1203 10738 1231 10744
rect 1443 10738 1471 10744
rect 1600 10738 1651 10744
rect 1781 10733 1831 10739
rect 2106 10728 2156 10733
rect 2286 10727 2336 10733
rect 2426 10728 2476 10733
rect 2696 10722 2746 10728
rect 2768 10722 2818 10728
rect 1252 10708 1280 10714
rect 1394 10708 1422 10715
rect 1529 10708 1579 10714
rect 1852 10709 1902 10715
rect 4595 10702 4596 10785
rect 4737 10764 4787 10770
rect 4809 10764 4859 10770
rect 5197 10764 5224 10770
rect 7955 10745 7995 10751
rect 8105 10745 8145 10751
rect 4737 10722 4787 10728
rect 4809 10722 4859 10728
rect 5197 10722 5224 10728
rect 7955 10704 7995 10710
rect 8105 10704 8145 10710
rect 2106 10686 2156 10691
rect 2286 10685 2336 10691
rect 2426 10686 2476 10691
rect 2697 10674 2747 10680
rect 2769 10674 2819 10680
rect 4737 10674 4787 10680
rect 4809 10674 4859 10680
rect 5197 10678 5224 10684
rect 1252 10666 1280 10672
rect 1394 10666 1422 10673
rect 1529 10666 1579 10672
rect 1852 10667 1902 10673
rect 7955 10662 7995 10668
rect 8105 10662 8145 10668
rect 2106 10644 2156 10649
rect 2286 10644 2336 10650
rect 2426 10644 2476 10649
rect 2697 10632 2747 10638
rect 2769 10632 2819 10638
rect 4737 10632 4787 10638
rect 4809 10632 4859 10638
rect 5197 10636 5224 10642
rect 7879 10638 7919 10643
rect 8105 10636 8145 10643
rect 5197 10611 5224 10617
rect 1203 10605 1231 10611
rect 1443 10605 1471 10611
rect 1600 10605 1651 10611
rect 1781 10600 1831 10606
rect 2106 10602 2156 10607
rect 2286 10602 2336 10608
rect 2426 10602 2476 10607
rect 7879 10596 7919 10601
rect 8105 10594 8145 10601
rect 2106 10577 2156 10583
rect 2426 10577 2476 10583
rect 5197 10569 5224 10575
rect 1203 10563 1231 10569
rect 1443 10563 1471 10569
rect 1600 10563 1651 10569
rect 1781 10558 1831 10564
rect 1252 10533 1280 10539
rect 1394 10533 1422 10540
rect 1529 10533 1579 10539
rect 1852 10534 1902 10540
rect 2106 10535 2156 10541
rect 2426 10535 2476 10541
rect 7879 10534 7919 10539
rect 8105 10534 8145 10541
rect 5197 10528 5224 10534
rect 1252 10491 1280 10497
rect 1394 10491 1422 10498
rect 1529 10491 1579 10497
rect 1852 10492 1902 10498
rect 7879 10492 7919 10497
rect 8105 10492 8145 10499
rect 5197 10486 5224 10492
rect 2106 10474 2156 10480
rect 2426 10474 2476 10480
rect 7955 10467 7995 10473
rect 8105 10467 8145 10473
rect 5197 10461 5224 10467
rect 1203 10430 1231 10436
rect 1443 10430 1471 10436
rect 1600 10430 1651 10436
rect 2106 10432 2156 10438
rect 2426 10432 2476 10438
rect 1781 10425 1831 10431
rect 7955 10425 7995 10431
rect 8105 10425 8145 10431
rect 5197 10419 5224 10425
rect 2106 10408 2156 10413
rect 2286 10407 2336 10413
rect 2426 10408 2476 10413
rect 1203 10388 1231 10394
rect 1443 10388 1471 10394
rect 1600 10388 1651 10394
rect 1781 10383 1831 10389
rect 5197 10378 5224 10384
rect 2106 10366 2156 10371
rect 2286 10365 2336 10371
rect 2426 10366 2476 10371
rect 1252 10358 1280 10364
rect 1394 10358 1422 10365
rect 1529 10358 1579 10364
rect 1852 10359 1902 10365
rect 5197 10336 5224 10342
rect 1252 10316 1280 10322
rect 1394 10316 1422 10323
rect 1529 10316 1579 10322
rect 1852 10317 1902 10323
rect 5197 10311 5224 10317
rect 5197 10269 5224 10275
rect 5197 10228 5224 10234
rect 5197 10186 5224 10192
rect 2697 10161 2747 10167
rect 2769 10161 2819 10167
rect 4737 10161 4787 10167
rect 4809 10161 4859 10167
rect 5197 10161 5224 10167
rect 2697 10119 2747 10125
rect 2769 10119 2819 10125
rect 4737 10119 4787 10125
rect 4809 10119 4859 10125
rect 5197 10119 5224 10125
rect 1203 9942 1231 9948
rect 1443 9942 1471 9948
rect 1600 9942 1651 9948
rect 1781 9937 1831 9943
rect 2104 9917 2154 9922
rect 2284 9917 2334 9923
rect 2424 9917 2474 9922
rect 2838 9916 2888 9922
rect 2910 9916 2960 9922
rect 4594 9916 4644 9922
rect 4666 9916 4716 9922
rect 1203 9900 1231 9906
rect 1443 9900 1471 9906
rect 1600 9900 1651 9906
rect 1781 9895 1831 9901
rect 1252 9870 1280 9876
rect 1394 9870 1422 9877
rect 1529 9870 1579 9876
rect 1852 9871 1902 9877
rect 2104 9875 2154 9880
rect 2284 9875 2334 9881
rect 2424 9875 2474 9880
rect 2838 9874 2888 9880
rect 2910 9874 2960 9880
rect 4594 9874 4644 9880
rect 4666 9874 4716 9880
rect 2104 9850 2154 9856
rect 2424 9850 2474 9856
rect 2910 9847 2960 9853
rect 4594 9847 4644 9853
rect 1252 9828 1280 9834
rect 1394 9828 1422 9835
rect 1529 9828 1579 9834
rect 1852 9829 1902 9835
rect 2104 9808 2154 9814
rect 2424 9808 2474 9814
rect 2910 9805 2960 9811
rect 4594 9805 4644 9811
rect 1203 9767 1231 9773
rect 1443 9767 1471 9773
rect 1600 9767 1651 9773
rect 1781 9762 1831 9768
rect 2910 9762 2960 9768
rect 4594 9762 4644 9768
rect 2104 9747 2154 9753
rect 2424 9747 2474 9753
rect 1203 9725 1231 9731
rect 1443 9725 1471 9731
rect 1600 9725 1651 9731
rect 1781 9720 1831 9726
rect 2910 9720 2960 9726
rect 4594 9720 4644 9726
rect 2104 9705 2154 9711
rect 2424 9705 2474 9711
rect 1252 9695 1280 9701
rect 1394 9695 1422 9702
rect 1529 9695 1579 9701
rect 1852 9696 1902 9702
rect 2838 9693 2888 9699
rect 2910 9693 2960 9699
rect 4594 9693 4644 9699
rect 4666 9693 4716 9699
rect 2104 9681 2154 9686
rect 2284 9680 2334 9686
rect 2424 9681 2474 9686
rect 1252 9653 1280 9659
rect 1394 9653 1422 9660
rect 1529 9653 1579 9659
rect 1852 9654 1902 9660
rect 2838 9651 2888 9657
rect 2910 9651 2960 9657
rect 4594 9651 4644 9657
rect 4666 9651 4716 9657
rect 2104 9639 2154 9644
rect 2284 9638 2334 9644
rect 2424 9639 2474 9644
rect 1203 9592 1231 9598
rect 1443 9592 1471 9598
rect 1600 9592 1651 9598
rect 2104 9597 2154 9602
rect 2284 9597 2334 9603
rect 2424 9597 2474 9602
rect 1781 9587 1831 9593
rect 2838 9592 2888 9598
rect 2910 9592 2960 9598
rect 4594 9592 4644 9598
rect 4666 9592 4716 9598
rect 1203 9550 1231 9556
rect 1443 9550 1471 9556
rect 1600 9550 1651 9556
rect 2104 9555 2154 9560
rect 2284 9555 2334 9561
rect 2424 9555 2474 9560
rect 1781 9545 1831 9551
rect 2838 9550 2888 9556
rect 2910 9550 2960 9556
rect 4594 9550 4644 9556
rect 4666 9550 4716 9556
rect 2104 9530 2154 9536
rect 2424 9530 2474 9536
rect 1252 9520 1280 9526
rect 1394 9520 1422 9527
rect 1529 9520 1579 9526
rect 1852 9521 1902 9527
rect 2910 9523 2960 9529
rect 4594 9523 4644 9529
rect 2104 9488 2154 9494
rect 2424 9488 2474 9494
rect 1252 9478 1280 9484
rect 1394 9478 1422 9485
rect 1529 9478 1579 9484
rect 1852 9479 1902 9485
rect 2910 9481 2960 9487
rect 4594 9481 4644 9487
rect 2910 9439 2960 9445
rect 4594 9439 4644 9445
rect 2104 9427 2154 9433
rect 2424 9427 2474 9433
rect 1203 9417 1231 9423
rect 1443 9417 1471 9423
rect 1600 9417 1651 9423
rect 1781 9412 1831 9418
rect 2910 9397 2960 9403
rect 4594 9397 4644 9403
rect 2104 9385 2154 9391
rect 2424 9385 2474 9391
rect 1203 9375 1231 9381
rect 1443 9375 1471 9381
rect 1600 9375 1651 9381
rect 1781 9370 1831 9376
rect 2838 9370 2888 9376
rect 2910 9370 2960 9376
rect 4594 9370 4644 9376
rect 4666 9370 4716 9376
rect 2104 9361 2154 9366
rect 2284 9360 2334 9366
rect 2424 9361 2474 9366
rect 1252 9345 1280 9351
rect 1394 9345 1422 9352
rect 1529 9345 1579 9351
rect 1852 9346 1902 9352
rect 2838 9328 2888 9334
rect 2910 9328 2960 9334
rect 4594 9328 4644 9334
rect 4666 9328 4716 9334
rect 2104 9319 2154 9324
rect 2284 9318 2334 9324
rect 2424 9319 2474 9324
rect 1252 9303 1280 9309
rect 1394 9303 1422 9310
rect 1529 9303 1579 9309
rect 1852 9304 1902 9310
rect 1199 9036 1227 9042
rect 1439 9036 1467 9042
rect 1596 9036 1647 9042
rect 1777 9031 1827 9037
rect 1199 8994 1227 9000
rect 1439 8994 1467 9000
rect 1596 8994 1647 9000
rect 1777 8989 1827 8995
rect 2107 8990 2157 8995
rect 2287 8990 2337 8996
rect 2427 8990 2477 8995
rect 2841 8983 2891 8989
rect 2913 8983 2963 8989
rect 1248 8964 1276 8970
rect 1390 8964 1418 8971
rect 1525 8964 1575 8970
rect 1848 8965 1898 8971
rect 2107 8948 2157 8953
rect 2287 8948 2337 8954
rect 2427 8948 2477 8953
rect 2841 8941 2891 8947
rect 2913 8941 2963 8947
rect 1248 8922 1276 8928
rect 1390 8922 1418 8929
rect 1525 8922 1575 8928
rect 1848 8923 1898 8929
rect 2107 8923 2157 8929
rect 2427 8923 2477 8929
rect 2913 8914 2963 8920
rect 2107 8881 2157 8887
rect 2427 8881 2477 8887
rect 2913 8872 2963 8878
rect 1199 8861 1227 8867
rect 1439 8861 1467 8867
rect 1596 8861 1647 8867
rect 1777 8856 1827 8862
rect 2913 8831 2963 8837
rect 1199 8819 1227 8825
rect 1439 8819 1467 8825
rect 1596 8819 1647 8825
rect 2107 8820 2157 8826
rect 2427 8820 2477 8826
rect 1777 8814 1827 8820
rect 1248 8789 1276 8795
rect 1390 8789 1418 8796
rect 1525 8789 1575 8795
rect 1848 8790 1898 8796
rect 2913 8789 2963 8795
rect 2107 8778 2157 8784
rect 2427 8778 2477 8784
rect 2841 8762 2891 8768
rect 2913 8762 2963 8768
rect 2107 8754 2157 8759
rect 1248 8747 1276 8753
rect 1390 8747 1418 8754
rect 1525 8747 1575 8753
rect 1848 8748 1898 8754
rect 2287 8753 2337 8759
rect 2427 8754 2477 8759
rect 2841 8720 2891 8726
rect 2913 8720 2963 8726
rect 2107 8712 2157 8717
rect 2287 8711 2337 8717
rect 2427 8712 2477 8717
rect 1199 8686 1227 8692
rect 1439 8686 1467 8692
rect 1596 8686 1647 8692
rect 1777 8681 1827 8687
rect 2107 8670 2157 8675
rect 2287 8670 2337 8676
rect 2427 8670 2477 8675
rect 2841 8659 2891 8665
rect 2913 8659 2963 8665
rect 1199 8644 1227 8650
rect 1439 8644 1467 8650
rect 1596 8644 1647 8650
rect 1777 8639 1827 8645
rect 2107 8628 2157 8633
rect 2287 8628 2337 8634
rect 2427 8628 2477 8633
rect 1248 8614 1276 8620
rect 1390 8614 1418 8621
rect 1525 8614 1575 8620
rect 1848 8615 1898 8621
rect 2841 8617 2891 8623
rect 2913 8617 2963 8623
rect 2107 8603 2157 8609
rect 2427 8603 2477 8609
rect 2913 8590 2963 8596
rect 1248 8572 1276 8578
rect 1390 8572 1418 8579
rect 1525 8572 1575 8578
rect 1848 8573 1898 8579
rect 2107 8561 2157 8567
rect 2427 8561 2477 8567
rect 2913 8548 2963 8554
rect 1199 8511 1227 8517
rect 1439 8511 1467 8517
rect 1596 8511 1647 8517
rect 1777 8506 1827 8512
rect 2913 8506 2963 8512
rect 2107 8500 2157 8506
rect 2427 8500 2477 8506
rect 1199 8469 1227 8475
rect 1439 8469 1467 8475
rect 1596 8469 1647 8475
rect 1777 8464 1827 8470
rect 2913 8464 2963 8470
rect 2107 8458 2157 8464
rect 2427 8458 2477 8464
rect 1248 8439 1276 8445
rect 1390 8439 1418 8446
rect 1525 8439 1575 8445
rect 1848 8440 1898 8446
rect 2107 8434 2157 8439
rect 2287 8433 2337 8439
rect 2427 8434 2477 8439
rect 2841 8437 2891 8443
rect 2913 8437 2963 8443
rect 1248 8397 1276 8403
rect 1390 8397 1418 8404
rect 1525 8397 1575 8403
rect 1848 8398 1898 8404
rect 2107 8392 2157 8397
rect 2287 8391 2337 8397
rect 2427 8392 2477 8397
rect 2841 8395 2891 8401
rect 2913 8395 2963 8401
rect 7469 7523 7472 7562
rect 7511 7523 7514 7562
rect 7565 7523 7568 7562
rect 7607 7523 7610 7562
rect 7661 7523 7664 7562
rect 7703 7523 7706 7562
rect 7757 7523 7760 7562
rect 7799 7523 7802 7562
rect 7853 7523 7856 7562
rect 7895 7523 7898 7562
rect 7949 7523 7952 7562
rect 7991 7523 7994 7562
rect 7469 7362 7472 7401
rect 7511 7362 7514 7401
rect 7565 7361 7568 7400
rect 7607 7361 7610 7400
rect 7661 7361 7664 7400
rect 7703 7361 7706 7400
rect 7757 7361 7760 7400
rect 7799 7361 7802 7400
rect 7853 7361 7856 7400
rect 7895 7361 7898 7400
rect 7949 7362 7952 7401
rect 7991 7362 7994 7401
rect 7469 7201 7472 7240
rect 7511 7201 7514 7240
rect 7565 7200 7568 7239
rect 7607 7200 7610 7239
rect 7661 7200 7664 7239
rect 7703 7200 7706 7239
rect 7757 7200 7760 7239
rect 7799 7200 7802 7239
rect 7853 7200 7856 7239
rect 7895 7200 7898 7239
rect 7949 7201 7952 7240
rect 7991 7201 7994 7240
rect 7469 7040 7472 7079
rect 7511 7040 7514 7079
rect 7565 7039 7568 7078
rect 7607 7039 7610 7078
rect 7661 7039 7664 7078
rect 7703 7039 7706 7078
rect 7757 7039 7760 7078
rect 7799 7039 7802 7078
rect 7853 7039 7856 7078
rect 7895 7039 7898 7078
rect 7949 7040 7952 7079
rect 7991 7040 7994 7079
rect 7469 6879 7472 6918
rect 7511 6879 7514 6918
rect 7565 6878 7568 6917
rect 7607 6878 7610 6917
rect 7661 6878 7664 6917
rect 7703 6878 7706 6917
rect 7757 6878 7760 6917
rect 7799 6878 7802 6917
rect 7853 6878 7856 6917
rect 7895 6878 7898 6917
rect 7949 6879 7952 6918
rect 7991 6879 7994 6918
rect 7737 6828 7741 6829
rect 7469 6718 7472 6757
rect 7511 6718 7514 6757
rect 7565 6717 7568 6756
rect 7607 6717 7610 6756
rect 7661 6717 7664 6756
rect 7703 6717 7706 6756
rect 7757 6717 7760 6756
rect 7799 6717 7802 6756
rect 7853 6717 7856 6756
rect 7895 6717 7898 6756
rect 7949 6718 7952 6757
rect 7991 6718 7994 6757
rect 7469 6557 7472 6596
rect 7511 6557 7514 6596
rect 7565 6556 7568 6595
rect 7607 6556 7610 6595
rect 7661 6556 7664 6595
rect 7703 6556 7706 6595
rect 7757 6556 7760 6595
rect 7799 6556 7802 6595
rect 7853 6556 7856 6595
rect 7895 6556 7898 6595
rect 7949 6557 7952 6596
rect 7991 6557 7994 6596
rect 7469 6396 7472 6435
rect 7511 6396 7514 6435
rect 7565 6395 7568 6434
rect 7607 6395 7610 6434
rect 7661 6395 7664 6434
rect 7703 6395 7706 6434
rect 7757 6395 7760 6434
rect 7799 6395 7802 6434
rect 7853 6395 7856 6434
rect 7895 6395 7898 6434
rect 7949 6396 7952 6435
rect 7991 6396 7994 6435
rect 7469 6235 7472 6274
rect 7511 6235 7514 6274
rect 7565 6234 7568 6273
rect 7607 6234 7610 6273
rect 7661 6234 7664 6273
rect 7703 6234 7706 6273
rect 7757 6234 7760 6273
rect 7799 6234 7802 6273
rect 7853 6234 7856 6273
rect 7895 6234 7898 6273
rect 7949 6235 7952 6274
rect 7991 6235 7994 6274
rect 7469 6074 7472 6113
rect 7511 6074 7514 6113
rect 7565 6074 7568 6113
rect 7607 6074 7610 6113
rect 7661 6074 7664 6113
rect 7703 6074 7706 6113
rect 7757 6074 7760 6113
rect 7799 6074 7802 6113
rect 7853 6074 7856 6113
rect 7895 6074 7898 6113
rect 7949 6074 7952 6113
rect 7991 6074 7994 6113
<< nwell >>
rect -14876 -21561 -14873 -21516
<< metal1 >>
rect -13106 14454 -12717 14571
rect -10247 14453 -9858 14570
rect -7388 14453 -6999 14570
rect -3198 14456 -2809 14573
rect 1014 14454 1403 14571
rect 3873 14454 4262 14571
rect 6733 14454 7122 14571
rect 9592 14454 9981 14571
rect 12451 14454 12840 14571
rect 15310 14453 15699 14570
rect 18169 14453 18558 14570
rect -12554 12222 -12231 13533
rect -9695 12563 -9372 13533
rect -6836 12992 -6513 13533
rect -5582 13312 -5565 13324
rect -6879 12961 -6496 12992
rect -6879 12736 -6836 12961
rect -6513 12736 -6496 12961
rect -6879 12718 -6496 12736
rect -5617 12656 -5565 13312
rect -5623 12645 -5558 12656
rect -5623 12608 -5617 12645
rect -5565 12608 -5558 12645
rect -5623 12605 -5558 12608
rect -9711 12512 -9361 12563
rect -9711 12287 -9695 12512
rect -9372 12287 -9361 12512
rect -9711 12274 -9361 12287
rect -12771 12183 -12231 12222
rect -12771 11860 -12737 12183
rect -12512 11860 -12231 12183
rect -14015 11852 -13676 11859
rect -14112 11843 -13676 11852
rect -14435 11520 -13890 11843
rect -13704 11520 -13676 11843
rect -12771 11842 -12477 11860
rect -5617 11837 -5565 12605
rect -5277 12214 -5236 13335
rect -2566 13135 -2450 13326
rect -2566 13022 170 13135
rect -2566 13002 189 13022
rect 37 12862 170 13002
rect 1566 12911 1889 13534
rect 2730 13326 2791 13340
rect 2728 13130 2846 13326
rect 2648 13039 2846 13130
rect 2648 13021 2829 13039
rect 3172 13023 3244 13409
rect 2648 12952 2721 13021
rect 4425 12911 4748 13533
rect 7284 12911 7607 13533
rect 8177 13272 8196 13273
rect 8890 13272 8962 13409
rect 8177 13237 8962 13272
rect 8177 13024 8196 13237
rect 10143 13218 10466 13533
rect 10067 13190 10466 13218
rect 10065 13170 10466 13190
rect 10047 13073 10482 13170
rect 10047 12867 10143 13073
rect 10466 12867 10482 13073
rect 10047 12800 10482 12867
rect 13002 12752 13325 13533
rect 12972 12708 13327 12752
rect 12972 12378 13002 12708
rect 13208 12378 13327 12708
rect 12972 12347 13327 12378
rect -5289 12211 -5236 12214
rect -5289 12170 -5283 12211
rect -5242 12170 -5236 12211
rect 15861 12189 16184 13533
rect -5289 12167 -5236 12170
rect -5637 11828 -5565 11837
rect -5637 11776 -5631 11828
rect -5579 11776 -5565 11828
rect -5637 11764 -5565 11776
rect -14112 11452 -13676 11520
rect -15468 10968 -15343 11357
rect -13098 8984 -12872 8988
rect -14435 8661 -13085 8984
rect -12877 8661 -12872 8984
rect -13098 8657 -12872 8661
rect -15467 8110 -15342 8499
rect -5617 8229 -5565 11764
rect -5277 11742 -5236 12167
rect 15841 12159 16200 12189
rect 15841 11953 15861 12159
rect 16184 11953 16200 12159
rect 15841 11936 16200 11953
rect 18720 11840 19043 13533
rect -5291 11732 -5229 11742
rect -5291 11691 -5278 11732
rect -5237 11691 -5229 11732
rect -5291 11683 -5229 11691
rect 18689 11717 19065 11840
rect -5625 8226 -5562 8229
rect -5625 8174 -5621 8226
rect -5569 8174 -5562 8226
rect -5625 8169 -5562 8174
rect -5277 8127 -5236 11683
rect 18689 11512 18720 11717
rect 19043 11512 19065 11717
rect 18689 11478 19065 11512
rect 20124 11771 20465 11803
rect 20124 11448 20154 11771
rect 20353 11448 20788 11771
rect 10956 11382 11398 11443
rect 20124 11399 20465 11448
rect 10956 11350 10980 11382
rect 11202 11350 11398 11382
rect 10956 8432 11398 11350
rect 21692 10898 21817 11287
rect 19283 8912 19515 8920
rect 19283 8589 19299 8912
rect 19508 8589 20787 8912
rect 19283 8583 19515 8589
rect 10953 8420 11400 8432
rect 10953 8311 10964 8420
rect 11392 8311 11400 8420
rect 10953 8300 11400 8311
rect -5282 8124 -5234 8127
rect -5282 8080 -5278 8124
rect -5237 8080 -5234 8124
rect -5282 8077 -5234 8080
rect -12707 6125 -12484 6133
rect -14434 5802 -12695 6125
rect -12487 5802 -12484 6125
rect -12707 5787 -12484 5802
rect -15468 5250 -15343 5639
rect -12256 3266 -12015 3276
rect -14435 2943 -12232 3266
rect -12024 2943 -12015 3266
rect -12256 2933 -12015 2943
rect -15466 2391 -15341 2780
rect -11800 407 -11573 414
rect -14434 84 -11791 407
rect -11583 84 -11573 407
rect -11800 74 -11573 84
rect -15467 -467 -15342 -78
rect -11364 -2452 -11139 -2446
rect -14435 -2775 -11357 -2452
rect -11149 -2775 -11139 -2452
rect -11364 -2783 -11139 -2775
rect -15468 -3327 -15343 -2938
rect -10932 -5311 -10707 -5300
rect -14435 -5634 -10692 -5311
rect -10932 -5645 -10707 -5634
rect -15467 -6185 -15342 -5796
rect 10956 -7830 11398 8300
rect 21691 8038 21816 8427
rect 18866 6053 19102 6066
rect 18866 5730 18874 6053
rect 19083 5730 20789 6053
rect 18866 5720 19102 5730
rect 21691 5178 21816 5567
rect 18465 3194 18693 3210
rect 18465 2871 18476 3194
rect 18685 2871 20787 3194
rect 18465 2860 18693 2871
rect 21692 2322 21817 2711
rect 18035 335 18277 347
rect 18035 12 18051 335
rect 18260 12 20787 335
rect 18035 -4 18277 12
rect 21690 -539 21815 -150
rect 17646 -2524 17873 -2513
rect 17646 -2847 17657 -2524
rect 17866 -2847 20788 -2524
rect 17646 -2860 17873 -2847
rect 21692 -3397 21817 -3008
rect 17206 -5383 17436 -5375
rect 17206 -5706 20788 -5383
rect 17206 -5716 17436 -5706
rect 21692 -6258 21817 -5869
rect 10864 -7841 11398 -7830
rect -10526 -8170 -10285 -8160
rect -14435 -8493 -10503 -8170
rect -10295 -8493 -10285 -8170
rect 10864 -8283 10882 -7841
rect 11324 -8204 11398 -7841
rect 11324 -8283 11340 -8204
rect 10864 -8300 11340 -8283
rect -10526 -8511 -10285 -8493
rect -15464 -9043 -15339 -8654
rect -10098 -11029 -9852 -11022
rect -14435 -11352 -9852 -11029
rect -10098 -11357 -9852 -11352
rect -15466 -11904 -15341 -11515
rect -9661 -13888 -9421 -13874
rect -14436 -14211 -9641 -13888
rect -9433 -14211 -9421 -13888
rect -9661 -14221 -9421 -14211
rect -15467 -14763 -15342 -14374
rect -9267 -16747 -9018 -16739
rect -14436 -17070 -9244 -16747
rect -9036 -17070 -9018 -16747
rect -9267 -17089 -9018 -17070
rect -15467 -17622 -15342 -17233
rect -8820 -19606 -8585 -19596
rect -14434 -19929 -8800 -19606
rect -8592 -19929 -8585 -19606
rect -8820 -19942 -8585 -19929
rect -15466 -20481 -15341 -20092
rect -8420 -22465 -8149 -22459
rect -14434 -22788 -8370 -22465
rect -8162 -22788 -8149 -22465
rect -8420 -22800 -8149 -22788
rect -15466 -23339 -15341 -22950
<< via1 >>
rect -6836 12736 -6513 12961
rect -5617 12608 -5565 12645
rect -9695 12287 -9372 12512
rect -12737 11860 -12512 12183
rect -13890 11520 -13704 11843
rect 10143 12867 10466 13073
rect 13002 12378 13208 12708
rect -5283 12170 -5242 12211
rect -5631 11776 -5579 11828
rect -13085 8661 -12877 8984
rect 15861 11953 16184 12159
rect -5278 11691 -5237 11732
rect -5621 8174 -5569 8226
rect 18720 11512 19043 11717
rect 20154 11448 20353 11771
rect 10980 11350 11202 11382
rect 19299 8589 19508 8912
rect 10964 8311 11392 8420
rect -5278 8080 -5237 8124
rect -12695 5802 -12487 6125
rect -12232 2943 -12024 3266
rect -11791 84 -11583 407
rect -11357 -2775 -11149 -2452
rect 18874 5730 19083 6053
rect 18476 2871 18685 3194
rect 18051 12 18260 335
rect 17657 -2847 17866 -2524
rect -10503 -8493 -10295 -8170
rect 10882 -8283 11324 -7841
rect -9641 -14211 -9433 -13888
rect -9244 -17070 -9036 -16747
rect -8800 -19929 -8592 -19606
rect -8370 -22788 -8162 -22465
<< metal2 >>
rect 21381 14165 21500 14166
rect -15126 14164 -13833 14165
rect -15139 14025 -13833 14164
rect 20201 14113 21500 14165
rect 20180 14037 21500 14113
rect -15139 13873 -14910 14025
rect -15094 13869 -14910 13873
rect -15050 13017 -14910 13869
rect 21284 13905 21500 14037
rect -14423 13388 -13848 13528
rect 20116 13395 20783 13535
rect -14423 12916 -14283 13388
rect 10028 13073 10508 13153
rect -6892 12987 -6483 13012
rect -6892 12961 -2695 12987
rect -6892 12736 -6836 12961
rect -6513 12762 -2695 12961
rect 10028 12944 10143 13073
rect 8858 12867 10143 12944
rect 10466 12944 10508 13073
rect 10466 12867 10513 12944
rect -6513 12736 -6483 12762
rect 8858 12738 10513 12867
rect 20642 12844 20782 13395
rect 21284 12982 21412 13905
rect 21336 12908 21412 12982
rect -6892 12702 -6483 12736
rect 12987 12708 13318 12737
rect -5622 12651 -5560 12653
rect -5622 12645 -2707 12651
rect -5622 12608 -5617 12645
rect -5565 12614 -2707 12645
rect -5565 12608 -5560 12614
rect -5622 12607 -5560 12608
rect -9704 12538 -9366 12549
rect -9745 12512 -2695 12538
rect 12987 12531 13002 12708
rect -9745 12313 -9695 12512
rect -9704 12287 -9695 12313
rect -9372 12313 -2695 12512
rect 8858 12378 13002 12531
rect 13208 12531 13318 12708
rect 13208 12378 13350 12531
rect 8858 12325 13350 12378
rect -9372 12287 -9366 12313
rect -9704 12281 -9366 12287
rect -5287 12211 -5239 12212
rect -12758 12183 -12494 12207
rect -12758 12089 -12737 12183
rect -12766 11864 -12737 12089
rect -12758 11860 -12737 11864
rect -12512 12089 -12494 12183
rect -5287 12170 -5283 12211
rect -5242 12209 -5239 12211
rect -5242 12171 -2708 12209
rect -5242 12170 -5239 12171
rect -5287 12169 -5239 12170
rect 15826 12159 16219 12168
rect 15826 12123 15861 12159
rect -12512 11864 -2735 12089
rect 8858 11953 15861 12123
rect 16184 11953 16219 12159
rect 8858 11917 16219 11953
rect 15826 11916 16219 11917
rect -12512 11860 -12494 11864
rect -13981 11843 -13692 11851
rect -12758 11847 -12494 11860
rect -13981 11655 -13890 11843
rect -13984 11520 -13890 11655
rect -13704 11655 -13692 11843
rect -5634 11828 -5572 11831
rect -5634 11776 -5631 11828
rect -5579 11822 -5572 11828
rect -5579 11781 -2740 11822
rect -5579 11776 -5572 11781
rect -5634 11772 -5572 11776
rect 19876 11771 20447 11846
rect -5287 11732 -5233 11735
rect -5287 11691 -5278 11732
rect -5237 11691 -2744 11732
rect 18706 11717 19056 11743
rect -5287 11687 -5233 11691
rect 18706 11689 18720 11717
rect -13704 11520 -2772 11655
rect -13984 11469 -2772 11520
rect 8858 11512 18720 11689
rect 19043 11689 19056 11717
rect 19043 11512 19065 11689
rect 8858 11484 19065 11512
rect 19876 11448 20154 11771
rect 20353 11448 20447 11771
rect 8876 11382 11209 11387
rect 8876 11350 10980 11382
rect 11202 11350 11209 11382
rect 8876 11344 11209 11350
rect 19876 11282 20447 11448
rect 19832 11278 20447 11282
rect 8858 11232 20447 11278
rect -13095 11003 -2743 11211
rect 8858 11042 20431 11232
rect -13095 8992 -12887 11003
rect 19298 10804 19507 10822
rect -12679 10515 -2695 10723
rect 8858 10595 19507 10804
rect -13102 8984 -12868 8992
rect -13102 8661 -13085 8984
rect -12877 8661 -12868 8984
rect -13102 8655 -12868 8661
rect -13095 8568 -12887 8655
rect -12679 6132 -12471 10515
rect -12701 6125 -12471 6132
rect -12701 5802 -12695 6125
rect -12487 5802 -12471 6125
rect -12701 5791 -12471 5802
rect -12679 5758 -12471 5791
rect -12245 10033 -2695 10241
rect 8858 10055 19093 10264
rect -12245 3284 -12037 10033
rect -11791 9563 -2695 9771
rect 8858 9567 18685 9776
rect -12266 3266 -12009 3284
rect -12266 2943 -12232 3266
rect -12024 2943 -12009 3266
rect -12266 2924 -12009 2943
rect -12245 2920 -12037 2924
rect -11791 422 -11583 9563
rect -11356 9137 -2695 9345
rect -11807 407 -11568 422
rect -11807 84 -11791 407
rect -11583 84 -11568 407
rect -11807 65 -11568 84
rect -11791 12 -11583 65
rect -11356 -2439 -11148 9137
rect 8858 9047 18276 9256
rect -10922 8730 -2695 8938
rect -11374 -2452 -11129 -2439
rect -11374 -2775 -11357 -2452
rect -11149 -2775 -11129 -2452
rect -11374 -2791 -11129 -2775
rect -11356 -2803 -11148 -2791
rect -10922 -5290 -10714 8730
rect 8858 8543 17863 8752
rect -10506 8315 -2695 8523
rect 10955 8421 11408 8429
rect 8886 8420 11415 8421
rect -10947 -5663 -10687 -5290
rect -10922 -5696 -10714 -5663
rect -10506 -8153 -10298 8315
rect 8886 8311 10964 8420
rect 11392 8311 11415 8420
rect 8886 8306 11415 8311
rect 10955 8304 11408 8306
rect -5624 8226 -5564 8227
rect -5624 8174 -5621 8226
rect -5569 8222 -5564 8226
rect -5569 8178 -2690 8222
rect -5569 8174 -5564 8178
rect -5624 8171 -5564 8174
rect -5281 8124 -5235 8125
rect -5281 8080 -5278 8124
rect -5237 8080 -2694 8124
rect -5281 8078 -5235 8080
rect -10081 7800 -2695 8008
rect 8890 7992 17439 8201
rect -10548 -8170 -10277 -8153
rect -10548 -8493 -10503 -8170
rect -10295 -8493 -10277 -8170
rect -10548 -8520 -10277 -8493
rect -10506 -8592 -10298 -8520
rect -10081 -11015 -9873 7800
rect -9655 7374 -2695 7582
rect -10114 -11363 -9840 -11015
rect -10081 -11444 -9873 -11363
rect -9655 -13844 -9447 7374
rect -9240 6870 -2695 7078
rect -9677 -13888 -9398 -13844
rect -9677 -14211 -9641 -13888
rect -9433 -14211 -9398 -13888
rect -9677 -14249 -9398 -14211
rect -9655 -14277 -9447 -14249
rect -9240 -16722 -9032 6870
rect -8805 6309 -2695 6517
rect -9289 -16747 -9006 -16722
rect -9289 -17070 -9244 -16747
rect -9036 -17070 -9006 -16747
rect -9289 -17100 -9006 -17070
rect -9240 -17156 -9032 -17100
rect -8805 -19580 -8597 6309
rect -8389 5839 -2695 6047
rect -8840 -19606 -8575 -19580
rect -8840 -19929 -8800 -19606
rect -8592 -19929 -8575 -19606
rect -8840 -19952 -8575 -19929
rect -8805 -19953 -8597 -19952
rect -8389 -22450 -8181 5839
rect -8408 -22465 -8141 -22450
rect -8408 -22788 -8370 -22465
rect -8162 -22788 -8141 -22465
rect -8408 -22803 -8141 -22788
rect -2235 -23386 -1901 5853
rect -1269 -23816 -1067 5843
rect -863 -23659 -661 5843
rect -863 -23815 -660 -23659
rect -466 -23660 -264 5843
rect -66 -23660 136 5843
rect -863 -23816 -661 -23815
rect -467 -23816 -264 -23660
rect -67 -23816 136 -23660
rect 339 -23816 541 5843
rect 740 -23659 942 5843
rect 739 -23815 942 -23659
rect 740 -23816 942 -23815
rect 1140 -23816 1342 5843
rect 1549 -23816 1751 5843
rect 1962 -23660 2164 5843
rect 2362 -23660 2564 5843
rect 2758 -23660 2960 5843
rect 1961 -23816 2164 -23660
rect 2361 -23816 2564 -23660
rect 2757 -23816 2960 -23660
rect 3163 -23659 3365 5843
rect 3163 -23815 3366 -23659
rect 3163 -23816 3365 -23815
rect 3572 -23816 3774 5843
rect 3973 -23661 4175 5843
rect 4377 -23660 4579 5843
rect 3973 -23816 4176 -23661
rect 4377 -23816 4580 -23660
rect 4786 -23662 4988 5843
rect 4786 -23816 4989 -23662
rect 5191 -23816 5393 5843
rect 5588 -23816 5790 5843
rect 6000 -23816 6202 5843
rect 3974 -23817 4176 -23816
rect 4787 -23818 4989 -23816
rect 6413 -23817 6615 5843
rect 6814 -23816 7016 5843
rect 7215 -23648 7417 5843
rect 7215 -23814 7419 -23648
rect 7624 -23650 7826 5843
rect 7624 -23816 7827 -23650
rect 8041 -23816 8243 5843
rect 8441 -23650 8643 5843
rect 8842 -23650 9044 5843
rect 9238 -23650 9440 5843
rect 8441 -23816 8644 -23650
rect 8839 -23816 9044 -23650
rect 9237 -23816 9440 -23650
rect 9643 -23650 9845 5843
rect 10049 -23650 10251 5843
rect 17230 -5151 17439 7992
rect 17654 -2504 17863 8543
rect 18067 344 18276 9047
rect 18476 3221 18685 9567
rect 18884 6071 19093 10055
rect 19298 8927 19507 10595
rect 19278 8912 19521 8927
rect 19278 8589 19299 8912
rect 19508 8589 19521 8912
rect 19278 8573 19521 8589
rect 19298 8506 19507 8573
rect 18860 6053 19111 6071
rect 18860 5730 18874 6053
rect 19083 5730 19111 6053
rect 18860 5714 19111 5730
rect 18456 3194 18708 3221
rect 18456 2871 18476 3194
rect 18685 2871 18708 3194
rect 18456 2850 18708 2871
rect 18476 2847 18685 2850
rect 18040 335 18276 344
rect 18040 12 18051 335
rect 18260 12 18276 335
rect 18040 2 18276 12
rect 18067 -69 18276 2
rect 17637 -2524 17880 -2504
rect 17637 -2847 17657 -2524
rect 17866 -2847 17880 -2524
rect 17637 -2875 17880 -2847
rect 17231 -5341 17439 -5151
rect 17231 -5353 17440 -5341
rect 17220 -5359 17440 -5353
rect 17194 -5727 17447 -5359
rect 17220 -5729 17429 -5727
rect 21338 -6998 21412 -6964
rect 20640 -7101 20780 -7023
rect 21272 -7038 21413 -6998
rect 20639 -7113 20780 -7101
rect 21274 -7107 21412 -7038
rect 20638 -7128 20780 -7113
rect 20638 -7218 20779 -7128
rect 21273 -7224 21413 -7107
rect 10871 -7841 11331 -7836
rect 10871 -8283 10882 -7841
rect 11324 -7914 11331 -7841
rect 11324 -8082 20786 -7914
rect 11324 -8211 20799 -8082
rect 11324 -8283 11331 -8211
rect 10871 -8293 11331 -8283
rect 9643 -23816 9847 -23650
rect 10049 -23816 10253 -23650
rect -15053 -24304 -14913 -24107
rect -14423 -24337 -14283 -23971
use sky130_hilas_TopLevelTextStructure  sky130_hilas_TopLevelTextStructure_0
timestamp 1629420194
transform 1 0 -2990 0 1 6624
box 218 -793 13243 6785
use sky130_hilas_RightProtection  sky130_hilas_RightProtection_0
timestamp 1629421669
transform 1 0 22518 0 1 -15744
box -2054 8715 -826 28728
use sky130_hilas_LeftProtection  sky130_hilas_LeftProtection_0
timestamp 1629421669
transform 1 0 -13278 0 1 -15672
box -2065 -8439 -833 28728
use sky130_hilas_TopProtection  sky130_hilas_TopProtection_0
timestamp 1629421669
transform 1 0 -13875 0 1 13286
box -2 -76 34131 1170
<< labels >>
rlabel metal1 21692 -6258 21817 -5869 0 IO07
port 1 nsew
rlabel metal1 21692 -3397 21817 -3008 0 IO08
port 2 nsew
rlabel metal1 21690 -539 21815 -150 0 IO09
port 3 nsew
rlabel metal1 21692 2322 21817 2711 0 IO10
port 4 nsew
rlabel metal1 21691 5178 21816 5567 0 IO11
port 5 nsew
rlabel metal1 21691 8038 21816 8427 0 IO12
port 6 nsew
rlabel metal1 21692 10898 21817 11287 0 IO13
port 7 nsew
rlabel metal1 -15468 10968 -15343 11357 0 IO25
port 8 nsew
rlabel metal1 -15467 8110 -15342 8499 0 IO26
port 9 nsew
rlabel metal1 -15468 5250 -15343 5639 0 IO27
port 10 nsew
rlabel metal1 -15466 2391 -15341 2780 0 IO28
port 11 nsew
rlabel metal1 -15467 -467 -15342 -78 0 IO29
port 12 nsew
rlabel metal1 -15468 -3327 -15343 -2938 0 IO30
port 13 nsew
rlabel metal1 -15467 -6185 -15342 -5796 0 IO31
port 14 nsew
rlabel metal1 -15464 -9043 -15339 -8654 0 IO32
port 15 nsew
rlabel metal1 -15466 -11904 -15341 -11515 0 IO33
port 16 nsew
rlabel metal1 -15467 -14763 -15342 -14374 0 IO34
port 17 nsew
rlabel metal1 -15467 -17622 -15342 -17233 0 IO35
port 18 nsew
rlabel metal1 -15466 -20481 -15341 -20092 0 IO36
port 19 nsew
rlabel metal1 -15466 -23339 -15341 -22950 0 IO37
port 20 nsew
rlabel metal2 -15139 13873 -14971 14164 0 VSSA1
port 21 nsew
rlabel metal1 -13106 14454 -12717 14571 0 ANALOG10
port 22 nsew
rlabel metal1 -10247 14453 -9858 14570 0 ANALOG09
port 23 nsew
rlabel metal1 -7388 14453 -6999 14570 0 ANALOG08
port 24 nsew
rlabel metal1 -3198 14456 -2809 14573 0 ANALOG07
port 25 nsew
rlabel metal1 1014 14454 1403 14571 0 ANALOG06
port 26 nsew
rlabel metal1 3873 14454 4262 14571 0 ANALOG05
port 27 nsew
rlabel metal1 6733 14454 7122 14571 0 ANALOG04
port 28 nsew
rlabel metal1 9592 14454 9981 14571 0 ANALOG03
port 29 nsew
rlabel metal1 12451 14454 12840 14571 0 ANALOG02
port 30 nsew
rlabel metal1 15310 14453 15699 14570 0 ANALOG01
port 31 nsew
rlabel metal1 18169 14453 18558 14570 0 ANALOG00
port 32 nsew
rlabel metal2 21381 13908 21500 14166 0 VSSA1
port 33 nsew
rlabel metal2 -14423 -24337 -14283 -24197 0 VDDA1
port 34 nsew
rlabel metal2 -15053 -24304 -14913 -24164 0 VSSA1
port 33 nsew
rlabel metal2 20639 -7218 20779 -7101 0 VDDA1
port 34 nsew
rlabel metal2 21273 -7224 21413 -7107 0 VSSA1
port 33 nsew
rlabel metal2 -1269 -23816 -1067 -23660 0 LADATAOUT00
port 36 nsew
rlabel metal2 -862 -23815 -660 -23659 0 LADATAOUT01
port 35 nsew
rlabel metal2 -467 -23816 -265 -23660 0 LADATAOUT02
port 37 nsew
rlabel metal2 -67 -23816 135 -23660 0 LADATAOUT03
port 38 nsew
rlabel metal2 339 -23816 541 -23660 0 LADATAOUT04
port 39 nsew
rlabel metal2 739 -23815 941 -23659 0 LADATAOUT05
port 40 nsew
rlabel metal2 1140 -23816 1342 -23660 0 LADATAOUT06
port 41 nsew
rlabel metal2 1549 -23816 1751 -23660 0 LADATAOUT07
port 42 nsew
rlabel metal2 1961 -23816 2163 -23660 0 LADATAOUT08
port 43 nsew
rlabel metal2 2361 -23816 2563 -23660 0 LADATAOUT09
port 44 nsew
rlabel metal2 2757 -23816 2959 -23660 0 LADATAOUT10
port 45 nsew
rlabel metal2 3164 -23815 3366 -23659 0 LADATAOUT11
port 46 nsew
rlabel metal2 3572 -23816 3774 -23660 0 LADATAOUT12
port 47 nsew
rlabel metal2 3974 -23817 4176 -23661 0 LADATAOUT13
port 48 nsew
rlabel metal2 4378 -23816 4580 -23660 0 LADATAOUT14
port 49 nsew
rlabel metal2 4787 -23818 4989 -23662 0 LADATAOUT15
port 50 nsew
rlabel metal2 5191 -23816 5393 -23660 0 LADATA16
port 51 nsew
rlabel metal2 5588 -23816 5790 -23660 0 LADATAOUT17
port 52 nsew
rlabel metal2 6000 -23815 6202 -23659 0 LADATAOUT18
port 53 nsew
rlabel metal2 6413 -23817 6615 -23661 0 LADATAOUT19
port 54 nsew
rlabel metal2 6814 -23816 7016 -23660 0 LADATAOUT20
port 55 nsew
rlabel metal2 7215 -23814 7419 -23648 0 LADATAOUT21
port 56 nsew
rlabel metal2 7624 -23816 7827 -23650 0 LADATAOUT22
port 57 nsew
rlabel metal2 8039 -23816 8242 -23650 0 LADATAOUT23
port 58 nsew
rlabel metal2 8441 -23816 8644 -23650 0 LADATAOUT24
port 59 nsew
rlabel metal2 8839 -23816 9042 -23650 0 LADATAIN00
port 60 nsew
rlabel metal2 9237 -23816 9440 -23650 0 LADATAIN01
port 61 nsew
rlabel metal2 9644 -23816 9847 -23650 0 LADATAIN02
port 62 nsew
rlabel metal2 10050 -23816 10253 -23650 0 LADATAIN03
port 63 nsew
rlabel metal2 20683 -8211 20799 -8085 0 VCCA
port 64 nsew
<< end >>
