magic
tech sky130A
timestamp 1628164971
<< nwell >>
rect -83 185 -27 382
<< psubdiff >>
rect -74 34 -45 63
rect -74 17 -68 34
rect -51 17 -45 34
rect -74 0 -45 17
rect -74 -17 -68 0
rect -51 -17 -45 0
rect -74 -30 -45 -17
<< nsubdiff >>
rect -73 298 -45 310
rect -73 281 -69 298
rect -52 281 -45 298
rect -73 264 -45 281
rect -73 247 -69 264
rect -52 247 -45 264
rect -73 218 -45 247
<< psubdiffcont >>
rect -68 17 -51 34
rect -68 -17 -51 0
<< nsubdiffcont >>
rect -69 281 -52 298
rect -69 247 -52 264
<< poly >>
rect -326 160 -247 175
rect -155 160 -76 175
rect -327 124 -248 139
rect -155 124 -76 139
<< locali >>
rect -69 298 -52 306
rect -69 239 -52 247
rect -68 0 -51 17
<< viali >>
rect -69 264 -52 281
rect -68 34 -51 51
rect -68 -34 -51 -17
<< metal1 >>
rect -75 288 -48 305
rect -77 285 -45 288
rect -77 259 -74 285
rect -48 259 -45 285
rect -77 256 -45 259
rect -75 238 -48 256
rect -28 111 -27 134
rect -74 51 -45 54
rect -74 34 -68 51
rect -51 34 -45 51
rect -74 23 -45 34
rect -74 -3 -72 23
rect -46 -3 -45 23
rect -74 -17 -45 -3
rect -74 -34 -68 -17
rect -51 -34 -45 -17
rect -74 -37 -45 -34
<< via1 >>
rect -74 281 -48 285
rect -74 264 -69 281
rect -69 264 -52 281
rect -52 264 -48 281
rect -74 259 -48 264
rect -72 -3 -46 23
<< metal2 >>
rect -380 392 -184 414
rect -95 400 -27 421
rect -380 315 -305 336
rect -210 317 -27 338
rect -380 314 -353 315
rect -77 285 -45 288
rect -77 259 -74 285
rect -48 282 -45 285
rect -48 261 -27 282
rect -48 259 -45 261
rect -77 256 -45 259
rect -380 215 -355 237
rect -380 159 -82 180
rect -380 119 -82 140
rect -380 61 -355 83
rect -75 23 -43 26
rect -75 -3 -72 23
rect -46 21 -43 23
rect -46 0 -27 21
rect -46 -3 -43 0
rect -75 -6 -43 -3
rect -380 -74 -309 -53
rect -214 -72 -27 -50
rect -380 -119 -181 -97
rect -96 -116 -27 -95
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_1
timestamp 1627744303
transform 0 -1 -53 1 0 169
box -9 -26 24 29
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1628164971
transform 1 0 -179 0 1 402
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628164971
transform 1 0 -108 0 1 408
box -14 -15 20 18
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_1
timestamp 1627744303
transform 1 0 -349 0 1 187
box 147 -22 266 265
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1628164971
transform 1 0 -296 0 1 324
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628164971
transform 1 0 -227 0 1 325
box -14 -15 20 18
use sky130_hilas_poly2m1  sky130_hilas_poly2m1_0
timestamp 1628164971
transform 1 0 -349 0 -1 185
box -9 -26 24 25
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_0
timestamp 1627744303
transform 1 0 -467 0 1 187
box 147 -22 266 265
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1628164971
transform 1 0 -349 0 1 221
box -9 -10 23 22
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_0
timestamp 1627744303
transform 0 -1 -54 1 0 115
box -9 -26 24 29
use sky130_hilas_li2m2  sky130_hilas_li2m2_7
timestamp 1628164971
transform 1 0 -177 0 1 -108
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_6
timestamp 1628164971
transform 1 0 -112 0 1 -108
box -14 -15 20 18
use sky130_hilas_nFETmed  sky130_hilas_nFETmed_0
timestamp 1627744303
transform 1 0 -171 0 1 -99
box -12 -44 70 228
use sky130_hilas_li2m2  sky130_hilas_li2m2_4
timestamp 1628164971
transform 1 0 -299 0 1 -64
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_5
timestamp 1628164971
transform 1 0 -229 0 1 -64
box -14 -15 20 18
use sky130_hilas_poly2m1  sky130_hilas_poly2m1_1
timestamp 1628164971
transform -1 0 -335 0 1 114
box -9 -26 24 25
use sky130_hilas_nFETmed  sky130_hilas_nFETmed_1
timestamp 1627744303
transform 1 0 -290 0 1 -99
box -12 -44 70 228
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1628164971
transform 1 0 -349 0 1 66
box -9 -10 23 22
<< labels >>
rlabel metal2 -380 215 -371 237 0 GATE1P
port 3 nsew analog default
rlabel metal2 -380 159 -372 180 0 GATE2P
port 2 nsew analog default
rlabel metal2 -380 119 -372 140 0 GATE2N
port 4 nsew analog default
rlabel metal2 -380 62 -372 83 0 GATE1N
port 1 nsew analog default
rlabel metal2 -37 400 -27 421 0 DRAIN2P
port 12 nsew analog default
rlabel metal2 -37 317 -27 338 0 DRAIN1P
port 11 nsew analog default
rlabel metal2 -380 314 -372 336 0 SOURCE1P
port 5 nsew analog default
rlabel metal2 -380 392 -372 414 0 SOURCE2P
port 6 nsew analog default
rlabel metal2 -380 -74 -373 -53 0 SOURCE1N
port 8 nsew analog default
rlabel metal2 -380 -119 -373 -97 0 SOURCE2N
port 7 nsew analog default
rlabel metal2 -34 -72 -27 -50 0 DRAIN1N
port 9 nsew analog default
rlabel metal2 -34 -116 -27 -95 0 DRAIN2N
port 10 nsew analog default
rlabel metal2 -38 0 -27 21 0 VGND
port 14 nsew
rlabel metal2 -36 261 -27 282 0 WELL
port 15 nsew
<< end >>
