magic
tech sky130A
timestamp 1627737364
<< error_s >>
rect -87 536 -60 543
rect 116 523 133 528
rect -87 494 -60 501
rect -87 470 -60 477
rect -87 428 -60 435
rect -87 388 -60 395
rect -87 346 -60 353
rect -87 322 -60 329
rect -87 280 -60 287
rect -87 240 -60 247
rect -87 198 -60 205
rect -87 174 -60 181
rect -87 132 -60 139
rect -87 92 -60 99
rect -87 50 -60 57
rect -87 26 -60 33
rect 92 20 116 25
rect -87 -16 -60 -9
<< metal1 >>
rect -41 -22 -7 550
rect 26 -21 53 549
<< metal2 >>
rect -136 507 118 530
rect -110 293 155 316
rect -136 211 155 233
rect -137 -6 134 17
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_1
timestamp 1627737364
transform 1 0 -113 0 1 131
box -59 -5 125 122
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_0
timestamp 1627737364
transform 1 0 -113 0 -1 100
box -59 -5 125 122
use sky130_hilas_pFETmirror02  sky130_hilas_pFETmirror02_0
timestamp 1627737364
transform 1 0 88 0 1 -111
box -61 89 67 373
use sky130_hilas_pFETmirror02  sky130_hilas_pFETmirror02_1
timestamp 1627737364
transform 1 0 88 0 -1 635
box -61 89 67 373
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1627737364
transform 1 0 98 0 1 3
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1627737364
transform 1 0 106 0 1 228
box -14 -15 20 18
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1627737364
transform 1 0 41 0 1 126
box -10 -8 13 21
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_2
timestamp 1627737364
transform 1 0 -113 0 1 427
box -59 -5 125 122
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_3
timestamp 1627737364
transform 1 0 -113 0 -1 396
box -59 -5 125 122
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1627737364
transform 1 0 102 0 1 522
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1627737364
transform 1 0 107 0 1 300
box -14 -15 20 18
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1627737364
transform 1 0 41 0 1 385
box -10 -8 13 21
<< labels >>
rlabel metal2 144 293 155 316 0 output1
rlabel space 144 211 155 234 0 output2
<< end >>
