* Copyright 2020 The Hilas PDK Authors
* 
* This file is part of HILAS.
* 
* HILAS is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published by
* the Free Software Foundation, version 3 of the License.
* 
* HILAS is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
* 
* You should have received a copy of the GNU Lesser General Public License
* along with HILAS.  If not, see <https://www.gnu.org/licenses/>.
* 
* Licensed under the Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
* https://www.gnu.org/licenses/lgpl-3.0.en.html
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
* SPDX-License-Identifier: LGPL-3.0
* 
* 

* NGSPICE file created from sky130_hilas_TACoreBlock.ext - technology: sky130A

.subckt sky130_hilas_TunCap01 VSUBS
X0 a_n2872_n666# w_n2902_n800# w_n2902_n800# sky130_fd_pr__cap_var w=590000u l=500000u
.ends

.subckt sky130_hilas_horizPcell01 VSUBS
X0 w_n578_94# a_n300_94# a_n344_162# w_n578_94# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
X1 a_n344_286# a_n578_238# a_n502_286# w_n578_94# sky130_fd_pr__pfet_g5v0d10v5 w=300000u l=500000u
X2 a_n344_162# a_n578_238# a_n508_162# w_n578_94# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
.ends

.subckt sky130_hilas_FGVaractorCapacitor VSUBS
X0 a_n1882_n672# w_n1914_n790# w_n1914_n790# sky130_fd_pr__cap_var w=1.11e+06u l=640000u
.ends


* Top level circuit sky130_hilas_TACoreBlock

Xsky130_hilas_TunCap01_0 VSUBS sky130_hilas_TunCap01
Xsky130_hilas_horizPcell01_0 VSUBS sky130_hilas_horizPcell01
Xsky130_hilas_FGVaractorCapacitor_0 VSUBS sky130_hilas_FGVaractorCapacitor
X0 a_n16_78# a_n42_20# a_n16_n38# VSUBS sky130_fd_pr__nfet_01v8 w=330000u l=290000u
.end

