magic
tech sky130A
magscale 1 2
timestamp 1627401095
<< error_s >>
rect 122 1496 166 1524
rect 636 1494 682 1522
rect 1338 1510 1382 1666
rect 1338 1498 1506 1510
rect 2332 1502 2386 1530
rect 0 1398 28 1434
rect 2564 1254 2592 1288
rect 766 1174 788 1252
rect 726 1172 792 1174
rect 766 1160 788 1172
rect 794 1146 816 1224
rect 1022 1148 1214 1174
rect 2206 1166 2310 1182
rect 2310 1157 2366 1166
rect 2914 1158 3014 1178
rect 2852 1157 2914 1158
rect 698 1144 820 1146
rect 794 1132 816 1144
rect 0 1096 28 1132
rect 994 1120 1242 1146
rect 968 1110 1244 1118
rect 968 1082 970 1090
rect 1024 1082 1216 1090
rect 1286 1080 1356 1088
rect 2206 1082 2310 1098
rect 2914 1074 3014 1094
rect 840 1036 946 1054
rect 786 1025 840 1036
rect 946 1025 1002 1036
rect 1198 1034 1302 1054
rect 2058 1036 2164 1054
rect 2352 1036 2456 1056
rect 1142 1028 1198 1034
rect 1016 1025 1198 1028
rect 2004 1025 2058 1036
rect 2456 1027 2510 1036
rect 2772 1034 2872 1056
rect 3056 1034 3156 1056
rect 2714 1027 2772 1034
rect 786 986 791 1025
rect 1016 1008 1164 1025
rect 1014 976 1164 1008
rect 2004 986 2009 1025
rect 2562 986 2588 994
rect 840 952 946 970
rect 1014 954 1068 976
rect 1112 948 1164 976
rect 1198 950 1302 970
rect 2058 952 2164 970
rect 2352 952 2456 972
rect 2562 966 2564 986
rect 2590 952 2592 966
rect 2772 950 2872 972
rect 3056 950 3156 972
rect 884 846 1216 872
rect 2206 864 2310 880
rect 2310 855 2366 864
rect 2914 856 3014 876
rect 2852 855 2914 856
rect 0 794 28 830
rect 884 828 1244 844
rect 880 818 1244 828
rect 880 816 1002 818
rect 880 808 1244 816
rect 908 788 974 800
rect 908 780 1216 788
rect 1286 778 1356 786
rect 2206 780 2310 796
rect 2914 772 3014 792
rect 840 734 946 752
rect 786 723 840 734
rect 946 723 1002 734
rect 1198 732 1302 752
rect 2058 734 2164 752
rect 2352 734 2456 754
rect 1142 726 1198 732
rect 1060 723 1198 726
rect 2004 723 2058 734
rect 2456 725 2510 734
rect 2772 732 2872 754
rect 3056 732 3156 754
rect 2714 725 2772 732
rect 786 684 791 723
rect 1060 708 1162 723
rect 1060 674 1168 708
rect 2004 684 2009 723
rect 2562 684 2588 692
rect 840 650 946 668
rect 1110 650 1168 674
rect 1198 648 1302 668
rect 2058 650 2164 668
rect 2352 650 2456 670
rect 2562 664 2564 684
rect 2590 650 2592 664
rect 2772 648 2872 670
rect 3056 648 3156 670
rect 892 546 1216 570
rect 2206 562 2310 578
rect 2310 553 2366 562
rect 2914 554 3014 574
rect 2852 553 2914 554
rect 892 518 1244 542
rect 974 516 1096 518
rect 974 506 1244 516
rect 1002 488 1068 500
rect 1002 478 1216 488
rect 1286 476 1356 484
rect 2206 478 2310 494
rect 840 432 946 450
rect 1026 446 1068 452
rect 1026 434 1066 446
rect 786 421 840 432
rect 946 421 1002 432
rect 1198 430 1302 450
rect 1142 424 1198 430
rect 1054 421 1198 424
rect 786 382 791 421
rect 1054 406 1160 421
rect 1060 400 1160 406
rect 1060 372 1166 400
rect 1338 386 1382 476
rect 2914 470 3014 490
rect 2058 432 2164 450
rect 2352 432 2456 452
rect 840 348 946 366
rect 1108 342 1166 372
rect 1274 366 1382 386
rect 2004 421 2058 432
rect 2456 423 2510 432
rect 2772 430 2872 452
rect 3056 430 3156 452
rect 2714 423 2772 430
rect 2004 382 2009 421
rect 2562 384 2588 390
rect 1198 346 1302 366
rect 1338 318 1382 366
rect 2058 348 2164 366
rect 2352 348 2456 368
rect 2562 362 2564 384
rect 2590 350 2592 362
rect 2772 346 2872 368
rect 3056 346 3156 368
rect 2352 342 2456 344
rect 2772 342 2872 344
rect 1382 308 1506 318
rect 2332 308 2386 336
rect 2206 262 2310 278
rect 2310 253 2366 262
rect 2914 254 3014 274
rect 2852 253 2914 254
rect 2206 178 2310 194
rect 2914 170 3014 190
rect 2058 132 2164 150
rect 2352 132 2456 152
rect 2004 121 2058 132
rect 2456 123 2510 132
rect 2772 130 2872 152
rect 3056 130 3156 152
rect 2714 123 2772 130
rect 2004 82 2009 121
rect 2058 48 2164 66
rect 2352 48 2456 68
rect 2772 46 2872 68
rect 3056 46 3156 68
<< nwell >>
rect 1338 1498 1382 1510
rect 1338 308 1382 318
<< metal1 >>
rect 122 1496 166 1512
rect 636 1494 682 1512
rect 734 1442 788 1500
rect 1338 1498 1382 1510
rect 2332 1502 2386 1512
rect 726 1388 732 1442
rect 786 1388 792 1442
rect 918 1404 972 1414
rect 734 1232 788 1388
rect 732 1226 788 1232
rect 786 1172 788 1226
rect 732 1166 788 1172
rect 734 1160 788 1166
rect 826 1306 880 1320
rect 826 896 880 1252
rect 918 1122 972 1350
rect 1108 1314 1166 1324
rect 1104 1308 1166 1314
rect 1162 1250 1166 1308
rect 1104 1244 1166 1250
rect 908 1068 914 1122
rect 968 1068 974 1122
rect 824 890 880 896
rect 878 836 880 890
rect 824 830 880 836
rect 826 596 880 830
rect 918 806 972 1068
rect 914 800 972 806
rect 968 746 972 800
rect 914 740 972 746
rect 918 736 972 740
rect 1012 1014 1066 1026
rect 1012 1008 1068 1014
rect 1012 954 1014 1008
rect 1012 948 1068 954
rect 1108 1000 1166 1244
rect 1108 948 1112 1000
rect 1164 948 1166 1000
rect 826 590 886 596
rect 826 536 832 590
rect 826 530 886 536
rect 826 520 880 530
rect 1012 506 1066 948
rect 1008 500 1066 506
rect 1062 446 1066 500
rect 1008 440 1066 446
rect 1012 434 1066 440
rect 1108 714 1166 948
rect 1108 708 1168 714
rect 1108 650 1110 708
rect 1108 644 1168 650
rect 1108 400 1166 644
rect 1108 336 1166 342
rect 1338 308 1382 318
rect 2332 308 2386 318
<< via1 >>
rect 732 1388 786 1442
rect 918 1350 972 1404
rect 732 1172 786 1226
rect 826 1252 880 1306
rect 1104 1250 1162 1308
rect 914 1068 968 1122
rect 824 836 878 890
rect 914 746 968 800
rect 1014 954 1068 1008
rect 1112 948 1164 1000
rect 832 536 886 590
rect 1008 446 1062 500
rect 1110 650 1168 708
rect 1108 342 1166 400
<< metal2 >>
rect 742 1480 1216 1482
rect 738 1450 1216 1480
rect 738 1448 792 1450
rect 732 1442 792 1448
rect 0 1398 22 1434
rect 686 1398 732 1434
rect 786 1398 792 1442
rect 732 1382 786 1388
rect 912 1350 918 1404
rect 972 1392 978 1404
rect 972 1360 1216 1392
rect 972 1350 978 1360
rect 820 1300 826 1306
rect 686 1264 826 1300
rect 820 1252 826 1264
rect 880 1300 886 1306
rect 880 1262 890 1300
rect 880 1252 886 1262
rect 1098 1250 1104 1308
rect 1162 1294 1168 1308
rect 1162 1262 1216 1294
rect 1162 1250 1168 1262
rect 2564 1254 2590 1288
rect 726 1172 732 1226
rect 786 1214 792 1226
rect 786 1182 1054 1214
rect 786 1172 792 1182
rect 1022 1180 1054 1182
rect 1022 1148 1214 1180
rect 0 1096 22 1132
rect 686 1128 958 1132
rect 686 1122 968 1128
rect 686 1096 914 1122
rect 968 1068 970 1090
rect 914 1062 970 1068
rect 924 1058 970 1062
rect 1024 1058 1216 1090
rect 1024 1008 1056 1058
rect 1008 998 1014 1008
rect 686 962 1014 998
rect 1008 954 1014 962
rect 1068 954 1074 1008
rect 1106 948 1112 1000
rect 1164 992 1170 1000
rect 1164 960 1216 992
rect 1164 948 1170 960
rect 2564 952 2590 986
rect 818 836 824 890
rect 878 878 884 890
rect 878 846 1216 878
rect 878 836 884 846
rect 0 794 22 830
rect 908 746 914 800
rect 968 788 974 800
rect 968 756 1216 788
rect 968 746 974 756
rect 1104 696 1110 708
rect 686 660 1110 696
rect 1104 650 1110 660
rect 1168 696 1174 708
rect 1168 690 1202 696
rect 1168 658 1216 690
rect 1168 650 1174 658
rect 2564 650 2590 684
rect 826 536 832 590
rect 886 578 892 590
rect 886 546 1216 578
rect 886 536 892 546
rect 1002 446 1008 500
rect 1062 488 1068 500
rect 1062 456 1216 488
rect 1062 446 1068 456
rect 1102 342 1108 400
rect 1166 390 1172 400
rect 1166 358 1216 390
rect 1166 342 1172 358
rect 2564 350 2590 384
use sky130_hilas_VinjNOR3  VinjNOR3_2
timestamp 1627400472
transform 1 0 1888 0 1 602
box 0 0 1376 328
use sky130_hilas_VinjNOR3  VinjNOR3_1
timestamp 1627400472
transform 1 0 1888 0 1 300
box 0 0 1376 328
use sky130_hilas_VinjNOR3  VinjNOR3_3
timestamp 1627400472
transform 1 0 1888 0 1 904
box 0 0 1376 328
use sky130_hilas_VinjNOR3  VinjNOR3_0
timestamp 1627400472
transform 1 0 1888 0 1 0
box 0 0 1376 328
use sky130_hilas_VinjInv2  VinjInv2_0
timestamp 1627400364
transform 1 0 672 0 1 904
box 0 0 722 328
use sky130_hilas_VinjInv2  VinjInv2_1
timestamp 1627400364
transform 1 0 672 0 1 602
box 0 0 722 328
use sky130_hilas_VinjInv2  VinjInv2_2
timestamp 1627400364
transform 1 0 672 0 1 300
box 0 0 722 328
<< labels >>
rlabel metal2 2564 1254 2590 1288 0 OUTPUT00
port 1 nsew
rlabel metal2 2564 952 2590 986 0 OUTPUT01
port 2 nsew
rlabel metal2 2564 650 2590 684 0 OUTPUT10
port 3 nsew
rlabel metal2 2564 350 2590 384 0 OUTPUT11
port 4 nsew
rlabel metal1 2332 1502 2386 1512 0 VGND
port 5 nsew
rlabel metal1 2332 308 2386 318 0 VGND
port 5 nsew
rlabel metal1 1338 308 1382 318 0 VINJ
port 6 nsew
rlabel metal1 1338 1498 1382 1510 0 VINJ
port 6 nsew
rlabel metal2 0 1398 22 1434 0 IN1
port 8 nsew
rlabel metal2 0 1096 22 1132 0 IN2
port 7 nsew
rlabel metal2 0 794 22 830 0 ENABLE
port 9 nsew
rlabel metal1 122 1496 166 1512 0 VINJ
port 6 nsew
rlabel metal1 636 1494 682 1512 0 VGND
port 5 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
