magic
tech sky130A
timestamp 1624408866
<< psubdiff >>
rect -2678 -72 2737 -55
rect -2678 -89 -2671 -72
rect 2691 -89 2737 -72
rect -2678 -103 2737 -89
<< psubdiffcont >>
rect -2671 -89 2691 -72
<< poly >>
rect -2746 369 -2636 377
rect -2746 338 -2724 369
rect -2645 349 -2636 369
rect -2645 338 2730 349
rect -2746 333 2730 338
rect 2714 311 2730 333
rect -2682 295 2730 311
rect -2682 273 -2666 295
rect -2682 257 2730 273
rect 2714 234 2730 257
rect -2682 218 2730 234
rect -2682 196 -2666 218
rect -2682 180 2730 196
rect 2714 158 2730 180
rect -2680 142 2730 158
rect -2680 121 -2664 142
rect -2680 105 2731 121
rect 2715 84 2731 105
rect -2677 68 2731 84
rect -2677 46 -2661 68
rect -2677 30 2730 46
rect 2714 7 2730 30
rect -2677 -1 2730 7
rect -2677 -10 -2645 -1
rect -2653 -19 -2645 -10
rect -2506 -9 2730 -1
rect -2506 -19 -2498 -9
rect -2653 -25 -2498 -19
<< polycont >>
rect -2724 338 -2645 369
rect -2645 -19 -2506 -1
<< locali >>
rect -2840 369 -2636 377
rect -2840 366 -2724 369
rect -2840 340 -2832 366
rect -2739 340 -2724 366
rect -2840 338 -2724 340
rect -2645 338 -2636 369
rect -2840 333 -2636 338
rect -2653 -1 -2498 7
rect -2653 -19 -2645 -1
rect -2506 -19 -2498 -1
rect -2653 -23 -2498 -19
rect -2657 -33 -2498 -23
rect -2657 -50 -2649 -33
rect -2504 -50 -2498 -33
rect -2657 -59 -2498 -50
rect -2682 -60 -2498 -59
rect -2682 -70 2714 -60
rect -2682 -72 -2661 -70
rect -2682 -89 -2671 -72
rect 2704 -87 2714 -70
rect 2699 -88 2714 -87
rect 2691 -89 2714 -88
rect -2682 -97 2714 -89
<< viali >>
rect -2832 340 -2739 366
rect -2649 -50 -2504 -33
rect -2661 -72 2704 -70
rect -2661 -88 2691 -72
rect 2691 -87 2704 -72
rect 2691 -88 2699 -87
<< metal1 >>
rect -2879 377 -2718 385
rect -2879 366 -2714 377
rect -2879 340 -2832 366
rect -2739 340 -2714 366
rect -2879 333 -2714 340
rect -2879 326 -2718 333
rect -2725 -23 -2565 -9
rect -2725 -33 -2498 -23
rect -2725 -50 -2649 -33
rect -2504 -50 -2498 -33
rect 2709 -50 2762 -49
rect -2725 -54 -2498 -50
rect 2675 -54 2762 -50
rect -2725 -70 2762 -54
rect -2725 -88 -2661 -70
rect 2704 -87 2762 -70
rect 2699 -88 2762 -87
rect -2725 -112 2762 -88
rect -2725 -113 -2565 -112
rect 2713 -113 2745 -112
<< labels >>
rlabel poly -2677 -10 -2651 7 0 VGND
rlabel metal1 -2725 -113 -2696 -9 0 VGND
port 1 nsew
rlabel metal1 -2879 326 -2850 385 0 Input
<< end >>
