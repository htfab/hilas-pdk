VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_li2m2
  CLASS BLOCK ;
  FOREIGN /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_li2m2 ;
  ORIGIN 0.140 0.150 ;
  SIZE 0.340 BY 0.330 ;
  OBS
      LAYER li1 ;
        RECT -0.130 -0.120 0.200 0.140 ;
      LAYER met1 ;
        RECT -0.140 -0.150 0.180 0.170 ;
      LAYER met2 ;
        RECT -0.140 -0.150 0.170 0.180 ;
  END
END /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_li2m2
END LIBRARY

