magic
tech sky130A
timestamp 1627255200
<< nwell >>
rect -1449 -440 -1275 -256
<< mvnsubdiff >>
rect -1394 -360 -1335 -331
rect -1394 -387 -1379 -360
rect -1351 -387 -1335 -360
rect -1394 -405 -1335 -387
<< mvnsubdiffcont >>
rect -1379 -387 -1351 -360
<< locali >>
rect -1406 -360 -1351 -352
rect -1406 -395 -1351 -387
<< viali >>
rect -1406 -387 -1379 -360
<< metal1 >>
rect -1412 -360 -1373 -255
rect -1412 -387 -1406 -360
rect -1379 -387 -1373 -360
rect -1412 -441 -1373 -387
<< end >>
