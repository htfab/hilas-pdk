magic
tech sky130A
timestamp 1627758336
<< error_s >>
rect -937 567 -887 578
rect -865 567 -815 578
rect 819 567 869 578
rect 891 567 941 578
rect -815 536 -783 537
rect 787 536 819 537
rect -937 525 -887 536
rect -865 525 -815 536
rect 819 525 869 536
rect 891 525 941 536
rect -865 505 -815 517
rect 819 505 869 517
rect -896 475 -892 505
rect -815 504 -786 505
rect 790 504 819 505
rect 896 475 900 505
rect -865 463 -815 475
rect 819 463 869 475
rect -865 423 -815 435
rect 819 423 869 435
rect -896 393 -892 423
rect -815 393 -786 394
rect 790 393 819 394
rect 896 393 900 423
rect -865 381 -815 393
rect 819 381 869 393
rect -937 362 -887 373
rect -865 362 -815 373
rect 819 362 869 373
rect 891 362 941 373
rect -815 361 -783 362
rect 787 361 819 362
rect -937 320 -887 331
rect -865 320 -815 331
rect 819 320 869 331
rect 891 320 941 331
rect -937 266 -887 277
rect -865 266 -815 277
rect 819 266 869 277
rect 891 266 941 277
rect -815 235 -783 236
rect 787 235 819 236
rect -937 224 -887 235
rect -865 224 -815 235
rect 819 224 869 235
rect 891 224 941 235
rect -865 204 -815 216
rect 819 204 869 216
rect -896 174 -892 204
rect -815 203 -786 204
rect 790 203 819 204
rect 896 174 900 204
rect -865 162 -815 174
rect 819 162 869 174
rect -865 123 -815 135
rect 819 123 869 135
rect -896 93 -892 123
rect -815 93 -786 94
rect 790 93 819 94
rect 896 93 900 123
rect -865 81 -815 93
rect 819 81 869 93
rect -937 62 -887 73
rect -865 62 -815 73
rect 819 62 869 73
rect 891 62 941 73
rect -815 61 -783 62
rect 787 61 819 62
rect -937 20 -887 31
rect -865 20 -815 31
rect 819 20 869 31
rect 891 20 941 31
<< metal1 >>
rect -968 597 -952 601
rect -984 595 -952 597
rect -927 596 -908 601
rect -887 596 -871 601
rect -984 569 -981 595
rect -955 569 -952 595
rect -693 592 -669 601
rect -475 591 -437 601
rect -300 595 -276 601
rect -72 588 -32 601
rect 36 591 76 601
rect 280 596 304 601
rect 441 591 479 601
rect 673 594 697 601
rect 875 596 891 601
rect 912 596 931 601
rect 956 597 972 601
rect 956 595 988 597
rect -984 567 -952 569
rect -32 565 36 587
rect 956 569 959 595
rect 985 569 988 595
rect 956 567 988 569
rect -968 -4 -952 2
rect -927 -3 -908 3
rect -887 -3 -871 3
rect -693 -4 -669 4
rect -475 -4 -437 5
rect -300 -4 -276 3
rect -72 -4 -32 8
rect 36 -4 76 8
rect 280 -4 304 3
rect 441 -4 479 11
rect 673 -4 697 2
rect 875 -3 891 3
rect 912 -3 931 3
rect 956 -3 972 3
<< via1 >>
rect -981 569 -955 595
rect 959 569 985 595
<< metal2 >>
rect -984 595 -699 597
rect -984 569 -981 595
rect -955 587 -699 595
rect 705 595 988 597
rect 705 587 959 595
rect -955 579 959 587
rect -955 569 -942 579
rect -743 569 725 579
rect 956 569 959 579
rect 985 569 988 595
rect -984 567 -942 569
rect 956 567 988 569
rect -1004 533 -990 552
rect 999 533 1008 551
rect -1004 490 -990 509
rect 999 490 1008 508
rect -1004 390 -989 409
rect 996 390 1009 408
rect -1004 347 -991 365
rect 995 347 1009 365
rect -1004 232 -997 250
rect 1000 232 1009 250
rect -1004 189 -997 207
rect 1000 189 1009 207
rect -334 134 342 152
rect -1004 90 -997 108
rect 1000 90 1009 108
rect -1004 47 -997 65
rect 1000 47 1009 65
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_1
timestamp 1627758336
transform -1 0 -260 0 1 378
box -264 -382 744 223
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_0
timestamp 1627758336
transform 1 0 264 0 1 378
box -264 -382 744 223
<< labels >>
rlabel metal1 441 591 479 601 0 GATE2
port 1 nsew analog default
rlabel metal1 -72 -4 -32 8 0 VTUN
port 2 nsew power default
rlabel metal1 36 -4 76 8 0 VTUN
port 2 nsew power default
rlabel metal1 36 591 76 601 0 VTUN
port 2 nsew power default
rlabel metal1 -72 588 -32 601 0 VTUN
port 2 nsew power default
rlabel metal1 -475 591 -437 601 0 GATE1
port 3 nsew analog default
rlabel metal1 -475 -4 -437 5 0 GATE1
port 3 nsew analog default
rlabel metal1 956 -3 972 3 0 VINJ
port 4 nsew power default
rlabel metal1 441 -4 479 11 0 GATE2
port 1 nsew analog default
rlabel metal1 912 596 931 601 0 SelectGate2
rlabel metal1 956 596 972 601 0 VINJ
port 6 nsew power default
rlabel metal1 -968 596 -952 601 0 VINJ
port 6 nsew power default
rlabel metal1 -927 596 -908 601 0 GATESELECT1
port 10 nsew analog default
rlabel metal1 -968 -4 -952 2 0 VINJ
port 6 nsew power default
rlabel metal1 -927 -3 -908 3 0 GATESELECT1
port 10 nsew analog default
rlabel metal1 -887 596 -871 601 0 COL1
port 12 nsew analog default
rlabel metal1 -887 -3 -871 3 0 COL1
port 12 nsew analog default
rlabel metal1 912 -3 931 3 0 GATESELECT2
port 11 nsew analog default
rlabel metal1 875 -3 891 3 0 COL2
port 13 nsew analog default
rlabel metal1 875 596 891 601 0 COL2
port 13 nsew analog default
rlabel metal2 -1004 490 -997 509 0 ROW1
port 14 nsew analog default
rlabel metal2 -1004 390 -997 409 0 ROW2
port 15 nsew analog default
rlabel metal2 -1004 533 -997 552 0 DRAIN1
port 16 nsew analog default
rlabel metal2 -1004 347 -997 365 0 DRAIN2
port 17 nsew analog default
rlabel metal2 -1004 232 -997 250 0 DRAIN3
port 18 nsew analog default
rlabel metal2 -1004 189 -997 207 0 ROW3
port 19 nsew analog default
rlabel metal2 -1004 90 -997 108 0 ROW4
port 20 nsew analog default
rlabel metal2 -1004 47 -997 65 0 DRAIN4
port 21 nsew analog default
rlabel metal2 999 533 1008 551 0 DRAIN1
port 16 nsew analog default
rlabel metal2 999 490 1008 508 0 ROW1
port 14 nsew analog default
rlabel metal2 1000 390 1009 408 0 ROW2
port 15 nsew
rlabel metal2 1000 347 1009 365 0 DRAIN2
port 17 nsew analog default
rlabel metal2 1000 232 1009 250 0 DRAIN3
port 18 nsew analog default
rlabel metal2 1000 189 1009 207 0 ROW3
port 19 nsew analog default
rlabel metal2 1000 90 1009 108 0 ROW4
port 20 nsew analog default
rlabel metal2 1000 47 1009 65 0 DRAIN4
port 21 nsew
rlabel metal1 -693 595 -669 601 0 VGND
port 22 nsew
rlabel metal1 -693 -4 -669 4 0 VGND
port 22 nsew
rlabel metal1 -300 -4 -276 3 0 VGND
port 22 nsew
rlabel metal1 -300 595 -276 601 0 VGND
port 22 nsew
rlabel metal1 280 -4 304 3 0 VGND
port 22 nsew
rlabel metal1 673 -4 697 2 0 VGND
port 22 nsew
rlabel metal1 280 596 304 601 0 VGND
port 22 nsew
rlabel metal1 673 594 697 601 0 VGND
port 22 nsew
<< end >>
