magic
tech sky130A
timestamp 1625574216
<< psubdiff >>
rect -2715 816 2607 820
rect -2715 799 -2677 816
rect 2586 799 2607 816
rect -2715 796 2607 799
rect -2715 793 -2691 796
rect -2715 33 -2711 793
rect -2694 33 -2691 793
rect 2742 794 2766 820
rect -2715 17 -2691 33
rect 2742 85 2746 794
rect 2763 85 2766 794
rect 2742 65 2766 85
<< psubdiffcont >>
rect -2677 799 2586 816
rect -2711 33 -2694 793
rect 2746 85 2763 794
<< poly >>
rect -642 963 70 968
rect -642 959 43 963
rect -642 942 -632 959
rect -615 946 43 959
rect 60 946 70 963
rect -615 942 70 946
rect -642 929 70 942
rect -642 925 43 929
rect -642 908 -632 925
rect -615 912 43 925
rect 60 912 70 929
rect -615 908 70 912
rect -642 895 70 908
rect -642 891 43 895
rect -642 874 -632 891
rect -615 878 43 891
rect 60 878 70 895
rect -615 874 70 878
rect -642 861 70 874
rect -642 857 43 861
rect -642 840 -632 857
rect -615 844 43 857
rect 60 844 70 861
rect -615 840 70 844
rect -642 833 70 840
rect 2621 812 2727 818
rect 2621 795 2630 812
rect 2718 795 2727 812
rect 2621 788 2727 795
rect -2682 772 2727 788
rect -2682 746 -2666 772
rect 2621 771 2727 772
rect -2682 730 2730 746
rect -2682 704 -2666 705
rect 2714 704 2730 730
rect -2682 688 2730 704
rect -2682 665 -2666 688
rect -2682 649 2730 665
rect 2714 624 2730 649
rect -2682 608 2730 624
rect -2682 586 -2666 608
rect -2682 570 2730 586
rect -2682 547 -2666 548
rect 2714 547 2730 570
rect -2682 531 2730 547
rect -2682 507 -2666 531
rect -2682 491 2730 507
rect -2682 469 -2666 470
rect 2714 469 2730 491
rect -2682 453 2730 469
rect -2682 427 -2666 453
rect -2682 411 2730 427
rect 2714 386 2730 411
rect -2682 370 2730 386
rect -2682 349 -2667 370
rect -2682 333 2730 349
rect 2714 311 2730 333
rect -2682 295 2730 311
rect -2682 273 -2666 295
rect -2682 257 2730 273
rect 2714 234 2730 257
rect -2682 218 2730 234
rect -2682 196 -2666 218
rect -2682 180 2730 196
rect 2714 158 2730 180
rect -2680 142 2730 158
rect -2680 121 -2664 142
rect -2680 105 2731 121
rect 2715 84 2731 105
rect -2677 68 2731 84
rect -2677 46 -2661 68
rect -2677 30 2730 46
rect 2714 7 2730 30
rect -62 -1 2730 7
rect -67 -18 -50 -1
rect -33 -18 -16 -1
rect 1 -18 18 -1
rect 35 -18 52 -1
rect 69 -18 86 -1
rect 103 -18 120 -1
rect 137 -9 2730 -1
rect 137 -18 174 -9
rect -62 -27 174 -18
<< polycont >>
rect -632 942 -615 959
rect 43 946 60 963
rect -632 908 -615 925
rect 43 912 60 929
rect -632 874 -615 891
rect 43 878 60 895
rect -632 840 -615 857
rect 43 844 60 861
rect 2630 795 2718 812
rect -50 -18 -33 -1
rect -16 -18 1 -1
rect 18 -18 35 -1
rect 52 -18 69 -1
rect 86 -18 103 -1
rect 120 -18 137 -1
<< locali >>
rect -635 959 -613 967
rect -635 855 -632 959
rect -640 840 -632 855
rect -615 855 -613 959
rect 39 963 63 971
rect -615 840 -607 855
rect -640 836 -607 840
rect 39 844 43 963
rect 60 844 63 963
rect 39 836 63 844
rect -2711 799 -2677 816
rect 2586 812 2763 816
rect 2586 799 2630 812
rect -2711 795 2630 799
rect -2711 793 -2677 795
rect -2694 778 -2677 793
rect -287 789 601 795
rect -287 778 -277 789
rect -2694 776 -277 778
rect 592 778 601 789
rect 2718 794 2763 812
rect 2718 778 2746 794
rect 592 776 2746 778
rect 2746 68 2763 85
rect -2711 16 -2694 33
<< viali >>
rect -632 925 -615 942
rect -632 891 -615 908
rect -632 857 -615 874
rect 43 929 60 946
rect 43 895 60 912
rect 43 861 60 878
rect -2677 778 -287 795
rect 601 778 2718 795
rect -67 -18 -50 -1
rect -33 -18 -16 -1
rect 1 -18 18 -1
rect 35 -18 52 -1
rect 69 -18 86 -1
rect 103 -18 120 -1
rect 137 -18 154 -1
<< metal1 >>
rect -643 968 -402 1032
rect -641 942 -600 968
rect -641 925 -632 942
rect -615 925 -600 942
rect -641 908 -600 925
rect -641 891 -632 908
rect -615 891 -600 908
rect -641 874 -600 891
rect 32 946 73 979
rect 32 929 43 946
rect 60 929 73 946
rect 32 912 73 929
rect 32 895 43 912
rect 60 895 73 912
rect 32 878 73 895
rect 32 875 43 878
rect -641 857 -632 874
rect -615 857 -600 874
rect -641 833 -600 857
rect -62 861 43 875
rect 60 875 73 878
rect 60 861 174 875
rect -2716 810 -279 816
rect -2716 795 -2667 810
rect -2716 778 -2677 795
rect -287 778 -279 810
rect -2716 775 -279 778
rect -62 25 174 861
rect 601 815 2630 816
rect 595 814 2630 815
rect 595 810 2724 814
rect 595 778 601 810
rect 2687 795 2724 810
rect 2718 778 2724 795
rect 595 776 2724 778
rect 595 775 2721 776
rect -74 -1 174 25
rect -74 -18 -67 -1
rect -50 -18 -33 -1
rect -16 -18 1 -1
rect 18 -18 35 -1
rect 52 -18 69 -1
rect 86 -18 103 -1
rect 120 -18 137 -1
rect 154 -18 174 -1
rect -74 -57 174 -18
<< via1 >>
rect -2667 795 -287 810
rect -2667 784 -287 795
rect 601 795 2687 810
rect 601 784 2687 795
<< metal2 >>
rect -2749 810 2798 820
rect -2749 784 -2667 810
rect -287 784 601 810
rect 2687 784 2798 810
rect -2749 681 2798 784
rect -2749 51 2798 191
<< labels >>
rlabel metal1 -642 983 -404 1022 0 INPUT
port 2 nsew
rlabel metal1 -74 -57 174 -30 0 OUTPUT
port 3 nsew
<< end >>
