magic
tech sky130A
timestamp 1629137242
<< checkpaint >>
rect 327 1153 1810 1460
rect 327 14 2280 1153
rect 357 -297 2280 14
rect 357 -435 1873 -297
<< error_s >>
rect 56 372 62 378
rect 161 372 167 378
rect 50 308 56 314
rect 167 308 173 314
rect 0 249 223 250
rect 426 225 501 243
rect 426 161 444 225
rect 483 161 501 225
rect 426 143 501 161
rect 421 94 516 112
rect 83 50 89 56
rect 136 50 142 56
rect 449 12 450 94
rect 482 77 516 94
rect 454 69 482 77
rect 454 58 495 69
rect 454 12 476 58
rect 482 40 516 58
rect 525 51 531 57
rect 630 51 636 57
rect 477 12 516 40
rect 449 11 516 12
rect 77 0 83 6
rect 142 0 148 6
rect 519 1 525 7
rect 636 1 642 7
<< nmos >>
rect 449 40 482 69
<< ndiff >>
rect 449 69 482 94
rect 449 34 482 40
rect 449 17 457 34
rect 474 17 482 34
rect 449 11 482 17
<< pdiff >>
rect 444 161 483 225
<< ndiffc >>
rect 457 17 474 34
<< poly >>
rect 436 40 449 69
rect 482 40 495 69
<< locali >>
rect 449 17 457 34
rect 474 17 482 34
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_0
timestamp 1629137126
transform 1 0 1477 0 1 333
box 0 0 173 190
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_0
timestamp 1629137207
transform 1 0 987 0 1 195
box 0 0 256 191
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_0
timestamp 1629137168
transform 1 0 957 0 1 644
box 0 0 223 186
<< end >>
