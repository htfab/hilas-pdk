magic
tech sky130A
timestamp 1628704392
<< error_p >>
rect 118 173 135 174
rect 142 162 143 203
rect 106 150 110 162
rect 142 150 147 162
rect 142 134 143 150
rect 142 102 143 133
rect 142 44 143 73
<< nmos >>
rect 25 203 58 232
rect 110 203 143 232
rect 25 73 58 102
rect 110 73 143 102
<< ndiff >>
rect 25 256 58 260
rect 25 239 33 256
rect 50 239 58 256
rect 25 232 58 239
rect 110 256 143 260
rect 110 239 118 256
rect 135 239 143 256
rect 110 232 143 239
rect 25 196 58 203
rect 25 179 33 196
rect 50 179 58 196
rect 25 173 58 179
rect 25 125 58 132
rect 25 108 33 125
rect 50 108 58 125
rect 25 102 58 108
rect 110 196 143 203
rect 110 179 118 196
rect 135 179 143 196
rect 110 173 143 179
rect 110 126 143 133
rect 110 109 118 126
rect 135 109 143 126
rect 110 102 143 109
rect 25 66 58 73
rect 25 49 32 66
rect 50 49 58 66
rect 25 45 58 49
rect 110 67 143 73
rect 110 50 117 67
rect 136 50 143 67
rect 110 44 143 50
<< ndiffc >>
rect 33 239 50 256
rect 118 239 135 256
rect 33 179 50 196
rect 33 108 50 125
rect 118 179 135 196
rect 118 109 135 126
rect 32 49 50 66
rect 117 50 136 67
<< psubdiff >>
rect 25 161 58 173
rect 25 144 33 161
rect 50 144 58 161
rect 25 132 58 144
rect 110 162 143 173
rect 110 145 118 162
rect 135 145 143 162
rect 110 134 143 145
rect 110 133 142 134
<< psubdiffcont >>
rect 33 144 50 161
rect 118 145 135 162
<< poly >>
rect 0 203 25 232
rect 58 203 71 232
rect 96 203 110 232
rect 143 203 166 232
rect 0 102 16 203
rect 150 102 166 203
rect 0 73 25 102
rect 58 73 71 102
rect 95 73 110 102
rect 143 73 166 102
rect 0 34 16 73
rect 0 26 59 34
rect 150 33 166 73
rect 0 9 32 26
rect 50 9 59 26
rect 0 3 59 9
rect 110 25 166 33
rect 110 8 119 25
rect 136 8 166 25
rect 110 3 166 8
<< polycont >>
rect 32 9 50 26
rect 119 8 136 25
<< locali >>
rect 28 256 55 275
rect 118 257 143 275
rect 110 256 143 257
rect 25 239 33 256
rect 50 239 58 256
rect 110 239 118 256
rect 135 239 143 256
rect 21 179 33 196
rect 50 179 62 196
rect 21 172 62 179
rect 106 179 118 196
rect 135 179 147 196
rect 106 172 147 179
rect 21 162 147 172
rect 21 161 118 162
rect 21 144 33 161
rect 50 145 118 161
rect 135 145 147 162
rect 50 144 147 145
rect 21 134 147 144
rect 21 125 62 134
rect 21 108 33 125
rect 50 108 62 125
rect 106 126 147 134
rect 106 109 118 126
rect 135 109 147 126
rect 24 49 32 66
rect 50 49 58 66
rect 109 50 117 67
rect 136 50 145 67
rect 109 49 145 50
rect 32 26 50 49
rect 32 0 50 9
rect 117 25 136 49
rect 117 8 119 25
rect 117 0 136 8
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
