magic
tech sky130A
timestamp 1628704325
<< checkpaint >>
rect -630 883 663 1018
rect -630 -293 821 883
rect -472 -428 821 -293
<< error_s >>
rect 68 542 107 545
rect 68 500 107 503
rect 67 446 106 449
rect 67 404 106 407
rect 67 350 106 353
rect 67 308 106 311
rect 67 254 106 257
rect 67 212 106 215
rect 67 158 106 161
rect 67 116 106 119
rect 68 62 107 65
rect 68 20 107 23
use sky130_hilas_pFETdevice01d  sky130_hilas_pFETdevice01d_0
timestamp 1628704241
transform 1 0 85 0 1 330
box -85 -128 106 58
use sky130_hilas_pFETdevice01a  sky130_hilas_pFETdevice01a_0
timestamp 1628285143
transform 1 0 86 0 1 42
box -80 -42 81 43
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_0
timestamp 1628704221
transform 1 0 86 0 1 522
box 0 0 172 121
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_6
timestamp 1628285143
transform 1 0 85 0 1 426
box -79 -78 82 43
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_4
timestamp 1628285143
transform 1 0 85 0 1 234
box -79 -78 82 43
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_0
timestamp 1628285143
transform 1 0 85 0 1 138
box -79 -78 82 43
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
