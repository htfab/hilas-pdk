magic
tech sky130A
timestamp 1628704321
<< checkpaint >>
rect 103 1263 1690 1266
rect -148 1249 1690 1263
rect -587 -575 1690 1249
rect -587 -616 1191 -575
rect -479 -630 990 -616
<< error_s >>
rect 783 402 784 403
<< nwell >>
rect 0 618 191 619
rect 0 58 560 618
rect 760 601 888 619
rect 0 40 43 58
rect 0 17 71 40
rect 0 15 43 17
rect 760 14 888 33
<< nsubdiff >>
rect 19 535 50 572
rect 19 518 25 535
rect 42 518 50 535
rect 19 501 50 518
rect 19 484 25 501
rect 42 484 50 501
rect 19 467 50 484
rect 19 450 25 467
rect 42 450 50 467
rect 19 433 50 450
rect 19 416 25 433
rect 42 416 50 433
rect 19 399 50 416
rect 19 382 25 399
rect 42 382 50 399
rect 19 367 50 382
rect 18 232 50 265
rect 18 215 26 232
rect 43 215 50 232
rect 18 198 50 215
rect 18 181 26 198
rect 43 181 50 198
rect 18 164 50 181
rect 18 147 26 164
rect 43 147 50 164
rect 18 130 50 147
rect 18 113 26 130
rect 43 113 50 130
rect 18 96 50 113
rect 18 79 26 96
rect 43 79 50 96
rect 18 64 50 79
<< nsubdiffcont >>
rect 25 518 42 535
rect 25 484 42 501
rect 25 450 42 467
rect 25 416 42 433
rect 25 382 42 399
rect 26 215 43 232
rect 26 181 43 198
rect 26 147 43 164
rect 26 113 43 130
rect 26 79 43 96
<< locali >>
rect 67 571 101 572
rect 42 547 101 571
rect 42 498 84 547
rect 765 472 767 489
rect 784 472 790 489
rect 765 435 790 472
rect 765 419 786 435
rect 765 402 767 419
rect 784 402 786 419
rect 765 400 786 402
rect 25 365 42 382
rect 26 71 43 79
<< viali >>
rect 25 535 42 552
rect 25 501 42 518
rect 84 530 101 547
rect 84 496 101 513
rect 25 467 42 484
rect 25 433 42 450
rect 25 399 42 416
rect 767 472 784 489
rect 767 402 784 419
rect 26 232 43 249
rect 26 198 43 215
rect 26 164 43 181
rect 26 130 43 147
rect 26 96 43 113
<< metal1 >>
rect 692 605 726 619
rect 759 604 786 619
rect 22 572 75 573
rect 22 571 101 572
rect 22 565 104 571
rect 22 552 34 565
rect 22 535 25 552
rect 93 547 104 565
rect 22 518 34 535
rect 101 541 104 547
rect 101 530 107 541
rect 22 501 25 518
rect 93 513 107 530
rect 22 493 34 501
rect 101 512 107 513
rect 101 496 104 512
rect 93 493 104 496
rect 22 487 104 493
rect 762 489 794 493
rect 22 484 86 487
rect 22 467 25 484
rect 42 467 86 484
rect 22 450 86 467
rect 22 433 25 450
rect 42 433 86 450
rect 22 416 86 433
rect 22 399 25 416
rect 42 399 86 416
rect 762 403 763 489
rect 789 403 794 489
rect 762 402 767 403
rect 784 402 794 403
rect 762 401 794 402
rect 765 400 794 401
rect 22 249 86 399
rect 22 232 26 249
rect 43 232 86 249
rect 22 215 86 232
rect 22 198 26 215
rect 43 198 86 215
rect 22 181 86 198
rect 22 164 26 181
rect 43 164 86 181
rect 22 147 86 164
rect 22 130 26 147
rect 43 130 86 147
rect 22 113 86 130
rect 22 96 26 113
rect 43 96 86 113
rect 22 69 86 96
rect 44 68 86 69
rect 692 14 726 33
rect 759 14 786 35
<< via1 >>
rect 34 552 93 565
rect 34 535 42 552
rect 42 547 93 552
rect 42 535 84 547
rect 34 530 84 535
rect 84 530 93 547
rect 34 518 93 530
rect 34 501 42 518
rect 42 513 93 518
rect 42 501 84 513
rect 34 496 84 501
rect 84 496 93 513
rect 34 493 93 496
rect 763 472 767 489
rect 767 472 784 489
rect 784 472 789 489
rect 763 419 789 472
rect 763 403 767 419
rect 767 403 784 419
rect 784 403 789 419
<< metal2 >>
rect 79 572 103 619
rect 439 592 464 618
rect 27 565 103 572
rect 27 493 34 565
rect 93 537 103 565
rect 93 514 481 537
rect 93 493 103 514
rect 27 490 103 493
rect 27 489 72 490
rect 458 478 481 514
rect 545 494 570 531
rect 760 489 793 493
rect 760 478 763 489
rect 188 445 407 467
rect 458 458 763 478
rect 484 457 763 458
rect 548 409 569 438
rect 760 403 763 457
rect 789 403 793 489
rect 760 400 793 403
rect 873 348 888 370
rect 443 325 468 348
rect 1 284 147 308
rect 287 284 315 308
rect 1 283 65 284
rect 873 266 888 288
rect 392 201 569 221
rect 235 166 251 184
rect 233 165 251 166
rect 211 152 251 165
rect 211 103 247 152
rect 363 120 569 141
rect 5 17 170 40
rect 283 16 309 41
<< rmetal2 >>
rect 72 489 103 490
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1628704305
transform 1 0 733 0 1 55
box 0 0 327 581
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_2
timestamp 1628704305
transform 1 0 -90 0 1 454
box 133 -454 320 165
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1628704305
transform 1 0 241 0 -1 179
box 133 -454 320 165
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_0
timestamp 1628704305
transform 1 0 85 0 1 454
box 133 -454 320 165
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628704305
transform 1 0 89 0 1 583
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628704305
transform 1 0 173 0 1 455
box 0 0 34 33
<< labels >>
rlabel metal1 692 14 726 20 0 VGND
port 3 nsew ground default
rlabel metal1 759 14 786 20 0 VPWR
port 4 nsew power default
rlabel metal1 692 614 726 619 0 VGND
port 3 nsew ground default
rlabel metal1 759 614 786 619 0 VPWR
port 4 nsew power default
rlabel metal2 287 284 310 308 0 VIN11
port 7 nsew analog default
rlabel metal2 443 325 468 348 0 VIN21
port 6 nsew analog default
rlabel metal2 283 16 306 41 0 VIN12
port 8 nsew analog default
rlabel metal2 439 592 464 618 0 VIN22
port 5 nsew analog default
rlabel metal2 873 266 888 288 0 VOUT_AMP1
port 2 nsew analog default
rlabel metal2 873 348 888 370 0 VOUT_AMP2
port 1 nsew analog default
rlabel metal2 79 611 103 619 0 VPWR
port 4 nsew power default
rlabel metal2 43 284 50 308 0 VBIAS1
port 10 nsew analog default
rlabel metal2 43 17 50 40 0 VBIAS2
port 9 nsew analog default
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
