magic
tech sky130A
timestamp 1628704233
<< metal2 >>
rect 0 528 797 546
rect 0 485 797 503
rect 3 385 797 403
rect 3 342 797 360
rect 2 280 29 308
rect 766 282 797 310
rect 3 227 797 244
rect 3 185 797 202
rect 3 87 797 104
rect 3 43 797 60
<< metal3 >>
rect 568 270 766 331
rect 568 269 764 270
rect 765 269 766 270
rect 568 256 766 269
<< metal4 >>
rect 116 320 217 321
rect 45 270 380 320
rect 45 269 152 270
rect 316 158 379 270
rect 316 128 531 158
rect 349 127 531 128
use sky130_hilas_m22m4  sky130_hilas_m22m4_0
timestamp 1607701799
transform 1 0 38 0 1 290
box -36 -36 43 39
use sky130_hilas_CapModule03  sky130_hilas_CapModule03_0
timestamp 1607813757
transform 1 0 538 0 1 247
box -392 -247 31 336
use sky130_hilas_m22m4  sky130_hilas_m22m4_1
timestamp 1607701799
transform 1 0 750 0 1 292
box -36 -36 43 39
<< labels >>
rlabel metal2 2 280 9 308 0 CAPTERM01
port 2 nsew analog default
rlabel metal2 782 282 797 310 0 CAPTERM02
port 1 nsew analog default
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
