magic
tech sky130A
timestamp 1627744303
<< error_p >>
rect -18 20 21 23
rect -18 -22 21 -19
<< nwell >>
rect -79 -78 82 43
<< pmos >>
rect -18 -19 21 20
<< pdiff >>
rect -45 9 -18 20
rect -45 -8 -41 9
rect -24 -8 -18 9
rect -45 -19 -18 -8
rect 21 9 48 20
rect 21 -8 27 9
rect 44 -8 48 9
rect 21 -19 48 -8
<< pdiffc >>
rect -41 -8 -24 9
rect 27 -8 44 9
<< poly >>
rect -79 18 -53 33
rect -18 20 21 33
rect -68 -27 -53 18
rect -18 -27 21 -19
rect -68 -42 71 -27
rect 56 -63 71 -42
rect 56 -78 82 -63
<< locali >>
rect -41 9 -24 17
rect -41 -16 -24 -8
rect 27 9 44 17
rect 27 -16 44 -8
<< end >>
