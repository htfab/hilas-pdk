* Copyright 2020 The Hilas PDK Authors
* 
* This file is part of HILAS.
* 
* HILAS is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published by
* the Free Software Foundation, version 3 of the License.
* 
* HILAS is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
* 
* You should have received a copy of the GNU Lesser General Public License
* along with HILAS.  If not, see <https://www.gnu.org/licenses/>.
* 
* Licensed under the Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
* https://www.gnu.org/licenses/lgpl-3.0.en.html
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
* SPDX-License-Identifier: LGPL-3.0
* 
* 

* NGSPICE file created from sky130_hilas_DAC5bit01.ext - technology: sky130A

.subckt sky130_hilas_pFETdevice01 w_n158_n156# a_n90_n38# $SUB a_42_n38# a_n158_36#
X0 a_42_n38# a_n158_36# a_n90_n38# w_n158_n156# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends

.subckt sky130_hilas_pFETdevice01aa a_n160_36# $SUB w_n160_n156#
X0 a_42_n38# a_n160_36# a_n92_n38# w_n160_n156# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends

.subckt sky130_hilas_pFETdevice01a a_n160_36# $SUB w_n160_n84#
X0 a_42_n38# a_n160_36# a_n92_n38# w_n160_n84# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends

.subckt sky130_hilas_DAC6TransistorStack01 sky130_hilas_pFETdevice01_3/a_n90_n38#
+ sky130_hilas_pFETdevice01_0/a_n90_n38# sky130_hilas_pFETdevice01_6/a_n158_36# sky130_hilas_pFETdevice01_0/a_42_n38#
+ sky130_hilas_pFETdevice01_4/a_42_n38# $SUB sky130_hilas_pFETdevice01_4/a_n158_36#
+ sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01a_0/a_n160_36#
+ sky130_hilas_pFETdevice01_3/a_n158_36# sky130_hilas_pFETdevice01_3/a_42_n38# sky130_hilas_pFETdevice01_6/a_n90_n38#
+ sky130_hilas_pFETdevice01aa_0/a_n160_36# sky130_hilas_pFETdevice01_4/a_n90_n38#
+ sky130_hilas_pFETdevice01_0/a_n158_36# sky130_hilas_pFETdevice01_6/a_42_n38#
Xsky130_hilas_pFETdevice01_0 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_0/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_0/a_42_n38# sky130_hilas_pFETdevice01_0/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01_3 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_3/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_3/a_42_n38# sky130_hilas_pFETdevice01_3/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01_4 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_4/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_4/a_42_n38# sky130_hilas_pFETdevice01_4/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01_6 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_6/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_6/a_42_n38# sky130_hilas_pFETdevice01_6/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01aa_0 sky130_hilas_pFETdevice01aa_0/a_n160_36# $SUB sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01aa
Xsky130_hilas_pFETdevice01a_0 sky130_hilas_pFETdevice01a_0/a_n160_36# $SUB sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01a
.ends

.subckt sky130_hilas_pFETdevice01d w_n158_n156# a_n90_n38# $SUB a_n36_n84# a_42_n38#
+ sky130_hilas_poly2m1_0/a_n18_n16#
X0 a_42_n38# a_n36_n84# a_n90_n38# w_n158_n156# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends

.subckt sky130_hilas_DAC6TransistorStack01b sky130_hilas_pFETdevice01_0/a_n90_n38#
+ sky130_hilas_pFETdevice01_6/a_n158_36# sky130_hilas_pFETdevice01d_0/a_n90_n38# sky130_hilas_pFETdevice01d_0/a_n36_n84#
+ sky130_hilas_pFETdevice01_0/a_42_n38# sky130_hilas_pFETdevice01_4/a_42_n38# $SUB
+ sky130_hilas_pFETdevice01_4/a_n158_36# sky130_hilas_pFETdevice01a_0/a_n160_36# sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01d_0/sky130_hilas_poly2m1_0/a_n18_n16# sky130_hilas_pFETdevice01_6/a_n90_n38#
+ sky130_hilas_pFETdevice01aa_0/a_n160_36# sky130_hilas_pFETdevice01_4/a_n90_n38#
+ sky130_hilas_pFETdevice01_0/a_n158_36# sky130_hilas_pFETdevice01d_0/a_42_n38# sky130_hilas_pFETdevice01_6/a_42_n38#
Xsky130_hilas_pFETdevice01d_0 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01d_0/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01d_0/a_n36_n84# sky130_hilas_pFETdevice01d_0/a_42_n38#
+ sky130_hilas_pFETdevice01d_0/sky130_hilas_poly2m1_0/a_n18_n16# sky130_hilas_pFETdevice01d
Xsky130_hilas_pFETdevice01_0 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_0/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_0/a_42_n38# sky130_hilas_pFETdevice01_0/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01_4 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_4/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_4/a_42_n38# sky130_hilas_pFETdevice01_4/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01_6 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_6/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_6/a_42_n38# sky130_hilas_pFETdevice01_6/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01aa_0 sky130_hilas_pFETdevice01aa_0/a_n160_36# $SUB sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01aa
Xsky130_hilas_pFETdevice01a_0 sky130_hilas_pFETdevice01a_0/a_n160_36# $SUB sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01a
.ends

.subckt sky130_hilas_pFETdevice01b w_n158_n156# $SUB a_n36_n84#
X0 a_42_n38# a_n36_n84# a_n90_n38# w_n158_n156# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends

.subckt sky130_hilas_DAC6TransistorStack01c sky130_hilas_pFETdevice01_3/a_n90_n38#
+ sky130_hilas_pFETdevice01b_1/a_n36_n84# sky130_hilas_pFETdevice01_0/a_n90_n38# sky130_hilas_pFETdevice01_6/a_n158_36#
+ sky130_hilas_pFETdevice01_0/a_42_n38# $SUB sky130_hilas_pFETdevice01a_0/a_n160_36#
+ sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_3/a_n158_36#
+ sky130_hilas_pFETdevice01_3/a_42_n38# sky130_hilas_pFETdevice01_6/a_n90_n38# sky130_hilas_pFETdevice01aa_0/a_n160_36#
+ sky130_hilas_pFETdevice01_0/a_n158_36# sky130_hilas_pFETdevice01_6/a_42_n38#
Xsky130_hilas_pFETdevice01b_1 sky130_hilas_pFETdevice01a_0/w_n160_n84# $SUB sky130_hilas_pFETdevice01b_1/a_n36_n84#
+ sky130_hilas_pFETdevice01b
Xsky130_hilas_pFETdevice01_0 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_0/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_0/a_42_n38# sky130_hilas_pFETdevice01_0/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01_3 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_3/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_3/a_42_n38# sky130_hilas_pFETdevice01_3/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01_6 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_6/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_6/a_42_n38# sky130_hilas_pFETdevice01_6/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01aa_0 sky130_hilas_pFETdevice01aa_0/a_n160_36# $SUB sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01aa
Xsky130_hilas_pFETdevice01a_0 sky130_hilas_pFETdevice01a_0/a_n160_36# $SUB sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01a
.ends

.subckt sky130_hilas_DAC6TransistorStack01a sky130_hilas_pFETdevice01aa_4/a_n160_36#
+ sky130_hilas_pFETdevice01aa_3/a_n160_36# $SUB sky130_hilas_pFETdevice01a_0/a_n160_36#
+ sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01aa_2/a_n160_36#
+ sky130_hilas_pFETdevice01aa_1/a_n160_36# sky130_hilas_pFETdevice01aa_0/a_n160_36#
Xsky130_hilas_pFETdevice01aa_0 sky130_hilas_pFETdevice01aa_0/a_n160_36# $SUB sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01aa
Xsky130_hilas_pFETdevice01aa_1 sky130_hilas_pFETdevice01aa_1/a_n160_36# $SUB sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01aa
Xsky130_hilas_pFETdevice01aa_2 sky130_hilas_pFETdevice01aa_2/a_n160_36# $SUB sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01aa
Xsky130_hilas_pFETdevice01aa_3 sky130_hilas_pFETdevice01aa_3/a_n160_36# $SUB sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01aa
Xsky130_hilas_pFETdevice01aa_4 sky130_hilas_pFETdevice01aa_4/a_n160_36# $SUB sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01aa
Xsky130_hilas_pFETdevice01a_0 sky130_hilas_pFETdevice01a_0/a_n160_36# $SUB sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01a
.ends

.subckt sky130_hilas_DAC5bit01 A0 A2 A3 A4 VPWR DRAIN
Xsky130_hilas_DAC6TransistorStack01_0[0] VPWR VPWR A4 DRAIN DRAIN $SUB sky130_hilas_poly2m2_11/a_n18_n16#
+ w_1238_2040# sky130_hilas_DAC6TransistorStack01a_0/sky130_hilas_pFETdevice01aa_0/a_n160_36#
+ A3 DRAIN VPWR A4 VPWR sky130_hilas_poly2m2_12/a_n18_n16# DRAIN sky130_hilas_DAC6TransistorStack01
Xsky130_hilas_DAC6TransistorStack01_0[1] VPWR VPWR A4 DRAIN DRAIN $SUB A3 w_1238_2040#
+ sky130_hilas_poly2m2_12/a_n18_n16# A4 DRAIN VPWR A3 VPWR sky130_hilas_poly2m2_11/a_n18_n16#
+ DRAIN sky130_hilas_DAC6TransistorStack01
Xsky130_hilas_DAC6TransistorStack01_0[2] VPWR VPWR A3 DRAIN DRAIN $SUB A4 w_1238_2040#
+ sky130_hilas_poly2m2_11/a_n18_n16# A4 DRAIN VPWR A4 VPWR A3 DRAIN sky130_hilas_DAC6TransistorStack01
Xsky130_hilas_DAC6TransistorStack01_2[0] VPWR VPWR A3 DRAIN DRAIN $SUB A4 w_1238_2040#
+ A4 A4 DRAIN VPWR A2 VPWR A3 DRAIN sky130_hilas_DAC6TransistorStack01
Xsky130_hilas_DAC6TransistorStack01_2[1] VPWR VPWR A2 DRAIN DRAIN $SUB A4 w_1238_2040#
+ A3 A3 DRAIN VPWR m2_764_1430# VPWR A4 DRAIN sky130_hilas_DAC6TransistorStack01
Xsky130_hilas_DAC6TransistorStack01_2[2] VPWR VPWR m2_764_1430# DRAIN DRAIN $SUB A3
+ w_1238_2040# A4 A2 DRAIN VPWR sky130_hilas_DAC6TransistorStack01a_1/sky130_hilas_pFETdevice01aa_2/a_n160_36#
+ VPWR A4 DRAIN sky130_hilas_DAC6TransistorStack01
Xsky130_hilas_DAC6TransistorStack01b_0 VPWR A4 VPWR A0 DRAIN DRAIN $SUB A4 A3 w_1238_2040#
+ A3 VPWR A4 VPWR A4 DRAIN DRAIN sky130_hilas_DAC6TransistorStack01b
Xsky130_hilas_DAC6TransistorStack01c_0 VPWR A3 VPWR A4 DRAIN $SUB A4 w_1238_2040#
+ A4 DRAIN VPWR A3 A4 DRAIN sky130_hilas_DAC6TransistorStack01c
Xsky130_hilas_DAC6TransistorStack01a_0 sky130_hilas_poly2m2_11/a_n18_n16# A4 $SUB
+ sky130_hilas_DAC6TransistorStack01a_0/sky130_hilas_pFETdevice01a_0/a_n160_36# w_1238_2040#
+ A3 sky130_hilas_poly2m2_12/a_n18_n16# sky130_hilas_DAC6TransistorStack01a_0/sky130_hilas_pFETdevice01aa_0/a_n160_36#
+ sky130_hilas_DAC6TransistorStack01a
Xsky130_hilas_DAC6TransistorStack01a_1 m2_764_1430# sky130_hilas_DAC6TransistorStack01a_1/sky130_hilas_pFETdevice01aa_3/a_n160_36#
+ $SUB A4 w_1238_2040# sky130_hilas_DAC6TransistorStack01a_1/sky130_hilas_pFETdevice01aa_2/a_n160_36#
+ A2 A3 sky130_hilas_DAC6TransistorStack01a
.ends

