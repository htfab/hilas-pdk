magic
tech sky130A
timestamp 1628704396
<< checkpaint >>
rect -620 1149 674 1164
rect -620 1096 688 1149
rect -620 1081 689 1096
rect -620 -547 703 1081
rect -620 -562 689 -547
rect -620 -615 688 -562
rect -620 -630 674 -615
<< poly >>
rect 196 505 216 534
rect 195 228 216 307
rect 196 0 216 29
<< metal1 >>
rect 118 257 141 277
rect 244 257 267 278
use sky130_hilas_WTAsinglestage01  sky130_hilas_WTAsinglestage01_3
timestamp 1628704379
transform 1 0 108 0 1 353
box 0 0 283 143
use sky130_hilas_WTAsinglestage01  sky130_hilas_WTAsinglestage01_2
timestamp 1628704379
transform 1 0 108 0 -1 458
box 0 0 283 143
use sky130_hilas_WTAsinglestage01  sky130_hilas_WTAsinglestage01_1
timestamp 1628704379
transform 1 0 108 0 -1 181
box 0 0 283 143
use sky130_hilas_WTAsinglestage01  sky130_hilas_WTAsinglestage01_0
timestamp 1628704379
transform 1 0 108 0 1 76
box 0 0 283 143
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
