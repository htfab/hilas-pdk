magic
tech sky130A
magscale 1 2
timestamp 1627400609
<< error_s >>
rect 136 1906 236 1928
rect 280 1906 380 1928
rect 380 1844 444 1845
rect 136 1822 236 1844
rect 280 1822 380 1844
rect 280 1782 380 1806
rect 218 1722 225 1782
rect 380 1781 438 1782
rect 280 1698 380 1722
rect 1460 1692 1494 1696
rect 656 1686 690 1690
rect 1460 1654 1494 1658
rect 656 1648 690 1652
rect 280 1618 380 1642
rect 218 1558 225 1618
rect 380 1558 438 1559
rect 280 1534 380 1558
rect 136 1496 236 1518
rect 280 1496 380 1518
rect 380 1495 444 1496
rect 654 1450 688 1454
rect 1458 1438 1492 1442
rect 136 1412 236 1434
rect 280 1412 380 1434
rect 654 1412 688 1416
rect 654 1382 688 1386
rect 820 1376 826 1432
rect 1458 1400 1492 1404
rect 136 1304 236 1326
rect 280 1304 380 1326
rect 380 1242 444 1243
rect 136 1220 236 1242
rect 280 1220 380 1242
rect 514 1210 826 1376
rect 1458 1370 1492 1374
rect 1458 1332 1492 1336
rect 1458 1302 1492 1306
rect 1458 1264 1492 1268
rect 536 1208 826 1210
rect 280 1180 380 1204
rect 218 1120 225 1180
rect 380 1179 438 1180
rect 536 1178 572 1208
rect 606 1196 638 1208
rect 648 1168 666 1208
rect 768 1196 800 1208
rect 820 1176 826 1208
rect 1592 1210 1668 1358
rect 1670 1210 1922 1464
rect 1592 1190 1922 1210
rect 2398 1210 2478 1350
rect 2398 1182 2566 1210
rect 1150 1154 2016 1176
rect 1150 1152 2014 1154
rect 434 1124 496 1138
rect 1150 1126 2044 1148
rect 1150 1124 2042 1126
rect 280 1096 380 1120
rect 424 1096 524 1110
rect 280 1018 380 1042
rect 218 958 225 1018
rect 2556 1000 2576 1018
rect 380 958 438 959
rect 280 934 380 958
rect 1054 956 1174 970
rect 462 948 496 950
rect 462 920 524 922
rect 136 896 236 918
rect 280 896 380 918
rect 380 895 444 896
rect 400 866 434 870
rect 432 842 434 852
rect 438 846 490 854
rect 428 838 434 842
rect 136 812 236 834
rect 280 812 380 834
rect 432 812 434 824
rect 536 762 600 934
rect 1082 928 1146 942
rect 536 2 622 762
rect 1592 0 1668 28
<< nwell >>
rect 454 1208 1046 1210
rect 454 1178 536 1208
rect 1592 1190 1668 1210
rect 2398 1182 2478 1210
rect 454 1176 572 1178
rect 454 824 536 1176
rect 432 594 536 824
rect 454 2 536 594
<< poly >>
rect 3074 1118 3114 1210
rect 3074 0 3114 50
<< locali >>
rect 426 42 462 220
<< metal1 >>
rect 606 1196 638 1210
rect 688 1196 726 1210
rect 768 1196 800 1210
rect 1592 1190 1668 1210
rect 2398 1182 2478 1210
rect 2918 1118 2964 1210
rect 3170 1118 3216 1210
rect 1092 946 1134 1094
rect 432 594 474 824
rect 1088 272 1120 572
rect 3170 340 3216 350
rect 3162 338 3218 340
rect 3162 334 3222 338
rect 3162 280 3164 334
rect 3218 280 3222 334
rect 3162 274 3222 280
rect 1592 0 1668 20
rect 2918 0 2964 50
rect 3170 0 3216 50
<< via1 >>
rect 3164 280 3218 334
<< metal2 >>
rect 1140 1110 2670 1148
rect 424 1074 534 1110
rect 1140 1106 2704 1110
rect 2628 1068 2704 1106
rect 432 922 462 1024
rect 2548 1000 2556 1018
rect 2526 960 2768 1000
rect 2996 938 3248 970
rect 432 890 1118 922
rect 432 790 484 842
rect 442 788 476 790
rect 2546 788 2788 828
rect 2996 752 3248 784
rect 420 702 534 738
rect 1074 694 1120 696
rect 1074 688 2588 694
rect 1074 654 2600 688
rect 1074 634 1122 654
rect 432 598 1122 634
rect 2562 614 2704 654
rect 432 594 1106 598
rect 1102 554 2592 558
rect 1102 514 2704 554
rect 1102 512 1166 514
rect 424 472 534 508
rect 424 470 456 472
rect 420 322 460 422
rect 2544 390 2744 422
rect 2996 384 3248 416
rect 3158 334 3224 336
rect 420 282 1130 322
rect 3158 318 3164 334
rect 1888 284 3164 318
rect 3158 280 3164 284
rect 3218 280 3224 334
rect 3158 278 3224 280
rect 418 180 474 234
rect 2546 194 2746 228
rect 3000 198 3248 230
rect 2546 192 2734 194
rect 428 138 460 140
rect 428 102 534 138
rect 2592 102 2702 104
rect 1076 58 2702 102
rect 1076 56 2594 58
rect 1076 54 1230 56
rect 1076 46 1124 54
rect 428 6 1124 46
rect 428 4 962 6
use sky130_hilas_m12m2  sky130_hilas_m12m2_4
timestamp 1607949437
transform 1 0 1100 0 1 528
box -18 -20 46 44
use sky130_hilas_m12m2  sky130_hilas_m12m2_5
timestamp 1607949437
transform 1 0 1068 0 1 292
box -18 -20 46 44
use sky130_hilas_m12m2  sky130_hilas_m12m2_2
timestamp 1607949437
transform 1 0 1100 0 1 904
box -18 -20 46 44
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1607949437
transform 1 0 1104 0 1 1114
box -18 -20 46 44
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1607089160
transform 1 0 452 0 1 34
box -28 -30 40 36
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1607089160
transform 1 0 442 0 1 204
box -28 -30 40 36
use sky130_hilas_m12m2  sky130_hilas_m12m2_3
timestamp 1607949437
transform 1 0 446 0 1 804
box -18 -20 46 44
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1607949437
transform 1 0 442 0 1 602
box -18 -20 46 44
use sky130_hilas_WTA4stage01  sky130_hilas_WTA4stage01_0
timestamp 1607370486
transform 1 0 2790 0 1 48
box -108 2 458 1070
use sky130_hilas_swc4x1BiasCell  sky130_hilas_swc4x1BiasCell_0
timestamp 1627063197
transform -1 0 2022 0 1 764
box 0 0 2022 1210
<< labels >>
rlabel metal2 3234 938 3248 970 0 OUTPUT1
port 4 nsew analog default
rlabel metal2 3238 752 3248 784 0 OUTPUT2
port 5 nsew analog default
rlabel metal2 3238 384 3248 416 0 OUTPUT3
port 6 nsew analog default
rlabel metal2 3238 198 3248 230 0 OUTPUT4
port 7 nsew analog default
rlabel metal1 3170 1198 3216 1210 0 VGND
port 1 nsew ground default
rlabel metal1 3170 0 3216 12 0 VGND
port 1 nsew ground default
rlabel metal2 432 984 462 1024 0 INPUT1
port 8 nsew analog default
rlabel metal2 432 790 484 842 0 INPUT2
port 9 nsew analog default
rlabel metal2 420 388 460 422 0 INPUT3
port 10 nsew analog default
rlabel metal2 418 180 474 234 0 INPUT4
port 11 nsew analog default
rlabel metal2 456 1074 480 1110 0 DRAIN1
port 12 nsew
rlabel metal2 456 702 480 738 0 DRAIN2
port 13 nsew
rlabel metal2 456 472 480 508 0 DRAIN3
port 14 nsew
rlabel metal2 456 102 480 138 0 DRAIN4
port 15 nsew
rlabel metal1 1594 1190 1666 1210 0 GATE1
port 16 nsew
rlabel metal1 2398 1182 2478 1210 0 VTUN
port 17 nsew
rlabel metal1 2918 0 2964 12 0 WTAMIDDLENODE
port 18 nsew
rlabel metal1 2918 1198 2964 1210 0 WTAMIDDLENODE
port 18 nsew
rlabel metal1 688 1196 726 1210 0 COLSEL1
port 19 nsew
rlabel metal1 606 1196 638 1210 0 VINJ
port 21 nsew
rlabel metal1 768 1196 800 1210 0 VPWR
port 20 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
