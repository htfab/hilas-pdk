magic
tech sky130A
timestamp 1629137234
<< checkpaint >>
rect -630 1742 4676 2340
rect -630 -10 4679 1742
rect -627 -608 4679 -10
rect 418 -630 4106 -608
<< error_s >>
rect 478 1199 484 1205
rect 583 1199 589 1205
rect 1449 1199 1455 1205
rect 1554 1199 1560 1205
rect 2528 1199 2534 1205
rect 2633 1199 2639 1205
rect 904 1189 910 1195
rect 957 1189 963 1195
rect 1075 1189 1081 1195
rect 1128 1189 1134 1195
rect 2954 1189 2960 1195
rect 3007 1189 3013 1195
rect 472 1135 478 1141
rect 589 1135 595 1141
rect 898 1139 904 1145
rect 963 1139 969 1145
rect 1069 1139 1075 1145
rect 1134 1139 1140 1145
rect 1443 1135 1449 1141
rect 1560 1135 1566 1141
rect 2522 1135 2528 1141
rect 2639 1135 2645 1141
rect 2948 1139 2954 1145
rect 3013 1139 3019 1145
rect 478 1082 484 1088
rect 583 1082 589 1088
rect 904 1080 910 1086
rect 957 1080 963 1086
rect 1075 1080 1081 1086
rect 1128 1080 1134 1086
rect 1449 1082 1455 1088
rect 1554 1082 1560 1088
rect 2528 1082 2534 1088
rect 2633 1082 2639 1088
rect 2954 1080 2960 1086
rect 3007 1080 3013 1086
rect 898 1030 904 1036
rect 963 1030 969 1036
rect 1069 1030 1075 1036
rect 1134 1030 1140 1036
rect 2948 1030 2954 1036
rect 3013 1030 3019 1036
rect 247 1022 260 1027
rect 261 1022 274 1026
rect 247 1019 274 1022
rect 472 1018 478 1024
rect 589 1018 595 1024
rect 1443 1018 1449 1024
rect 1560 1018 1566 1024
rect 1764 1022 1777 1026
rect 1778 1022 1791 1027
rect 1764 1019 1791 1022
rect 2522 1018 2528 1024
rect 2639 1018 2645 1024
rect 478 897 484 903
rect 583 897 589 903
rect 1449 897 1455 903
rect 1554 897 1560 903
rect 2528 897 2534 903
rect 2633 897 2639 903
rect 904 891 910 897
rect 957 891 963 897
rect 1075 891 1081 897
rect 1128 891 1134 897
rect 2954 891 2960 897
rect 3007 891 3013 897
rect 898 841 904 847
rect 963 841 969 847
rect 1069 841 1075 847
rect 1134 841 1140 847
rect 2948 841 2954 847
rect 3013 841 3019 847
rect 472 833 478 839
rect 589 833 595 839
rect 1443 833 1449 839
rect 1560 833 1566 839
rect 2522 833 2528 839
rect 2639 833 2645 839
rect 478 781 484 787
rect 583 781 589 787
rect 1449 781 1455 787
rect 1554 781 1560 787
rect 904 774 910 780
rect 957 774 963 780
rect 1075 774 1081 780
rect 1128 774 1134 780
rect 1989 778 1990 790
rect 2528 781 2534 787
rect 2633 781 2639 787
rect 2003 764 2004 776
rect 2954 774 2960 780
rect 3007 774 3013 780
rect 898 724 904 730
rect 963 724 969 730
rect 1069 724 1075 730
rect 1134 724 1140 730
rect 2948 724 2954 730
rect 3013 724 3019 730
rect 472 717 478 723
rect 589 717 595 723
rect 1443 717 1449 723
rect 1560 717 1566 723
rect 2522 717 2528 723
rect 2639 717 2645 723
rect 152 677 154 685
rect 2202 677 2203 685
rect 65 664 66 672
rect 146 664 147 672
rect 1908 666 1909 672
rect 1908 658 1910 666
rect 1989 664 1990 672
rect 481 601 487 607
rect 586 601 592 607
rect 1452 601 1458 607
rect 1557 601 1563 607
rect 2530 601 2536 607
rect 2635 601 2641 607
rect 907 591 913 597
rect 960 591 966 597
rect 1078 591 1084 597
rect 1131 591 1137 597
rect 2956 591 2962 597
rect 3009 591 3015 597
rect 475 537 481 543
rect 592 537 598 543
rect 901 541 907 547
rect 966 541 972 547
rect 1072 541 1078 547
rect 1137 541 1143 547
rect 1446 537 1452 543
rect 1563 537 1569 543
rect 2524 537 2530 543
rect 2641 537 2647 543
rect 2950 541 2956 547
rect 3015 541 3021 547
rect 481 484 487 490
rect 586 484 592 490
rect 907 482 913 488
rect 960 482 966 488
rect 1078 482 1084 488
rect 1131 482 1137 488
rect 1452 484 1458 490
rect 1557 484 1563 490
rect 2530 484 2536 490
rect 2635 484 2641 490
rect 2956 482 2962 488
rect 3009 482 3015 488
rect 901 432 907 438
rect 966 432 972 438
rect 1072 432 1078 438
rect 1137 432 1143 438
rect 2950 432 2956 438
rect 3015 432 3021 438
rect 250 424 263 429
rect 264 424 277 428
rect 250 421 277 424
rect 475 420 481 426
rect 592 420 598 426
rect 1446 420 1452 426
rect 1563 420 1569 426
rect 1767 424 1780 428
rect 1781 424 1794 429
rect 1767 421 1794 424
rect 2524 420 2530 426
rect 2641 420 2647 426
rect 481 299 487 305
rect 586 299 592 305
rect 1452 299 1458 305
rect 1557 299 1563 305
rect 2530 299 2536 305
rect 2635 299 2641 305
rect 907 293 913 299
rect 960 293 966 299
rect 1078 293 1084 299
rect 1131 293 1137 299
rect 2956 293 2962 299
rect 3009 293 3015 299
rect 901 243 907 249
rect 966 243 972 249
rect 1072 243 1078 249
rect 1137 243 1143 249
rect 2950 243 2956 249
rect 3015 243 3021 249
rect 475 235 481 241
rect 592 235 598 241
rect 1446 235 1452 241
rect 1563 235 1569 241
rect 2524 235 2530 241
rect 2641 235 2647 241
rect 481 183 487 189
rect 586 183 592 189
rect 1452 183 1458 189
rect 1557 183 1563 189
rect 907 176 913 182
rect 960 176 966 182
rect 1078 176 1084 182
rect 1131 176 1137 182
rect 1991 180 1993 192
rect 2530 183 2536 189
rect 2635 183 2641 189
rect 1991 132 1992 180
rect 2005 166 2007 178
rect 2956 176 2962 182
rect 3009 176 3015 182
rect 2005 146 2006 166
rect 901 126 907 132
rect 966 126 972 132
rect 1072 126 1078 132
rect 1137 126 1143 132
rect 2950 126 2956 132
rect 3015 126 3021 132
rect 475 119 481 125
rect 592 119 598 125
rect 1446 119 1452 125
rect 1563 119 1569 125
rect 2524 119 2530 125
rect 2641 119 2647 125
use sky130_hilas_WTA4Stage01  sky130_hilas_WTA4Stage01_1
timestamp 1628285143
transform 1 0 3124 0 1 700
box -2078 -102 350 989
use sky130_hilas_WTA4Stage01  sky130_hilas_WTA4Stage01_0
timestamp 1628285143
transform 1 0 3126 0 1 102
box -2078 -102 350 989
use sky130_hilas_swc4x2cell  sky130_hilas_swc4x2cell_1
timestamp 1629137207
transform 1 0 1017 0 1 661
box -1017 -41 3029 1049
use sky130_hilas_swc4x2cell  sky130_hilas_swc4x2cell_0
timestamp 1629137207
transform 1 0 1020 0 1 63
box -1017 -41 3029 1049
<< end >>
