VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_hilas_TA2Cell_1FG_Strong
  CLASS CORE ;
  FOREIGN sky130_hilas_TA2Cell_1FG_Strong ;
  ORIGIN 0.000 0.000 ;
  SIZE 46.940 BY 23.320 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 25.760 14.880 26.180 15.030 ;
        RECT 26.790 14.880 27.210 15.030 ;
        RECT 25.760 14.740 27.210 14.880 ;
    END
  END VTUN
  PIN PROG
    PORT
      LAYER met1 ;
        RECT 18.520 14.970 18.730 15.030 ;
    END
  END PROG
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT 30.490 14.950 30.720 15.030 ;
    END
  END GATE1
  PIN VIN11
    PORT
      LAYER met1 ;
        RECT 17.640 14.920 17.850 15.030 ;
    END
  END VIN11
  PIN VINJ
    PORT
      LAYER met2 ;
        RECT 15.200 14.890 15.520 15.010 ;
        RECT 37.470 14.890 37.790 15.010 ;
        RECT 15.200 14.710 37.790 14.890 ;
    END
    PORT
      LAYER met1 ;
        RECT 37.450 15.010 37.730 15.030 ;
        RECT 37.450 14.950 37.790 15.010 ;
        RECT 37.470 14.710 37.790 14.950 ;
      LAYER via ;
        RECT 37.500 14.730 37.760 14.990 ;
    END
    PORT
      LAYER met1 ;
        RECT 37.450 8.980 37.730 9.030 ;
    END
  END VINJ
  PIN VIN22
    PORT
      LAYER met2 ;
        RECT 38.570 14.760 38.880 15.000 ;
    END
  END VIN22
  PIN VIN21
    PORT
      LAYER met2 ;
        RECT 38.650 12.090 38.970 12.330 ;
    END
  END VIN21
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 41.800 14.880 42.080 15.030 ;
    END
    PORT
      LAYER met1 ;
        RECT 41.810 8.980 42.080 9.190 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 41.570 16.460 41.890 16.540 ;
        RECT 40.580 16.280 41.890 16.460 ;
        RECT 40.580 16.110 41.760 16.280 ;
        RECT 40.630 15.960 40.950 16.110 ;
    END
    PORT
      LAYER met2 ;
        RECT 39.610 9.330 39.930 9.480 ;
        RECT 23.420 9.180 39.930 9.330 ;
        RECT 23.420 9.030 23.740 9.180 ;
        RECT 29.220 9.030 29.540 9.180 ;
    END
  END VGND
  PIN OUTPUT2
    PORT
      LAYER met2 ;
        RECT 42.990 11.500 43.100 11.720 ;
    END
  END OUTPUT2
  PIN OUTPUT1
    PORT
      LAYER met2 ;
        RECT 42.990 12.320 43.100 12.550 ;
    END
  END OUTPUT1
  PIN GATESEL1
    PORT
      LAYER met1 ;
        RECT 15.520 15.030 15.940 19.320 ;
        RECT 15.360 15.010 15.960 15.030 ;
        RECT 15.200 14.970 15.960 15.010 ;
        RECT 15.200 14.710 15.940 14.970 ;
        RECT 15.520 13.270 15.940 14.710 ;
      LAYER via ;
        RECT 15.230 14.730 15.490 14.990 ;
    END
  END GATESEL1
  PIN GATESEL2
    PORT
      LAYER met1 ;
        RECT 37.010 8.980 37.200 9.030 ;
    END
    PORT
      LAYER met1 ;
        RECT 37.010 14.950 37.200 15.030 ;
    END
  END GATESEL2
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 15.000 14.350 15.080 14.530 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 15.000 9.480 15.080 9.660 ;
    END
  END DRAIN2
  PIN VIN12
    PORT
      LAYER met1 ;
        RECT 17.650 8.990 17.880 9.110 ;
    END
  END VIN12
  PIN GATE2
    PORT
      LAYER met1 ;
        RECT 18.110 14.950 18.300 15.030 ;
    END
  END GATE2
  PIN RUN
    PORT
      LAYER met1 ;
        RECT 19.600 14.960 19.780 15.030 ;
    END
  END RUN
  OBS
      LAYER nwell ;
        RECT 0.040 22.980 1.770 23.320 ;
        RECT 44.920 22.980 46.650 23.320 ;
        RECT 0.040 21.420 1.790 22.980 ;
        RECT 0.060 19.790 1.790 21.420 ;
        RECT 44.900 21.420 46.650 22.980 ;
        RECT 44.900 19.790 46.630 21.420 ;
        RECT 0.000 16.620 3.310 19.790 ;
        RECT 43.390 19.400 46.690 19.790 ;
        RECT 19.850 19.360 22.560 19.400 ;
        RECT 43.390 19.360 46.930 19.400 ;
        RECT 19.850 17.710 22.570 19.360 ;
        RECT 38.630 19.310 41.930 19.320 ;
        RECT 40.970 19.280 41.160 19.310 ;
        RECT 43.390 17.710 46.940 19.360 ;
        RECT 0.000 12.800 3.310 15.970 ;
        RECT 15.140 15.030 15.700 17.090 ;
        RECT 15.000 15.020 18.310 15.030 ;
        RECT 15.140 14.670 15.700 15.020 ;
        RECT 15.520 13.280 15.940 13.350 ;
        RECT 19.850 13.130 22.570 14.780 ;
        RECT 30.990 14.670 31.550 17.090 ;
        RECT 43.390 16.620 46.690 17.710 ;
        RECT 43.800 15.970 45.080 16.620 ;
        RECT 37.970 15.020 39.310 15.030 ;
        RECT 37.470 14.710 37.790 15.010 ;
        RECT 41.820 14.850 43.100 15.030 ;
        RECT 43.390 14.780 46.690 15.970 ;
        RECT 43.390 13.130 46.940 14.780 ;
        RECT 19.850 13.090 22.560 13.130 ;
        RECT 43.390 13.090 46.930 13.130 ;
        RECT 43.390 12.800 46.690 13.090 ;
        RECT 43.800 9.470 45.080 12.310 ;
        RECT 41.820 8.980 43.100 9.170 ;
        RECT 37.970 7.550 38.420 7.780 ;
        RECT 36.630 7.420 38.490 7.490 ;
        RECT 40.260 3.050 42.120 6.040 ;
        RECT 40.260 0.000 42.120 2.990 ;
      LAYER li1 ;
        RECT 0.820 21.590 1.370 22.020 ;
        RECT 45.320 21.590 45.870 22.020 ;
        RECT 0.820 19.860 1.370 20.290 ;
        RECT 45.320 19.860 45.870 20.290 ;
        RECT 0.400 19.060 0.600 19.410 ;
        RECT 1.880 19.160 2.410 19.330 ;
        RECT 44.280 19.160 44.810 19.330 ;
        RECT 0.390 19.030 0.600 19.060 ;
        RECT 46.090 19.060 46.290 19.410 ;
        RECT 46.090 19.030 46.300 19.060 ;
        RECT 0.390 18.450 0.610 19.030 ;
        RECT 0.390 18.440 0.600 18.450 ;
        RECT 0.770 18.270 0.960 18.280 ;
        RECT 0.760 17.980 0.960 18.270 ;
        RECT 0.700 17.650 0.970 17.980 ;
        RECT 1.160 17.170 1.330 18.780 ;
        RECT 7.310 18.770 7.500 19.000 ;
        RECT 1.150 16.980 1.330 17.170 ;
        RECT 1.990 17.080 2.160 18.770 ;
        RECT 2.580 18.580 2.910 18.750 ;
        RECT 3.930 18.580 4.280 18.750 ;
        RECT 7.590 18.720 8.470 18.890 ;
        RECT 7.780 18.330 7.970 18.440 ;
        RECT 7.670 18.210 7.970 18.330 ;
        RECT 8.300 18.330 8.470 18.720 ;
        RECT 7.670 18.160 7.890 18.210 ;
        RECT 8.300 18.160 8.690 18.330 ;
        RECT 20.150 18.230 20.380 18.920 ;
        RECT 44.520 18.230 44.750 18.920 ;
        RECT 2.580 17.790 2.910 17.960 ;
        RECT 3.930 17.790 4.280 17.960 ;
        RECT 39.750 17.940 40.070 17.980 ;
        RECT 39.750 17.750 40.080 17.940 ;
        RECT 39.750 17.720 40.070 17.750 ;
        RECT 6.380 17.370 6.700 17.410 ;
        RECT 7.630 17.370 8.710 17.540 ;
        RECT 9.040 17.370 10.120 17.540 ;
        RECT 6.370 17.180 6.700 17.370 ;
        RECT 2.580 17.000 2.910 17.170 ;
        RECT 3.930 17.000 4.270 17.170 ;
        RECT 6.380 17.150 6.700 17.180 ;
        RECT 44.530 17.080 44.700 18.230 ;
        RECT 45.360 17.170 45.530 18.780 ;
        RECT 46.080 18.450 46.300 19.030 ;
        RECT 46.090 18.440 46.300 18.450 ;
        RECT 45.730 18.270 45.920 18.280 ;
        RECT 45.730 17.980 45.930 18.270 ;
        RECT 45.720 17.650 46.010 17.980 ;
        RECT 7.310 16.780 7.500 17.010 ;
        RECT 45.360 16.980 45.540 17.170 ;
        RECT 7.610 16.580 7.690 16.750 ;
        RECT 8.170 16.430 8.380 16.860 ;
        RECT 8.190 16.410 8.360 16.430 ;
        RECT 6.370 15.680 6.690 15.720 ;
        RECT 7.320 15.710 7.510 15.940 ;
        RECT 7.640 15.840 7.690 16.010 ;
        RECT 7.780 15.890 7.970 16.120 ;
        RECT 8.780 16.010 8.950 16.580 ;
        RECT 13.060 16.430 13.250 16.750 ;
        RECT 33.440 16.430 33.630 16.750 ;
        RECT 13.060 16.340 13.340 16.430 ;
        RECT 9.700 16.200 13.340 16.340 ;
        RECT 33.350 16.340 33.630 16.430 ;
        RECT 44.360 16.540 44.690 16.710 ;
        RECT 44.800 16.630 45.130 16.800 ;
        RECT 33.350 16.200 36.990 16.340 ;
        RECT 44.360 16.260 44.720 16.540 ;
        RECT 9.700 16.160 13.250 16.200 ;
        RECT 8.060 15.980 8.110 15.990 ;
        RECT 8.690 15.980 8.770 15.990 ;
        RECT 8.060 15.940 8.770 15.980 ;
        RECT 8.060 15.900 8.790 15.940 ;
        RECT 8.020 15.780 8.860 15.900 ;
        RECT 13.060 15.740 13.250 16.160 ;
        RECT 33.440 16.160 36.990 16.200 ;
        RECT 33.440 15.740 33.630 16.160 ;
        RECT 42.290 16.010 42.610 16.050 ;
        RECT 42.290 15.820 42.620 16.010 ;
        RECT 42.290 15.790 42.610 15.820 ;
        RECT 42.690 15.800 42.890 16.130 ;
        RECT 43.280 15.940 43.480 16.130 ;
        RECT 44.010 16.090 44.720 16.260 ;
        RECT 43.950 15.970 44.270 16.010 ;
        RECT 1.150 15.420 1.330 15.610 ;
        RECT 0.700 14.610 0.970 14.940 ;
        RECT 0.760 14.320 0.960 14.610 ;
        RECT 0.770 14.310 0.960 14.320 ;
        RECT 0.390 14.140 0.600 14.150 ;
        RECT 0.390 13.560 0.610 14.140 ;
        RECT 1.160 13.810 1.330 15.420 ;
        RECT 1.990 13.820 2.160 15.510 ;
        RECT 2.580 15.420 2.910 15.590 ;
        RECT 3.930 15.420 4.270 15.590 ;
        RECT 6.360 15.490 6.690 15.680 ;
        RECT 6.370 15.460 6.690 15.490 ;
        RECT 42.970 15.610 43.160 15.620 ;
        RECT 43.170 15.610 43.520 15.940 ;
        RECT 43.950 15.780 44.280 15.970 ;
        RECT 43.950 15.750 44.270 15.780 ;
        RECT 7.630 15.050 8.710 15.220 ;
        RECT 9.030 15.050 10.270 15.220 ;
        RECT 39.750 15.180 40.070 15.220 ;
        RECT 34.470 15.120 34.700 15.160 ;
        RECT 39.750 14.990 40.080 15.180 ;
        RECT 42.060 15.100 42.230 15.430 ;
        RECT 42.240 15.360 42.560 15.400 ;
        RECT 42.240 15.170 42.570 15.360 ;
        RECT 42.240 15.140 42.560 15.170 ;
        RECT 42.690 15.140 42.890 15.470 ;
        RECT 42.970 15.280 43.520 15.610 ;
        RECT 39.750 14.960 40.070 14.990 ;
        RECT 43.170 14.950 43.520 15.280 ;
        RECT 2.580 14.630 2.910 14.800 ;
        RECT 3.930 14.630 4.280 14.800 ;
        RECT 9.360 14.730 9.530 14.790 ;
        RECT 44.010 14.770 44.710 15.650 ;
        RECT 45.360 15.420 45.540 15.610 ;
        RECT 7.770 14.430 7.960 14.540 ;
        RECT 9.340 14.520 9.550 14.730 ;
        RECT 9.360 14.450 9.530 14.520 ;
        RECT 7.670 14.310 7.960 14.430 ;
        RECT 8.230 14.420 8.690 14.430 ;
        RECT 7.670 14.260 7.880 14.310 ;
        RECT 8.230 14.270 8.700 14.420 ;
        RECT 43.350 14.380 43.540 14.610 ;
        RECT 44.530 14.350 44.700 14.770 ;
        RECT 8.230 14.260 8.690 14.270 ;
        RECT 2.580 13.840 2.910 14.010 ;
        RECT 3.930 13.840 4.280 14.010 ;
        RECT 7.340 13.920 7.530 14.030 ;
        RECT 8.230 13.920 8.420 14.260 ;
        RECT 7.340 13.800 8.420 13.920 ;
        RECT 7.460 13.740 8.420 13.800 ;
        RECT 20.150 13.570 20.380 14.260 ;
        RECT 42.060 13.840 42.230 14.170 ;
        RECT 42.240 14.100 42.560 14.130 ;
        RECT 42.240 13.910 42.570 14.100 ;
        RECT 42.240 13.870 42.560 13.910 ;
        RECT 42.690 13.800 42.890 14.130 ;
        RECT 43.170 13.990 43.520 14.320 ;
        RECT 44.000 14.260 44.700 14.350 ;
        RECT 44.000 14.170 44.750 14.260 ;
        RECT 42.970 13.660 43.520 13.990 ;
        RECT 42.970 13.650 43.160 13.660 ;
        RECT 0.390 13.530 0.600 13.560 ;
        RECT 0.400 13.180 0.600 13.530 ;
        RECT 42.290 13.450 42.610 13.480 ;
        RECT 1.880 13.260 2.410 13.430 ;
        RECT 42.290 13.260 42.620 13.450 ;
        RECT 42.290 13.220 42.610 13.260 ;
        RECT 42.690 13.140 42.890 13.470 ;
        RECT 43.170 13.330 43.520 13.660 ;
        RECT 44.000 13.750 44.320 13.790 ;
        RECT 44.000 13.560 44.330 13.750 ;
        RECT 44.520 13.570 44.750 14.170 ;
        RECT 45.360 13.810 45.530 15.420 ;
        RECT 45.720 14.610 46.010 14.940 ;
        RECT 45.730 14.320 45.930 14.610 ;
        RECT 45.730 14.310 45.920 14.320 ;
        RECT 46.090 14.140 46.300 14.150 ;
        RECT 46.080 13.560 46.300 14.140 ;
        RECT 44.000 13.530 44.320 13.560 ;
        RECT 46.090 13.530 46.300 13.560 ;
        RECT 43.280 13.140 43.480 13.330 ;
        RECT 44.280 13.260 44.810 13.430 ;
        RECT 46.090 13.180 46.290 13.530 ;
        RECT 42.290 13.010 42.610 13.050 ;
        RECT 42.290 12.820 42.620 13.010 ;
        RECT 42.290 12.790 42.610 12.820 ;
        RECT 42.690 12.800 42.890 13.130 ;
        RECT 43.280 12.940 43.480 13.130 ;
        RECT 43.990 13.030 44.310 13.070 ;
        RECT 42.970 12.610 43.160 12.620 ;
        RECT 43.170 12.610 43.520 12.940 ;
        RECT 43.990 12.840 44.320 13.030 ;
        RECT 43.990 12.810 44.310 12.840 ;
        RECT 42.060 12.100 42.230 12.430 ;
        RECT 42.240 12.360 42.560 12.400 ;
        RECT 42.240 12.170 42.570 12.360 ;
        RECT 42.240 12.140 42.560 12.170 ;
        RECT 42.690 12.140 42.890 12.470 ;
        RECT 42.970 12.280 43.520 12.610 ;
        RECT 43.170 12.020 43.520 12.280 ;
        RECT 43.170 11.950 43.540 12.020 ;
        RECT 43.350 11.790 43.540 11.950 ;
        RECT 44.000 11.890 44.700 12.070 ;
        RECT 42.060 10.840 42.230 11.170 ;
        RECT 42.240 11.100 42.560 11.130 ;
        RECT 42.240 10.910 42.570 11.100 ;
        RECT 42.240 10.870 42.560 10.910 ;
        RECT 42.690 10.800 42.890 11.130 ;
        RECT 43.170 10.990 43.520 11.320 ;
        RECT 42.970 10.660 43.520 10.990 ;
        RECT 44.010 10.820 44.710 11.470 ;
        RECT 42.970 10.650 43.160 10.660 ;
        RECT 37.720 10.550 38.040 10.590 ;
        RECT 37.710 10.360 38.040 10.550 ;
        RECT 37.720 10.350 38.040 10.360 ;
        RECT 37.710 10.330 38.040 10.350 ;
        RECT 42.290 10.450 42.610 10.480 ;
        RECT 37.710 10.020 37.880 10.330 ;
        RECT 42.290 10.260 42.620 10.450 ;
        RECT 42.290 10.220 42.610 10.260 ;
        RECT 42.690 10.140 42.890 10.470 ;
        RECT 43.170 10.330 43.520 10.660 ;
        RECT 43.910 10.590 44.710 10.820 ;
        RECT 43.910 10.560 44.230 10.590 ;
        RECT 43.280 10.140 43.480 10.330 ;
        RECT 44.010 9.980 44.720 10.150 ;
        RECT 37.870 9.720 38.190 9.760 ;
        RECT 37.860 9.530 38.190 9.720 ;
        RECT 44.360 9.700 44.720 9.980 ;
        RECT 44.360 9.530 44.690 9.700 ;
        RECT 37.870 9.500 38.190 9.530 ;
        RECT 44.800 9.440 45.130 9.610 ;
        RECT 37.060 8.900 37.380 8.930 ;
        RECT 37.060 8.710 37.390 8.900 ;
        RECT 37.060 8.670 37.380 8.710 ;
        RECT 37.040 6.950 37.220 8.010 ;
        RECT 37.790 7.620 38.110 7.650 ;
        RECT 37.790 7.550 38.120 7.620 ;
        RECT 37.650 7.430 38.120 7.550 ;
        RECT 37.650 7.420 38.110 7.430 ;
        RECT 37.770 7.390 38.110 7.420 ;
        RECT 37.770 7.320 37.820 7.390 ;
        RECT 37.690 6.990 37.860 7.320 ;
        RECT 38.090 6.790 38.170 6.870 ;
        RECT 38.230 6.790 38.420 6.910 ;
        RECT 38.090 6.700 38.420 6.790 ;
        RECT 38.230 6.680 38.420 6.700 ;
        RECT 40.670 3.520 40.850 5.570 ;
        RECT 41.400 5.310 41.730 5.480 ;
        RECT 41.480 3.530 41.650 5.310 ;
        RECT 40.670 0.470 40.850 2.520 ;
        RECT 41.400 2.260 41.730 2.430 ;
        RECT 41.480 0.480 41.650 2.260 ;
      LAYER mcon ;
        RECT 1.100 21.670 1.370 21.940 ;
        RECT 45.320 21.670 45.590 21.940 ;
        RECT 1.100 19.940 1.370 20.210 ;
        RECT 45.320 19.940 45.590 20.210 ;
        RECT 2.230 19.160 2.410 19.330 ;
        RECT 0.420 18.860 0.590 19.030 ;
        RECT 7.320 18.800 7.490 18.970 ;
        RECT 0.770 18.020 0.950 18.210 ;
        RECT 7.790 18.240 7.960 18.410 ;
        RECT 20.180 18.710 20.350 18.880 ;
        RECT 20.180 18.260 20.350 18.430 ;
        RECT 44.550 18.710 44.720 18.880 ;
        RECT 46.100 18.860 46.270 19.030 ;
        RECT 44.550 18.260 44.720 18.430 ;
        RECT 39.810 17.760 39.980 17.930 ;
        RECT 6.470 17.190 6.640 17.360 ;
        RECT 45.740 18.020 45.920 18.210 ;
        RECT 7.320 16.810 7.490 16.980 ;
        RECT 7.330 15.740 7.500 15.910 ;
        RECT 7.790 15.920 7.960 16.090 ;
        RECT 13.160 16.230 13.330 16.400 ;
        RECT 33.360 16.230 33.530 16.400 ;
        RECT 42.350 15.830 42.520 16.000 ;
        RECT 0.770 14.380 0.950 14.570 ;
        RECT 6.460 15.500 6.630 15.670 ;
        RECT 44.010 15.790 44.180 15.960 ;
        RECT 39.810 15.000 39.980 15.170 ;
        RECT 42.300 15.180 42.470 15.350 ;
        RECT 43.290 15.440 43.460 15.610 ;
        RECT 7.780 14.340 7.950 14.510 ;
        RECT 43.360 14.410 43.530 14.580 ;
        RECT 7.350 13.830 7.520 14.000 ;
        RECT 20.180 14.060 20.350 14.230 ;
        RECT 42.300 13.920 42.470 14.090 ;
        RECT 0.420 13.560 0.590 13.730 ;
        RECT 20.180 13.610 20.350 13.780 ;
        RECT 43.290 13.660 43.460 13.830 ;
        RECT 44.550 14.060 44.720 14.230 ;
        RECT 2.230 13.260 2.410 13.430 ;
        RECT 42.350 13.270 42.520 13.440 ;
        RECT 45.740 14.380 45.920 14.570 ;
        RECT 44.060 13.570 44.230 13.740 ;
        RECT 44.550 13.610 44.720 13.780 ;
        RECT 46.100 13.560 46.270 13.730 ;
        RECT 42.350 12.830 42.520 13.000 ;
        RECT 44.050 12.850 44.220 13.020 ;
        RECT 42.300 12.180 42.470 12.350 ;
        RECT 43.290 12.440 43.460 12.610 ;
        RECT 43.360 11.820 43.530 11.990 ;
        RECT 42.300 10.920 42.470 11.090 ;
        RECT 43.290 10.660 43.460 10.830 ;
        RECT 37.810 10.370 37.980 10.540 ;
        RECT 42.350 10.270 42.520 10.440 ;
        RECT 43.970 10.600 44.140 10.770 ;
        RECT 37.960 9.540 38.130 9.710 ;
        RECT 37.120 8.720 37.290 8.890 ;
        RECT 37.850 7.440 38.020 7.610 ;
        RECT 38.240 6.710 38.410 6.880 ;
      LAYER met1 ;
        RECT 0.360 19.090 0.520 19.730 ;
        RECT 0.360 18.540 0.630 19.090 ;
        RECT 0.350 18.490 0.630 18.540 ;
        RECT 0.350 18.400 0.520 18.490 ;
        RECT 0.360 16.710 0.520 18.400 ;
        RECT 0.770 18.280 0.960 19.730 ;
        RECT 1.040 19.400 1.430 22.990 ;
        RECT 45.260 19.400 45.650 22.990 ;
        RECT 2.170 18.920 2.480 19.360 ;
        RECT 5.120 19.270 5.280 19.320 ;
        RECT 5.530 19.260 5.720 19.320 ;
        RECT 7.400 19.030 7.610 19.320 ;
        RECT 7.290 18.740 7.610 19.030 ;
        RECT 0.740 18.250 0.960 18.280 ;
        RECT 0.730 17.980 0.980 18.250 ;
        RECT 0.730 17.970 0.970 17.980 ;
        RECT 0.740 17.730 0.970 17.970 ;
        RECT 0.770 16.710 0.930 17.730 ;
        RECT 1.120 16.920 1.360 17.300 ;
        RECT 6.390 17.120 6.710 17.440 ;
        RECT 7.400 17.040 7.610 18.740 ;
        RECT 7.870 18.470 8.060 19.320 ;
        RECT 7.760 18.180 8.060 18.470 ;
        RECT 7.290 16.750 7.610 17.040 ;
        RECT 5.760 16.500 6.020 16.560 ;
        RECT 7.400 16.530 7.610 16.750 ;
        RECT 5.760 16.240 6.120 16.500 ;
        RECT 5.880 16.080 6.120 16.240 ;
        RECT 7.870 16.150 8.060 18.180 ;
        RECT 8.280 16.860 8.490 19.320 ;
        RECT 8.160 16.350 8.490 16.860 ;
        RECT 7.420 15.970 7.610 16.020 ;
        RECT 0.360 14.190 0.520 15.880 ;
        RECT 0.770 14.860 0.930 15.880 ;
        RECT 1.120 15.290 1.360 15.670 ;
        RECT 6.380 15.430 6.700 15.750 ;
        RECT 7.300 15.680 7.610 15.970 ;
        RECT 7.760 15.860 8.060 16.150 ;
        RECT 0.740 14.620 0.970 14.860 ;
        RECT 0.730 14.610 0.970 14.620 ;
        RECT 0.730 14.340 0.980 14.610 ;
        RECT 0.740 14.310 0.960 14.340 ;
        RECT 0.350 14.100 0.520 14.190 ;
        RECT 0.350 14.050 0.630 14.100 ;
        RECT 0.360 13.500 0.630 14.050 ;
        RECT 0.360 12.860 0.520 13.500 ;
        RECT 0.770 12.860 0.960 14.310 ;
        RECT 7.420 14.060 7.610 15.680 ;
        RECT 7.870 14.570 8.060 15.860 ;
        RECT 7.750 14.280 8.060 14.570 ;
        RECT 7.100 13.770 7.110 13.780 ;
        RECT 7.320 13.770 7.610 14.060 ;
        RECT 2.170 13.230 2.480 13.670 ;
        RECT 5.120 13.270 5.280 13.320 ;
        RECT 5.530 13.270 5.720 13.320 ;
        RECT 7.410 13.270 7.640 13.770 ;
        RECT 7.870 13.270 8.060 14.280 ;
        RECT 8.280 13.270 8.490 16.350 ;
        RECT 9.360 14.790 9.540 19.320 ;
        RECT 13.230 16.460 13.460 19.320 ;
        RECT 20.130 18.180 20.390 18.970 ;
        RECT 13.130 16.170 13.460 16.460 ;
        RECT 9.300 14.450 9.590 14.790 ;
        RECT 9.360 13.270 9.540 14.450 ;
        RECT 13.230 13.270 13.460 16.170 ;
        RECT 20.130 13.520 20.390 14.310 ;
        RECT 30.750 13.270 31.170 19.320 ;
        RECT 33.230 16.460 33.460 19.320 ;
        RECT 33.230 16.170 33.560 16.460 ;
        RECT 33.230 13.270 33.460 16.170 ;
        RECT 34.450 13.270 34.680 19.320 ;
        RECT 40.970 19.280 41.160 19.320 ;
        RECT 39.740 17.690 40.060 18.010 ;
        RECT 40.660 16.530 40.920 16.850 ;
        RECT 41.410 16.570 41.690 19.320 ;
        RECT 44.210 18.970 44.520 19.360 ;
        RECT 44.210 18.920 44.760 18.970 ;
        RECT 44.500 18.180 44.760 18.920 ;
        RECT 45.730 18.280 45.920 19.730 ;
        RECT 46.170 19.090 46.330 19.730 ;
        RECT 46.060 18.540 46.330 19.090 ;
        RECT 46.060 18.490 46.340 18.540 ;
        RECT 46.170 18.400 46.340 18.490 ;
        RECT 45.730 18.250 45.950 18.280 ;
        RECT 45.710 17.980 45.960 18.250 ;
        RECT 45.720 17.970 45.960 17.980 ;
        RECT 45.720 17.730 45.950 17.970 ;
        RECT 45.330 16.920 45.570 17.300 ;
        RECT 45.760 16.710 45.920 17.730 ;
        RECT 46.170 16.710 46.330 18.400 ;
        RECT 41.410 16.250 41.860 16.570 ;
        RECT 40.660 15.930 40.920 16.250 ;
        RECT 39.740 14.930 40.060 15.250 ;
        RECT 41.410 15.030 41.690 16.250 ;
        RECT 42.280 16.000 42.600 16.080 ;
        RECT 42.280 15.760 42.850 16.000 ;
        RECT 42.510 15.430 42.850 15.760 ;
        RECT 42.230 15.110 42.850 15.430 ;
        RECT 41.140 14.890 41.690 15.030 ;
        RECT 40.970 13.270 41.160 13.320 ;
        RECT 41.410 13.270 41.690 14.890 ;
        RECT 42.510 14.160 42.850 15.110 ;
        RECT 42.230 13.840 42.850 14.160 ;
        RECT 42.510 13.510 42.850 13.840 ;
        RECT 42.280 13.190 42.850 13.510 ;
        RECT 42.510 13.080 42.850 13.190 ;
        RECT 42.280 12.760 42.850 13.080 ;
        RECT 42.510 12.430 42.850 12.760 ;
        RECT 42.230 12.110 42.850 12.430 ;
        RECT 42.510 11.160 42.850 12.110 ;
        RECT 42.230 10.840 42.850 11.160 ;
        RECT 37.730 10.300 38.050 10.620 ;
        RECT 42.510 10.510 42.850 10.840 ;
        RECT 42.280 10.280 42.850 10.510 ;
        RECT 43.180 15.670 43.450 15.990 ;
        RECT 43.940 15.720 44.260 16.040 ;
        RECT 43.180 15.380 43.490 15.670 ;
        RECT 43.180 14.640 43.450 15.380 ;
        RECT 45.330 15.290 45.570 15.670 ;
        RECT 45.760 14.860 45.920 15.880 ;
        RECT 43.180 14.350 43.560 14.640 ;
        RECT 45.720 14.620 45.950 14.860 ;
        RECT 45.720 14.610 45.960 14.620 ;
        RECT 43.180 13.890 43.450 14.350 ;
        RECT 45.710 14.340 45.960 14.610 ;
        RECT 45.730 14.310 45.950 14.340 ;
        RECT 43.180 13.600 43.490 13.890 ;
        RECT 43.990 13.670 44.310 13.820 ;
        RECT 44.500 13.670 44.760 14.310 ;
        RECT 43.180 12.670 43.450 13.600 ;
        RECT 43.990 13.520 44.760 13.670 ;
        RECT 43.990 13.500 44.520 13.520 ;
        RECT 44.210 13.230 44.520 13.500 ;
        RECT 43.980 12.780 44.300 13.100 ;
        RECT 45.730 12.860 45.920 14.310 ;
        RECT 46.170 14.190 46.330 15.880 ;
        RECT 46.170 14.100 46.340 14.190 ;
        RECT 46.060 14.050 46.340 14.100 ;
        RECT 46.060 13.500 46.330 14.050 ;
        RECT 46.170 12.860 46.330 13.500 ;
        RECT 43.180 12.380 43.490 12.670 ;
        RECT 43.180 12.050 43.450 12.380 ;
        RECT 43.180 11.760 43.560 12.050 ;
        RECT 43.180 10.890 43.450 11.760 ;
        RECT 43.180 10.600 43.490 10.890 ;
        RECT 43.180 10.290 43.450 10.600 ;
        RECT 43.900 10.530 44.220 10.850 ;
        RECT 42.280 10.190 42.600 10.280 ;
        RECT 37.880 9.470 38.200 9.790 ;
        RECT 23.420 9.030 23.740 9.330 ;
        RECT 29.220 9.030 29.540 9.330 ;
        RECT 39.610 9.180 39.930 9.480 ;
        RECT 39.610 9.150 40.040 9.180 ;
        RECT 40.640 9.170 41.150 9.180 ;
        RECT 40.640 9.150 41.480 9.170 ;
        RECT 39.610 9.120 41.480 9.150 ;
        RECT 39.760 9.070 41.480 9.120 ;
        RECT 39.790 9.040 41.480 9.070 ;
        RECT 39.820 9.020 41.480 9.040 ;
        RECT 39.890 9.010 40.850 9.020 ;
        RECT 41.140 8.980 41.480 9.020 ;
        RECT 37.050 8.640 37.370 8.960 ;
        RECT 38.130 8.530 38.340 8.740 ;
        RECT 38.130 8.210 38.460 8.530 ;
        RECT 37.780 7.360 38.100 7.680 ;
        RECT 38.130 6.970 38.340 8.210 ;
        RECT 38.210 6.650 38.440 6.940 ;
      LAYER via ;
        RECT 2.190 18.950 2.450 19.210 ;
        RECT 6.420 17.150 6.680 17.410 ;
        RECT 5.760 16.270 6.020 16.530 ;
        RECT 6.410 15.460 6.670 15.720 ;
        RECT 2.190 13.380 2.450 13.640 ;
        RECT 39.770 17.720 40.030 17.980 ;
        RECT 40.660 16.560 40.920 16.820 ;
        RECT 44.240 18.950 44.500 19.210 ;
        RECT 41.600 16.280 41.860 16.540 ;
        RECT 40.660 15.960 40.920 16.220 ;
        RECT 39.770 14.960 40.030 15.220 ;
        RECT 42.310 15.790 42.570 16.050 ;
        RECT 42.260 15.140 42.520 15.400 ;
        RECT 42.260 13.870 42.520 14.130 ;
        RECT 42.310 13.220 42.570 13.480 ;
        RECT 42.310 12.790 42.570 13.050 ;
        RECT 42.260 12.140 42.520 12.400 ;
        RECT 42.260 10.870 42.520 11.130 ;
        RECT 37.760 10.330 38.020 10.590 ;
        RECT 42.310 10.220 42.570 10.480 ;
        RECT 43.970 15.750 44.230 16.010 ;
        RECT 44.020 13.640 44.280 13.790 ;
        RECT 44.020 13.530 44.500 13.640 ;
        RECT 44.240 13.380 44.500 13.530 ;
        RECT 44.010 12.810 44.270 13.070 ;
        RECT 43.930 10.560 44.190 10.820 ;
        RECT 37.910 9.500 38.170 9.760 ;
        RECT 23.450 9.050 23.710 9.310 ;
        RECT 29.250 9.050 29.510 9.310 ;
        RECT 39.640 9.200 39.900 9.460 ;
        RECT 37.080 8.670 37.340 8.930 ;
        RECT 38.200 8.240 38.460 8.500 ;
        RECT 37.810 7.390 38.070 7.650 ;
      LAYER met2 ;
        RECT 2.170 19.240 2.480 19.250 ;
        RECT 0.000 19.060 2.480 19.240 ;
        RECT 2.170 18.920 2.480 19.060 ;
        RECT 44.210 19.240 44.520 19.250 ;
        RECT 44.210 19.060 46.690 19.240 ;
        RECT 44.210 18.920 44.520 19.060 ;
        RECT 7.170 18.820 7.490 18.840 ;
        RECT 4.760 18.640 4.840 18.820 ;
        RECT 7.170 18.640 16.280 18.820 ;
        RECT 30.400 18.640 39.520 18.820 ;
        RECT 39.740 17.800 40.050 18.020 ;
        RECT 39.740 17.690 41.930 17.800 ;
        RECT 39.900 17.580 41.930 17.690 ;
        RECT 6.400 17.280 6.710 17.450 ;
        RECT 6.400 17.120 16.280 17.280 ;
        RECT 6.570 17.090 16.280 17.120 ;
        RECT 40.630 16.560 40.950 16.820 ;
        RECT 5.730 16.270 6.050 16.530 ;
        RECT 6.120 16.360 16.280 16.400 ;
        RECT 6.110 16.170 16.280 16.360 ;
        RECT 42.280 15.800 42.590 16.090 ;
        RECT 43.940 15.800 44.250 16.050 ;
        RECT 6.390 15.430 6.700 15.760 ;
        RECT 41.560 15.720 44.250 15.800 ;
        RECT 41.560 15.570 44.100 15.720 ;
        RECT 6.560 15.230 16.280 15.420 ;
        RECT 39.740 15.040 40.050 15.260 ;
        RECT 41.790 15.040 42.120 15.210 ;
        RECT 42.230 15.110 42.540 15.440 ;
        RECT 39.740 15.000 42.120 15.040 ;
        RECT 39.740 14.930 41.930 15.000 ;
        RECT 39.890 14.830 41.930 14.930 ;
        RECT 39.680 14.130 39.900 14.150 ;
        RECT 4.760 13.770 4.840 13.950 ;
        RECT 7.070 13.940 7.230 13.960 ;
        RECT 39.460 13.940 39.620 13.960 ;
        RECT 7.070 13.890 16.280 13.940 ;
        RECT 7.190 13.790 16.280 13.890 ;
        RECT 30.400 13.890 39.620 13.940 ;
        RECT 30.400 13.790 39.500 13.890 ;
        RECT 39.630 13.790 39.900 14.130 ;
        RECT 41.790 14.060 42.120 14.270 ;
        RECT 42.230 13.830 42.540 14.160 ;
        RECT 43.990 13.670 44.300 13.830 ;
        RECT 2.170 13.530 2.480 13.670 ;
        RECT 43.990 13.660 44.520 13.670 ;
        RECT 0.000 13.350 2.480 13.530 ;
        RECT 41.820 13.530 44.520 13.660 ;
        RECT 2.170 13.340 2.480 13.350 ;
        RECT 37.890 13.290 38.240 13.510 ;
        RECT 41.820 13.430 46.690 13.530 ;
        RECT 39.700 13.220 39.900 13.230 ;
        RECT 26.510 12.800 34.500 13.000 ;
        RECT 39.700 12.890 39.920 13.220 ;
        RECT 42.280 13.180 42.590 13.430 ;
        RECT 44.210 13.350 46.690 13.430 ;
        RECT 44.210 13.340 44.520 13.350 ;
        RECT 39.720 12.880 39.920 12.890 ;
        RECT 42.280 12.830 42.590 13.090 ;
        RECT 43.980 12.830 44.290 13.110 ;
        RECT 33.100 12.120 33.320 12.130 ;
        RECT 26.520 11.870 33.350 12.120 ;
        RECT 34.280 12.080 34.500 12.800 ;
        RECT 41.560 12.610 44.470 12.830 ;
        RECT 26.520 10.950 30.030 11.140 ;
        RECT 29.800 10.350 30.030 10.950 ;
        RECT 33.060 10.700 33.350 11.870 ;
        RECT 34.250 12.040 34.500 12.080 ;
        RECT 34.250 11.400 34.510 12.040 ;
        RECT 41.790 12.000 42.120 12.210 ;
        RECT 42.230 12.110 42.540 12.440 ;
        RECT 34.250 11.190 38.380 11.400 ;
        RECT 38.170 11.050 38.380 11.190 ;
        RECT 41.790 11.060 42.120 11.270 ;
        RECT 38.170 10.840 40.180 11.050 ;
        RECT 42.230 10.830 42.540 11.160 ;
        RECT 33.060 10.480 35.950 10.700 ;
        RECT 43.900 10.670 44.210 10.860 ;
        RECT 33.060 10.470 33.350 10.480 ;
        RECT 37.740 10.470 38.050 10.630 ;
        RECT 29.800 10.200 30.020 10.350 ;
        RECT 37.310 10.250 38.190 10.470 ;
        RECT 41.550 10.440 44.260 10.670 ;
        RECT 34.170 10.200 40.170 10.250 ;
        RECT 29.800 10.050 40.170 10.200 ;
        RECT 42.280 10.180 42.590 10.440 ;
        RECT 29.800 10.040 40.040 10.050 ;
        RECT 29.800 9.980 34.560 10.040 ;
        RECT 37.890 9.610 38.200 9.800 ;
        RECT 37.850 9.360 38.400 9.610 ;
        RECT 37.050 8.630 37.360 8.960 ;
        RECT 38.030 8.330 38.500 8.580 ;
        RECT 38.170 8.240 38.490 8.330 ;
        RECT 37.550 7.780 37.980 7.790 ;
        RECT 37.550 7.550 38.420 7.780 ;
        RECT 37.780 7.350 38.090 7.550 ;
  END
END sky130_hilas_TA2Cell_1FG_Strong

MACRO sky130_hilas_TA2Cell_NoFG
  CLASS CORE ;
  FOREIGN sky130_hilas_TA2Cell_NoFG ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.500 BY 24.010 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN COLSEL1
    PORT
      LAYER met1 ;
        RECT 10.570 14.950 10.760 15.030 ;
    END
  END COLSEL1
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 11.870 9.000 12.130 9.250 ;
    END
  END VIN12
  PIN VIN21
    PORT
      LAYER met2 ;
        RECT 13.470 12.090 13.720 12.320 ;
    END
  END VIN21
  PIN VIN22
    PORT
      LAYER met2 ;
        RECT 13.300 15.040 13.610 15.260 ;
        RECT 13.300 14.930 15.490 15.040 ;
        RECT 13.430 14.830 15.490 14.930 ;
        RECT 13.430 14.760 13.680 14.830 ;
    END
  END VIN22
  PIN OUTPUT1
    PORT
      LAYER met2 ;
        RECT 17.770 11.500 17.920 11.720 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    PORT
      LAYER met2 ;
        RECT 17.770 12.320 17.920 12.540 ;
    END
  END OUTPUT2
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 15.960 8.980 16.300 9.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.960 14.890 16.300 15.030 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 16.630 8.980 16.900 9.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 16.630 14.880 16.900 15.030 ;
    END
  END VPWR
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 0.000 14.350 0.070 14.530 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 0.000 9.500 0.080 9.650 ;
    END
  END DRAIN2
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 0.350 14.960 0.770 15.030 ;
    END
  END VTUN
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT 4.050 14.950 4.280 15.030 ;
    END
  END GATE1
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 11.010 14.950 11.290 15.030 ;
    END
  END VINJ
  PIN VIN11
    PORT
      LAYER met2 ;
        RECT 11.910 11.680 12.190 11.920 ;
    END
  END VIN11
  OBS
      LAYER nwell ;
        RECT 13.520 21.020 15.380 24.010 ;
        RECT 18.480 22.980 20.210 23.320 ;
        RECT 18.460 21.420 20.210 22.980 ;
        RECT 13.520 19.320 15.380 20.960 ;
        RECT 18.460 19.790 20.190 21.420 ;
        RECT 16.950 19.400 20.250 19.790 ;
        RECT 16.950 19.360 20.490 19.400 ;
        RECT 12.190 19.310 15.490 19.320 ;
        RECT 13.520 17.970 15.380 19.310 ;
        RECT 16.950 17.710 20.500 19.360 ;
        RECT 4.550 14.670 5.110 17.090 ;
        RECT 16.950 16.620 20.250 17.710 ;
        RECT 9.890 16.520 11.750 16.590 ;
        RECT 11.230 16.230 11.680 16.460 ;
        RECT 18.620 15.970 19.900 16.620 ;
        RECT 16.950 15.030 20.250 15.970 ;
        RECT 16.650 14.850 20.250 15.030 ;
        RECT 16.950 14.780 20.250 14.850 ;
        RECT 11.450 13.290 13.110 13.510 ;
        RECT 16.950 13.130 20.500 14.780 ;
        RECT 16.950 13.090 20.490 13.130 ;
        RECT 16.950 12.800 20.250 13.090 ;
        RECT 11.910 11.680 12.190 11.920 ;
        RECT 18.620 9.470 19.900 12.310 ;
        RECT 16.640 8.980 17.920 9.170 ;
        RECT 12.790 7.550 13.240 7.780 ;
        RECT 11.450 7.420 13.310 7.490 ;
        RECT 15.080 3.050 16.940 6.040 ;
        RECT 15.080 0.000 16.940 2.990 ;
      LAYER li1 ;
        RECT 13.930 21.490 14.110 23.540 ;
        RECT 14.740 21.750 14.910 23.530 ;
        RECT 14.660 21.580 14.990 21.750 ;
        RECT 18.880 21.590 19.430 22.020 ;
        RECT 13.930 18.440 14.110 20.490 ;
        RECT 14.740 18.700 14.910 20.480 ;
        RECT 18.880 19.860 19.430 20.290 ;
        RECT 17.840 19.160 18.370 19.330 ;
        RECT 19.650 19.060 19.850 19.410 ;
        RECT 19.650 19.030 19.860 19.060 ;
        RECT 14.660 18.530 14.990 18.700 ;
        RECT 18.080 18.230 18.310 18.920 ;
        RECT 13.310 17.940 13.630 17.980 ;
        RECT 13.310 17.750 13.640 17.940 ;
        RECT 13.310 17.720 13.630 17.750 ;
        RECT 11.490 17.310 11.680 17.330 ;
        RECT 11.350 17.220 11.680 17.310 ;
        RECT 11.350 17.140 11.430 17.220 ;
        RECT 11.490 17.100 11.680 17.220 ;
        RECT 18.090 17.080 18.260 18.230 ;
        RECT 18.920 17.170 19.090 18.780 ;
        RECT 19.640 18.450 19.860 19.030 ;
        RECT 19.650 18.440 19.860 18.450 ;
        RECT 19.290 18.270 19.480 18.280 ;
        RECT 19.290 17.980 19.490 18.270 ;
        RECT 19.280 17.650 19.570 17.980 ;
        RECT 7.000 16.430 7.190 16.750 ;
        RECT 6.910 16.340 7.190 16.430 ;
        RECT 10.300 16.340 10.480 17.060 ;
        RECT 10.950 16.690 11.120 17.020 ;
        RECT 18.920 16.980 19.100 17.170 ;
        RECT 11.030 16.620 11.080 16.690 ;
        RECT 11.030 16.590 11.370 16.620 ;
        RECT 10.910 16.580 11.370 16.590 ;
        RECT 10.910 16.460 11.380 16.580 ;
        RECT 11.050 16.390 11.380 16.460 ;
        RECT 19.180 16.540 19.510 16.710 ;
        RECT 19.620 16.630 19.950 16.800 ;
        RECT 11.050 16.360 11.370 16.390 ;
        RECT 6.910 16.200 10.550 16.340 ;
        RECT 19.180 16.260 19.540 16.540 ;
        RECT 7.000 16.160 10.550 16.200 ;
        RECT 7.000 15.740 7.190 16.160 ;
        RECT 10.300 16.000 10.480 16.160 ;
        RECT 17.110 16.010 17.430 16.050 ;
        RECT 17.110 15.820 17.440 16.010 ;
        RECT 17.110 15.790 17.430 15.820 ;
        RECT 17.510 15.800 17.710 16.130 ;
        RECT 18.100 15.940 18.300 16.130 ;
        RECT 18.830 16.090 19.540 16.260 ;
        RECT 18.770 15.970 19.090 16.010 ;
        RECT 17.790 15.610 17.980 15.620 ;
        RECT 17.990 15.610 18.340 15.940 ;
        RECT 18.770 15.780 19.100 15.970 ;
        RECT 18.770 15.750 19.090 15.780 ;
        RECT 10.320 15.300 10.640 15.340 ;
        RECT 8.030 15.120 8.260 15.160 ;
        RECT 10.320 15.110 10.650 15.300 ;
        RECT 13.310 15.180 13.630 15.220 ;
        RECT 10.320 15.080 10.640 15.110 ;
        RECT 13.310 14.990 13.640 15.180 ;
        RECT 16.880 15.100 17.050 15.430 ;
        RECT 17.060 15.360 17.380 15.400 ;
        RECT 17.060 15.170 17.390 15.360 ;
        RECT 17.060 15.140 17.380 15.170 ;
        RECT 17.510 15.140 17.710 15.470 ;
        RECT 17.790 15.280 18.340 15.610 ;
        RECT 13.310 14.960 13.630 14.990 ;
        RECT 17.990 14.950 18.340 15.280 ;
        RECT 18.090 14.610 18.260 14.950 ;
        RECT 18.830 14.940 19.530 15.650 ;
        RECT 18.830 14.770 19.570 14.940 ;
        RECT 11.130 14.480 11.450 14.510 ;
        RECT 11.120 14.290 11.450 14.480 ;
        RECT 18.090 14.380 18.360 14.610 ;
        RECT 18.090 14.320 18.260 14.380 ;
        RECT 18.920 14.350 19.090 14.770 ;
        RECT 19.280 14.610 19.570 14.770 ;
        RECT 19.290 14.350 19.490 14.610 ;
        RECT 11.130 14.250 11.450 14.290 ;
        RECT 10.970 13.680 11.140 13.990 ;
        RECT 16.880 13.840 17.050 14.170 ;
        RECT 17.060 14.100 17.380 14.130 ;
        RECT 17.060 13.910 17.390 14.100 ;
        RECT 17.060 13.870 17.380 13.910 ;
        RECT 17.510 13.800 17.710 14.130 ;
        RECT 17.990 13.990 18.340 14.320 ;
        RECT 18.820 14.170 19.520 14.350 ;
        RECT 10.970 13.660 11.300 13.680 ;
        RECT 10.980 13.650 11.300 13.660 ;
        RECT 17.790 13.660 18.340 13.990 ;
        RECT 18.920 13.810 19.090 14.170 ;
        RECT 19.650 14.140 19.860 14.150 ;
        RECT 17.790 13.650 17.980 13.660 ;
        RECT 10.970 13.460 11.300 13.650 ;
        RECT 10.980 13.420 11.300 13.460 ;
        RECT 17.110 13.450 17.430 13.480 ;
        RECT 17.110 13.260 17.440 13.450 ;
        RECT 17.110 13.220 17.430 13.260 ;
        RECT 17.510 13.140 17.710 13.470 ;
        RECT 17.990 13.430 18.340 13.660 ;
        RECT 18.820 13.750 19.140 13.790 ;
        RECT 18.820 13.560 19.150 13.750 ;
        RECT 19.640 13.560 19.860 14.140 ;
        RECT 18.820 13.530 19.140 13.560 ;
        RECT 19.650 13.530 19.860 13.560 ;
        RECT 17.840 13.260 18.370 13.430 ;
        RECT 18.100 13.140 18.300 13.260 ;
        RECT 19.650 13.180 19.850 13.530 ;
        RECT 17.110 13.010 17.430 13.050 ;
        RECT 17.110 12.820 17.440 13.010 ;
        RECT 17.110 12.790 17.430 12.820 ;
        RECT 17.510 12.800 17.710 13.130 ;
        RECT 18.100 12.940 18.300 13.130 ;
        RECT 18.810 13.030 19.130 13.070 ;
        RECT 17.790 12.610 17.980 12.620 ;
        RECT 17.990 12.610 18.340 12.940 ;
        RECT 18.810 12.840 19.140 13.030 ;
        RECT 18.810 12.810 19.130 12.840 ;
        RECT 2.830 11.450 3.290 12.460 ;
        RECT 16.880 12.100 17.050 12.430 ;
        RECT 17.060 12.360 17.380 12.400 ;
        RECT 17.060 12.170 17.390 12.360 ;
        RECT 17.060 12.140 17.380 12.170 ;
        RECT 17.510 12.140 17.710 12.470 ;
        RECT 17.790 12.280 18.340 12.610 ;
        RECT 17.990 12.020 18.340 12.280 ;
        RECT 17.990 11.950 18.360 12.020 ;
        RECT 18.170 11.790 18.360 11.950 ;
        RECT 18.820 11.890 19.520 12.070 ;
        RECT 16.880 10.840 17.050 11.170 ;
        RECT 17.060 11.100 17.380 11.130 ;
        RECT 17.060 10.910 17.390 11.100 ;
        RECT 17.060 10.870 17.380 10.910 ;
        RECT 17.510 10.800 17.710 11.130 ;
        RECT 17.990 10.990 18.340 11.320 ;
        RECT 17.790 10.660 18.340 10.990 ;
        RECT 18.830 10.820 19.530 11.470 ;
        RECT 17.790 10.650 17.980 10.660 ;
        RECT 12.540 10.550 12.860 10.590 ;
        RECT 12.530 10.360 12.860 10.550 ;
        RECT 12.540 10.350 12.860 10.360 ;
        RECT 12.530 10.330 12.860 10.350 ;
        RECT 17.110 10.450 17.430 10.480 ;
        RECT 12.530 10.020 12.700 10.330 ;
        RECT 17.110 10.260 17.440 10.450 ;
        RECT 17.110 10.220 17.430 10.260 ;
        RECT 17.510 10.140 17.710 10.470 ;
        RECT 17.990 10.330 18.340 10.660 ;
        RECT 18.730 10.590 19.530 10.820 ;
        RECT 18.730 10.560 19.050 10.590 ;
        RECT 18.100 10.140 18.300 10.330 ;
        RECT 18.830 9.980 19.540 10.150 ;
        RECT 12.690 9.720 13.010 9.760 ;
        RECT 12.680 9.530 13.010 9.720 ;
        RECT 19.180 9.700 19.540 9.980 ;
        RECT 19.180 9.530 19.510 9.700 ;
        RECT 12.690 9.500 13.010 9.530 ;
        RECT 19.620 9.440 19.950 9.610 ;
        RECT 11.880 8.900 12.200 8.930 ;
        RECT 11.880 8.710 12.210 8.900 ;
        RECT 11.880 8.670 12.200 8.710 ;
        RECT 11.860 6.950 12.040 8.010 ;
        RECT 12.610 7.620 12.930 7.650 ;
        RECT 12.610 7.550 12.940 7.620 ;
        RECT 12.470 7.430 12.940 7.550 ;
        RECT 12.470 7.420 12.930 7.430 ;
        RECT 12.590 7.390 12.930 7.420 ;
        RECT 12.590 7.320 12.640 7.390 ;
        RECT 12.510 6.990 12.680 7.320 ;
        RECT 12.910 6.790 12.990 6.870 ;
        RECT 13.050 6.790 13.240 6.910 ;
        RECT 12.910 6.700 13.240 6.790 ;
        RECT 13.050 6.680 13.240 6.700 ;
        RECT 15.490 3.520 15.670 5.570 ;
        RECT 16.220 5.310 16.550 5.480 ;
        RECT 16.300 3.530 16.470 5.310 ;
        RECT 15.490 0.470 15.670 2.520 ;
        RECT 16.220 2.260 16.550 2.430 ;
        RECT 16.300 0.480 16.470 2.260 ;
      LAYER mcon ;
        RECT 18.880 21.670 19.150 21.940 ;
        RECT 18.880 19.940 19.150 20.210 ;
        RECT 18.110 18.710 18.280 18.880 ;
        RECT 19.660 18.860 19.830 19.030 ;
        RECT 18.110 18.260 18.280 18.430 ;
        RECT 13.370 17.760 13.540 17.930 ;
        RECT 11.500 17.130 11.670 17.300 ;
        RECT 19.300 18.020 19.480 18.210 ;
        RECT 6.920 16.230 7.090 16.400 ;
        RECT 11.110 16.400 11.280 16.570 ;
        RECT 17.170 15.830 17.340 16.000 ;
        RECT 18.830 15.790 19.000 15.960 ;
        RECT 10.380 15.120 10.550 15.290 ;
        RECT 13.370 15.000 13.540 15.170 ;
        RECT 17.120 15.180 17.290 15.350 ;
        RECT 18.110 15.440 18.280 15.610 ;
        RECT 18.920 15.420 19.100 15.610 ;
        RECT 11.220 14.300 11.390 14.470 ;
        RECT 18.180 14.410 18.350 14.580 ;
        RECT 19.300 14.380 19.480 14.570 ;
        RECT 17.120 13.920 17.290 14.090 ;
        RECT 18.110 14.060 18.280 14.230 ;
        RECT 11.070 13.470 11.240 13.640 ;
        RECT 18.110 13.610 18.280 13.830 ;
        RECT 17.170 13.270 17.340 13.440 ;
        RECT 18.880 13.570 19.050 13.740 ;
        RECT 19.660 13.560 19.830 13.730 ;
        RECT 17.170 12.830 17.340 13.000 ;
        RECT 18.870 12.850 19.040 13.020 ;
        RECT 2.860 12.200 3.030 12.370 ;
        RECT 17.120 12.180 17.290 12.350 ;
        RECT 18.110 12.440 18.280 12.610 ;
        RECT 18.180 11.820 18.350 11.990 ;
        RECT 2.860 11.510 3.030 11.680 ;
        RECT 17.120 10.920 17.290 11.090 ;
        RECT 18.110 10.660 18.280 10.830 ;
        RECT 12.630 10.370 12.800 10.540 ;
        RECT 17.170 10.270 17.340 10.440 ;
        RECT 18.790 10.600 18.960 10.770 ;
        RECT 12.780 9.540 12.950 9.710 ;
        RECT 11.940 8.720 12.110 8.890 ;
        RECT 12.670 7.440 12.840 7.610 ;
        RECT 13.060 6.710 13.230 6.880 ;
      LAYER met1 ;
        RECT 18.820 19.400 19.210 22.990 ;
        RECT 4.310 13.270 4.730 19.320 ;
        RECT 6.790 16.460 7.020 19.320 ;
        RECT 6.790 16.170 7.120 16.460 ;
        RECT 6.790 13.270 7.020 16.170 ;
        RECT 8.010 13.270 8.240 19.320 ;
        RECT 14.530 19.280 14.720 19.320 ;
        RECT 13.300 17.690 13.620 18.010 ;
        RECT 11.470 17.070 11.700 17.360 ;
        RECT 11.040 16.330 11.360 16.650 ;
        RECT 11.390 15.800 11.600 17.040 ;
        RECT 14.220 16.530 14.480 16.850 ;
        RECT 14.970 16.570 15.250 19.320 ;
        RECT 17.770 18.970 18.080 19.360 ;
        RECT 17.770 18.920 18.320 18.970 ;
        RECT 18.060 18.180 18.320 18.920 ;
        RECT 19.290 18.280 19.480 19.730 ;
        RECT 19.730 19.090 19.890 19.730 ;
        RECT 19.620 18.540 19.890 19.090 ;
        RECT 19.620 18.490 19.900 18.540 ;
        RECT 19.730 18.400 19.900 18.490 ;
        RECT 19.290 18.250 19.510 18.280 ;
        RECT 19.270 17.980 19.520 18.250 ;
        RECT 19.280 17.970 19.520 17.980 ;
        RECT 19.280 17.730 19.510 17.970 ;
        RECT 18.890 16.920 19.130 17.300 ;
        RECT 19.320 16.710 19.480 17.730 ;
        RECT 19.730 16.710 19.890 18.400 ;
        RECT 14.970 16.250 15.420 16.570 ;
        RECT 14.220 15.930 14.480 16.250 ;
        RECT 11.390 15.480 11.720 15.800 ;
        RECT 10.310 15.050 10.630 15.370 ;
        RECT 11.390 15.270 11.600 15.480 ;
        RECT 13.300 14.930 13.620 15.250 ;
        RECT 11.140 14.220 11.460 14.540 ;
        RECT 10.990 13.390 11.310 13.710 ;
        RECT 14.530 13.270 14.720 13.320 ;
        RECT 14.970 13.270 15.250 16.250 ;
        RECT 17.100 16.000 17.420 16.080 ;
        RECT 17.100 15.760 17.670 16.000 ;
        RECT 17.330 15.430 17.670 15.760 ;
        RECT 17.050 15.110 17.670 15.430 ;
        RECT 17.330 14.160 17.670 15.110 ;
        RECT 17.050 13.840 17.670 14.160 ;
        RECT 16.000 13.370 16.260 13.630 ;
        RECT 17.330 13.510 17.670 13.840 ;
        RECT 18.000 15.670 18.270 15.990 ;
        RECT 18.760 15.720 19.080 16.040 ;
        RECT 18.000 15.380 18.310 15.670 ;
        RECT 18.000 14.640 18.270 15.380 ;
        RECT 18.890 15.290 19.130 15.670 ;
        RECT 19.320 14.860 19.480 15.880 ;
        RECT 18.000 14.350 18.380 14.640 ;
        RECT 19.280 14.620 19.510 14.860 ;
        RECT 19.280 14.610 19.520 14.620 ;
        RECT 18.000 14.310 18.270 14.350 ;
        RECT 19.270 14.340 19.520 14.610 ;
        RECT 19.290 14.310 19.510 14.340 ;
        RECT 18.000 13.670 18.320 14.310 ;
        RECT 17.100 13.190 17.670 13.510 ;
        RECT 17.770 13.520 18.320 13.670 ;
        RECT 17.770 13.230 18.270 13.520 ;
        RECT 18.810 13.500 19.130 13.820 ;
        RECT 17.330 13.080 17.670 13.190 ;
        RECT 17.100 12.760 17.670 13.080 ;
        RECT 2.790 11.450 3.170 12.460 ;
        RECT 17.330 12.430 17.670 12.760 ;
        RECT 17.050 12.110 17.670 12.430 ;
        RECT 17.330 11.160 17.670 12.110 ;
        RECT 17.050 10.840 17.670 11.160 ;
        RECT 12.550 10.300 12.870 10.620 ;
        RECT 17.330 10.510 17.670 10.840 ;
        RECT 17.100 10.280 17.670 10.510 ;
        RECT 18.000 12.670 18.270 13.230 ;
        RECT 18.800 12.780 19.120 13.100 ;
        RECT 19.290 12.860 19.480 14.310 ;
        RECT 19.730 14.190 19.890 15.880 ;
        RECT 19.730 14.100 19.900 14.190 ;
        RECT 19.620 14.050 19.900 14.100 ;
        RECT 19.620 13.500 19.890 14.050 ;
        RECT 19.730 12.860 19.890 13.500 ;
        RECT 18.000 12.380 18.310 12.670 ;
        RECT 18.000 12.050 18.270 12.380 ;
        RECT 18.000 11.760 18.380 12.050 ;
        RECT 18.000 10.890 18.270 11.760 ;
        RECT 18.000 10.600 18.310 10.890 ;
        RECT 18.000 10.290 18.270 10.600 ;
        RECT 18.720 10.530 19.040 10.850 ;
        RECT 17.100 10.190 17.420 10.280 ;
        RECT 12.700 9.470 13.020 9.790 ;
        RECT 11.870 8.640 12.190 8.960 ;
        RECT 12.950 8.530 13.160 8.740 ;
        RECT 12.950 8.210 13.280 8.530 ;
        RECT 12.600 7.360 12.920 7.680 ;
        RECT 12.950 6.970 13.160 8.210 ;
        RECT 13.030 6.650 13.260 6.940 ;
      LAYER via ;
        RECT 13.330 17.720 13.590 17.980 ;
        RECT 11.070 16.360 11.330 16.620 ;
        RECT 14.220 16.560 14.480 16.820 ;
        RECT 17.800 18.950 18.060 19.210 ;
        RECT 15.160 16.280 15.420 16.540 ;
        RECT 14.220 15.960 14.480 16.220 ;
        RECT 11.460 15.510 11.720 15.770 ;
        RECT 10.340 15.080 10.600 15.340 ;
        RECT 13.330 14.960 13.590 15.220 ;
        RECT 11.170 14.250 11.430 14.510 ;
        RECT 11.020 13.420 11.280 13.680 ;
        RECT 17.130 15.790 17.390 16.050 ;
        RECT 17.080 15.140 17.340 15.400 ;
        RECT 17.080 13.870 17.340 14.130 ;
        RECT 18.790 15.750 19.050 16.010 ;
        RECT 17.130 13.220 17.390 13.480 ;
        RECT 17.800 13.380 18.060 13.640 ;
        RECT 18.840 13.530 19.100 13.790 ;
        RECT 17.130 12.790 17.390 13.050 ;
        RECT 2.830 11.490 3.120 12.420 ;
        RECT 17.080 12.140 17.340 12.400 ;
        RECT 17.080 10.870 17.340 11.130 ;
        RECT 12.580 10.330 12.840 10.590 ;
        RECT 17.130 10.220 17.390 10.480 ;
        RECT 18.830 12.810 19.090 13.070 ;
        RECT 18.750 10.560 19.010 10.820 ;
        RECT 12.730 9.500 12.990 9.760 ;
        RECT 11.900 8.670 12.160 8.930 ;
        RECT 13.020 8.240 13.280 8.500 ;
        RECT 12.630 7.390 12.890 7.650 ;
      LAYER met2 ;
        RECT 17.770 19.240 18.080 19.250 ;
        RECT 17.770 19.060 20.250 19.240 ;
        RECT 17.770 18.920 18.080 19.060 ;
        RECT 3.960 18.640 13.080 18.820 ;
        RECT 13.300 17.800 13.610 18.020 ;
        RECT 13.300 17.690 15.490 17.800 ;
        RECT 13.460 17.580 15.490 17.690 ;
        RECT 11.040 16.460 11.350 16.660 ;
        RECT 14.190 16.560 14.510 16.820 ;
        RECT 15.130 16.460 15.450 16.540 ;
        RECT 10.810 16.230 11.680 16.460 ;
        RECT 14.140 16.280 15.450 16.460 ;
        RECT 10.810 16.220 11.240 16.230 ;
        RECT 14.140 16.110 15.320 16.280 ;
        RECT 14.190 15.960 14.510 16.110 ;
        RECT 17.100 15.800 17.410 16.090 ;
        RECT 18.760 15.800 19.070 16.050 ;
        RECT 11.430 15.680 11.750 15.770 ;
        RECT 16.380 15.720 19.070 15.800 ;
        RECT 11.290 15.430 11.760 15.680 ;
        RECT 16.380 15.570 18.920 15.720 ;
        RECT 10.310 15.050 10.620 15.380 ;
        RECT 16.610 15.000 16.940 15.210 ;
        RECT 17.050 15.110 17.360 15.440 ;
        RECT 11.110 14.400 11.660 14.650 ;
        RECT 11.150 14.210 11.460 14.400 ;
        RECT 13.020 13.940 13.180 13.960 ;
        RECT 3.960 13.890 13.180 13.940 ;
        RECT 3.960 13.790 13.060 13.890 ;
        RECT 10.570 13.540 11.450 13.790 ;
        RECT 14.490 13.780 14.740 14.150 ;
        RECT 16.610 14.060 16.940 14.270 ;
        RECT 17.050 13.830 17.360 14.160 ;
        RECT 15.960 13.580 16.300 13.670 ;
        RECT 17.770 13.660 18.080 13.670 ;
        RECT 18.810 13.660 19.120 13.830 ;
        RECT 11.000 13.380 11.310 13.540 ;
        RECT 11.450 13.290 13.110 13.510 ;
        RECT 13.610 13.390 16.300 13.580 ;
        RECT 16.640 13.530 19.290 13.660 ;
        RECT 16.640 13.430 20.250 13.530 ;
        RECT 13.610 12.820 13.800 13.390 ;
        RECT 15.960 13.340 16.300 13.390 ;
        RECT 14.520 12.930 14.730 13.220 ;
        RECT 17.100 13.180 17.410 13.430 ;
        RECT 17.770 13.350 20.250 13.430 ;
        RECT 17.770 13.340 18.080 13.350 ;
        RECT 17.100 12.830 17.410 13.090 ;
        RECT 18.800 12.830 19.110 13.110 ;
        RECT 2.820 12.630 13.800 12.820 ;
        RECT 2.820 12.450 3.010 12.630 ;
        RECT 16.380 12.610 19.290 12.830 ;
        RECT 2.800 11.460 3.150 12.450 ;
        RECT 16.610 12.000 16.940 12.210 ;
        RECT 17.050 12.110 17.360 12.440 ;
        RECT 16.610 11.060 16.940 11.270 ;
        RECT 12.960 10.850 14.730 11.050 ;
        RECT 17.050 10.830 17.360 11.160 ;
        RECT 11.390 10.360 11.550 10.760 ;
        RECT 18.720 10.670 19.030 10.860 ;
        RECT 12.560 10.470 12.870 10.630 ;
        RECT 12.130 10.250 13.010 10.470 ;
        RECT 16.370 10.440 19.080 10.670 ;
        RECT 12.130 10.220 14.730 10.250 ;
        RECT 12.670 10.040 14.730 10.220 ;
        RECT 17.100 10.180 17.410 10.440 ;
        RECT 12.710 9.610 13.020 9.800 ;
        RECT 12.670 9.360 13.220 9.610 ;
        RECT 11.870 8.630 12.180 8.960 ;
        RECT 12.850 8.330 13.320 8.580 ;
        RECT 12.990 8.240 13.310 8.330 ;
        RECT 12.370 7.780 12.800 7.790 ;
        RECT 12.370 7.550 13.240 7.780 ;
        RECT 12.600 7.350 12.910 7.550 ;
  END
END sky130_hilas_TA2Cell_NoFG

MACRO sky130_hilas_pFETLarge
  CLASS CORE ;
  FOREIGN sky130_hilas_pFETLarge ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.640 BY 5.990 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA 6.540500 ;
    PORT
      LAYER met2 ;
        RECT 0.430 0.830 0.740 0.960 ;
        RECT 0.000 0.630 0.740 0.830 ;
        RECT 0.000 0.490 0.600 0.630 ;
        RECT 0.000 0.160 0.750 0.490 ;
        RECT 0.000 0.010 0.600 0.160 ;
    END
  END GATE
  PIN SOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 4.358700 ;
    PORT
      LAYER met2 ;
        RECT 1.010 5.610 1.320 5.750 ;
        RECT 2.100 5.610 2.410 5.750 ;
        RECT 3.200 5.610 3.510 5.740 ;
        RECT 0.330 5.600 3.510 5.610 ;
        RECT 0.240 5.410 3.510 5.600 ;
        RECT 0.240 5.270 3.390 5.410 ;
        RECT 0.240 2.820 0.560 5.270 ;
        RECT 1.000 2.820 1.310 2.970 ;
        RECT 2.100 2.820 2.410 2.970 ;
        RECT 3.200 2.820 3.510 2.970 ;
        RECT 0.240 2.640 3.510 2.820 ;
        RECT 0.240 2.490 3.400 2.640 ;
        RECT 0.240 1.450 0.560 2.490 ;
        RECT 1.000 1.450 1.310 1.600 ;
        RECT 2.100 1.450 2.410 1.600 ;
        RECT 3.200 1.450 3.510 1.600 ;
        RECT 0.240 1.270 3.510 1.450 ;
        RECT 0.240 1.130 3.400 1.270 ;
    END
  END SOURCE
  PIN DRAIN
    USE ANALOG ;
    ANTENNADIFFAREA 4.311400 ;
    PORT
      LAYER met2 ;
        RECT 1.560 4.890 1.870 5.070 ;
        RECT 2.650 4.890 2.960 5.050 ;
        RECT 3.760 4.890 4.070 5.040 ;
        RECT 1.430 4.590 4.370 4.890 ;
        RECT 3.620 4.550 4.370 4.590 ;
        RECT 3.990 4.420 4.370 4.550 ;
        RECT 4.020 3.700 4.370 4.420 ;
        RECT 1.560 3.550 1.870 3.700 ;
        RECT 2.650 3.550 2.960 3.700 ;
        RECT 3.750 3.550 4.370 3.700 ;
        RECT 1.420 3.220 4.370 3.550 ;
        RECT 4.020 0.930 4.370 3.220 ;
        RECT 1.560 0.780 1.870 0.920 ;
        RECT 2.650 0.780 2.960 0.920 ;
        RECT 3.750 0.780 4.370 0.930 ;
        RECT 1.430 0.460 4.370 0.780 ;
        RECT 1.430 0.450 4.140 0.460 ;
    END
  END DRAIN
  PIN WELL
    USE ANALOG ;
    ANTENNADIFFAREA 0.213200 ;
    PORT
      LAYER nwell ;
        RECT 0.780 5.880 4.170 5.970 ;
        RECT 0.780 0.270 4.640 5.880 ;
        RECT 4.020 0.180 4.640 0.270 ;
      LAYER met1 ;
        RECT 4.140 5.790 4.400 5.990 ;
        RECT 4.140 4.980 4.450 5.790 ;
        RECT 4.140 0.000 4.400 4.980 ;
    END
  END WELL
  OBS
      LAYER li1 ;
        RECT 1.020 5.710 1.190 5.740 ;
        RECT 1.020 5.670 1.340 5.710 ;
        RECT 1.020 5.480 1.350 5.670 ;
        RECT 1.020 5.450 1.340 5.480 ;
        RECT 1.020 3.250 1.190 5.450 ;
        RECT 1.570 5.030 1.740 5.740 ;
        RECT 2.120 5.710 2.290 5.740 ;
        RECT 2.110 5.670 2.430 5.710 ;
        RECT 2.110 5.480 2.440 5.670 ;
        RECT 2.110 5.450 2.430 5.480 ;
        RECT 1.570 4.990 1.890 5.030 ;
        RECT 1.570 4.800 1.900 4.990 ;
        RECT 1.570 4.770 1.890 4.800 ;
        RECT 1.570 3.660 1.740 4.770 ;
        RECT 1.570 3.620 1.890 3.660 ;
        RECT 1.570 3.430 1.900 3.620 ;
        RECT 1.570 3.400 1.890 3.430 ;
        RECT 1.570 3.240 1.740 3.400 ;
        RECT 2.120 3.240 2.290 5.450 ;
        RECT 2.670 5.010 2.840 5.740 ;
        RECT 3.220 5.700 3.390 5.740 ;
        RECT 3.210 5.660 3.530 5.700 ;
        RECT 3.210 5.470 3.540 5.660 ;
        RECT 3.210 5.440 3.530 5.470 ;
        RECT 2.660 4.970 2.980 5.010 ;
        RECT 2.660 4.780 2.990 4.970 ;
        RECT 2.660 4.750 2.980 4.780 ;
        RECT 2.670 3.660 2.840 4.750 ;
        RECT 2.660 3.620 2.980 3.660 ;
        RECT 2.660 3.430 2.990 3.620 ;
        RECT 2.660 3.400 2.980 3.430 ;
        RECT 2.670 3.240 2.840 3.400 ;
        RECT 3.220 3.240 3.390 5.440 ;
        RECT 3.770 5.000 3.940 5.740 ;
        RECT 3.770 4.960 4.090 5.000 ;
        RECT 3.770 4.770 4.100 4.960 ;
        RECT 4.250 4.920 4.420 5.680 ;
        RECT 3.770 4.740 4.090 4.770 ;
        RECT 3.770 3.660 3.940 4.740 ;
        RECT 3.760 3.620 4.080 3.660 ;
        RECT 3.760 3.430 4.090 3.620 ;
        RECT 3.760 3.400 4.080 3.430 ;
        RECT 3.770 3.240 3.940 3.400 ;
        RECT 0.960 3.160 1.120 3.190 ;
        RECT 0.960 2.930 1.130 3.160 ;
        RECT 1.510 3.150 1.670 3.190 ;
        RECT 0.960 2.890 1.330 2.930 ;
        RECT 1.510 2.910 1.680 3.150 ;
        RECT 2.060 2.930 2.230 3.220 ;
        RECT 2.610 3.150 2.770 3.190 ;
        RECT 3.160 3.150 3.320 3.190 ;
        RECT 3.710 3.170 3.870 3.190 ;
        RECT 0.960 2.810 1.340 2.890 ;
        RECT 1.510 2.810 1.740 2.910 ;
        RECT 2.060 2.890 2.430 2.930 ;
        RECT 2.610 2.910 2.780 3.150 ;
        RECT 3.160 2.930 3.330 3.150 ;
        RECT 2.060 2.810 2.440 2.890 ;
        RECT 2.610 2.810 2.840 2.910 ;
        RECT 3.160 2.890 3.530 2.930 ;
        RECT 3.710 2.910 3.880 3.170 ;
        RECT 3.160 2.810 3.540 2.890 ;
        RECT 3.710 2.810 3.940 2.910 ;
        RECT 1.010 2.700 1.340 2.810 ;
        RECT 1.010 2.670 1.330 2.700 ;
        RECT 1.020 1.560 1.190 2.670 ;
        RECT 1.010 1.520 1.330 1.560 ;
        RECT 1.010 1.330 1.340 1.520 ;
        RECT 1.010 1.300 1.330 1.330 ;
        RECT 0.190 0.940 0.700 1.020 ;
        RECT 0.190 0.920 0.710 0.940 ;
        RECT 0.190 0.880 0.760 0.920 ;
        RECT 0.190 0.690 0.770 0.880 ;
        RECT 0.200 0.660 0.760 0.690 ;
        RECT 0.200 0.450 0.710 0.660 ;
        RECT 0.200 0.410 0.770 0.450 ;
        RECT 1.020 0.420 1.190 1.300 ;
        RECT 1.570 0.880 1.740 2.810 ;
        RECT 2.110 2.700 2.440 2.810 ;
        RECT 2.110 2.670 2.430 2.700 ;
        RECT 2.120 1.560 2.290 2.670 ;
        RECT 2.110 1.520 2.430 1.560 ;
        RECT 2.110 1.330 2.440 1.520 ;
        RECT 2.110 1.300 2.430 1.330 ;
        RECT 1.570 0.840 1.890 0.880 ;
        RECT 1.570 0.650 1.900 0.840 ;
        RECT 1.570 0.620 1.890 0.650 ;
        RECT 1.570 0.410 1.740 0.620 ;
        RECT 2.120 0.410 2.290 1.300 ;
        RECT 2.670 0.880 2.840 2.810 ;
        RECT 3.210 2.700 3.540 2.810 ;
        RECT 3.210 2.670 3.530 2.700 ;
        RECT 3.220 1.560 3.390 2.670 ;
        RECT 3.210 1.520 3.530 1.560 ;
        RECT 3.210 1.330 3.540 1.520 ;
        RECT 3.210 1.300 3.530 1.330 ;
        RECT 2.660 0.840 2.980 0.880 ;
        RECT 2.660 0.650 2.990 0.840 ;
        RECT 2.660 0.620 2.980 0.650 ;
        RECT 2.670 0.410 2.840 0.620 ;
        RECT 3.220 0.410 3.390 1.300 ;
        RECT 3.770 0.890 3.940 2.810 ;
        RECT 3.760 0.850 4.080 0.890 ;
        RECT 3.760 0.660 4.090 0.850 ;
        RECT 3.760 0.630 4.080 0.660 ;
        RECT 3.770 0.410 3.940 0.630 ;
        RECT 0.200 0.220 0.780 0.410 ;
        RECT 0.200 0.190 0.770 0.220 ;
        RECT 0.200 0.010 0.710 0.190 ;
      LAYER mcon ;
        RECT 1.080 5.490 1.250 5.660 ;
        RECT 2.170 5.490 2.340 5.660 ;
        RECT 1.630 4.810 1.800 4.980 ;
        RECT 1.630 3.440 1.800 3.610 ;
        RECT 3.270 5.480 3.440 5.650 ;
        RECT 2.720 4.790 2.890 4.960 ;
        RECT 2.720 3.440 2.890 3.610 ;
        RECT 4.250 5.510 4.420 5.680 ;
        RECT 4.250 5.150 4.420 5.320 ;
        RECT 3.830 4.780 4.000 4.950 ;
        RECT 3.820 3.440 3.990 3.610 ;
        RECT 1.070 2.710 1.240 2.880 ;
        RECT 1.070 1.340 1.240 1.510 ;
        RECT 0.500 0.700 0.670 0.870 ;
        RECT 2.170 2.710 2.340 2.880 ;
        RECT 2.170 1.340 2.340 1.510 ;
        RECT 1.630 0.660 1.800 0.830 ;
        RECT 3.270 2.710 3.440 2.880 ;
        RECT 3.270 1.340 3.440 1.510 ;
        RECT 2.720 0.660 2.890 0.830 ;
        RECT 3.820 0.670 3.990 0.840 ;
        RECT 0.510 0.230 0.680 0.400 ;
      LAYER met1 ;
        RECT 1.010 5.420 1.330 5.740 ;
        RECT 2.100 5.420 2.420 5.740 ;
        RECT 3.200 5.410 3.520 5.730 ;
        RECT 1.560 4.740 1.880 5.060 ;
        RECT 2.650 4.720 2.970 5.040 ;
        RECT 3.760 4.710 4.080 5.030 ;
        RECT 1.560 3.370 1.880 3.690 ;
        RECT 2.650 3.370 2.970 3.690 ;
        RECT 3.750 3.370 4.070 3.690 ;
        RECT 1.000 2.640 1.320 2.960 ;
        RECT 2.100 2.640 2.420 2.960 ;
        RECT 3.200 2.640 3.520 2.960 ;
        RECT 1.000 1.270 1.320 1.590 ;
        RECT 2.100 1.270 2.420 1.590 ;
        RECT 3.200 1.270 3.520 1.590 ;
        RECT 0.430 0.630 0.750 0.950 ;
        RECT 1.560 0.590 1.880 0.910 ;
        RECT 2.650 0.590 2.970 0.910 ;
        RECT 3.750 0.600 4.070 0.920 ;
        RECT 0.440 0.160 0.760 0.480 ;
      LAYER via ;
        RECT 1.040 5.450 1.300 5.710 ;
        RECT 2.130 5.450 2.390 5.710 ;
        RECT 3.230 5.440 3.490 5.700 ;
        RECT 1.590 4.770 1.850 5.030 ;
        RECT 2.680 4.750 2.940 5.010 ;
        RECT 3.790 4.740 4.050 5.000 ;
        RECT 1.590 3.400 1.850 3.660 ;
        RECT 2.680 3.400 2.940 3.660 ;
        RECT 3.780 3.400 4.040 3.660 ;
        RECT 1.030 2.670 1.290 2.930 ;
        RECT 2.130 2.670 2.390 2.930 ;
        RECT 3.230 2.670 3.490 2.930 ;
        RECT 1.030 1.300 1.290 1.560 ;
        RECT 2.130 1.300 2.390 1.560 ;
        RECT 3.230 1.300 3.490 1.560 ;
        RECT 0.460 0.660 0.720 0.920 ;
        RECT 1.590 0.620 1.850 0.880 ;
        RECT 2.680 0.620 2.940 0.880 ;
        RECT 3.780 0.630 4.040 0.890 ;
        RECT 0.470 0.190 0.730 0.450 ;
  END
END sky130_hilas_pFETLarge

MACRO sky130_hilas_VinjInv2
  CLASS CORE ;
  FOREIGN sky130_hilas_VinjInv2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.610 BY 1.640 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 0.000 0.000 1.980 1.640 ;
      LAYER li1 ;
        RECT 0.620 1.210 0.790 1.350 ;
        RECT 0.620 1.040 0.810 1.210 ;
        RECT 0.620 0.940 0.790 1.040 ;
        RECT 0.190 0.560 0.360 0.660 ;
        RECT 0.170 0.390 0.360 0.560 ;
        RECT 0.190 0.330 0.360 0.390 ;
        RECT 0.610 0.600 0.780 0.660 ;
        RECT 0.610 0.330 0.860 0.600 ;
        RECT 1.350 0.580 1.600 0.660 ;
        RECT 1.350 0.410 2.650 0.580 ;
        RECT 3.210 0.570 3.380 1.200 ;
        RECT 0.620 0.310 0.860 0.330 ;
        RECT 1.430 0.320 1.600 0.410 ;
        RECT 3.130 0.400 3.460 0.570 ;
      LAYER mcon ;
        RECT 0.640 1.040 0.810 1.210 ;
        RECT 3.210 0.680 3.380 0.850 ;
        RECT 0.650 0.360 0.820 0.530 ;
        RECT 1.990 0.410 2.160 0.580 ;
      LAYER met1 ;
        RECT 0.610 1.260 0.830 1.600 ;
        RECT 0.610 1.000 0.840 1.260 ;
        RECT 0.080 0.320 0.390 0.670 ;
        RECT 0.610 0.600 0.830 1.000 ;
        RECT 0.610 0.290 0.860 0.600 ;
        RECT 1.910 0.360 2.230 0.620 ;
        RECT 0.610 0.090 0.830 0.290 ;
        RECT 3.180 0.090 3.410 1.600 ;
      LAYER via ;
        RECT 0.110 0.350 0.370 0.610 ;
        RECT 1.940 0.360 2.200 0.620 ;
      LAYER met2 ;
        RECT 0.000 1.030 3.610 1.210 ;
        RECT 0.080 0.510 0.400 0.610 ;
        RECT 0.070 0.350 0.400 0.510 ;
        RECT 1.910 0.540 2.230 0.620 ;
        RECT 1.910 0.360 3.610 0.540 ;
  END
END sky130_hilas_VinjInv2

MACRO sky130_hilas_capacitorSize03
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize03 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.720 BY 7.900 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.420 2.410 5.790 2.690 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.020 2.370 0.290 2.650 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 0.000 4.850 5.780 5.030 ;
        RECT 0.000 4.420 5.780 4.600 ;
        RECT 0.030 3.420 5.780 3.600 ;
        RECT 0.030 3.110 5.780 3.170 ;
        RECT 0.030 2.990 5.820 3.110 ;
        RECT 0.600 2.670 0.970 2.990 ;
        RECT 5.450 2.710 5.820 2.990 ;
        RECT 0.030 1.840 5.780 2.010 ;
        RECT 0.030 1.420 5.780 1.590 ;
        RECT 0.030 0.440 5.780 0.610 ;
        RECT 0.030 0.000 5.780 0.170 ;
      LAYER via2 ;
        RECT 0.650 2.730 0.930 3.010 ;
        RECT 5.500 2.770 5.780 3.050 ;
      LAYER met3 ;
        RECT 5.880 5.040 8.720 7.900 ;
        RECT 5.880 3.260 8.720 4.890 ;
        RECT 0.380 2.470 1.170 3.220 ;
        RECT 1.450 2.900 1.720 2.910 ;
        RECT 5.230 2.900 8.720 3.260 ;
        RECT 1.450 2.510 8.720 2.900 ;
        RECT 1.450 2.150 5.590 2.510 ;
        RECT 5.880 2.030 8.720 2.510 ;
      LAYER via3 ;
        RECT 0.570 2.620 1.000 3.100 ;
        RECT 5.420 2.660 5.850 3.140 ;
      LAYER met4 ;
        RECT 7.000 6.560 7.450 6.570 ;
        RECT 6.980 6.070 7.500 6.560 ;
        RECT 0.470 2.770 1.130 3.190 ;
        RECT 2.580 2.780 3.020 3.620 ;
        RECT 7.000 3.550 7.450 3.560 ;
        RECT 1.160 2.770 2.170 2.780 ;
        RECT 2.570 2.770 3.030 2.780 ;
        RECT 0.450 2.270 3.030 2.770 ;
        RECT 5.320 2.570 5.980 3.230 ;
        RECT 6.980 3.060 7.500 3.550 ;
        RECT 0.450 2.260 1.520 2.270 ;
        RECT 2.570 1.610 3.030 2.270 ;
        RECT 2.570 1.110 3.050 1.610 ;
        RECT 3.020 0.810 3.050 1.110 ;
  END
END sky130_hilas_capacitorSize03

MACRO sky130_hilas_swc4x1BiasCell
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x1BiasCell ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.250 BY 10.910 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN ROW1
    PORT
      LAYER met2 ;
        RECT 9.990 5.740 10.080 5.920 ;
    END
  END ROW1
  PIN ROW2
    PORT
      LAYER met2 ;
        RECT 9.990 4.650 10.080 4.830 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.010 4.650 7.640 4.830 ;
    END
  END ROW2
  PIN ROW3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.010 2.540 0.480 2.700 ;
        RECT 0.020 2.530 0.480 2.540 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.970 2.500 10.080 2.680 ;
    END
  END ROW3
  PIN ROW4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.010 1.550 7.640 1.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.970 1.400 10.080 1.580 ;
    END
  END ROW4
  PIN VTUN
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 0.360 0.410 0.760 6.910 ;
    END
  END VTUN
  PIN GATE1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 4.410 0.410 4.790 0.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.410 6.540 4.790 6.910 ;
    END
  END GATE1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 9.560 6.570 9.720 6.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 9.560 0.600 9.720 0.670 ;
    END
  END VINJ
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 8.750 6.570 8.910 6.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.750 0.600 8.910 0.670 ;
    END
  END VPWR
  PIN COLSEL1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 9.120 0.600 9.310 0.670 ;
    END
  END COLSEL1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 2.540 2.110 2.870 2.140 ;
        RECT 6.570 2.110 6.890 2.170 ;
        RECT 2.540 1.940 6.890 2.110 ;
        RECT 2.540 1.880 2.870 1.940 ;
        RECT 6.570 1.890 6.890 1.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.600 2.200 6.850 6.910 ;
        RECT 6.590 2.170 6.870 2.200 ;
        RECT 6.580 1.890 6.880 2.170 ;
        RECT 6.590 1.870 6.870 1.890 ;
        RECT 6.600 0.410 6.850 1.870 ;
      LAYER via ;
        RECT 6.600 1.900 6.860 2.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.570 2.170 2.840 6.910 ;
        RECT 2.550 1.860 2.860 2.170 ;
        RECT 2.570 0.410 2.840 1.860 ;
      LAYER via ;
        RECT 2.570 1.880 2.840 2.140 ;
    END
  END VGND
  PIN DRAIN3
    PORT
      LAYER met2 ;
        RECT 9.970 2.930 10.080 3.110 ;
    END
  END DRAIN3
  PIN DRAIN4
    PORT
      LAYER met2 ;
        RECT 9.970 0.970 10.080 1.150 ;
    END
  END DRAIN4
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 9.990 6.170 10.080 6.350 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 9.990 4.220 10.080 4.400 ;
    END
  END DRAIN2
  OBS
      LAYER nwell ;
        RECT 14.520 10.850 16.250 10.910 ;
        RECT 10.410 5.410 12.970 7.320 ;
        RECT 0.580 5.180 1.170 5.340 ;
        RECT 4.320 5.120 5.430 5.390 ;
        RECT 7.520 4.200 7.610 4.280 ;
        RECT 8.960 3.700 9.130 3.760 ;
        RECT 8.960 3.690 9.310 3.700 ;
        RECT 8.960 3.590 9.130 3.690 ;
        RECT 9.300 3.590 9.310 3.690 ;
        RECT 10.410 2.170 12.970 5.160 ;
        RECT 13.330 4.410 16.250 10.850 ;
        RECT 18.520 7.280 20.250 9.120 ;
        RECT 13.330 4.360 15.560 4.410 ;
        RECT 0.580 1.940 1.170 2.090 ;
        RECT 4.320 1.920 5.430 2.110 ;
        RECT 10.410 0.000 12.970 1.910 ;
      LAYER li1 ;
        RECT 14.910 7.800 15.460 8.230 ;
        RECT 18.940 7.730 19.490 8.160 ;
        RECT 10.650 6.970 10.970 7.010 ;
        RECT 10.650 6.850 10.980 6.970 ;
        RECT 10.650 6.750 11.090 6.850 ;
        RECT 10.750 6.680 11.090 6.750 ;
        RECT 12.370 6.580 12.570 6.930 ;
        RECT 10.650 6.420 10.970 6.460 ;
        RECT 10.650 6.230 10.980 6.420 ;
        RECT 10.650 6.200 11.090 6.230 ;
        RECT 10.750 6.060 11.090 6.200 ;
        RECT 11.640 5.960 11.840 6.560 ;
        RECT 12.370 6.550 12.580 6.580 ;
        RECT 12.360 5.960 12.580 6.550 ;
        RECT 2.620 4.890 2.790 5.420 ;
        RECT 6.640 4.860 6.810 5.390 ;
        RECT 10.750 4.370 11.090 4.510 ;
        RECT 10.650 4.340 11.090 4.370 ;
        RECT 2.630 2.960 2.800 4.130 ;
        RECT 6.650 3.000 6.820 4.190 ;
        RECT 10.650 4.150 10.980 4.340 ;
        RECT 10.650 4.110 10.970 4.150 ;
        RECT 11.640 4.010 11.840 4.610 ;
        RECT 12.360 4.020 12.580 4.610 ;
        RECT 12.370 3.990 12.580 4.020 ;
        RECT 10.750 3.820 11.090 3.890 ;
        RECT 8.870 3.590 9.310 3.760 ;
        RECT 10.650 3.720 11.090 3.820 ;
        RECT 10.650 3.610 10.980 3.720 ;
        RECT 10.650 3.510 11.090 3.610 ;
        RECT 10.750 3.440 11.090 3.510 ;
        RECT 12.370 3.340 12.570 3.990 ;
        RECT 10.650 3.180 10.970 3.220 ;
        RECT 10.650 2.990 10.980 3.180 ;
        RECT 10.650 2.960 11.090 2.990 ;
        RECT 10.750 2.820 11.090 2.960 ;
        RECT 11.640 2.720 11.840 3.320 ;
        RECT 12.370 3.310 12.580 3.340 ;
        RECT 12.360 2.720 12.580 3.310 ;
        RECT 10.750 1.120 11.090 1.260 ;
        RECT 10.650 1.090 11.090 1.120 ;
        RECT 10.650 0.900 10.980 1.090 ;
        RECT 10.650 0.860 10.970 0.900 ;
        RECT 11.640 0.760 11.840 1.360 ;
        RECT 12.360 0.770 12.580 1.360 ;
        RECT 12.370 0.740 12.580 0.770 ;
        RECT 10.750 0.570 11.090 0.640 ;
        RECT 10.650 0.470 11.090 0.570 ;
        RECT 10.650 0.350 10.980 0.470 ;
        RECT 12.370 0.390 12.570 0.740 ;
        RECT 10.650 0.310 10.970 0.350 ;
      LAYER mcon ;
        RECT 14.910 7.880 15.180 8.150 ;
        RECT 18.940 7.810 19.210 8.080 ;
        RECT 10.710 6.790 10.880 6.960 ;
        RECT 10.710 6.240 10.880 6.410 ;
        RECT 11.650 6.350 11.820 6.520 ;
        RECT 12.380 6.380 12.550 6.550 ;
        RECT 2.620 5.250 2.790 5.420 ;
        RECT 6.640 5.220 6.810 5.390 ;
        RECT 2.630 3.960 2.800 4.130 ;
        RECT 2.630 3.320 2.800 3.490 ;
        RECT 6.650 4.020 6.820 4.190 ;
        RECT 10.710 4.160 10.880 4.330 ;
        RECT 11.650 4.050 11.820 4.220 ;
        RECT 12.380 4.020 12.550 4.190 ;
        RECT 9.130 3.590 9.310 3.760 ;
        RECT 6.650 3.360 6.820 3.530 ;
        RECT 10.710 3.550 10.880 3.780 ;
        RECT 10.710 3.000 10.880 3.170 ;
        RECT 11.650 3.110 11.820 3.280 ;
        RECT 12.380 3.140 12.550 3.310 ;
        RECT 10.710 0.910 10.880 1.080 ;
        RECT 11.650 0.800 11.820 0.970 ;
        RECT 12.380 0.770 12.550 0.940 ;
        RECT 10.710 0.360 10.880 0.530 ;
      LAYER met1 ;
        RECT 10.640 6.720 10.960 7.040 ;
        RECT 9.120 6.570 9.310 6.640 ;
        RECT 11.640 6.580 11.800 7.310 ;
        RECT 11.640 6.560 11.840 6.580 ;
        RECT 10.640 6.170 10.960 6.490 ;
        RECT 11.620 6.320 11.850 6.560 ;
        RECT 11.640 6.270 11.850 6.320 ;
        RECT 12.010 6.270 12.200 7.260 ;
        RECT 12.450 6.610 12.610 7.310 ;
        RECT 11.640 5.410 11.800 6.270 ;
        RECT 12.030 6.150 12.200 6.270 ;
        RECT 12.040 5.410 12.200 6.150 ;
        RECT 12.340 6.060 12.610 6.610 ;
        RECT 12.340 6.010 12.620 6.060 ;
        RECT 12.450 5.920 12.620 6.010 ;
        RECT 12.450 5.410 12.610 5.920 ;
        RECT 10.640 4.080 10.960 4.400 ;
        RECT 11.640 4.300 11.800 5.160 ;
        RECT 12.040 4.420 12.200 5.160 ;
        RECT 12.450 4.650 12.610 5.160 ;
        RECT 12.450 4.560 12.620 4.650 ;
        RECT 12.030 4.300 12.200 4.420 ;
        RECT 11.640 4.250 11.850 4.300 ;
        RECT 11.620 4.010 11.850 4.250 ;
        RECT 11.640 3.990 11.840 4.010 ;
        RECT 9.100 3.760 9.340 3.790 ;
        RECT 8.910 3.670 9.340 3.760 ;
        RECT 8.750 3.660 9.340 3.670 ;
        RECT 9.560 3.660 9.720 3.670 ;
        RECT 8.910 3.590 9.340 3.660 ;
        RECT 9.100 3.560 9.340 3.590 ;
        RECT 9.200 3.460 9.310 3.560 ;
        RECT 10.640 3.480 10.960 3.850 ;
        RECT 11.640 3.340 11.800 3.990 ;
        RECT 11.640 3.320 11.840 3.340 ;
        RECT 10.640 2.930 10.960 3.250 ;
        RECT 11.620 3.080 11.850 3.320 ;
        RECT 11.640 3.030 11.850 3.080 ;
        RECT 12.010 3.030 12.200 4.300 ;
        RECT 12.340 4.510 12.620 4.560 ;
        RECT 12.340 3.960 12.610 4.510 ;
        RECT 13.980 4.360 14.360 10.860 ;
        RECT 14.850 7.340 15.240 9.200 ;
        RECT 18.880 7.270 19.270 9.130 ;
        RECT 12.450 3.370 12.610 3.960 ;
        RECT 11.640 2.170 11.800 3.030 ;
        RECT 12.030 2.910 12.200 3.030 ;
        RECT 12.040 2.170 12.200 2.910 ;
        RECT 12.340 2.820 12.610 3.370 ;
        RECT 12.340 2.770 12.620 2.820 ;
        RECT 12.450 2.680 12.620 2.770 ;
        RECT 12.450 2.170 12.610 2.680 ;
        RECT 10.640 0.830 10.960 1.150 ;
        RECT 11.640 1.050 11.800 1.910 ;
        RECT 12.040 1.170 12.200 1.910 ;
        RECT 12.450 1.400 12.610 1.910 ;
        RECT 12.450 1.310 12.620 1.400 ;
        RECT 12.030 1.050 12.200 1.170 ;
        RECT 11.640 1.000 11.850 1.050 ;
        RECT 11.620 0.760 11.850 1.000 ;
        RECT 11.640 0.740 11.840 0.760 ;
        RECT 10.640 0.280 10.960 0.600 ;
        RECT 11.640 0.010 11.800 0.740 ;
        RECT 12.010 0.060 12.200 1.050 ;
        RECT 12.340 1.260 12.620 1.310 ;
        RECT 12.340 0.710 12.610 1.260 ;
        RECT 12.450 0.010 12.610 0.710 ;
      LAYER via ;
        RECT 10.670 6.750 10.930 7.010 ;
        RECT 10.670 6.200 10.930 6.460 ;
        RECT 10.670 4.110 10.930 4.370 ;
        RECT 10.670 3.510 10.930 3.820 ;
        RECT 10.670 2.960 10.930 3.220 ;
        RECT 10.670 0.860 10.930 1.120 ;
        RECT 10.670 0.310 10.930 0.570 ;
      LAYER met2 ;
        RECT 10.640 6.760 10.950 7.050 ;
        RECT 10.640 6.720 12.970 6.760 ;
        RECT 10.790 6.580 12.970 6.720 ;
        RECT 10.640 6.330 10.950 6.500 ;
        RECT 10.410 6.150 10.500 6.330 ;
        RECT 10.640 6.170 12.970 6.330 ;
        RECT 10.800 6.150 12.970 6.170 ;
        RECT 0.010 5.730 7.620 5.920 ;
        RECT 10.410 4.240 10.500 4.420 ;
        RECT 10.800 4.400 12.970 4.420 ;
        RECT 10.640 4.240 12.970 4.400 ;
        RECT 7.520 4.210 7.610 4.240 ;
        RECT 7.520 4.100 7.640 4.210 ;
        RECT 10.640 4.070 10.950 4.240 ;
        RECT 10.790 3.850 12.970 3.990 ;
        RECT 10.640 3.810 12.970 3.850 ;
        RECT 10.640 3.520 10.950 3.810 ;
        RECT 10.640 3.480 12.970 3.520 ;
        RECT 10.790 3.340 12.970 3.480 ;
        RECT 7.490 2.950 7.640 3.120 ;
        RECT 10.640 3.090 10.950 3.260 ;
        RECT 10.410 2.910 10.500 3.090 ;
        RECT 10.640 2.930 12.970 3.090 ;
        RECT 10.800 2.910 12.970 2.930 ;
        RECT 0.780 2.510 7.640 2.680 ;
        RECT 10.410 0.990 10.500 1.170 ;
        RECT 10.800 1.150 12.970 1.170 ;
        RECT 10.640 0.990 12.970 1.150 ;
        RECT 10.640 0.820 10.950 0.990 ;
        RECT 10.790 0.600 12.970 0.740 ;
        RECT 10.640 0.560 12.970 0.600 ;
        RECT 10.640 0.270 10.950 0.560 ;
  END
END sky130_hilas_swc4x1BiasCell

MACRO sky130_hilas_FGtrans2x1cell
  CLASS CORE ;
  FOREIGN sky130_hilas_FGtrans2x1cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.570 BY 10.520 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN COLSEL1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 16.850 6.460 17.040 6.520 ;
    END
    PORT
      LAYER met1 ;
        RECT 16.850 0.470 17.040 0.520 ;
    END
  END COLSEL1
  PIN VINJ
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 17.290 0.470 17.450 0.520 ;
    END
  END VINJ
  PIN DRAIN1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 17.730 5.840 17.810 6.020 ;
    END
  END DRAIN1
  PIN DRAIN2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 17.730 0.970 17.810 1.150 ;
    END
  END DRAIN2
  PIN PROG
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 14.080 4.060 14.290 6.520 ;
        RECT 14.080 3.550 14.410 4.060 ;
        RECT 14.080 0.470 14.290 3.550 ;
    END
  END PROG
  PIN RUN
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 13.030 1.990 13.210 6.520 ;
        RECT 12.980 1.650 13.270 1.990 ;
        RECT 13.030 0.470 13.210 1.650 ;
    END
  END RUN
  PIN VIN2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 14.960 3.170 15.150 3.220 ;
        RECT 14.960 2.880 15.270 3.170 ;
        RECT 14.960 1.260 15.150 2.880 ;
        RECT 14.960 0.970 15.250 1.260 ;
        RECT 14.930 0.470 15.160 0.970 ;
    END
  END VIN2
  PIN VIN1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 14.960 6.230 15.170 6.520 ;
        RECT 14.960 5.940 15.280 6.230 ;
        RECT 14.960 4.240 15.170 5.940 ;
        RECT 14.960 3.950 15.280 4.240 ;
        RECT 14.960 3.730 15.170 3.950 ;
    END
  END VIN1
  PIN GATE1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 14.510 5.670 14.700 6.520 ;
        RECT 14.510 5.380 14.810 5.670 ;
        RECT 14.510 3.350 14.700 5.380 ;
        RECT 14.510 3.060 14.810 3.350 ;
        RECT 14.510 1.770 14.700 3.060 ;
        RECT 14.510 1.480 14.820 1.770 ;
        RECT 14.510 0.470 14.700 1.480 ;
    END
  END GATE1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 9.110 3.660 9.340 6.520 ;
        RECT 9.110 3.370 9.440 3.660 ;
        RECT 9.110 0.470 9.340 3.370 ;
    END
  END VGND
  PIN VTUN
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 6.630 0.470 7.050 6.520 ;
    END
  END VTUN
  PIN DRAIN2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 15.340 1.140 15.500 1.160 ;
        RECT 6.290 1.090 15.500 1.140 ;
        RECT 6.290 0.990 15.380 1.090 ;
    END
  END DRAIN2
  PIN DRAIN1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 15.080 6.020 15.400 6.040 ;
        RECT 6.290 5.840 15.400 6.020 ;
    END
  END DRAIN1
  PIN COL1
    PORT
      LAYER met2 ;
        RECT 6.290 3.560 16.450 3.600 ;
        RECT 6.290 3.370 16.460 3.560 ;
    END
  END COL1
  PIN ROW1
    PORT
      LAYER met2 ;
        RECT 15.860 4.480 16.170 4.650 ;
        RECT 6.290 4.320 16.170 4.480 ;
        RECT 6.290 4.290 16.000 4.320 ;
    END
  END ROW1
  PIN ROW2
    PORT
      LAYER met2 ;
        RECT 6.290 2.430 16.010 2.620 ;
    END
  END ROW2
  OBS
      LAYER nwell ;
        RECT 20.800 10.180 22.530 10.520 ;
        RECT 20.780 8.620 22.530 10.180 ;
        RECT 20.780 6.990 22.510 8.620 ;
        RECT 0.010 6.560 2.720 6.600 ;
        RECT 0.000 4.910 2.720 6.560 ;
        RECT 0.000 0.330 2.720 1.980 ;
        RECT 6.870 1.870 7.430 4.290 ;
        RECT 19.260 3.820 22.570 6.990 ;
        RECT 6.630 0.480 7.050 0.550 ;
        RECT 0.010 0.290 2.720 0.330 ;
        RECT 19.260 0.000 22.570 3.170 ;
      LAYER li1 ;
        RECT 21.200 8.790 21.750 9.220 ;
        RECT 21.200 7.060 21.750 7.490 ;
        RECT 20.160 6.360 20.690 6.530 ;
        RECT 21.970 6.260 22.170 6.610 ;
        RECT 21.970 6.230 22.180 6.260 ;
        RECT 2.190 5.430 2.420 6.120 ;
        RECT 14.100 5.920 14.980 6.090 ;
        RECT 15.070 5.970 15.260 6.200 ;
        RECT 14.100 5.530 14.270 5.920 ;
        RECT 18.290 5.780 18.640 5.950 ;
        RECT 19.660 5.780 19.990 5.950 ;
        RECT 13.880 5.360 14.270 5.530 ;
        RECT 14.600 5.530 14.790 5.640 ;
        RECT 14.600 5.410 14.900 5.530 ;
        RECT 14.680 5.360 14.900 5.410 ;
        RECT 18.290 4.990 18.640 5.160 ;
        RECT 19.660 4.990 19.990 5.160 ;
        RECT 12.450 4.570 13.530 4.740 ;
        RECT 13.860 4.570 14.940 4.740 ;
        RECT 15.870 4.570 16.190 4.610 ;
        RECT 15.870 4.380 16.200 4.570 ;
        RECT 15.870 4.350 16.190 4.380 ;
        RECT 9.320 3.630 9.510 3.950 ;
        RECT 9.230 3.540 9.510 3.630 ;
        RECT 9.230 3.400 12.870 3.540 ;
        RECT 9.320 3.360 12.870 3.400 ;
        RECT 9.320 2.940 9.510 3.360 ;
        RECT 13.620 3.210 13.790 3.780 ;
        RECT 14.190 3.630 14.400 4.060 ;
        RECT 15.070 3.980 15.260 4.210 ;
        RECT 18.300 4.200 18.640 4.370 ;
        RECT 19.660 4.200 19.990 4.370 ;
        RECT 20.410 4.280 20.580 5.970 ;
        RECT 21.240 4.370 21.410 5.980 ;
        RECT 21.960 5.650 22.180 6.230 ;
        RECT 21.970 5.640 22.180 5.650 ;
        RECT 21.610 5.470 21.800 5.480 ;
        RECT 21.610 5.180 21.810 5.470 ;
        RECT 21.600 4.850 21.870 5.180 ;
        RECT 21.240 4.180 21.420 4.370 ;
        RECT 14.880 3.780 14.960 3.950 ;
        RECT 14.210 3.610 14.380 3.630 ;
        RECT 13.800 3.180 13.880 3.190 ;
        RECT 14.460 3.180 14.510 3.190 ;
        RECT 13.800 3.140 14.510 3.180 ;
        RECT 13.780 3.100 14.510 3.140 ;
        RECT 13.710 2.980 14.550 3.100 ;
        RECT 14.600 3.090 14.790 3.320 ;
        RECT 14.880 3.040 14.930 3.210 ;
        RECT 15.060 2.910 15.250 3.140 ;
        RECT 15.880 2.880 16.200 2.920 ;
        RECT 15.880 2.690 16.210 2.880 ;
        RECT 15.880 2.660 16.200 2.690 ;
        RECT 18.300 2.620 18.640 2.790 ;
        RECT 19.660 2.620 19.990 2.790 ;
        RECT 12.300 2.250 13.540 2.420 ;
        RECT 13.860 2.250 14.940 2.420 ;
        RECT 13.040 1.930 13.210 1.990 ;
        RECT 13.020 1.720 13.230 1.930 ;
        RECT 18.290 1.830 18.640 2.000 ;
        RECT 19.660 1.830 19.990 2.000 ;
        RECT 13.040 1.650 13.210 1.720 ;
        RECT 14.610 1.630 14.800 1.740 ;
        RECT 13.880 1.620 14.340 1.630 ;
        RECT 13.870 1.470 14.340 1.620 ;
        RECT 14.610 1.510 14.900 1.630 ;
        RECT 13.880 1.460 14.340 1.470 ;
        RECT 14.690 1.460 14.900 1.510 ;
        RECT 2.190 0.770 2.420 1.460 ;
        RECT 14.150 1.120 14.340 1.460 ;
        RECT 15.040 1.120 15.230 1.230 ;
        RECT 14.150 1.000 15.230 1.120 ;
        RECT 18.290 1.040 18.640 1.210 ;
        RECT 19.660 1.040 19.990 1.210 ;
        RECT 20.410 1.020 20.580 2.710 ;
        RECT 21.240 2.620 21.420 2.810 ;
        RECT 21.240 1.010 21.410 2.620 ;
        RECT 21.600 1.810 21.870 2.140 ;
        RECT 21.610 1.520 21.810 1.810 ;
        RECT 21.610 1.510 21.800 1.520 ;
        RECT 21.970 1.340 22.180 1.350 ;
        RECT 14.150 0.940 15.110 1.000 ;
        RECT 21.960 0.760 22.180 1.340 ;
        RECT 21.970 0.730 22.180 0.760 ;
        RECT 20.160 0.460 20.690 0.630 ;
        RECT 21.970 0.380 22.170 0.730 ;
      LAYER mcon ;
        RECT 21.200 8.870 21.470 9.140 ;
        RECT 21.200 7.140 21.470 7.410 ;
        RECT 2.220 5.910 2.390 6.080 ;
        RECT 2.220 5.460 2.390 5.630 ;
        RECT 15.080 6.000 15.250 6.170 ;
        RECT 21.980 6.060 22.150 6.230 ;
        RECT 14.610 5.440 14.780 5.610 ;
        RECT 15.930 4.390 16.100 4.560 ;
        RECT 21.620 5.220 21.800 5.410 ;
        RECT 15.080 4.010 15.250 4.180 ;
        RECT 9.240 3.430 9.410 3.600 ;
        RECT 14.610 3.120 14.780 3.290 ;
        RECT 15.070 2.940 15.240 3.110 ;
        RECT 15.940 2.700 16.110 2.870 ;
        RECT 14.620 1.540 14.790 1.710 ;
        RECT 2.220 1.260 2.390 1.430 ;
        RECT 2.220 0.810 2.390 0.980 ;
        RECT 15.050 1.030 15.220 1.200 ;
        RECT 21.620 1.580 21.800 1.770 ;
        RECT 21.980 0.760 22.150 0.930 ;
      LAYER met1 ;
        RECT 21.140 6.600 21.530 10.190 ;
        RECT 17.290 6.470 17.450 6.520 ;
        RECT 2.180 5.380 2.440 6.170 ;
        RECT 20.090 6.120 20.400 6.560 ;
        RECT 21.610 5.480 21.800 6.930 ;
        RECT 22.050 6.290 22.210 6.930 ;
        RECT 21.940 5.740 22.210 6.290 ;
        RECT 21.940 5.690 22.220 5.740 ;
        RECT 22.050 5.600 22.220 5.690 ;
        RECT 21.610 5.450 21.830 5.480 ;
        RECT 21.590 5.180 21.840 5.450 ;
        RECT 21.600 5.170 21.840 5.180 ;
        RECT 21.600 4.930 21.830 5.170 ;
        RECT 15.860 4.320 16.180 4.640 ;
        RECT 21.210 4.120 21.450 4.500 ;
        RECT 21.640 3.910 21.800 4.930 ;
        RECT 22.050 3.910 22.210 5.600 ;
        RECT 16.550 3.700 16.810 3.760 ;
        RECT 16.450 3.440 16.810 3.700 ;
        RECT 16.450 3.280 16.690 3.440 ;
        RECT 15.870 2.630 16.190 2.950 ;
        RECT 21.210 2.490 21.450 2.870 ;
        RECT 21.640 2.060 21.800 3.080 ;
        RECT 21.600 1.820 21.830 2.060 ;
        RECT 21.600 1.810 21.840 1.820 ;
        RECT 21.590 1.540 21.840 1.810 ;
        RECT 21.610 1.510 21.830 1.540 ;
        RECT 2.180 0.720 2.440 1.510 ;
        RECT 15.460 0.970 15.470 0.980 ;
        RECT 20.090 0.430 20.400 0.870 ;
        RECT 21.610 0.060 21.800 1.510 ;
        RECT 22.050 1.390 22.210 3.080 ;
        RECT 22.050 1.300 22.220 1.390 ;
        RECT 21.940 1.250 22.220 1.300 ;
        RECT 21.940 0.700 22.210 1.250 ;
        RECT 22.050 0.060 22.210 0.700 ;
      LAYER via ;
        RECT 20.120 6.150 20.380 6.410 ;
        RECT 15.890 4.350 16.150 4.610 ;
        RECT 16.550 3.470 16.810 3.730 ;
        RECT 15.900 2.660 16.160 2.920 ;
        RECT 20.120 0.580 20.380 0.840 ;
      LAYER met2 ;
        RECT 20.090 6.440 20.400 6.450 ;
        RECT 20.090 6.260 22.570 6.440 ;
        RECT 20.090 6.120 20.400 6.260 ;
        RECT 16.520 3.470 16.840 3.730 ;
        RECT 15.870 2.630 16.180 2.960 ;
        RECT 20.090 0.730 20.400 0.870 ;
        RECT 20.090 0.550 22.570 0.730 ;
        RECT 20.090 0.540 20.400 0.550 ;
  END
END sky130_hilas_FGtrans2x1cell

MACRO sky130_hilas_capacitorSize01
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.090 BY 7.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 10.060 2.380 10.420 2.660 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.020 2.370 0.290 2.650 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 0.000 4.850 10.420 5.030 ;
        RECT 0.000 4.420 10.420 4.600 ;
        RECT 0.030 3.420 10.420 3.600 ;
        RECT 8.510 3.170 10.420 3.180 ;
        RECT 0.030 3.080 10.420 3.170 ;
        RECT 0.030 2.990 10.460 3.080 ;
        RECT 0.600 2.670 0.970 2.990 ;
        RECT 10.090 2.680 10.460 2.990 ;
        RECT 0.030 1.840 10.420 2.010 ;
        RECT 0.030 1.420 10.420 1.590 ;
        RECT 0.030 0.440 10.420 0.610 ;
        RECT 0.030 0.000 10.420 0.170 ;
      LAYER via2 ;
        RECT 0.650 2.730 0.930 3.010 ;
        RECT 10.140 2.740 10.420 3.020 ;
      LAYER met3 ;
        RECT 5.890 7.840 8.710 7.870 ;
        RECT 0.380 2.470 1.170 3.220 ;
        RECT 5.890 2.060 13.090 7.840 ;
        RECT 8.680 2.040 13.090 2.060 ;
      LAYER via3 ;
        RECT 0.570 2.620 1.000 3.100 ;
        RECT 10.060 2.630 10.490 3.110 ;
      LAYER met4 ;
        RECT 0.470 2.770 1.130 3.190 ;
        RECT 6.780 3.140 9.820 3.610 ;
        RECT 1.160 2.770 2.170 2.780 ;
        RECT 0.450 2.270 3.800 2.770 ;
        RECT 9.960 2.540 10.620 3.200 ;
        RECT 0.450 2.260 1.520 2.270 ;
        RECT 3.160 1.150 3.790 2.270 ;
        RECT 3.160 0.850 5.310 1.150 ;
        RECT 3.490 0.840 5.310 0.850 ;
  END
END sky130_hilas_capacitorSize01

MACRO sky130_hilas_Tgate4Double01
  CLASS CORE ;
  FOREIGN sky130_hilas_Tgate4Double01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.710 BY 6.950 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.740 6.460 0.940 6.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.570 0.450 6.760 0.490 ;
    END
  END VGND
  PIN INPUT1_1
    PORT
      LAYER met2 ;
        RECT 0.000 6.190 0.050 6.390 ;
    END
  END INPUT1_1
  PIN SELECT1
    PORT
      LAYER met2 ;
        RECT 0.000 5.210 0.060 5.410 ;
    END
  END SELECT1
  PIN SELECT2
    PORT
      LAYER met2 ;
        RECT 0.000 4.560 0.060 4.760 ;
    END
  END SELECT2
  PIN INPUT2_2
    PORT
      LAYER met2 ;
        RECT 0.000 4.060 0.050 4.260 ;
    END
  END INPUT2_2
  PIN INPUT1_2
    PORT
      LAYER met2 ;
        RECT 0.000 3.580 0.050 3.780 ;
    END
  END INPUT1_2
  PIN SELECT3
    PORT
      LAYER met2 ;
        RECT 0.000 2.190 0.060 2.390 ;
    END
  END SELECT3
  PIN INPUT2_3
    PORT
      LAYER met2 ;
        RECT 0.000 2.690 0.050 2.890 ;
    END
  END INPUT2_3
  PIN SELECT4
    PORT
      LAYER met2 ;
        RECT 0.000 1.540 0.060 1.740 ;
    END
  END SELECT4
  PIN INPUT2_4
    PORT
      LAYER met2 ;
        RECT 0.000 1.040 0.050 1.240 ;
    END
  END INPUT2_4
  PIN INPUT1_4
    PORT
      LAYER met2 ;
        RECT 0.000 0.560 0.050 0.760 ;
    END
  END INPUT1_4
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 6.570 6.460 6.760 6.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.740 0.450 0.940 0.490 ;
    END
  END VPWR
  PIN OUTPUT4
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 7.020 1.560 7.080 1.740 ;
        RECT 2.630 1.410 8.400 1.560 ;
        RECT 2.630 1.360 8.610 1.410 ;
        RECT 5.220 1.090 5.530 1.360 ;
        RECT 8.300 1.080 8.610 1.360 ;
    END
  END OUTPUT4
  PIN OUTPUT3
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 5.220 2.570 5.530 2.840 ;
        RECT 8.300 2.570 8.610 2.850 ;
        RECT 2.630 2.520 8.610 2.570 ;
        RECT 2.630 2.370 8.400 2.520 ;
        RECT 7.020 2.190 7.080 2.370 ;
    END
  END OUTPUT3
  PIN OUTPUT2
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 7.020 4.580 7.080 4.760 ;
        RECT 2.630 4.430 8.400 4.580 ;
        RECT 2.630 4.380 8.610 4.430 ;
        RECT 5.220 4.110 5.530 4.380 ;
        RECT 8.300 4.100 8.610 4.380 ;
    END
  END OUTPUT2
  PIN OUTPUT1
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 5.220 5.590 5.530 5.860 ;
        RECT 8.300 5.590 8.610 5.870 ;
        RECT 2.630 5.540 8.610 5.590 ;
        RECT 2.630 5.390 8.400 5.540 ;
        RECT 7.010 5.210 7.080 5.390 ;
    END
  END OUTPUT1
  PIN INPUT2_1
    PORT
      LAYER met2 ;
        RECT 0.000 5.710 0.050 5.910 ;
    END
  END INPUT2_1
  PIN INPUT1_3
    PORT
      LAYER met2 ;
        RECT 0.000 3.170 0.050 3.370 ;
    END
  END INPUT1_3
  OBS
      LAYER nwell ;
        RECT 2.750 5.280 6.220 6.800 ;
        RECT 2.750 2.260 6.220 4.690 ;
        RECT 2.750 0.150 6.220 1.670 ;
      LAYER li1 ;
        RECT 2.960 6.520 3.170 6.950 ;
        RECT 2.980 6.500 3.150 6.520 ;
        RECT 3.480 6.380 3.670 6.490 ;
        RECT 3.480 6.260 3.900 6.380 ;
        RECT 3.380 6.210 3.900 6.260 ;
        RECT 4.250 6.210 8.470 6.390 ;
        RECT 8.850 6.220 9.200 6.390 ;
        RECT 9.300 6.380 9.490 6.490 ;
        RECT 9.300 6.260 9.630 6.380 ;
        RECT 3.380 6.130 3.570 6.210 ;
        RECT 3.360 6.100 3.570 6.130 ;
        RECT 3.350 6.090 3.570 6.100 ;
        RECT 3.230 6.040 3.570 6.090 ;
        RECT 3.100 6.010 3.570 6.040 ;
        RECT 3.060 5.980 3.570 6.010 ;
        RECT 3.880 6.150 4.200 6.190 ;
        RECT 3.060 5.920 3.550 5.980 ;
        RECT 3.880 5.960 4.210 6.150 ;
        RECT 4.740 6.090 5.070 6.210 ;
        RECT 6.800 6.150 7.120 6.190 ;
        RECT 9.380 6.180 9.630 6.260 ;
        RECT 4.450 5.990 4.640 6.080 ;
        RECT 3.880 5.930 4.200 5.960 ;
        RECT 3.060 5.870 3.400 5.920 ;
        RECT 3.060 5.850 3.320 5.870 ;
        RECT 4.340 5.850 4.640 5.990 ;
        RECT 5.900 5.870 6.090 6.100 ;
        RECT 6.800 5.960 7.130 6.150 ;
        RECT 6.800 5.930 7.120 5.960 ;
        RECT 7.610 5.870 7.800 6.090 ;
        RECT 7.510 5.860 7.800 5.870 ;
        RECT 3.060 5.830 3.290 5.850 ;
        RECT 3.060 5.790 3.270 5.830 ;
        RECT 3.060 5.510 3.230 5.790 ;
        RECT 3.740 5.750 3.920 5.790 ;
        RECT 3.570 5.580 3.920 5.750 ;
        RECT 4.340 5.500 4.510 5.850 ;
        RECT 5.120 5.820 5.290 5.840 ;
        RECT 5.120 5.780 5.550 5.820 ;
        RECT 5.120 5.590 5.560 5.780 ;
        RECT 5.120 5.560 5.550 5.590 ;
        RECT 5.120 5.540 5.290 5.560 ;
        RECT 5.810 5.500 5.980 5.850 ;
        RECT 6.770 5.500 6.940 5.800 ;
        RECT 7.510 5.490 7.680 5.860 ;
        RECT 8.230 5.830 8.400 5.840 ;
        RECT 8.230 5.790 8.630 5.830 ;
        RECT 8.230 5.600 8.640 5.790 ;
        RECT 8.840 5.760 9.030 5.870 ;
        RECT 8.840 5.640 9.180 5.760 ;
        RECT 8.230 5.570 8.630 5.600 ;
        RECT 8.890 5.590 9.180 5.640 ;
        RECT 8.230 5.540 8.400 5.570 ;
        RECT 9.460 5.500 9.630 6.180 ;
        RECT 3.060 4.180 3.230 4.460 ;
        RECT 3.570 4.220 3.920 4.390 ;
        RECT 3.740 4.180 3.920 4.220 ;
        RECT 3.060 4.140 3.270 4.180 ;
        RECT 3.060 4.120 3.290 4.140 ;
        RECT 4.340 4.120 4.510 4.470 ;
        RECT 5.120 4.410 5.290 4.430 ;
        RECT 5.120 4.380 5.550 4.410 ;
        RECT 5.120 4.190 5.560 4.380 ;
        RECT 5.120 4.150 5.550 4.190 ;
        RECT 5.120 4.130 5.290 4.150 ;
        RECT 5.810 4.120 5.980 4.470 ;
        RECT 6.770 4.170 6.940 4.470 ;
        RECT 3.060 4.100 3.320 4.120 ;
        RECT 3.060 4.050 3.400 4.100 ;
        RECT 3.060 3.990 3.550 4.050 ;
        RECT 3.880 4.010 4.200 4.040 ;
        RECT 3.060 3.960 3.570 3.990 ;
        RECT 3.100 3.930 3.570 3.960 ;
        RECT 2.960 3.500 3.170 3.930 ;
        RECT 3.230 3.880 3.570 3.930 ;
        RECT 3.350 3.870 3.570 3.880 ;
        RECT 3.360 3.840 3.570 3.870 ;
        RECT 3.380 3.760 3.570 3.840 ;
        RECT 3.880 3.820 4.210 4.010 ;
        RECT 4.340 3.980 4.640 4.120 ;
        RECT 7.510 4.110 7.680 4.480 ;
        RECT 8.230 4.400 8.400 4.430 ;
        RECT 8.230 4.370 8.630 4.400 ;
        RECT 8.230 4.180 8.640 4.370 ;
        RECT 8.890 4.330 9.180 4.380 ;
        RECT 8.840 4.210 9.180 4.330 ;
        RECT 8.230 4.140 8.630 4.180 ;
        RECT 8.230 4.130 8.400 4.140 ;
        RECT 7.510 4.100 7.800 4.110 ;
        RECT 8.840 4.100 9.030 4.210 ;
        RECT 4.450 3.890 4.640 3.980 ;
        RECT 3.880 3.780 4.200 3.820 ;
        RECT 4.740 3.760 5.070 3.880 ;
        RECT 5.900 3.870 6.090 4.100 ;
        RECT 6.800 4.010 7.120 4.040 ;
        RECT 6.800 3.820 7.130 4.010 ;
        RECT 7.610 3.880 7.800 4.100 ;
        RECT 6.800 3.780 7.120 3.820 ;
        RECT 9.460 3.790 9.630 4.470 ;
        RECT 3.380 3.710 3.900 3.760 ;
        RECT 3.480 3.590 3.900 3.710 ;
        RECT 2.980 3.480 3.150 3.500 ;
        RECT 3.480 3.480 3.670 3.590 ;
        RECT 4.250 3.580 8.470 3.760 ;
        RECT 8.850 3.580 9.200 3.750 ;
        RECT 9.380 3.710 9.630 3.790 ;
        RECT 9.300 3.590 9.630 3.710 ;
        RECT 9.300 3.480 9.490 3.590 ;
        RECT 2.980 3.450 3.150 3.470 ;
        RECT 2.960 3.020 3.170 3.450 ;
        RECT 3.480 3.360 3.670 3.470 ;
        RECT 3.480 3.240 3.900 3.360 ;
        RECT 3.380 3.190 3.900 3.240 ;
        RECT 4.250 3.190 8.470 3.370 ;
        RECT 8.850 3.200 9.200 3.370 ;
        RECT 9.300 3.360 9.490 3.470 ;
        RECT 9.300 3.240 9.630 3.360 ;
        RECT 3.380 3.110 3.570 3.190 ;
        RECT 3.360 3.080 3.570 3.110 ;
        RECT 3.350 3.070 3.570 3.080 ;
        RECT 3.230 3.020 3.570 3.070 ;
        RECT 3.100 2.990 3.570 3.020 ;
        RECT 3.060 2.960 3.570 2.990 ;
        RECT 3.880 3.130 4.200 3.170 ;
        RECT 3.060 2.900 3.550 2.960 ;
        RECT 3.880 2.940 4.210 3.130 ;
        RECT 4.740 3.070 5.070 3.190 ;
        RECT 6.800 3.130 7.120 3.170 ;
        RECT 9.380 3.160 9.630 3.240 ;
        RECT 4.450 2.970 4.640 3.060 ;
        RECT 3.880 2.910 4.200 2.940 ;
        RECT 3.060 2.850 3.400 2.900 ;
        RECT 3.060 2.830 3.320 2.850 ;
        RECT 4.340 2.830 4.640 2.970 ;
        RECT 5.900 2.850 6.090 3.080 ;
        RECT 6.800 2.940 7.130 3.130 ;
        RECT 6.800 2.910 7.120 2.940 ;
        RECT 7.610 2.850 7.800 3.070 ;
        RECT 7.510 2.840 7.800 2.850 ;
        RECT 3.060 2.810 3.290 2.830 ;
        RECT 3.060 2.770 3.270 2.810 ;
        RECT 3.060 2.490 3.230 2.770 ;
        RECT 3.740 2.730 3.920 2.770 ;
        RECT 3.570 2.560 3.920 2.730 ;
        RECT 4.340 2.480 4.510 2.830 ;
        RECT 5.120 2.800 5.290 2.820 ;
        RECT 5.120 2.760 5.550 2.800 ;
        RECT 5.120 2.570 5.560 2.760 ;
        RECT 5.120 2.540 5.550 2.570 ;
        RECT 5.120 2.520 5.290 2.540 ;
        RECT 5.810 2.480 5.980 2.830 ;
        RECT 6.770 2.480 6.940 2.780 ;
        RECT 7.510 2.470 7.680 2.840 ;
        RECT 8.230 2.810 8.400 2.820 ;
        RECT 8.230 2.770 8.630 2.810 ;
        RECT 8.230 2.580 8.640 2.770 ;
        RECT 8.840 2.740 9.030 2.850 ;
        RECT 8.840 2.620 9.180 2.740 ;
        RECT 8.230 2.550 8.630 2.580 ;
        RECT 8.890 2.570 9.180 2.620 ;
        RECT 8.230 2.520 8.400 2.550 ;
        RECT 9.460 2.480 9.630 3.160 ;
        RECT 3.060 1.160 3.230 1.440 ;
        RECT 3.570 1.200 3.920 1.370 ;
        RECT 3.740 1.160 3.920 1.200 ;
        RECT 3.060 1.120 3.270 1.160 ;
        RECT 3.060 1.100 3.290 1.120 ;
        RECT 4.340 1.100 4.510 1.450 ;
        RECT 5.120 1.390 5.290 1.410 ;
        RECT 5.120 1.360 5.550 1.390 ;
        RECT 5.120 1.170 5.560 1.360 ;
        RECT 5.120 1.130 5.550 1.170 ;
        RECT 5.120 1.110 5.290 1.130 ;
        RECT 5.810 1.100 5.980 1.450 ;
        RECT 6.770 1.150 6.940 1.450 ;
        RECT 3.060 1.080 3.320 1.100 ;
        RECT 3.060 1.030 3.400 1.080 ;
        RECT 3.060 0.970 3.550 1.030 ;
        RECT 3.880 0.990 4.200 1.020 ;
        RECT 3.060 0.940 3.570 0.970 ;
        RECT 3.100 0.910 3.570 0.940 ;
        RECT 3.230 0.860 3.570 0.910 ;
        RECT 3.350 0.850 3.570 0.860 ;
        RECT 3.360 0.820 3.570 0.850 ;
        RECT 3.380 0.740 3.570 0.820 ;
        RECT 3.880 0.800 4.210 0.990 ;
        RECT 4.340 0.960 4.640 1.100 ;
        RECT 7.510 1.090 7.680 1.460 ;
        RECT 8.230 1.380 8.400 1.410 ;
        RECT 8.230 1.350 8.630 1.380 ;
        RECT 8.230 1.160 8.640 1.350 ;
        RECT 8.890 1.310 9.180 1.360 ;
        RECT 8.840 1.190 9.180 1.310 ;
        RECT 8.230 1.120 8.630 1.160 ;
        RECT 8.230 1.110 8.400 1.120 ;
        RECT 7.510 1.080 7.800 1.090 ;
        RECT 8.840 1.080 9.030 1.190 ;
        RECT 4.450 0.870 4.640 0.960 ;
        RECT 3.880 0.760 4.200 0.800 ;
        RECT 4.740 0.740 5.070 0.860 ;
        RECT 5.900 0.850 6.090 1.080 ;
        RECT 6.800 0.990 7.120 1.020 ;
        RECT 6.800 0.800 7.130 0.990 ;
        RECT 7.610 0.860 7.800 1.080 ;
        RECT 6.800 0.760 7.120 0.800 ;
        RECT 9.460 0.770 9.630 1.450 ;
        RECT 3.380 0.690 3.900 0.740 ;
        RECT 3.480 0.570 3.900 0.690 ;
        RECT 3.480 0.460 3.670 0.570 ;
        RECT 4.250 0.560 8.470 0.740 ;
        RECT 8.850 0.560 9.200 0.730 ;
        RECT 9.380 0.690 9.630 0.770 ;
        RECT 9.300 0.570 9.630 0.690 ;
        RECT 9.300 0.460 9.490 0.570 ;
        RECT 2.980 0.430 3.150 0.450 ;
        RECT 2.960 0.000 3.170 0.430 ;
      LAYER mcon ;
        RECT 3.490 6.290 3.660 6.460 ;
        RECT 9.310 6.290 9.480 6.460 ;
        RECT 3.940 5.970 4.110 6.140 ;
        RECT 4.460 5.880 4.630 6.050 ;
        RECT 5.910 5.900 6.080 6.070 ;
        RECT 6.860 5.970 7.030 6.140 ;
        RECT 7.620 5.890 7.790 6.060 ;
        RECT 5.290 5.600 5.460 5.770 ;
        RECT 8.370 5.610 8.540 5.780 ;
        RECT 8.850 5.670 9.020 5.840 ;
        RECT 5.290 4.200 5.460 4.370 ;
        RECT 8.370 4.190 8.540 4.360 ;
        RECT 8.850 4.130 9.020 4.300 ;
        RECT 3.940 3.830 4.110 4.000 ;
        RECT 4.460 3.920 4.630 4.090 ;
        RECT 5.910 3.900 6.080 4.070 ;
        RECT 6.860 3.830 7.030 4.000 ;
        RECT 7.620 3.910 7.790 4.080 ;
        RECT 3.490 3.510 3.660 3.680 ;
        RECT 9.310 3.510 9.480 3.680 ;
        RECT 2.980 3.300 3.150 3.470 ;
        RECT 3.490 3.270 3.660 3.440 ;
        RECT 9.310 3.270 9.480 3.440 ;
        RECT 3.940 2.950 4.110 3.120 ;
        RECT 4.460 2.860 4.630 3.030 ;
        RECT 5.910 2.880 6.080 3.050 ;
        RECT 6.860 2.950 7.030 3.120 ;
        RECT 7.620 2.870 7.790 3.040 ;
        RECT 5.290 2.580 5.460 2.750 ;
        RECT 8.370 2.590 8.540 2.760 ;
        RECT 8.850 2.650 9.020 2.820 ;
        RECT 5.290 1.180 5.460 1.350 ;
        RECT 8.370 1.170 8.540 1.340 ;
        RECT 8.850 1.110 9.020 1.280 ;
        RECT 3.940 0.810 4.110 0.980 ;
        RECT 4.460 0.900 4.630 1.070 ;
        RECT 5.910 0.880 6.080 1.050 ;
        RECT 6.860 0.810 7.030 0.980 ;
        RECT 7.620 0.890 7.790 1.060 ;
        RECT 3.490 0.490 3.660 0.660 ;
        RECT 9.310 0.490 9.480 0.660 ;
        RECT 2.980 0.280 3.150 0.450 ;
      LAYER met1 ;
        RECT 2.960 6.790 3.180 6.950 ;
        RECT 2.960 6.730 3.300 6.790 ;
        RECT 2.950 6.470 3.300 6.730 ;
        RECT 3.370 6.520 3.570 6.800 ;
        RECT 2.950 6.440 3.180 6.470 ;
        RECT 3.370 6.230 3.690 6.520 ;
        RECT 4.430 6.390 4.690 6.710 ;
        RECT 5.850 6.400 6.110 6.720 ;
        RECT 7.600 6.420 7.860 6.740 ;
        RECT 8.640 6.560 8.900 6.730 ;
        RECT 8.640 6.410 8.910 6.560 ;
        RECT 3.370 5.280 3.570 6.230 ;
        RECT 3.870 5.900 4.190 6.220 ;
        RECT 4.350 6.110 4.520 6.290 ;
        RECT 5.800 6.130 5.970 6.310 ;
        RECT 4.350 6.020 4.660 6.110 ;
        RECT 5.800 6.040 6.110 6.130 ;
        RECT 4.430 5.820 4.660 6.020 ;
        RECT 5.220 5.530 5.540 5.850 ;
        RECT 5.880 5.840 6.110 6.040 ;
        RECT 6.790 5.900 7.110 6.220 ;
        RECT 7.520 6.120 7.690 6.350 ;
        RECT 7.520 6.010 7.820 6.120 ;
        RECT 7.590 5.830 7.820 6.010 ;
        RECT 8.720 5.900 8.910 6.410 ;
        RECT 9.200 6.520 9.390 6.800 ;
        RECT 9.200 6.230 9.510 6.520 ;
        RECT 8.300 5.540 8.620 5.860 ;
        RECT 8.720 5.810 9.050 5.900 ;
        RECT 8.820 5.610 9.050 5.810 ;
        RECT 9.200 5.280 9.390 6.230 ;
        RECT 2.960 3.770 3.180 3.930 ;
        RECT 2.960 3.710 3.300 3.770 ;
        RECT 2.950 3.240 3.300 3.710 ;
        RECT 2.960 3.180 3.300 3.240 ;
        RECT 3.370 3.740 3.570 4.690 ;
        RECT 3.870 3.750 4.190 4.070 ;
        RECT 4.430 3.950 4.660 4.150 ;
        RECT 5.220 4.120 5.540 4.440 ;
        RECT 4.350 3.860 4.660 3.950 ;
        RECT 5.880 3.930 6.110 4.130 ;
        RECT 3.370 3.210 3.690 3.740 ;
        RECT 4.350 3.690 4.520 3.860 ;
        RECT 5.800 3.840 6.110 3.930 ;
        RECT 5.800 3.700 5.970 3.840 ;
        RECT 6.790 3.750 7.110 4.070 ;
        RECT 7.590 3.960 7.820 4.140 ;
        RECT 8.300 4.110 8.620 4.430 ;
        RECT 8.820 4.160 9.050 4.360 ;
        RECT 7.520 3.850 7.820 3.960 ;
        RECT 8.720 4.070 9.050 4.160 ;
        RECT 7.520 3.720 7.690 3.850 ;
        RECT 4.350 3.680 4.690 3.690 ;
        RECT 4.430 3.270 4.690 3.680 ;
        RECT 5.800 3.660 6.110 3.700 ;
        RECT 5.850 3.290 6.110 3.660 ;
        RECT 7.520 3.620 7.860 3.720 ;
        RECT 8.720 3.710 8.910 4.070 ;
        RECT 7.600 3.330 7.860 3.620 ;
        RECT 4.350 3.260 4.690 3.270 ;
        RECT 2.960 3.020 3.180 3.180 ;
        RECT 3.370 2.260 3.570 3.210 ;
        RECT 3.870 2.880 4.190 3.200 ;
        RECT 4.350 3.090 4.520 3.260 ;
        RECT 5.800 3.250 6.110 3.290 ;
        RECT 5.800 3.110 5.970 3.250 ;
        RECT 7.520 3.230 7.860 3.330 ;
        RECT 8.640 3.240 8.910 3.710 ;
        RECT 4.350 3.000 4.660 3.090 ;
        RECT 5.800 3.020 6.110 3.110 ;
        RECT 4.430 2.800 4.660 3.000 ;
        RECT 5.220 2.510 5.540 2.830 ;
        RECT 5.880 2.820 6.110 3.020 ;
        RECT 6.790 2.880 7.110 3.200 ;
        RECT 7.520 3.100 7.690 3.230 ;
        RECT 7.520 2.990 7.820 3.100 ;
        RECT 7.590 2.810 7.820 2.990 ;
        RECT 8.720 2.880 8.910 3.240 ;
        RECT 9.200 3.740 9.390 4.690 ;
        RECT 9.200 3.210 9.510 3.740 ;
        RECT 8.300 2.520 8.620 2.840 ;
        RECT 8.720 2.790 9.050 2.880 ;
        RECT 8.820 2.590 9.050 2.790 ;
        RECT 9.200 2.260 9.390 3.210 ;
        RECT 3.370 0.720 3.570 1.670 ;
        RECT 3.870 0.730 4.190 1.050 ;
        RECT 4.430 0.930 4.660 1.130 ;
        RECT 5.220 1.100 5.540 1.420 ;
        RECT 4.350 0.840 4.660 0.930 ;
        RECT 5.880 0.910 6.110 1.110 ;
        RECT 2.950 0.480 3.180 0.510 ;
        RECT 2.950 0.220 3.300 0.480 ;
        RECT 2.960 0.160 3.300 0.220 ;
        RECT 3.370 0.430 3.690 0.720 ;
        RECT 4.350 0.660 4.520 0.840 ;
        RECT 5.800 0.820 6.110 0.910 ;
        RECT 5.800 0.640 5.970 0.820 ;
        RECT 6.790 0.730 7.110 1.050 ;
        RECT 7.590 0.940 7.820 1.120 ;
        RECT 8.300 1.090 8.620 1.410 ;
        RECT 8.820 1.140 9.050 1.340 ;
        RECT 7.520 0.830 7.820 0.940 ;
        RECT 8.720 1.050 9.050 1.140 ;
        RECT 7.520 0.600 7.690 0.830 ;
        RECT 2.960 0.000 3.180 0.160 ;
        RECT 3.370 0.150 3.570 0.430 ;
        RECT 4.430 0.240 4.690 0.560 ;
        RECT 5.850 0.230 6.110 0.550 ;
        RECT 8.720 0.540 8.910 1.050 ;
        RECT 7.600 0.210 7.860 0.530 ;
        RECT 8.640 0.390 8.910 0.540 ;
        RECT 9.200 0.720 9.390 1.670 ;
        RECT 9.200 0.430 9.510 0.720 ;
        RECT 8.640 0.220 8.900 0.390 ;
        RECT 9.200 0.150 9.390 0.430 ;
      LAYER via ;
        RECT 3.040 6.500 3.300 6.760 ;
        RECT 4.430 6.420 4.690 6.680 ;
        RECT 5.850 6.430 6.110 6.690 ;
        RECT 7.600 6.450 7.860 6.710 ;
        RECT 8.640 6.440 8.900 6.700 ;
        RECT 3.900 5.930 4.160 6.190 ;
        RECT 6.820 5.930 7.080 6.190 ;
        RECT 5.250 5.560 5.510 5.820 ;
        RECT 8.330 5.570 8.590 5.830 ;
        RECT 3.040 3.480 3.300 3.740 ;
        RECT 3.040 3.210 3.300 3.470 ;
        RECT 5.250 4.150 5.510 4.410 ;
        RECT 3.900 3.780 4.160 4.040 ;
        RECT 8.330 4.140 8.590 4.400 ;
        RECT 6.820 3.780 7.080 4.040 ;
        RECT 4.430 3.290 4.690 3.660 ;
        RECT 5.850 3.280 6.110 3.670 ;
        RECT 3.900 2.910 4.160 3.170 ;
        RECT 7.600 3.260 7.860 3.690 ;
        RECT 8.640 3.270 8.900 3.680 ;
        RECT 6.820 2.910 7.080 3.170 ;
        RECT 5.250 2.540 5.510 2.800 ;
        RECT 8.330 2.550 8.590 2.810 ;
        RECT 5.250 1.130 5.510 1.390 ;
        RECT 3.900 0.760 4.160 1.020 ;
        RECT 8.330 1.120 8.590 1.380 ;
        RECT 3.040 0.190 3.300 0.450 ;
        RECT 6.820 0.760 7.080 1.020 ;
        RECT 4.430 0.270 4.690 0.530 ;
        RECT 5.850 0.260 6.110 0.520 ;
        RECT 7.600 0.240 7.860 0.500 ;
        RECT 8.640 0.250 8.900 0.510 ;
      LAYER met2 ;
        RECT 3.010 6.570 3.330 6.760 ;
        RECT 4.400 6.570 4.720 6.680 ;
        RECT 5.820 6.570 6.140 6.690 ;
        RECT 7.570 6.570 7.890 6.710 ;
        RECT 8.610 6.570 8.930 6.700 ;
        RECT 2.630 6.500 3.330 6.570 ;
        RECT 2.630 6.370 3.240 6.500 ;
        RECT 4.330 6.370 9.710 6.570 ;
        RECT 3.870 6.070 4.180 6.230 ;
        RECT 6.790 6.070 7.100 6.230 ;
        RECT 2.630 5.900 7.100 6.070 ;
        RECT 2.630 5.870 7.000 5.900 ;
        RECT 2.630 4.070 7.000 4.100 ;
        RECT 2.630 3.900 7.100 4.070 ;
        RECT 3.870 3.740 4.180 3.900 ;
        RECT 6.790 3.740 7.100 3.900 ;
        RECT 3.010 3.600 3.330 3.740 ;
        RECT 4.400 3.600 4.720 3.660 ;
        RECT 5.820 3.600 6.140 3.670 ;
        RECT 7.570 3.600 7.890 3.690 ;
        RECT 8.610 3.600 8.930 3.680 ;
        RECT 2.630 3.480 3.330 3.600 ;
        RECT 2.630 3.470 3.240 3.480 ;
        RECT 2.630 3.350 3.330 3.470 ;
        RECT 4.330 3.350 9.710 3.600 ;
        RECT 3.010 3.210 3.330 3.350 ;
        RECT 4.400 3.290 4.720 3.350 ;
        RECT 5.820 3.280 6.140 3.350 ;
        RECT 7.570 3.260 7.890 3.350 ;
        RECT 8.610 3.270 8.930 3.350 ;
        RECT 3.870 3.050 4.180 3.210 ;
        RECT 6.790 3.050 7.100 3.210 ;
        RECT 2.630 2.880 7.100 3.050 ;
        RECT 2.630 2.850 7.000 2.880 ;
        RECT 2.630 1.050 7.000 1.080 ;
        RECT 2.630 0.880 7.100 1.050 ;
        RECT 3.870 0.720 4.180 0.880 ;
        RECT 6.790 0.720 7.100 0.880 ;
        RECT 2.630 0.450 3.240 0.580 ;
        RECT 2.630 0.380 3.330 0.450 ;
        RECT 4.330 0.380 9.710 0.580 ;
        RECT 3.010 0.190 3.330 0.380 ;
        RECT 4.400 0.270 4.720 0.380 ;
        RECT 5.820 0.260 6.140 0.380 ;
        RECT 7.570 0.240 7.890 0.380 ;
        RECT 8.610 0.250 8.930 0.380 ;
  END
END sky130_hilas_Tgate4Double01

MACRO sky130_hilas_cellAttempt01
  CLASS CORE ;
  FOREIGN sky130_hilas_cellAttempt01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.240 BY 10.900 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 0.350 0.410 0.750 6.910 ;
    END
  END VTUN
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 9.550 6.630 9.710 6.680 ;
    END
  END VINJ
  PIN COLSEL1
    PORT
      LAYER met1 ;
        RECT 9.110 6.630 9.300 6.680 ;
    END
  END COLSEL1
  PIN COL1
    PORT
      LAYER met1 ;
        RECT 8.740 6.640 8.900 6.680 ;
    END
  END COL1
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT 4.400 6.580 4.780 6.910 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.400 0.410 4.780 1.010 ;
    END
  END GATE1
  PIN ROW4
    PORT
      LAYER met2 ;
        RECT 0.000 1.400 7.620 1.580 ;
    END
  END ROW4
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 2.750 2.190 3.070 2.200 ;
        RECT 6.680 2.190 7.000 2.250 ;
        RECT 2.750 2.010 7.000 2.190 ;
        RECT 2.750 1.940 3.070 2.010 ;
        RECT 6.680 1.960 7.000 2.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.720 5.520 6.960 6.910 ;
        RECT 6.700 4.860 6.970 5.520 ;
        RECT 6.720 2.270 6.960 4.860 ;
        RECT 6.710 1.950 6.970 2.270 ;
        RECT 6.720 0.410 6.960 1.950 ;
      LAYER via ;
        RECT 6.710 1.980 6.970 2.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.790 5.500 3.030 6.910 ;
        RECT 2.780 4.840 3.040 5.500 ;
        RECT 2.790 2.230 3.030 4.840 ;
        RECT 2.780 1.910 3.040 2.230 ;
        RECT 2.790 0.410 3.030 1.910 ;
      LAYER via ;
        RECT 2.780 1.940 3.040 2.200 ;
    END
  END VGND
  PIN DRAIN4
    PORT
      LAYER met2 ;
        RECT 0.000 0.980 7.600 1.150 ;
    END
  END DRAIN4
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 0.000 6.170 7.630 6.350 ;
    END
  END DRAIN1
  PIN ROW1
    PORT
      LAYER met2 ;
        RECT 0.000 5.730 7.630 5.910 ;
    END
  END ROW1
  PIN ROW3
    PORT
      LAYER met2 ;
        RECT 0.000 2.500 7.630 2.680 ;
    END
  END ROW3
  PIN DRAIN3
    PORT
      LAYER met2 ;
        RECT 0.000 2.930 7.620 3.110 ;
    END
  END DRAIN3
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 0.000 4.200 7.630 4.380 ;
    END
  END DRAIN2
  PIN ROW2
    PORT
      LAYER met2 ;
        RECT 0.000 4.630 7.630 4.810 ;
    END
  END ROW2
  OBS
      LAYER nwell ;
        RECT 14.510 10.850 16.240 10.900 ;
        RECT 0.000 5.570 0.070 5.750 ;
        RECT 10.400 5.410 12.960 7.320 ;
        RECT 0.570 5.220 1.160 5.330 ;
        RECT 4.310 5.160 5.420 5.390 ;
        RECT 8.950 3.730 9.300 3.740 ;
        RECT 8.950 3.570 9.120 3.730 ;
        RECT 9.290 3.570 9.300 3.730 ;
        RECT 0.570 1.940 1.160 2.130 ;
        RECT 4.310 1.920 5.420 2.190 ;
        RECT 10.400 2.170 12.960 5.140 ;
        RECT 13.320 4.410 16.240 10.850 ;
        RECT 18.510 7.320 20.240 9.160 ;
        RECT 13.320 4.360 15.550 4.410 ;
        RECT 10.400 0.000 12.960 1.910 ;
      LAYER li1 ;
        RECT 14.900 7.840 15.450 8.270 ;
        RECT 18.930 7.770 19.480 8.200 ;
        RECT 10.640 6.970 10.960 7.010 ;
        RECT 10.640 6.850 10.970 6.970 ;
        RECT 10.640 6.750 11.080 6.850 ;
        RECT 10.740 6.680 11.080 6.750 ;
        RECT 12.360 6.580 12.560 6.930 ;
        RECT 10.640 6.420 10.960 6.460 ;
        RECT 10.640 6.230 10.970 6.420 ;
        RECT 10.640 6.200 11.080 6.230 ;
        RECT 10.740 6.060 11.080 6.200 ;
        RECT 11.630 5.960 11.830 6.560 ;
        RECT 12.360 6.550 12.570 6.580 ;
        RECT 12.350 5.960 12.570 6.550 ;
        RECT 2.820 4.930 2.990 5.460 ;
        RECT 6.760 4.920 6.930 5.450 ;
        RECT 10.740 4.350 11.080 4.490 ;
        RECT 10.640 4.320 11.080 4.350 ;
        RECT 2.830 3.220 3.000 4.230 ;
        RECT 10.640 4.130 10.970 4.320 ;
        RECT 10.640 4.090 10.960 4.130 ;
        RECT 6.760 3.080 6.930 4.090 ;
        RECT 11.630 3.990 11.830 4.590 ;
        RECT 12.350 4.000 12.570 4.590 ;
        RECT 12.360 3.970 12.570 4.000 ;
        RECT 10.740 3.800 11.080 3.870 ;
        RECT 8.860 3.570 9.300 3.740 ;
        RECT 10.640 3.700 11.080 3.800 ;
        RECT 10.640 3.610 10.970 3.700 ;
        RECT 10.640 3.510 11.080 3.610 ;
        RECT 10.740 3.440 11.080 3.510 ;
        RECT 12.360 3.340 12.560 3.970 ;
        RECT 10.640 3.180 10.960 3.220 ;
        RECT 10.640 2.990 10.970 3.180 ;
        RECT 10.640 2.960 11.080 2.990 ;
        RECT 10.740 2.820 11.080 2.960 ;
        RECT 11.630 2.720 11.830 3.320 ;
        RECT 12.360 3.310 12.570 3.340 ;
        RECT 12.350 2.720 12.570 3.310 ;
        RECT 10.740 1.120 11.080 1.260 ;
        RECT 10.640 1.090 11.080 1.120 ;
        RECT 10.640 0.900 10.970 1.090 ;
        RECT 10.640 0.860 10.960 0.900 ;
        RECT 11.630 0.760 11.830 1.360 ;
        RECT 12.350 0.770 12.570 1.360 ;
        RECT 12.360 0.740 12.570 0.770 ;
        RECT 10.740 0.570 11.080 0.640 ;
        RECT 10.640 0.470 11.080 0.570 ;
        RECT 10.640 0.350 10.970 0.470 ;
        RECT 12.360 0.390 12.560 0.740 ;
        RECT 10.640 0.310 10.960 0.350 ;
      LAYER mcon ;
        RECT 14.900 7.920 15.170 8.190 ;
        RECT 18.930 7.850 19.200 8.120 ;
        RECT 10.700 6.790 10.870 6.960 ;
        RECT 10.700 6.240 10.870 6.410 ;
        RECT 11.640 6.350 11.810 6.520 ;
        RECT 12.370 6.380 12.540 6.550 ;
        RECT 2.820 5.290 2.990 5.460 ;
        RECT 6.760 5.280 6.930 5.450 ;
        RECT 10.700 4.140 10.870 4.310 ;
        RECT 2.830 3.830 3.000 4.000 ;
        RECT 2.830 3.470 3.000 3.640 ;
        RECT 11.640 4.030 11.810 4.200 ;
        RECT 12.370 4.000 12.540 4.170 ;
        RECT 6.760 3.690 6.930 3.860 ;
        RECT 9.120 3.570 9.300 3.740 ;
        RECT 10.700 3.550 10.870 3.760 ;
        RECT 6.760 3.330 6.930 3.500 ;
        RECT 10.700 3.000 10.870 3.170 ;
        RECT 11.640 3.110 11.810 3.280 ;
        RECT 12.370 3.140 12.540 3.310 ;
        RECT 10.700 0.910 10.870 1.080 ;
        RECT 11.640 0.800 11.810 0.970 ;
        RECT 12.370 0.770 12.540 0.940 ;
        RECT 10.700 0.360 10.870 0.530 ;
      LAYER met1 ;
        RECT 10.630 6.720 10.950 7.040 ;
        RECT 11.630 6.580 11.790 7.310 ;
        RECT 11.630 6.560 11.830 6.580 ;
        RECT 10.630 6.170 10.950 6.490 ;
        RECT 11.610 6.320 11.840 6.560 ;
        RECT 11.630 6.270 11.840 6.320 ;
        RECT 12.000 6.270 12.190 7.260 ;
        RECT 12.440 6.610 12.600 7.310 ;
        RECT 11.630 5.410 11.790 6.270 ;
        RECT 12.020 6.150 12.190 6.270 ;
        RECT 12.030 5.410 12.190 6.150 ;
        RECT 12.330 6.060 12.600 6.610 ;
        RECT 12.330 6.010 12.610 6.060 ;
        RECT 12.440 5.920 12.610 6.010 ;
        RECT 12.440 5.410 12.600 5.920 ;
        RECT 10.630 4.060 10.950 4.380 ;
        RECT 11.630 4.280 11.790 5.140 ;
        RECT 12.030 4.400 12.190 5.140 ;
        RECT 12.440 4.630 12.600 5.140 ;
        RECT 12.440 4.540 12.610 4.630 ;
        RECT 12.020 4.280 12.190 4.400 ;
        RECT 11.630 4.230 11.840 4.280 ;
        RECT 11.610 3.990 11.840 4.230 ;
        RECT 11.630 3.970 11.830 3.990 ;
        RECT 9.170 3.770 9.300 3.790 ;
        RECT 9.090 3.750 9.330 3.770 ;
        RECT 8.890 3.560 9.330 3.750 ;
        RECT 9.090 3.540 9.330 3.560 ;
        RECT 9.190 3.500 9.300 3.540 ;
        RECT 10.630 3.480 10.950 3.830 ;
        RECT 11.630 3.340 11.790 3.970 ;
        RECT 11.630 3.320 11.830 3.340 ;
        RECT 10.630 2.930 10.950 3.250 ;
        RECT 11.610 3.080 11.840 3.320 ;
        RECT 11.630 3.030 11.840 3.080 ;
        RECT 12.000 3.030 12.190 4.280 ;
        RECT 12.330 4.490 12.610 4.540 ;
        RECT 12.330 3.940 12.600 4.490 ;
        RECT 13.970 4.360 14.350 10.860 ;
        RECT 14.840 7.380 15.230 9.240 ;
        RECT 18.870 7.310 19.260 9.170 ;
        RECT 12.440 3.370 12.600 3.940 ;
        RECT 11.630 2.170 11.790 3.030 ;
        RECT 12.020 2.910 12.190 3.030 ;
        RECT 12.030 2.170 12.190 2.910 ;
        RECT 12.330 2.820 12.600 3.370 ;
        RECT 12.330 2.770 12.610 2.820 ;
        RECT 12.440 2.680 12.610 2.770 ;
        RECT 12.440 2.170 12.600 2.680 ;
        RECT 10.630 0.830 10.950 1.150 ;
        RECT 11.630 1.050 11.790 1.910 ;
        RECT 12.030 1.170 12.190 1.910 ;
        RECT 12.440 1.400 12.600 1.910 ;
        RECT 12.440 1.310 12.610 1.400 ;
        RECT 12.020 1.050 12.190 1.170 ;
        RECT 11.630 1.000 11.840 1.050 ;
        RECT 11.610 0.760 11.840 1.000 ;
        RECT 11.630 0.740 11.830 0.760 ;
        RECT 10.630 0.280 10.950 0.600 ;
        RECT 11.630 0.010 11.790 0.740 ;
        RECT 12.000 0.060 12.190 1.050 ;
        RECT 12.330 1.260 12.610 1.310 ;
        RECT 12.330 0.710 12.600 1.260 ;
        RECT 12.440 0.010 12.600 0.710 ;
      LAYER via ;
        RECT 10.660 6.750 10.920 7.010 ;
        RECT 10.660 6.200 10.920 6.460 ;
        RECT 10.660 4.090 10.920 4.350 ;
        RECT 10.660 3.510 10.920 3.800 ;
        RECT 10.660 2.960 10.920 3.220 ;
        RECT 10.660 0.860 10.920 1.120 ;
        RECT 10.660 0.310 10.920 0.570 ;
      LAYER met2 ;
        RECT 10.630 6.760 10.940 7.050 ;
        RECT 10.630 6.720 12.960 6.760 ;
        RECT 10.780 6.580 12.960 6.720 ;
        RECT 10.630 6.330 10.940 6.500 ;
        RECT 10.400 6.150 10.490 6.330 ;
        RECT 10.630 6.170 12.960 6.330 ;
        RECT 10.790 6.150 12.960 6.170 ;
        RECT 10.400 4.220 10.490 4.400 ;
        RECT 10.790 4.380 12.960 4.400 ;
        RECT 10.630 4.220 12.960 4.380 ;
        RECT 10.630 4.050 10.940 4.220 ;
        RECT 10.780 3.830 12.960 3.970 ;
        RECT 10.630 3.790 12.960 3.830 ;
        RECT 10.630 3.520 10.940 3.790 ;
        RECT 10.630 3.480 12.960 3.520 ;
        RECT 10.780 3.340 12.960 3.480 ;
        RECT 10.630 3.090 10.940 3.260 ;
        RECT 10.400 2.910 10.490 3.090 ;
        RECT 10.630 2.930 12.960 3.090 ;
        RECT 10.790 2.910 12.960 2.930 ;
        RECT 10.400 0.990 10.490 1.170 ;
        RECT 10.790 1.150 12.960 1.170 ;
        RECT 10.630 0.990 12.960 1.150 ;
        RECT 10.630 0.820 10.940 0.990 ;
        RECT 10.780 0.600 12.960 0.740 ;
        RECT 10.630 0.560 12.960 0.600 ;
        RECT 10.630 0.270 10.940 0.560 ;
  END
END sky130_hilas_cellAttempt01

MACRO sky130_hilas_StepUpDigital
  CLASS CORE ;
  FOREIGN sky130_hilas_StepUpDigital ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.360 BY 2.180 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 0.220 0.000 2.720 1.750 ;
        RECT 3.810 0.580 5.580 2.170 ;
        RECT 6.590 1.680 8.360 1.750 ;
        RECT 6.590 0.000 8.360 0.090 ;
      LAYER li1 ;
        RECT 0.160 1.750 0.330 1.790 ;
        RECT 0.160 1.730 1.310 1.750 ;
        RECT 0.160 1.560 1.350 1.730 ;
        RECT 1.800 1.700 2.260 1.730 ;
        RECT 3.570 1.700 3.920 1.800 ;
        RECT 1.800 1.560 2.910 1.700 ;
        RECT 2.090 1.530 2.910 1.560 ;
        RECT 3.150 1.530 4.320 1.700 ;
        RECT 4.570 1.530 5.330 1.700 ;
        RECT 2.090 1.390 2.350 1.530 ;
        RECT 0.560 1.060 0.890 1.230 ;
        RECT 1.170 1.220 2.350 1.390 ;
        RECT 5.100 1.520 5.330 1.530 ;
        RECT 1.170 1.070 1.950 1.220 ;
        RECT 2.090 1.080 2.350 1.220 ;
        RECT 2.650 1.290 2.940 1.320 ;
        RECT 2.650 1.120 2.980 1.290 ;
        RECT 2.650 1.080 2.940 1.120 ;
        RECT 3.560 1.080 3.890 1.340 ;
        RECT 5.100 1.080 5.370 1.520 ;
        RECT 0.000 0.880 0.620 1.050 ;
        RECT 0.630 0.600 0.810 1.060 ;
        RECT 1.170 0.780 1.350 1.070 ;
        RECT 1.590 0.720 1.800 1.050 ;
        RECT 2.090 0.910 2.420 1.080 ;
        RECT 2.660 0.910 4.820 1.080 ;
        RECT 2.090 0.860 2.320 0.910 ;
        RECT 5.070 0.900 5.400 1.080 ;
        RECT 5.750 0.940 5.920 1.000 ;
        RECT 2.150 0.630 2.320 0.860 ;
        RECT 5.730 0.720 5.950 0.940 ;
        RECT 5.750 0.670 5.920 0.720 ;
        RECT 2.150 0.620 2.530 0.630 ;
        RECT 0.630 0.430 1.590 0.600 ;
        RECT 2.060 0.560 2.530 0.620 ;
        RECT 2.060 0.510 2.870 0.560 ;
        RECT 2.060 0.450 2.880 0.510 ;
        RECT 2.140 0.390 2.880 0.450 ;
        RECT 2.140 0.340 2.530 0.390 ;
      LAYER mcon ;
        RECT 3.630 1.570 3.840 1.780 ;
        RECT 1.670 1.140 1.840 1.310 ;
        RECT 2.710 1.100 2.880 1.270 ;
        RECT 5.140 1.200 5.310 1.370 ;
        RECT 0.630 0.800 0.800 0.970 ;
        RECT 0.630 0.440 0.800 0.610 ;
      LAYER met1 ;
        RECT 0.560 0.000 0.850 1.750 ;
        RECT 1.600 1.110 1.920 1.390 ;
        RECT 1.560 1.090 1.920 1.110 ;
        RECT 1.560 0.780 1.840 1.090 ;
        RECT 2.090 0.490 2.400 2.180 ;
        RECT 3.570 1.530 3.920 1.820 ;
        RECT 5.100 1.750 5.340 2.170 ;
        RECT 4.870 1.690 5.340 1.750 ;
        RECT 3.720 1.510 3.920 1.530 ;
        RECT 2.650 1.320 2.960 1.330 ;
        RECT 2.640 1.050 2.960 1.320 ;
        RECT 2.650 1.040 2.940 1.050 ;
        RECT 5.100 0.490 5.340 1.690 ;
        RECT 7.880 1.680 8.120 1.750 ;
        RECT 5.670 0.670 6.080 1.000 ;
      LAYER via ;
        RECT 1.630 1.100 1.890 1.360 ;
        RECT 1.570 0.820 1.830 1.080 ;
        RECT 3.610 1.540 3.870 1.800 ;
        RECT 2.670 1.060 2.930 1.320 ;
        RECT 5.710 0.700 5.970 0.960 ;
      LAYER met2 ;
        RECT 1.600 1.310 1.920 1.360 ;
        RECT 2.630 1.320 2.950 1.330 ;
        RECT 2.630 1.310 2.960 1.320 ;
        RECT 0.290 1.110 2.960 1.310 ;
        RECT 1.600 1.100 1.920 1.110 ;
        RECT 1.530 1.030 1.870 1.090 ;
        RECT 2.630 1.060 2.960 1.110 ;
        RECT 2.630 1.040 2.950 1.060 ;
        RECT 3.610 1.030 3.870 1.830 ;
        RECT 1.530 0.810 3.970 1.030 ;
        RECT 5.680 0.670 6.140 0.990 ;
  END
END sky130_hilas_StepUpDigital

MACRO sky130_hilas_VinjNOR3
  CLASS CORE ;
  FOREIGN sky130_hilas_VinjNOR3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.880 BY 1.640 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 0.010 0.000 3.450 1.640 ;
      LAYER li1 ;
        RECT 0.630 1.210 0.800 1.350 ;
        RECT 1.360 1.230 1.530 1.310 ;
        RECT 2.170 1.230 2.340 1.310 ;
        RECT 3.710 1.270 3.880 1.390 ;
        RECT 0.630 1.040 0.820 1.210 ;
        RECT 0.630 0.940 0.800 1.040 ;
        RECT 1.360 0.660 1.570 1.230 ;
        RECT 2.130 0.980 2.340 1.230 ;
        RECT 2.730 1.050 2.900 1.150 ;
        RECT 3.670 1.100 3.880 1.270 ;
        RECT 5.600 1.200 5.860 1.270 ;
        RECT 6.400 1.200 6.580 1.330 ;
        RECT 3.710 1.060 3.880 1.100 ;
        RECT 2.130 0.660 2.300 0.980 ;
        RECT 2.700 0.880 2.900 1.050 ;
        RECT 2.730 0.780 2.900 0.880 ;
        RECT 4.270 1.020 5.140 1.190 ;
        RECT 5.600 1.020 6.580 1.200 ;
        RECT 0.200 0.560 0.370 0.660 ;
        RECT 0.180 0.390 0.370 0.560 ;
        RECT 0.200 0.330 0.370 0.390 ;
        RECT 0.620 0.600 0.790 0.660 ;
        RECT 0.620 0.330 0.870 0.600 ;
        RECT 1.360 0.410 1.610 0.660 ;
        RECT 0.630 0.310 0.870 0.330 ;
        RECT 1.440 0.320 1.610 0.410 ;
        RECT 2.090 0.410 2.300 0.660 ;
        RECT 4.270 0.580 4.440 1.020 ;
        RECT 5.600 0.580 5.860 1.020 ;
        RECT 6.400 0.910 6.580 1.020 ;
        RECT 2.810 0.410 4.440 0.580 ;
        RECT 4.890 0.410 5.860 0.580 ;
        RECT 6.310 0.410 6.650 0.580 ;
        RECT 2.090 0.330 2.260 0.410 ;
        RECT 3.580 0.370 3.750 0.410 ;
      LAYER mcon ;
        RECT 0.650 1.040 0.820 1.210 ;
        RECT 0.660 0.360 0.830 0.530 ;
        RECT 5.630 0.700 5.810 0.880 ;
      LAYER met1 ;
        RECT 0.620 1.260 0.840 1.600 ;
        RECT 0.620 1.000 0.850 1.260 ;
        RECT 0.090 0.320 0.400 0.670 ;
        RECT 0.620 0.600 0.840 1.000 ;
        RECT 2.640 0.840 2.970 1.100 ;
        RECT 3.610 1.060 4.040 1.350 ;
        RECT 0.620 0.290 0.870 0.600 ;
        RECT 3.480 0.310 3.870 0.580 ;
        RECT 0.620 0.090 0.840 0.290 ;
        RECT 5.590 0.090 5.860 1.610 ;
        RECT 6.410 0.320 6.720 0.640 ;
      LAYER via ;
        RECT 0.120 0.350 0.380 0.610 ;
        RECT 2.680 0.840 2.940 1.100 ;
        RECT 3.670 1.090 3.930 1.350 ;
        RECT 3.540 0.310 3.800 0.570 ;
        RECT 6.440 0.350 6.700 0.610 ;
      LAYER met2 ;
        RECT 0.000 1.290 4.040 1.450 ;
        RECT 2.640 1.020 2.970 1.100 ;
        RECT 3.620 1.060 4.040 1.290 ;
        RECT 2.370 1.000 2.970 1.020 ;
        RECT 0.010 0.840 2.970 1.000 ;
        RECT 0.090 0.510 0.410 0.610 ;
        RECT 0.010 0.350 0.410 0.510 ;
        RECT 3.500 0.490 3.870 0.570 ;
        RECT 3.500 0.480 4.530 0.490 ;
        RECT 6.410 0.480 6.720 0.640 ;
        RECT 3.500 0.310 6.880 0.480 ;
  END
END sky130_hilas_VinjNOR3

MACRO sky130_hilas_VinjDiodeProtect01
  CLASS CORE ;
  FOREIGN sky130_hilas_VinjDiodeProtect01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.590 BY 10.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN OUTPUT 
    ANTENNADIFFAREA 58.685200 ;
    PORT
      LAYER met1 ;
        RECT 14.350 10.250 14.700 10.410 ;
        RECT 14.340 9.300 14.710 10.250 ;
        RECT 13.990 8.930 16.460 9.300 ;
        RECT 12.550 7.470 16.460 8.930 ;
        RECT 2.840 7.460 16.460 7.470 ;
        RECT 2.170 6.900 16.460 7.460 ;
        RECT 2.170 2.600 25.520 6.900 ;
        RECT 2.170 2.320 16.460 2.600 ;
        RECT 12.550 0.770 16.460 2.320 ;
        RECT 12.530 0.000 16.480 0.770 ;
    END
  END OUTPUT 
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.000 7.380 28.590 8.780 ;
        RECT 0.470 7.370 1.400 7.380 ;
        RECT 0.720 6.260 0.890 7.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.440 8.130 2.810 8.760 ;
        RECT 23.780 8.280 27.910 8.680 ;
        RECT 23.780 8.190 27.920 8.280 ;
        RECT 0.470 6.170 1.420 8.130 ;
        RECT 2.170 8.110 2.750 8.130 ;
        RECT 27.390 7.290 27.920 8.190 ;
        RECT 0.700 0.500 1.420 6.170 ;
      LAYER via ;
        RECT 0.660 8.280 2.690 8.610 ;
        RECT 24.050 8.280 27.040 8.630 ;
        RECT 0.600 7.420 1.300 8.040 ;
        RECT 27.480 7.480 27.830 8.240 ;
    END
  END VGND
  PIN VINJ
    ANTENNADIFFAREA 9.088799 ;
    PORT
      LAYER nwell ;
        RECT 14.870 1.910 26.920 7.850 ;
      LAYER met2 ;
        RECT 26.340 2.480 26.980 5.490 ;
        RECT 0.000 1.080 28.590 2.480 ;
        RECT 25.440 0.950 28.070 1.080 ;
        RECT 25.440 0.440 27.990 0.950 ;
        RECT 25.440 0.370 26.060 0.440 ;
    END
  END VINJ
  PIN INPUT
    PORT
      LAYER met1 ;
        RECT 7.710 10.280 11.610 10.870 ;
        RECT 7.710 8.930 8.000 10.280 ;
    END
  END INPUT
  OBS
      LAYER li1 ;
        RECT 7.730 8.930 7.980 10.390 ;
        RECT 7.770 8.920 7.940 8.930 ;
        RECT 14.410 8.900 14.660 10.380 ;
        RECT 0.550 8.180 27.930 8.690 ;
        RECT 0.550 6.250 1.350 8.180 ;
        RECT 1.930 7.730 2.100 7.810 ;
        RECT 13.170 7.730 13.400 7.820 ;
        RECT 1.930 7.720 13.400 7.730 ;
        RECT 0.550 1.670 1.060 6.250 ;
        RECT 1.920 2.250 13.400 7.720 ;
        RECT 1.850 2.080 13.400 2.250 ;
        RECT 1.920 2.020 2.110 2.080 ;
        RECT 13.170 1.840 13.400 2.080 ;
        RECT 1.800 1.670 3.600 1.680 ;
        RECT 13.960 1.670 14.470 8.180 ;
        RECT 15.230 7.290 26.480 7.460 ;
        RECT 15.230 2.420 15.400 7.290 ;
        RECT 15.790 6.960 25.900 6.970 ;
        RECT 15.790 2.730 25.920 6.960 ;
        RECT 26.310 5.530 26.480 7.290 ;
        RECT 15.790 2.650 25.900 2.730 ;
        RECT 15.220 2.350 15.400 2.420 ;
        RECT 26.310 2.350 26.920 5.530 ;
        RECT 15.220 2.180 26.920 2.350 ;
        RECT 26.380 2.070 26.920 2.180 ;
        RECT 27.380 1.830 27.930 8.180 ;
        RECT 27.370 1.670 27.930 1.830 ;
        RECT 0.550 1.330 27.930 1.670 ;
        RECT 0.580 1.160 27.930 1.330 ;
        RECT 0.580 1.140 1.270 1.160 ;
        RECT 1.780 1.150 3.580 1.160 ;
      LAYER mcon ;
        RECT 7.770 9.870 7.940 10.040 ;
        RECT 7.770 9.510 7.940 9.680 ;
        RECT 7.770 9.140 7.940 9.310 ;
        RECT 14.450 10.190 14.620 10.360 ;
        RECT 14.450 9.830 14.620 10.000 ;
        RECT 14.450 9.470 14.620 9.640 ;
        RECT 14.450 9.110 14.620 9.280 ;
        RECT 0.630 8.520 2.490 8.530 ;
        RECT 0.630 8.350 2.500 8.520 ;
        RECT 23.990 8.340 27.150 8.520 ;
        RECT 0.670 6.260 0.850 8.160 ;
        RECT 1.070 6.250 1.250 8.160 ;
        RECT 2.260 7.220 13.240 7.390 ;
        RECT 2.260 6.600 13.240 6.770 ;
        RECT 2.270 5.980 13.250 6.150 ;
        RECT 2.290 5.400 13.270 5.570 ;
        RECT 2.300 4.810 13.280 4.980 ;
        RECT 2.300 4.210 13.280 4.380 ;
        RECT 2.250 3.610 13.230 3.780 ;
        RECT 2.260 3.000 13.240 3.170 ;
        RECT 2.250 2.400 13.230 2.570 ;
        RECT 15.990 6.460 25.440 6.630 ;
        RECT 15.980 5.710 25.370 5.880 ;
        RECT 16.010 4.990 25.410 5.160 ;
        RECT 16.020 4.330 25.390 4.500 ;
        RECT 16.010 3.680 25.460 3.850 ;
        RECT 16.020 3.040 25.410 3.210 ;
        RECT 27.560 7.360 27.760 8.290 ;
        RECT 26.490 2.120 26.840 5.420 ;
      LAYER met1 ;
        RECT 26.290 5.480 26.860 5.490 ;
        RECT 26.290 2.060 26.910 5.480 ;
        RECT 26.290 2.050 26.860 2.060 ;
        RECT 25.460 0.420 26.020 0.920 ;
        RECT 25.470 0.200 26.020 0.420 ;
      LAYER via ;
        RECT 26.450 2.190 26.870 5.360 ;
        RECT 25.480 0.370 26.000 0.890 ;
  END
END sky130_hilas_VinjDiodeProtect01

MACRO sky130_hilas_LevelShift4InputUp
  CLASS CORE ;
  FOREIGN sky130_hilas_LevelShift4InputUp ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.890 BY 7.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 7.850 6.950 8.090 7.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 7.850 0.000 8.090 0.050 ;
    END
  END VPWR
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 0.530 0.000 0.820 0.120 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.220 5.960 2.720 7.440 ;
        RECT 0.190 5.760 2.720 5.960 ;
        RECT 0.220 0.440 2.720 5.760 ;
      LAYER met1 ;
        RECT 0.560 7.000 0.850 7.440 ;
        RECT 0.530 6.910 0.850 7.000 ;
        RECT 0.560 0.440 0.850 6.910 ;
    END
  END VINJ
  PIN OUTPUT1
    PORT
      LAYER met2 ;
        RECT 0.190 6.360 0.350 6.560 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    PORT
      LAYER met2 ;
        RECT 0.190 4.610 0.360 4.810 ;
    END
  END OUTPUT2
  PIN OUTPUT3
    PORT
      LAYER met2 ;
        RECT 0.190 2.860 0.380 3.060 ;
    END
  END OUTPUT3
  PIN OUTPUT4
    PORT
      LAYER met2 ;
        RECT 0.190 1.110 0.350 1.310 ;
    END
  END OUTPUT4
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 4.840 0.000 5.150 0.060 ;
    END
    PORT
      LAYER nwell ;
        RECT 3.810 6.270 5.580 7.860 ;
      LAYER met1 ;
        RECT 5.100 7.440 5.340 7.860 ;
        RECT 4.870 7.380 5.340 7.440 ;
        RECT 5.100 7.000 5.340 7.380 ;
        RECT 4.840 6.940 5.340 7.000 ;
        RECT 5.100 6.180 5.340 6.940 ;
    END
  END VGND
  PIN INPUT1
    PORT
      LAYER met2 ;
        RECT 8.790 5.430 8.890 5.750 ;
    END
  END INPUT1
  PIN INPUT2
    PORT
      LAYER met2 ;
        RECT 8.790 3.680 8.890 4.000 ;
    END
  END INPUT2
  PIN INPUT3
    PORT
      LAYER met2 ;
        RECT 8.790 1.930 8.890 2.250 ;
    END
  END INPUT3
  PIN INPUT4
    PORT
      LAYER met2 ;
        RECT 8.790 0.180 8.890 0.500 ;
    END
  END INPUT4
  OBS
      LAYER nwell ;
        RECT 6.590 7.370 8.360 7.440 ;
        RECT 3.810 4.520 5.580 6.110 ;
        RECT 6.590 5.620 8.360 5.780 ;
        RECT 3.810 2.770 5.580 4.360 ;
        RECT 6.590 3.870 8.360 4.030 ;
        RECT 3.810 1.020 5.580 2.610 ;
        RECT 6.590 2.120 8.360 2.280 ;
        RECT 6.590 0.440 8.360 0.530 ;
      LAYER li1 ;
        RECT 0.160 7.440 0.330 7.480 ;
        RECT 0.160 7.420 1.310 7.440 ;
        RECT 0.160 7.250 1.350 7.420 ;
        RECT 1.800 7.390 2.260 7.420 ;
        RECT 3.570 7.390 3.920 7.490 ;
        RECT 1.800 7.250 2.910 7.390 ;
        RECT 2.090 7.220 2.910 7.250 ;
        RECT 3.150 7.220 4.320 7.390 ;
        RECT 4.570 7.220 5.330 7.390 ;
        RECT 2.090 7.080 2.350 7.220 ;
        RECT 0.560 6.750 0.890 6.920 ;
        RECT 1.170 6.910 2.350 7.080 ;
        RECT 5.100 7.210 5.330 7.220 ;
        RECT 1.170 6.760 1.950 6.910 ;
        RECT 2.090 6.770 2.350 6.910 ;
        RECT 2.650 6.980 2.940 7.010 ;
        RECT 2.650 6.810 2.980 6.980 ;
        RECT 2.650 6.770 2.940 6.810 ;
        RECT 3.560 6.770 3.890 7.030 ;
        RECT 5.100 6.770 5.370 7.210 ;
        RECT 0.000 6.570 0.620 6.740 ;
        RECT 0.630 6.290 0.810 6.750 ;
        RECT 1.170 6.470 1.350 6.760 ;
        RECT 1.590 6.410 1.800 6.740 ;
        RECT 2.090 6.600 2.420 6.770 ;
        RECT 2.660 6.600 4.820 6.770 ;
        RECT 2.090 6.550 2.320 6.600 ;
        RECT 5.070 6.590 5.400 6.770 ;
        RECT 5.750 6.630 5.920 6.690 ;
        RECT 2.150 6.320 2.320 6.550 ;
        RECT 5.730 6.410 5.950 6.630 ;
        RECT 5.750 6.360 5.920 6.410 ;
        RECT 2.150 6.310 2.530 6.320 ;
        RECT 0.630 6.120 1.590 6.290 ;
        RECT 2.060 6.250 2.530 6.310 ;
        RECT 2.060 6.200 2.870 6.250 ;
        RECT 2.060 6.140 2.880 6.200 ;
        RECT 2.140 6.080 2.880 6.140 ;
        RECT 2.140 6.030 2.530 6.080 ;
        RECT 0.160 5.690 0.330 5.730 ;
        RECT 0.160 5.670 1.310 5.690 ;
        RECT 0.160 5.500 1.350 5.670 ;
        RECT 1.800 5.640 2.260 5.670 ;
        RECT 3.570 5.640 3.920 5.740 ;
        RECT 1.800 5.500 2.910 5.640 ;
        RECT 2.090 5.470 2.910 5.500 ;
        RECT 3.150 5.470 4.320 5.640 ;
        RECT 4.570 5.470 5.330 5.640 ;
        RECT 2.090 5.330 2.350 5.470 ;
        RECT 0.560 5.000 0.890 5.170 ;
        RECT 1.170 5.160 2.350 5.330 ;
        RECT 5.100 5.460 5.330 5.470 ;
        RECT 1.170 5.010 1.950 5.160 ;
        RECT 2.090 5.020 2.350 5.160 ;
        RECT 2.650 5.230 2.940 5.260 ;
        RECT 2.650 5.060 2.980 5.230 ;
        RECT 2.650 5.020 2.940 5.060 ;
        RECT 3.560 5.020 3.890 5.280 ;
        RECT 5.100 5.020 5.370 5.460 ;
        RECT 0.000 4.820 0.620 4.990 ;
        RECT 0.630 4.540 0.810 5.000 ;
        RECT 1.170 4.720 1.350 5.010 ;
        RECT 1.590 4.660 1.800 4.990 ;
        RECT 2.090 4.850 2.420 5.020 ;
        RECT 2.660 4.850 4.820 5.020 ;
        RECT 2.090 4.800 2.320 4.850 ;
        RECT 5.070 4.840 5.400 5.020 ;
        RECT 5.750 4.880 5.920 4.940 ;
        RECT 2.150 4.570 2.320 4.800 ;
        RECT 5.730 4.660 5.950 4.880 ;
        RECT 5.750 4.610 5.920 4.660 ;
        RECT 2.150 4.560 2.530 4.570 ;
        RECT 0.630 4.370 1.590 4.540 ;
        RECT 2.060 4.500 2.530 4.560 ;
        RECT 2.060 4.450 2.870 4.500 ;
        RECT 2.060 4.390 2.880 4.450 ;
        RECT 2.140 4.330 2.880 4.390 ;
        RECT 2.140 4.280 2.530 4.330 ;
        RECT 0.160 3.940 0.330 3.980 ;
        RECT 0.160 3.920 1.310 3.940 ;
        RECT 0.160 3.750 1.350 3.920 ;
        RECT 1.800 3.890 2.260 3.920 ;
        RECT 3.570 3.890 3.920 3.990 ;
        RECT 1.800 3.750 2.910 3.890 ;
        RECT 2.090 3.720 2.910 3.750 ;
        RECT 3.150 3.720 4.320 3.890 ;
        RECT 4.570 3.720 5.330 3.890 ;
        RECT 2.090 3.580 2.350 3.720 ;
        RECT 0.560 3.250 0.890 3.420 ;
        RECT 1.170 3.410 2.350 3.580 ;
        RECT 5.100 3.710 5.330 3.720 ;
        RECT 1.170 3.260 1.950 3.410 ;
        RECT 2.090 3.270 2.350 3.410 ;
        RECT 2.650 3.480 2.940 3.510 ;
        RECT 2.650 3.310 2.980 3.480 ;
        RECT 2.650 3.270 2.940 3.310 ;
        RECT 3.560 3.270 3.890 3.530 ;
        RECT 5.100 3.270 5.370 3.710 ;
        RECT 0.000 3.070 0.620 3.240 ;
        RECT 0.630 2.790 0.810 3.250 ;
        RECT 1.170 2.970 1.350 3.260 ;
        RECT 1.590 2.910 1.800 3.240 ;
        RECT 2.090 3.100 2.420 3.270 ;
        RECT 2.660 3.100 4.820 3.270 ;
        RECT 2.090 3.050 2.320 3.100 ;
        RECT 5.070 3.090 5.400 3.270 ;
        RECT 5.750 3.130 5.920 3.190 ;
        RECT 2.150 2.820 2.320 3.050 ;
        RECT 5.730 2.910 5.950 3.130 ;
        RECT 5.750 2.860 5.920 2.910 ;
        RECT 2.150 2.810 2.530 2.820 ;
        RECT 0.630 2.620 1.590 2.790 ;
        RECT 2.060 2.750 2.530 2.810 ;
        RECT 2.060 2.700 2.870 2.750 ;
        RECT 2.060 2.640 2.880 2.700 ;
        RECT 2.140 2.580 2.880 2.640 ;
        RECT 2.140 2.530 2.530 2.580 ;
        RECT 0.160 2.190 0.330 2.230 ;
        RECT 0.160 2.170 1.310 2.190 ;
        RECT 0.160 2.000 1.350 2.170 ;
        RECT 1.800 2.140 2.260 2.170 ;
        RECT 3.570 2.140 3.920 2.240 ;
        RECT 1.800 2.000 2.910 2.140 ;
        RECT 2.090 1.970 2.910 2.000 ;
        RECT 3.150 1.970 4.320 2.140 ;
        RECT 4.570 1.970 5.330 2.140 ;
        RECT 2.090 1.830 2.350 1.970 ;
        RECT 0.560 1.500 0.890 1.670 ;
        RECT 1.170 1.660 2.350 1.830 ;
        RECT 5.100 1.960 5.330 1.970 ;
        RECT 1.170 1.510 1.950 1.660 ;
        RECT 2.090 1.520 2.350 1.660 ;
        RECT 2.650 1.730 2.940 1.760 ;
        RECT 2.650 1.560 2.980 1.730 ;
        RECT 2.650 1.520 2.940 1.560 ;
        RECT 3.560 1.520 3.890 1.780 ;
        RECT 5.100 1.520 5.370 1.960 ;
        RECT 0.000 1.320 0.620 1.490 ;
        RECT 0.630 1.040 0.810 1.500 ;
        RECT 1.170 1.220 1.350 1.510 ;
        RECT 1.590 1.160 1.800 1.490 ;
        RECT 2.090 1.350 2.420 1.520 ;
        RECT 2.660 1.350 4.820 1.520 ;
        RECT 2.090 1.300 2.320 1.350 ;
        RECT 5.070 1.340 5.400 1.520 ;
        RECT 5.750 1.380 5.920 1.440 ;
        RECT 2.150 1.070 2.320 1.300 ;
        RECT 5.730 1.160 5.950 1.380 ;
        RECT 5.750 1.110 5.920 1.160 ;
        RECT 2.150 1.060 2.530 1.070 ;
        RECT 0.630 0.870 1.590 1.040 ;
        RECT 2.060 1.000 2.530 1.060 ;
        RECT 2.060 0.950 2.870 1.000 ;
        RECT 2.060 0.890 2.880 0.950 ;
        RECT 2.140 0.830 2.880 0.890 ;
        RECT 2.140 0.780 2.530 0.830 ;
      LAYER mcon ;
        RECT 3.630 7.260 3.840 7.470 ;
        RECT 1.670 6.830 1.840 7.000 ;
        RECT 2.710 6.790 2.880 6.960 ;
        RECT 5.140 6.890 5.310 7.060 ;
        RECT 0.630 6.490 0.800 6.660 ;
        RECT 0.630 6.130 0.800 6.300 ;
        RECT 3.630 5.510 3.840 5.720 ;
        RECT 1.670 5.080 1.840 5.250 ;
        RECT 2.710 5.040 2.880 5.210 ;
        RECT 5.140 5.140 5.310 5.310 ;
        RECT 0.630 4.740 0.800 4.910 ;
        RECT 0.630 4.380 0.800 4.550 ;
        RECT 3.630 3.760 3.840 3.970 ;
        RECT 1.670 3.330 1.840 3.500 ;
        RECT 2.710 3.290 2.880 3.460 ;
        RECT 5.140 3.390 5.310 3.560 ;
        RECT 0.630 2.990 0.800 3.160 ;
        RECT 0.630 2.630 0.800 2.800 ;
        RECT 3.630 2.010 3.840 2.220 ;
        RECT 1.670 1.580 1.840 1.750 ;
        RECT 2.710 1.540 2.880 1.710 ;
        RECT 5.140 1.640 5.310 1.810 ;
        RECT 0.630 1.240 0.800 1.410 ;
        RECT 0.630 0.880 0.800 1.050 ;
      LAYER met1 ;
        RECT 1.600 6.800 1.920 7.080 ;
        RECT 1.560 6.780 1.920 6.800 ;
        RECT 1.560 6.470 1.840 6.780 ;
        RECT 2.090 6.180 2.400 7.870 ;
        RECT 3.570 7.220 3.920 7.510 ;
        RECT 7.880 7.370 8.120 7.440 ;
        RECT 3.720 7.200 3.920 7.220 ;
        RECT 2.650 7.010 2.960 7.020 ;
        RECT 2.640 6.740 2.960 7.010 ;
        RECT 2.650 6.730 2.940 6.740 ;
        RECT 5.670 6.360 6.080 6.690 ;
        RECT 1.600 5.050 1.920 5.330 ;
        RECT 1.560 5.030 1.920 5.050 ;
        RECT 1.560 4.720 1.840 5.030 ;
        RECT 2.090 4.430 2.400 6.120 ;
        RECT 3.570 5.470 3.920 5.760 ;
        RECT 5.100 5.690 5.340 6.110 ;
        RECT 4.870 5.630 5.340 5.690 ;
        RECT 3.720 5.450 3.920 5.470 ;
        RECT 2.650 5.260 2.960 5.270 ;
        RECT 2.640 4.990 2.960 5.260 ;
        RECT 2.650 4.980 2.940 4.990 ;
        RECT 5.100 4.430 5.340 5.630 ;
        RECT 7.880 5.620 8.120 5.690 ;
        RECT 5.670 4.610 6.080 4.940 ;
        RECT 1.600 3.300 1.920 3.580 ;
        RECT 1.560 3.280 1.920 3.300 ;
        RECT 1.560 2.970 1.840 3.280 ;
        RECT 2.090 2.680 2.400 4.370 ;
        RECT 3.570 3.720 3.920 4.010 ;
        RECT 5.100 3.940 5.340 4.360 ;
        RECT 4.870 3.880 5.340 3.940 ;
        RECT 3.720 3.700 3.920 3.720 ;
        RECT 2.650 3.510 2.960 3.520 ;
        RECT 2.640 3.240 2.960 3.510 ;
        RECT 2.650 3.230 2.940 3.240 ;
        RECT 5.100 2.680 5.340 3.880 ;
        RECT 7.880 3.870 8.120 3.940 ;
        RECT 5.670 2.860 6.080 3.190 ;
        RECT 1.600 1.550 1.920 1.830 ;
        RECT 1.560 1.530 1.920 1.550 ;
        RECT 1.560 1.220 1.840 1.530 ;
        RECT 2.090 0.930 2.400 2.620 ;
        RECT 3.570 1.970 3.920 2.260 ;
        RECT 5.100 2.190 5.340 2.610 ;
        RECT 4.870 2.130 5.340 2.190 ;
        RECT 3.720 1.950 3.920 1.970 ;
        RECT 2.650 1.760 2.960 1.770 ;
        RECT 2.640 1.490 2.960 1.760 ;
        RECT 2.650 1.480 2.940 1.490 ;
        RECT 5.100 0.930 5.340 2.130 ;
        RECT 7.880 2.120 8.120 2.190 ;
        RECT 5.670 1.110 6.080 1.440 ;
      LAYER via ;
        RECT 1.630 6.790 1.890 7.050 ;
        RECT 1.570 6.510 1.830 6.770 ;
        RECT 3.610 7.230 3.870 7.490 ;
        RECT 2.670 6.750 2.930 7.010 ;
        RECT 5.710 6.390 5.970 6.650 ;
        RECT 1.630 5.040 1.890 5.300 ;
        RECT 1.570 4.760 1.830 5.020 ;
        RECT 3.610 5.480 3.870 5.740 ;
        RECT 2.670 5.000 2.930 5.260 ;
        RECT 5.710 4.640 5.970 4.900 ;
        RECT 1.630 3.290 1.890 3.550 ;
        RECT 1.570 3.010 1.830 3.270 ;
        RECT 3.610 3.730 3.870 3.990 ;
        RECT 2.670 3.250 2.930 3.510 ;
        RECT 5.710 2.890 5.970 3.150 ;
        RECT 1.630 1.540 1.890 1.800 ;
        RECT 1.570 1.260 1.830 1.520 ;
        RECT 3.610 1.980 3.870 2.240 ;
        RECT 2.670 1.500 2.930 1.760 ;
        RECT 5.710 1.140 5.970 1.400 ;
      LAYER met2 ;
        RECT 1.600 7.000 1.920 7.050 ;
        RECT 2.630 7.010 2.950 7.020 ;
        RECT 2.630 7.000 2.960 7.010 ;
        RECT 0.290 6.800 2.960 7.000 ;
        RECT 1.600 6.790 1.920 6.800 ;
        RECT 1.530 6.720 1.870 6.780 ;
        RECT 2.630 6.750 2.960 6.800 ;
        RECT 2.630 6.730 2.950 6.750 ;
        RECT 3.610 6.720 3.870 7.520 ;
        RECT 1.530 6.500 3.970 6.720 ;
        RECT 5.680 6.360 6.140 6.680 ;
        RECT 1.600 5.250 1.920 5.300 ;
        RECT 2.630 5.260 2.950 5.270 ;
        RECT 2.630 5.250 2.960 5.260 ;
        RECT 0.290 5.050 2.960 5.250 ;
        RECT 1.600 5.040 1.920 5.050 ;
        RECT 1.530 4.970 1.870 5.030 ;
        RECT 2.630 5.000 2.960 5.050 ;
        RECT 2.630 4.980 2.950 5.000 ;
        RECT 3.610 4.970 3.870 5.770 ;
        RECT 1.530 4.750 3.970 4.970 ;
        RECT 5.680 4.610 6.140 4.930 ;
        RECT 1.600 3.500 1.920 3.550 ;
        RECT 2.630 3.510 2.950 3.520 ;
        RECT 2.630 3.500 2.960 3.510 ;
        RECT 0.290 3.300 2.960 3.500 ;
        RECT 1.600 3.290 1.920 3.300 ;
        RECT 1.530 3.220 1.870 3.280 ;
        RECT 2.630 3.250 2.960 3.300 ;
        RECT 2.630 3.230 2.950 3.250 ;
        RECT 3.610 3.220 3.870 4.020 ;
        RECT 1.530 3.000 3.970 3.220 ;
        RECT 5.680 2.860 6.140 3.180 ;
        RECT 1.600 1.750 1.920 1.800 ;
        RECT 2.630 1.760 2.950 1.770 ;
        RECT 2.630 1.750 2.960 1.760 ;
        RECT 0.290 1.550 2.960 1.750 ;
        RECT 1.600 1.540 1.920 1.550 ;
        RECT 1.530 1.470 1.870 1.530 ;
        RECT 2.630 1.500 2.960 1.550 ;
        RECT 2.630 1.480 2.950 1.500 ;
        RECT 3.610 1.470 3.870 2.270 ;
        RECT 1.530 1.250 3.970 1.470 ;
        RECT 5.680 1.110 6.140 1.430 ;
  END
END sky130_hilas_LevelShift4InputUp

MACRO sky130_hilas_WTA4Stage01
  CLASS CORE ;
  FOREIGN sky130_hilas_WTA4Stage01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.920 BY 14.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 25.990 5.730 26.220 6.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.990 0.140 26.220 0.390 ;
    END
  END VGND
  PIN OUTPUT1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 25.120 4.830 26.380 4.990 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.476800 ;
    ANTENNADIFFAREA 0.725100 ;
    PORT
      LAYER met2 ;
        RECT 24.480 4.810 24.790 5.070 ;
        RECT 24.330 4.650 26.920 4.810 ;
        RECT 24.330 4.480 24.640 4.650 ;
        RECT 24.330 4.220 24.640 4.390 ;
        RECT 24.330 4.060 26.920 4.220 ;
        RECT 24.480 3.800 24.790 4.060 ;
        RECT 25.120 3.900 26.380 4.060 ;
    END
  END OUTPUT2
  PIN OUTPUT3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 25.120 2.060 26.380 2.220 ;
    END
  END OUTPUT3
  PIN OUTPUT4
    USE ANALOG ;
    ANTENNAGATEAREA 0.476800 ;
    ANTENNADIFFAREA 0.725100 ;
    PORT
      LAYER met2 ;
        RECT 24.480 2.040 24.790 2.300 ;
        RECT 24.330 1.880 26.920 2.040 ;
        RECT 24.330 1.730 24.640 1.880 ;
        RECT 25.930 1.730 26.260 1.820 ;
        RECT 19.580 1.560 26.260 1.730 ;
        RECT 24.330 1.450 24.640 1.560 ;
        RECT 25.930 1.530 26.260 1.560 ;
        RECT 24.330 1.290 26.920 1.450 ;
        RECT 24.480 1.030 24.790 1.290 ;
        RECT 25.140 1.130 26.380 1.290 ;
    END
  END OUTPUT4
  PIN INPUT1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 12.300 4.840 12.450 5.260 ;
        RECT 12.300 4.750 15.570 4.840 ;
        RECT 15.640 4.750 15.960 4.950 ;
        RECT 12.300 4.690 15.960 4.750 ;
        RECT 15.430 4.590 15.730 4.690 ;
    END
  END INPUT1
  PIN INPUT2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 12.370 4.360 12.690 4.450 ;
        RECT 12.280 4.190 12.690 4.360 ;
        RECT 12.280 4.090 12.600 4.190 ;
        RECT 15.510 3.610 15.740 3.620 ;
        RECT 15.510 3.580 23.080 3.610 ;
        RECT 12.350 3.310 12.670 3.440 ;
        RECT 15.510 3.410 23.140 3.580 ;
        RECT 15.510 3.310 15.750 3.410 ;
        RECT 12.300 3.130 15.750 3.310 ;
        RECT 22.950 3.210 23.660 3.410 ;
        RECT 12.300 3.110 15.670 3.130 ;
    END
  END INPUT2
  PIN INPUT3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 15.640 2.930 15.960 3.070 ;
        RECT 15.640 2.910 23.100 2.930 ;
        RECT 15.640 2.810 23.660 2.910 ;
        RECT 15.650 2.710 23.660 2.810 ;
        RECT 15.650 2.700 15.970 2.710 ;
        RECT 12.240 1.750 12.440 2.250 ;
        RECT 15.510 1.750 15.830 1.890 ;
        RECT 12.240 1.630 15.830 1.750 ;
        RECT 12.240 1.550 15.790 1.630 ;
    END
  END INPUT3
  PIN INPUT4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 12.350 1.310 12.660 1.490 ;
        RECT 12.230 1.160 12.660 1.310 ;
        RECT 12.230 1.040 12.510 1.160 ;
        RECT 12.240 0.520 12.810 0.700 ;
        RECT 23.100 0.650 23.650 0.660 ;
        RECT 12.400 0.370 12.710 0.520 ;
        RECT 12.280 0.240 12.710 0.370 ;
        RECT 15.520 0.430 23.650 0.650 ;
        RECT 15.520 0.420 23.110 0.430 ;
        RECT 15.520 0.410 16.290 0.420 ;
        RECT 15.520 0.240 15.760 0.410 ;
        RECT 12.280 0.160 15.760 0.240 ;
        RECT 12.390 0.000 15.760 0.160 ;
    END
  END INPUT4
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 12.260 5.720 12.990 5.900 ;
    END
  END DRAIN1
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT 18.100 6.090 18.480 6.190 ;
    END
  END GATE1
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 22.130 5.910 22.530 6.190 ;
    END
  END VTUN
  PIN WTAMIDDLENODE
    PORT
      LAYER met1 ;
        RECT 24.730 0.140 24.960 0.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 24.730 5.730 24.960 6.190 ;
    END
  END WTAMIDDLENODE
  PIN COLSEL1
    ANTENNADIFFAREA 1.047900 ;
    PORT
      LAYER met2 ;
        RECT 13.360 6.070 13.680 6.130 ;
        RECT 17.380 6.070 17.710 6.100 ;
        RECT 13.360 5.900 17.710 6.070 ;
        RECT 13.360 5.850 13.680 5.900 ;
        RECT 15.660 5.880 15.980 5.900 ;
        RECT 17.380 5.880 17.710 5.900 ;
        RECT 15.660 5.740 23.490 5.880 ;
        RECT 15.840 5.690 23.490 5.740 ;
        RECT 15.840 5.680 23.660 5.690 ;
        RECT 12.610 5.670 23.660 5.680 ;
        RECT 12.610 5.510 20.240 5.670 ;
        RECT 23.280 5.480 23.660 5.670 ;
    END
  END COLSEL1
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 13.980 6.120 14.140 6.190 ;
    END
  END VPWR
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 13.170 6.120 13.330 6.190 ;
    END
  END VINJ
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 12.230 3.770 12.810 3.950 ;
    END
  END DRAIN2
  PIN DRAIN3
    PORT
      LAYER met2 ;
        RECT 12.260 2.480 12.810 2.660 ;
    END
  END DRAIN3
  OBS
      LAYER nwell ;
        RECT 4.000 14.810 5.730 14.870 ;
        RECT 0.000 11.240 1.730 13.080 ;
        RECT 4.000 8.370 6.920 14.810 ;
        RECT 7.280 9.370 9.840 11.280 ;
        RECT 4.690 8.320 6.920 8.370 ;
        RECT 7.280 6.130 9.840 9.120 ;
        RECT 14.820 9.080 15.930 9.350 ;
        RECT 19.080 9.140 19.670 9.300 ;
        RECT 12.640 8.160 12.730 8.240 ;
        RECT 11.120 7.660 11.290 7.720 ;
        RECT 10.940 7.650 11.290 7.660 ;
        RECT 10.940 7.550 10.950 7.650 ;
        RECT 11.120 7.550 11.290 7.650 ;
        RECT 12.410 6.180 15.370 6.190 ;
        RECT 12.410 6.030 12.820 6.180 ;
        RECT 18.100 6.090 18.480 6.190 ;
        RECT 12.410 6.020 13.000 6.030 ;
        RECT 7.280 3.960 9.840 5.870 ;
        RECT 12.410 4.260 12.820 6.020 ;
        RECT 14.820 5.880 15.930 6.070 ;
        RECT 22.130 6.050 22.530 6.190 ;
        RECT 19.080 5.900 19.670 6.050 ;
        RECT 12.300 3.840 12.820 4.260 ;
        RECT 12.300 3.640 12.810 3.840 ;
        RECT 12.300 3.110 12.820 3.640 ;
        RECT 12.410 0.150 12.820 3.110 ;
      LAYER li1 ;
        RECT 0.760 11.690 1.310 12.120 ;
        RECT 4.790 11.760 5.340 12.190 ;
        RECT 9.280 10.930 9.600 10.970 ;
        RECT 7.680 10.540 7.880 10.890 ;
        RECT 9.270 10.810 9.600 10.930 ;
        RECT 9.160 10.710 9.600 10.810 ;
        RECT 9.160 10.640 9.500 10.710 ;
        RECT 7.670 10.510 7.880 10.540 ;
        RECT 7.670 9.920 7.890 10.510 ;
        RECT 8.410 9.920 8.610 10.520 ;
        RECT 9.280 10.380 9.600 10.420 ;
        RECT 9.270 10.190 9.600 10.380 ;
        RECT 9.160 10.160 9.600 10.190 ;
        RECT 9.160 10.020 9.500 10.160 ;
        RECT 13.440 8.820 13.610 9.350 ;
        RECT 17.460 8.850 17.630 9.380 ;
        RECT 7.670 7.980 7.890 8.570 ;
        RECT 7.670 7.950 7.880 7.980 ;
        RECT 8.410 7.970 8.610 8.570 ;
        RECT 9.160 8.330 9.500 8.470 ;
        RECT 9.160 8.300 9.600 8.330 ;
        RECT 9.270 8.110 9.600 8.300 ;
        RECT 9.280 8.070 9.600 8.110 ;
        RECT 7.680 7.300 7.880 7.950 ;
        RECT 9.160 7.780 9.500 7.850 ;
        RECT 9.160 7.680 9.600 7.780 ;
        RECT 9.270 7.570 9.600 7.680 ;
        RECT 9.160 7.470 9.600 7.570 ;
        RECT 10.940 7.550 11.380 7.720 ;
        RECT 9.160 7.400 9.500 7.470 ;
        RECT 7.670 7.270 7.880 7.300 ;
        RECT 7.670 6.680 7.890 7.270 ;
        RECT 8.410 6.680 8.610 7.280 ;
        RECT 9.280 7.140 9.600 7.180 ;
        RECT 9.270 6.950 9.600 7.140 ;
        RECT 13.430 6.960 13.600 8.150 ;
        RECT 9.160 6.920 9.600 6.950 ;
        RECT 17.450 6.920 17.620 8.090 ;
        RECT 9.160 6.780 9.500 6.920 ;
        RECT 7.670 4.730 7.890 5.320 ;
        RECT 7.670 4.700 7.880 4.730 ;
        RECT 8.410 4.720 8.610 5.320 ;
        RECT 25.280 5.280 25.490 5.300 ;
        RECT 9.160 5.080 9.500 5.220 ;
        RECT 25.260 5.110 25.930 5.280 ;
        RECT 9.160 5.050 9.600 5.080 ;
        RECT 9.270 4.860 9.600 5.050 ;
        RECT 9.280 4.820 9.600 4.860 ;
        RECT 24.490 4.990 24.810 5.030 ;
        RECT 24.490 4.900 24.820 4.990 ;
        RECT 25.260 4.900 25.510 5.110 ;
        RECT 24.490 4.880 25.990 4.900 ;
        RECT 24.490 4.780 26.070 4.880 ;
        RECT 24.340 4.730 26.070 4.780 ;
        RECT 7.680 4.350 7.880 4.700 ;
        RECT 9.160 4.530 9.500 4.600 ;
        RECT 24.340 4.560 25.010 4.730 ;
        RECT 25.180 4.710 25.510 4.730 ;
        RECT 25.730 4.710 26.070 4.730 ;
        RECT 9.160 4.430 9.600 4.530 ;
        RECT 24.340 4.520 24.660 4.560 ;
        RECT 9.270 4.310 9.600 4.430 ;
        RECT 9.280 4.270 9.600 4.310 ;
        RECT 24.340 4.310 24.660 4.350 ;
        RECT 24.670 4.310 25.010 4.560 ;
        RECT 25.260 4.540 25.430 4.710 ;
        RECT 25.820 4.540 25.990 4.710 ;
        RECT 25.180 4.330 25.510 4.540 ;
        RECT 25.730 4.330 26.070 4.540 ;
        RECT 24.340 4.140 25.010 4.310 ;
        RECT 25.260 4.160 25.430 4.330 ;
        RECT 25.820 4.160 25.990 4.330 ;
        RECT 25.180 4.140 25.510 4.160 ;
        RECT 25.730 4.140 26.070 4.160 ;
        RECT 24.340 4.090 26.070 4.140 ;
        RECT 24.490 3.990 26.070 4.090 ;
        RECT 24.490 3.970 25.990 3.990 ;
        RECT 24.490 3.880 24.820 3.970 ;
        RECT 24.490 3.840 24.810 3.880 ;
        RECT 25.260 3.760 25.510 3.970 ;
        RECT 26.390 3.910 26.900 4.960 ;
        RECT 25.260 3.590 25.930 3.760 ;
        RECT 25.280 3.570 25.490 3.590 ;
        RECT 25.280 2.510 25.490 2.530 ;
        RECT 25.260 2.340 25.930 2.510 ;
        RECT 24.490 2.220 24.810 2.260 ;
        RECT 24.490 2.130 24.820 2.220 ;
        RECT 25.260 2.130 25.510 2.340 ;
        RECT 24.490 2.110 25.990 2.130 ;
        RECT 24.490 2.010 26.070 2.110 ;
        RECT 24.340 1.960 26.070 2.010 ;
        RECT 24.340 1.790 25.010 1.960 ;
        RECT 25.180 1.940 25.510 1.960 ;
        RECT 25.730 1.940 26.070 1.960 ;
        RECT 24.340 1.750 24.660 1.790 ;
        RECT 24.340 1.540 24.660 1.580 ;
        RECT 24.670 1.540 25.010 1.790 ;
        RECT 25.260 1.770 25.430 1.940 ;
        RECT 25.820 1.770 25.990 1.940 ;
        RECT 25.180 1.560 25.510 1.770 ;
        RECT 25.730 1.560 26.070 1.770 ;
        RECT 12.360 1.410 12.680 1.450 ;
        RECT 12.360 1.240 12.690 1.410 ;
        RECT 24.340 1.370 25.010 1.540 ;
        RECT 25.260 1.390 25.430 1.560 ;
        RECT 25.820 1.390 25.990 1.560 ;
        RECT 25.180 1.370 25.510 1.390 ;
        RECT 25.730 1.370 26.070 1.390 ;
        RECT 24.340 1.320 26.070 1.370 ;
        RECT 12.270 1.220 12.690 1.240 ;
        RECT 24.490 1.220 26.070 1.320 ;
        RECT 12.270 1.190 12.680 1.220 ;
        RECT 24.490 1.200 25.990 1.220 ;
        RECT 12.270 0.490 12.450 1.190 ;
        RECT 24.490 1.110 24.820 1.200 ;
        RECT 24.490 1.070 24.810 1.110 ;
        RECT 25.260 0.990 25.510 1.200 ;
        RECT 26.390 1.140 26.900 2.190 ;
        RECT 25.260 0.820 25.930 0.990 ;
        RECT 25.280 0.800 25.490 0.820 ;
        RECT 12.270 0.450 12.730 0.490 ;
        RECT 12.270 0.320 12.740 0.450 ;
        RECT 12.410 0.260 12.740 0.320 ;
        RECT 12.410 0.230 12.730 0.260 ;
      LAYER mcon ;
        RECT 1.040 11.770 1.310 12.040 ;
        RECT 5.070 11.840 5.340 12.110 ;
        RECT 9.370 10.750 9.540 10.920 ;
        RECT 7.700 10.340 7.870 10.510 ;
        RECT 8.430 10.310 8.600 10.480 ;
        RECT 9.370 10.200 9.540 10.370 ;
        RECT 13.440 9.180 13.610 9.350 ;
        RECT 17.460 9.210 17.630 9.380 ;
        RECT 7.700 7.980 7.870 8.150 ;
        RECT 8.430 8.010 8.600 8.180 ;
        RECT 9.370 8.120 9.540 8.290 ;
        RECT 13.430 7.980 13.600 8.150 ;
        RECT 9.370 7.510 9.540 7.740 ;
        RECT 13.430 7.320 13.600 7.490 ;
        RECT 7.700 7.100 7.870 7.270 ;
        RECT 8.430 7.070 8.600 7.240 ;
        RECT 9.370 6.960 9.540 7.130 ;
        RECT 17.450 7.920 17.620 8.090 ;
        RECT 17.450 7.280 17.620 7.450 ;
        RECT 7.700 4.730 7.870 4.900 ;
        RECT 25.300 5.110 25.470 5.280 ;
        RECT 8.430 4.760 8.600 4.930 ;
        RECT 9.370 4.870 9.540 5.040 ;
        RECT 24.550 4.810 24.720 4.980 ;
        RECT 24.400 4.570 24.570 4.740 ;
        RECT 9.370 4.320 9.540 4.490 ;
        RECT 26.560 4.540 26.730 4.710 ;
        RECT 24.400 4.130 24.570 4.300 ;
        RECT 26.560 4.160 26.730 4.330 ;
        RECT 24.550 3.890 24.720 4.060 ;
        RECT 25.300 3.590 25.470 3.760 ;
        RECT 25.300 2.340 25.470 2.510 ;
        RECT 24.550 2.040 24.720 2.210 ;
        RECT 24.400 1.800 24.570 1.970 ;
        RECT 26.560 1.770 26.730 1.940 ;
        RECT 12.420 1.230 12.590 1.400 ;
        RECT 24.400 1.360 24.570 1.530 ;
        RECT 26.560 1.390 26.730 1.560 ;
        RECT 24.550 1.120 24.720 1.290 ;
        RECT 25.300 0.820 25.470 0.990 ;
        RECT 12.470 0.270 12.640 0.440 ;
      LAYER met1 ;
        RECT 0.980 11.230 1.370 13.090 ;
        RECT 5.010 11.300 5.400 13.160 ;
        RECT 5.890 8.320 6.270 14.820 ;
        RECT 7.640 10.570 7.800 11.270 ;
        RECT 7.640 10.020 7.910 10.570 ;
        RECT 7.630 9.970 7.910 10.020 ;
        RECT 8.050 10.230 8.240 11.220 ;
        RECT 8.450 10.540 8.610 11.270 ;
        RECT 9.290 10.680 9.610 11.000 ;
        RECT 8.410 10.520 8.610 10.540 ;
        RECT 10.530 10.530 10.690 10.600 ;
        RECT 10.940 10.530 11.130 10.600 ;
        RECT 11.340 10.530 11.500 10.600 ;
        RECT 8.400 10.280 8.630 10.520 ;
        RECT 8.400 10.230 8.610 10.280 ;
        RECT 8.050 10.110 8.220 10.230 ;
        RECT 7.630 9.880 7.800 9.970 ;
        RECT 7.640 9.370 7.800 9.880 ;
        RECT 8.050 9.370 8.210 10.110 ;
        RECT 8.450 9.370 8.610 10.230 ;
        RECT 9.290 10.130 9.610 10.450 ;
        RECT 7.640 8.610 7.800 9.120 ;
        RECT 7.630 8.520 7.800 8.610 ;
        RECT 7.630 8.470 7.910 8.520 ;
        RECT 7.640 7.920 7.910 8.470 ;
        RECT 8.050 8.380 8.210 9.120 ;
        RECT 8.050 8.260 8.220 8.380 ;
        RECT 8.450 8.260 8.610 9.120 ;
        RECT 7.640 7.330 7.800 7.920 ;
        RECT 7.640 6.780 7.910 7.330 ;
        RECT 7.630 6.730 7.910 6.780 ;
        RECT 8.050 6.990 8.240 8.260 ;
        RECT 8.400 8.210 8.610 8.260 ;
        RECT 8.400 7.970 8.630 8.210 ;
        RECT 9.290 8.040 9.610 8.360 ;
        RECT 8.410 7.950 8.610 7.970 ;
        RECT 8.450 7.300 8.610 7.950 ;
        RECT 9.290 7.440 9.610 7.810 ;
        RECT 10.910 7.720 11.150 7.750 ;
        RECT 10.910 7.630 11.340 7.720 ;
        RECT 10.530 7.620 10.690 7.630 ;
        RECT 10.910 7.620 11.500 7.630 ;
        RECT 10.910 7.550 11.340 7.620 ;
        RECT 10.910 7.520 11.150 7.550 ;
        RECT 10.940 7.420 11.050 7.520 ;
        RECT 8.410 7.280 8.610 7.300 ;
        RECT 8.400 7.040 8.630 7.280 ;
        RECT 8.400 6.990 8.610 7.040 ;
        RECT 8.050 6.870 8.220 6.990 ;
        RECT 7.630 6.640 7.800 6.730 ;
        RECT 7.640 6.130 7.800 6.640 ;
        RECT 8.050 6.130 8.210 6.870 ;
        RECT 8.450 6.130 8.610 6.990 ;
        RECT 9.290 6.890 9.610 7.210 ;
        RECT 13.400 6.190 13.650 10.870 ;
        RECT 15.460 10.500 15.840 10.870 ;
        RECT 13.400 6.160 13.770 6.190 ;
        RECT 13.380 6.130 13.770 6.160 ;
        RECT 17.410 6.130 17.680 10.870 ;
        RECT 13.370 6.120 13.770 6.130 ;
        RECT 7.640 5.360 7.800 5.870 ;
        RECT 7.630 5.270 7.800 5.360 ;
        RECT 7.630 5.220 7.910 5.270 ;
        RECT 7.640 4.670 7.910 5.220 ;
        RECT 8.050 5.130 8.210 5.870 ;
        RECT 8.050 5.010 8.220 5.130 ;
        RECT 8.450 5.010 8.610 5.870 ;
        RECT 13.370 5.850 13.670 6.120 ;
        RECT 13.380 5.830 13.660 5.850 ;
        RECT 7.640 3.970 7.800 4.670 ;
        RECT 8.050 4.020 8.240 5.010 ;
        RECT 8.400 4.960 8.610 5.010 ;
        RECT 8.400 4.720 8.630 4.960 ;
        RECT 9.290 4.790 9.610 5.110 ;
        RECT 8.410 4.700 8.610 4.720 ;
        RECT 8.450 3.970 8.610 4.700 ;
        RECT 10.530 4.560 10.690 4.630 ;
        RECT 10.940 4.560 11.130 4.630 ;
        RECT 11.340 4.560 11.500 4.630 ;
        RECT 9.290 4.240 9.610 4.560 ;
        RECT 12.400 4.260 12.660 4.480 ;
        RECT 13.400 4.370 13.650 5.830 ;
        RECT 15.690 5.710 15.950 6.030 ;
        RECT 17.390 5.820 17.700 6.130 ;
        RECT 15.600 4.980 15.810 5.610 ;
        RECT 15.600 4.870 15.930 4.980 ;
        RECT 15.670 4.660 15.930 4.870 ;
        RECT 15.460 4.370 15.840 4.650 ;
        RECT 17.410 4.370 17.680 5.820 ;
        RECT 19.490 4.370 19.890 10.870 ;
        RECT 24.480 4.810 24.800 5.060 ;
        RECT 24.330 4.740 24.800 4.810 ;
        RECT 24.330 4.490 24.650 4.740 ;
        RECT 12.300 4.160 12.660 4.260 ;
        RECT 12.300 3.470 12.510 4.160 ;
        RECT 24.330 4.130 24.650 4.380 ;
        RECT 24.330 4.060 24.800 4.130 ;
        RECT 24.480 3.810 24.800 4.060 ;
        RECT 25.270 3.530 25.500 5.340 ;
        RECT 26.530 3.670 26.760 5.200 ;
        RECT 12.300 3.150 12.640 3.470 ;
        RECT 12.300 3.110 12.510 3.150 ;
        RECT 15.670 3.000 15.930 3.100 ;
        RECT 15.580 2.780 15.930 3.000 ;
        RECT 24.190 2.950 24.420 3.150 ;
        RECT 25.450 2.950 25.680 3.160 ;
        RECT 15.580 1.920 15.740 2.780 ;
        RECT 24.480 2.040 24.800 2.290 ;
        RECT 24.330 1.970 24.800 2.040 ;
        RECT 15.540 1.600 15.800 1.920 ;
        RECT 24.330 1.720 24.650 1.970 ;
        RECT 15.580 1.500 15.740 1.600 ;
        RECT 12.350 1.160 12.670 1.480 ;
        RECT 24.330 1.360 24.650 1.610 ;
        RECT 24.330 1.290 24.800 1.360 ;
        RECT 24.480 1.040 24.800 1.290 ;
        RECT 25.270 0.760 25.500 2.570 ;
        RECT 25.990 1.840 26.220 1.890 ;
        RECT 25.950 1.830 26.230 1.840 ;
        RECT 25.950 1.510 26.250 1.830 ;
        RECT 26.530 0.900 26.760 2.430 ;
        RECT 12.400 0.200 12.720 0.520 ;
        RECT 18.100 0.140 18.480 0.240 ;
      LAYER via ;
        RECT 9.320 10.710 9.580 10.970 ;
        RECT 9.320 10.160 9.580 10.420 ;
        RECT 9.320 8.070 9.580 8.330 ;
        RECT 9.320 7.470 9.580 7.780 ;
        RECT 9.320 6.920 9.580 7.180 ;
        RECT 13.390 5.860 13.650 6.120 ;
        RECT 9.320 4.820 9.580 5.080 ;
        RECT 9.320 4.270 9.580 4.530 ;
        RECT 12.400 4.190 12.660 4.450 ;
        RECT 15.690 5.740 15.950 6.000 ;
        RECT 17.410 5.840 17.680 6.100 ;
        RECT 15.670 4.690 15.930 4.950 ;
        RECT 24.510 4.780 24.770 5.030 ;
        RECT 24.360 4.770 24.770 4.780 ;
        RECT 24.360 4.520 24.620 4.770 ;
        RECT 24.360 4.100 24.620 4.350 ;
        RECT 24.360 4.090 24.770 4.100 ;
        RECT 24.510 3.840 24.770 4.090 ;
        RECT 12.380 3.180 12.640 3.440 ;
        RECT 15.670 2.810 15.930 3.070 ;
        RECT 24.510 2.010 24.770 2.260 ;
        RECT 15.540 1.630 15.800 1.890 ;
        RECT 24.360 2.000 24.770 2.010 ;
        RECT 24.360 1.750 24.620 2.000 ;
        RECT 12.380 1.190 12.640 1.450 ;
        RECT 24.360 1.330 24.620 1.580 ;
        RECT 24.360 1.320 24.770 1.330 ;
        RECT 24.510 1.070 24.770 1.320 ;
        RECT 25.960 1.540 26.230 1.810 ;
        RECT 12.430 0.230 12.690 0.490 ;
      LAYER met2 ;
        RECT 9.300 10.720 9.610 11.010 ;
        RECT 7.280 10.680 9.610 10.720 ;
        RECT 7.280 10.540 9.460 10.680 ;
        RECT 9.300 10.290 9.610 10.460 ;
        RECT 7.280 10.130 9.610 10.290 ;
        RECT 7.280 10.110 9.450 10.130 ;
        RECT 9.750 10.110 9.840 10.290 ;
        RECT 10.170 10.130 10.260 10.310 ;
        RECT 10.170 9.700 10.260 9.880 ;
        RECT 12.630 9.690 20.240 9.880 ;
        RECT 10.170 8.610 10.260 8.790 ;
        RECT 12.610 8.610 20.240 8.790 ;
        RECT 7.280 8.360 9.450 8.380 ;
        RECT 7.280 8.200 9.610 8.360 ;
        RECT 9.750 8.200 9.840 8.380 ;
        RECT 9.300 8.030 9.610 8.200 ;
        RECT 10.170 8.180 10.260 8.360 ;
        RECT 12.640 8.170 12.730 8.200 ;
        RECT 12.610 8.060 12.730 8.170 ;
        RECT 7.280 7.810 9.460 7.950 ;
        RECT 7.280 7.770 9.610 7.810 ;
        RECT 9.300 7.480 9.610 7.770 ;
        RECT 7.280 7.440 9.610 7.480 ;
        RECT 7.280 7.300 9.460 7.440 ;
        RECT 9.300 7.050 9.610 7.220 ;
        RECT 7.280 6.890 9.610 7.050 ;
        RECT 7.280 6.870 9.450 6.890 ;
        RECT 9.750 6.870 9.840 7.050 ;
        RECT 10.170 6.890 10.280 7.070 ;
        RECT 12.610 6.910 12.760 7.080 ;
        RECT 10.170 6.460 10.280 6.640 ;
        RECT 12.610 6.470 19.470 6.640 ;
        RECT 19.770 6.500 20.240 6.660 ;
        RECT 19.770 6.490 20.230 6.500 ;
        RECT 10.170 5.360 10.280 5.540 ;
        RECT 22.770 5.470 22.910 5.480 ;
        RECT 22.770 5.140 22.920 5.470 ;
        RECT 7.280 5.110 9.450 5.130 ;
        RECT 7.280 4.950 9.610 5.110 ;
        RECT 9.750 4.950 9.840 5.130 ;
        RECT 9.300 4.780 9.610 4.950 ;
        RECT 10.170 4.930 10.280 5.110 ;
        RECT 22.770 4.940 23.980 5.140 ;
        RECT 24.090 4.710 24.210 4.920 ;
        RECT 7.280 4.560 9.460 4.700 ;
        RECT 7.280 4.520 9.610 4.560 ;
        RECT 9.300 4.230 9.610 4.520 ;
        RECT 22.880 4.280 24.080 4.380 ;
        RECT 22.870 4.200 24.080 4.280 ;
        RECT 23.800 4.080 24.080 4.200 ;
        RECT 23.800 4.060 23.830 4.080 ;
        RECT 24.090 3.950 24.210 4.160 ;
        RECT 22.860 2.090 23.860 2.250 ;
        RECT 24.090 1.940 24.210 2.150 ;
        RECT 22.870 1.110 23.870 1.280 ;
        RECT 24.090 1.180 24.210 1.390 ;
        RECT 22.870 1.100 23.810 1.110 ;
  END
END sky130_hilas_WTA4Stage01

MACRO sky130_hilas_Trans4small
  CLASS CORE ;
  FOREIGN sky130_hilas_Trans4small ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.400 BY 6.460 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN NFET_SOURCE1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 5.710 0.070 5.750 ;
        RECT 0.000 5.480 0.140 5.710 ;
    END
  END NFET_SOURCE1
  PIN NFET_GATE1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 5.070 0.160 5.240 ;
    END
  END NFET_GATE1
  PIN NFET_SOURCE2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 4.560 0.140 4.730 ;
    END
  END NFET_SOURCE2
  PIN NFET_GATE2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 4.150 0.170 4.320 ;
    END
  END NFET_GATE2
  PIN NFET_SOURCE3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 3.780 0.140 3.810 ;
        RECT 0.000 3.640 0.210 3.780 ;
    END
  END NFET_SOURCE3
  PIN NFET_GATE3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 3.230 0.160 3.400 ;
    END
  END NFET_GATE3
  PIN PFET_SOURCE1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 2.620 0.140 2.810 ;
    END
  END PFET_SOURCE1
  PIN PFET_GATE1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 2.200 0.140 2.390 ;
    END
  END PFET_GATE1
  PIN PFET_SOURCE2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 1.830 0.140 1.850 ;
        RECT 0.000 1.660 0.070 1.830 ;
    END
  END PFET_SOURCE2
  PIN PFET_GATE2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 1.410 0.140 1.430 ;
        RECT 0.000 1.240 0.070 1.410 ;
    END
  END PFET_GATE2
  PIN PFET_SOURCE3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 0.840 0.140 0.890 ;
        RECT 0.000 0.700 0.070 0.840 ;
    END
  END PFET_SOURCE3
  PIN PFET_GATE3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 0.450 0.140 0.470 ;
        RECT 0.000 0.280 0.150 0.450 ;
    END
  END PFET_GATE3
  PIN WELL
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 1.280 0.740 3.310 3.710 ;
        RECT 2.100 0.630 2.640 0.740 ;
        RECT 1.920 0.180 2.640 0.630 ;
        RECT 0.070 0.000 2.640 0.180 ;
      LAYER met2 ;
        RECT 1.850 1.790 2.170 1.990 ;
        RECT 1.850 1.710 2.800 1.790 ;
        RECT 1.760 1.590 2.800 1.710 ;
        RECT 1.760 1.380 2.070 1.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.850 1.950 2.170 1.990 ;
        RECT 1.620 1.720 2.170 1.950 ;
        RECT 1.850 1.700 2.170 1.720 ;
        RECT 1.760 1.670 2.170 1.700 ;
        RECT 1.760 1.380 2.080 1.670 ;
        RECT 2.180 1.270 2.400 5.880 ;
        RECT 2.160 1.200 2.400 1.270 ;
        RECT 2.160 1.100 2.500 1.200 ;
        RECT 2.180 0.970 2.500 1.100 ;
        RECT 2.180 0.000 2.400 0.970 ;
      LAYER via ;
        RECT 1.880 1.700 2.140 1.960 ;
        RECT 1.790 1.410 2.050 1.670 ;
    END
  END WELL
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 1.850 5.080 2.160 5.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.850 5.080 2.170 5.400 ;
        RECT 2.580 5.330 2.800 5.880 ;
        RECT 2.580 5.040 2.900 5.330 ;
        RECT 2.580 0.000 2.800 5.040 ;
      LAYER via ;
        RECT 1.880 5.110 2.140 5.370 ;
    END
  END VGND
  PIN PFET_DRAIN3
    USE ANALOG ;
    ANTENNAGATEAREA 0.163800 ;
    PORT
      LAYER met2 ;
        RECT 1.850 0.830 2.170 1.000 ;
        RECT 1.850 0.680 2.800 0.830 ;
        RECT 1.990 0.630 2.800 0.680 ;
    END
  END PFET_DRAIN3
  PIN PFET_DRAIN1
    USE ANALOG ;
    ANTENNAGATEAREA 0.163800 ;
    ANTENNADIFFAREA 0.117600 ;
    PORT
      LAYER met2 ;
        RECT 1.850 2.750 2.170 2.980 ;
        RECT 1.850 2.700 2.800 2.750 ;
        RECT 1.760 2.550 2.800 2.700 ;
        RECT 1.760 2.370 2.070 2.550 ;
    END
  END PFET_DRAIN1
  PIN NFET_DRAIN3
    USE ANALOG ;
    ANTENNAGATEAREA 0.113400 ;
    ANTENNADIFFAREA 0.117600 ;
    PORT
      LAYER met2 ;
        RECT 1.980 3.690 2.800 3.820 ;
        RECT 1.760 3.650 2.800 3.690 ;
        RECT 1.760 3.360 2.070 3.650 ;
    END
  END NFET_DRAIN3
  PIN NFET_DRAIN2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.980 4.570 2.800 4.740 ;
    END
  END NFET_DRAIN2
  PIN NFET_DRAIN1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.980 5.490 2.800 5.660 ;
    END
  END NFET_DRAIN1
  OBS
      LAYER li1 ;
        RECT 1.850 6.320 2.170 6.360 ;
        RECT 2.940 6.330 3.260 6.370 ;
        RECT 1.850 6.250 2.180 6.320 ;
        RECT 1.850 6.100 2.220 6.250 ;
        RECT 2.020 5.920 2.220 6.100 ;
        RECT 2.610 5.920 2.810 6.250 ;
        RECT 2.940 6.140 3.270 6.330 ;
        RECT 2.940 6.110 3.260 6.140 ;
        RECT 1.470 5.610 1.800 5.780 ;
        RECT 0.310 5.410 0.630 5.450 ;
        RECT 0.310 5.220 0.640 5.410 ;
        RECT 1.860 5.330 2.180 5.370 ;
        RECT 2.950 5.340 3.270 5.380 ;
        RECT 1.860 5.260 2.190 5.330 ;
        RECT 2.200 5.260 2.370 5.310 ;
        RECT 2.690 5.260 2.880 5.300 ;
        RECT 1.860 5.230 2.370 5.260 ;
        RECT 2.620 5.230 2.880 5.260 ;
        RECT 0.310 5.190 0.630 5.220 ;
        RECT 0.330 5.120 0.540 5.190 ;
        RECT 1.860 5.110 2.880 5.230 ;
        RECT 2.950 5.150 3.280 5.340 ;
        RECT 2.950 5.120 3.270 5.150 ;
        RECT 2.030 5.070 2.880 5.110 ;
        RECT 2.030 4.980 2.820 5.070 ;
        RECT 2.030 4.930 2.380 4.980 ;
        RECT 2.620 4.930 2.820 4.980 ;
        RECT 2.200 4.920 2.380 4.930 ;
        RECT 1.480 4.620 1.810 4.790 ;
        RECT 0.290 4.490 0.610 4.530 ;
        RECT 0.290 4.300 0.620 4.490 ;
        RECT 1.860 4.340 2.180 4.380 ;
        RECT 2.950 4.350 3.270 4.390 ;
        RECT 0.290 4.270 0.610 4.300 ;
        RECT 1.860 4.270 2.190 4.340 ;
        RECT 1.860 4.120 2.230 4.270 ;
        RECT 2.030 3.940 2.230 4.120 ;
        RECT 2.620 3.940 2.820 4.270 ;
        RECT 2.950 4.160 3.280 4.350 ;
        RECT 2.950 4.130 3.270 4.160 ;
        RECT 1.480 3.650 1.810 3.800 ;
        RECT 1.480 3.630 2.090 3.650 ;
        RECT 1.770 3.610 2.090 3.630 ;
        RECT 0.270 3.500 0.590 3.540 ;
        RECT 0.270 3.310 0.600 3.500 ;
        RECT 1.770 3.440 2.100 3.610 ;
        RECT 3.070 3.510 3.390 3.550 ;
        RECT 1.770 3.390 2.250 3.440 ;
        RECT 0.270 3.280 0.590 3.310 ;
        RECT 1.940 3.260 2.250 3.390 ;
        RECT 1.920 3.240 2.250 3.260 ;
        RECT 2.080 3.110 2.250 3.240 ;
        RECT 2.760 3.110 2.930 3.440 ;
        RECT 3.070 3.320 3.400 3.510 ;
        RECT 3.070 3.290 3.390 3.320 ;
        RECT 1.700 2.910 2.130 2.930 ;
        RECT 1.680 2.740 2.130 2.910 ;
        RECT 1.700 2.720 2.130 2.740 ;
        RECT 1.770 2.620 2.090 2.660 ;
        RECT 1.770 2.450 2.100 2.620 ;
        RECT 3.070 2.520 3.390 2.560 ;
        RECT 1.770 2.400 2.250 2.450 ;
        RECT 1.940 2.270 2.250 2.400 ;
        RECT 1.920 2.250 2.250 2.270 ;
        RECT 2.080 2.120 2.250 2.250 ;
        RECT 2.760 2.120 2.930 2.450 ;
        RECT 3.070 2.330 3.400 2.520 ;
        RECT 3.070 2.300 3.390 2.330 ;
        RECT 1.700 1.920 2.130 1.940 ;
        RECT 1.680 1.750 2.130 1.920 ;
        RECT 1.700 1.730 2.130 1.750 ;
        RECT 1.770 1.630 2.090 1.670 ;
        RECT 1.770 1.460 2.100 1.630 ;
        RECT 3.070 1.530 3.390 1.570 ;
        RECT 1.770 1.410 2.250 1.460 ;
        RECT 1.940 1.280 2.250 1.410 ;
        RECT 1.920 1.270 2.250 1.280 ;
        RECT 1.920 1.260 2.410 1.270 ;
        RECT 2.080 1.180 2.410 1.260 ;
        RECT 2.080 1.100 2.470 1.180 ;
        RECT 2.760 1.130 2.930 1.460 ;
        RECT 3.070 1.340 3.400 1.530 ;
        RECT 3.070 1.310 3.390 1.340 ;
        RECT 2.240 0.990 2.470 1.100 ;
        RECT 1.700 0.930 2.130 0.950 ;
        RECT 1.680 0.760 2.130 0.930 ;
        RECT 1.700 0.740 2.130 0.760 ;
      LAYER mcon ;
        RECT 1.910 6.140 2.080 6.310 ;
        RECT 3.000 6.150 3.170 6.320 ;
        RECT 0.370 5.230 0.540 5.400 ;
        RECT 1.920 5.150 2.090 5.320 ;
        RECT 2.700 5.100 2.870 5.270 ;
        RECT 3.010 5.160 3.180 5.330 ;
        RECT 0.350 4.310 0.520 4.480 ;
        RECT 1.920 4.160 2.090 4.330 ;
        RECT 3.010 4.170 3.180 4.340 ;
        RECT 0.330 3.320 0.500 3.490 ;
        RECT 1.830 3.430 2.000 3.600 ;
        RECT 3.130 3.330 3.300 3.500 ;
        RECT 1.830 2.440 2.000 2.610 ;
        RECT 3.130 2.340 3.300 2.510 ;
        RECT 1.830 1.450 2.000 1.620 ;
        RECT 2.270 1.000 2.440 1.170 ;
        RECT 3.130 1.350 3.300 1.520 ;
      LAYER met1 ;
        RECT 1.840 6.070 2.160 6.390 ;
        RECT 2.930 6.080 3.250 6.400 ;
        RECT 0.300 5.160 0.620 5.480 ;
        RECT 2.940 5.090 3.260 5.410 ;
        RECT 0.280 4.240 0.600 4.560 ;
        RECT 1.850 4.090 2.170 4.410 ;
        RECT 2.940 4.100 3.260 4.420 ;
        RECT 0.260 3.250 0.580 3.570 ;
        RECT 1.760 3.360 2.080 3.680 ;
        RECT 3.060 3.260 3.380 3.580 ;
        RECT 1.850 2.940 2.170 2.980 ;
        RECT 1.620 2.710 2.170 2.940 ;
        RECT 1.850 2.690 2.170 2.710 ;
        RECT 1.760 2.660 2.170 2.690 ;
        RECT 1.760 2.370 2.080 2.660 ;
        RECT 3.060 2.270 3.380 2.590 ;
        RECT 3.060 1.280 3.380 1.600 ;
        RECT 1.850 0.960 2.170 1.000 ;
        RECT 1.620 0.730 2.170 0.960 ;
        RECT 1.850 0.680 2.170 0.730 ;
      LAYER via ;
        RECT 1.870 6.100 2.130 6.360 ;
        RECT 2.960 6.110 3.220 6.370 ;
        RECT 0.330 5.190 0.590 5.450 ;
        RECT 2.970 5.120 3.230 5.380 ;
        RECT 0.310 4.270 0.570 4.530 ;
        RECT 1.880 4.120 2.140 4.380 ;
        RECT 2.970 4.130 3.230 4.390 ;
        RECT 0.290 3.280 0.550 3.540 ;
        RECT 1.790 3.390 2.050 3.650 ;
        RECT 3.090 3.290 3.350 3.550 ;
        RECT 1.880 2.690 2.140 2.950 ;
        RECT 1.790 2.400 2.050 2.660 ;
        RECT 3.090 2.300 3.350 2.560 ;
        RECT 3.090 1.310 3.350 1.570 ;
        RECT 1.880 0.710 2.140 0.970 ;
      LAYER met2 ;
        RECT 1.170 5.990 1.770 6.160 ;
        RECT 1.840 6.070 2.150 6.400 ;
        RECT 2.930 6.170 3.240 6.410 ;
        RECT 2.930 6.080 3.250 6.170 ;
        RECT 3.030 6.000 3.250 6.080 ;
        RECT 0.300 5.160 0.610 5.490 ;
        RECT 2.940 5.180 3.250 5.420 ;
        RECT 1.180 5.000 1.780 5.170 ;
        RECT 2.940 5.090 3.260 5.180 ;
        RECT 3.040 5.010 3.260 5.090 ;
        RECT 0.280 4.240 0.590 4.570 ;
        RECT 1.180 4.010 1.780 4.180 ;
        RECT 1.850 4.090 2.160 4.420 ;
        RECT 2.940 4.190 3.250 4.430 ;
        RECT 2.940 4.100 3.260 4.190 ;
        RECT 3.040 4.020 3.260 4.100 ;
        RECT 0.260 3.250 0.570 3.580 ;
        RECT 1.280 3.240 1.650 3.430 ;
        RECT 3.060 3.260 3.370 3.590 ;
        RECT 1.280 2.820 1.660 3.010 ;
        RECT 1.280 2.250 1.650 2.440 ;
        RECT 3.060 2.270 3.370 2.600 ;
        RECT 1.280 1.830 1.660 2.020 ;
        RECT 1.280 1.260 1.650 1.450 ;
        RECT 3.060 1.280 3.370 1.610 ;
        RECT 1.280 0.840 1.660 1.030 ;
  END
END sky130_hilas_Trans4small

MACRO sky130_hilas_FGBiasWeakGate2x1cell
  CLASS CORE ;
  FOREIGN sky130_hilas_FGBiasWeakGate2x1cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.540 BY 10.520 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DRAIN1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 5.840 9.120 6.020 ;
    END
  END DRAIN1
  PIN VIN11
    PORT
      LAYER met2 ;
        RECT 2.080 5.430 2.390 5.630 ;
        RECT 1.790 5.420 2.390 5.430 ;
        RECT 0.000 5.300 2.390 5.420 ;
        RECT 0.000 5.260 2.250 5.300 ;
        RECT 0.000 5.240 1.940 5.260 ;
    END
  END VIN11
  PIN ROW1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 9.340 5.000 9.650 5.220 ;
        RECT 9.340 4.990 11.530 5.000 ;
        RECT 0.000 4.780 11.530 4.990 ;
        RECT 0.000 4.770 10.220 4.780 ;
    END
  END ROW1
  PIN ROW2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 9.340 2.240 9.650 2.460 ;
        RECT 0.000 2.030 11.530 2.240 ;
        RECT 0.000 2.020 10.220 2.030 ;
    END
  END ROW2
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 11.010 0.470 11.290 6.520 ;
    END
  END VINJ
  PIN COLSEL1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 10.570 6.460 10.760 6.520 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.570 0.470 10.760 0.530 ;
    END
  END COLSEL1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2.830 5.550 3.060 6.520 ;
        RECT 2.830 5.300 3.070 5.550 ;
        RECT 2.830 3.660 3.060 5.300 ;
        RECT 2.830 3.370 3.160 3.660 ;
        RECT 2.830 0.470 3.060 3.370 ;
    END
  END VGND
  PIN GATE1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 4.050 0.470 4.280 6.520 ;
    END
  END GATE1
  PIN VTUN
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 0.350 0.480 0.770 6.520 ;
    END
  END VTUN
  PIN DRAIN2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 9.060 1.140 9.220 1.160 ;
        RECT 0.000 1.090 9.220 1.140 ;
        RECT 0.000 0.990 9.100 1.090 ;
    END
  END DRAIN2
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 1.500 1.950 1.710 ;
    END
  END VIN12
  PIN COMMONSOURCE
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 3.800 10.550 4.020 ;
        RECT 10.230 3.760 10.550 3.800 ;
    END
  END COMMONSOURCE
  OBS
      LAYER nwell ;
        RECT 14.520 10.180 16.250 10.520 ;
        RECT 14.500 8.620 16.250 10.180 ;
        RECT 14.500 6.990 16.230 8.620 ;
        RECT 12.990 6.600 16.290 6.990 ;
        RECT 12.990 6.560 16.530 6.600 ;
        RECT 12.990 4.910 16.540 6.560 ;
        RECT 0.590 1.870 1.150 4.290 ;
        RECT 12.990 3.820 16.290 4.910 ;
        RECT 12.990 1.980 16.290 3.170 ;
        RECT 12.990 0.330 16.540 1.980 ;
        RECT 12.990 0.290 16.530 0.330 ;
        RECT 12.990 0.000 16.290 0.290 ;
      LAYER li1 ;
        RECT 14.920 8.790 15.470 9.220 ;
        RECT 14.920 7.060 15.470 7.490 ;
        RECT 13.880 6.360 14.410 6.530 ;
        RECT 1.870 5.510 6.930 6.340 ;
        RECT 15.690 6.260 15.890 6.610 ;
        RECT 15.690 6.230 15.900 6.260 ;
        RECT 1.940 5.430 2.420 5.510 ;
        RECT 14.120 5.430 14.350 6.120 ;
        RECT 2.090 5.330 2.420 5.430 ;
        RECT 2.270 5.180 2.420 5.330 ;
        RECT 9.350 5.140 9.670 5.180 ;
        RECT 9.350 4.950 9.680 5.140 ;
        RECT 9.350 4.920 9.670 4.950 ;
        RECT 14.130 4.280 14.300 5.430 ;
        RECT 14.960 4.370 15.130 5.980 ;
        RECT 15.680 5.650 15.900 6.230 ;
        RECT 15.690 5.640 15.900 5.650 ;
        RECT 15.330 5.470 15.520 5.480 ;
        RECT 15.330 5.180 15.530 5.470 ;
        RECT 15.320 4.850 15.610 5.180 ;
        RECT 14.960 4.180 15.140 4.370 ;
        RECT 3.040 3.630 3.230 3.950 ;
        RECT 2.950 3.540 3.230 3.630 ;
        RECT 2.950 3.400 6.590 3.540 ;
        RECT 3.040 3.360 6.590 3.400 ;
        RECT 3.040 2.940 3.230 3.360 ;
        RECT 9.350 2.380 9.670 2.420 ;
        RECT 4.070 2.320 4.300 2.360 ;
        RECT 9.350 2.190 9.680 2.380 ;
        RECT 9.350 2.160 9.670 2.190 ;
        RECT 2.060 1.860 2.380 1.900 ;
        RECT 2.060 1.670 2.390 1.860 ;
        RECT 2.060 1.640 2.380 1.670 ;
        RECT 2.240 1.500 2.260 1.640 ;
        RECT 1.910 1.420 2.260 1.500 ;
        RECT 14.130 1.460 14.300 2.710 ;
        RECT 14.960 2.620 15.140 2.810 ;
        RECT 1.910 0.570 6.960 1.420 ;
        RECT 14.120 0.770 14.350 1.460 ;
        RECT 14.960 1.010 15.130 2.620 ;
        RECT 15.320 1.810 15.610 2.140 ;
        RECT 15.330 1.520 15.530 1.810 ;
        RECT 15.330 1.510 15.520 1.520 ;
        RECT 15.690 1.340 15.900 1.350 ;
        RECT 15.680 0.760 15.900 1.340 ;
        RECT 15.690 0.730 15.900 0.760 ;
        RECT 13.880 0.460 14.410 0.630 ;
        RECT 15.690 0.380 15.890 0.730 ;
      LAYER mcon ;
        RECT 14.920 8.870 15.190 9.140 ;
        RECT 14.920 7.140 15.190 7.410 ;
        RECT 2.150 5.370 2.320 5.540 ;
        RECT 14.150 5.910 14.320 6.080 ;
        RECT 15.700 6.060 15.870 6.230 ;
        RECT 14.150 5.460 14.320 5.630 ;
        RECT 9.410 4.960 9.580 5.130 ;
        RECT 15.340 5.220 15.520 5.410 ;
        RECT 2.960 3.430 3.130 3.600 ;
        RECT 9.410 2.200 9.580 2.370 ;
        RECT 2.120 1.680 2.290 1.850 ;
        RECT 14.150 1.260 14.320 1.430 ;
        RECT 15.340 1.580 15.520 1.770 ;
        RECT 14.150 0.810 14.320 0.980 ;
        RECT 15.700 0.760 15.870 0.930 ;
      LAYER met1 ;
        RECT 14.860 6.600 15.250 10.190 ;
        RECT 13.810 6.170 14.120 6.560 ;
        RECT 13.810 6.120 14.360 6.170 ;
        RECT 2.080 5.300 2.400 5.620 ;
        RECT 14.100 5.380 14.360 6.120 ;
        RECT 15.330 5.480 15.520 6.930 ;
        RECT 15.770 6.290 15.930 6.930 ;
        RECT 15.660 5.740 15.930 6.290 ;
        RECT 15.660 5.690 15.940 5.740 ;
        RECT 15.770 5.600 15.940 5.690 ;
        RECT 15.330 5.450 15.550 5.480 ;
        RECT 9.340 4.890 9.660 5.210 ;
        RECT 15.310 5.180 15.560 5.450 ;
        RECT 15.320 5.170 15.560 5.180 ;
        RECT 15.320 4.930 15.550 5.170 ;
        RECT 14.930 4.120 15.170 4.500 ;
        RECT 10.260 3.730 10.520 4.050 ;
        RECT 15.360 3.910 15.520 4.930 ;
        RECT 15.770 3.910 15.930 5.600 ;
        RECT 10.260 3.130 10.520 3.450 ;
        RECT 14.930 2.490 15.170 2.870 ;
        RECT 9.340 2.130 9.660 2.450 ;
        RECT 15.360 2.060 15.520 3.080 ;
        RECT 2.050 1.610 2.370 1.930 ;
        RECT 15.320 1.820 15.550 2.060 ;
        RECT 15.320 1.810 15.560 1.820 ;
        RECT 15.310 1.540 15.560 1.810 ;
        RECT 15.330 1.510 15.550 1.540 ;
        RECT 14.100 0.870 14.360 1.510 ;
        RECT 13.810 0.720 14.360 0.870 ;
        RECT 13.810 0.430 14.120 0.720 ;
        RECT 15.330 0.060 15.520 1.510 ;
        RECT 15.770 1.390 15.930 3.080 ;
        RECT 15.770 1.300 15.940 1.390 ;
        RECT 15.660 1.250 15.940 1.300 ;
        RECT 15.660 0.700 15.930 1.250 ;
        RECT 15.770 0.060 15.930 0.700 ;
      LAYER via ;
        RECT 13.840 6.150 14.100 6.410 ;
        RECT 2.110 5.330 2.370 5.590 ;
        RECT 9.370 4.920 9.630 5.180 ;
        RECT 10.260 3.760 10.520 4.020 ;
        RECT 10.260 3.160 10.520 3.420 ;
        RECT 9.370 2.160 9.630 2.420 ;
        RECT 2.080 1.640 2.340 1.900 ;
        RECT 13.840 0.580 14.100 0.840 ;
      LAYER met2 ;
        RECT 13.810 6.440 14.120 6.450 ;
        RECT 13.810 6.260 16.290 6.440 ;
        RECT 13.810 6.120 14.120 6.260 ;
        RECT 10.180 3.420 10.440 3.660 ;
        RECT 10.180 3.310 10.550 3.420 ;
        RECT 10.230 3.160 10.550 3.310 ;
        RECT 2.050 1.610 2.360 1.940 ;
        RECT 13.810 0.730 14.120 0.870 ;
        RECT 13.810 0.550 16.290 0.730 ;
        RECT 13.810 0.540 14.120 0.550 ;
  END
END sky130_hilas_FGBiasWeakGate2x1cell

MACRO sky130_hilas_swc4x2cell
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x2cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 45.720 BY 14.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 27.250 5.950 27.630 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.250 0.000 27.630 0.150 ;
    END
  END GATE2
  PIN VTUN
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 22.120 0.000 22.520 0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.200 0.000 23.600 0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.200 5.950 23.600 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 22.120 5.920 22.520 6.050 ;
    END
  END VTUN
  PIN GATE1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 18.090 5.950 18.470 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 18.090 0.000 18.470 0.090 ;
    END
  END GATE1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 32.400 0.010 32.560 0.070 ;
    END
  END VINJ
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 13.000 6.000 32.740 6.180 ;
        RECT 13.000 5.860 17.490 6.000 ;
        RECT 13.240 5.830 17.490 5.860 ;
        RECT 13.240 5.780 13.560 5.830 ;
        RECT 17.170 5.760 17.490 5.830 ;
        RECT 28.230 5.870 32.740 6.000 ;
        RECT 28.230 5.830 32.480 5.870 ;
        RECT 28.230 5.760 28.550 5.830 ;
        RECT 32.160 5.780 32.480 5.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.280 9.340 13.520 10.730 ;
        RECT 13.270 8.680 13.540 9.340 ;
        RECT 13.280 6.150 13.520 8.680 ;
        RECT 13.010 6.090 13.520 6.150 ;
        RECT 13.010 6.010 13.530 6.090 ;
        RECT 13.000 5.860 13.530 6.010 ;
        RECT 13.160 5.770 13.530 5.860 ;
        RECT 13.160 5.710 13.520 5.770 ;
        RECT 13.280 4.230 13.520 5.710 ;
      LAYER via ;
        RECT 13.040 6.060 13.300 6.140 ;
        RECT 13.040 5.880 13.530 6.060 ;
        RECT 13.270 5.800 13.530 5.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.160 0.000 13.320 0.060 ;
    END
  END VINJ
  PIN GATESELECT1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 13.570 6.000 13.760 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.570 0.010 13.760 0.070 ;
    END
  END GATESELECT1
  PIN GATESELECT2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 31.960 0.010 32.150 0.070 ;
    END
  END GATESELECT2
  PIN COL1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 13.970 6.000 14.130 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.970 0.010 14.130 0.070 ;
    END
  END COL1
  PIN COL2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 31.590 0.010 31.750 0.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.590 6.000 31.750 6.050 ;
    END
  END COL2
  PIN ROW1
    PORT
      LAYER met2 ;
        RECT 12.620 5.220 20.240 5.400 ;
        RECT 12.800 5.110 12.870 5.220 ;
    END
    PORT
      LAYER met2 ;
        RECT 25.480 5.220 33.100 5.400 ;
        RECT 32.830 5.110 32.920 5.220 ;
    END
  END ROW1
  PIN ROW2
    PORT
      LAYER met2 ;
        RECT 12.800 4.000 12.860 4.180 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.860 4.000 32.920 4.180 ;
    END
  END ROW2
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 12.800 5.540 12.860 5.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.830 5.540 32.920 5.720 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 12.800 3.570 12.930 3.750 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.860 3.570 32.920 3.750 ;
    END
  END DRAIN2
  PIN DRAIN3
    PORT
      LAYER met2 ;
        RECT 12.800 2.300 12.870 2.480 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.830 2.300 32.920 2.480 ;
    END
  END DRAIN3
  PIN ROW3
    PORT
      LAYER met2 ;
        RECT 12.800 1.870 12.870 2.050 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.830 1.870 32.920 2.050 ;
    END
  END ROW3
  PIN ROW4
    PORT
      LAYER met2 ;
        RECT 12.800 0.770 12.870 0.950 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.830 0.770 32.920 0.950 ;
    END
  END ROW4
  PIN DRAIN4
    PORT
      LAYER met2 ;
        RECT 12.800 0.340 12.870 0.520 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.830 0.340 32.920 0.520 ;
    END
  END DRAIN4
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 15.910 5.960 16.150 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.910 0.000 16.150 0.080 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.840 0.000 20.080 0.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.490 6.050 19.890 10.730 ;
        RECT 19.490 5.990 20.080 6.050 ;
        RECT 19.490 4.230 19.890 5.990 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.640 0.000 25.880 0.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.570 0.000 29.810 0.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.830 6.050 26.230 10.730 ;
        RECT 25.640 6.000 26.230 6.050 ;
        RECT 25.830 4.230 26.230 6.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.570 5.980 29.810 6.050 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 4.000 14.670 5.730 14.720 ;
        RECT 39.990 14.670 41.720 14.720 ;
        RECT 0.000 11.140 1.730 12.980 ;
        RECT 4.000 8.230 6.920 14.670 ;
        RECT 7.280 9.230 9.840 11.140 ;
        RECT 20.170 9.390 20.240 9.570 ;
        RECT 25.480 9.390 25.550 9.570 ;
        RECT 35.880 9.230 38.440 11.140 ;
        RECT 14.820 8.980 15.930 9.210 ;
        RECT 19.080 9.040 19.670 9.150 ;
        RECT 26.050 9.040 26.640 9.150 ;
        RECT 29.790 8.980 30.900 9.210 ;
        RECT 4.690 8.180 6.920 8.230 ;
        RECT 7.280 5.990 9.840 8.960 ;
        RECT 10.940 7.550 11.290 7.560 ;
        RECT 10.940 7.390 10.950 7.550 ;
        RECT 11.120 7.390 11.290 7.550 ;
        RECT 34.430 7.550 34.780 7.560 ;
        RECT 34.430 7.390 34.600 7.550 ;
        RECT 34.770 7.390 34.780 7.550 ;
        RECT 14.820 5.740 15.930 6.010 ;
        RECT 19.080 5.760 19.670 5.950 ;
        RECT 26.050 5.760 26.640 5.950 ;
        RECT 29.790 5.740 30.900 6.010 ;
        RECT 32.640 5.870 32.730 6.170 ;
        RECT 35.880 5.990 38.440 8.960 ;
        RECT 38.800 8.230 41.720 14.670 ;
        RECT 43.990 11.140 45.720 12.980 ;
        RECT 38.800 8.180 41.030 8.230 ;
        RECT 7.280 3.820 9.840 5.730 ;
        RECT 35.880 3.820 38.440 5.730 ;
        RECT 12.800 3.690 12.930 3.750 ;
        RECT 12.800 3.570 12.870 3.690 ;
      LAYER li1 ;
        RECT 0.760 11.590 1.310 12.020 ;
        RECT 4.790 11.660 5.340 12.090 ;
        RECT 40.380 11.660 40.930 12.090 ;
        RECT 44.410 11.590 44.960 12.020 ;
        RECT 9.280 10.790 9.600 10.830 ;
        RECT 7.680 10.400 7.880 10.750 ;
        RECT 9.270 10.670 9.600 10.790 ;
        RECT 9.160 10.570 9.600 10.670 ;
        RECT 36.120 10.790 36.440 10.830 ;
        RECT 36.120 10.670 36.450 10.790 ;
        RECT 36.120 10.570 36.560 10.670 ;
        RECT 9.160 10.500 9.500 10.570 ;
        RECT 36.220 10.500 36.560 10.570 ;
        RECT 7.670 10.370 7.880 10.400 ;
        RECT 37.840 10.400 38.040 10.750 ;
        RECT 7.670 9.780 7.890 10.370 ;
        RECT 8.410 9.780 8.610 10.380 ;
        RECT 9.280 10.240 9.600 10.280 ;
        RECT 9.270 10.050 9.600 10.240 ;
        RECT 9.160 10.020 9.600 10.050 ;
        RECT 36.120 10.240 36.440 10.280 ;
        RECT 36.120 10.050 36.450 10.240 ;
        RECT 36.120 10.020 36.560 10.050 ;
        RECT 9.160 9.880 9.500 10.020 ;
        RECT 36.220 9.880 36.560 10.020 ;
        RECT 37.110 9.780 37.310 10.380 ;
        RECT 37.840 10.370 38.050 10.400 ;
        RECT 37.830 9.780 38.050 10.370 ;
        RECT 13.310 8.740 13.480 9.270 ;
        RECT 17.250 8.750 17.420 9.280 ;
        RECT 28.300 8.750 28.470 9.280 ;
        RECT 32.240 8.740 32.410 9.270 ;
        RECT 7.670 7.820 7.890 8.410 ;
        RECT 7.670 7.790 7.880 7.820 ;
        RECT 8.410 7.810 8.610 8.410 ;
        RECT 9.160 8.170 9.500 8.310 ;
        RECT 36.220 8.170 36.560 8.310 ;
        RECT 9.160 8.140 9.600 8.170 ;
        RECT 9.270 7.950 9.600 8.140 ;
        RECT 36.120 8.140 36.560 8.170 ;
        RECT 9.280 7.910 9.600 7.950 ;
        RECT 7.680 7.160 7.880 7.790 ;
        RECT 9.160 7.620 9.500 7.690 ;
        RECT 9.160 7.520 9.600 7.620 ;
        RECT 9.270 7.430 9.600 7.520 ;
        RECT 9.160 7.330 9.600 7.430 ;
        RECT 10.940 7.390 11.380 7.560 ;
        RECT 9.160 7.260 9.500 7.330 ;
        RECT 7.670 7.130 7.880 7.160 ;
        RECT 7.670 6.540 7.890 7.130 ;
        RECT 8.410 6.540 8.610 7.140 ;
        RECT 9.280 7.000 9.600 7.040 ;
        RECT 9.270 6.810 9.600 7.000 ;
        RECT 13.310 6.900 13.480 7.910 ;
        RECT 17.240 7.040 17.410 8.050 ;
        RECT 28.310 7.040 28.480 8.050 ;
        RECT 36.120 7.950 36.450 8.140 ;
        RECT 36.120 7.910 36.440 7.950 ;
        RECT 32.240 6.900 32.410 7.910 ;
        RECT 37.110 7.810 37.310 8.410 ;
        RECT 37.830 7.820 38.050 8.410 ;
        RECT 37.840 7.790 38.050 7.820 ;
        RECT 36.220 7.620 36.560 7.690 ;
        RECT 34.340 7.390 34.780 7.560 ;
        RECT 36.120 7.520 36.560 7.620 ;
        RECT 36.120 7.430 36.450 7.520 ;
        RECT 36.120 7.330 36.560 7.430 ;
        RECT 36.220 7.260 36.560 7.330 ;
        RECT 37.840 7.160 38.040 7.790 ;
        RECT 36.120 7.000 36.440 7.040 ;
        RECT 9.160 6.780 9.600 6.810 ;
        RECT 36.120 6.810 36.450 7.000 ;
        RECT 36.120 6.780 36.560 6.810 ;
        RECT 9.160 6.640 9.500 6.780 ;
        RECT 36.220 6.640 36.560 6.780 ;
        RECT 37.110 6.540 37.310 7.140 ;
        RECT 37.840 7.130 38.050 7.160 ;
        RECT 37.830 6.540 38.050 7.130 ;
        RECT 7.670 4.590 7.890 5.180 ;
        RECT 7.670 4.560 7.880 4.590 ;
        RECT 8.410 4.580 8.610 5.180 ;
        RECT 9.160 4.940 9.500 5.080 ;
        RECT 36.220 4.940 36.560 5.080 ;
        RECT 9.160 4.910 9.600 4.940 ;
        RECT 9.270 4.720 9.600 4.910 ;
        RECT 9.280 4.680 9.600 4.720 ;
        RECT 36.120 4.910 36.560 4.940 ;
        RECT 36.120 4.720 36.450 4.910 ;
        RECT 36.120 4.680 36.440 4.720 ;
        RECT 37.110 4.580 37.310 5.180 ;
        RECT 37.830 4.590 38.050 5.180 ;
        RECT 7.680 4.210 7.880 4.560 ;
        RECT 37.840 4.560 38.050 4.590 ;
        RECT 9.160 4.390 9.500 4.460 ;
        RECT 36.220 4.390 36.560 4.460 ;
        RECT 9.160 4.290 9.600 4.390 ;
        RECT 9.270 4.170 9.600 4.290 ;
        RECT 9.280 4.130 9.600 4.170 ;
        RECT 36.120 4.290 36.560 4.390 ;
        RECT 36.120 4.170 36.450 4.290 ;
        RECT 37.840 4.210 38.040 4.560 ;
        RECT 36.120 4.130 36.440 4.170 ;
      LAYER mcon ;
        RECT 1.040 11.670 1.310 11.940 ;
        RECT 5.070 11.740 5.340 12.010 ;
        RECT 40.380 11.740 40.650 12.010 ;
        RECT 44.410 11.670 44.680 11.940 ;
        RECT 9.370 10.610 9.540 10.780 ;
        RECT 36.180 10.610 36.350 10.780 ;
        RECT 7.700 10.200 7.870 10.370 ;
        RECT 8.430 10.170 8.600 10.340 ;
        RECT 9.370 10.060 9.540 10.230 ;
        RECT 36.180 10.060 36.350 10.230 ;
        RECT 37.120 10.170 37.290 10.340 ;
        RECT 37.850 10.200 38.020 10.370 ;
        RECT 13.310 9.100 13.480 9.270 ;
        RECT 17.250 9.110 17.420 9.280 ;
        RECT 28.300 9.110 28.470 9.280 ;
        RECT 32.240 9.100 32.410 9.270 ;
        RECT 7.700 7.820 7.870 7.990 ;
        RECT 8.430 7.850 8.600 8.020 ;
        RECT 9.370 7.960 9.540 8.130 ;
        RECT 9.370 7.370 9.540 7.580 ;
        RECT 13.310 7.510 13.480 7.680 ;
        RECT 13.310 7.150 13.480 7.320 ;
        RECT 7.700 6.960 7.870 7.130 ;
        RECT 8.430 6.930 8.600 7.100 ;
        RECT 9.370 6.820 9.540 6.990 ;
        RECT 17.240 7.650 17.410 7.820 ;
        RECT 17.240 7.290 17.410 7.460 ;
        RECT 36.180 7.960 36.350 8.130 ;
        RECT 28.310 7.650 28.480 7.820 ;
        RECT 28.310 7.290 28.480 7.460 ;
        RECT 37.120 7.850 37.290 8.020 ;
        RECT 37.850 7.820 38.020 7.990 ;
        RECT 32.240 7.510 32.410 7.680 ;
        RECT 34.600 7.390 34.780 7.560 ;
        RECT 36.180 7.370 36.350 7.580 ;
        RECT 32.240 7.150 32.410 7.320 ;
        RECT 36.180 6.820 36.350 6.990 ;
        RECT 37.120 6.930 37.290 7.100 ;
        RECT 37.850 6.960 38.020 7.130 ;
        RECT 7.700 4.590 7.870 4.760 ;
        RECT 8.430 4.620 8.600 4.790 ;
        RECT 9.370 4.730 9.540 4.900 ;
        RECT 36.180 4.730 36.350 4.900 ;
        RECT 37.120 4.620 37.290 4.790 ;
        RECT 37.850 4.590 38.020 4.760 ;
        RECT 9.370 4.180 9.540 4.350 ;
        RECT 36.180 4.180 36.350 4.350 ;
      LAYER met1 ;
        RECT 0.980 11.130 1.370 12.990 ;
        RECT 5.010 11.200 5.400 13.060 ;
        RECT 5.890 8.180 6.270 14.680 ;
        RECT 7.640 10.430 7.800 11.130 ;
        RECT 7.640 9.880 7.910 10.430 ;
        RECT 7.630 9.830 7.910 9.880 ;
        RECT 8.050 10.090 8.240 11.080 ;
        RECT 8.450 10.400 8.610 11.130 ;
        RECT 9.290 10.540 9.610 10.860 ;
        RECT 10.530 10.450 10.690 10.500 ;
        RECT 10.940 10.450 11.130 10.500 ;
        RECT 11.340 10.460 11.500 10.500 ;
        RECT 15.460 10.400 15.840 10.730 ;
        RECT 8.410 10.380 8.610 10.400 ;
        RECT 8.400 10.140 8.630 10.380 ;
        RECT 8.400 10.090 8.610 10.140 ;
        RECT 8.050 9.970 8.220 10.090 ;
        RECT 7.630 9.740 7.800 9.830 ;
        RECT 7.640 9.230 7.800 9.740 ;
        RECT 8.050 9.230 8.210 9.970 ;
        RECT 8.450 9.230 8.610 10.090 ;
        RECT 9.290 9.990 9.610 10.310 ;
        RECT 17.210 9.320 17.450 10.730 ;
        RECT 28.270 9.320 28.510 10.730 ;
        RECT 29.880 10.400 30.260 10.730 ;
        RECT 32.200 9.340 32.440 10.730 ;
        RECT 36.110 10.540 36.430 10.860 ;
        RECT 34.220 10.460 34.380 10.500 ;
        RECT 34.590 10.450 34.780 10.500 ;
        RECT 35.030 10.450 35.190 10.500 ;
        RECT 37.110 10.400 37.270 11.130 ;
        RECT 37.110 10.380 37.310 10.400 ;
        RECT 36.110 9.990 36.430 10.310 ;
        RECT 37.090 10.140 37.320 10.380 ;
        RECT 37.110 10.090 37.320 10.140 ;
        RECT 37.480 10.090 37.670 11.080 ;
        RECT 37.920 10.430 38.080 11.130 ;
        RECT 7.640 8.450 7.800 8.960 ;
        RECT 7.630 8.360 7.800 8.450 ;
        RECT 7.630 8.310 7.910 8.360 ;
        RECT 7.640 7.760 7.910 8.310 ;
        RECT 8.050 8.220 8.210 8.960 ;
        RECT 8.050 8.100 8.220 8.220 ;
        RECT 8.450 8.100 8.610 8.960 ;
        RECT 17.200 8.660 17.460 9.320 ;
        RECT 28.260 8.660 28.520 9.320 ;
        RECT 32.180 8.680 32.450 9.340 ;
        RECT 37.110 9.230 37.270 10.090 ;
        RECT 37.500 9.970 37.670 10.090 ;
        RECT 37.510 9.230 37.670 9.970 ;
        RECT 37.810 9.880 38.080 10.430 ;
        RECT 37.810 9.830 38.090 9.880 ;
        RECT 37.920 9.740 38.090 9.830 ;
        RECT 37.920 9.230 38.080 9.740 ;
        RECT 7.640 7.190 7.800 7.760 ;
        RECT 7.640 6.640 7.910 7.190 ;
        RECT 7.630 6.590 7.910 6.640 ;
        RECT 8.050 6.850 8.240 8.100 ;
        RECT 8.400 8.050 8.610 8.100 ;
        RECT 8.400 7.810 8.630 8.050 ;
        RECT 9.290 7.880 9.610 8.200 ;
        RECT 8.410 7.790 8.610 7.810 ;
        RECT 8.450 7.160 8.610 7.790 ;
        RECT 9.290 7.300 9.610 7.650 ;
        RECT 10.940 7.590 11.070 7.610 ;
        RECT 10.910 7.570 11.150 7.590 ;
        RECT 10.910 7.380 11.350 7.570 ;
        RECT 10.910 7.360 11.150 7.380 ;
        RECT 10.940 7.320 11.050 7.360 ;
        RECT 8.410 7.140 8.610 7.160 ;
        RECT 8.400 6.900 8.630 7.140 ;
        RECT 8.400 6.850 8.610 6.900 ;
        RECT 8.050 6.730 8.220 6.850 ;
        RECT 7.630 6.500 7.800 6.590 ;
        RECT 7.640 5.990 7.800 6.500 ;
        RECT 8.050 5.990 8.210 6.730 ;
        RECT 8.450 5.990 8.610 6.850 ;
        RECT 9.290 6.750 9.610 7.070 ;
        RECT 17.210 6.050 17.450 8.660 ;
        RECT 28.270 6.050 28.510 8.660 ;
        RECT 32.200 6.160 32.440 8.680 ;
        RECT 36.110 7.880 36.430 8.200 ;
        RECT 37.110 8.100 37.270 8.960 ;
        RECT 37.510 8.220 37.670 8.960 ;
        RECT 37.920 8.450 38.080 8.960 ;
        RECT 37.920 8.360 38.090 8.450 ;
        RECT 37.500 8.100 37.670 8.220 ;
        RECT 37.110 8.050 37.320 8.100 ;
        RECT 37.090 7.810 37.320 8.050 ;
        RECT 37.110 7.790 37.310 7.810 ;
        RECT 34.650 7.590 34.780 7.610 ;
        RECT 34.570 7.570 34.810 7.590 ;
        RECT 34.370 7.380 34.810 7.570 ;
        RECT 34.570 7.360 34.810 7.380 ;
        RECT 34.670 7.320 34.780 7.360 ;
        RECT 36.110 7.300 36.430 7.650 ;
        RECT 37.110 7.160 37.270 7.790 ;
        RECT 37.110 7.140 37.310 7.160 ;
        RECT 36.110 6.750 36.430 7.070 ;
        RECT 37.090 6.900 37.320 7.140 ;
        RECT 37.110 6.850 37.320 6.900 ;
        RECT 37.480 6.850 37.670 8.100 ;
        RECT 37.810 8.310 38.090 8.360 ;
        RECT 37.810 7.760 38.080 8.310 ;
        RECT 39.450 8.180 39.830 14.680 ;
        RECT 40.320 11.200 40.710 13.060 ;
        RECT 44.350 11.130 44.740 12.990 ;
        RECT 37.920 7.190 38.080 7.760 ;
        RECT 32.200 6.090 32.730 6.160 ;
        RECT 17.200 5.730 17.460 6.050 ;
        RECT 7.640 5.220 7.800 5.730 ;
        RECT 7.630 5.130 7.800 5.220 ;
        RECT 7.630 5.080 7.910 5.130 ;
        RECT 7.640 4.530 7.910 5.080 ;
        RECT 8.050 4.990 8.210 5.730 ;
        RECT 8.050 4.870 8.220 4.990 ;
        RECT 8.450 4.870 8.610 5.730 ;
        RECT 7.640 3.830 7.800 4.530 ;
        RECT 8.050 3.880 8.240 4.870 ;
        RECT 8.400 4.820 8.610 4.870 ;
        RECT 8.400 4.580 8.630 4.820 ;
        RECT 9.290 4.650 9.610 4.970 ;
        RECT 8.410 4.560 8.610 4.580 ;
        RECT 8.450 3.830 8.610 4.560 ;
        RECT 9.290 4.100 9.610 4.420 ;
        RECT 15.460 4.230 15.840 4.830 ;
        RECT 17.210 4.230 17.450 5.730 ;
        RECT 22.520 5.690 23.200 5.910 ;
        RECT 28.260 5.730 28.520 6.050 ;
        RECT 31.960 6.000 32.150 6.050 ;
        RECT 32.190 5.880 32.730 6.090 ;
        RECT 37.110 5.990 37.270 6.850 ;
        RECT 37.500 6.730 37.670 6.850 ;
        RECT 37.510 5.990 37.670 6.730 ;
        RECT 37.810 6.640 38.080 7.190 ;
        RECT 37.810 6.590 38.090 6.640 ;
        RECT 37.920 6.500 38.090 6.590 ;
        RECT 37.920 5.990 38.080 6.500 ;
        RECT 32.190 5.770 32.560 5.880 ;
        RECT 28.270 4.230 28.510 5.730 ;
        RECT 32.200 5.710 32.560 5.770 ;
        RECT 29.880 4.230 30.260 4.830 ;
        RECT 32.200 4.230 32.440 5.710 ;
        RECT 36.110 4.650 36.430 4.970 ;
        RECT 37.110 4.870 37.270 5.730 ;
        RECT 37.510 4.990 37.670 5.730 ;
        RECT 37.920 5.220 38.080 5.730 ;
        RECT 37.920 5.130 38.090 5.220 ;
        RECT 37.500 4.870 37.670 4.990 ;
        RECT 37.110 4.820 37.320 4.870 ;
        RECT 37.090 4.580 37.320 4.820 ;
        RECT 37.110 4.560 37.310 4.580 ;
        RECT 36.110 4.100 36.430 4.420 ;
        RECT 37.110 3.830 37.270 4.560 ;
        RECT 37.480 3.880 37.670 4.870 ;
        RECT 37.810 5.080 38.090 5.130 ;
        RECT 37.810 4.530 38.080 5.080 ;
        RECT 37.920 3.830 38.080 4.530 ;
      LAYER via ;
        RECT 9.320 10.570 9.580 10.830 ;
        RECT 9.320 10.020 9.580 10.280 ;
        RECT 36.140 10.570 36.400 10.830 ;
        RECT 36.140 10.020 36.400 10.280 ;
        RECT 9.320 7.910 9.580 8.170 ;
        RECT 9.320 7.330 9.580 7.620 ;
        RECT 9.320 6.780 9.580 7.040 ;
        RECT 36.140 7.910 36.400 8.170 ;
        RECT 36.140 7.330 36.400 7.620 ;
        RECT 36.140 6.780 36.400 7.040 ;
        RECT 32.440 6.060 32.700 6.150 ;
        RECT 17.200 5.760 17.460 6.020 ;
        RECT 9.320 4.680 9.580 4.940 ;
        RECT 9.320 4.130 9.580 4.390 ;
        RECT 28.260 5.760 28.520 6.020 ;
        RECT 32.190 5.890 32.700 6.060 ;
        RECT 32.190 5.800 32.450 5.890 ;
        RECT 36.140 4.680 36.400 4.940 ;
        RECT 36.140 4.130 36.400 4.390 ;
      LAYER met2 ;
        RECT 9.300 10.580 9.610 10.870 ;
        RECT 7.280 10.540 9.610 10.580 ;
        RECT 36.110 10.580 36.420 10.870 ;
        RECT 36.110 10.540 38.440 10.580 ;
        RECT 7.280 10.400 9.460 10.540 ;
        RECT 36.260 10.400 38.440 10.540 ;
        RECT 9.300 10.150 9.610 10.320 ;
        RECT 7.280 9.990 9.610 10.150 ;
        RECT 7.280 9.970 9.450 9.990 ;
        RECT 9.750 9.970 9.840 10.150 ;
        RECT 12.610 9.990 20.240 10.170 ;
        RECT 25.480 9.990 33.110 10.170 ;
        RECT 36.110 10.150 36.420 10.320 ;
        RECT 35.880 9.970 35.970 10.150 ;
        RECT 36.110 9.990 38.440 10.150 ;
        RECT 36.270 9.970 38.440 9.990 ;
        RECT 12.610 9.550 20.240 9.730 ;
        RECT 25.480 9.550 33.110 9.730 ;
        RECT 12.610 8.450 20.240 8.630 ;
        RECT 25.480 8.450 33.110 8.630 ;
        RECT 7.280 8.200 9.450 8.220 ;
        RECT 7.280 8.040 9.610 8.200 ;
        RECT 9.750 8.040 9.840 8.220 ;
        RECT 9.300 7.870 9.610 8.040 ;
        RECT 12.610 8.020 20.240 8.200 ;
        RECT 25.480 8.020 33.110 8.200 ;
        RECT 35.880 8.040 35.970 8.220 ;
        RECT 36.270 8.200 38.440 8.220 ;
        RECT 36.110 8.040 38.440 8.200 ;
        RECT 36.110 7.870 36.420 8.040 ;
        RECT 7.280 7.650 9.460 7.790 ;
        RECT 36.260 7.650 38.440 7.790 ;
        RECT 7.280 7.610 9.610 7.650 ;
        RECT 9.300 7.340 9.610 7.610 ;
        RECT 7.280 7.300 9.610 7.340 ;
        RECT 36.110 7.610 38.440 7.650 ;
        RECT 36.110 7.340 36.420 7.610 ;
        RECT 36.110 7.300 38.440 7.340 ;
        RECT 7.280 7.160 9.460 7.300 ;
        RECT 36.260 7.160 38.440 7.300 ;
        RECT 9.300 6.910 9.610 7.080 ;
        RECT 7.280 6.750 9.610 6.910 ;
        RECT 7.280 6.730 9.450 6.750 ;
        RECT 9.750 6.730 9.840 6.910 ;
        RECT 12.620 6.750 20.240 6.930 ;
        RECT 25.480 6.750 33.100 6.930 ;
        RECT 36.110 6.910 36.420 7.080 ;
        RECT 35.880 6.730 35.970 6.910 ;
        RECT 36.110 6.750 38.440 6.910 ;
        RECT 36.270 6.730 38.440 6.750 ;
        RECT 12.610 6.320 20.240 6.500 ;
        RECT 25.480 6.320 33.110 6.500 ;
        RECT 7.280 4.970 9.450 4.990 ;
        RECT 7.280 4.810 9.610 4.970 ;
        RECT 9.750 4.810 9.840 4.990 ;
        RECT 9.300 4.640 9.610 4.810 ;
        RECT 12.640 4.800 20.240 4.970 ;
        RECT 25.480 4.800 33.080 4.970 ;
        RECT 35.880 4.810 35.970 4.990 ;
        RECT 36.270 4.970 38.440 4.990 ;
        RECT 36.110 4.810 38.440 4.970 ;
        RECT 36.110 4.640 36.420 4.810 ;
        RECT 7.280 4.420 9.460 4.560 ;
        RECT 36.260 4.420 38.440 4.560 ;
        RECT 7.280 4.380 9.610 4.420 ;
        RECT 9.300 4.090 9.610 4.380 ;
        RECT 36.110 4.380 38.440 4.420 ;
        RECT 36.110 4.090 36.420 4.380 ;
        RECT 19.500 1.380 26.260 1.560 ;
  END
END sky130_hilas_swc4x2cell

MACRO sky130_hilas_polyresistorGND
  CLASS CORE ;
  FOREIGN sky130_hilas_polyresistorGND ;
  ORIGIN 0.000 0.000 ;
  SIZE 55.470 BY 10.890 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN INPUT
    PORT
      LAYER met1 ;
        RECT 21.060 10.250 23.470 10.890 ;
        RECT 21.080 8.900 21.490 10.250 ;
    END
  END INPUT
  PIN OUTPUT
    ANTENNADIFFAREA 16.452000 ;
    PORT
      LAYER met2 ;
        RECT 0.000 7.380 55.470 8.770 ;
    END
  END OUTPUT
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 27.810 9.590 28.220 10.360 ;
        RECT 27.540 9.320 28.220 9.590 ;
        RECT 27.540 8.890 29.230 9.320 ;
        RECT 0.330 8.710 24.700 8.730 ;
        RECT 0.270 8.320 24.700 8.710 ;
        RECT 0.270 0.070 0.680 8.320 ;
        RECT 26.870 0.820 29.230 8.890 ;
        RECT 33.500 8.720 54.860 8.730 ;
        RECT 33.440 8.330 54.860 8.720 ;
        RECT 33.440 8.320 54.700 8.330 ;
        RECT 26.750 0.000 29.230 0.820 ;
      LAYER via ;
        RECT 0.820 8.410 24.620 8.670 ;
        RECT 33.500 8.410 54.360 8.670 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 21.140 9.120 21.360 10.240 ;
        RECT 21.090 8.930 21.420 9.120 ;
        RECT 27.880 8.930 28.120 10.280 ;
        RECT 0.380 8.460 55.120 8.730 ;
        RECT 0.380 8.330 24.720 8.460 ;
        RECT 33.410 8.330 55.120 8.460 ;
        RECT 0.380 0.730 0.550 8.330 ;
        RECT 54.950 1.250 55.120 8.330 ;
        RECT 26.820 0.390 29.180 0.560 ;
      LAYER mcon ;
        RECT 21.170 10.040 21.340 10.210 ;
        RECT 21.170 9.680 21.340 9.850 ;
        RECT 21.170 9.320 21.340 9.490 ;
        RECT 21.170 8.960 21.340 9.130 ;
        RECT 27.920 9.870 28.090 10.040 ;
        RECT 27.920 9.510 28.090 9.680 ;
        RECT 27.920 9.150 28.090 9.320 ;
        RECT 0.720 8.350 24.620 8.520 ;
        RECT 33.500 8.350 54.670 8.520 ;
        RECT 27.190 0.390 27.360 0.560 ;
        RECT 27.560 0.390 27.730 0.560 ;
        RECT 27.920 0.390 28.090 0.560 ;
        RECT 28.280 0.390 28.450 0.560 ;
        RECT 28.640 0.390 28.820 0.560 ;
        RECT 29.010 0.390 29.180 0.560 ;
      LAYER met2 ;
        RECT 0.000 1.080 55.470 2.480 ;
  END
END sky130_hilas_polyresistorGND

MACRO sky130_hilas_swc4x2cellOverlap
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x2cellOverlap ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.570 BY 10.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VERT1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 5.970 5.990 6.130 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.970 0.010 6.130 0.080 ;
    END
  END VERT1
  PIN HORIZ1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.800 4.940 4.880 5.120 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.670 4.940 22.780 5.120 ;
    END
  END HORIZ1
  PIN DRAIN1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.800 5.370 4.880 5.550 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.660 5.370 22.770 5.550 ;
    END
  END DRAIN1
  PIN HORIZ2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.800 3.940 4.880 4.120 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.670 3.940 22.780 4.120 ;
    END
  END HORIZ2
  PIN DRAIN2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.800 3.510 4.880 3.690 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.670 3.510 22.780 3.690 ;
    END
  END DRAIN2
  PIN DRAIN3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.800 2.360 4.870 2.540 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.660 2.360 22.770 2.540 ;
    END
  END DRAIN3
  PIN HORIZ3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.800 1.930 4.870 2.110 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.660 1.930 22.770 2.110 ;
    END
  END HORIZ3
  PIN HORIZ4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.800 0.940 4.870 1.120 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.660 0.940 22.770 1.120 ;
    END
  END HORIZ4
  PIN DRAIN4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.800 0.510 4.870 0.690 ;
    END
  END DRAIN4
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 5.160 5.990 5.320 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.160 0.010 5.320 0.080 ;
    END
    PORT
      LAYER met1 ;
        RECT 22.250 0.010 22.410 0.080 ;
    END
    PORT
      LAYER met1 ;
        RECT 22.250 5.980 22.410 6.050 ;
    END
  END VINJ
  PIN GATESELECT1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 5.570 5.990 5.760 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.570 0.010 5.760 0.080 ;
    END
  END GATESELECT1
  PIN VERT2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 21.440 5.980 21.600 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.440 0.010 21.600 0.080 ;
    END
  END VERT2
  PIN GATESELECT2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 21.810 5.980 22.000 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.810 0.010 22.000 0.080 ;
    END
  END GATESELECT2
  PIN DRAIN
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 22.660 0.510 22.770 0.690 ;
    END
  END DRAIN
  PIN GATE2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 18.090 0.000 18.330 6.050 ;
    END
  END GATE2
  PIN GATE1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 9.240 0.000 9.490 6.050 ;
    END
  END GATE1
  PIN VTUN
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 12.850 0.000 13.150 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 14.430 0.000 14.730 6.050 ;
    END
  END VTUN
  OBS
      LAYER nwell ;
        RECT 0.240 10.800 4.240 10.870 ;
        RECT 0.000 8.890 4.240 10.800 ;
        RECT 0.240 8.730 4.240 8.890 ;
        RECT 0.000 5.880 4.240 8.730 ;
        RECT 0.240 5.730 4.240 5.880 ;
        RECT 0.000 4.820 4.240 5.730 ;
        RECT 23.330 10.800 27.330 10.870 ;
        RECT 23.330 8.890 27.570 10.800 ;
        RECT 23.330 8.730 27.330 8.890 ;
        RECT 23.330 5.880 27.570 8.730 ;
        RECT 23.330 5.730 27.330 5.880 ;
        RECT 23.330 4.820 27.570 5.730 ;
        RECT 0.000 3.820 2.560 4.820 ;
        RECT 25.010 3.820 27.570 4.820 ;
      LAYER li1 ;
        RECT 0.580 10.410 3.890 10.540 ;
        RECT 0.400 10.060 3.890 10.410 ;
        RECT 0.390 9.560 3.890 10.060 ;
        RECT 0.390 9.440 0.610 9.560 ;
        RECT 1.130 9.440 1.330 9.560 ;
        RECT 1.880 9.540 2.220 9.560 ;
        RECT 10.390 9.550 10.560 10.440 ;
        RECT 17.010 9.550 17.180 10.440 ;
        RECT 23.680 10.410 26.990 10.540 ;
        RECT 23.680 10.060 27.170 10.410 ;
        RECT 23.680 9.560 27.180 10.060 ;
        RECT 25.350 9.540 25.690 9.560 ;
        RECT 26.240 9.440 26.440 9.560 ;
        RECT 26.960 9.440 27.180 9.560 ;
        RECT 0.580 8.180 3.890 9.070 ;
        RECT 0.390 8.090 3.890 8.180 ;
        RECT 0.390 7.600 0.610 8.090 ;
        RECT 1.130 7.600 1.330 8.090 ;
        RECT 1.880 7.940 2.220 8.080 ;
        RECT 10.390 8.030 10.560 8.920 ;
        RECT 17.010 8.030 17.180 8.920 ;
        RECT 23.680 8.180 26.990 9.070 ;
        RECT 23.680 8.090 27.180 8.180 ;
        RECT 25.350 7.940 25.690 8.080 ;
        RECT 1.880 7.910 2.320 7.940 ;
        RECT 1.990 7.720 2.320 7.910 ;
        RECT 2.000 7.680 2.320 7.720 ;
        RECT 25.250 7.910 25.690 7.940 ;
        RECT 25.250 7.720 25.580 7.910 ;
        RECT 25.250 7.680 25.570 7.720 ;
        RECT 26.240 7.600 26.440 8.090 ;
        RECT 26.960 7.600 27.180 8.090 ;
        RECT 0.390 7.560 3.890 7.600 ;
        RECT 0.400 7.390 3.890 7.560 ;
        RECT 23.680 7.560 27.180 7.600 ;
        RECT 0.400 7.220 4.100 7.390 ;
        RECT 0.400 7.050 3.890 7.220 ;
        RECT 0.390 6.620 3.890 7.050 ;
        RECT 0.390 6.430 0.610 6.620 ;
        RECT 1.130 6.430 1.330 6.620 ;
        RECT 1.880 6.530 2.220 6.620 ;
        RECT 10.390 6.580 10.560 7.470 ;
        RECT 17.010 6.580 17.180 7.470 ;
        RECT 23.680 7.390 27.170 7.560 ;
        RECT 23.470 7.220 27.170 7.390 ;
        RECT 23.680 7.050 27.170 7.220 ;
        RECT 23.680 6.620 27.180 7.050 ;
        RECT 25.350 6.530 25.690 6.620 ;
        RECT 26.240 6.430 26.440 6.620 ;
        RECT 26.960 6.430 27.180 6.620 ;
        RECT 0.580 5.180 3.890 6.130 ;
        RECT 0.390 5.150 3.890 5.180 ;
        RECT 0.390 4.590 0.610 5.150 ;
        RECT 0.390 4.560 0.600 4.590 ;
        RECT 1.130 4.580 1.330 5.150 ;
        RECT 1.880 4.940 2.220 5.080 ;
        RECT 10.390 5.040 10.560 5.930 ;
        RECT 17.010 5.040 17.180 5.930 ;
        RECT 23.680 5.180 26.990 6.130 ;
        RECT 23.680 5.150 27.180 5.180 ;
        RECT 25.350 4.940 25.690 5.080 ;
        RECT 1.880 4.910 2.320 4.940 ;
        RECT 1.990 4.720 2.320 4.910 ;
        RECT 2.000 4.680 2.320 4.720 ;
        RECT 25.250 4.910 25.690 4.940 ;
        RECT 25.250 4.720 25.580 4.910 ;
        RECT 25.250 4.680 25.570 4.720 ;
        RECT 26.240 4.580 26.440 5.150 ;
        RECT 26.960 4.590 27.180 5.150 ;
        RECT 0.400 4.210 0.600 4.560 ;
        RECT 26.970 4.560 27.180 4.590 ;
        RECT 1.880 4.390 2.220 4.460 ;
        RECT 25.350 4.390 25.690 4.460 ;
        RECT 1.880 4.290 2.320 4.390 ;
        RECT 1.990 4.170 2.320 4.290 ;
        RECT 2.000 4.130 2.320 4.170 ;
        RECT 25.250 4.290 25.690 4.390 ;
        RECT 25.250 4.170 25.580 4.290 ;
        RECT 26.970 4.210 27.170 4.560 ;
        RECT 25.250 4.130 25.570 4.170 ;
      LAYER mcon ;
        RECT 2.150 10.440 2.320 10.480 ;
        RECT 2.090 10.310 2.320 10.440 ;
        RECT 2.090 10.270 2.260 10.310 ;
        RECT 0.420 9.860 0.590 10.030 ;
        RECT 1.150 9.830 1.320 10.000 ;
        RECT 2.090 9.790 2.260 9.890 ;
        RECT 2.090 9.720 2.320 9.790 ;
        RECT 2.150 9.620 2.320 9.720 ;
        RECT 10.390 10.240 10.560 10.410 ;
        RECT 17.010 10.240 17.180 10.410 ;
        RECT 25.250 10.440 25.420 10.480 ;
        RECT 25.250 10.310 25.480 10.440 ;
        RECT 25.310 10.270 25.480 10.310 ;
        RECT 25.310 9.790 25.480 9.890 ;
        RECT 26.250 9.830 26.420 10.000 ;
        RECT 26.980 9.860 27.150 10.030 ;
        RECT 25.250 9.720 25.480 9.790 ;
        RECT 25.250 9.620 25.420 9.720 ;
        RECT 2.150 8.840 2.320 9.010 ;
        RECT 2.150 8.150 2.320 8.320 ;
        RECT 10.390 8.720 10.560 8.890 ;
        RECT 0.420 7.590 0.590 7.760 ;
        RECT 17.010 8.720 17.180 8.890 ;
        RECT 25.250 8.840 25.420 9.010 ;
        RECT 25.250 8.150 25.420 8.320 ;
        RECT 1.150 7.620 1.320 7.790 ;
        RECT 2.090 7.730 2.260 7.900 ;
        RECT 25.310 7.730 25.480 7.900 ;
        RECT 26.250 7.620 26.420 7.790 ;
        RECT 2.150 7.430 2.320 7.540 ;
        RECT 2.090 7.370 2.320 7.430 ;
        RECT 26.980 7.590 27.150 7.760 ;
        RECT 2.090 7.180 2.260 7.370 ;
        RECT 3.660 7.220 3.840 7.390 ;
        RECT 10.390 7.270 10.560 7.440 ;
        RECT 0.420 6.850 0.590 7.020 ;
        RECT 1.150 6.820 1.320 6.990 ;
        RECT 2.090 6.850 2.260 6.880 ;
        RECT 2.090 6.710 2.320 6.850 ;
        RECT 2.150 6.680 2.320 6.710 ;
        RECT 17.010 7.270 17.180 7.440 ;
        RECT 25.250 7.430 25.420 7.540 ;
        RECT 23.730 7.220 23.910 7.390 ;
        RECT 25.250 7.370 25.480 7.430 ;
        RECT 25.310 7.180 25.480 7.370 ;
        RECT 25.310 6.850 25.480 6.880 ;
        RECT 25.250 6.710 25.480 6.850 ;
        RECT 26.250 6.820 26.420 6.990 ;
        RECT 26.980 6.850 27.150 7.020 ;
        RECT 25.250 6.680 25.420 6.710 ;
        RECT 2.150 5.900 2.320 6.070 ;
        RECT 2.150 5.210 2.320 5.380 ;
        RECT 10.390 5.730 10.560 5.900 ;
        RECT 0.420 4.590 0.590 4.760 ;
        RECT 17.010 5.730 17.180 5.900 ;
        RECT 25.250 5.900 25.420 6.070 ;
        RECT 25.250 5.210 25.420 5.380 ;
        RECT 1.150 4.620 1.320 4.790 ;
        RECT 2.090 4.730 2.260 4.900 ;
        RECT 25.310 4.730 25.480 4.900 ;
        RECT 26.250 4.620 26.420 4.790 ;
        RECT 26.980 4.590 27.150 4.760 ;
        RECT 2.090 4.180 2.260 4.350 ;
        RECT 25.310 4.180 25.480 4.350 ;
      LAYER met1 ;
        RECT 0.360 10.090 0.520 10.790 ;
        RECT 0.360 9.540 0.630 10.090 ;
        RECT 0.350 9.490 0.630 9.540 ;
        RECT 0.770 9.750 0.960 10.740 ;
        RECT 1.170 10.060 1.330 10.790 ;
        RECT 2.120 10.520 2.360 10.540 ;
        RECT 2.010 10.200 2.360 10.520 ;
        RECT 1.130 10.040 1.330 10.060 ;
        RECT 1.120 9.800 1.350 10.040 ;
        RECT 2.120 9.970 2.360 10.200 ;
        RECT 2.010 9.900 2.360 9.970 ;
        RECT 1.120 9.750 1.330 9.800 ;
        RECT 0.770 9.630 0.940 9.750 ;
        RECT 0.350 9.400 0.520 9.490 ;
        RECT 0.360 8.890 0.520 9.400 ;
        RECT 0.770 8.890 0.930 9.630 ;
        RECT 1.170 8.890 1.330 9.750 ;
        RECT 2.010 9.650 2.350 9.900 ;
        RECT 2.120 9.640 2.350 9.650 ;
        RECT 2.110 9.420 2.350 9.640 ;
        RECT 10.360 9.340 10.590 10.630 ;
        RECT 0.360 8.220 0.520 8.730 ;
        RECT 0.350 8.130 0.520 8.220 ;
        RECT 0.350 8.080 0.630 8.130 ;
        RECT 0.360 7.530 0.630 8.080 ;
        RECT 0.770 7.990 0.930 8.730 ;
        RECT 0.770 7.870 0.940 7.990 ;
        RECT 1.170 7.870 1.330 8.730 ;
        RECT 2.120 8.430 2.360 9.070 ;
        RECT 2.120 8.170 2.350 8.430 ;
        RECT 2.110 7.970 2.350 8.170 ;
        RECT 0.360 7.080 0.520 7.530 ;
        RECT 0.360 6.530 0.630 7.080 ;
        RECT 0.350 6.480 0.630 6.530 ;
        RECT 0.770 6.740 0.960 7.870 ;
        RECT 1.120 7.820 1.330 7.870 ;
        RECT 2.010 7.950 2.350 7.970 ;
        RECT 1.120 7.580 1.350 7.820 ;
        RECT 2.010 7.650 2.330 7.950 ;
        RECT 10.360 7.820 10.590 9.110 ;
        RECT 1.130 7.560 1.330 7.580 ;
        RECT 1.170 7.050 1.330 7.560 ;
        RECT 2.120 7.510 2.360 7.600 ;
        RECT 2.010 7.100 2.360 7.510 ;
        RECT 3.660 7.420 3.790 7.440 ;
        RECT 3.630 7.190 3.870 7.420 ;
        RECT 3.660 7.150 3.770 7.190 ;
        RECT 1.130 7.030 1.330 7.050 ;
        RECT 1.120 6.790 1.350 7.030 ;
        RECT 2.120 6.960 2.360 7.100 ;
        RECT 1.120 6.740 1.330 6.790 ;
        RECT 0.770 6.620 0.940 6.740 ;
        RECT 0.350 6.390 0.520 6.480 ;
        RECT 0.360 5.880 0.520 6.390 ;
        RECT 0.770 5.880 0.930 6.620 ;
        RECT 1.170 5.880 1.330 6.740 ;
        RECT 2.010 6.640 2.350 6.960 ;
        RECT 2.110 6.480 2.350 6.640 ;
        RECT 10.360 6.370 10.590 7.660 ;
        RECT 0.360 5.220 0.520 5.730 ;
        RECT 0.350 5.130 0.520 5.220 ;
        RECT 0.350 5.080 0.630 5.130 ;
        RECT 0.360 4.530 0.630 5.080 ;
        RECT 0.770 4.990 0.930 5.730 ;
        RECT 0.770 4.870 0.940 4.990 ;
        RECT 1.170 4.870 1.330 5.730 ;
        RECT 2.120 5.490 2.360 6.130 ;
        RECT 2.120 5.230 2.350 5.490 ;
        RECT 2.110 5.010 2.350 5.230 ;
        RECT 0.360 3.830 0.520 4.530 ;
        RECT 0.770 3.880 0.960 4.870 ;
        RECT 1.120 4.820 1.330 4.870 ;
        RECT 1.120 4.580 1.350 4.820 ;
        RECT 2.010 4.650 2.330 4.970 ;
        RECT 10.360 4.830 10.590 6.120 ;
        RECT 1.130 4.560 1.330 4.580 ;
        RECT 1.170 3.830 1.330 4.560 ;
        RECT 2.010 4.100 2.330 4.420 ;
        RECT 10.960 4.280 11.230 10.330 ;
        RECT 16.340 4.280 16.610 10.330 ;
        RECT 16.980 9.340 17.210 10.630 ;
        RECT 25.210 10.520 25.450 10.540 ;
        RECT 25.210 10.200 25.560 10.520 ;
        RECT 25.210 9.970 25.450 10.200 ;
        RECT 26.240 10.060 26.400 10.790 ;
        RECT 26.240 10.040 26.440 10.060 ;
        RECT 25.210 9.900 25.560 9.970 ;
        RECT 25.220 9.650 25.560 9.900 ;
        RECT 26.220 9.800 26.450 10.040 ;
        RECT 26.240 9.750 26.450 9.800 ;
        RECT 26.610 9.750 26.800 10.740 ;
        RECT 27.050 10.090 27.210 10.790 ;
        RECT 25.220 9.640 25.450 9.650 ;
        RECT 25.220 9.420 25.460 9.640 ;
        RECT 16.980 7.820 17.210 9.110 ;
        RECT 25.210 8.430 25.450 9.070 ;
        RECT 26.240 8.890 26.400 9.750 ;
        RECT 26.630 9.630 26.800 9.750 ;
        RECT 26.640 8.890 26.800 9.630 ;
        RECT 26.940 9.540 27.210 10.090 ;
        RECT 26.940 9.490 27.220 9.540 ;
        RECT 27.050 9.400 27.220 9.490 ;
        RECT 27.050 8.890 27.210 9.400 ;
        RECT 25.220 8.170 25.450 8.430 ;
        RECT 25.220 7.970 25.460 8.170 ;
        RECT 25.220 7.950 25.560 7.970 ;
        RECT 16.980 6.370 17.210 7.660 ;
        RECT 25.240 7.650 25.560 7.950 ;
        RECT 26.240 7.870 26.400 8.730 ;
        RECT 26.640 7.990 26.800 8.730 ;
        RECT 27.050 8.220 27.210 8.730 ;
        RECT 27.050 8.130 27.220 8.220 ;
        RECT 26.630 7.870 26.800 7.990 ;
        RECT 26.240 7.820 26.450 7.870 ;
        RECT 25.210 7.510 25.450 7.600 ;
        RECT 26.220 7.580 26.450 7.820 ;
        RECT 26.240 7.560 26.440 7.580 ;
        RECT 23.780 7.420 23.910 7.440 ;
        RECT 23.700 7.190 23.940 7.420 ;
        RECT 23.800 7.150 23.910 7.190 ;
        RECT 25.210 7.100 25.560 7.510 ;
        RECT 25.210 6.960 25.450 7.100 ;
        RECT 26.240 7.050 26.400 7.560 ;
        RECT 26.240 7.030 26.440 7.050 ;
        RECT 25.220 6.640 25.560 6.960 ;
        RECT 26.220 6.790 26.450 7.030 ;
        RECT 26.240 6.740 26.450 6.790 ;
        RECT 26.610 6.740 26.800 7.870 ;
        RECT 26.940 8.080 27.220 8.130 ;
        RECT 26.940 7.530 27.210 8.080 ;
        RECT 27.050 7.080 27.210 7.530 ;
        RECT 25.220 6.480 25.460 6.640 ;
        RECT 16.980 4.830 17.210 6.120 ;
        RECT 25.210 5.490 25.450 6.130 ;
        RECT 26.240 5.880 26.400 6.740 ;
        RECT 26.630 6.620 26.800 6.740 ;
        RECT 26.640 5.880 26.800 6.620 ;
        RECT 26.940 6.530 27.210 7.080 ;
        RECT 26.940 6.480 27.220 6.530 ;
        RECT 27.050 6.390 27.220 6.480 ;
        RECT 27.050 5.880 27.210 6.390 ;
        RECT 25.220 5.230 25.450 5.490 ;
        RECT 25.220 5.010 25.460 5.230 ;
        RECT 25.240 4.650 25.560 4.970 ;
        RECT 26.240 4.870 26.400 5.730 ;
        RECT 26.640 4.990 26.800 5.730 ;
        RECT 27.050 5.220 27.210 5.730 ;
        RECT 27.050 5.130 27.220 5.220 ;
        RECT 26.630 4.870 26.800 4.990 ;
        RECT 26.240 4.820 26.450 4.870 ;
        RECT 26.220 4.580 26.450 4.820 ;
        RECT 26.240 4.560 26.440 4.580 ;
        RECT 25.240 4.100 25.560 4.420 ;
        RECT 26.240 3.830 26.400 4.560 ;
        RECT 26.610 3.880 26.800 4.870 ;
        RECT 26.940 5.080 27.220 5.130 ;
        RECT 26.940 4.530 27.210 5.080 ;
        RECT 27.050 3.830 27.210 4.530 ;
      LAYER via ;
        RECT 2.040 10.230 2.300 10.490 ;
        RECT 2.040 9.680 2.300 9.940 ;
        RECT 2.040 7.680 2.300 7.940 ;
        RECT 2.040 7.130 2.300 7.480 ;
        RECT 2.040 6.670 2.300 6.930 ;
        RECT 2.040 4.680 2.300 4.940 ;
        RECT 2.040 4.130 2.300 4.390 ;
        RECT 25.270 10.230 25.530 10.490 ;
        RECT 25.270 9.680 25.530 9.940 ;
        RECT 25.270 7.680 25.530 7.940 ;
        RECT 25.270 7.130 25.530 7.480 ;
        RECT 25.270 6.670 25.530 6.930 ;
        RECT 25.270 4.680 25.530 4.940 ;
        RECT 25.270 4.130 25.530 4.390 ;
      LAYER met2 ;
        RECT 2.020 10.240 2.330 10.530 ;
        RECT 0.000 10.200 2.330 10.240 ;
        RECT 25.240 10.240 25.550 10.530 ;
        RECT 25.240 10.200 27.570 10.240 ;
        RECT 0.000 10.060 2.180 10.200 ;
        RECT 25.390 10.060 27.570 10.200 ;
        RECT 2.020 9.810 2.330 9.980 ;
        RECT 0.000 9.650 2.330 9.810 ;
        RECT 0.000 9.630 2.170 9.650 ;
        RECT 2.470 9.630 2.560 9.810 ;
        RECT 5.360 9.760 12.240 9.830 ;
        RECT 5.330 9.650 12.240 9.760 ;
        RECT 15.330 9.760 22.210 9.830 ;
        RECT 25.240 9.810 25.550 9.980 ;
        RECT 15.330 9.650 22.240 9.760 ;
        RECT 25.010 9.630 25.100 9.810 ;
        RECT 25.240 9.650 27.570 9.810 ;
        RECT 25.400 9.630 27.570 9.650 ;
        RECT 3.230 9.220 12.240 9.400 ;
        RECT 15.330 9.220 24.340 9.400 ;
        RECT 5.360 8.340 12.240 8.400 ;
        RECT 5.330 8.220 12.240 8.340 ;
        RECT 15.330 8.340 22.210 8.400 ;
        RECT 15.330 8.220 22.240 8.340 ;
        RECT 0.000 7.970 2.170 7.990 ;
        RECT 0.000 7.810 2.330 7.970 ;
        RECT 2.470 7.810 2.560 7.990 ;
        RECT 5.370 7.900 12.240 7.970 ;
        RECT 2.020 7.640 2.330 7.810 ;
        RECT 5.330 7.790 12.240 7.900 ;
        RECT 15.330 7.900 22.200 7.970 ;
        RECT 15.330 7.790 22.240 7.900 ;
        RECT 25.010 7.810 25.100 7.990 ;
        RECT 25.400 7.970 27.570 7.990 ;
        RECT 25.240 7.810 27.570 7.970 ;
        RECT 25.240 7.640 25.550 7.810 ;
        RECT 0.000 7.520 2.180 7.560 ;
        RECT 25.390 7.520 27.570 7.560 ;
        RECT 0.000 7.380 2.330 7.520 ;
        RECT 2.020 7.230 2.330 7.380 ;
        RECT 0.000 7.090 2.330 7.230 ;
        RECT 25.240 7.380 27.570 7.520 ;
        RECT 25.240 7.230 25.550 7.380 ;
        RECT 25.240 7.090 27.570 7.230 ;
        RECT 0.000 7.050 2.180 7.090 ;
        RECT 25.390 7.050 27.570 7.090 ;
        RECT 2.020 6.800 2.330 6.970 ;
        RECT 0.000 6.640 2.330 6.800 ;
        RECT 0.000 6.620 2.170 6.640 ;
        RECT 2.470 6.620 2.560 6.800 ;
        RECT 5.330 6.640 12.240 6.810 ;
        RECT 15.330 6.640 22.240 6.810 ;
        RECT 25.240 6.800 25.550 6.970 ;
        RECT 25.010 6.620 25.100 6.800 ;
        RECT 25.240 6.640 27.570 6.800 ;
        RECT 25.400 6.620 27.570 6.640 ;
        RECT 5.330 6.220 12.240 6.390 ;
        RECT 15.330 6.220 22.240 6.390 ;
        RECT 5.330 5.240 12.240 5.410 ;
        RECT 15.330 5.240 22.240 5.410 ;
        RECT 0.000 4.970 2.170 4.990 ;
        RECT 0.000 4.810 2.330 4.970 ;
        RECT 2.470 4.810 2.560 4.990 ;
        RECT 2.020 4.640 2.330 4.810 ;
        RECT 5.330 4.800 12.240 4.970 ;
        RECT 15.330 4.800 22.240 4.970 ;
        RECT 25.010 4.810 25.100 4.990 ;
        RECT 25.400 4.970 27.570 4.990 ;
        RECT 25.240 4.810 27.570 4.970 ;
        RECT 25.240 4.640 25.550 4.810 ;
        RECT 0.000 4.420 2.180 4.560 ;
        RECT 25.390 4.420 27.570 4.560 ;
        RECT 0.000 4.380 2.330 4.420 ;
        RECT 2.020 4.090 2.330 4.380 ;
        RECT 25.240 4.380 27.570 4.420 ;
        RECT 25.240 4.090 25.550 4.380 ;
        RECT 7.200 3.610 7.320 3.690 ;
        RECT 20.290 3.550 20.410 3.690 ;
  END
END sky130_hilas_swc4x2cellOverlap

MACRO sky130_hilas_FGBias2x1cell
  CLASS CORE ;
  FOREIGN sky130_hilas_FGBias2x1cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.540 BY 10.520 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VTUN
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 0.350 0.470 0.770 6.520 ;
    END
  END VTUN
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2.830 3.660 3.060 6.520 ;
        RECT 2.830 3.370 3.160 3.660 ;
        RECT 2.830 0.470 3.060 3.370 ;
    END
  END VGND
  PIN GATE_CONTROL
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 4.050 0.470 4.280 6.520 ;
    END
  END GATE_CONTROL
  PIN DRAIN1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 5.840 9.120 6.020 ;
    END
  END DRAIN1
  PIN DRAIN4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 9.060 1.140 9.220 1.160 ;
        RECT 0.000 1.090 9.220 1.140 ;
        RECT 0.000 0.990 9.100 1.090 ;
    END
  END DRAIN4
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 11.170 3.660 11.490 3.740 ;
        RECT 10.180 3.480 11.490 3.660 ;
        RECT 10.180 3.310 11.360 3.480 ;
        RECT 10.230 3.160 10.550 3.310 ;
    END
  END VINJ
  PIN OUTPUT1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 9.340 5.000 9.650 5.220 ;
        RECT 9.340 4.890 11.530 5.000 ;
        RECT 9.500 4.780 11.530 4.890 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 9.340 2.240 9.650 2.460 ;
        RECT 9.340 2.130 11.530 2.240 ;
        RECT 9.490 2.030 11.530 2.130 ;
    END
  END OUTPUT2
  PIN GATECOL
    PORT
      LAYER met1 ;
        RECT 10.570 6.480 10.760 6.520 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.570 0.470 10.760 0.520 ;
    END
  END GATECOL
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 11.010 3.770 11.290 6.520 ;
        RECT 11.010 3.450 11.460 3.770 ;
        RECT 11.010 0.470 11.290 3.450 ;
      LAYER via ;
        RECT 11.200 3.480 11.460 3.740 ;
    END
  END VINJ
  OBS
      LAYER nwell ;
        RECT 14.520 10.180 16.250 10.520 ;
        RECT 14.500 8.620 16.250 10.180 ;
        RECT 14.500 6.990 16.230 8.620 ;
        RECT 12.990 6.600 16.290 6.990 ;
        RECT 12.990 6.560 16.530 6.600 ;
        RECT 8.230 6.510 11.530 6.520 ;
        RECT 10.570 6.480 10.760 6.510 ;
        RECT 12.990 4.910 16.540 6.560 ;
        RECT 0.590 1.870 1.150 4.290 ;
        RECT 12.990 3.820 16.290 4.910 ;
        RECT 12.990 1.980 16.290 3.170 ;
        RECT 12.990 0.330 16.540 1.980 ;
        RECT 12.990 0.290 16.530 0.330 ;
        RECT 12.990 0.000 16.290 0.290 ;
      LAYER li1 ;
        RECT 14.920 8.790 15.470 9.220 ;
        RECT 14.920 7.060 15.470 7.490 ;
        RECT 13.880 6.360 14.410 6.530 ;
        RECT 15.690 6.260 15.890 6.610 ;
        RECT 15.690 6.230 15.900 6.260 ;
        RECT 14.120 5.430 14.350 6.120 ;
        RECT 9.350 5.140 9.670 5.180 ;
        RECT 9.350 4.950 9.680 5.140 ;
        RECT 9.350 4.920 9.670 4.950 ;
        RECT 14.130 4.280 14.300 5.430 ;
        RECT 14.960 4.370 15.130 5.980 ;
        RECT 15.680 5.650 15.900 6.230 ;
        RECT 15.690 5.640 15.900 5.650 ;
        RECT 15.330 5.470 15.520 5.480 ;
        RECT 15.330 5.180 15.530 5.470 ;
        RECT 15.320 4.850 15.610 5.180 ;
        RECT 14.960 4.180 15.140 4.370 ;
        RECT 3.040 3.630 3.230 3.950 ;
        RECT 2.950 3.540 3.230 3.630 ;
        RECT 2.950 3.400 6.590 3.540 ;
        RECT 3.040 3.360 6.590 3.400 ;
        RECT 3.040 2.940 3.230 3.360 ;
        RECT 9.350 2.380 9.670 2.420 ;
        RECT 4.070 2.320 4.300 2.360 ;
        RECT 9.350 2.190 9.680 2.380 ;
        RECT 9.350 2.160 9.670 2.190 ;
        RECT 14.130 1.460 14.300 2.710 ;
        RECT 14.960 2.620 15.140 2.810 ;
        RECT 14.120 0.770 14.350 1.460 ;
        RECT 14.960 1.010 15.130 2.620 ;
        RECT 15.320 1.810 15.610 2.140 ;
        RECT 15.330 1.520 15.530 1.810 ;
        RECT 15.330 1.510 15.520 1.520 ;
        RECT 15.690 1.340 15.900 1.350 ;
        RECT 15.680 0.760 15.900 1.340 ;
        RECT 15.690 0.730 15.900 0.760 ;
        RECT 13.880 0.460 14.410 0.630 ;
        RECT 15.690 0.380 15.890 0.730 ;
      LAYER mcon ;
        RECT 14.920 8.870 15.190 9.140 ;
        RECT 14.920 7.140 15.190 7.410 ;
        RECT 14.150 5.910 14.320 6.080 ;
        RECT 15.700 6.060 15.870 6.230 ;
        RECT 14.150 5.460 14.320 5.630 ;
        RECT 9.410 4.960 9.580 5.130 ;
        RECT 15.340 5.220 15.520 5.410 ;
        RECT 2.960 3.430 3.130 3.600 ;
        RECT 9.410 2.200 9.580 2.370 ;
        RECT 14.150 1.260 14.320 1.430 ;
        RECT 15.340 1.580 15.520 1.770 ;
        RECT 14.150 0.810 14.320 0.980 ;
        RECT 15.700 0.760 15.870 0.930 ;
      LAYER met1 ;
        RECT 14.860 6.600 15.250 10.190 ;
        RECT 13.810 6.170 14.120 6.560 ;
        RECT 13.810 6.120 14.360 6.170 ;
        RECT 14.100 5.380 14.360 6.120 ;
        RECT 15.330 5.480 15.520 6.930 ;
        RECT 15.770 6.290 15.930 6.930 ;
        RECT 15.660 5.740 15.930 6.290 ;
        RECT 15.660 5.690 15.940 5.740 ;
        RECT 15.770 5.600 15.940 5.690 ;
        RECT 15.330 5.450 15.550 5.480 ;
        RECT 9.340 4.890 9.660 5.210 ;
        RECT 15.310 5.180 15.560 5.450 ;
        RECT 15.320 5.170 15.560 5.180 ;
        RECT 15.320 4.930 15.550 5.170 ;
        RECT 14.930 4.120 15.170 4.500 ;
        RECT 10.260 3.730 10.520 4.050 ;
        RECT 15.360 3.910 15.520 4.930 ;
        RECT 15.770 3.910 15.930 5.600 ;
        RECT 10.260 3.130 10.520 3.450 ;
        RECT 14.930 2.490 15.170 2.870 ;
        RECT 9.340 2.130 9.660 2.450 ;
        RECT 15.360 2.060 15.520 3.080 ;
        RECT 15.320 1.820 15.550 2.060 ;
        RECT 15.320 1.810 15.560 1.820 ;
        RECT 15.310 1.540 15.560 1.810 ;
        RECT 15.330 1.510 15.550 1.540 ;
        RECT 14.100 0.870 14.360 1.510 ;
        RECT 13.810 0.720 14.360 0.870 ;
        RECT 13.810 0.430 14.120 0.720 ;
        RECT 15.330 0.060 15.520 1.510 ;
        RECT 15.770 1.390 15.930 3.080 ;
        RECT 15.770 1.300 15.940 1.390 ;
        RECT 15.660 1.250 15.940 1.300 ;
        RECT 15.660 0.700 15.930 1.250 ;
        RECT 15.770 0.060 15.930 0.700 ;
      LAYER via ;
        RECT 13.840 6.150 14.100 6.410 ;
        RECT 9.370 4.920 9.630 5.180 ;
        RECT 10.260 3.760 10.520 4.020 ;
        RECT 10.260 3.160 10.520 3.420 ;
        RECT 9.370 2.160 9.630 2.420 ;
        RECT 13.840 0.580 14.100 0.840 ;
      LAYER met2 ;
        RECT 13.810 6.440 14.120 6.450 ;
        RECT 13.810 6.260 16.290 6.440 ;
        RECT 13.810 6.120 14.120 6.260 ;
        RECT 10.230 3.760 10.550 4.020 ;
        RECT 13.810 0.730 14.120 0.870 ;
        RECT 13.810 0.550 16.290 0.730 ;
        RECT 13.810 0.540 14.120 0.550 ;
  END
END sky130_hilas_FGBias2x1cell

MACRO sky130_hilas_drainSelect01
  CLASS CORE ;
  FOREIGN sky130_hilas_drainSelect01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.000 BY 6.110 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DRAIN3
    PORT
      LAYER met2 ;
        RECT 0.000 2.590 0.570 2.600 ;
        RECT 0.000 2.580 1.270 2.590 ;
        RECT 0.000 2.420 2.000 2.580 ;
    END
  END DRAIN3
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.580 6.040 0.830 6.110 ;
    END
  END VINJ
  PIN DRAIN_MUX
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 3.570 6.040 3.800 6.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.570 0.060 3.800 0.140 ;
    END
  END DRAIN_MUX
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 4.920 0.060 5.110 0.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.920 6.060 5.110 6.110 ;
    END
  END VGND
  PIN SELECT2
    ANTENNADIFFAREA 0.322600 ;
    PORT
      LAYER met2 ;
        RECT 4.070 4.000 4.390 4.050 ;
        RECT 5.570 4.000 5.720 4.080 ;
        RECT 6.480 4.000 6.800 4.080 ;
        RECT 4.070 3.810 6.800 4.000 ;
        RECT 4.070 3.790 4.390 3.810 ;
        RECT 6.480 3.760 6.800 3.810 ;
    END
  END SELECT2
  PIN SELECT1
    ANTENNADIFFAREA 0.322600 ;
    PORT
      LAYER met2 ;
        RECT 4.070 5.440 4.390 5.460 ;
        RECT 6.480 5.440 6.800 5.490 ;
        RECT 4.070 5.250 6.800 5.440 ;
        RECT 4.070 5.200 4.390 5.250 ;
        RECT 5.640 5.180 5.720 5.250 ;
        RECT 6.480 5.170 6.800 5.250 ;
    END
  END SELECT1
  PIN SELECT3
    ANTENNADIFFAREA 0.322600 ;
    PORT
      LAYER met2 ;
        RECT 4.070 2.240 4.390 2.260 ;
        RECT 6.480 2.240 6.800 2.290 ;
        RECT 4.070 2.050 6.800 2.240 ;
        RECT 4.070 2.000 4.390 2.050 ;
        RECT 5.640 1.980 5.720 2.050 ;
        RECT 6.480 1.970 6.800 2.050 ;
    END
  END SELECT3
  PIN SELECT4
    ANTENNADIFFAREA 0.322600 ;
    PORT
      LAYER met2 ;
        RECT 4.070 0.800 4.390 0.850 ;
        RECT 5.630 0.800 5.720 0.870 ;
        RECT 6.480 0.800 6.800 0.880 ;
        RECT 4.070 0.610 6.800 0.800 ;
        RECT 4.070 0.590 4.390 0.610 ;
        RECT 6.480 0.560 6.800 0.610 ;
    END
  END SELECT4
  OBS
      LAYER nwell ;
        RECT 2.320 4.630 5.740 5.870 ;
        RECT 0.000 4.620 5.740 4.630 ;
        RECT 2.320 3.380 5.740 4.620 ;
        RECT 2.320 1.430 5.740 2.670 ;
        RECT 0.000 1.410 5.740 1.430 ;
        RECT 2.320 0.180 5.740 1.410 ;
      LAYER li1 ;
        RECT 2.540 5.010 2.710 5.540 ;
        RECT 2.540 4.240 2.720 5.010 ;
        RECT 2.540 3.710 2.710 4.240 ;
        RECT 2.940 3.760 3.110 5.490 ;
        RECT 6.630 5.420 6.870 5.450 ;
        RECT 3.640 5.250 4.600 5.420 ;
        RECT 5.050 5.250 6.390 5.420 ;
        RECT 6.630 5.250 7.200 5.420 ;
        RECT 3.920 5.240 4.090 5.250 ;
        RECT 6.630 5.210 6.870 5.250 ;
        RECT 7.510 5.120 7.680 5.540 ;
        RECT 4.120 4.800 4.460 4.980 ;
        RECT 7.580 4.900 7.750 4.940 ;
        RECT 3.640 4.630 6.390 4.800 ;
        RECT 6.850 4.630 7.220 4.800 ;
        RECT 3.640 4.450 6.390 4.620 ;
        RECT 6.850 4.450 7.220 4.620 ;
        RECT 7.320 4.510 7.510 4.740 ;
        RECT 7.580 4.730 7.810 4.900 ;
        RECT 7.580 4.520 7.750 4.730 ;
        RECT 4.120 4.270 4.460 4.450 ;
        RECT 7.580 4.350 7.810 4.520 ;
        RECT 7.580 4.310 7.750 4.350 ;
        RECT 3.920 4.000 4.090 4.010 ;
        RECT 6.630 4.000 6.870 4.040 ;
        RECT 3.640 3.830 4.600 4.000 ;
        RECT 5.050 3.830 6.390 4.000 ;
        RECT 6.630 3.830 7.200 4.000 ;
        RECT 6.630 3.800 6.870 3.830 ;
        RECT 7.510 3.710 7.680 4.130 ;
        RECT 2.540 1.810 2.710 2.340 ;
        RECT 2.540 1.040 2.720 1.810 ;
        RECT 2.540 0.510 2.710 1.040 ;
        RECT 2.940 0.560 3.110 2.290 ;
        RECT 6.630 2.220 6.870 2.250 ;
        RECT 3.640 2.050 4.600 2.220 ;
        RECT 5.050 2.050 6.390 2.220 ;
        RECT 6.630 2.050 7.200 2.220 ;
        RECT 3.920 2.040 4.090 2.050 ;
        RECT 6.630 2.010 6.870 2.050 ;
        RECT 7.510 1.920 7.680 2.340 ;
        RECT 4.120 1.600 4.460 1.780 ;
        RECT 7.580 1.700 7.750 1.740 ;
        RECT 3.640 1.430 6.390 1.600 ;
        RECT 6.850 1.430 7.220 1.600 ;
        RECT 3.640 1.250 6.390 1.420 ;
        RECT 6.850 1.250 7.220 1.420 ;
        RECT 7.320 1.310 7.510 1.540 ;
        RECT 7.580 1.530 7.810 1.700 ;
        RECT 7.580 1.320 7.750 1.530 ;
        RECT 4.120 1.070 4.460 1.250 ;
        RECT 7.580 1.150 7.810 1.320 ;
        RECT 7.580 1.110 7.750 1.150 ;
        RECT 3.920 0.800 4.090 0.810 ;
        RECT 6.630 0.800 6.870 0.840 ;
        RECT 3.640 0.630 4.600 0.800 ;
        RECT 5.050 0.630 6.390 0.800 ;
        RECT 6.630 0.630 7.200 0.800 ;
        RECT 6.630 0.600 6.870 0.630 ;
        RECT 7.510 0.510 7.680 0.930 ;
      LAYER mcon ;
        RECT 2.540 5.370 2.710 5.540 ;
        RECT 5.920 5.250 6.090 5.420 ;
        RECT 6.670 5.250 6.840 5.420 ;
        RECT 7.510 5.370 7.680 5.540 ;
        RECT 2.940 4.920 3.110 5.090 ;
        RECT 7.330 4.540 7.500 4.710 ;
        RECT 7.640 4.730 7.810 4.900 ;
        RECT 2.540 4.070 2.710 4.240 ;
        RECT 2.940 4.160 3.110 4.330 ;
        RECT 7.640 4.350 7.810 4.520 ;
        RECT 3.920 3.840 4.090 4.010 ;
        RECT 5.920 3.830 6.090 4.000 ;
        RECT 6.670 3.830 6.840 4.000 ;
        RECT 2.540 2.170 2.710 2.340 ;
        RECT 5.920 2.050 6.090 2.220 ;
        RECT 6.670 2.050 6.840 2.220 ;
        RECT 7.510 2.170 7.680 2.340 ;
        RECT 2.940 1.720 3.110 1.890 ;
        RECT 7.330 1.340 7.500 1.510 ;
        RECT 7.640 1.530 7.810 1.700 ;
        RECT 2.540 0.870 2.710 1.040 ;
        RECT 2.940 0.960 3.110 1.130 ;
        RECT 7.640 1.150 7.810 1.320 ;
        RECT 3.920 0.640 4.090 0.810 ;
        RECT 5.920 0.630 6.090 0.800 ;
        RECT 6.670 0.630 6.840 0.800 ;
      LAYER met1 ;
        RECT 2.900 5.600 3.150 5.820 ;
        RECT 2.510 5.530 3.150 5.600 ;
        RECT 2.500 5.170 3.150 5.530 ;
        RECT 4.050 5.440 4.390 5.490 ;
        RECT 3.830 5.420 4.390 5.440 ;
        RECT 3.830 5.250 4.510 5.420 ;
        RECT 3.830 5.210 4.390 5.250 ;
        RECT 4.050 5.170 4.390 5.210 ;
        RECT 0.580 4.620 0.830 4.630 ;
        RECT 2.510 4.080 3.150 5.170 ;
        RECT 2.500 3.720 3.150 4.080 ;
        RECT 4.050 4.040 4.390 4.080 ;
        RECT 3.830 4.000 4.390 4.040 ;
        RECT 3.830 3.830 4.510 4.000 ;
        RECT 3.830 3.810 4.390 3.830 ;
        RECT 4.050 3.760 4.390 3.810 ;
        RECT 2.510 3.650 3.150 3.720 ;
        RECT 2.900 3.430 3.150 3.650 ;
        RECT 5.890 3.430 6.120 5.820 ;
        RECT 7.240 5.600 7.430 5.820 ;
        RECT 6.480 5.460 6.850 5.480 ;
        RECT 6.480 5.200 6.900 5.460 ;
        RECT 6.480 5.190 6.850 5.200 ;
        RECT 7.240 5.110 7.710 5.600 ;
        RECT 7.240 4.770 7.430 5.110 ;
        RECT 7.240 4.480 7.530 4.770 ;
        RECT 7.570 4.670 7.890 4.950 ;
        RECT 7.240 4.140 7.430 4.480 ;
        RECT 7.570 4.300 7.890 4.580 ;
        RECT 6.480 4.050 6.850 4.060 ;
        RECT 6.480 3.790 6.900 4.050 ;
        RECT 6.480 3.770 6.850 3.790 ;
        RECT 7.240 3.650 7.710 4.140 ;
        RECT 7.240 3.430 7.430 3.650 ;
        RECT 2.900 2.400 3.150 2.620 ;
        RECT 2.510 2.330 3.150 2.400 ;
        RECT 2.500 1.970 3.150 2.330 ;
        RECT 4.050 2.240 4.390 2.290 ;
        RECT 3.830 2.220 4.390 2.240 ;
        RECT 3.830 2.050 4.510 2.220 ;
        RECT 3.830 2.010 4.390 2.050 ;
        RECT 4.050 1.970 4.390 2.010 ;
        RECT 0.580 1.420 0.830 1.430 ;
        RECT 2.510 0.880 3.150 1.970 ;
        RECT 2.500 0.520 3.150 0.880 ;
        RECT 4.050 0.840 4.390 0.880 ;
        RECT 3.830 0.800 4.390 0.840 ;
        RECT 3.830 0.630 4.510 0.800 ;
        RECT 3.830 0.610 4.390 0.630 ;
        RECT 4.050 0.560 4.390 0.610 ;
        RECT 2.510 0.450 3.150 0.520 ;
        RECT 2.900 0.230 3.150 0.450 ;
        RECT 5.890 0.230 6.120 2.620 ;
        RECT 7.240 2.400 7.430 2.620 ;
        RECT 6.480 2.260 6.850 2.280 ;
        RECT 6.480 2.000 6.900 2.260 ;
        RECT 6.480 1.990 6.850 2.000 ;
        RECT 7.240 1.910 7.710 2.400 ;
        RECT 7.240 1.570 7.430 1.910 ;
        RECT 7.240 1.280 7.530 1.570 ;
        RECT 7.570 1.470 7.890 1.750 ;
        RECT 7.240 0.940 7.430 1.280 ;
        RECT 7.570 1.100 7.890 1.380 ;
        RECT 6.480 0.850 6.850 0.860 ;
        RECT 6.480 0.590 6.900 0.850 ;
        RECT 6.480 0.570 6.850 0.590 ;
        RECT 7.240 0.450 7.710 0.940 ;
        RECT 7.240 0.230 7.430 0.450 ;
      LAYER via ;
        RECT 4.100 5.200 4.360 5.460 ;
        RECT 4.100 3.790 4.360 4.050 ;
        RECT 6.510 5.200 6.770 5.460 ;
        RECT 7.600 4.680 7.860 4.940 ;
        RECT 7.600 4.310 7.860 4.570 ;
        RECT 6.510 3.790 6.770 4.050 ;
        RECT 4.100 2.000 4.360 2.260 ;
        RECT 4.100 0.590 4.360 0.850 ;
        RECT 6.510 2.000 6.770 2.260 ;
        RECT 7.600 1.480 7.860 1.740 ;
        RECT 7.600 1.110 7.860 1.370 ;
        RECT 6.510 0.590 6.770 0.850 ;
      LAYER met2 ;
        RECT 0.000 5.680 1.780 5.860 ;
        RECT 7.560 4.730 8.000 4.960 ;
        RECT 7.560 4.660 7.900 4.730 ;
        RECT 7.560 4.520 7.900 4.590 ;
        RECT 7.560 4.290 8.000 4.520 ;
        RECT 0.000 3.380 1.780 3.540 ;
        RECT 7.560 1.530 8.000 1.760 ;
        RECT 7.560 1.460 7.900 1.530 ;
        RECT 7.560 1.320 7.900 1.390 ;
        RECT 7.560 1.090 8.000 1.320 ;
        RECT 0.000 0.160 1.780 0.330 ;
  END
END sky130_hilas_drainSelect01

MACRO sky130_hilas_DAC5bit01
  CLASS CORE ;
  FOREIGN sky130_hilas_DAC5bit01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.580 BY 7.990 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 8.350 0.980 8.670 1.110 ;
        RECT 0.000 0.850 8.670 0.980 ;
        RECT 0.000 0.780 8.540 0.850 ;
    END
  END A0
  PIN A1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 11.710 2.100 11.860 5.840 ;
        RECT 0.000 1.900 11.870 2.100 ;
        RECT 0.000 1.890 0.140 1.900 ;
    END
  END A1
  PIN A2
    USE ANALOG ;
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER met2 ;
        RECT 10.110 3.080 10.310 5.680 ;
        RECT 0.000 2.870 10.310 3.080 ;
        RECT 0.320 2.670 0.640 2.870 ;
    END
  END A2
  PIN A3
    USE ANALOG ;
    ANTENNAGATEAREA 0.307500 ;
    PORT
      LAYER met2 ;
        RECT 0.000 4.950 2.060 5.010 ;
        RECT 3.480 4.950 3.700 5.410 ;
        RECT 8.400 4.960 8.650 5.720 ;
        RECT 8.400 4.950 8.680 4.960 ;
        RECT 0.000 4.800 8.680 4.950 ;
        RECT 0.260 4.560 0.620 4.800 ;
        RECT 1.900 4.650 8.680 4.800 ;
    END
  END A3
  PIN A4
    USE ANALOG ;
    ANTENNAGATEAREA 6.324800 ;
    ANTENNADIFFAREA 0.522900 ;
    PORT
      LAYER met2 ;
        RECT 0.320 5.960 0.640 6.190 ;
        RECT 2.030 5.960 2.350 6.230 ;
        RECT 5.230 5.960 5.550 6.230 ;
        RECT 6.840 5.960 7.160 6.240 ;
        RECT 0.000 5.920 7.160 5.960 ;
        RECT 0.000 5.770 7.050 5.920 ;
        RECT 8.460 5.910 8.780 6.230 ;
        RECT 10.070 5.920 10.390 6.240 ;
        RECT 11.680 5.920 12.000 6.240 ;
        RECT 0.000 5.750 0.290 5.770 ;
        RECT 3.750 5.150 4.070 5.470 ;
    END
  END A4
  PIN VPWR
    USE ANALOG ;
    ANTENNADIFFAREA 2.316600 ;
    PORT
      LAYER met2 ;
        RECT 12.970 5.960 13.280 5.980 ;
        RECT 13.640 5.960 13.950 5.980 ;
        RECT 12.710 5.680 13.950 5.960 ;
        RECT 12.970 5.650 13.280 5.680 ;
        RECT 13.460 5.670 13.950 5.680 ;
        RECT 13.640 5.650 13.950 5.670 ;
    END
  END VPWR
  PIN OUT
    USE ANALOG ;
    ANTENNADIFFAREA 0.947700 ;
    PORT
      LAYER met1 ;
        RECT 3.110 0.230 3.340 0.360 ;
        RECT 4.730 0.230 4.960 0.360 ;
        RECT 6.330 0.230 6.560 0.360 ;
        RECT 7.950 0.230 8.180 0.360 ;
        RECT 9.550 0.230 9.780 0.360 ;
        RECT 11.170 0.230 11.400 0.360 ;
        RECT 12.770 0.230 13.000 0.360 ;
        RECT 14.380 0.230 14.610 0.360 ;
        RECT 3.040 0.000 16.580 0.230 ;
    END
  END OUT
  OBS
      LAYER nwell ;
        RECT 0.270 7.030 1.880 7.990 ;
        RECT 1.890 7.030 16.370 7.990 ;
        RECT 0.270 5.820 16.370 7.030 ;
        RECT 0.270 5.110 6.710 5.820 ;
        RECT 6.770 5.360 16.370 5.820 ;
        RECT 8.320 5.110 16.370 5.360 ;
        RECT 0.270 2.940 16.370 5.110 ;
        RECT 0.270 1.980 1.880 2.830 ;
        RECT 1.890 1.980 16.370 2.830 ;
      LAYER li1 ;
        RECT 2.260 6.440 2.430 6.770 ;
        RECT 2.940 6.440 3.110 6.770 ;
        RECT 3.870 6.440 4.040 6.770 ;
        RECT 4.550 6.440 4.720 6.770 ;
        RECT 5.480 6.440 5.650 6.770 ;
        RECT 6.160 6.440 6.330 6.770 ;
        RECT 6.770 6.290 6.980 6.720 ;
        RECT 7.090 6.440 7.260 6.770 ;
        RECT 7.770 6.440 7.940 6.770 ;
        RECT 8.700 6.440 8.870 6.770 ;
        RECT 9.380 6.440 9.550 6.770 ;
        RECT 10.310 6.440 10.480 6.770 ;
        RECT 10.990 6.440 11.160 6.770 ;
        RECT 11.920 6.440 12.090 6.770 ;
        RECT 12.600 6.440 12.770 6.770 ;
        RECT 13.530 6.440 13.700 6.770 ;
        RECT 14.210 6.440 14.380 6.770 ;
        RECT 6.790 6.270 6.960 6.290 ;
        RECT 0.370 5.720 0.580 6.150 ;
        RECT 2.080 5.810 2.290 6.190 ;
        RECT 5.280 5.810 5.490 6.190 ;
        RECT 2.080 5.760 2.430 5.810 ;
        RECT 2.100 5.740 2.430 5.760 ;
        RECT 0.390 5.700 0.560 5.720 ;
        RECT 2.260 5.480 2.430 5.740 ;
        RECT 2.940 5.480 3.110 5.810 ;
        RECT 3.870 5.480 4.040 5.810 ;
        RECT 4.550 5.480 4.720 5.810 ;
        RECT 5.280 5.760 5.650 5.810 ;
        RECT 5.300 5.740 5.470 5.760 ;
        RECT 5.480 5.480 5.650 5.760 ;
        RECT 6.160 5.480 6.330 5.810 ;
        RECT 6.890 5.770 7.100 6.200 ;
        RECT 7.150 5.980 7.320 6.310 ;
        RECT 7.830 5.980 8.000 6.310 ;
        RECT 8.510 5.810 8.720 6.190 ;
        RECT 10.120 5.810 10.330 6.200 ;
        RECT 11.730 5.810 11.940 6.200 ;
        RECT 12.980 5.900 13.300 5.940 ;
        RECT 13.650 5.900 13.970 5.940 ;
        RECT 6.910 5.750 7.080 5.770 ;
        RECT 8.510 5.760 8.870 5.810 ;
        RECT 8.530 5.740 8.870 5.760 ;
        RECT 8.700 5.480 8.870 5.740 ;
        RECT 9.380 5.480 9.550 5.810 ;
        RECT 10.120 5.770 10.480 5.810 ;
        RECT 10.140 5.750 10.480 5.770 ;
        RECT 10.310 5.480 10.480 5.750 ;
        RECT 10.990 5.480 11.160 5.810 ;
        RECT 11.730 5.770 12.090 5.810 ;
        RECT 11.750 5.750 12.090 5.770 ;
        RECT 11.920 5.480 12.090 5.750 ;
        RECT 12.600 5.480 12.770 5.810 ;
        RECT 12.980 5.800 13.310 5.900 ;
        RECT 13.650 5.810 13.980 5.900 ;
        RECT 12.950 5.710 13.310 5.800 ;
        RECT 13.530 5.710 13.980 5.810 ;
        RECT 12.950 5.680 13.300 5.710 ;
        RECT 13.530 5.680 13.970 5.710 ;
        RECT 3.600 5.400 4.030 5.420 ;
        RECT 3.580 5.230 4.030 5.400 ;
        RECT 8.370 5.290 8.540 5.310 ;
        RECT 3.600 5.210 4.030 5.230 ;
        RECT 3.980 5.020 4.150 5.030 ;
        RECT 8.350 5.020 8.560 5.290 ;
        RECT 12.950 5.020 13.160 5.680 ;
        RECT 13.530 5.480 13.790 5.680 ;
        RECT 14.210 5.480 14.380 5.810 ;
        RECT 13.620 5.020 13.790 5.480 ;
        RECT 2.370 4.850 13.800 5.020 ;
        RECT 0.350 4.410 0.560 4.840 ;
        RECT 2.260 4.790 13.800 4.850 ;
        RECT 2.260 4.520 2.540 4.790 ;
        RECT 2.940 4.520 3.110 4.790 ;
        RECT 3.870 4.520 4.150 4.790 ;
        RECT 4.550 4.520 4.720 4.790 ;
        RECT 5.480 4.520 5.740 4.790 ;
        RECT 6.160 4.520 6.330 4.790 ;
        RECT 7.090 4.520 7.360 4.790 ;
        RECT 7.770 4.520 7.940 4.790 ;
        RECT 0.370 4.390 0.540 4.410 ;
        RECT 2.370 3.890 2.540 4.520 ;
        RECT 3.030 3.890 3.200 4.460 ;
        RECT 3.980 3.890 4.150 4.520 ;
        RECT 4.660 3.890 4.830 4.420 ;
        RECT 5.570 3.890 5.740 4.520 ;
        RECT 6.260 3.890 6.430 4.500 ;
        RECT 7.190 3.890 7.360 4.520 ;
        RECT 7.880 3.890 8.050 4.450 ;
        RECT 8.810 3.890 8.980 4.790 ;
        RECT 10.310 4.520 10.580 4.790 ;
        RECT 10.990 4.520 11.160 4.790 ;
        RECT 11.920 4.520 12.190 4.790 ;
        RECT 12.600 4.520 12.770 4.790 ;
        RECT 13.530 4.520 13.800 4.790 ;
        RECT 14.210 4.660 14.380 4.850 ;
        RECT 14.210 4.520 14.480 4.660 ;
        RECT 9.480 3.890 9.650 4.500 ;
        RECT 9.930 4.000 10.140 4.430 ;
        RECT 9.950 3.980 10.120 4.000 ;
        RECT 10.410 3.890 10.580 4.520 ;
        RECT 11.100 3.890 11.270 4.500 ;
        RECT 12.020 3.890 12.190 4.520 ;
        RECT 12.700 3.890 12.870 4.480 ;
        RECT 13.630 3.890 13.800 4.520 ;
        RECT 14.310 3.890 14.480 4.520 ;
        RECT 0.370 3.460 0.580 3.890 ;
        RECT 2.260 3.560 2.540 3.890 ;
        RECT 2.940 3.560 3.200 3.890 ;
        RECT 3.870 3.560 4.150 3.890 ;
        RECT 4.550 3.560 4.830 3.890 ;
        RECT 5.480 3.560 5.740 3.890 ;
        RECT 6.160 3.560 6.430 3.890 ;
        RECT 7.090 3.560 7.360 3.890 ;
        RECT 7.770 3.560 8.050 3.890 ;
        RECT 8.700 3.560 8.980 3.890 ;
        RECT 9.380 3.560 9.650 3.890 ;
        RECT 10.310 3.560 10.580 3.890 ;
        RECT 10.990 3.560 11.270 3.890 ;
        RECT 11.920 3.560 12.190 3.890 ;
        RECT 12.600 3.560 12.870 3.890 ;
        RECT 13.530 3.560 13.800 3.890 ;
        RECT 14.210 3.560 14.480 3.890 ;
        RECT 0.390 3.440 0.560 3.460 ;
        RECT 0.370 2.520 0.580 2.950 ;
        RECT 0.390 2.500 0.560 2.520 ;
        RECT 2.370 1.230 2.540 3.560 ;
        RECT 3.030 0.330 3.200 3.560 ;
        RECT 3.980 1.230 4.150 3.560 ;
        RECT 4.660 0.330 4.830 3.560 ;
        RECT 5.570 1.230 5.740 3.560 ;
        RECT 6.260 0.330 6.430 3.560 ;
        RECT 7.190 1.230 7.360 3.560 ;
        RECT 7.880 0.330 8.050 3.560 ;
        RECT 8.810 1.250 8.980 3.560 ;
        RECT 9.480 0.330 9.650 3.560 ;
        RECT 10.410 1.260 10.580 3.560 ;
        RECT 11.100 0.330 11.270 3.560 ;
        RECT 12.020 1.250 12.190 3.560 ;
        RECT 12.700 0.330 12.870 3.560 ;
        RECT 13.630 1.220 13.800 3.560 ;
        RECT 14.310 0.330 14.480 3.560 ;
        RECT 3.030 0.100 3.320 0.330 ;
        RECT 4.660 0.100 4.940 0.330 ;
        RECT 6.260 0.100 6.540 0.330 ;
        RECT 7.880 0.100 8.160 0.330 ;
        RECT 9.480 0.100 9.760 0.330 ;
        RECT 11.100 0.100 11.380 0.330 ;
        RECT 12.700 0.100 12.980 0.330 ;
        RECT 14.310 0.100 14.590 0.330 ;
        RECT 3.030 0.000 3.200 0.100 ;
        RECT 4.660 0.000 4.830 0.100 ;
        RECT 6.260 0.000 6.430 0.100 ;
        RECT 7.880 0.000 8.050 0.100 ;
        RECT 9.480 0.000 9.650 0.100 ;
        RECT 11.100 0.000 11.270 0.100 ;
        RECT 12.700 0.000 12.870 0.100 ;
        RECT 14.310 0.000 14.480 0.100 ;
      LAYER mcon ;
        RECT 13.040 5.720 13.210 5.890 ;
        RECT 13.710 5.720 13.880 5.890 ;
        RECT 8.370 5.140 8.540 5.310 ;
        RECT 3.140 0.130 3.310 0.300 ;
        RECT 4.760 0.130 4.930 0.300 ;
        RECT 6.360 0.130 6.530 0.300 ;
        RECT 7.980 0.130 8.150 0.300 ;
        RECT 9.580 0.130 9.750 0.300 ;
        RECT 11.200 0.130 11.370 0.300 ;
        RECT 12.800 0.130 12.970 0.300 ;
        RECT 14.410 0.130 14.580 0.300 ;
      LAYER met1 ;
        RECT 6.770 6.500 6.990 6.720 ;
        RECT 6.760 6.240 6.990 6.500 ;
        RECT 0.320 5.870 0.640 6.190 ;
        RECT 2.030 5.910 2.350 6.230 ;
        RECT 5.230 5.910 5.550 6.230 ;
        RECT 6.760 6.210 7.160 6.240 ;
        RECT 6.840 5.920 7.160 6.210 ;
        RECT 0.360 5.640 0.590 5.870 ;
        RECT 2.070 5.680 2.300 5.910 ;
        RECT 5.270 5.680 5.500 5.910 ;
        RECT 6.880 5.690 7.110 5.920 ;
        RECT 8.460 5.910 8.780 6.230 ;
        RECT 10.070 5.920 10.390 6.240 ;
        RECT 11.680 5.920 12.000 6.240 ;
        RECT 8.500 5.680 8.730 5.910 ;
        RECT 10.110 5.690 10.340 5.920 ;
        RECT 11.720 5.690 11.950 5.920 ;
        RECT 12.970 5.650 13.290 5.970 ;
        RECT 13.640 5.650 13.960 5.970 ;
        RECT 3.750 5.430 4.070 5.470 ;
        RECT 3.520 5.200 4.070 5.430 ;
        RECT 3.750 5.150 4.070 5.200 ;
        RECT 8.340 5.080 8.570 5.370 ;
        RECT 0.300 4.560 0.620 4.880 ;
        RECT 8.350 4.860 8.570 5.080 ;
        RECT 0.340 4.330 0.570 4.560 ;
        RECT 9.930 4.210 10.150 4.430 ;
        RECT 0.320 3.610 0.640 3.930 ;
        RECT 9.920 3.920 10.150 4.210 ;
        RECT 0.360 3.380 0.590 3.610 ;
        RECT 6.740 3.550 10.190 3.720 ;
        RECT 0.320 2.670 0.640 2.990 ;
        RECT 0.360 2.440 0.590 2.670 ;
        RECT 8.290 1.140 8.470 2.560 ;
        RECT 9.990 1.710 10.190 3.550 ;
        RECT 8.290 1.020 8.640 1.140 ;
        RECT 8.380 0.820 8.640 1.020 ;
      LAYER via ;
        RECT 0.350 5.900 0.610 6.160 ;
        RECT 2.060 5.940 2.320 6.200 ;
        RECT 5.260 5.940 5.520 6.200 ;
        RECT 6.870 5.950 7.130 6.210 ;
        RECT 8.490 5.940 8.750 6.200 ;
        RECT 10.100 5.950 10.360 6.210 ;
        RECT 11.710 5.950 11.970 6.210 ;
        RECT 13.000 5.680 13.260 5.940 ;
        RECT 13.670 5.680 13.930 5.940 ;
        RECT 3.780 5.180 4.040 5.440 ;
        RECT 0.330 4.590 0.590 4.850 ;
        RECT 0.350 3.640 0.610 3.900 ;
        RECT 0.350 2.700 0.610 2.960 ;
        RECT 8.380 0.850 8.640 1.110 ;
      LAYER met2 ;
        RECT 0.320 3.610 0.640 3.930 ;
  END
END sky130_hilas_DAC5bit01

MACRO sky130_hilas_capacitorSize04
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize04 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.150 BY 7.320 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAP1TERM02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.400 3.900 5.750 4.180 ;
    END
  END CAP1TERM02
  PIN CAP2TERM02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.400 0.900 5.760 1.180 ;
    END
  END CAP2TERM02
  PIN CAP2TERM01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 0.900 0.280 1.180 ;
    END
  END CAP2TERM01
  PIN CAP1TERM01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 3.900 0.270 4.180 ;
    END
  END CAP1TERM01
  OBS
      LAYER met2 ;
        RECT 0.000 4.850 5.750 5.030 ;
        RECT 0.000 4.420 5.800 4.600 ;
        RECT 0.560 4.200 0.930 4.420 ;
        RECT 5.430 4.200 5.800 4.420 ;
        RECT 0.000 3.420 5.750 3.600 ;
        RECT 0.000 2.990 5.750 3.170 ;
        RECT 0.000 1.840 5.750 2.010 ;
        RECT 0.590 1.590 0.960 1.600 ;
        RECT 5.430 1.590 5.800 1.600 ;
        RECT 0.000 1.420 5.800 1.590 ;
        RECT 0.590 1.200 0.960 1.420 ;
        RECT 5.430 1.200 5.800 1.420 ;
        RECT 0.000 0.440 5.750 0.610 ;
        RECT 0.000 0.000 5.750 0.170 ;
      LAYER via2 ;
        RECT 0.610 4.260 0.890 4.540 ;
        RECT 5.480 4.260 5.760 4.540 ;
        RECT 0.640 1.260 0.920 1.540 ;
        RECT 5.480 1.260 5.760 1.540 ;
      LAYER met3 ;
        RECT 5.850 5.040 8.150 7.320 ;
        RECT 0.340 4.000 1.130 4.750 ;
        RECT 3.840 3.640 4.870 4.390 ;
        RECT 5.210 4.310 6.000 4.750 ;
        RECT 5.210 4.000 8.150 4.310 ;
        RECT 5.850 2.030 8.150 4.000 ;
        RECT 0.370 1.000 1.160 1.750 ;
        RECT 3.830 0.650 4.890 1.380 ;
        RECT 5.210 1.000 6.000 1.750 ;
      LAYER via3 ;
        RECT 0.530 4.150 0.960 4.630 ;
        RECT 5.400 4.150 5.830 4.630 ;
        RECT 0.560 1.150 0.990 1.630 ;
        RECT 5.400 1.150 5.830 1.630 ;
      LAYER met4 ;
        RECT 6.700 6.270 7.150 6.280 ;
        RECT 6.680 5.780 7.200 6.270 ;
        RECT 0.430 4.110 1.090 4.720 ;
        RECT 0.240 3.700 3.030 4.110 ;
        RECT 5.300 4.060 5.960 4.720 ;
        RECT 6.700 3.260 7.150 3.270 ;
        RECT 6.680 2.770 7.200 3.260 ;
        RECT 0.460 1.100 1.120 1.720 ;
        RECT 0.460 1.060 2.670 1.100 ;
        RECT 5.300 1.060 5.960 1.720 ;
        RECT 0.550 0.690 2.670 1.060 ;
  END
END sky130_hilas_capacitorSize04

MACRO sky130_hilas_capacitorArray01
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorArray01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.700 BY 14.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM2
    USE ANALOG ;
    PORT
      LAYER met3 ;
        RECT 35.230 2.200 36.380 3.840 ;
        RECT 35.680 2.190 36.380 2.200 ;
    END
  END CAPTERM2
  PIN CAPTERM1
    USE ANALOG ;
    ANTENNADIFFAREA 1.012300 ;
    PORT
      LAYER met3 ;
        RECT 11.250 5.740 11.630 6.030 ;
        RECT 11.170 4.490 11.710 5.740 ;
    END
  END CAPTERM1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 5.390 6.010 5.710 6.020 ;
        RECT 8.760 6.010 9.080 6.100 ;
        RECT 9.320 6.010 9.640 6.070 ;
        RECT 5.390 5.930 9.640 6.010 ;
        RECT 10.740 6.020 11.250 6.050 ;
        RECT 10.740 5.930 11.670 6.020 ;
        RECT 5.390 5.830 11.670 5.930 ;
        RECT 5.390 5.760 5.710 5.830 ;
        RECT 8.880 5.740 11.670 5.830 ;
        RECT 11.170 5.720 11.670 5.740 ;
      LAYER via2 ;
        RECT 11.300 5.720 11.580 6.000 ;
    END
  END VINJ
  PIN GATESELECT
    PORT
      LAYER met1 ;
        RECT 9.120 6.000 9.310 6.050 ;
    END
  END GATESELECT
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 0.360 5.910 0.760 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.360 0.000 0.750 0.120 ;
    END
  END VTUN
  PIN GATE
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 4.420 5.970 4.790 6.050 ;
        RECT 4.410 5.920 4.790 5.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.400 0.130 4.410 0.150 ;
        RECT 4.400 0.010 4.790 0.130 ;
        RECT 4.400 0.000 4.410 0.010 ;
    END
  END GATE
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 0.000 3.510 0.120 3.690 ;
    END
    PORT
      LAYER met2 ;
        RECT 35.690 3.690 36.700 3.700 ;
        RECT 8.940 3.510 36.700 3.690 ;
    END
  END DRAIN2
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 0.010 5.370 0.120 5.550 ;
    END
    PORT
      LAYER met2 ;
        RECT 8.980 5.400 36.700 5.550 ;
        RECT 2.640 5.370 36.700 5.400 ;
        RECT 2.640 5.220 10.260 5.370 ;
    END
  END DRAIN1
  PIN DRAIN4
    PORT
      LAYER met2 ;
        RECT 8.810 0.520 36.700 0.690 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.020 0.520 0.120 0.690 ;
    END
  END DRAIN4
  PIN DRAIN3
    PORT
      LAYER met4 ;
        RECT 10.070 2.300 10.730 2.680 ;
        RECT 13.710 2.300 16.900 2.330 ;
        RECT 19.350 2.300 19.650 2.330 ;
        RECT 10.070 2.020 22.570 2.300 ;
        RECT 10.370 2.000 22.570 2.020 ;
        RECT 13.710 1.630 14.010 2.000 ;
        RECT 16.600 1.660 16.900 2.000 ;
        RECT 19.350 1.660 19.650 2.000 ;
        RECT 16.600 1.630 19.650 1.660 ;
        RECT 22.270 1.630 22.570 2.000 ;
        RECT 13.710 1.330 22.570 1.630 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.020 2.360 0.120 2.530 ;
    END
  END DRAIN3
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2.990 6.050 3.390 10.730 ;
        RECT 2.800 5.990 3.390 6.050 ;
        RECT 2.990 4.230 3.390 5.990 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.730 5.980 6.970 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.800 0.000 3.040 0.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.730 0.000 6.970 0.070 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 17.150 14.670 18.880 14.720 ;
        RECT 2.640 9.390 2.710 9.570 ;
        RECT 13.040 9.230 15.600 11.140 ;
        RECT 3.210 9.040 3.800 9.150 ;
        RECT 6.950 8.980 8.060 9.210 ;
        RECT 11.590 7.550 11.940 7.560 ;
        RECT 11.590 7.390 11.760 7.550 ;
        RECT 11.930 7.390 11.940 7.550 ;
        RECT 13.040 6.050 15.600 8.960 ;
        RECT 15.960 8.230 18.880 14.670 ;
        RECT 21.150 11.140 22.880 12.980 ;
        RECT 15.960 8.180 18.190 8.230 ;
        RECT 10.070 6.040 35.420 6.050 ;
        RECT 3.210 5.760 3.800 5.950 ;
        RECT 6.950 5.740 8.060 6.010 ;
        RECT 10.080 5.970 35.420 6.040 ;
        RECT 0.010 5.370 0.120 5.550 ;
        RECT 0.000 3.510 0.120 3.690 ;
        RECT 0.020 0.520 0.120 0.690 ;
        RECT 10.060 0.060 35.420 5.970 ;
        RECT 10.070 0.010 35.420 0.060 ;
        RECT 12.000 0.000 35.420 0.010 ;
      LAYER li1 ;
        RECT 17.540 11.660 18.090 12.090 ;
        RECT 21.570 11.590 22.120 12.020 ;
        RECT 13.280 10.790 13.600 10.830 ;
        RECT 13.280 10.670 13.610 10.790 ;
        RECT 13.280 10.570 13.720 10.670 ;
        RECT 13.380 10.500 13.720 10.570 ;
        RECT 15.000 10.400 15.200 10.750 ;
        RECT 13.280 10.240 13.600 10.280 ;
        RECT 13.280 10.050 13.610 10.240 ;
        RECT 13.280 10.020 13.720 10.050 ;
        RECT 13.380 9.880 13.720 10.020 ;
        RECT 14.270 9.780 14.470 10.380 ;
        RECT 15.000 10.370 15.210 10.400 ;
        RECT 14.990 9.780 15.210 10.370 ;
        RECT 5.460 8.750 5.630 9.280 ;
        RECT 9.400 8.740 9.570 9.270 ;
        RECT 13.380 8.170 13.720 8.310 ;
        RECT 13.280 8.140 13.720 8.170 ;
        RECT 5.470 7.040 5.640 8.050 ;
        RECT 13.280 7.950 13.610 8.140 ;
        RECT 13.280 7.910 13.600 7.950 ;
        RECT 9.400 6.900 9.570 7.910 ;
        RECT 14.270 7.810 14.470 8.410 ;
        RECT 14.990 7.820 15.210 8.410 ;
        RECT 15.000 7.790 15.210 7.820 ;
        RECT 13.380 7.620 13.720 7.690 ;
        RECT 11.500 7.390 11.940 7.560 ;
        RECT 13.280 7.520 13.720 7.620 ;
        RECT 13.280 7.430 13.610 7.520 ;
        RECT 13.280 7.330 13.720 7.430 ;
        RECT 13.380 7.260 13.720 7.330 ;
        RECT 15.000 7.160 15.200 7.790 ;
        RECT 13.280 7.000 13.600 7.040 ;
        RECT 13.280 6.810 13.610 7.000 ;
        RECT 13.280 6.780 13.720 6.810 ;
        RECT 13.380 6.640 13.720 6.780 ;
        RECT 14.270 6.540 14.470 7.140 ;
        RECT 15.000 7.130 15.210 7.160 ;
        RECT 14.990 6.540 15.210 7.130 ;
        RECT 13.380 4.940 13.720 5.080 ;
        RECT 13.280 4.910 13.720 4.940 ;
        RECT 13.280 4.720 13.610 4.910 ;
        RECT 13.280 4.680 13.600 4.720 ;
        RECT 14.270 4.580 14.470 5.180 ;
        RECT 14.990 4.590 15.210 5.180 ;
        RECT 15.000 4.560 15.210 4.590 ;
        RECT 13.380 4.390 13.720 4.460 ;
        RECT 13.280 4.290 13.720 4.390 ;
        RECT 13.280 4.170 13.610 4.290 ;
        RECT 15.000 4.210 15.200 4.560 ;
        RECT 13.280 4.130 13.600 4.170 ;
      LAYER mcon ;
        RECT 17.540 11.740 17.810 12.010 ;
        RECT 21.570 11.670 21.840 11.940 ;
        RECT 13.340 10.610 13.510 10.780 ;
        RECT 13.340 10.060 13.510 10.230 ;
        RECT 14.280 10.170 14.450 10.340 ;
        RECT 15.010 10.200 15.180 10.370 ;
        RECT 5.460 9.110 5.630 9.280 ;
        RECT 9.400 9.100 9.570 9.270 ;
        RECT 13.340 7.960 13.510 8.130 ;
        RECT 5.470 7.650 5.640 7.820 ;
        RECT 5.470 7.290 5.640 7.460 ;
        RECT 14.280 7.850 14.450 8.020 ;
        RECT 15.010 7.820 15.180 7.990 ;
        RECT 9.400 7.510 9.570 7.680 ;
        RECT 11.760 7.390 11.940 7.560 ;
        RECT 13.340 7.370 13.510 7.580 ;
        RECT 9.400 7.150 9.570 7.320 ;
        RECT 13.340 6.820 13.510 6.990 ;
        RECT 14.280 6.930 14.450 7.100 ;
        RECT 15.010 6.960 15.180 7.130 ;
        RECT 13.340 4.730 13.510 4.900 ;
        RECT 14.280 4.620 14.450 4.790 ;
        RECT 15.010 4.590 15.180 4.760 ;
        RECT 13.340 4.180 13.510 4.350 ;
      LAYER met1 ;
        RECT 5.430 9.320 5.670 10.730 ;
        RECT 7.040 10.400 7.420 10.730 ;
        RECT 9.360 9.340 9.600 10.730 ;
        RECT 13.270 10.540 13.590 10.860 ;
        RECT 11.380 10.460 11.540 10.500 ;
        RECT 11.750 10.450 11.940 10.500 ;
        RECT 12.190 10.450 12.350 10.500 ;
        RECT 14.270 10.400 14.430 11.130 ;
        RECT 14.270 10.380 14.470 10.400 ;
        RECT 13.270 9.990 13.590 10.310 ;
        RECT 14.250 10.140 14.480 10.380 ;
        RECT 14.270 10.090 14.480 10.140 ;
        RECT 14.640 10.090 14.830 11.080 ;
        RECT 15.080 10.430 15.240 11.130 ;
        RECT 5.420 8.660 5.680 9.320 ;
        RECT 9.340 8.680 9.610 9.340 ;
        RECT 14.270 9.230 14.430 10.090 ;
        RECT 14.660 9.970 14.830 10.090 ;
        RECT 14.670 9.230 14.830 9.970 ;
        RECT 14.970 9.880 15.240 10.430 ;
        RECT 14.970 9.830 15.250 9.880 ;
        RECT 15.080 9.740 15.250 9.830 ;
        RECT 15.080 9.230 15.240 9.740 ;
        RECT 5.430 6.050 5.670 8.660 ;
        RECT 5.420 5.730 5.680 6.050 ;
        RECT 8.790 5.810 9.050 6.130 ;
        RECT 9.360 6.090 9.600 8.680 ;
        RECT 13.270 7.880 13.590 8.200 ;
        RECT 14.270 8.100 14.430 8.960 ;
        RECT 14.670 8.220 14.830 8.960 ;
        RECT 15.080 8.450 15.240 8.960 ;
        RECT 15.080 8.360 15.250 8.450 ;
        RECT 14.660 8.100 14.830 8.220 ;
        RECT 14.270 8.050 14.480 8.100 ;
        RECT 14.250 7.810 14.480 8.050 ;
        RECT 14.270 7.790 14.470 7.810 ;
        RECT 11.810 7.590 11.940 7.610 ;
        RECT 11.730 7.570 11.970 7.590 ;
        RECT 11.530 7.380 11.970 7.570 ;
        RECT 11.730 7.360 11.970 7.380 ;
        RECT 11.830 7.320 11.940 7.360 ;
        RECT 13.270 7.300 13.590 7.650 ;
        RECT 14.270 7.160 14.430 7.790 ;
        RECT 14.270 7.140 14.470 7.160 ;
        RECT 13.270 6.750 13.590 7.070 ;
        RECT 14.250 6.900 14.480 7.140 ;
        RECT 14.270 6.850 14.480 6.900 ;
        RECT 14.640 6.850 14.830 8.100 ;
        RECT 14.970 8.310 15.250 8.360 ;
        RECT 14.970 7.760 15.240 8.310 ;
        RECT 16.610 8.180 16.990 14.680 ;
        RECT 17.480 11.200 17.870 13.060 ;
        RECT 21.510 11.130 21.900 12.990 ;
        RECT 15.080 7.190 15.240 7.760 ;
        RECT 9.350 6.050 9.610 6.090 ;
        RECT 9.350 6.000 9.720 6.050 ;
        RECT 9.350 5.770 9.610 6.000 ;
        RECT 14.270 5.990 14.430 6.850 ;
        RECT 14.660 6.730 14.830 6.850 ;
        RECT 14.670 5.990 14.830 6.730 ;
        RECT 14.970 6.640 15.240 7.190 ;
        RECT 14.970 6.590 15.250 6.640 ;
        RECT 15.080 6.500 15.250 6.590 ;
        RECT 15.080 5.990 15.240 6.500 ;
        RECT 5.430 4.230 5.670 5.730 ;
        RECT 7.040 4.230 7.420 4.830 ;
        RECT 9.360 4.230 9.600 5.770 ;
        RECT 13.270 4.650 13.590 4.970 ;
        RECT 14.270 4.870 14.430 5.730 ;
        RECT 14.670 4.990 14.830 5.730 ;
        RECT 15.080 5.220 15.240 5.730 ;
        RECT 15.080 5.130 15.250 5.220 ;
        RECT 14.660 4.870 14.830 4.990 ;
        RECT 14.270 4.820 14.480 4.870 ;
        RECT 14.250 4.580 14.480 4.820 ;
        RECT 14.270 4.560 14.470 4.580 ;
        RECT 13.270 4.100 13.590 4.420 ;
        RECT 14.270 3.830 14.430 4.560 ;
        RECT 14.640 3.880 14.830 4.870 ;
        RECT 14.970 5.080 15.250 5.130 ;
        RECT 14.970 4.530 15.240 5.080 ;
        RECT 15.080 3.830 15.240 4.530 ;
        RECT 8.750 0.010 8.910 0.070 ;
        RECT 9.120 0.010 9.310 0.070 ;
        RECT 9.560 0.010 9.720 0.070 ;
      LAYER via ;
        RECT 13.300 10.570 13.560 10.830 ;
        RECT 13.300 10.020 13.560 10.280 ;
        RECT 5.420 5.760 5.680 6.020 ;
        RECT 8.790 5.840 9.050 6.100 ;
        RECT 13.300 7.910 13.560 8.170 ;
        RECT 13.300 7.330 13.560 7.620 ;
        RECT 13.300 6.780 13.560 7.040 ;
        RECT 9.350 5.800 9.610 6.060 ;
        RECT 13.300 4.680 13.560 4.940 ;
        RECT 13.300 4.130 13.560 4.390 ;
      LAYER met2 ;
        RECT 13.270 10.580 13.580 10.870 ;
        RECT 13.270 10.540 15.600 10.580 ;
        RECT 13.420 10.400 15.600 10.540 ;
        RECT 2.640 9.990 10.270 10.170 ;
        RECT 13.270 10.150 13.580 10.320 ;
        RECT 13.040 9.970 13.130 10.150 ;
        RECT 13.270 9.990 15.600 10.150 ;
        RECT 13.430 9.970 15.600 9.990 ;
        RECT 2.640 9.550 10.270 9.730 ;
        RECT 2.640 8.450 10.270 8.630 ;
        RECT 2.640 8.020 10.270 8.200 ;
        RECT 13.040 8.040 13.130 8.220 ;
        RECT 13.430 8.200 15.600 8.220 ;
        RECT 13.270 8.040 15.600 8.200 ;
        RECT 13.270 7.870 13.580 8.040 ;
        RECT 13.420 7.650 15.600 7.790 ;
        RECT 13.270 7.610 15.600 7.650 ;
        RECT 13.270 7.340 13.580 7.610 ;
        RECT 13.270 7.300 15.600 7.340 ;
        RECT 13.420 7.160 15.600 7.300 ;
        RECT 2.640 6.750 10.260 6.930 ;
        RECT 13.270 6.910 13.580 7.080 ;
        RECT 13.040 6.730 13.130 6.910 ;
        RECT 13.270 6.750 15.600 6.910 ;
        RECT 13.430 6.730 15.600 6.750 ;
        RECT 2.640 6.320 10.270 6.500 ;
        RECT 8.920 4.970 36.700 5.120 ;
        RECT 2.640 4.940 36.700 4.970 ;
        RECT 2.640 4.800 10.240 4.940 ;
        RECT 13.040 4.810 13.130 4.940 ;
        RECT 13.270 4.810 15.600 4.940 ;
        RECT 10.240 4.250 10.610 4.650 ;
        RECT 13.270 4.640 13.580 4.810 ;
        RECT 13.420 4.420 15.600 4.560 ;
        RECT 13.270 4.380 15.600 4.420 ;
        RECT 13.270 4.120 13.580 4.380 ;
        RECT 8.980 3.940 36.700 4.120 ;
        RECT 36.010 2.790 36.700 3.200 ;
        RECT 10.200 2.530 10.570 2.560 ;
        RECT 8.770 2.360 36.700 2.530 ;
        RECT 10.200 2.160 10.570 2.360 ;
        RECT 8.870 1.940 36.700 2.110 ;
        RECT 11.290 1.290 11.660 1.690 ;
        RECT 8.850 0.960 36.700 1.130 ;
      LAYER via2 ;
        RECT 10.290 4.310 10.570 4.590 ;
        RECT 36.080 2.850 36.370 3.130 ;
        RECT 10.250 2.220 10.530 2.500 ;
        RECT 11.340 1.350 11.620 1.630 ;
      LAYER met3 ;
        RECT 10.020 4.050 10.810 4.800 ;
        RECT 9.980 1.960 10.770 2.710 ;
        RECT 11.070 1.090 11.860 1.840 ;
        RECT 11.460 0.790 11.640 1.090 ;
      LAYER via3 ;
        RECT 10.210 4.200 10.640 4.680 ;
        RECT 10.170 2.110 10.600 2.590 ;
        RECT 11.260 1.240 11.690 1.720 ;
      LAYER met4 ;
        RECT 12.790 5.380 16.890 5.680 ;
        RECT 11.100 4.770 13.800 4.880 ;
        RECT 10.110 4.110 10.770 4.770 ;
        RECT 11.100 4.470 14.010 4.770 ;
        RECT 13.500 4.130 14.010 4.470 ;
        RECT 16.510 4.180 16.890 5.380 ;
        RECT 19.350 4.210 22.630 4.510 ;
        RECT 10.410 3.750 11.770 4.050 ;
        RECT 11.470 3.190 11.770 3.750 ;
        RECT 19.350 3.190 19.650 4.210 ;
        RECT 22.330 3.190 22.630 4.210 ;
        RECT 11.470 2.890 22.630 3.190 ;
        RECT 25.030 4.190 33.920 4.490 ;
        RECT 11.160 1.150 11.820 1.810 ;
        RECT 25.030 1.670 25.330 4.190 ;
        RECT 27.860 4.160 30.970 4.190 ;
        RECT 27.860 1.670 28.160 4.160 ;
        RECT 30.670 1.670 30.970 4.160 ;
        RECT 33.620 1.670 33.920 4.190 ;
        RECT 25.030 1.370 33.980 1.670 ;
        RECT 30.670 1.360 33.980 1.370 ;
        RECT 11.340 0.790 11.850 1.090 ;
        RECT 11.550 0.550 11.850 0.790 ;
        RECT 33.680 0.550 33.980 1.360 ;
        RECT 11.550 0.250 33.980 0.550 ;
  END
END sky130_hilas_capacitorArray01

MACRO sky130_hilas_pFETmed
  CLASS CORE ;
  FOREIGN sky130_hilas_pFETmed ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.190 BY 2.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 0.000 0.000 1.190 2.870 ;
      LAYER li1 ;
        RECT 0.240 0.150 0.410 2.640 ;
        RECT 0.790 0.140 0.960 2.640 ;
  END
END sky130_hilas_pFETmed

MACRO sky130_hilas_swc4x1cellOverlap2
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x1cellOverlap2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.240 BY 7.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 8.000 6.980 12.000 7.050 ;
        RECT 8.000 5.070 12.240 6.980 ;
        RECT 8.000 4.910 12.000 5.070 ;
        RECT 8.000 2.060 12.240 4.910 ;
        RECT 8.000 1.910 12.000 2.060 ;
        RECT 8.000 1.000 12.240 1.910 ;
        RECT 9.680 0.000 12.240 1.000 ;
      LAYER li1 ;
        RECT 1.680 5.730 1.850 6.620 ;
        RECT 8.350 6.590 11.660 6.720 ;
        RECT 8.350 6.240 11.840 6.590 ;
        RECT 8.350 5.740 11.850 6.240 ;
        RECT 10.020 5.720 10.360 5.740 ;
        RECT 10.910 5.620 11.110 5.740 ;
        RECT 11.630 5.620 11.850 5.740 ;
        RECT 1.680 4.210 1.850 5.100 ;
        RECT 8.350 4.360 11.660 5.250 ;
        RECT 8.350 4.270 11.850 4.360 ;
        RECT 10.020 4.120 10.360 4.260 ;
        RECT 9.920 4.090 10.360 4.120 ;
        RECT 9.920 3.900 10.250 4.090 ;
        RECT 9.920 3.860 10.240 3.900 ;
        RECT 10.910 3.780 11.110 4.270 ;
        RECT 11.630 3.780 11.850 4.270 ;
        RECT 8.350 3.740 11.850 3.780 ;
        RECT 1.680 2.760 1.850 3.650 ;
        RECT 8.350 3.570 11.840 3.740 ;
        RECT 8.140 3.400 11.840 3.570 ;
        RECT 8.350 3.230 11.840 3.400 ;
        RECT 8.350 2.800 11.850 3.230 ;
        RECT 10.020 2.710 10.360 2.800 ;
        RECT 10.910 2.610 11.110 2.800 ;
        RECT 11.630 2.610 11.850 2.800 ;
        RECT 1.680 1.220 1.850 2.110 ;
        RECT 8.350 1.360 11.660 2.310 ;
        RECT 8.350 1.330 11.850 1.360 ;
        RECT 10.020 1.120 10.360 1.260 ;
        RECT 9.920 1.090 10.360 1.120 ;
        RECT 9.920 0.900 10.250 1.090 ;
        RECT 9.920 0.860 10.240 0.900 ;
        RECT 10.910 0.760 11.110 1.330 ;
        RECT 11.630 0.770 11.850 1.330 ;
        RECT 11.640 0.740 11.850 0.770 ;
        RECT 10.020 0.570 10.360 0.640 ;
        RECT 9.920 0.470 10.360 0.570 ;
        RECT 9.920 0.350 10.250 0.470 ;
        RECT 11.640 0.390 11.840 0.740 ;
        RECT 9.920 0.310 10.240 0.350 ;
      LAYER mcon ;
        RECT 1.680 6.420 1.850 6.590 ;
        RECT 9.920 6.620 10.090 6.660 ;
        RECT 9.920 6.490 10.150 6.620 ;
        RECT 9.980 6.450 10.150 6.490 ;
        RECT 9.980 5.970 10.150 6.070 ;
        RECT 10.920 6.010 11.090 6.180 ;
        RECT 11.650 6.040 11.820 6.210 ;
        RECT 9.920 5.900 10.150 5.970 ;
        RECT 9.920 5.800 10.090 5.900 ;
        RECT 1.680 4.900 1.850 5.070 ;
        RECT 9.920 5.020 10.090 5.190 ;
        RECT 9.920 4.330 10.090 4.500 ;
        RECT 9.980 3.910 10.150 4.080 ;
        RECT 10.920 3.800 11.090 3.970 ;
        RECT 11.650 3.770 11.820 3.940 ;
        RECT 1.680 3.450 1.850 3.620 ;
        RECT 9.920 3.610 10.090 3.720 ;
        RECT 8.400 3.400 8.580 3.570 ;
        RECT 9.920 3.550 10.150 3.610 ;
        RECT 9.980 3.360 10.150 3.550 ;
        RECT 9.980 3.030 10.150 3.060 ;
        RECT 9.920 2.890 10.150 3.030 ;
        RECT 10.920 3.000 11.090 3.170 ;
        RECT 11.650 3.030 11.820 3.200 ;
        RECT 9.920 2.860 10.090 2.890 ;
        RECT 1.680 1.910 1.850 2.080 ;
        RECT 9.920 2.080 10.090 2.250 ;
        RECT 9.920 1.390 10.090 1.560 ;
        RECT 9.980 0.910 10.150 1.080 ;
        RECT 10.920 0.800 11.090 0.970 ;
        RECT 11.650 0.770 11.820 0.940 ;
        RECT 9.980 0.360 10.150 0.530 ;
      LAYER met1 ;
        RECT 1.010 0.460 1.280 6.510 ;
        RECT 1.650 5.520 1.880 6.810 ;
        RECT 9.880 6.700 10.120 6.720 ;
        RECT 9.880 6.380 10.230 6.700 ;
        RECT 9.880 6.150 10.120 6.380 ;
        RECT 10.910 6.240 11.070 6.970 ;
        RECT 10.910 6.220 11.110 6.240 ;
        RECT 9.880 6.080 10.230 6.150 ;
        RECT 9.890 5.830 10.230 6.080 ;
        RECT 10.890 5.980 11.120 6.220 ;
        RECT 10.910 5.930 11.120 5.980 ;
        RECT 11.280 5.930 11.470 6.920 ;
        RECT 11.720 6.270 11.880 6.970 ;
        RECT 9.890 5.820 10.120 5.830 ;
        RECT 9.890 5.600 10.130 5.820 ;
        RECT 1.650 4.000 1.880 5.290 ;
        RECT 9.880 4.610 10.120 5.250 ;
        RECT 10.910 5.070 11.070 5.930 ;
        RECT 11.300 5.810 11.470 5.930 ;
        RECT 11.310 5.070 11.470 5.810 ;
        RECT 11.610 5.720 11.880 6.270 ;
        RECT 11.610 5.670 11.890 5.720 ;
        RECT 11.720 5.580 11.890 5.670 ;
        RECT 11.720 5.070 11.880 5.580 ;
        RECT 9.890 4.350 10.120 4.610 ;
        RECT 9.890 4.150 10.130 4.350 ;
        RECT 9.890 4.130 10.230 4.150 ;
        RECT 1.650 2.550 1.880 3.840 ;
        RECT 9.910 3.830 10.230 4.130 ;
        RECT 10.910 4.050 11.070 4.910 ;
        RECT 11.310 4.170 11.470 4.910 ;
        RECT 11.720 4.400 11.880 4.910 ;
        RECT 11.720 4.310 11.890 4.400 ;
        RECT 11.300 4.050 11.470 4.170 ;
        RECT 10.910 4.000 11.120 4.050 ;
        RECT 9.880 3.690 10.120 3.780 ;
        RECT 10.890 3.760 11.120 4.000 ;
        RECT 10.910 3.740 11.110 3.760 ;
        RECT 8.450 3.600 8.580 3.620 ;
        RECT 8.370 3.370 8.610 3.600 ;
        RECT 8.470 3.330 8.580 3.370 ;
        RECT 9.880 3.280 10.230 3.690 ;
        RECT 9.880 3.140 10.120 3.280 ;
        RECT 10.910 3.230 11.070 3.740 ;
        RECT 10.910 3.210 11.110 3.230 ;
        RECT 9.890 2.820 10.230 3.140 ;
        RECT 10.890 2.970 11.120 3.210 ;
        RECT 10.910 2.920 11.120 2.970 ;
        RECT 11.280 2.920 11.470 4.050 ;
        RECT 11.610 4.260 11.890 4.310 ;
        RECT 11.610 3.710 11.880 4.260 ;
        RECT 11.720 3.260 11.880 3.710 ;
        RECT 9.890 2.660 10.130 2.820 ;
        RECT 1.650 1.010 1.880 2.300 ;
        RECT 9.880 1.670 10.120 2.310 ;
        RECT 10.910 2.060 11.070 2.920 ;
        RECT 11.300 2.800 11.470 2.920 ;
        RECT 11.310 2.060 11.470 2.800 ;
        RECT 11.610 2.710 11.880 3.260 ;
        RECT 11.610 2.660 11.890 2.710 ;
        RECT 11.720 2.570 11.890 2.660 ;
        RECT 11.720 2.060 11.880 2.570 ;
        RECT 9.890 1.410 10.120 1.670 ;
        RECT 9.890 1.190 10.130 1.410 ;
        RECT 9.910 0.830 10.230 1.150 ;
        RECT 10.910 1.050 11.070 1.910 ;
        RECT 11.310 1.170 11.470 1.910 ;
        RECT 11.720 1.400 11.880 1.910 ;
        RECT 11.720 1.310 11.890 1.400 ;
        RECT 11.300 1.050 11.470 1.170 ;
        RECT 10.910 1.000 11.120 1.050 ;
        RECT 10.890 0.760 11.120 1.000 ;
        RECT 10.910 0.740 11.110 0.760 ;
        RECT 9.910 0.280 10.230 0.600 ;
        RECT 10.910 0.010 11.070 0.740 ;
        RECT 11.280 0.060 11.470 1.050 ;
        RECT 11.610 1.260 11.890 1.310 ;
        RECT 11.610 0.710 11.880 1.260 ;
        RECT 11.720 0.010 11.880 0.710 ;
      LAYER via ;
        RECT 9.940 6.410 10.200 6.670 ;
        RECT 9.940 5.860 10.200 6.120 ;
        RECT 9.940 3.860 10.200 4.120 ;
        RECT 9.940 3.310 10.200 3.660 ;
        RECT 9.940 2.850 10.200 3.110 ;
        RECT 9.940 0.860 10.200 1.120 ;
        RECT 9.940 0.310 10.200 0.570 ;
      LAYER met2 ;
        RECT 9.910 6.420 10.220 6.710 ;
        RECT 9.910 6.380 12.240 6.420 ;
        RECT 10.060 6.240 12.240 6.380 ;
        RECT 0.000 5.940 6.880 6.010 ;
        RECT 9.910 5.990 10.220 6.160 ;
        RECT 0.000 5.830 6.910 5.940 ;
        RECT 9.680 5.810 9.770 5.990 ;
        RECT 9.910 5.830 12.240 5.990 ;
        RECT 10.070 5.810 12.240 5.830 ;
        RECT 0.000 5.400 9.010 5.580 ;
        RECT 0.000 4.520 6.880 4.580 ;
        RECT 0.000 4.400 6.910 4.520 ;
        RECT 0.000 4.080 6.870 4.150 ;
        RECT 0.000 3.970 6.910 4.080 ;
        RECT 9.680 3.990 9.770 4.170 ;
        RECT 10.070 4.150 12.240 4.170 ;
        RECT 9.910 3.990 12.240 4.150 ;
        RECT 9.910 3.820 10.220 3.990 ;
        RECT 10.060 3.700 12.240 3.740 ;
        RECT 9.910 3.560 12.240 3.700 ;
        RECT 9.910 3.410 10.220 3.560 ;
        RECT 9.910 3.270 12.240 3.410 ;
        RECT 10.060 3.230 12.240 3.270 ;
        RECT 0.000 2.820 6.910 2.990 ;
        RECT 9.910 2.980 10.220 3.150 ;
        RECT 9.680 2.800 9.770 2.980 ;
        RECT 9.910 2.820 12.240 2.980 ;
        RECT 10.070 2.800 12.240 2.820 ;
        RECT 0.000 2.400 6.910 2.570 ;
        RECT 0.000 1.420 6.910 1.590 ;
        RECT 0.000 0.980 6.910 1.150 ;
        RECT 9.680 0.990 9.770 1.170 ;
        RECT 10.070 1.150 12.240 1.170 ;
        RECT 9.910 0.990 12.240 1.150 ;
        RECT 9.910 0.820 10.220 0.990 ;
        RECT 10.060 0.600 12.240 0.740 ;
        RECT 9.910 0.560 12.240 0.600 ;
        RECT 9.910 0.270 10.220 0.560 ;
  END
END sky130_hilas_swc4x1cellOverlap2

MACRO sky130_hilas_TA2SignalBiasCell
  CLASS CORE ;
  FOREIGN sky130_hilas_TA2SignalBiasCell ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.810 BY 24.010 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VOUT_AMP2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 9.630 12.320 9.780 12.540 ;
    END
  END VOUT_AMP2
  PIN VOUT_AMP1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 9.630 11.500 9.780 11.720 ;
    END
  END VOUT_AMP1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 7.820 8.980 8.160 9.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 7.820 14.890 8.160 15.030 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 8.490 8.980 8.760 9.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.490 14.880 8.760 15.030 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.900 15.020 2.810 15.030 ;
        RECT 0.900 9.420 6.500 15.020 ;
        RECT 10.480 9.470 11.760 12.310 ;
        RECT 0.900 9.240 1.330 9.420 ;
        RECT 0.900 9.010 1.610 9.240 ;
        RECT 0.900 8.990 1.330 9.010 ;
      LAYER met2 ;
        RECT 8.960 15.800 9.270 16.090 ;
        RECT 10.620 15.800 10.930 16.050 ;
        RECT 8.240 15.720 10.930 15.800 ;
        RECT 8.240 15.570 10.780 15.720 ;
        RECT 8.910 15.110 9.220 15.440 ;
        RECT 1.690 15.000 1.930 15.030 ;
        RECT 1.690 14.670 2.100 15.000 ;
        RECT 1.690 14.650 1.930 14.670 ;
        RECT 1.220 14.560 1.930 14.650 ;
        RECT 1.170 14.210 1.930 14.560 ;
        RECT 2.970 14.400 3.520 14.650 ;
        RECT 3.010 14.210 3.320 14.400 ;
        RECT 1.170 13.980 5.710 14.210 ;
        RECT 1.170 13.790 1.930 13.980 ;
        RECT 0.680 13.740 1.930 13.790 ;
        RECT 0.680 13.730 1.620 13.740 ;
        RECT 0.680 13.540 1.560 13.730 ;
        RECT 5.480 13.620 5.710 13.980 ;
        RECT 8.910 13.830 9.220 14.160 ;
        RECT 8.500 13.660 8.830 13.770 ;
        RECT 10.670 13.660 10.980 13.830 ;
        RECT 8.500 13.620 11.150 13.660 ;
        RECT 1.110 13.380 1.420 13.540 ;
        RECT 5.480 13.430 11.150 13.620 ;
        RECT 5.480 13.420 8.830 13.430 ;
        RECT 5.740 13.410 8.830 13.420 ;
        RECT 8.500 12.840 8.830 13.410 ;
        RECT 8.960 13.180 9.270 13.430 ;
        RECT 8.960 12.830 9.270 13.090 ;
        RECT 10.660 12.830 10.970 13.110 ;
        RECT 8.240 12.610 11.150 12.830 ;
        RECT 8.910 12.110 9.220 12.440 ;
        RECT 8.910 10.830 9.220 11.160 ;
        RECT 10.580 10.670 10.890 10.860 ;
        RECT 8.230 10.440 10.940 10.670 ;
        RECT 8.960 10.180 9.270 10.440 ;
    END
  END VPWR
  PIN VIN22
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.290 14.760 5.540 15.020 ;
    END
  END VIN22
  PIN VIN21
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.330 12.090 5.580 12.320 ;
    END
  END VIN21
  PIN VIN11
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 3.770 11.680 4.050 11.920 ;
    END
  END VIN11
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 3.730 9.000 3.990 9.250 ;
    END
  END VIN12
  PIN VBIAS2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.950 9.010 2.600 9.240 ;
    END
  END VBIAS2
  PIN VBIAS1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.910 11.680 2.370 11.920 ;
        RECT 0.910 11.670 1.550 11.680 ;
    END
  END VBIAS1
  OBS
      LAYER nwell ;
        RECT 3.630 21.020 7.240 24.010 ;
        RECT 3.630 17.970 7.240 20.960 ;
        RECT 0.000 16.520 3.610 16.590 ;
        RECT 1.340 16.230 1.790 16.460 ;
        RECT 3.090 16.230 3.540 16.460 ;
        RECT 8.500 14.850 9.780 15.030 ;
        RECT 10.480 13.930 11.760 16.770 ;
        RECT 8.500 8.980 9.780 9.170 ;
        RECT 4.650 7.550 5.100 7.780 ;
        RECT 3.310 7.420 5.170 7.490 ;
        RECT 6.940 3.050 8.800 6.040 ;
        RECT 6.940 0.000 8.800 2.990 ;
      LAYER li1 ;
        RECT 4.040 21.490 4.220 23.540 ;
        RECT 4.850 21.750 5.020 23.530 ;
        RECT 4.770 21.580 5.100 21.750 ;
        RECT 5.790 21.490 5.970 23.540 ;
        RECT 6.600 21.750 6.770 23.530 ;
        RECT 6.520 21.580 6.850 21.750 ;
        RECT 4.040 18.440 4.220 20.490 ;
        RECT 4.850 18.700 5.020 20.480 ;
        RECT 4.770 18.530 5.100 18.700 ;
        RECT 5.790 18.440 5.970 20.490 ;
        RECT 6.600 18.700 6.770 20.480 ;
        RECT 6.520 18.530 6.850 18.700 ;
        RECT 1.600 17.310 1.790 17.330 ;
        RECT 3.350 17.310 3.540 17.330 ;
        RECT 1.460 17.220 1.790 17.310 ;
        RECT 1.460 17.140 1.540 17.220 ;
        RECT 1.600 17.100 1.790 17.220 ;
        RECT 3.210 17.220 3.540 17.310 ;
        RECT 3.210 17.140 3.290 17.220 ;
        RECT 3.350 17.100 3.540 17.220 ;
        RECT 0.410 16.000 0.590 17.060 ;
        RECT 1.060 16.690 1.230 17.020 ;
        RECT 1.140 16.620 1.190 16.690 ;
        RECT 1.140 16.590 1.480 16.620 ;
        RECT 1.020 16.580 1.480 16.590 ;
        RECT 1.020 16.460 1.490 16.580 ;
        RECT 1.160 16.390 1.490 16.460 ;
        RECT 1.160 16.360 1.480 16.390 ;
        RECT 2.160 16.000 2.340 17.060 ;
        RECT 2.810 16.690 2.980 17.020 ;
        RECT 2.890 16.620 2.940 16.690 ;
        RECT 2.890 16.590 3.230 16.620 ;
        RECT 2.770 16.580 3.230 16.590 ;
        RECT 2.770 16.460 3.240 16.580 ;
        RECT 2.910 16.390 3.240 16.460 ;
        RECT 11.040 16.540 11.370 16.710 ;
        RECT 11.480 16.630 11.810 16.800 ;
        RECT 2.910 16.360 3.230 16.390 ;
        RECT 11.040 16.260 11.400 16.540 ;
        RECT 8.970 16.010 9.290 16.050 ;
        RECT 8.970 15.820 9.300 16.010 ;
        RECT 8.970 15.790 9.290 15.820 ;
        RECT 9.370 15.800 9.570 16.130 ;
        RECT 9.960 15.940 10.160 16.130 ;
        RECT 10.690 16.090 11.400 16.260 ;
        RECT 10.630 15.970 10.950 16.010 ;
        RECT 9.650 15.610 9.840 15.620 ;
        RECT 9.850 15.610 10.200 15.940 ;
        RECT 10.630 15.780 10.960 15.970 ;
        RECT 10.630 15.750 10.950 15.780 ;
        RECT 0.430 15.300 0.750 15.340 ;
        RECT 2.180 15.300 2.500 15.340 ;
        RECT 0.430 15.110 0.760 15.300 ;
        RECT 2.180 15.110 2.510 15.300 ;
        RECT 0.430 15.080 0.750 15.110 ;
        RECT 2.180 15.080 2.500 15.110 ;
        RECT 8.740 15.100 8.910 15.430 ;
        RECT 8.920 15.360 9.240 15.400 ;
        RECT 8.920 15.170 9.250 15.360 ;
        RECT 8.920 15.140 9.240 15.170 ;
        RECT 9.370 15.140 9.570 15.470 ;
        RECT 9.650 15.280 10.200 15.610 ;
        RECT 1.800 14.920 2.120 14.960 ;
        RECT 9.850 14.950 10.200 15.280 ;
        RECT 1.800 14.730 2.130 14.920 ;
        RECT 10.690 14.770 11.390 15.650 ;
        RECT 1.800 14.700 2.120 14.730 ;
        RECT 1.570 14.550 1.910 14.560 ;
        RECT 1.320 14.510 1.910 14.550 ;
        RECT 1.240 14.480 1.910 14.510 ;
        RECT 2.990 14.480 3.310 14.510 ;
        RECT 1.230 14.360 1.910 14.480 ;
        RECT 1.150 14.140 1.910 14.360 ;
        RECT 2.980 14.290 3.310 14.480 ;
        RECT 10.030 14.380 10.220 14.610 ;
        RECT 2.990 14.250 3.310 14.290 ;
        RECT 1.150 13.990 1.740 14.140 ;
        RECT 1.080 13.970 1.740 13.990 ;
        RECT 1.080 13.820 1.910 13.970 ;
        RECT 1.080 13.680 1.320 13.820 ;
        RECT 1.740 13.800 1.910 13.820 ;
        RECT 2.830 13.680 3.000 13.990 ;
        RECT 8.740 13.840 8.910 14.170 ;
        RECT 8.920 14.100 9.240 14.130 ;
        RECT 8.920 13.910 9.250 14.100 ;
        RECT 8.920 13.870 9.240 13.910 ;
        RECT 9.370 13.800 9.570 14.130 ;
        RECT 9.850 13.990 10.200 14.320 ;
        RECT 10.680 14.170 11.380 14.350 ;
        RECT 1.080 13.660 1.410 13.680 ;
        RECT 1.090 13.650 1.410 13.660 ;
        RECT 1.080 13.460 1.410 13.650 ;
        RECT 1.090 13.420 1.410 13.460 ;
        RECT 2.640 13.420 3.160 13.680 ;
        RECT 1.150 12.490 1.320 13.420 ;
        RECT 8.550 13.190 8.800 13.730 ;
        RECT 9.650 13.660 10.200 13.990 ;
        RECT 9.650 13.650 9.840 13.660 ;
        RECT 8.970 13.450 9.290 13.480 ;
        RECT 8.970 13.260 9.300 13.450 ;
        RECT 8.970 13.220 9.290 13.260 ;
        RECT 8.550 12.840 8.760 13.190 ;
        RECT 9.370 13.140 9.570 13.470 ;
        RECT 9.850 13.330 10.200 13.660 ;
        RECT 10.680 13.750 11.000 13.790 ;
        RECT 10.680 13.560 11.010 13.750 ;
        RECT 10.680 13.530 11.000 13.560 ;
        RECT 9.960 13.140 10.160 13.330 ;
        RECT 8.970 13.010 9.290 13.050 ;
        RECT 8.970 12.820 9.300 13.010 ;
        RECT 8.970 12.790 9.290 12.820 ;
        RECT 9.370 12.800 9.570 13.130 ;
        RECT 9.960 12.940 10.160 13.130 ;
        RECT 10.670 13.030 10.990 13.070 ;
        RECT 9.650 12.610 9.840 12.620 ;
        RECT 9.850 12.610 10.200 12.940 ;
        RECT 10.670 12.840 11.000 13.030 ;
        RECT 10.670 12.810 10.990 12.840 ;
        RECT 8.740 12.100 8.910 12.430 ;
        RECT 8.920 12.360 9.240 12.400 ;
        RECT 8.920 12.170 9.250 12.360 ;
        RECT 8.920 12.140 9.240 12.170 ;
        RECT 9.370 12.140 9.570 12.470 ;
        RECT 9.650 12.280 10.200 12.610 ;
        RECT 9.850 12.020 10.200 12.280 ;
        RECT 9.850 11.950 10.220 12.020 ;
        RECT 10.030 11.790 10.220 11.950 ;
        RECT 10.680 11.890 11.380 12.070 ;
        RECT 1.160 9.550 1.330 11.330 ;
        RECT 8.740 10.840 8.910 11.170 ;
        RECT 8.920 11.100 9.240 11.130 ;
        RECT 8.920 10.910 9.250 11.100 ;
        RECT 8.920 10.870 9.240 10.910 ;
        RECT 9.370 10.800 9.570 11.130 ;
        RECT 9.850 10.990 10.200 11.320 ;
        RECT 9.650 10.660 10.200 10.990 ;
        RECT 10.690 10.820 11.390 11.470 ;
        RECT 9.650 10.650 9.840 10.660 ;
        RECT 4.400 10.550 4.720 10.590 ;
        RECT 4.390 10.360 4.720 10.550 ;
        RECT 4.400 10.350 4.720 10.360 ;
        RECT 4.390 10.330 4.720 10.350 ;
        RECT 8.970 10.450 9.290 10.480 ;
        RECT 4.390 10.020 4.560 10.330 ;
        RECT 8.970 10.260 9.300 10.450 ;
        RECT 8.970 10.220 9.290 10.260 ;
        RECT 9.370 10.140 9.570 10.470 ;
        RECT 9.850 10.330 10.200 10.660 ;
        RECT 10.590 10.590 11.390 10.820 ;
        RECT 10.590 10.560 10.910 10.590 ;
        RECT 9.960 10.140 10.160 10.330 ;
        RECT 10.690 9.980 11.400 10.150 ;
        RECT 4.550 9.720 4.870 9.760 ;
        RECT 4.540 9.530 4.870 9.720 ;
        RECT 11.040 9.700 11.400 9.980 ;
        RECT 11.040 9.530 11.370 9.700 ;
        RECT 4.550 9.500 4.870 9.530 ;
        RECT 11.480 9.440 11.810 9.610 ;
        RECT 3.740 8.900 4.060 8.930 ;
        RECT 3.740 8.710 4.070 8.900 ;
        RECT 3.740 8.670 4.060 8.710 ;
        RECT 3.720 6.950 3.900 8.010 ;
        RECT 4.470 7.620 4.790 7.650 ;
        RECT 4.470 7.550 4.800 7.620 ;
        RECT 4.330 7.430 4.800 7.550 ;
        RECT 4.330 7.420 4.790 7.430 ;
        RECT 4.450 7.390 4.790 7.420 ;
        RECT 4.450 7.320 4.500 7.390 ;
        RECT 4.370 6.990 4.540 7.320 ;
        RECT 4.770 6.790 4.850 6.870 ;
        RECT 4.910 6.790 5.100 6.910 ;
        RECT 4.770 6.700 5.100 6.790 ;
        RECT 4.910 6.680 5.100 6.700 ;
        RECT 7.350 3.520 7.530 5.570 ;
        RECT 8.080 5.310 8.410 5.480 ;
        RECT 8.160 3.530 8.330 5.310 ;
        RECT 7.350 0.470 7.530 2.520 ;
        RECT 8.080 2.260 8.410 2.430 ;
        RECT 8.160 0.480 8.330 2.260 ;
      LAYER mcon ;
        RECT 1.610 17.130 1.780 17.300 ;
        RECT 3.360 17.130 3.530 17.300 ;
        RECT 1.220 16.400 1.390 16.570 ;
        RECT 2.970 16.400 3.140 16.570 ;
        RECT 9.030 15.830 9.200 16.000 ;
        RECT 10.690 15.790 10.860 15.960 ;
        RECT 0.490 15.120 0.660 15.290 ;
        RECT 2.240 15.120 2.410 15.290 ;
        RECT 8.980 15.180 9.150 15.350 ;
        RECT 9.970 15.440 10.140 15.610 ;
        RECT 1.860 14.740 2.030 14.910 ;
        RECT 1.150 14.190 1.320 14.360 ;
        RECT 1.330 14.300 1.500 14.470 ;
        RECT 1.740 14.140 1.910 14.310 ;
        RECT 3.080 14.300 3.250 14.470 ;
        RECT 10.040 14.410 10.210 14.580 ;
        RECT 1.150 13.850 1.320 14.020 ;
        RECT 8.980 13.920 9.150 14.090 ;
        RECT 1.150 13.640 1.320 13.680 ;
        RECT 1.150 13.510 1.350 13.640 ;
        RECT 1.180 13.470 1.350 13.510 ;
        RECT 2.700 13.460 2.870 13.630 ;
        RECT 2.930 13.470 3.100 13.640 ;
        RECT 8.570 13.560 8.740 13.730 ;
        RECT 9.970 13.660 10.140 13.830 ;
        RECT 1.150 13.170 1.320 13.340 ;
        RECT 1.150 12.830 1.320 13.000 ;
        RECT 9.030 13.270 9.200 13.440 ;
        RECT 10.740 13.570 10.910 13.740 ;
        RECT 8.570 12.860 8.740 13.030 ;
        RECT 9.030 12.830 9.200 13.000 ;
        RECT 10.730 12.850 10.900 13.020 ;
        RECT 8.980 12.180 9.150 12.350 ;
        RECT 9.970 12.440 10.140 12.610 ;
        RECT 10.040 11.820 10.210 11.990 ;
        RECT 1.160 11.160 1.330 11.330 ;
        RECT 1.160 10.820 1.330 10.990 ;
        RECT 8.980 10.920 9.150 11.090 ;
        RECT 9.970 10.660 10.140 10.830 ;
        RECT 1.160 10.480 1.330 10.650 ;
        RECT 4.490 10.370 4.660 10.540 ;
        RECT 1.160 10.140 1.330 10.310 ;
        RECT 9.030 10.270 9.200 10.440 ;
        RECT 10.650 10.600 10.820 10.770 ;
        RECT 1.160 9.800 1.330 9.970 ;
        RECT 4.640 9.540 4.810 9.710 ;
        RECT 3.800 8.720 3.970 8.890 ;
        RECT 4.530 7.440 4.700 7.610 ;
        RECT 4.920 6.710 5.090 6.880 ;
      LAYER met1 ;
        RECT 1.580 17.070 1.810 17.360 ;
        RECT 3.330 17.070 3.560 17.360 ;
        RECT 1.150 16.330 1.470 16.650 ;
        RECT 1.500 15.800 1.710 17.040 ;
        RECT 2.900 16.330 3.220 16.650 ;
        RECT 3.250 15.800 3.460 17.040 ;
        RECT 8.960 16.000 9.280 16.080 ;
        RECT 1.500 15.480 1.830 15.800 ;
        RECT 3.250 15.480 3.580 15.800 ;
        RECT 8.960 15.760 9.530 16.000 ;
        RECT 0.420 15.050 0.740 15.370 ;
        RECT 1.500 15.270 1.710 15.480 ;
        RECT 2.170 15.050 2.490 15.370 ;
        RECT 3.250 15.270 3.460 15.480 ;
        RECT 9.190 15.430 9.530 15.760 ;
        RECT 8.910 15.110 9.530 15.430 ;
        RECT 1.790 14.670 2.110 14.990 ;
        RECT 1.120 14.560 1.650 14.570 ;
        RECT 1.120 14.550 1.910 14.560 ;
        RECT 1.120 14.250 1.940 14.550 ;
        RECT 1.120 13.960 1.970 14.250 ;
        RECT 3.000 14.220 3.320 14.540 ;
        RECT 9.190 14.160 9.530 15.110 ;
        RECT 1.120 13.710 1.940 13.960 ;
        RECT 8.910 13.840 9.530 14.160 ;
        RECT 1.100 13.390 1.760 13.710 ;
        RECT 2.630 13.390 3.170 13.710 ;
        RECT 1.120 9.530 1.760 13.390 ;
        RECT 8.520 12.850 8.840 13.770 ;
        RECT 9.190 13.510 9.530 13.840 ;
        RECT 8.960 13.190 9.530 13.510 ;
        RECT 9.190 13.080 9.530 13.190 ;
        RECT 8.550 12.840 8.840 12.850 ;
        RECT 8.960 12.760 9.530 13.080 ;
        RECT 9.190 12.430 9.530 12.760 ;
        RECT 8.910 12.110 9.530 12.430 ;
        RECT 9.190 11.160 9.530 12.110 ;
        RECT 8.910 10.840 9.530 11.160 ;
        RECT 4.410 10.300 4.730 10.620 ;
        RECT 9.190 10.510 9.530 10.840 ;
        RECT 8.960 10.280 9.530 10.510 ;
        RECT 9.860 15.670 10.130 15.990 ;
        RECT 10.620 15.720 10.940 16.040 ;
        RECT 9.860 15.380 10.170 15.670 ;
        RECT 9.860 14.640 10.130 15.380 ;
        RECT 9.860 14.350 10.240 14.640 ;
        RECT 9.860 13.890 10.130 14.350 ;
        RECT 9.860 13.600 10.170 13.890 ;
        RECT 9.860 12.670 10.130 13.600 ;
        RECT 10.670 13.500 10.990 13.820 ;
        RECT 10.660 12.780 10.980 13.100 ;
        RECT 9.860 12.380 10.170 12.670 ;
        RECT 9.860 12.050 10.130 12.380 ;
        RECT 9.860 11.760 10.240 12.050 ;
        RECT 9.860 10.890 10.130 11.760 ;
        RECT 9.860 10.600 10.170 10.890 ;
        RECT 9.860 10.290 10.130 10.600 ;
        RECT 10.580 10.530 10.900 10.850 ;
        RECT 8.960 10.190 9.280 10.280 ;
        RECT 1.340 9.520 1.760 9.530 ;
        RECT 4.560 9.470 4.880 9.790 ;
        RECT 3.730 8.640 4.050 8.960 ;
        RECT 4.810 8.530 5.020 8.740 ;
        RECT 4.810 8.210 5.140 8.530 ;
        RECT 4.460 7.360 4.780 7.680 ;
        RECT 4.810 6.970 5.020 8.210 ;
        RECT 4.890 6.650 5.120 6.940 ;
      LAYER via ;
        RECT 1.180 16.360 1.440 16.620 ;
        RECT 2.930 16.360 3.190 16.620 ;
        RECT 1.570 15.510 1.830 15.770 ;
        RECT 3.320 15.510 3.580 15.770 ;
        RECT 8.990 15.790 9.250 16.050 ;
        RECT 0.450 15.080 0.710 15.340 ;
        RECT 2.200 15.080 2.460 15.340 ;
        RECT 8.940 15.140 9.200 15.400 ;
        RECT 1.820 14.700 2.080 14.960 ;
        RECT 1.280 14.490 1.540 14.510 ;
        RECT 1.240 13.770 1.830 14.490 ;
        RECT 3.030 14.250 3.290 14.510 ;
        RECT 8.940 13.870 9.200 14.130 ;
        RECT 1.130 13.420 1.390 13.680 ;
        RECT 2.660 13.420 3.140 13.680 ;
        RECT 8.530 12.870 8.790 13.730 ;
        RECT 8.990 13.220 9.250 13.480 ;
        RECT 8.990 12.790 9.250 13.050 ;
        RECT 8.940 12.140 9.200 12.400 ;
        RECT 8.940 10.870 9.200 11.130 ;
        RECT 4.440 10.330 4.700 10.590 ;
        RECT 8.990 10.220 9.250 10.480 ;
        RECT 10.650 15.750 10.910 16.010 ;
        RECT 10.700 13.530 10.960 13.790 ;
        RECT 10.690 12.810 10.950 13.070 ;
        RECT 10.610 10.560 10.870 10.820 ;
        RECT 4.590 9.500 4.850 9.760 ;
        RECT 3.760 8.670 4.020 8.930 ;
        RECT 4.880 8.240 5.140 8.500 ;
        RECT 4.490 7.390 4.750 7.650 ;
      LAYER met2 ;
        RECT 1.150 16.460 1.460 16.660 ;
        RECT 2.900 16.460 3.210 16.660 ;
        RECT 0.920 16.230 1.790 16.460 ;
        RECT 2.670 16.230 3.540 16.460 ;
        RECT 0.920 16.220 1.350 16.230 ;
        RECT 2.670 16.220 3.100 16.230 ;
        RECT 1.540 15.680 1.860 15.770 ;
        RECT 3.290 15.680 3.610 15.770 ;
        RECT 1.400 15.430 1.870 15.680 ;
        RECT 3.150 15.430 3.620 15.680 ;
        RECT 0.420 15.050 0.730 15.380 ;
        RECT 2.170 15.050 2.480 15.380 ;
        RECT 8.470 15.000 8.800 15.210 ;
        RECT 2.430 13.540 3.310 13.790 ;
        RECT 6.350 13.780 6.600 14.150 ;
        RECT 8.470 14.060 8.800 14.270 ;
        RECT 2.630 13.510 3.170 13.540 ;
        RECT 2.630 13.390 4.970 13.510 ;
        RECT 2.780 13.290 4.970 13.390 ;
        RECT 6.380 12.930 6.590 13.220 ;
        RECT 8.470 12.000 8.800 12.210 ;
        RECT 8.470 11.060 8.800 11.270 ;
        RECT 4.820 10.850 6.590 11.050 ;
        RECT 3.250 10.500 3.410 10.680 ;
        RECT 3.230 10.490 3.410 10.500 ;
        RECT 3.010 10.360 3.410 10.490 ;
        RECT 4.420 10.470 4.730 10.630 ;
        RECT 3.010 9.870 3.370 10.360 ;
        RECT 3.990 10.250 4.870 10.470 ;
        RECT 3.990 10.220 6.590 10.250 ;
        RECT 4.530 10.040 6.590 10.220 ;
        RECT 4.570 9.610 4.880 9.800 ;
        RECT 4.530 9.360 5.080 9.610 ;
        RECT 3.730 8.630 4.040 8.960 ;
        RECT 4.710 8.330 5.180 8.580 ;
        RECT 4.850 8.240 5.170 8.330 ;
        RECT 4.230 7.780 4.660 7.790 ;
        RECT 4.230 7.550 5.100 7.780 ;
        RECT 4.460 7.350 4.770 7.550 ;
  END
END sky130_hilas_TA2SignalBiasCell

MACRO sky130_hilas_Tgate4Single01
  CLASS CORE ;
  FOREIGN sky130_hilas_Tgate4Single01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.390 BY 10.470 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPWR
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 0.740 2.260 0.940 2.300 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.740 8.270 0.940 8.310 ;
    END
  END VPWR
  PIN INPUT1_2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 5.390 0.050 5.590 ;
    END
  END INPUT1_2
  PIN SELECT2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.000 6.370 0.060 6.570 ;
    END
  END SELECT2
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 4.250 8.250 4.440 8.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.250 2.260 4.440 2.320 ;
    END
  END VGND
  PIN OUTPUT2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.690 6.370 4.760 6.570 ;
    END
  END OUTPUT2
  PIN OUTPUT4
    PORT
      LAYER met2 ;
        RECT 4.690 3.170 4.760 3.370 ;
    END
  END OUTPUT4
  PIN OUTPUT3
    PORT
      LAYER met2 ;
        RECT 4.690 3.900 4.760 4.100 ;
    END
  END OUTPUT3
  PIN OUTPUT1
    PORT
      LAYER met2 ;
        RECT 4.690 7.100 4.760 7.300 ;
    END
  END OUTPUT1
  PIN INPUT1_4
    PORT
      LAYER met2 ;
        RECT 0.000 2.190 0.050 2.390 ;
    END
  END INPUT1_4
  PIN SELECT4
    PORT
      LAYER met2 ;
        RECT 0.000 3.170 0.060 3.370 ;
    END
  END SELECT4
  PIN SELECT3
    PORT
      LAYER met2 ;
        RECT 0.000 3.900 0.060 4.100 ;
    END
  END SELECT3
  PIN INPUT1_3
    PORT
      LAYER met2 ;
        RECT 0.000 4.880 0.050 5.080 ;
    END
  END INPUT1_3
  PIN SELECT1
    PORT
      LAYER met2 ;
        RECT 0.000 7.100 0.060 7.300 ;
    END
  END SELECT1
  PIN INPUT1_1
    PORT
      LAYER met2 ;
        RECT 0.000 8.080 0.050 8.280 ;
    END
  END INPUT1_1
  OBS
      LAYER nwell ;
        RECT 5.040 9.790 6.180 10.380 ;
        RECT 4.550 8.950 6.180 9.790 ;
        RECT 2.750 7.930 5.510 8.700 ;
        RECT 0.120 7.520 0.130 7.900 ;
        RECT 2.750 7.760 4.740 7.930 ;
        RECT 2.750 7.140 4.730 7.760 ;
        RECT 5.040 7.140 6.180 7.180 ;
        RECT 2.750 7.090 6.180 7.140 ;
        RECT 5.040 6.590 6.180 7.090 ;
        RECT 4.550 6.580 6.180 6.590 ;
        RECT 2.750 5.750 6.180 6.580 ;
        RECT 2.750 5.740 4.740 5.750 ;
        RECT 2.750 4.730 5.510 5.740 ;
        RECT 2.750 4.720 4.740 4.730 ;
        RECT 2.750 3.890 6.180 4.720 ;
        RECT 4.550 3.880 6.180 3.890 ;
        RECT 5.040 3.380 6.180 3.880 ;
        RECT 2.750 3.330 6.180 3.380 ;
        RECT 2.750 2.710 4.730 3.330 ;
        RECT 5.040 3.290 6.180 3.330 ;
        RECT 2.750 2.540 4.740 2.710 ;
        RECT 2.750 1.770 5.510 2.540 ;
        RECT 4.550 0.680 6.180 1.520 ;
        RECT 5.040 0.090 6.180 0.680 ;
      LAYER li1 ;
        RECT 2.940 9.880 3.580 10.060 ;
        RECT 3.960 9.890 4.310 10.060 ;
        RECT 4.410 10.050 4.600 10.160 ;
        RECT 4.410 9.930 4.740 10.050 ;
        RECT 4.490 9.850 4.740 9.930 ;
        RECT 5.040 9.880 6.180 10.060 ;
        RECT 3.340 9.500 3.510 9.510 ;
        RECT 3.340 9.460 3.740 9.500 ;
        RECT 3.340 9.270 3.750 9.460 ;
        RECT 3.950 9.430 4.140 9.540 ;
        RECT 3.950 9.310 4.290 9.430 ;
        RECT 3.340 9.240 3.740 9.270 ;
        RECT 4.000 9.260 4.290 9.310 ;
        RECT 3.340 9.210 3.510 9.240 ;
        RECT 4.570 9.170 4.740 9.850 ;
        RECT 5.080 9.500 5.250 9.510 ;
        RECT 5.080 9.460 5.410 9.500 ;
        RECT 5.080 9.270 5.420 9.460 ;
        RECT 6.060 9.440 6.250 9.550 ;
        RECT 5.940 9.430 6.250 9.440 ;
        RECT 5.690 9.320 6.250 9.430 ;
        RECT 5.080 9.240 5.410 9.270 ;
        RECT 5.690 9.260 6.070 9.320 ;
        RECT 5.080 9.210 5.250 9.240 ;
        RECT 2.960 8.380 3.170 8.810 ;
        RECT 2.980 8.360 3.150 8.380 ;
        RECT 3.480 8.240 3.670 8.350 ;
        RECT 3.480 8.120 3.900 8.240 ;
        RECT 3.380 8.070 3.900 8.120 ;
        RECT 4.250 8.070 5.510 8.250 ;
        RECT 3.380 7.990 3.570 8.070 ;
        RECT 3.360 7.960 3.570 7.990 ;
        RECT 3.350 7.950 3.570 7.960 ;
        RECT 4.740 7.950 5.070 8.070 ;
        RECT 3.230 7.900 3.570 7.950 ;
        RECT 3.100 7.870 3.570 7.900 ;
        RECT 3.060 7.840 3.570 7.870 ;
        RECT 3.060 7.780 3.550 7.840 ;
        RECT 3.060 7.730 3.400 7.780 ;
        RECT 3.060 7.710 3.320 7.730 ;
        RECT 3.060 7.690 3.290 7.710 ;
        RECT 3.060 7.650 3.270 7.690 ;
        RECT 3.060 7.370 3.230 7.650 ;
        RECT 2.940 6.680 3.580 6.860 ;
        RECT 3.960 6.690 4.310 6.860 ;
        RECT 4.410 6.850 4.600 6.960 ;
        RECT 4.410 6.730 4.740 6.850 ;
        RECT 4.490 6.650 4.740 6.730 ;
        RECT 5.040 6.680 6.180 6.860 ;
        RECT 3.340 6.300 3.510 6.310 ;
        RECT 3.060 6.020 3.230 6.300 ;
        RECT 3.340 6.260 3.740 6.300 ;
        RECT 3.340 6.070 3.750 6.260 ;
        RECT 3.950 6.230 4.140 6.340 ;
        RECT 3.950 6.110 4.290 6.230 ;
        RECT 3.340 6.040 3.740 6.070 ;
        RECT 4.000 6.060 4.290 6.110 ;
        RECT 3.060 5.980 3.270 6.020 ;
        RECT 3.340 6.010 3.510 6.040 ;
        RECT 3.060 5.960 3.290 5.980 ;
        RECT 4.570 5.970 4.740 6.650 ;
        RECT 5.080 6.300 5.250 6.310 ;
        RECT 5.080 6.260 5.410 6.300 ;
        RECT 5.080 6.070 5.420 6.260 ;
        RECT 6.060 6.240 6.250 6.350 ;
        RECT 5.940 6.230 6.250 6.240 ;
        RECT 5.690 6.120 6.250 6.230 ;
        RECT 5.080 6.040 5.410 6.070 ;
        RECT 5.690 6.060 6.070 6.120 ;
        RECT 5.080 6.010 5.250 6.040 ;
        RECT 3.060 5.940 3.320 5.960 ;
        RECT 3.060 5.890 3.400 5.940 ;
        RECT 3.060 5.830 3.550 5.890 ;
        RECT 3.060 5.800 3.570 5.830 ;
        RECT 3.100 5.770 3.570 5.800 ;
        RECT 3.230 5.720 3.570 5.770 ;
        RECT 3.350 5.710 3.570 5.720 ;
        RECT 3.360 5.680 3.570 5.710 ;
        RECT 2.960 4.860 3.170 5.610 ;
        RECT 3.380 5.600 3.570 5.680 ;
        RECT 4.740 5.600 5.070 5.720 ;
        RECT 3.380 5.550 3.900 5.600 ;
        RECT 3.480 5.430 3.900 5.550 ;
        RECT 3.480 5.320 3.670 5.430 ;
        RECT 4.250 5.420 5.510 5.600 ;
        RECT 3.480 5.040 3.670 5.150 ;
        RECT 3.480 4.920 3.900 5.040 ;
        RECT 3.380 4.870 3.900 4.920 ;
        RECT 4.250 4.870 5.510 5.050 ;
        RECT 3.380 4.790 3.570 4.870 ;
        RECT 3.360 4.760 3.570 4.790 ;
        RECT 3.350 4.750 3.570 4.760 ;
        RECT 4.740 4.750 5.070 4.870 ;
        RECT 3.230 4.700 3.570 4.750 ;
        RECT 3.100 4.670 3.570 4.700 ;
        RECT 3.060 4.640 3.570 4.670 ;
        RECT 3.060 4.580 3.550 4.640 ;
        RECT 3.060 4.530 3.400 4.580 ;
        RECT 3.060 4.510 3.320 4.530 ;
        RECT 3.060 4.490 3.290 4.510 ;
        RECT 3.060 4.450 3.270 4.490 ;
        RECT 3.060 4.170 3.230 4.450 ;
        RECT 3.340 4.430 3.510 4.460 ;
        RECT 3.340 4.400 3.740 4.430 ;
        RECT 3.340 4.210 3.750 4.400 ;
        RECT 4.000 4.360 4.290 4.410 ;
        RECT 3.950 4.240 4.290 4.360 ;
        RECT 3.340 4.170 3.740 4.210 ;
        RECT 3.340 4.160 3.510 4.170 ;
        RECT 3.950 4.130 4.140 4.240 ;
        RECT 4.570 3.820 4.740 4.500 ;
        RECT 5.080 4.430 5.250 4.460 ;
        RECT 5.080 4.400 5.410 4.430 ;
        RECT 5.080 4.210 5.420 4.400 ;
        RECT 5.690 4.350 6.070 4.410 ;
        RECT 5.690 4.240 6.250 4.350 ;
        RECT 5.940 4.230 6.250 4.240 ;
        RECT 5.080 4.170 5.410 4.210 ;
        RECT 5.080 4.160 5.250 4.170 ;
        RECT 6.060 4.120 6.250 4.230 ;
        RECT 2.940 3.610 3.580 3.790 ;
        RECT 3.960 3.610 4.310 3.780 ;
        RECT 4.490 3.740 4.740 3.820 ;
        RECT 4.410 3.620 4.740 3.740 ;
        RECT 4.410 3.510 4.600 3.620 ;
        RECT 5.040 3.610 6.180 3.790 ;
        RECT 3.060 2.820 3.230 3.100 ;
        RECT 3.060 2.780 3.270 2.820 ;
        RECT 3.060 2.760 3.290 2.780 ;
        RECT 3.060 2.740 3.320 2.760 ;
        RECT 3.060 2.690 3.400 2.740 ;
        RECT 3.060 2.630 3.550 2.690 ;
        RECT 3.060 2.600 3.570 2.630 ;
        RECT 3.100 2.570 3.570 2.600 ;
        RECT 3.230 2.520 3.570 2.570 ;
        RECT 3.350 2.510 3.570 2.520 ;
        RECT 3.360 2.480 3.570 2.510 ;
        RECT 3.380 2.400 3.570 2.480 ;
        RECT 4.740 2.400 5.070 2.520 ;
        RECT 3.380 2.350 3.900 2.400 ;
        RECT 3.480 2.230 3.900 2.350 ;
        RECT 3.480 2.120 3.670 2.230 ;
        RECT 4.250 2.220 5.510 2.400 ;
        RECT 2.980 2.090 3.150 2.110 ;
        RECT 2.960 1.660 3.170 2.090 ;
        RECT 3.340 1.230 3.510 1.260 ;
        RECT 3.340 1.200 3.740 1.230 ;
        RECT 3.340 1.010 3.750 1.200 ;
        RECT 4.000 1.160 4.290 1.210 ;
        RECT 3.950 1.040 4.290 1.160 ;
        RECT 3.340 0.970 3.740 1.010 ;
        RECT 3.340 0.960 3.510 0.970 ;
        RECT 3.950 0.930 4.140 1.040 ;
        RECT 4.570 0.620 4.740 1.300 ;
        RECT 5.080 1.230 5.250 1.260 ;
        RECT 5.080 1.200 5.410 1.230 ;
        RECT 5.080 1.010 5.420 1.200 ;
        RECT 5.690 1.150 6.070 1.210 ;
        RECT 5.690 1.040 6.250 1.150 ;
        RECT 5.940 1.030 6.250 1.040 ;
        RECT 5.080 0.970 5.410 1.010 ;
        RECT 5.080 0.960 5.250 0.970 ;
        RECT 6.060 0.920 6.250 1.030 ;
        RECT 2.940 0.410 3.580 0.590 ;
        RECT 3.960 0.410 4.310 0.580 ;
        RECT 4.490 0.540 4.740 0.620 ;
        RECT 4.410 0.420 4.740 0.540 ;
        RECT 4.410 0.310 4.600 0.420 ;
        RECT 5.040 0.410 6.180 0.590 ;
      LAYER mcon ;
        RECT 4.420 9.960 4.590 10.130 ;
        RECT 3.480 9.280 3.650 9.450 ;
        RECT 3.960 9.340 4.130 9.510 ;
        RECT 5.150 9.280 5.320 9.450 ;
        RECT 6.070 9.350 6.240 9.520 ;
        RECT 3.490 8.150 3.660 8.320 ;
        RECT 4.420 6.760 4.590 6.930 ;
        RECT 3.480 6.080 3.650 6.250 ;
        RECT 3.960 6.140 4.130 6.310 ;
        RECT 5.150 6.080 5.320 6.250 ;
        RECT 6.070 6.150 6.240 6.320 ;
        RECT 2.980 5.140 3.150 5.330 ;
        RECT 3.490 5.350 3.660 5.520 ;
        RECT 3.490 4.950 3.660 5.120 ;
        RECT 3.480 4.220 3.650 4.390 ;
        RECT 3.960 4.160 4.130 4.330 ;
        RECT 5.150 4.220 5.320 4.390 ;
        RECT 6.070 4.150 6.240 4.320 ;
        RECT 4.420 3.540 4.590 3.710 ;
        RECT 3.490 2.150 3.660 2.320 ;
        RECT 2.980 1.940 3.150 2.110 ;
        RECT 3.480 1.020 3.650 1.190 ;
        RECT 3.960 0.960 4.130 1.130 ;
        RECT 5.150 1.020 5.320 1.190 ;
        RECT 6.070 0.950 6.240 1.120 ;
        RECT 4.420 0.340 4.590 0.510 ;
      LAYER met1 ;
        RECT 3.750 10.300 4.010 10.400 ;
        RECT 3.650 10.230 4.010 10.300 ;
        RECT 3.650 9.980 4.020 10.230 ;
        RECT 3.830 9.570 4.020 9.980 ;
        RECT 4.310 10.190 4.500 10.470 ;
        RECT 4.310 9.900 4.620 10.190 ;
        RECT 5.980 10.090 6.240 10.390 ;
        RECT 5.960 10.070 6.240 10.090 ;
        RECT 3.410 9.210 3.730 9.530 ;
        RECT 3.830 9.480 4.160 9.570 ;
        RECT 3.930 9.280 4.160 9.480 ;
        RECT 4.310 8.950 4.500 9.900 ;
        RECT 5.960 9.580 6.150 10.070 ;
        RECT 5.080 9.210 5.400 9.530 ;
        RECT 5.960 9.500 6.270 9.580 ;
        RECT 5.940 9.290 6.270 9.500 ;
        RECT 5.940 9.210 6.170 9.290 ;
        RECT 2.960 8.650 3.180 8.810 ;
        RECT 2.960 8.590 3.300 8.650 ;
        RECT 2.950 8.330 3.300 8.590 ;
        RECT 3.370 8.380 3.570 8.700 ;
        RECT 6.880 8.660 7.070 8.700 ;
        RECT 2.950 8.300 3.180 8.330 ;
        RECT 3.370 8.090 3.690 8.380 ;
        RECT 3.370 7.090 3.570 8.090 ;
        RECT 3.750 7.100 4.010 7.200 ;
        RECT 3.650 7.030 4.010 7.100 ;
        RECT 3.650 6.780 4.020 7.030 ;
        RECT 3.370 6.330 3.570 6.580 ;
        RECT 3.830 6.370 4.020 6.780 ;
        RECT 4.310 6.990 4.500 7.270 ;
        RECT 4.310 6.700 4.620 6.990 ;
        RECT 5.980 6.890 6.240 7.190 ;
        RECT 6.880 7.090 7.070 7.140 ;
        RECT 5.960 6.870 6.240 6.890 ;
        RECT 3.370 6.010 3.730 6.330 ;
        RECT 3.830 6.280 4.160 6.370 ;
        RECT 3.930 6.080 4.160 6.280 ;
        RECT 2.960 5.450 3.180 5.610 ;
        RECT 3.370 5.580 3.570 6.010 ;
        RECT 4.310 5.750 4.500 6.700 ;
        RECT 5.960 6.380 6.150 6.870 ;
        RECT 6.880 6.530 7.070 6.580 ;
        RECT 5.080 6.010 5.400 6.330 ;
        RECT 5.960 6.300 6.270 6.380 ;
        RECT 5.940 6.090 6.270 6.300 ;
        RECT 5.940 6.010 6.170 6.090 ;
        RECT 2.960 5.390 3.300 5.450 ;
        RECT 2.950 5.080 3.300 5.390 ;
        RECT 2.960 5.020 3.300 5.080 ;
        RECT 3.370 5.290 3.690 5.580 ;
        RECT 6.880 5.460 7.070 5.500 ;
        RECT 3.370 5.180 3.570 5.290 ;
        RECT 2.960 4.860 3.180 5.020 ;
        RECT 3.370 4.890 3.690 5.180 ;
        RECT 6.880 4.970 7.070 5.010 ;
        RECT 3.370 4.460 3.570 4.890 ;
        RECT 3.370 4.140 3.730 4.460 ;
        RECT 3.930 4.190 4.160 4.390 ;
        RECT 3.370 3.890 3.570 4.140 ;
        RECT 3.830 4.100 4.160 4.190 ;
        RECT 3.830 3.690 4.020 4.100 ;
        RECT 3.650 3.440 4.020 3.690 ;
        RECT 4.310 3.770 4.500 4.720 ;
        RECT 5.080 4.140 5.400 4.460 ;
        RECT 5.940 4.380 6.170 4.460 ;
        RECT 5.940 4.170 6.270 4.380 ;
        RECT 5.960 4.090 6.270 4.170 ;
        RECT 4.310 3.480 4.620 3.770 ;
        RECT 5.960 3.600 6.150 4.090 ;
        RECT 6.880 3.890 7.070 3.940 ;
        RECT 5.960 3.580 6.240 3.600 ;
        RECT 3.370 2.380 3.570 3.380 ;
        RECT 3.650 3.370 4.010 3.440 ;
        RECT 3.750 3.270 4.010 3.370 ;
        RECT 4.310 3.200 4.500 3.480 ;
        RECT 5.980 3.280 6.240 3.580 ;
        RECT 6.880 3.330 7.070 3.380 ;
        RECT 2.950 2.140 3.180 2.170 ;
        RECT 2.950 1.880 3.300 2.140 ;
        RECT 2.960 1.820 3.300 1.880 ;
        RECT 3.370 2.090 3.690 2.380 ;
        RECT 2.960 1.660 3.180 1.820 ;
        RECT 3.370 1.770 3.570 2.090 ;
        RECT 6.880 1.770 7.070 1.810 ;
        RECT 3.410 0.940 3.730 1.260 ;
        RECT 3.930 0.990 4.160 1.190 ;
        RECT 3.830 0.900 4.160 0.990 ;
        RECT 3.830 0.490 4.020 0.900 ;
        RECT 3.650 0.240 4.020 0.490 ;
        RECT 4.310 0.570 4.500 1.520 ;
        RECT 5.080 0.940 5.400 1.260 ;
        RECT 5.940 1.180 6.170 1.260 ;
        RECT 5.940 0.970 6.270 1.180 ;
        RECT 5.960 0.890 6.270 0.970 ;
        RECT 4.310 0.280 4.620 0.570 ;
        RECT 5.960 0.400 6.150 0.890 ;
        RECT 5.960 0.380 6.240 0.400 ;
        RECT 3.650 0.170 4.010 0.240 ;
        RECT 3.750 0.070 4.010 0.170 ;
        RECT 4.310 0.000 4.500 0.280 ;
        RECT 5.980 0.080 6.240 0.380 ;
      LAYER via ;
        RECT 3.750 10.110 4.010 10.370 ;
        RECT 5.980 10.100 6.240 10.360 ;
        RECT 3.440 9.240 3.700 9.500 ;
        RECT 5.110 9.240 5.370 9.500 ;
        RECT 3.040 8.360 3.300 8.620 ;
        RECT 3.750 6.910 4.010 7.170 ;
        RECT 5.980 6.900 6.240 7.160 ;
        RECT 3.440 6.040 3.700 6.300 ;
        RECT 5.110 6.040 5.370 6.300 ;
        RECT 3.040 5.050 3.300 5.420 ;
        RECT 3.440 4.170 3.700 4.430 ;
        RECT 3.750 3.300 4.010 3.560 ;
        RECT 5.110 4.170 5.370 4.430 ;
        RECT 5.980 3.310 6.240 3.570 ;
        RECT 3.040 1.850 3.300 2.110 ;
        RECT 3.440 0.970 3.700 1.230 ;
        RECT 3.750 0.100 4.010 0.360 ;
        RECT 5.110 0.970 5.370 1.230 ;
        RECT 5.980 0.110 6.240 0.370 ;
      LAYER met2 ;
        RECT 3.720 10.240 4.040 10.370 ;
        RECT 5.950 10.240 6.270 10.360 ;
        RECT 2.940 10.040 4.820 10.240 ;
        RECT 5.810 10.100 6.270 10.240 ;
        RECT 5.810 10.040 6.180 10.100 ;
        RECT 3.410 9.260 3.720 9.540 ;
        RECT 2.940 9.210 3.720 9.260 ;
        RECT 4.550 9.260 4.770 9.270 ;
        RECT 5.080 9.260 5.390 9.540 ;
        RECT 2.940 9.060 3.510 9.210 ;
        RECT 4.550 9.060 6.180 9.260 ;
        RECT 4.550 9.050 4.770 9.060 ;
        RECT 3.010 8.430 3.330 8.620 ;
        RECT 2.630 8.360 3.330 8.430 ;
        RECT 2.630 8.230 3.240 8.360 ;
        RECT 7.320 8.230 7.390 8.430 ;
        RECT 3.500 7.450 4.620 7.460 ;
        RECT 2.630 7.250 4.620 7.450 ;
        RECT 3.500 7.240 4.620 7.250 ;
        RECT 3.720 7.040 4.040 7.170 ;
        RECT 5.950 7.040 6.270 7.160 ;
        RECT 2.940 6.840 4.820 7.040 ;
        RECT 5.810 6.900 6.270 7.040 ;
        RECT 5.810 6.840 6.180 6.900 ;
        RECT 3.500 6.420 4.620 6.430 ;
        RECT 2.630 6.220 4.620 6.420 ;
        RECT 3.410 6.210 4.620 6.220 ;
        RECT 3.410 6.060 3.720 6.210 ;
        RECT 2.940 6.010 3.720 6.060 ;
        RECT 4.550 6.060 4.770 6.070 ;
        RECT 5.080 6.060 5.390 6.340 ;
        RECT 2.940 5.860 3.510 6.010 ;
        RECT 4.550 5.860 6.180 6.060 ;
        RECT 4.550 5.850 4.770 5.860 ;
        RECT 2.630 5.420 3.240 5.440 ;
        RECT 2.630 5.240 3.330 5.420 ;
        RECT 7.320 5.240 7.390 5.440 ;
        RECT 3.010 5.230 3.330 5.240 ;
        RECT 2.630 5.050 3.330 5.230 ;
        RECT 2.630 5.030 3.240 5.050 ;
        RECT 7.320 5.030 7.390 5.230 ;
        RECT 4.550 4.610 4.770 4.620 ;
        RECT 2.940 4.460 3.510 4.610 ;
        RECT 2.940 4.410 3.720 4.460 ;
        RECT 3.410 4.260 3.720 4.410 ;
        RECT 4.550 4.410 6.180 4.610 ;
        RECT 4.550 4.400 4.770 4.410 ;
        RECT 3.410 4.250 4.620 4.260 ;
        RECT 2.630 4.050 4.620 4.250 ;
        RECT 5.080 4.130 5.390 4.410 ;
        RECT 3.500 4.040 4.620 4.050 ;
        RECT 2.940 3.430 4.820 3.630 ;
        RECT 5.810 3.570 6.180 3.630 ;
        RECT 5.810 3.430 6.270 3.570 ;
        RECT 3.720 3.300 4.040 3.430 ;
        RECT 5.950 3.310 6.270 3.430 ;
        RECT 3.500 3.220 4.620 3.230 ;
        RECT 2.630 3.020 4.620 3.220 ;
        RECT 3.500 3.010 4.620 3.020 ;
        RECT 2.630 2.110 3.240 2.240 ;
        RECT 2.630 2.040 3.330 2.110 ;
        RECT 7.320 2.040 7.390 2.240 ;
        RECT 3.010 1.850 3.330 2.040 ;
        RECT 4.550 1.410 4.770 1.420 ;
        RECT 2.940 1.260 3.510 1.410 ;
        RECT 2.940 1.210 3.720 1.260 ;
        RECT 3.410 0.930 3.720 1.210 ;
        RECT 4.550 1.210 6.180 1.410 ;
        RECT 4.550 1.200 4.770 1.210 ;
        RECT 5.080 0.930 5.390 1.210 ;
        RECT 2.940 0.230 4.820 0.430 ;
        RECT 5.810 0.370 6.180 0.430 ;
        RECT 5.810 0.230 6.270 0.370 ;
        RECT 3.720 0.100 4.040 0.230 ;
        RECT 5.950 0.110 6.270 0.230 ;
  END
END sky130_hilas_Tgate4Single01

MACRO sky130_hilas_VinjDecode2to4
  CLASS CORE ;
  FOREIGN sky130_hilas_VinjDecode2to4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.320 BY 7.560 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN OUTPUT00
    PORT
      LAYER met2 ;
        RECT 12.820 6.270 12.950 6.440 ;
    END
  END OUTPUT00
  PIN OUTPUT01
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 12.940 5.010 13.310 5.090 ;
        RECT 12.940 5.000 13.970 5.010 ;
        RECT 15.850 5.000 16.160 5.160 ;
        RECT 12.940 4.930 16.320 5.000 ;
        RECT 12.820 4.830 16.320 4.930 ;
        RECT 12.820 4.760 12.950 4.830 ;
    END
  END OUTPUT01
  PIN OUTPUT10
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 12.940 3.500 13.310 3.580 ;
        RECT 12.940 3.490 13.970 3.500 ;
        RECT 15.850 3.490 16.160 3.650 ;
        RECT 12.940 3.420 16.320 3.490 ;
        RECT 12.820 3.320 16.320 3.420 ;
        RECT 12.820 3.250 12.950 3.320 ;
    END
  END OUTPUT10
  PIN OUTPUT11
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 12.940 1.990 13.310 2.070 ;
        RECT 12.940 1.980 13.970 1.990 ;
        RECT 15.850 1.980 16.160 2.140 ;
        RECT 12.940 1.920 16.320 1.980 ;
        RECT 12.820 1.810 16.320 1.920 ;
        RECT 12.820 1.750 12.950 1.810 ;
    END
  END OUTPUT11
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 11.660 7.510 11.930 7.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.660 1.540 11.930 1.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.180 7.470 3.410 7.560 ;
    END
  END VGND
  PIN VINJ
    ANTENNADIFFAREA 0.691200 ;
    PORT
      LAYER met1 ;
        RECT 6.540 1.590 6.770 6.120 ;
        RECT 6.690 1.540 6.910 1.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.690 7.490 6.910 7.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.610 7.480 0.830 7.560 ;
    END
  END VINJ
  PIN IN2
    PORT
      LAYER met2 ;
        RECT 0.000 5.480 0.110 5.660 ;
    END
  END IN2
  PIN IN1
    PORT
      LAYER met2 ;
        RECT 0.000 6.990 0.110 7.170 ;
    END
  END IN1
  PIN ENABLE
    PORT
      LAYER met2 ;
        RECT 0.000 3.970 0.110 4.150 ;
    END
  END ENABLE
  OBS
      LAYER nwell ;
        RECT 6.690 7.490 6.910 7.550 ;
        RECT 3.360 1.500 5.340 6.160 ;
        RECT 6.690 1.540 6.910 1.590 ;
        RECT 9.450 0.000 12.890 6.160 ;
      LAYER li1 ;
        RECT 3.980 5.730 4.150 5.870 ;
        RECT 10.070 5.730 10.240 5.870 ;
        RECT 10.800 5.750 10.970 5.830 ;
        RECT 11.610 5.750 11.780 5.830 ;
        RECT 13.150 5.790 13.320 5.910 ;
        RECT 3.980 5.560 4.170 5.730 ;
        RECT 3.980 5.460 4.150 5.560 ;
        RECT 3.550 5.080 3.720 5.180 ;
        RECT 3.530 4.910 3.720 5.080 ;
        RECT 3.550 4.850 3.720 4.910 ;
        RECT 3.970 5.120 4.140 5.180 ;
        RECT 3.970 4.850 4.220 5.120 ;
        RECT 4.710 5.100 4.960 5.180 ;
        RECT 4.710 4.930 6.010 5.100 ;
        RECT 6.570 5.090 6.740 5.720 ;
        RECT 10.070 5.560 10.260 5.730 ;
        RECT 10.070 5.460 10.240 5.560 ;
        RECT 10.800 5.180 11.010 5.750 ;
        RECT 11.570 5.500 11.780 5.750 ;
        RECT 12.170 5.570 12.340 5.670 ;
        RECT 13.110 5.620 13.320 5.790 ;
        RECT 15.040 5.720 15.300 5.790 ;
        RECT 15.840 5.720 16.020 5.850 ;
        RECT 13.150 5.580 13.320 5.620 ;
        RECT 11.570 5.180 11.740 5.500 ;
        RECT 12.140 5.400 12.340 5.570 ;
        RECT 12.170 5.300 12.340 5.400 ;
        RECT 13.710 5.540 14.580 5.710 ;
        RECT 15.040 5.540 16.020 5.720 ;
        RECT 3.980 4.830 4.220 4.850 ;
        RECT 4.790 4.840 4.960 4.930 ;
        RECT 6.490 4.920 6.820 5.090 ;
        RECT 9.640 5.080 9.810 5.180 ;
        RECT 9.620 4.910 9.810 5.080 ;
        RECT 9.640 4.850 9.810 4.910 ;
        RECT 10.060 5.120 10.230 5.180 ;
        RECT 10.060 4.850 10.310 5.120 ;
        RECT 10.800 4.930 11.050 5.180 ;
        RECT 10.070 4.830 10.310 4.850 ;
        RECT 10.880 4.840 11.050 4.930 ;
        RECT 11.530 4.930 11.740 5.180 ;
        RECT 13.710 5.100 13.880 5.540 ;
        RECT 15.040 5.100 15.300 5.540 ;
        RECT 15.840 5.430 16.020 5.540 ;
        RECT 12.250 4.930 13.880 5.100 ;
        RECT 14.330 4.930 15.300 5.100 ;
        RECT 15.750 4.930 16.090 5.100 ;
        RECT 11.530 4.850 11.700 4.930 ;
        RECT 13.020 4.890 13.190 4.930 ;
        RECT 3.980 4.220 4.150 4.360 ;
        RECT 10.070 4.220 10.240 4.360 ;
        RECT 10.800 4.240 10.970 4.320 ;
        RECT 11.610 4.240 11.780 4.320 ;
        RECT 13.150 4.280 13.320 4.400 ;
        RECT 3.980 4.050 4.170 4.220 ;
        RECT 3.980 3.950 4.150 4.050 ;
        RECT 3.550 3.570 3.720 3.670 ;
        RECT 3.530 3.400 3.720 3.570 ;
        RECT 3.550 3.340 3.720 3.400 ;
        RECT 3.970 3.610 4.140 3.670 ;
        RECT 3.970 3.340 4.220 3.610 ;
        RECT 4.710 3.590 4.960 3.670 ;
        RECT 4.710 3.420 6.010 3.590 ;
        RECT 6.570 3.580 6.740 4.210 ;
        RECT 10.070 4.050 10.260 4.220 ;
        RECT 10.070 3.950 10.240 4.050 ;
        RECT 10.800 3.670 11.010 4.240 ;
        RECT 11.570 3.990 11.780 4.240 ;
        RECT 12.170 4.060 12.340 4.160 ;
        RECT 13.110 4.110 13.320 4.280 ;
        RECT 15.040 4.210 15.300 4.280 ;
        RECT 15.840 4.210 16.020 4.340 ;
        RECT 13.150 4.070 13.320 4.110 ;
        RECT 11.570 3.670 11.740 3.990 ;
        RECT 12.140 3.890 12.340 4.060 ;
        RECT 12.170 3.790 12.340 3.890 ;
        RECT 13.710 4.030 14.580 4.200 ;
        RECT 15.040 4.030 16.020 4.210 ;
        RECT 3.980 3.320 4.220 3.340 ;
        RECT 4.790 3.330 4.960 3.420 ;
        RECT 6.490 3.410 6.820 3.580 ;
        RECT 9.640 3.570 9.810 3.670 ;
        RECT 9.620 3.400 9.810 3.570 ;
        RECT 9.640 3.340 9.810 3.400 ;
        RECT 10.060 3.610 10.230 3.670 ;
        RECT 10.060 3.340 10.310 3.610 ;
        RECT 10.800 3.420 11.050 3.670 ;
        RECT 10.070 3.320 10.310 3.340 ;
        RECT 10.880 3.330 11.050 3.420 ;
        RECT 11.530 3.420 11.740 3.670 ;
        RECT 13.710 3.590 13.880 4.030 ;
        RECT 15.040 3.590 15.300 4.030 ;
        RECT 15.840 3.920 16.020 4.030 ;
        RECT 12.250 3.420 13.880 3.590 ;
        RECT 14.330 3.420 15.300 3.590 ;
        RECT 15.750 3.420 16.090 3.590 ;
        RECT 11.530 3.340 11.700 3.420 ;
        RECT 13.020 3.380 13.190 3.420 ;
        RECT 3.980 2.710 4.150 2.850 ;
        RECT 10.070 2.710 10.240 2.850 ;
        RECT 10.800 2.730 10.970 2.810 ;
        RECT 11.610 2.730 11.780 2.810 ;
        RECT 13.150 2.770 13.320 2.890 ;
        RECT 3.980 2.540 4.170 2.710 ;
        RECT 3.980 2.440 4.150 2.540 ;
        RECT 3.550 2.060 3.720 2.160 ;
        RECT 3.530 1.890 3.720 2.060 ;
        RECT 3.550 1.830 3.720 1.890 ;
        RECT 3.970 2.100 4.140 2.160 ;
        RECT 3.970 1.830 4.220 2.100 ;
        RECT 4.710 2.080 4.960 2.160 ;
        RECT 4.710 1.910 6.010 2.080 ;
        RECT 6.570 2.070 6.740 2.700 ;
        RECT 10.070 2.540 10.260 2.710 ;
        RECT 10.070 2.440 10.240 2.540 ;
        RECT 10.800 2.160 11.010 2.730 ;
        RECT 11.570 2.480 11.780 2.730 ;
        RECT 12.170 2.550 12.340 2.650 ;
        RECT 13.110 2.600 13.320 2.770 ;
        RECT 15.040 2.700 15.300 2.770 ;
        RECT 15.840 2.700 16.020 2.830 ;
        RECT 13.150 2.560 13.320 2.600 ;
        RECT 11.570 2.160 11.740 2.480 ;
        RECT 12.140 2.380 12.340 2.550 ;
        RECT 12.170 2.280 12.340 2.380 ;
        RECT 13.710 2.520 14.580 2.690 ;
        RECT 15.040 2.520 16.020 2.700 ;
        RECT 3.980 1.810 4.220 1.830 ;
        RECT 4.790 1.820 4.960 1.910 ;
        RECT 6.490 1.900 6.820 2.070 ;
        RECT 9.640 2.060 9.810 2.160 ;
        RECT 9.620 1.890 9.810 2.060 ;
        RECT 9.640 1.830 9.810 1.890 ;
        RECT 10.060 2.100 10.230 2.160 ;
        RECT 10.060 1.830 10.310 2.100 ;
        RECT 10.800 1.910 11.050 2.160 ;
        RECT 10.070 1.810 10.310 1.830 ;
        RECT 10.880 1.820 11.050 1.910 ;
        RECT 11.530 1.910 11.740 2.160 ;
        RECT 13.710 2.080 13.880 2.520 ;
        RECT 15.040 2.080 15.300 2.520 ;
        RECT 15.840 2.410 16.020 2.520 ;
        RECT 12.250 1.910 13.880 2.080 ;
        RECT 14.330 1.910 15.300 2.080 ;
        RECT 15.750 1.910 16.090 2.080 ;
        RECT 11.530 1.830 11.700 1.910 ;
        RECT 13.020 1.870 13.190 1.910 ;
        RECT 10.070 1.210 10.240 1.350 ;
        RECT 10.800 1.230 10.970 1.310 ;
        RECT 11.610 1.230 11.780 1.310 ;
        RECT 13.150 1.270 13.320 1.390 ;
        RECT 10.070 1.040 10.260 1.210 ;
        RECT 10.070 0.940 10.240 1.040 ;
        RECT 10.800 0.660 11.010 1.230 ;
        RECT 11.570 0.980 11.780 1.230 ;
        RECT 12.170 1.050 12.340 1.150 ;
        RECT 13.110 1.100 13.320 1.270 ;
        RECT 15.040 1.200 15.300 1.270 ;
        RECT 15.840 1.200 16.020 1.330 ;
        RECT 13.150 1.060 13.320 1.100 ;
        RECT 11.570 0.660 11.740 0.980 ;
        RECT 12.140 0.880 12.340 1.050 ;
        RECT 12.170 0.780 12.340 0.880 ;
        RECT 13.710 1.020 14.580 1.190 ;
        RECT 15.040 1.020 16.020 1.200 ;
        RECT 9.640 0.560 9.810 0.660 ;
        RECT 9.620 0.390 9.810 0.560 ;
        RECT 9.640 0.330 9.810 0.390 ;
        RECT 10.060 0.600 10.230 0.660 ;
        RECT 10.060 0.330 10.310 0.600 ;
        RECT 10.800 0.410 11.050 0.660 ;
        RECT 10.070 0.310 10.310 0.330 ;
        RECT 10.880 0.320 11.050 0.410 ;
        RECT 11.530 0.410 11.740 0.660 ;
        RECT 13.710 0.580 13.880 1.020 ;
        RECT 15.040 0.580 15.300 1.020 ;
        RECT 15.840 0.910 16.020 1.020 ;
        RECT 12.250 0.410 13.880 0.580 ;
        RECT 14.330 0.410 15.300 0.580 ;
        RECT 15.750 0.410 16.090 0.580 ;
        RECT 11.530 0.330 11.700 0.410 ;
        RECT 13.020 0.370 13.190 0.410 ;
      LAYER mcon ;
        RECT 4.000 5.560 4.170 5.730 ;
        RECT 10.090 5.560 10.260 5.730 ;
        RECT 6.570 5.200 6.740 5.370 ;
        RECT 4.010 4.880 4.180 5.050 ;
        RECT 5.350 4.930 5.520 5.100 ;
        RECT 10.100 4.880 10.270 5.050 ;
        RECT 15.070 5.220 15.250 5.400 ;
        RECT 4.000 4.050 4.170 4.220 ;
        RECT 10.090 4.050 10.260 4.220 ;
        RECT 6.570 3.690 6.740 3.860 ;
        RECT 4.010 3.370 4.180 3.540 ;
        RECT 5.350 3.420 5.520 3.590 ;
        RECT 10.100 3.370 10.270 3.540 ;
        RECT 15.070 3.710 15.250 3.890 ;
        RECT 4.000 2.540 4.170 2.710 ;
        RECT 10.090 2.540 10.260 2.710 ;
        RECT 6.570 2.180 6.740 2.350 ;
        RECT 4.010 1.860 4.180 2.030 ;
        RECT 5.350 1.910 5.520 2.080 ;
        RECT 10.100 1.860 10.270 2.030 ;
        RECT 15.070 2.200 15.250 2.380 ;
        RECT 10.090 1.040 10.260 1.210 ;
        RECT 10.100 0.360 10.270 0.530 ;
        RECT 15.070 0.700 15.250 0.880 ;
      LAYER met1 ;
        RECT 3.670 7.210 3.940 7.500 ;
        RECT 3.630 6.940 3.960 7.210 ;
        RECT 3.670 6.160 3.940 6.940 ;
        RECT 3.660 5.830 3.940 6.160 ;
        RECT 4.130 6.120 4.400 6.600 ;
        RECT 3.670 5.800 3.940 5.830 ;
        RECT 3.440 4.840 3.750 5.190 ;
        RECT 3.440 3.330 3.750 3.680 ;
        RECT 3.970 2.980 4.400 6.120 ;
        RECT 4.590 5.610 4.860 7.070 ;
        RECT 5.540 6.570 5.830 6.620 ;
        RECT 5.520 6.220 5.830 6.570 ;
        RECT 4.540 5.340 4.870 5.610 ;
        RECT 4.590 4.030 4.860 5.340 ;
        RECT 5.540 5.140 5.830 6.220 ;
        RECT 10.060 5.780 10.280 6.120 ;
        RECT 10.060 5.520 10.290 5.780 ;
        RECT 5.270 5.130 5.830 5.140 ;
        RECT 4.570 3.700 4.860 4.030 ;
        RECT 4.590 3.680 4.860 3.700 ;
        RECT 5.060 4.880 5.830 5.130 ;
        RECT 5.060 4.740 5.340 4.880 ;
        RECT 5.060 3.630 5.330 4.740 ;
        RECT 5.540 3.630 5.830 4.880 ;
        RECT 9.530 4.840 9.840 5.190 ;
        RECT 10.060 5.120 10.280 5.520 ;
        RECT 12.080 5.360 12.410 5.620 ;
        RECT 13.050 5.580 13.480 5.870 ;
        RECT 10.060 4.810 10.310 5.120 ;
        RECT 12.920 4.830 13.310 5.100 ;
        RECT 10.060 4.270 10.280 4.810 ;
        RECT 10.060 4.010 10.290 4.270 ;
        RECT 5.060 3.570 5.830 3.630 ;
        RECT 5.060 3.370 5.840 3.570 ;
        RECT 3.970 2.650 4.430 2.980 ;
        RECT 3.970 2.600 4.400 2.650 ;
        RECT 3.970 2.500 4.200 2.600 ;
        RECT 5.060 2.530 5.330 3.370 ;
        RECT 3.440 1.820 3.750 2.170 ;
        RECT 3.970 2.100 4.190 2.500 ;
        RECT 5.040 2.200 5.330 2.530 ;
        RECT 5.060 2.170 5.330 2.200 ;
        RECT 5.540 3.220 5.840 3.370 ;
        RECT 9.530 3.330 9.840 3.680 ;
        RECT 10.060 3.610 10.280 4.010 ;
        RECT 12.080 3.850 12.410 4.110 ;
        RECT 13.050 4.070 13.480 4.360 ;
        RECT 10.060 3.300 10.310 3.610 ;
        RECT 12.920 3.320 13.310 3.590 ;
        RECT 5.540 2.120 5.830 3.220 ;
        RECT 10.060 2.760 10.280 3.300 ;
        RECT 10.060 2.500 10.290 2.760 ;
        RECT 3.970 1.790 4.220 2.100 ;
        RECT 5.270 1.860 5.830 2.120 ;
        RECT 3.970 1.590 4.190 1.790 ;
        RECT 5.540 1.680 5.830 1.860 ;
        RECT 9.530 1.820 9.840 2.170 ;
        RECT 10.060 2.100 10.280 2.500 ;
        RECT 12.080 2.340 12.410 2.600 ;
        RECT 13.050 2.560 13.480 2.850 ;
        RECT 10.060 1.790 10.310 2.100 ;
        RECT 12.920 1.810 13.310 2.080 ;
        RECT 10.060 1.260 10.280 1.790 ;
        RECT 10.060 1.000 10.290 1.260 ;
        RECT 9.530 0.320 9.840 0.670 ;
        RECT 10.060 0.600 10.280 1.000 ;
        RECT 12.080 0.840 12.410 1.100 ;
        RECT 13.050 1.060 13.480 1.350 ;
        RECT 10.060 0.290 10.310 0.600 ;
        RECT 12.920 0.310 13.310 0.580 ;
        RECT 10.060 0.090 10.280 0.290 ;
        RECT 15.030 0.090 15.300 6.130 ;
        RECT 15.850 4.840 16.160 5.160 ;
        RECT 15.850 3.330 16.160 3.650 ;
        RECT 15.850 1.820 16.160 2.140 ;
        RECT 15.850 0.320 16.160 0.640 ;
      LAYER via ;
        RECT 3.660 6.940 3.930 7.210 ;
        RECT 4.590 6.750 4.860 7.020 ;
        RECT 3.660 5.860 3.930 6.130 ;
        RECT 4.130 6.260 4.400 6.530 ;
        RECT 3.470 4.870 3.730 5.130 ;
        RECT 5.520 6.250 5.810 6.540 ;
        RECT 4.570 5.340 4.840 5.610 ;
        RECT 4.120 4.180 4.390 4.450 ;
        RECT 3.470 3.360 3.730 3.620 ;
        RECT 4.570 3.730 4.840 4.000 ;
        RECT 5.300 5.040 5.560 5.140 ;
        RECT 5.070 5.000 5.560 5.040 ;
        RECT 5.070 4.880 5.820 5.000 ;
        RECT 5.070 4.770 5.340 4.880 ;
        RECT 5.560 4.740 5.820 4.880 ;
        RECT 9.560 4.870 9.820 5.130 ;
        RECT 12.120 5.360 12.380 5.620 ;
        RECT 13.110 5.610 13.370 5.870 ;
        RECT 12.980 4.830 13.240 5.090 ;
        RECT 5.300 3.540 5.560 3.630 ;
        RECT 5.300 3.370 5.840 3.540 ;
        RECT 4.160 2.680 4.430 2.950 ;
        RECT 3.470 1.850 3.730 2.110 ;
        RECT 5.040 2.230 5.310 2.500 ;
        RECT 5.550 3.250 5.840 3.370 ;
        RECT 9.560 3.360 9.820 3.620 ;
        RECT 12.120 3.850 12.380 4.110 ;
        RECT 13.110 4.100 13.370 4.360 ;
        RECT 12.980 3.320 13.240 3.580 ;
        RECT 5.300 2.000 5.560 2.120 ;
        RECT 5.300 1.860 5.830 2.000 ;
        RECT 5.540 1.710 5.830 1.860 ;
        RECT 9.560 1.850 9.820 2.110 ;
        RECT 12.120 2.340 12.380 2.600 ;
        RECT 13.110 2.590 13.370 2.850 ;
        RECT 12.980 1.810 13.240 2.070 ;
        RECT 9.560 0.350 9.820 0.610 ;
        RECT 12.120 0.840 12.380 1.100 ;
        RECT 13.110 1.090 13.370 1.350 ;
        RECT 12.980 0.310 13.240 0.570 ;
        RECT 15.880 4.870 16.140 5.130 ;
        RECT 15.880 3.360 16.140 3.620 ;
        RECT 15.880 1.850 16.140 2.110 ;
        RECT 15.880 0.350 16.140 0.610 ;
      LAYER met2 ;
        RECT 3.710 7.400 6.080 7.410 ;
        RECT 3.690 7.250 6.080 7.400 ;
        RECT 3.690 7.240 3.960 7.250 ;
        RECT 3.660 7.170 3.960 7.240 ;
        RECT 3.430 6.990 3.960 7.170 ;
        RECT 3.660 6.910 3.930 6.990 ;
        RECT 4.560 6.960 4.890 7.020 ;
        RECT 4.560 6.800 6.080 6.960 ;
        RECT 4.560 6.750 4.890 6.800 ;
        RECT 4.100 6.500 4.430 6.530 ;
        RECT 3.430 6.320 4.450 6.500 ;
        RECT 4.100 6.310 4.450 6.320 ;
        RECT 5.490 6.470 5.840 6.540 ;
        RECT 5.490 6.310 6.080 6.470 ;
        RECT 4.100 6.260 4.430 6.310 ;
        RECT 5.490 6.250 5.840 6.310 ;
        RECT 3.630 6.070 3.960 6.130 ;
        RECT 3.630 5.910 5.270 6.070 ;
        RECT 3.630 5.860 3.960 5.910 ;
        RECT 5.110 5.900 5.270 5.910 ;
        RECT 5.110 5.740 6.070 5.900 ;
        RECT 9.440 5.810 13.480 5.970 ;
        RECT 3.360 5.550 6.970 5.730 ;
        RECT 3.430 5.480 4.840 5.550 ;
        RECT 12.080 5.540 12.410 5.620 ;
        RECT 13.060 5.580 13.480 5.810 ;
        RECT 11.810 5.520 12.410 5.540 ;
        RECT 4.570 5.450 4.840 5.480 ;
        RECT 4.570 5.310 4.850 5.450 ;
        RECT 4.620 5.290 4.850 5.310 ;
        RECT 5.120 5.290 6.080 5.450 ;
        RECT 9.450 5.360 12.410 5.520 ;
        RECT 5.120 5.140 5.280 5.290 ;
        RECT 3.440 5.030 3.760 5.130 ;
        RECT 5.120 5.060 5.590 5.140 ;
        RECT 5.120 5.040 6.970 5.060 ;
        RECT 3.430 4.990 3.760 5.030 ;
        RECT 5.040 4.990 6.970 5.040 ;
        RECT 9.530 5.030 9.850 5.130 ;
        RECT 3.430 4.880 6.970 4.990 ;
        RECT 3.430 4.810 5.370 4.880 ;
        RECT 5.040 4.770 5.370 4.810 ;
        RECT 5.530 4.800 6.080 4.880 ;
        RECT 9.450 4.870 9.850 5.030 ;
        RECT 5.530 4.740 5.850 4.800 ;
        RECT 4.090 4.390 4.420 4.450 ;
        RECT 4.090 4.230 6.080 4.390 ;
        RECT 9.440 4.300 13.480 4.460 ;
        RECT 4.090 4.220 4.420 4.230 ;
        RECT 3.360 4.040 6.970 4.220 ;
        RECT 12.080 4.030 12.410 4.110 ;
        RECT 13.060 4.070 13.480 4.300 ;
        RECT 11.810 4.010 12.410 4.030 ;
        RECT 4.540 3.940 4.870 4.000 ;
        RECT 4.540 3.780 6.080 3.940 ;
        RECT 9.450 3.850 12.410 4.010 ;
        RECT 4.540 3.730 4.870 3.780 ;
        RECT 3.440 3.520 3.760 3.620 ;
        RECT 3.430 3.480 3.760 3.520 ;
        RECT 5.270 3.550 5.590 3.630 ;
        RECT 5.270 3.480 6.970 3.550 ;
        RECT 9.530 3.520 9.850 3.620 ;
        RECT 3.430 3.370 6.970 3.480 ;
        RECT 3.430 3.300 6.080 3.370 ;
        RECT 9.450 3.360 9.850 3.520 ;
        RECT 5.520 3.290 6.080 3.300 ;
        RECT 5.520 3.250 5.870 3.290 ;
        RECT 4.130 2.890 4.460 2.950 ;
        RECT 4.130 2.730 6.080 2.890 ;
        RECT 9.440 2.790 13.480 2.950 ;
        RECT 4.130 2.710 4.460 2.730 ;
        RECT 3.360 2.530 6.970 2.710 ;
        RECT 12.080 2.520 12.410 2.600 ;
        RECT 13.060 2.560 13.480 2.790 ;
        RECT 11.810 2.500 12.410 2.520 ;
        RECT 5.010 2.440 5.340 2.500 ;
        RECT 5.010 2.280 6.080 2.440 ;
        RECT 9.450 2.340 12.410 2.500 ;
        RECT 5.010 2.230 5.340 2.280 ;
        RECT 3.440 2.010 3.760 2.110 ;
        RECT 3.430 1.850 3.760 2.010 ;
        RECT 5.270 2.040 5.590 2.120 ;
        RECT 5.270 1.860 6.970 2.040 ;
        RECT 9.530 2.010 9.850 2.110 ;
        RECT 5.510 1.790 6.080 1.860 ;
        RECT 9.450 1.850 9.850 2.010 ;
        RECT 5.510 1.710 5.860 1.790 ;
        RECT 9.440 1.290 13.480 1.450 ;
        RECT 12.080 1.020 12.410 1.100 ;
        RECT 13.060 1.060 13.480 1.290 ;
        RECT 11.810 1.000 12.410 1.020 ;
        RECT 9.450 0.840 12.410 1.000 ;
        RECT 9.530 0.510 9.850 0.610 ;
        RECT 9.450 0.350 9.850 0.510 ;
        RECT 12.940 0.490 13.310 0.570 ;
        RECT 12.940 0.480 13.970 0.490 ;
        RECT 15.850 0.480 16.160 0.640 ;
        RECT 12.940 0.310 16.320 0.480 ;
  END
END sky130_hilas_VinjDecode2to4

MACRO sky130_hilas_TA2Cell_1FG
  CLASS CORE ;
  FOREIGN sky130_hilas_TA2Cell_1FG ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.900 BY 23.320 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 17.820 10.230 18.300 10.240 ;
        RECT 17.820 9.990 18.710 10.230 ;
    END
  END VIN12
  PIN VIN11
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 17.870 13.750 18.710 13.950 ;
    END
  END VIN11
  PIN VIN21
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 32.610 12.090 32.930 12.330 ;
    END
  END VIN21
  PIN VIN22
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 32.530 14.760 32.840 15.000 ;
    END
  END VIN22
  PIN VPWR
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 35.760 14.880 36.040 15.030 ;
    END
    PORT
      LAYER met1 ;
        RECT 35.770 8.980 36.040 9.190 ;
    END
  END VPWR
  PIN VGND
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 35.530 16.460 35.850 16.540 ;
        RECT 34.540 16.280 35.850 16.460 ;
        RECT 34.540 16.110 35.720 16.280 ;
        RECT 34.590 15.960 34.910 16.110 ;
    END
    PORT
      LAYER met2 ;
        RECT 23.150 9.330 23.470 9.340 ;
        RECT 33.590 9.330 33.920 9.470 ;
        RECT 23.150 9.170 33.920 9.330 ;
        RECT 23.150 9.160 23.840 9.170 ;
        RECT 23.150 9.040 23.470 9.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.440 14.940 17.670 15.020 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.230 14.940 23.460 15.030 ;
    END
  END VGND
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 6.890 15.040 7.200 15.260 ;
        RECT 5.010 14.860 16.540 15.040 ;
        RECT 31.410 14.860 31.730 14.980 ;
        RECT 5.010 14.830 31.730 14.860 ;
        RECT 6.320 14.820 31.730 14.830 ;
        RECT 9.210 14.680 31.730 14.820 ;
        RECT 14.180 14.410 14.490 14.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.410 8.980 31.690 9.030 ;
    END
    PORT
      LAYER met1 ;
        RECT 9.210 14.980 9.490 15.030 ;
        RECT 9.210 14.700 9.530 14.980 ;
      LAYER via ;
        RECT 9.240 14.710 9.500 14.970 ;
    END
  END VINJ
  PIN OUTPUT1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 36.950 12.320 37.060 12.550 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 36.950 11.500 37.060 11.720 ;
    END
  END OUTPUT2
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 8.970 14.350 9.040 14.530 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 8.970 9.480 9.050 9.660 ;
    END
  END DRAIN2
  PIN COLSEL2
    PORT
      LAYER met1 ;
        RECT 9.740 14.970 9.930 15.030 ;
    END
  END COLSEL2
  PIN GATE2
    PORT
      LAYER met1 ;
        RECT 16.220 14.940 16.450 15.020 ;
    END
  END GATE2
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT 24.450 14.950 24.680 15.030 ;
    END
  END GATE1
  PIN COLSEL1
    PORT
      LAYER met1 ;
        RECT 30.970 14.950 31.160 15.030 ;
    END
    PORT
      LAYER met1 ;
        RECT 30.970 8.980 31.160 9.030 ;
    END
  END COLSEL1
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 19.730 14.870 21.170 15.030 ;
    END
  END VTUN
  OBS
      LAYER nwell ;
        RECT 0.290 22.980 2.020 23.320 ;
        RECT 38.880 22.980 40.610 23.320 ;
        RECT 0.290 21.420 2.040 22.980 ;
        RECT 0.310 19.790 2.040 21.420 ;
        RECT 38.860 21.420 40.610 22.980 ;
        RECT 38.860 19.790 40.590 21.420 ;
        RECT 0.250 19.400 3.550 19.790 ;
        RECT 0.010 19.360 3.550 19.400 ;
        RECT 0.000 17.710 3.550 19.360 ;
        RECT 37.350 19.400 40.650 19.790 ;
        RECT 37.350 19.360 40.890 19.400 ;
        RECT 32.590 19.310 35.890 19.320 ;
        RECT 34.930 19.280 35.120 19.310 ;
        RECT 0.250 16.620 3.550 17.710 ;
        RECT 37.350 17.710 40.900 19.360 ;
        RECT 0.250 14.780 3.550 15.970 ;
        RECT 8.970 15.020 10.950 15.030 ;
        RECT 0.000 13.130 3.550 14.780 ;
        RECT 15.390 14.670 15.950 17.090 ;
        RECT 24.950 14.670 25.510 17.090 ;
        RECT 37.350 16.620 40.650 17.710 ;
        RECT 37.760 15.970 39.040 16.620 ;
        RECT 31.930 15.020 33.400 15.030 ;
        RECT 35.780 14.850 37.060 15.030 ;
        RECT 37.350 14.780 40.650 15.970 ;
        RECT 8.970 14.350 9.040 14.530 ;
        RECT 0.010 13.090 3.550 13.130 ;
        RECT 0.250 12.800 3.550 13.090 ;
        RECT 37.350 13.130 40.900 14.780 ;
        RECT 37.350 13.090 40.890 13.130 ;
        RECT 37.350 12.800 40.650 13.090 ;
        RECT 8.970 9.480 9.050 9.660 ;
        RECT 37.760 9.470 39.040 12.310 ;
        RECT 35.780 8.980 37.060 9.170 ;
        RECT 31.930 7.550 32.380 7.780 ;
        RECT 30.590 7.420 32.450 7.490 ;
        RECT 34.220 3.050 36.080 6.040 ;
        RECT 34.220 0.000 36.080 2.990 ;
      LAYER li1 ;
        RECT 1.070 21.590 1.620 22.020 ;
        RECT 39.280 21.590 39.830 22.020 ;
        RECT 1.070 19.860 1.620 20.290 ;
        RECT 39.280 19.860 39.830 20.290 ;
        RECT 0.650 19.060 0.850 19.410 ;
        RECT 2.130 19.160 2.660 19.330 ;
        RECT 38.240 19.160 38.770 19.330 ;
        RECT 0.640 19.030 0.850 19.060 ;
        RECT 0.640 18.450 0.860 19.030 ;
        RECT 0.640 18.440 0.850 18.450 ;
        RECT 1.020 18.270 1.210 18.280 ;
        RECT 1.010 17.980 1.210 18.270 ;
        RECT 0.930 17.650 1.220 17.980 ;
        RECT 1.410 17.170 1.580 18.780 ;
        RECT 2.190 18.230 2.420 18.920 ;
        RECT 9.610 18.310 14.670 19.140 ;
        RECT 40.050 19.060 40.250 19.410 ;
        RECT 40.050 19.030 40.260 19.060 ;
        RECT 14.120 18.230 14.600 18.310 ;
        RECT 38.480 18.230 38.710 18.920 ;
        RECT 1.400 16.980 1.580 17.170 ;
        RECT 2.240 17.080 2.410 18.230 ;
        RECT 14.120 18.130 14.450 18.230 ;
        RECT 14.120 17.980 14.270 18.130 ;
        RECT 6.870 17.940 7.190 17.980 ;
        RECT 6.860 17.750 7.190 17.940 ;
        RECT 6.870 17.720 7.190 17.750 ;
        RECT 33.710 17.940 34.030 17.980 ;
        RECT 33.710 17.750 34.040 17.940 ;
        RECT 33.710 17.720 34.030 17.750 ;
        RECT 38.490 17.080 38.660 18.230 ;
        RECT 39.320 17.170 39.490 18.780 ;
        RECT 40.040 18.450 40.260 19.030 ;
        RECT 40.050 18.440 40.260 18.450 ;
        RECT 39.690 18.270 39.880 18.280 ;
        RECT 39.690 17.980 39.890 18.270 ;
        RECT 39.680 17.650 39.970 17.980 ;
        RECT 39.320 16.980 39.500 17.170 ;
        RECT 13.310 16.430 13.500 16.750 ;
        RECT 27.400 16.430 27.590 16.750 ;
        RECT 13.310 16.340 13.590 16.430 ;
        RECT 9.950 16.200 13.590 16.340 ;
        RECT 27.310 16.340 27.590 16.430 ;
        RECT 38.320 16.540 38.650 16.710 ;
        RECT 38.760 16.630 39.090 16.800 ;
        RECT 27.310 16.200 30.950 16.340 ;
        RECT 38.320 16.260 38.680 16.540 ;
        RECT 9.950 16.160 13.500 16.200 ;
        RECT 13.310 15.740 13.500 16.160 ;
        RECT 27.400 16.160 30.950 16.200 ;
        RECT 27.400 15.740 27.590 16.160 ;
        RECT 36.250 16.010 36.570 16.050 ;
        RECT 36.250 15.820 36.580 16.010 ;
        RECT 36.250 15.790 36.570 15.820 ;
        RECT 36.650 15.800 36.850 16.130 ;
        RECT 37.240 15.940 37.440 16.130 ;
        RECT 37.970 16.090 38.680 16.260 ;
        RECT 37.910 15.970 38.230 16.010 ;
        RECT 36.930 15.610 37.120 15.620 ;
        RECT 37.130 15.610 37.480 15.940 ;
        RECT 37.910 15.780 38.240 15.970 ;
        RECT 37.910 15.750 38.230 15.780 ;
        RECT 1.400 15.420 1.580 15.610 ;
        RECT 0.930 14.610 1.220 14.940 ;
        RECT 1.010 14.320 1.210 14.610 ;
        RECT 1.020 14.310 1.210 14.320 ;
        RECT 0.640 14.140 0.850 14.150 ;
        RECT 0.640 13.560 0.860 14.140 ;
        RECT 1.410 13.810 1.580 15.420 ;
        RECT 2.240 14.260 2.410 15.510 ;
        RECT 6.870 15.180 7.190 15.220 ;
        RECT 6.860 14.990 7.190 15.180 ;
        RECT 33.710 15.180 34.030 15.220 ;
        RECT 12.240 15.120 12.470 15.160 ;
        RECT 28.430 15.120 28.660 15.160 ;
        RECT 6.870 14.960 7.190 14.990 ;
        RECT 33.710 14.990 34.040 15.180 ;
        RECT 36.020 15.100 36.190 15.430 ;
        RECT 36.200 15.360 36.520 15.400 ;
        RECT 36.200 15.170 36.530 15.360 ;
        RECT 36.200 15.140 36.520 15.170 ;
        RECT 36.650 15.140 36.850 15.470 ;
        RECT 36.930 15.280 37.480 15.610 ;
        RECT 33.710 14.960 34.030 14.990 ;
        RECT 37.130 14.950 37.480 15.280 ;
        RECT 37.970 14.770 38.670 15.650 ;
        RECT 39.320 15.420 39.500 15.610 ;
        RECT 14.160 14.660 14.480 14.700 ;
        RECT 14.150 14.470 14.480 14.660 ;
        RECT 14.160 14.440 14.480 14.470 ;
        RECT 14.280 14.300 14.300 14.440 ;
        RECT 37.310 14.380 37.500 14.610 ;
        RECT 38.490 14.350 38.660 14.770 ;
        RECT 2.190 13.570 2.420 14.260 ;
        RECT 14.280 14.220 14.630 14.300 ;
        RECT 0.640 13.530 0.850 13.560 ;
        RECT 0.650 13.180 0.850 13.530 ;
        RECT 2.130 13.260 2.660 13.430 ;
        RECT 9.580 13.370 14.630 14.220 ;
        RECT 36.020 13.840 36.190 14.170 ;
        RECT 36.200 14.100 36.520 14.130 ;
        RECT 36.200 13.910 36.530 14.100 ;
        RECT 36.200 13.870 36.520 13.910 ;
        RECT 36.650 13.800 36.850 14.130 ;
        RECT 37.130 13.990 37.480 14.320 ;
        RECT 37.960 14.260 38.660 14.350 ;
        RECT 37.960 14.170 38.710 14.260 ;
        RECT 36.930 13.660 37.480 13.990 ;
        RECT 36.930 13.650 37.120 13.660 ;
        RECT 36.250 13.450 36.570 13.480 ;
        RECT 36.250 13.260 36.580 13.450 ;
        RECT 36.250 13.220 36.570 13.260 ;
        RECT 36.650 13.140 36.850 13.470 ;
        RECT 37.130 13.330 37.480 13.660 ;
        RECT 37.960 13.750 38.280 13.790 ;
        RECT 37.960 13.560 38.290 13.750 ;
        RECT 38.480 13.570 38.710 14.170 ;
        RECT 39.320 13.810 39.490 15.420 ;
        RECT 39.680 14.610 39.970 14.940 ;
        RECT 39.690 14.320 39.890 14.610 ;
        RECT 39.690 14.310 39.880 14.320 ;
        RECT 40.050 14.140 40.260 14.150 ;
        RECT 40.040 13.560 40.260 14.140 ;
        RECT 37.960 13.530 38.280 13.560 ;
        RECT 40.050 13.530 40.260 13.560 ;
        RECT 37.240 13.140 37.440 13.330 ;
        RECT 38.240 13.260 38.770 13.430 ;
        RECT 40.050 13.180 40.250 13.530 ;
        RECT 36.250 13.010 36.570 13.050 ;
        RECT 36.250 12.820 36.580 13.010 ;
        RECT 36.250 12.790 36.570 12.820 ;
        RECT 36.650 12.800 36.850 13.130 ;
        RECT 37.240 12.940 37.440 13.130 ;
        RECT 37.950 13.030 38.270 13.070 ;
        RECT 36.930 12.610 37.120 12.620 ;
        RECT 37.130 12.610 37.480 12.940 ;
        RECT 37.950 12.840 38.280 13.030 ;
        RECT 37.950 12.810 38.270 12.840 ;
        RECT 17.460 11.450 17.660 12.460 ;
        RECT 23.210 11.450 23.500 12.460 ;
        RECT 36.020 12.100 36.190 12.430 ;
        RECT 36.200 12.360 36.520 12.400 ;
        RECT 36.200 12.170 36.530 12.360 ;
        RECT 36.200 12.140 36.520 12.170 ;
        RECT 36.650 12.140 36.850 12.470 ;
        RECT 36.930 12.280 37.480 12.610 ;
        RECT 37.130 12.020 37.480 12.280 ;
        RECT 37.130 11.950 37.500 12.020 ;
        RECT 37.310 11.790 37.500 11.950 ;
        RECT 37.960 11.890 38.660 12.070 ;
        RECT 36.020 10.840 36.190 11.170 ;
        RECT 36.200 11.100 36.520 11.130 ;
        RECT 36.200 10.910 36.530 11.100 ;
        RECT 36.200 10.870 36.520 10.910 ;
        RECT 36.650 10.800 36.850 11.130 ;
        RECT 37.130 10.990 37.480 11.320 ;
        RECT 36.930 10.660 37.480 10.990 ;
        RECT 37.970 10.820 38.670 11.470 ;
        RECT 36.930 10.650 37.120 10.660 ;
        RECT 31.680 10.550 32.000 10.590 ;
        RECT 31.670 10.360 32.000 10.550 ;
        RECT 31.680 10.350 32.000 10.360 ;
        RECT 31.670 10.330 32.000 10.350 ;
        RECT 36.250 10.450 36.570 10.480 ;
        RECT 31.670 10.020 31.840 10.330 ;
        RECT 36.250 10.260 36.580 10.450 ;
        RECT 36.250 10.220 36.570 10.260 ;
        RECT 36.650 10.140 36.850 10.470 ;
        RECT 37.130 10.330 37.480 10.660 ;
        RECT 37.870 10.590 38.670 10.820 ;
        RECT 37.870 10.560 38.190 10.590 ;
        RECT 37.240 10.140 37.440 10.330 ;
        RECT 37.970 9.980 38.680 10.150 ;
        RECT 31.830 9.720 32.150 9.760 ;
        RECT 31.820 9.530 32.150 9.720 ;
        RECT 38.320 9.700 38.680 9.980 ;
        RECT 38.320 9.530 38.650 9.700 ;
        RECT 31.830 9.500 32.150 9.530 ;
        RECT 38.760 9.440 39.090 9.610 ;
        RECT 31.020 8.900 31.340 8.930 ;
        RECT 31.020 8.710 31.350 8.900 ;
        RECT 31.020 8.670 31.340 8.710 ;
        RECT 31.000 6.950 31.180 8.010 ;
        RECT 31.750 7.620 32.070 7.650 ;
        RECT 31.750 7.550 32.080 7.620 ;
        RECT 31.610 7.430 32.080 7.550 ;
        RECT 31.610 7.420 32.070 7.430 ;
        RECT 31.730 7.390 32.070 7.420 ;
        RECT 31.730 7.320 31.780 7.390 ;
        RECT 31.650 6.990 31.820 7.320 ;
        RECT 32.050 6.790 32.130 6.870 ;
        RECT 32.190 6.790 32.380 6.910 ;
        RECT 32.050 6.700 32.380 6.790 ;
        RECT 32.190 6.680 32.380 6.700 ;
        RECT 34.630 3.520 34.810 5.570 ;
        RECT 35.360 5.310 35.690 5.480 ;
        RECT 35.440 3.530 35.610 5.310 ;
        RECT 34.630 0.470 34.810 2.520 ;
        RECT 35.360 2.260 35.690 2.430 ;
        RECT 35.440 0.480 35.610 2.260 ;
      LAYER mcon ;
        RECT 1.350 21.670 1.620 21.940 ;
        RECT 39.280 21.670 39.550 21.940 ;
        RECT 1.350 19.940 1.620 20.210 ;
        RECT 39.280 19.940 39.550 20.210 ;
        RECT 2.480 19.160 2.660 19.330 ;
        RECT 0.670 18.860 0.840 19.030 ;
        RECT 1.020 18.020 1.200 18.210 ;
        RECT 2.220 18.710 2.390 18.880 ;
        RECT 2.220 18.260 2.390 18.430 ;
        RECT 14.220 18.170 14.390 18.340 ;
        RECT 38.510 18.710 38.680 18.880 ;
        RECT 40.060 18.860 40.230 19.030 ;
        RECT 38.510 18.260 38.680 18.430 ;
        RECT 6.960 17.760 7.130 17.930 ;
        RECT 33.770 17.760 33.940 17.930 ;
        RECT 39.700 18.020 39.880 18.210 ;
        RECT 13.410 16.230 13.580 16.400 ;
        RECT 27.320 16.230 27.490 16.400 ;
        RECT 36.310 15.830 36.480 16.000 ;
        RECT 37.970 15.790 38.140 15.960 ;
        RECT 1.020 14.380 1.200 14.570 ;
        RECT 6.960 15.000 7.130 15.170 ;
        RECT 33.770 15.000 33.940 15.170 ;
        RECT 36.260 15.180 36.430 15.350 ;
        RECT 37.250 15.440 37.420 15.610 ;
        RECT 14.250 14.480 14.420 14.650 ;
        RECT 37.320 14.410 37.490 14.580 ;
        RECT 2.220 14.060 2.390 14.230 ;
        RECT 0.670 13.560 0.840 13.730 ;
        RECT 2.220 13.610 2.390 13.780 ;
        RECT 2.480 13.260 2.660 13.430 ;
        RECT 36.260 13.920 36.430 14.090 ;
        RECT 37.250 13.660 37.420 13.830 ;
        RECT 38.510 14.060 38.680 14.230 ;
        RECT 36.310 13.270 36.480 13.440 ;
        RECT 39.700 14.380 39.880 14.570 ;
        RECT 38.020 13.570 38.190 13.740 ;
        RECT 38.510 13.610 38.680 13.780 ;
        RECT 40.060 13.560 40.230 13.730 ;
        RECT 36.310 12.830 36.480 13.000 ;
        RECT 38.010 12.850 38.180 13.020 ;
        RECT 17.470 12.220 17.640 12.390 ;
        RECT 17.480 11.500 17.650 11.670 ;
        RECT 23.260 12.220 23.430 12.390 ;
        RECT 36.260 12.180 36.430 12.350 ;
        RECT 37.250 12.440 37.420 12.610 ;
        RECT 37.320 11.820 37.490 11.990 ;
        RECT 23.260 11.500 23.430 11.670 ;
        RECT 36.260 10.920 36.430 11.090 ;
        RECT 37.250 10.660 37.420 10.830 ;
        RECT 31.770 10.370 31.940 10.540 ;
        RECT 36.310 10.270 36.480 10.440 ;
        RECT 37.930 10.600 38.100 10.770 ;
        RECT 31.920 9.540 32.090 9.710 ;
        RECT 31.080 8.720 31.250 8.890 ;
        RECT 31.810 7.440 31.980 7.610 ;
        RECT 32.200 6.710 32.370 6.880 ;
      LAYER met1 ;
        RECT 0.610 19.090 0.770 19.730 ;
        RECT 0.610 18.540 0.880 19.090 ;
        RECT 0.600 18.490 0.880 18.540 ;
        RECT 0.600 18.400 0.770 18.490 ;
        RECT 0.610 16.710 0.770 18.400 ;
        RECT 1.020 18.280 1.210 19.730 ;
        RECT 1.290 19.400 1.680 22.990 ;
        RECT 39.220 19.400 39.610 22.990 ;
        RECT 2.420 18.970 2.730 19.360 ;
        RECT 0.990 18.250 1.210 18.280 ;
        RECT 2.180 18.920 2.730 18.970 ;
        RECT 0.980 17.980 1.230 18.250 ;
        RECT 2.180 18.180 2.440 18.920 ;
        RECT 0.980 17.970 1.220 17.980 ;
        RECT 0.990 17.730 1.220 17.970 ;
        RECT 1.020 16.710 1.180 17.730 ;
        RECT 1.370 16.920 1.610 17.300 ;
        RECT 0.610 14.190 0.770 15.880 ;
        RECT 1.020 14.860 1.180 15.880 ;
        RECT 1.370 15.290 1.610 15.670 ;
        RECT 0.990 14.620 1.220 14.860 ;
        RECT 0.980 14.610 1.220 14.620 ;
        RECT 0.980 14.340 1.230 14.610 ;
        RECT 0.990 14.310 1.210 14.340 ;
        RECT 0.600 14.100 0.770 14.190 ;
        RECT 0.600 14.050 0.880 14.100 ;
        RECT 0.610 13.500 0.880 14.050 ;
        RECT 0.610 12.860 0.770 13.500 ;
        RECT 1.020 12.860 1.210 14.310 ;
        RECT 2.180 13.670 2.440 14.310 ;
        RECT 2.180 13.520 2.730 13.670 ;
        RECT 2.420 13.230 2.730 13.520 ;
        RECT 5.250 13.270 5.530 19.320 ;
        RECT 5.780 19.260 5.970 19.320 ;
        RECT 6.880 17.690 7.200 18.010 ;
        RECT 6.020 16.530 6.280 16.850 ;
        RECT 6.020 15.930 6.280 16.250 ;
        RECT 6.880 14.930 7.200 15.250 ;
        RECT 5.780 13.270 5.970 13.330 ;
        RECT 12.260 13.270 12.490 19.320 ;
        RECT 13.480 18.350 13.710 19.320 ;
        RECT 13.470 18.100 13.710 18.350 ;
        RECT 14.140 18.100 14.460 18.420 ;
        RECT 13.480 16.460 13.710 18.100 ;
        RECT 13.380 16.170 13.710 16.460 ;
        RECT 13.480 13.270 13.710 16.170 ;
        RECT 14.170 14.410 14.490 14.730 ;
        RECT 15.770 13.280 16.190 19.320 ;
        RECT 24.710 13.270 25.130 19.320 ;
        RECT 27.190 16.460 27.420 19.320 ;
        RECT 27.190 16.170 27.520 16.460 ;
        RECT 27.190 13.270 27.420 16.170 ;
        RECT 28.410 13.270 28.640 19.320 ;
        RECT 34.930 19.280 35.120 19.320 ;
        RECT 33.700 17.690 34.020 18.010 ;
        RECT 34.620 16.530 34.880 16.850 ;
        RECT 35.370 16.570 35.650 19.320 ;
        RECT 38.170 18.970 38.480 19.360 ;
        RECT 38.170 18.920 38.720 18.970 ;
        RECT 38.460 18.180 38.720 18.920 ;
        RECT 39.690 18.280 39.880 19.730 ;
        RECT 40.130 19.090 40.290 19.730 ;
        RECT 40.020 18.540 40.290 19.090 ;
        RECT 40.020 18.490 40.300 18.540 ;
        RECT 40.130 18.400 40.300 18.490 ;
        RECT 39.690 18.250 39.910 18.280 ;
        RECT 39.670 17.980 39.920 18.250 ;
        RECT 39.680 17.970 39.920 17.980 ;
        RECT 39.680 17.730 39.910 17.970 ;
        RECT 39.290 16.920 39.530 17.300 ;
        RECT 39.720 16.710 39.880 17.730 ;
        RECT 40.130 16.710 40.290 18.400 ;
        RECT 35.370 16.250 35.820 16.570 ;
        RECT 34.620 15.930 34.880 16.250 ;
        RECT 31.410 14.980 31.690 15.030 ;
        RECT 31.410 14.680 31.730 14.980 ;
        RECT 33.700 14.930 34.020 15.250 ;
        RECT 35.370 15.030 35.650 16.250 ;
        RECT 36.240 16.000 36.560 16.080 ;
        RECT 36.240 15.760 36.810 16.000 ;
        RECT 36.470 15.430 36.810 15.760 ;
        RECT 36.190 15.110 36.810 15.430 ;
        RECT 35.100 14.890 35.650 15.030 ;
        RECT 34.930 13.270 35.120 13.320 ;
        RECT 35.370 13.270 35.650 14.890 ;
        RECT 36.470 14.160 36.810 15.110 ;
        RECT 36.190 13.840 36.810 14.160 ;
        RECT 36.470 13.510 36.810 13.840 ;
        RECT 36.240 13.190 36.810 13.510 ;
        RECT 36.470 13.080 36.810 13.190 ;
        RECT 36.240 12.760 36.810 13.080 ;
        RECT 36.470 12.430 36.810 12.760 ;
        RECT 17.470 12.210 17.640 12.390 ;
        RECT 23.260 12.210 23.430 12.390 ;
        RECT 36.190 12.110 36.810 12.430 ;
        RECT 17.450 11.620 17.770 11.920 ;
        RECT 17.450 11.510 17.690 11.620 ;
        RECT 23.150 11.550 23.470 11.870 ;
        RECT 17.480 11.500 17.650 11.510 ;
        RECT 17.670 11.450 17.690 11.510 ;
        RECT 23.260 11.500 23.430 11.550 ;
        RECT 36.470 11.160 36.810 12.110 ;
        RECT 36.190 10.840 36.810 11.160 ;
        RECT 31.690 10.300 32.010 10.620 ;
        RECT 36.470 10.510 36.810 10.840 ;
        RECT 36.240 10.280 36.810 10.510 ;
        RECT 37.140 15.670 37.410 15.990 ;
        RECT 37.900 15.720 38.220 16.040 ;
        RECT 37.140 15.380 37.450 15.670 ;
        RECT 37.140 14.640 37.410 15.380 ;
        RECT 39.290 15.290 39.530 15.670 ;
        RECT 39.720 14.860 39.880 15.880 ;
        RECT 37.140 14.350 37.520 14.640 ;
        RECT 39.680 14.620 39.910 14.860 ;
        RECT 39.680 14.610 39.920 14.620 ;
        RECT 37.140 13.890 37.410 14.350 ;
        RECT 39.670 14.340 39.920 14.610 ;
        RECT 39.690 14.310 39.910 14.340 ;
        RECT 37.140 13.600 37.450 13.890 ;
        RECT 37.950 13.670 38.270 13.820 ;
        RECT 38.460 13.670 38.720 14.310 ;
        RECT 37.140 12.670 37.410 13.600 ;
        RECT 37.950 13.520 38.720 13.670 ;
        RECT 37.950 13.500 38.480 13.520 ;
        RECT 38.170 13.230 38.480 13.500 ;
        RECT 37.940 12.780 38.260 13.100 ;
        RECT 39.690 12.860 39.880 14.310 ;
        RECT 40.130 14.190 40.290 15.880 ;
        RECT 40.130 14.100 40.300 14.190 ;
        RECT 40.020 14.050 40.300 14.100 ;
        RECT 40.020 13.500 40.290 14.050 ;
        RECT 40.130 12.860 40.290 13.500 ;
        RECT 37.140 12.380 37.450 12.670 ;
        RECT 37.140 12.050 37.410 12.380 ;
        RECT 37.140 11.760 37.520 12.050 ;
        RECT 37.140 10.890 37.410 11.760 ;
        RECT 37.140 10.600 37.450 10.890 ;
        RECT 37.140 10.290 37.410 10.600 ;
        RECT 37.860 10.530 38.180 10.850 ;
        RECT 36.240 10.190 36.560 10.280 ;
        RECT 31.840 9.470 32.160 9.790 ;
        RECT 23.150 9.040 23.470 9.340 ;
        RECT 33.590 9.180 33.920 9.470 ;
        RECT 33.580 9.150 34.000 9.180 ;
        RECT 34.600 9.170 35.100 9.180 ;
        RECT 34.600 9.150 35.440 9.170 ;
        RECT 33.580 9.040 35.440 9.150 ;
        RECT 33.860 9.010 34.760 9.040 ;
        RECT 35.100 8.980 35.440 9.040 ;
        RECT 31.010 8.640 31.330 8.960 ;
        RECT 32.090 8.530 32.300 8.740 ;
        RECT 32.090 8.210 32.420 8.530 ;
        RECT 31.740 7.360 32.060 7.680 ;
        RECT 32.090 6.970 32.300 8.210 ;
        RECT 32.170 6.650 32.400 6.940 ;
      LAYER via ;
        RECT 2.440 18.950 2.700 19.210 ;
        RECT 2.440 13.380 2.700 13.640 ;
        RECT 6.910 17.720 7.170 17.980 ;
        RECT 6.020 16.560 6.280 16.820 ;
        RECT 6.020 15.960 6.280 16.220 ;
        RECT 6.910 14.960 7.170 15.220 ;
        RECT 14.170 18.130 14.430 18.390 ;
        RECT 14.200 14.440 14.460 14.700 ;
        RECT 33.730 17.720 33.990 17.980 ;
        RECT 34.620 16.560 34.880 16.820 ;
        RECT 38.200 18.950 38.460 19.210 ;
        RECT 35.560 16.280 35.820 16.540 ;
        RECT 34.620 15.960 34.880 16.220 ;
        RECT 31.440 14.700 31.700 14.960 ;
        RECT 33.730 14.960 33.990 15.220 ;
        RECT 36.270 15.790 36.530 16.050 ;
        RECT 36.220 15.140 36.480 15.400 ;
        RECT 36.220 13.870 36.480 14.130 ;
        RECT 36.270 13.220 36.530 13.480 ;
        RECT 36.270 12.790 36.530 13.050 ;
        RECT 36.220 12.140 36.480 12.400 ;
        RECT 17.480 11.640 17.740 11.900 ;
        RECT 23.180 11.580 23.440 11.840 ;
        RECT 36.220 10.870 36.480 11.130 ;
        RECT 31.720 10.330 31.980 10.590 ;
        RECT 36.270 10.220 36.530 10.480 ;
        RECT 37.930 15.750 38.190 16.010 ;
        RECT 37.980 13.640 38.240 13.790 ;
        RECT 37.980 13.530 38.460 13.640 ;
        RECT 38.200 13.380 38.460 13.530 ;
        RECT 37.970 12.810 38.230 13.070 ;
        RECT 37.890 10.560 38.150 10.820 ;
        RECT 31.870 9.500 32.130 9.760 ;
        RECT 23.180 9.060 23.440 9.320 ;
        RECT 33.620 9.190 33.890 9.450 ;
        RECT 31.040 8.670 31.300 8.930 ;
        RECT 32.160 8.240 32.420 8.500 ;
        RECT 31.770 7.390 32.030 7.650 ;
      LAYER met2 ;
        RECT 2.420 19.240 2.730 19.250 ;
        RECT 0.250 19.060 2.730 19.240 ;
        RECT 2.420 18.920 2.730 19.060 ;
        RECT 38.170 19.240 38.480 19.250 ;
        RECT 38.170 19.060 40.650 19.240 ;
        RECT 38.170 18.920 38.480 19.060 ;
        RECT 7.420 18.640 16.540 18.820 ;
        RECT 24.360 18.640 33.480 18.820 ;
        RECT 14.150 18.230 14.460 18.430 ;
        RECT 14.150 18.220 14.750 18.230 ;
        RECT 14.150 18.100 16.540 18.220 ;
        RECT 14.290 18.060 16.540 18.100 ;
        RECT 14.600 18.040 16.540 18.060 ;
        RECT 6.890 17.800 7.200 18.020 ;
        RECT 5.010 17.790 7.200 17.800 ;
        RECT 33.700 17.800 34.010 18.020 ;
        RECT 5.010 17.580 16.540 17.790 ;
        RECT 33.700 17.690 35.890 17.800 ;
        RECT 33.860 17.580 35.890 17.690 ;
        RECT 6.320 17.570 16.540 17.580 ;
        RECT 5.990 16.600 16.540 16.820 ;
        RECT 5.990 16.560 6.310 16.600 ;
        RECT 34.590 16.560 34.910 16.820 ;
        RECT 6.100 16.220 6.360 16.460 ;
        RECT 5.990 16.110 6.360 16.220 ;
        RECT 5.990 15.960 6.310 16.110 ;
        RECT 36.240 15.800 36.550 16.090 ;
        RECT 37.900 15.800 38.210 16.050 ;
        RECT 35.520 15.720 38.210 15.800 ;
        RECT 35.520 15.570 38.060 15.720 ;
        RECT 33.700 15.040 34.010 15.260 ;
        RECT 35.750 15.040 36.080 15.210 ;
        RECT 36.190 15.110 36.500 15.440 ;
        RECT 33.700 15.000 36.080 15.040 ;
        RECT 33.700 14.930 35.890 15.000 ;
        RECT 33.850 14.830 35.890 14.930 ;
        RECT 14.590 14.300 16.540 14.510 ;
        RECT 33.640 14.130 33.860 14.150 ;
        RECT 7.320 13.940 7.480 13.960 ;
        RECT 33.420 13.940 33.580 13.960 ;
        RECT 7.320 13.890 16.540 13.940 ;
        RECT 7.440 13.790 16.540 13.890 ;
        RECT 24.360 13.890 33.580 13.940 ;
        RECT 24.360 13.790 33.460 13.890 ;
        RECT 33.590 13.790 33.860 14.130 ;
        RECT 35.750 14.060 36.080 14.270 ;
        RECT 36.190 13.830 36.500 14.160 ;
        RECT 37.950 13.670 38.260 13.830 ;
        RECT 2.420 13.530 2.730 13.670 ;
        RECT 37.950 13.660 38.480 13.670 ;
        RECT 0.250 13.350 2.730 13.530 ;
        RECT 35.780 13.530 38.480 13.660 ;
        RECT 2.420 13.340 2.730 13.350 ;
        RECT 18.320 13.280 28.460 13.500 ;
        RECT 31.850 13.290 32.200 13.510 ;
        RECT 35.780 13.430 40.650 13.530 ;
        RECT 18.270 12.310 27.280 12.530 ;
        RECT 17.450 11.870 17.770 11.920 ;
        RECT 17.450 11.620 23.470 11.870 ;
        RECT 23.150 11.550 23.470 11.620 ;
        RECT 18.320 10.530 23.980 10.750 ;
        RECT 23.760 10.200 23.980 10.530 ;
        RECT 27.060 10.700 27.280 12.310 ;
        RECT 28.240 12.080 28.460 13.280 ;
        RECT 33.660 13.220 33.860 13.230 ;
        RECT 33.660 12.890 33.880 13.220 ;
        RECT 36.240 13.180 36.550 13.430 ;
        RECT 38.170 13.350 40.650 13.430 ;
        RECT 38.170 13.340 38.480 13.350 ;
        RECT 33.680 12.880 33.880 12.890 ;
        RECT 36.240 12.830 36.550 13.090 ;
        RECT 37.940 12.830 38.250 13.110 ;
        RECT 35.520 12.610 38.430 12.830 ;
        RECT 28.210 12.040 28.460 12.080 ;
        RECT 28.210 11.400 28.470 12.040 ;
        RECT 35.750 12.000 36.080 12.210 ;
        RECT 36.190 12.110 36.500 12.440 ;
        RECT 28.210 11.190 32.340 11.400 ;
        RECT 32.130 11.050 32.340 11.190 ;
        RECT 35.750 11.060 36.080 11.270 ;
        RECT 32.130 10.840 34.150 11.050 ;
        RECT 36.190 10.830 36.500 11.160 ;
        RECT 27.060 10.480 29.910 10.700 ;
        RECT 37.860 10.670 38.170 10.860 ;
        RECT 31.700 10.470 32.010 10.630 ;
        RECT 31.270 10.250 32.150 10.470 ;
        RECT 35.510 10.440 38.220 10.670 ;
        RECT 28.130 10.200 34.150 10.250 ;
        RECT 23.760 10.040 34.150 10.200 ;
        RECT 36.240 10.180 36.550 10.440 ;
        RECT 23.760 9.980 28.520 10.040 ;
        RECT 31.850 9.610 32.160 9.800 ;
        RECT 31.810 9.360 32.360 9.610 ;
        RECT 31.010 8.630 31.320 8.960 ;
        RECT 31.990 8.330 32.460 8.580 ;
        RECT 32.130 8.240 32.450 8.330 ;
        RECT 31.510 7.780 31.940 7.790 ;
        RECT 31.510 7.550 32.380 7.780 ;
        RECT 31.740 7.350 32.050 7.550 ;
  END
END sky130_hilas_TA2Cell_1FG

MACRO sky130_hilas_swc4x1cellOverlap
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x1cellOverlap ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 10.510 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 14.520 9.060 16.250 10.510 ;
        RECT 7.740 6.980 10.460 7.510 ;
        RECT 14.490 7.220 16.250 9.060 ;
        RECT 7.740 5.070 12.970 6.980 ;
        RECT 7.740 4.910 10.460 5.070 ;
        RECT 7.740 4.420 12.970 4.910 ;
        RECT 14.520 4.460 16.250 7.220 ;
        RECT 7.730 2.060 12.970 4.420 ;
        RECT 7.730 1.910 10.450 2.060 ;
        RECT 7.730 0.920 12.970 1.910 ;
        RECT 10.410 0.000 12.970 0.920 ;
      LAYER li1 ;
        RECT 14.910 7.670 15.460 8.100 ;
        RECT 8.140 5.940 10.090 7.110 ;
        RECT 10.650 6.630 10.970 6.670 ;
        RECT 10.650 6.510 10.980 6.630 ;
        RECT 10.650 6.410 11.090 6.510 ;
        RECT 10.750 6.340 11.090 6.410 ;
        RECT 12.370 6.240 12.570 6.590 ;
        RECT 10.650 6.080 10.970 6.120 ;
        RECT 10.650 5.890 10.980 6.080 ;
        RECT 10.650 5.860 11.090 5.890 ;
        RECT 10.750 5.720 11.090 5.860 ;
        RECT 11.640 5.620 11.840 6.220 ;
        RECT 12.370 6.210 12.580 6.240 ;
        RECT 12.360 5.620 12.580 6.210 ;
        RECT 8.140 4.410 10.090 5.580 ;
        RECT 10.750 4.120 11.090 4.260 ;
        RECT 10.650 4.090 11.090 4.120 ;
        RECT 8.130 2.850 10.080 4.020 ;
        RECT 10.650 3.900 10.980 4.090 ;
        RECT 10.650 3.860 10.970 3.900 ;
        RECT 11.640 3.760 11.840 4.360 ;
        RECT 12.360 3.770 12.580 4.360 ;
        RECT 12.370 3.740 12.580 3.770 ;
        RECT 10.650 3.640 10.970 3.660 ;
        RECT 10.650 3.330 11.090 3.640 ;
        RECT 10.650 3.310 10.970 3.330 ;
        RECT 12.370 3.230 12.570 3.740 ;
        RECT 10.650 3.070 10.970 3.110 ;
        RECT 10.650 2.880 10.980 3.070 ;
        RECT 10.650 2.850 11.090 2.880 ;
        RECT 10.750 2.710 11.090 2.850 ;
        RECT 11.640 2.610 11.840 3.210 ;
        RECT 12.370 3.200 12.580 3.230 ;
        RECT 12.360 2.610 12.580 3.200 ;
        RECT 8.130 1.310 10.080 2.480 ;
        RECT 10.750 1.120 11.090 1.260 ;
        RECT 10.650 1.090 11.090 1.120 ;
        RECT 10.650 0.900 10.980 1.090 ;
        RECT 10.650 0.860 10.970 0.900 ;
        RECT 11.640 0.760 11.840 1.360 ;
        RECT 12.360 0.770 12.580 1.360 ;
        RECT 12.370 0.740 12.580 0.770 ;
        RECT 10.750 0.570 11.090 0.640 ;
        RECT 10.650 0.470 11.090 0.570 ;
        RECT 10.650 0.350 10.980 0.470 ;
        RECT 12.370 0.390 12.570 0.740 ;
        RECT 10.650 0.310 10.970 0.350 ;
      LAYER mcon ;
        RECT 14.910 7.750 15.180 8.020 ;
        RECT 8.620 6.770 8.790 6.940 ;
        RECT 8.620 6.430 8.790 6.600 ;
        RECT 10.710 6.450 10.880 6.620 ;
        RECT 8.620 6.090 8.790 6.260 ;
        RECT 10.710 5.900 10.880 6.070 ;
        RECT 11.650 6.010 11.820 6.180 ;
        RECT 12.380 6.040 12.550 6.210 ;
        RECT 8.620 5.240 8.790 5.410 ;
        RECT 8.620 4.900 8.790 5.070 ;
        RECT 8.620 4.560 8.790 4.730 ;
        RECT 10.710 3.910 10.880 4.080 ;
        RECT 8.610 3.680 8.780 3.850 ;
        RECT 11.650 3.800 11.820 3.970 ;
        RECT 12.380 3.770 12.550 3.940 ;
        RECT 8.610 3.340 8.780 3.510 ;
        RECT 9.130 3.400 9.310 3.570 ;
        RECT 10.710 3.360 10.880 3.610 ;
        RECT 8.610 3.000 8.780 3.170 ;
        RECT 10.710 2.890 10.880 3.060 ;
        RECT 11.650 3.000 11.820 3.170 ;
        RECT 12.380 3.030 12.550 3.200 ;
        RECT 8.610 2.140 8.780 2.310 ;
        RECT 8.610 1.800 8.780 1.970 ;
        RECT 8.610 1.460 8.780 1.630 ;
        RECT 10.710 0.910 10.880 1.080 ;
        RECT 11.650 0.800 11.820 0.970 ;
        RECT 12.380 0.770 12.550 0.940 ;
        RECT 10.710 0.360 10.880 0.530 ;
      LAYER met1 ;
        RECT 14.850 7.210 15.240 9.070 ;
        RECT 8.580 6.520 8.840 7.000 ;
        RECT 0.360 0.460 0.760 6.450 ;
        RECT 8.570 6.000 8.840 6.520 ;
        RECT 10.640 6.380 10.960 6.700 ;
        RECT 11.640 6.240 11.800 6.970 ;
        RECT 11.640 6.220 11.840 6.240 ;
        RECT 8.570 5.550 8.830 6.000 ;
        RECT 10.640 5.830 10.960 6.150 ;
        RECT 11.620 5.980 11.850 6.220 ;
        RECT 11.640 5.930 11.850 5.980 ;
        RECT 12.010 5.930 12.200 6.920 ;
        RECT 12.450 6.270 12.610 6.970 ;
        RECT 8.580 4.990 8.840 5.470 ;
        RECT 11.640 5.070 11.800 5.930 ;
        RECT 12.030 5.810 12.200 5.930 ;
        RECT 12.040 5.070 12.200 5.810 ;
        RECT 12.340 5.720 12.610 6.270 ;
        RECT 12.340 5.670 12.620 5.720 ;
        RECT 12.450 5.580 12.620 5.670 ;
        RECT 12.450 5.070 12.610 5.580 ;
        RECT 8.570 4.470 8.840 4.990 ;
        RECT 8.570 4.020 8.830 4.470 ;
        RECT 8.570 3.430 8.830 3.910 ;
        RECT 10.640 3.830 10.960 4.150 ;
        RECT 11.640 4.050 11.800 4.910 ;
        RECT 12.040 4.170 12.200 4.910 ;
        RECT 12.450 4.400 12.610 4.910 ;
        RECT 12.450 4.310 12.620 4.400 ;
        RECT 12.030 4.050 12.200 4.170 ;
        RECT 11.640 4.000 11.850 4.050 ;
        RECT 11.620 3.760 11.850 4.000 ;
        RECT 11.640 3.740 11.840 3.760 ;
        RECT 9.180 3.600 9.310 3.620 ;
        RECT 8.560 2.910 8.830 3.430 ;
        RECT 9.100 3.370 9.340 3.600 ;
        RECT 9.200 3.330 9.310 3.370 ;
        RECT 10.640 3.280 10.960 3.690 ;
        RECT 11.640 3.230 11.800 3.740 ;
        RECT 11.640 3.210 11.840 3.230 ;
        RECT 8.560 2.460 8.820 2.910 ;
        RECT 10.640 2.820 10.960 3.140 ;
        RECT 11.620 2.970 11.850 3.210 ;
        RECT 11.640 2.920 11.850 2.970 ;
        RECT 12.010 2.920 12.200 4.050 ;
        RECT 12.340 4.260 12.620 4.310 ;
        RECT 12.340 3.710 12.610 4.260 ;
        RECT 12.450 3.260 12.610 3.710 ;
        RECT 8.570 1.890 8.830 2.370 ;
        RECT 11.640 2.060 11.800 2.920 ;
        RECT 12.030 2.800 12.200 2.920 ;
        RECT 12.040 2.060 12.200 2.800 ;
        RECT 12.340 2.710 12.610 3.260 ;
        RECT 12.340 2.660 12.620 2.710 ;
        RECT 12.450 2.570 12.620 2.660 ;
        RECT 12.450 2.060 12.610 2.570 ;
        RECT 8.560 1.370 8.830 1.890 ;
        RECT 8.560 0.920 8.820 1.370 ;
        RECT 10.640 0.830 10.960 1.150 ;
        RECT 11.640 1.050 11.800 1.910 ;
        RECT 12.040 1.170 12.200 1.910 ;
        RECT 12.450 1.400 12.610 1.910 ;
        RECT 12.450 1.310 12.620 1.400 ;
        RECT 12.030 1.050 12.200 1.170 ;
        RECT 11.640 1.000 11.850 1.050 ;
        RECT 11.620 0.760 11.850 1.000 ;
        RECT 11.640 0.740 11.840 0.760 ;
        RECT 10.640 0.280 10.960 0.600 ;
        RECT 11.640 0.010 11.800 0.740 ;
        RECT 12.010 0.060 12.200 1.050 ;
        RECT 12.340 1.260 12.620 1.310 ;
        RECT 12.340 0.710 12.610 1.260 ;
        RECT 12.450 0.010 12.610 0.710 ;
      LAYER via ;
        RECT 10.670 6.410 10.930 6.670 ;
        RECT 10.670 5.860 10.930 6.120 ;
        RECT 10.670 3.860 10.930 4.120 ;
        RECT 10.670 3.310 10.930 3.660 ;
        RECT 10.670 2.850 10.930 3.110 ;
        RECT 10.670 0.860 10.930 1.120 ;
        RECT 10.670 0.310 10.930 0.570 ;
      LAYER met2 ;
        RECT 10.640 6.420 10.950 6.710 ;
        RECT 10.640 6.380 12.970 6.420 ;
        RECT 10.790 6.240 12.970 6.380 ;
        RECT 0.000 5.940 7.610 6.010 ;
        RECT 10.640 5.990 10.950 6.160 ;
        RECT 0.000 5.830 7.640 5.940 ;
        RECT 10.410 5.810 10.500 5.990 ;
        RECT 10.640 5.830 12.970 5.990 ;
        RECT 10.800 5.810 12.970 5.830 ;
        RECT 0.000 5.400 9.740 5.580 ;
        RECT 0.000 4.520 7.610 4.580 ;
        RECT 0.000 4.400 7.640 4.520 ;
        RECT 0.000 4.080 7.600 4.150 ;
        RECT 0.000 3.970 7.640 4.080 ;
        RECT 10.410 3.990 10.500 4.170 ;
        RECT 10.800 4.150 12.970 4.170 ;
        RECT 10.640 3.990 12.970 4.150 ;
        RECT 10.640 3.820 10.950 3.990 ;
        RECT 10.790 3.700 12.970 3.740 ;
        RECT 10.640 3.560 12.970 3.700 ;
        RECT 10.640 3.410 10.950 3.560 ;
        RECT 10.640 3.270 12.970 3.410 ;
        RECT 10.790 3.230 12.970 3.270 ;
        RECT 0.020 2.820 7.640 2.990 ;
        RECT 10.640 2.980 10.950 3.150 ;
        RECT 10.410 2.800 10.500 2.980 ;
        RECT 10.640 2.820 12.970 2.980 ;
        RECT 10.800 2.800 12.970 2.820 ;
        RECT 0.020 2.400 7.640 2.570 ;
        RECT 0.020 1.420 7.640 1.590 ;
        RECT 0.800 1.330 2.340 1.420 ;
        RECT 0.020 0.980 7.640 1.150 ;
        RECT 10.410 0.990 10.500 1.170 ;
        RECT 10.800 1.150 12.970 1.170 ;
        RECT 10.640 0.990 12.970 1.150 ;
        RECT 10.640 0.820 10.950 0.990 ;
        RECT 10.790 0.600 12.970 0.740 ;
        RECT 10.640 0.560 12.970 0.600 ;
        RECT 10.640 0.270 10.950 0.560 ;
  END
END sky130_hilas_swc4x1cellOverlap

MACRO sky130_hilas_capacitorSize02
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize02 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.610 BY 7.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 7.660 2.390 7.970 2.670 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.020 2.370 0.290 2.650 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 0.000 4.850 7.970 5.030 ;
        RECT 0.000 4.420 7.970 4.600 ;
        RECT 0.030 3.420 7.970 3.600 ;
        RECT 0.030 3.090 7.970 3.170 ;
        RECT 0.030 2.990 8.090 3.090 ;
        RECT 0.600 2.670 0.970 2.990 ;
        RECT 7.720 2.690 8.090 2.990 ;
        RECT 0.030 1.840 7.970 2.010 ;
        RECT 0.030 1.420 7.970 1.590 ;
        RECT 0.030 0.440 7.970 0.610 ;
        RECT 0.030 0.000 7.970 0.170 ;
      LAYER via2 ;
        RECT 0.650 2.730 0.930 3.010 ;
        RECT 7.770 2.750 8.050 3.030 ;
      LAYER met3 ;
        RECT 5.380 7.840 7.690 7.870 ;
        RECT 0.380 2.470 1.170 3.220 ;
        RECT 5.380 2.060 9.610 7.840 ;
        RECT 7.660 2.040 9.610 2.060 ;
      LAYER via3 ;
        RECT 0.570 2.620 1.000 3.100 ;
        RECT 7.690 2.640 8.120 3.120 ;
      LAYER met4 ;
        RECT 0.470 2.770 1.130 3.190 ;
        RECT 5.760 3.140 8.770 3.610 ;
        RECT 1.160 2.770 2.170 2.780 ;
        RECT 0.450 2.270 3.800 2.770 ;
        RECT 7.590 2.550 8.250 3.140 ;
        RECT 0.450 2.260 1.520 2.270 ;
        RECT 3.160 1.150 3.790 2.270 ;
        RECT 3.160 0.850 5.310 1.150 ;
        RECT 3.490 0.840 5.310 0.850 ;
  END
END sky130_hilas_capacitorSize02

MACRO sky130_hilas_nFETLarge
  CLASS CORE ;
  FOREIGN sky130_hilas_nFETLarge ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.570 BY 6.030 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    USE ANALOG ;
    ANTENNAGATEAREA 2.642500 ;
    PORT
      LAYER met2 ;
        RECT 0.430 0.820 0.740 0.950 ;
        RECT 0.000 0.620 0.740 0.820 ;
        RECT 0.000 0.480 0.600 0.620 ;
        RECT 0.000 0.150 0.750 0.480 ;
        RECT 0.000 0.000 0.600 0.150 ;
    END
  END GATE
  PIN SOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 1.343400 ;
    PORT
      LAYER met2 ;
        RECT 1.010 5.600 1.320 5.740 ;
        RECT 2.100 5.600 2.410 5.740 ;
        RECT 3.200 5.600 3.510 5.730 ;
        RECT 0.330 5.590 3.510 5.600 ;
        RECT 0.240 5.400 3.510 5.590 ;
        RECT 0.240 5.260 3.390 5.400 ;
        RECT 0.240 2.810 0.560 5.260 ;
        RECT 1.000 2.810 1.310 2.960 ;
        RECT 2.100 2.810 2.410 2.960 ;
        RECT 3.200 2.810 3.510 2.960 ;
        RECT 0.240 2.630 3.510 2.810 ;
        RECT 0.240 2.480 3.400 2.630 ;
        RECT 0.240 1.440 0.560 2.480 ;
        RECT 1.000 1.440 1.310 1.590 ;
        RECT 2.100 1.440 2.410 1.590 ;
        RECT 3.200 1.440 3.510 1.590 ;
        RECT 0.240 1.260 3.510 1.440 ;
        RECT 0.240 1.120 3.400 1.260 ;
    END
  END SOURCE
  PIN DRAIN
    USE ANALOG ;
    ANTENNADIFFAREA 2.723900 ;
    PORT
      LAYER met2 ;
        RECT 1.560 4.880 1.870 5.060 ;
        RECT 2.650 4.880 2.960 5.040 ;
        RECT 3.760 4.880 4.070 5.030 ;
        RECT 1.430 4.580 4.370 4.880 ;
        RECT 3.620 4.540 4.370 4.580 ;
        RECT 3.990 4.410 4.370 4.540 ;
        RECT 4.020 3.690 4.370 4.410 ;
        RECT 1.560 3.540 1.870 3.690 ;
        RECT 2.650 3.540 2.960 3.690 ;
        RECT 3.750 3.540 4.370 3.690 ;
        RECT 1.420 3.210 4.370 3.540 ;
        RECT 4.020 0.920 4.370 3.210 ;
        RECT 1.560 0.770 1.870 0.910 ;
        RECT 2.650 0.770 2.960 0.910 ;
        RECT 3.750 0.770 4.370 0.920 ;
        RECT 1.430 0.450 4.370 0.770 ;
        RECT 1.430 0.440 4.140 0.450 ;
    END
  END DRAIN
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.180 2.450 0.450 2.480 ;
        RECT 0.180 1.920 0.460 2.450 ;
        RECT 0.000 1.620 0.460 1.920 ;
        RECT 0.000 1.600 0.470 1.620 ;
        RECT 0.180 1.170 0.470 1.600 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.020 5.660 1.340 5.700 ;
        RECT 2.110 5.660 2.430 5.700 ;
        RECT 1.020 5.470 1.350 5.660 ;
        RECT 2.110 5.470 2.440 5.660 ;
        RECT 1.020 5.440 1.340 5.470 ;
        RECT 2.110 5.440 2.430 5.470 ;
        RECT 1.570 4.980 1.890 5.020 ;
        RECT 2.600 5.000 2.770 5.890 ;
        RECT 3.150 5.690 3.320 5.890 ;
        RECT 3.150 5.650 3.530 5.690 ;
        RECT 3.150 5.460 3.540 5.650 ;
        RECT 3.150 5.430 3.530 5.460 ;
        RECT 1.570 4.790 1.900 4.980 ;
        RECT 2.600 4.960 2.980 5.000 ;
        RECT 1.570 4.760 1.890 4.790 ;
        RECT 2.600 4.770 2.990 4.960 ;
        RECT 2.600 4.740 2.980 4.770 ;
        RECT 2.600 3.650 2.770 4.740 ;
        RECT 1.570 3.610 1.890 3.650 ;
        RECT 2.600 3.610 2.980 3.650 ;
        RECT 1.570 3.420 1.900 3.610 ;
        RECT 2.600 3.490 2.990 3.610 ;
        RECT 3.150 3.490 3.320 5.430 ;
        RECT 3.700 4.990 3.870 5.890 ;
        RECT 3.700 4.950 4.090 4.990 ;
        RECT 3.700 4.760 4.100 4.950 ;
        RECT 3.700 4.730 4.090 4.760 ;
        RECT 3.700 3.650 3.870 4.730 ;
        RECT 3.700 3.610 4.080 3.650 ;
        RECT 3.700 3.490 4.090 3.610 ;
        RECT 4.250 3.490 4.420 5.890 ;
        RECT 4.800 3.490 4.970 5.890 ;
        RECT 5.350 3.490 5.520 5.890 ;
        RECT 2.660 3.420 2.990 3.490 ;
        RECT 3.760 3.420 4.090 3.490 ;
        RECT 1.570 3.390 1.890 3.420 ;
        RECT 2.660 3.390 2.980 3.420 ;
        RECT 3.760 3.390 4.080 3.420 ;
        RECT 0.950 2.920 1.120 3.180 ;
        RECT 0.950 2.880 1.330 2.920 ;
        RECT 0.950 2.800 1.340 2.880 ;
        RECT 1.500 2.800 1.670 3.180 ;
        RECT 2.050 2.920 2.220 3.180 ;
        RECT 2.050 2.880 2.430 2.920 ;
        RECT 2.050 2.800 2.440 2.880 ;
        RECT 1.010 2.690 1.340 2.800 ;
        RECT 2.110 2.690 2.440 2.800 ;
        RECT 1.010 2.660 1.330 2.690 ;
        RECT 2.110 2.660 2.430 2.690 ;
        RECT 0.240 1.200 0.410 2.420 ;
        RECT 1.010 1.510 1.330 1.550 ;
        RECT 2.110 1.510 2.430 1.550 ;
        RECT 1.010 1.320 1.340 1.510 ;
        RECT 2.110 1.320 2.440 1.510 ;
        RECT 1.010 1.290 1.330 1.320 ;
        RECT 2.110 1.290 2.430 1.320 ;
        RECT 0.190 0.910 0.700 1.010 ;
        RECT 0.190 0.870 0.760 0.910 ;
        RECT 2.600 0.870 2.770 3.180 ;
        RECT 3.150 2.920 3.320 3.180 ;
        RECT 3.150 2.880 3.530 2.920 ;
        RECT 3.150 2.690 3.540 2.880 ;
        RECT 3.150 2.660 3.530 2.690 ;
        RECT 3.150 1.550 3.320 2.660 ;
        RECT 3.150 1.510 3.530 1.550 ;
        RECT 3.150 1.320 3.540 1.510 ;
        RECT 3.150 1.290 3.530 1.320 ;
        RECT 0.190 0.680 0.770 0.870 ;
        RECT 1.570 0.830 1.890 0.870 ;
        RECT 2.600 0.830 2.980 0.870 ;
        RECT 0.200 0.650 0.760 0.680 ;
        RECT 0.200 0.440 0.710 0.650 ;
        RECT 1.570 0.640 1.900 0.830 ;
        RECT 2.600 0.710 2.990 0.830 ;
        RECT 3.150 0.710 3.320 1.290 ;
        RECT 3.700 0.880 3.870 3.180 ;
        RECT 3.700 0.840 4.080 0.880 ;
        RECT 3.700 0.710 4.090 0.840 ;
        RECT 4.250 0.710 4.420 3.110 ;
        RECT 4.800 0.710 4.970 3.110 ;
        RECT 5.350 0.710 5.520 3.110 ;
        RECT 2.660 0.640 2.990 0.710 ;
        RECT 3.760 0.650 4.090 0.710 ;
        RECT 1.570 0.610 1.890 0.640 ;
        RECT 2.660 0.610 2.980 0.640 ;
        RECT 3.760 0.620 4.080 0.650 ;
        RECT 0.200 0.400 0.770 0.440 ;
        RECT 0.200 0.210 0.780 0.400 ;
        RECT 0.200 0.180 0.770 0.210 ;
        RECT 0.200 0.000 0.710 0.180 ;
      LAYER mcon ;
        RECT 1.080 5.480 1.250 5.650 ;
        RECT 2.170 5.480 2.340 5.650 ;
        RECT 3.270 5.470 3.440 5.640 ;
        RECT 1.630 4.800 1.800 4.970 ;
        RECT 2.720 4.780 2.890 4.950 ;
        RECT 1.630 3.430 1.800 3.600 ;
        RECT 2.720 3.430 2.890 3.600 ;
        RECT 3.830 4.770 4.000 4.940 ;
        RECT 3.820 3.430 3.990 3.600 ;
        RECT 1.070 2.700 1.240 2.870 ;
        RECT 2.170 2.700 2.340 2.870 ;
        RECT 0.240 2.250 0.410 2.420 ;
        RECT 0.240 1.890 0.410 2.060 ;
        RECT 1.070 1.330 1.240 1.500 ;
        RECT 2.170 1.330 2.340 1.500 ;
        RECT 3.270 2.700 3.440 2.870 ;
        RECT 3.270 1.330 3.440 1.500 ;
        RECT 0.500 0.690 0.670 0.860 ;
        RECT 1.630 0.650 1.800 0.820 ;
        RECT 2.720 0.650 2.890 0.820 ;
        RECT 3.820 0.660 3.990 0.830 ;
        RECT 0.510 0.220 0.680 0.390 ;
      LAYER met1 ;
        RECT 1.010 5.410 1.330 5.730 ;
        RECT 2.100 5.410 2.420 5.730 ;
        RECT 3.200 5.400 3.520 5.720 ;
        RECT 1.560 4.730 1.880 5.050 ;
        RECT 2.650 4.710 2.970 5.030 ;
        RECT 3.760 4.700 4.080 5.020 ;
        RECT 1.560 3.360 1.880 3.680 ;
        RECT 2.650 3.360 2.970 3.680 ;
        RECT 3.750 3.360 4.070 3.680 ;
        RECT 1.000 2.630 1.320 2.950 ;
        RECT 2.100 2.630 2.420 2.950 ;
        RECT 3.200 2.630 3.520 2.950 ;
        RECT 1.000 1.260 1.320 1.580 ;
        RECT 2.100 1.260 2.420 1.580 ;
        RECT 3.200 1.260 3.520 1.580 ;
        RECT 0.430 0.620 0.750 0.940 ;
        RECT 1.560 0.580 1.880 0.900 ;
        RECT 2.650 0.580 2.970 0.900 ;
        RECT 3.750 0.590 4.070 0.910 ;
        RECT 0.440 0.150 0.760 0.470 ;
      LAYER via ;
        RECT 1.040 5.440 1.300 5.700 ;
        RECT 2.130 5.440 2.390 5.700 ;
        RECT 3.230 5.430 3.490 5.690 ;
        RECT 1.590 4.760 1.850 5.020 ;
        RECT 2.680 4.740 2.940 5.000 ;
        RECT 3.790 4.730 4.050 4.990 ;
        RECT 1.590 3.390 1.850 3.650 ;
        RECT 2.680 3.390 2.940 3.650 ;
        RECT 3.780 3.390 4.040 3.650 ;
        RECT 1.030 2.660 1.290 2.920 ;
        RECT 2.130 2.660 2.390 2.920 ;
        RECT 3.230 2.660 3.490 2.920 ;
        RECT 1.030 1.290 1.290 1.550 ;
        RECT 2.130 1.290 2.390 1.550 ;
        RECT 3.230 1.290 3.490 1.550 ;
        RECT 0.460 0.650 0.720 0.910 ;
        RECT 1.590 0.610 1.850 0.870 ;
        RECT 2.680 0.610 2.940 0.870 ;
        RECT 3.780 0.620 4.040 0.880 ;
        RECT 0.470 0.180 0.730 0.440 ;
  END
END sky130_hilas_nFETLarge

END LIBRARY