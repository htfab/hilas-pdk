magic
tech sky130A
timestamp 1629137141
<< error_p >>
rect 67 131 96 147
rect 146 131 175 147
rect 225 131 254 147
rect 304 131 333 147
rect 67 97 68 98
rect 95 97 96 98
rect 146 97 147 98
rect 174 97 175 98
rect 225 97 226 98
rect 253 97 254 98
rect 304 97 305 98
rect 332 97 333 98
rect 17 68 35 97
rect 66 96 97 97
rect 145 96 176 97
rect 224 96 255 97
rect 303 96 334 97
rect 67 89 96 96
rect 146 89 175 96
rect 225 89 254 96
rect 304 89 333 96
rect 67 75 77 89
rect 324 75 333 89
rect 67 69 96 75
rect 146 69 175 75
rect 225 69 254 75
rect 304 69 333 75
rect 66 68 97 69
rect 145 68 176 69
rect 224 68 255 69
rect 303 68 334 69
rect 366 68 383 97
rect 67 67 68 68
rect 95 67 96 68
rect 146 67 147 68
rect 174 67 175 68
rect 225 67 226 68
rect 253 67 254 68
rect 304 67 305 68
rect 332 67 333 68
rect 67 18 96 33
rect 146 18 175 33
rect 225 18 254 33
rect 304 18 333 33
<< nwell >>
rect 0 0 400 164
<< mvpmos >>
rect 35 97 366 131
rect 35 68 67 97
rect 96 68 146 97
rect 175 68 225 97
rect 254 68 304 97
rect 333 68 366 97
rect 35 33 366 68
<< mvpdiff >>
rect 67 91 96 97
rect 67 74 73 91
rect 90 74 96 91
rect 67 68 96 74
rect 146 91 175 97
rect 146 74 152 91
rect 169 74 175 91
rect 146 68 175 74
rect 225 91 254 97
rect 225 74 231 91
rect 248 74 254 91
rect 225 68 254 74
rect 304 91 333 97
rect 304 74 310 91
rect 327 74 333 91
rect 304 68 333 74
<< mvpdiffc >>
rect 73 74 90 91
rect 152 74 169 91
rect 231 74 248 91
rect 310 74 327 91
<< poly >>
rect 19 131 381 145
rect 19 33 35 131
rect 366 33 381 131
rect 19 19 381 33
<< locali >>
rect 35 125 366 131
rect 35 108 192 125
rect 209 108 366 125
rect 35 91 366 108
rect 35 74 73 91
rect 90 74 152 91
rect 169 74 231 91
rect 248 74 310 91
rect 327 74 366 91
rect 35 56 366 74
rect 35 39 192 56
rect 209 39 366 56
rect 35 33 366 39
<< viali >>
rect 192 108 209 125
rect 192 39 209 56
<< metal1 >>
rect 188 125 212 131
rect 188 108 192 125
rect 209 108 212 125
rect 188 67 212 108
rect 189 56 212 67
rect 189 39 192 56
rect 209 41 212 56
rect 209 39 213 41
rect 189 19 213 39
<< end >>
