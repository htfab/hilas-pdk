magic
tech sky130A
magscale 1 2
timestamp 1632256312
<< error_s >>
rect 120 292 180 306
rect 220 292 286 306
rect 120 284 170 292
rect 180 284 200 290
rect 108 282 200 284
rect 220 282 224 284
rect 108 280 224 282
rect 108 256 200 280
rect 220 256 224 280
rect 146 254 166 256
rect 180 254 220 256
rect 232 254 266 292
rect 298 256 338 270
rect 120 222 170 254
rect 180 224 200 254
rect 286 228 348 256
rect 232 222 348 228
rect 120 204 180 222
rect 220 214 336 222
rect 220 204 368 214
rect 232 196 368 204
rect 236 186 274 188
rect 276 186 368 196
rect 232 174 266 186
rect 286 184 368 186
rect 232 160 286 174
rect 294 160 300 184
rect 56 134 88 150
rect 170 148 232 160
rect 90 134 122 144
rect 56 102 122 134
rect 146 136 154 144
rect 146 102 156 136
rect 170 123 190 148
rect 180 106 190 123
rect 202 106 220 148
rect 224 145 232 148
rect 236 120 254 160
rect 286 159 348 160
rect 294 152 300 159
rect 294 140 340 152
rect 298 122 338 138
rect 286 112 348 122
rect 232 106 348 112
rect 170 102 348 106
rect 56 92 348 102
rect 56 86 94 92
rect 120 90 348 92
rect 56 84 88 86
rect 60 64 66 84
rect 120 80 336 90
rect 108 72 336 80
rect 108 70 310 72
rect 108 52 311 70
rect 170 50 286 52
rect 120 0 274 50
<< nmos >>
rect 170 254 224 256
rect 170 50 224 52
<< ndiff >>
rect 108 254 170 256
rect 224 254 286 256
rect 108 50 170 52
rect 224 50 286 52
<< psubdiff >>
rect 286 236 368 256
rect 286 202 310 236
rect 344 202 368 236
rect 286 184 368 202
rect 286 104 368 122
rect 286 70 310 104
rect 344 70 368 104
rect 286 50 368 70
<< psubdiffcont >>
rect 310 202 344 236
rect 310 70 344 104
<< poly >>
rect 170 280 224 282
rect 26 148 224 168
rect 26 138 170 148
rect 26 122 80 138
rect 170 24 224 26
<< locali >>
rect 276 236 346 252
rect 276 202 310 236
rect 344 202 346 236
rect 236 186 274 188
rect 276 186 346 202
rect 236 120 346 186
rect 276 104 346 120
rect 276 70 310 104
rect 344 70 346 104
rect 276 54 346 70
<< metal2 >>
rect 0 64 66 106
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1632251332
transform 1 0 294 0 1 140
box 0 0 46 58
use sky130_hilas_nFET03  sky130_hilas_nFET03_0
timestamp 1632251436
transform 1 0 170 0 1 64
box 0 0 178 122
use sky130_hilas_nFET03  sky130_hilas_nFET03_1
timestamp 1632251436
transform 1 0 170 0 1 196
box 0 0 178 122
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1632251356
transform 1 0 88 0 1 86
box 0 0 68 66
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1632251356
transform 1 0 98 0 1 216
box 0 0 68 66
use sky130_hilas_poly2li  sky130_hilas_poly2li_0
timestamp 1632251374
transform 1 0 44 0 1 84
box 0 0 54 66
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
