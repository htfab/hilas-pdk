* NGSPICE file created from /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_DAC6bit01.ext - technology: sky130A

.subckt sky130_hilas_pFETdevice01 w_n158_n156# a_n90_n38# $SUB a_42_n38# a_n158_36#
X0 a_42_n38# a_n158_36# a_n90_n38# w_n158_n156# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends

.subckt sky130_hilas_pFETdevice01aa a_n160_36# $SUB a_n92_n38# a_42_n38# w_n160_n156#
X0 a_42_n38# a_n160_36# a_n92_n38# w_n160_n156# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends

.subckt sky130_hilas_pFETdevice01a a_n160_36# $SUB a_n92_n38# a_42_n38# w_n160_n84#
X0 a_42_n38# a_n160_36# a_n92_n38# w_n160_n84# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends

.subckt sky130_hilas_DAC6TransistorStack01 sky130_hilas_pFETdevice01_3/a_n90_n38#
+ sky130_hilas_pFETdevice01a_0/a_42_n38# sky130_hilas_pFETdevice01a_0/a_n92_n38# sky130_hilas_pFETdevice01_0/a_n90_n38#
+ sky130_hilas_pFETdevice01aa_0/a_n92_n38# sky130_hilas_pFETdevice01_6/a_n158_36#
+ sky130_hilas_pFETdevice01_0/a_42_n38# sky130_hilas_pFETdevice01_4/a_42_n38# sky130_hilas_pFETdevice01aa_0/a_42_n38#
+ $SUB sky130_hilas_pFETdevice01_4/a_n158_36# sky130_hilas_pFETdevice01a_0/a_n160_36#
+ sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_3/a_n158_36#
+ sky130_hilas_pFETdevice01_3/a_42_n38# sky130_hilas_pFETdevice01_6/a_n90_n38# sky130_hilas_pFETdevice01aa_0/a_n160_36#
+ sky130_hilas_pFETdevice01_4/a_n90_n38# sky130_hilas_pFETdevice01_0/a_n158_36# sky130_hilas_pFETdevice01_6/a_42_n38#
Xsky130_hilas_pFETdevice01_0 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_0/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_0/a_42_n38# sky130_hilas_pFETdevice01_0/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01_3 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_3/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_3/a_42_n38# sky130_hilas_pFETdevice01_3/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01_4 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_4/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_4/a_42_n38# sky130_hilas_pFETdevice01_4/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01_6 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_6/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_6/a_42_n38# sky130_hilas_pFETdevice01_6/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01aa_0 sky130_hilas_pFETdevice01aa_0/a_n160_36# $SUB sky130_hilas_pFETdevice01aa_0/a_n92_n38#
+ sky130_hilas_pFETdevice01aa_0/a_42_n38# sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01aa
Xsky130_hilas_pFETdevice01a_0 sky130_hilas_pFETdevice01a_0/a_n160_36# $SUB sky130_hilas_pFETdevice01a_0/a_n92_n38#
+ sky130_hilas_pFETdevice01a_0/a_42_n38# sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01a
.ends

.subckt sky130_hilas_DAC6TransistorStack01a sky130_hilas_pFETdevice01aa_4/a_n160_36#
+ sky130_hilas_pFETdevice01aa_3/a_n160_36# $SUB sky130_hilas_pFETdevice01a_0/a_n160_36#
+ sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01aa_2/a_n160_36#
+ sky130_hilas_pFETdevice01aa_1/a_n160_36# sky130_hilas_pFETdevice01aa_0/a_n160_36#
Xsky130_hilas_pFETdevice01aa_0 sky130_hilas_pFETdevice01aa_0/a_n160_36# $SUB sky130_hilas_pFETdevice01aa_0/a_n92_n38#
+ sky130_hilas_pFETdevice01aa_0/a_42_n38# sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01aa
Xsky130_hilas_pFETdevice01aa_1 sky130_hilas_pFETdevice01aa_1/a_n160_36# $SUB sky130_hilas_pFETdevice01aa_1/a_n92_n38#
+ sky130_hilas_pFETdevice01aa_1/a_42_n38# sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01aa
Xsky130_hilas_pFETdevice01aa_2 sky130_hilas_pFETdevice01aa_2/a_n160_36# $SUB sky130_hilas_pFETdevice01aa_2/a_n92_n38#
+ sky130_hilas_pFETdevice01aa_2/a_42_n38# sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01aa
Xsky130_hilas_pFETdevice01aa_3 sky130_hilas_pFETdevice01aa_3/a_n160_36# $SUB sky130_hilas_pFETdevice01aa_3/a_n92_n38#
+ sky130_hilas_pFETdevice01aa_3/a_42_n38# sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01aa
Xsky130_hilas_pFETdevice01aa_4 sky130_hilas_pFETdevice01aa_4/a_n160_36# $SUB sky130_hilas_pFETdevice01aa_4/a_n92_n38#
+ sky130_hilas_pFETdevice01aa_4/a_42_n38# sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01aa
Xsky130_hilas_pFETdevice01a_0 sky130_hilas_pFETdevice01a_0/a_n160_36# $SUB sky130_hilas_pFETdevice01a_0/a_n92_n38#
+ sky130_hilas_pFETdevice01a_0/a_42_n38# sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01a
.ends

.subckt sky130_hilas_DAC_bit6_01 $SUB
Xsky130_hilas_DAC6TransistorStack01_0 sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_3/a_n90_n38#
+ sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01a_0/a_42_n38# sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01a_0/a_n92_n38#
+ sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_0/a_n90_n38# sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01aa_0/a_n92_n38#
+ sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_6/a_n158_36# sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_0/a_42_n38#
+ sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_4/a_42_n38# sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01aa_0/a_42_n38#
+ $SUB sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_6/a_n158_36#
+ sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_6/a_n158_36# sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_6/a_n158_36# sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_3/a_42_n38#
+ sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_6/a_n90_n38# sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_6/a_n158_36#
+ sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_4/a_n90_n38# sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_6/a_n158_36#
+ sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_6/a_42_n38# sky130_hilas_DAC6TransistorStack01
Xsky130_hilas_DAC6TransistorStack01_1 sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_3/a_n90_n38#
+ sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01a_0/a_42_n38# sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01a_0/a_n92_n38#
+ sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_0/a_n90_n38# sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01aa_0/a_n92_n38#
+ sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_6/a_n158_36# sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_0/a_42_n38#
+ sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_4/a_42_n38# sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01aa_0/a_42_n38#
+ $SUB sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_6/a_n158_36#
+ sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_6/a_n158_36# sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_6/a_n158_36# sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_3/a_42_n38#
+ sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_6/a_n90_n38# sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_6/a_n158_36#
+ sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_4/a_n90_n38# sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_6/a_n158_36#
+ sky130_hilas_DAC6TransistorStack01_1/sky130_hilas_pFETdevice01_6/a_42_n38# sky130_hilas_DAC6TransistorStack01
Xsky130_hilas_DAC6TransistorStack01a_0 sky130_hilas_poly2m2_11/a_n18_n16# m2_836_2204#
+ $SUB sky130_hilas_DAC6TransistorStack01a_0/sky130_hilas_pFETdevice01a_0/a_n160_36#
+ sky130_hilas_DAC6TransistorStack01a_0/sky130_hilas_pFETdevice01a_0/w_n160_n84# m2_836_1962#
+ sky130_hilas_poly2m2_12/a_n18_n16# sky130_hilas_DAC6TransistorStack01a_0/sky130_hilas_pFETdevice01aa_0/a_n160_36#
+ sky130_hilas_DAC6TransistorStack01a
Xsky130_hilas_DAC6TransistorStack01a_1 sky130_hilas_DAC6TransistorStack01a_1/sky130_hilas_pFETdevice01aa_4/a_n160_36#
+ sky130_hilas_DAC6TransistorStack01a_1/sky130_hilas_pFETdevice01aa_3/a_n160_36# $SUB
+ sky130_hilas_DAC6TransistorStack01a_1/sky130_hilas_pFETdevice01a_0/a_n160_36# sky130_hilas_DAC6TransistorStack01a_1/sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_DAC6TransistorStack01a_1/sky130_hilas_pFETdevice01aa_2/a_n160_36# sky130_hilas_DAC6TransistorStack01a_1/sky130_hilas_pFETdevice01aa_1/a_n160_36#
+ sky130_hilas_DAC6TransistorStack01a_1/sky130_hilas_pFETdevice01aa_0/a_n160_36# sky130_hilas_DAC6TransistorStack01a
.ends

.subckt sky130_hilas_pFETdevice01d w_n158_n156# a_n90_n38# $SUB a_n36_n84# a_42_n38#
+ sky130_hilas_poly2m1_0/a_n18_n16#
X0 a_42_n38# a_n36_n84# a_n90_n38# w_n158_n156# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends

.subckt sky130_hilas_DAC6TransistorStack01b sky130_hilas_pFETdevice01_0/a_n90_n38#
+ sky130_hilas_pFETdevice01_6/a_n158_36# sky130_hilas_pFETdevice01d_0/a_n90_n38# sky130_hilas_pFETdevice01d_0/a_n36_n84#
+ sky130_hilas_pFETdevice01_0/a_42_n38# sky130_hilas_pFETdevice01_4/a_42_n38# $SUB
+ sky130_hilas_pFETdevice01_4/a_n158_36# sky130_hilas_pFETdevice01a_0/a_n160_36# sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01d_0/sky130_hilas_poly2m1_0/a_n18_n16# sky130_hilas_pFETdevice01_6/a_n90_n38#
+ sky130_hilas_pFETdevice01aa_0/a_n160_36# sky130_hilas_pFETdevice01_4/a_n90_n38#
+ sky130_hilas_pFETdevice01_0/a_n158_36# sky130_hilas_pFETdevice01d_0/a_42_n38# sky130_hilas_pFETdevice01_6/a_42_n38#
Xsky130_hilas_pFETdevice01d_0 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01d_0/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01d_0/a_n36_n84# sky130_hilas_pFETdevice01d_0/a_42_n38#
+ sky130_hilas_pFETdevice01d_0/sky130_hilas_poly2m1_0/a_n18_n16# sky130_hilas_pFETdevice01d
Xsky130_hilas_pFETdevice01_0 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_0/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_0/a_42_n38# sky130_hilas_pFETdevice01_0/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01_4 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_4/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_4/a_42_n38# sky130_hilas_pFETdevice01_4/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01_6 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_6/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_6/a_42_n38# sky130_hilas_pFETdevice01_6/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01aa_0 sky130_hilas_pFETdevice01aa_0/a_n160_36# $SUB sky130_hilas_pFETdevice01aa_0/a_n92_n38#
+ sky130_hilas_pFETdevice01aa_0/a_42_n38# sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01aa
Xsky130_hilas_pFETdevice01a_0 sky130_hilas_pFETdevice01a_0/a_n160_36# $SUB sky130_hilas_pFETdevice01a_0/a_n92_n38#
+ sky130_hilas_pFETdevice01a_0/a_42_n38# sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01a
.ends

.subckt sky130_hilas_pFETdevice01b w_n158_n156# $SUB a_n36_n84#
X0 a_42_n38# a_n36_n84# a_n90_n38# w_n158_n156# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends

.subckt sky130_hilas_DAC6TransistorStack01c sky130_hilas_pFETdevice01_3/a_n90_n38#
+ sky130_hilas_pFETdevice01b_1/a_n36_n84# sky130_hilas_pFETdevice01_0/a_n90_n38# sky130_hilas_pFETdevice01_6/a_n158_36#
+ sky130_hilas_pFETdevice01_0/a_42_n38# $SUB sky130_hilas_pFETdevice01a_0/a_n160_36#
+ sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_3/a_n158_36#
+ sky130_hilas_pFETdevice01_3/a_42_n38# sky130_hilas_pFETdevice01_6/a_n90_n38# sky130_hilas_pFETdevice01aa_0/a_n160_36#
+ sky130_hilas_pFETdevice01_0/a_n158_36# sky130_hilas_pFETdevice01_6/a_42_n38#
Xsky130_hilas_pFETdevice01b_1 sky130_hilas_pFETdevice01a_0/w_n160_n84# $SUB sky130_hilas_pFETdevice01b_1/a_n36_n84#
+ sky130_hilas_pFETdevice01b
Xsky130_hilas_pFETdevice01_0 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_0/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_0/a_42_n38# sky130_hilas_pFETdevice01_0/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01_3 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_3/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_3/a_42_n38# sky130_hilas_pFETdevice01_3/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01_6 sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01_6/a_n90_n38#
+ $SUB sky130_hilas_pFETdevice01_6/a_42_n38# sky130_hilas_pFETdevice01_6/a_n158_36#
+ sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01aa_0 sky130_hilas_pFETdevice01aa_0/a_n160_36# $SUB sky130_hilas_pFETdevice01aa_0/a_n92_n38#
+ sky130_hilas_pFETdevice01aa_0/a_42_n38# sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01aa
Xsky130_hilas_pFETdevice01a_0 sky130_hilas_pFETdevice01a_0/a_n160_36# $SUB sky130_hilas_pFETdevice01a_0/a_n92_n38#
+ sky130_hilas_pFETdevice01a_0/a_42_n38# sky130_hilas_pFETdevice01a_0/w_n160_n84#
+ sky130_hilas_pFETdevice01a
.ends

.subckt sky130_hilas_DAC5bit01 A0 A2 A3 A4 Vdd Drain $SUB
Xsky130_hilas_DAC6TransistorStack01_0[0] Vdd sky130_hilas_DAC6TransistorStack01_0[0]/sky130_hilas_pFETdevice01a_0/a_42_n38#
+ sky130_hilas_DAC6TransistorStack01_0[0]/sky130_hilas_pFETdevice01a_0/a_n92_n38#
+ Vdd sky130_hilas_DAC6TransistorStack01_0[0]/sky130_hilas_pFETdevice01aa_0/a_n92_n38#
+ A4 Drain Drain sky130_hilas_DAC6TransistorStack01_0[0]/sky130_hilas_pFETdevice01aa_0/a_42_n38#
+ $SUB sky130_hilas_poly2m2_11/a_n18_n16# sky130_hilas_DAC6TransistorStack01a_0/sky130_hilas_pFETdevice01aa_0/a_n160_36#
+ w_1238_2040# A3 Drain Vdd A4 Vdd sky130_hilas_poly2m2_12/a_n18_n16# Drain sky130_hilas_DAC6TransistorStack01
Xsky130_hilas_DAC6TransistorStack01_0[1] Vdd sky130_hilas_DAC6TransistorStack01_0[1]/sky130_hilas_pFETdevice01a_0/a_42_n38#
+ sky130_hilas_DAC6TransistorStack01_0[1]/sky130_hilas_pFETdevice01a_0/a_n92_n38#
+ Vdd sky130_hilas_DAC6TransistorStack01_0[1]/sky130_hilas_pFETdevice01aa_0/a_n92_n38#
+ A4 Drain Drain sky130_hilas_DAC6TransistorStack01_0[1]/sky130_hilas_pFETdevice01aa_0/a_42_n38#
+ $SUB A3 sky130_hilas_poly2m2_12/a_n18_n16# w_1238_2040# A4 Drain Vdd A3 Vdd sky130_hilas_poly2m2_11/a_n18_n16#
+ Drain sky130_hilas_DAC6TransistorStack01
Xsky130_hilas_DAC6TransistorStack01_0[2] Vdd sky130_hilas_DAC6TransistorStack01_0[2]/sky130_hilas_pFETdevice01a_0/a_42_n38#
+ sky130_hilas_DAC6TransistorStack01_0[2]/sky130_hilas_pFETdevice01a_0/a_n92_n38#
+ Vdd sky130_hilas_DAC6TransistorStack01_0[2]/sky130_hilas_pFETdevice01aa_0/a_n92_n38#
+ A3 Drain Drain sky130_hilas_DAC6TransistorStack01_0[2]/sky130_hilas_pFETdevice01aa_0/a_42_n38#
+ $SUB A4 sky130_hilas_poly2m2_11/a_n18_n16# w_1238_2040# A4 Drain Vdd A4 Vdd A3 Drain
+ sky130_hilas_DAC6TransistorStack01
Xsky130_hilas_DAC6TransistorStack01_2[0] Vdd sky130_hilas_DAC6TransistorStack01_2[0]/sky130_hilas_pFETdevice01a_0/a_42_n38#
+ sky130_hilas_DAC6TransistorStack01_2[0]/sky130_hilas_pFETdevice01a_0/a_n92_n38#
+ Vdd sky130_hilas_DAC6TransistorStack01_2[0]/sky130_hilas_pFETdevice01aa_0/a_n92_n38#
+ A3 Drain Drain sky130_hilas_DAC6TransistorStack01_2[0]/sky130_hilas_pFETdevice01aa_0/a_42_n38#
+ $SUB A4 A4 w_1238_2040# A4 Drain Vdd A2 Vdd A3 Drain sky130_hilas_DAC6TransistorStack01
Xsky130_hilas_DAC6TransistorStack01_2[1] Vdd sky130_hilas_DAC6TransistorStack01_2[1]/sky130_hilas_pFETdevice01a_0/a_42_n38#
+ sky130_hilas_DAC6TransistorStack01_2[1]/sky130_hilas_pFETdevice01a_0/a_n92_n38#
+ Vdd sky130_hilas_DAC6TransistorStack01_2[1]/sky130_hilas_pFETdevice01aa_0/a_n92_n38#
+ A2 Drain Drain sky130_hilas_DAC6TransistorStack01_2[1]/sky130_hilas_pFETdevice01aa_0/a_42_n38#
+ $SUB A4 A3 w_1238_2040# A3 Drain Vdd m2_764_1430# Vdd A4 Drain sky130_hilas_DAC6TransistorStack01
Xsky130_hilas_DAC6TransistorStack01_2[2] Vdd sky130_hilas_DAC6TransistorStack01_2[2]/sky130_hilas_pFETdevice01a_0/a_42_n38#
+ sky130_hilas_DAC6TransistorStack01_2[2]/sky130_hilas_pFETdevice01a_0/a_n92_n38#
+ Vdd sky130_hilas_DAC6TransistorStack01_2[2]/sky130_hilas_pFETdevice01aa_0/a_n92_n38#
+ m2_764_1430# Drain Drain sky130_hilas_DAC6TransistorStack01_2[2]/sky130_hilas_pFETdevice01aa_0/a_42_n38#
+ $SUB A3 A4 w_1238_2040# A2 Drain Vdd sky130_hilas_DAC6TransistorStack01a_1/sky130_hilas_pFETdevice01aa_2/a_n160_36#
+ Vdd A4 Drain sky130_hilas_DAC6TransistorStack01
Xsky130_hilas_DAC6TransistorStack01b_0 Vdd A4 Vdd A0 Drain Drain $SUB A4 A3 w_1238_2040#
+ A3 Vdd A4 Vdd A4 Drain Drain sky130_hilas_DAC6TransistorStack01b
Xsky130_hilas_DAC6TransistorStack01c_0 Vdd A3 Vdd A4 Drain $SUB A4 w_1238_2040# A4
+ Drain Vdd A3 A4 Drain sky130_hilas_DAC6TransistorStack01c
Xsky130_hilas_DAC6TransistorStack01a_0 sky130_hilas_poly2m2_11/a_n18_n16# A4 $SUB
+ sky130_hilas_DAC6TransistorStack01a_0/sky130_hilas_pFETdevice01a_0/a_n160_36# w_1238_2040#
+ A3 sky130_hilas_poly2m2_12/a_n18_n16# sky130_hilas_DAC6TransistorStack01a_0/sky130_hilas_pFETdevice01aa_0/a_n160_36#
+ sky130_hilas_DAC6TransistorStack01a
Xsky130_hilas_DAC6TransistorStack01a_1 m2_764_1430# sky130_hilas_DAC6TransistorStack01a_1/sky130_hilas_pFETdevice01aa_3/a_n160_36#
+ $SUB A4 w_1238_2040# sky130_hilas_DAC6TransistorStack01a_1/sky130_hilas_pFETdevice01aa_2/a_n160_36#
+ A2 A3 sky130_hilas_DAC6TransistorStack01a
.ends


* Top level circuit /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_DAC6bit01

Xsky130_hilas_DAC_bit6_01_0 $SUB sky130_hilas_DAC_bit6_01
Xsky130_hilas_DAC5bit01_0 sky130_hilas_DAC5bit01_0/A0 sky130_hilas_DAC5bit01_0/A2
+ sky130_hilas_DAC5bit01_0/A3 sky130_hilas_DAC5bit01_0/A4 sky130_hilas_DAC5bit01_0/Vdd
+ sky130_hilas_DAC5bit01_0/Drain $SUB sky130_hilas_DAC5bit01
.end

