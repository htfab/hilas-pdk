magic
tech sky130A
timestamp 1628707329
<< error_p >>
rect 11 206 13 256
rect 53 206 55 256
rect 146 206 149 256
rect 188 206 191 256
rect 11 127 13 177
rect 53 127 55 177
rect 146 127 149 177
rect 188 127 191 177
rect 254 69 304 75
rect 326 69 376 75
rect 254 27 304 33
rect 326 27 376 33
<< nwell >>
rect 112 0 443 317
<< mvnmos >>
rect 13 206 53 256
rect 13 127 53 177
<< mvpmos >>
rect 149 206 188 256
rect 149 127 188 177
rect 252 100 303 284
rect 254 33 304 69
rect 326 33 376 69
<< mvndiff >>
rect 13 279 53 284
rect 13 262 24 279
rect 42 262 53 279
rect 13 256 53 262
rect 13 200 53 206
rect 13 183 23 200
rect 42 183 53 200
rect 13 177 53 183
rect 13 121 53 127
rect 13 104 24 121
rect 42 104 53 121
rect 13 100 53 104
<< mvpdiff >>
rect 149 279 188 284
rect 149 262 160 279
rect 177 262 188 279
rect 149 256 188 262
rect 220 263 252 284
rect 220 246 227 263
rect 244 246 252 263
rect 220 229 252 246
rect 220 212 227 229
rect 244 212 252 229
rect 149 200 188 206
rect 149 183 160 200
rect 177 183 188 200
rect 149 177 188 183
rect 220 195 252 212
rect 220 178 227 195
rect 244 178 252 195
rect 220 161 252 178
rect 220 144 227 161
rect 244 144 252 161
rect 220 127 252 144
rect 149 121 188 127
rect 149 104 160 121
rect 177 104 188 121
rect 149 100 188 104
rect 220 110 227 127
rect 244 110 252 127
rect 220 100 252 110
rect 303 262 331 284
rect 303 245 310 262
rect 327 245 331 262
rect 303 228 331 245
rect 303 211 310 228
rect 327 211 331 228
rect 303 194 331 211
rect 303 177 310 194
rect 327 177 331 194
rect 303 160 331 177
rect 303 143 310 160
rect 327 143 331 160
rect 303 126 331 143
rect 303 109 310 126
rect 327 109 331 126
rect 303 100 331 109
rect 220 63 254 69
rect 220 46 229 63
rect 247 46 254 63
rect 220 33 254 46
rect 304 33 326 69
rect 376 63 410 69
rect 376 46 383 63
rect 403 46 410 63
rect 376 33 410 46
<< mvndiffc >>
rect 24 262 42 279
rect 23 183 42 200
rect 24 104 42 121
<< mvpdiffc >>
rect 160 262 177 279
rect 227 246 244 263
rect 227 212 244 229
rect 160 183 177 200
rect 227 178 244 195
rect 227 144 244 161
rect 160 104 177 121
rect 227 110 244 127
rect 310 245 327 262
rect 310 211 327 228
rect 310 177 327 194
rect 310 143 327 160
rect 310 109 327 126
rect 229 46 247 63
rect 383 46 403 63
<< mvnsubdiff >>
rect 376 127 410 141
rect 376 109 383 127
rect 403 109 410 127
rect 376 97 410 109
<< mvnsubdiffcont >>
rect 383 109 403 127
<< poly >>
rect 252 284 303 297
rect 0 206 13 256
rect 53 206 149 256
rect 188 206 201 256
rect 0 127 13 177
rect 53 127 149 177
rect 188 127 201 177
rect 343 206 378 214
rect 343 189 355 206
rect 372 189 378 206
rect 343 181 378 189
rect 343 180 372 181
rect 343 151 370 180
rect 68 92 134 94
rect 252 92 303 100
rect 0 77 304 92
rect 347 85 370 151
rect 347 83 376 85
rect 254 69 304 77
rect 326 69 376 83
rect 254 18 304 33
rect 326 18 376 33
<< polycont >>
rect 355 189 372 206
<< locali >>
rect 16 262 24 279
rect 42 262 50 279
rect 152 262 160 279
rect 177 262 185 279
rect 227 263 244 271
rect 227 229 244 246
rect 15 183 23 200
rect 42 183 50 200
rect 152 183 160 200
rect 177 183 185 200
rect 227 195 244 212
rect 227 161 244 178
rect 227 127 244 144
rect 15 104 24 121
rect 42 104 50 121
rect 152 104 160 121
rect 177 104 185 121
rect 227 102 244 110
rect 310 228 327 245
rect 310 194 327 211
rect 346 206 373 214
rect 346 189 355 206
rect 372 189 373 206
rect 346 181 373 189
rect 310 160 327 177
rect 347 177 367 181
rect 347 158 348 177
rect 366 158 367 177
rect 347 152 367 158
rect 347 151 366 152
rect 310 126 327 143
rect 383 134 404 135
rect 310 101 327 109
rect 382 127 404 134
rect 382 109 383 127
rect 403 109 404 127
rect 382 93 404 109
rect 382 76 384 93
rect 401 76 404 93
rect 383 73 404 76
rect 383 63 403 73
rect 220 46 229 63
rect 247 46 255 63
rect 383 38 403 46
<< viali >>
rect 310 262 328 281
rect 348 158 366 177
rect 384 76 401 93
rect 202 46 220 63
<< metal1 >>
rect 307 281 331 287
rect 307 262 310 281
rect 328 262 331 281
rect 307 249 331 262
rect 350 206 366 308
rect 346 182 369 206
rect 346 181 370 182
rect 345 177 370 181
rect 345 158 348 177
rect 366 158 370 177
rect 345 154 370 158
rect 347 151 369 154
rect 195 84 226 87
rect 195 58 198 84
rect 224 58 226 84
rect 195 46 202 58
rect 220 46 226 58
rect 195 43 226 46
rect 347 6 366 151
rect 391 139 407 308
rect 391 130 408 139
rect 380 125 408 130
rect 380 93 407 125
rect 380 76 384 93
rect 401 76 407 93
rect 380 70 407 76
rect 391 6 407 70
<< via1 >>
rect 198 63 224 84
rect 198 58 202 63
rect 202 58 220 63
rect 220 58 224 63
<< metal2 >>
rect 195 84 226 87
rect 195 58 198 84
rect 224 73 226 84
rect 224 58 443 73
rect 195 55 443 58
rect 195 54 226 55
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
