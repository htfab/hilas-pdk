magic
tech sky130A
timestamp 1627737364
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_2
timestamp 1627737364
transform 1 0 12 0 1 13
box 147 -22 266 265
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_1
timestamp 1627737364
transform 1 0 -43 0 1 13
box 147 -22 266 265
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_0
timestamp 1627737364
transform 1 0 -98 0 1 13
box 147 -22 266 265
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_4
timestamp 1627737364
transform 1 0 -153 0 1 13
box 147 -22 266 265
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_3
timestamp 1627737364
transform 1 0 67 0 1 13
box 147 -22 266 265
<< end >>
