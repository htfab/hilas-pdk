magic
tech sky130A
timestamp 1627737364
<< metal1 >>
rect -2053 27123 -1982 27519
rect -898 26641 -826 27030
rect -2054 24263 -1984 24659
rect -898 23782 -826 24171
rect -2052 21404 -1982 21800
rect -898 20922 -826 21311
rect -2054 18545 -1984 18941
rect -898 18065 -826 18454
rect -2054 15685 -1984 16081
rect -899 15205 -827 15594
rect -2053 12827 -1983 13223
rect -898 12346 -826 12735
rect -2053 9967 -1983 10363
rect -898 9486 -826 9875
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_12
timestamp 1627735001
transform 0 1 -1755 1 0 26614
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_11
timestamp 1627735001
transform 0 1 -1755 1 0 23755
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_10
timestamp 1627735001
transform 0 1 -1755 1 0 20896
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_5
timestamp 1627735001
transform 0 1 -1755 1 0 18037
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_8
timestamp 1627735001
transform 0 1 -1755 1 0 15178
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_7
timestamp 1627735001
transform 0 1 -1755 1 0 12319
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_9
timestamp 1627735001
transform 0 1 -1755 1 0 9460
box -745 -229 2114 858
<< labels >>
rlabel metal1 -898 9486 -826 9875 0 IO7
port 1 nsew
rlabel metal1 -898 12346 -826 12735 0 IO8
port 2 nsew
rlabel metal1 -899 15205 -827 15594 0 IO9
port 3 nsew
rlabel metal1 -898 18065 -826 18454 0 IO10
port 4 nsew
rlabel metal1 -898 20922 -826 21311 0 IO11
port 5 nsew
rlabel metal1 -898 23782 -826 24171 0 IO12
port 7 nsew
rlabel metal1 -898 26641 -826 27030 0 IO13
port 6 nsew
rlabel metal1 -2053 9967 -1983 10363 0 PIN1
port 8 nsew
rlabel metal1 -2053 12827 -1983 13223 0 PIN2
port 9 nsew
rlabel metal1 -2054 15685 -1984 16081 0 PIN3
port 10 nsew
rlabel metal1 -2054 18545 -1984 18941 0 PIN4
port 11 nsew
rlabel metal1 -2052 21404 -1982 21800 0 PIN5
port 12 nsew
rlabel metal1 -2054 24263 -1984 24659 0 PIN6
port 13 nsew
rlabel metal1 -2053 27123 -1983 27519 0 PIN7
port 14 nsew
<< end >>
