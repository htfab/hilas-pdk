magic
tech sky130A
timestamp 1628704378
<< checkpaint >>
rect -591 731 703 746
rect -605 678 703 731
rect -606 663 703 678
rect -620 -547 703 663
rect -620 -562 689 -547
rect -620 -615 688 -562
rect -620 -630 674 -615
<< nmos >>
rect 90 42 110 101
rect 196 42 216 101
<< ndiff >>
rect 224 101 254 109
rect 61 97 90 101
rect 61 80 67 97
rect 84 80 90 97
rect 61 63 90 80
rect 61 46 67 63
rect 84 46 90 63
rect 61 42 90 46
rect 110 97 140 101
rect 110 80 117 97
rect 134 80 140 97
rect 110 63 140 80
rect 110 46 117 63
rect 134 46 140 63
rect 110 42 140 46
rect 167 97 196 101
rect 167 80 173 97
rect 190 80 196 97
rect 167 63 196 80
rect 167 46 173 63
rect 190 46 196 63
rect 167 42 196 46
rect 216 97 254 101
rect 216 80 230 97
rect 247 80 254 97
rect 216 63 254 80
rect 216 46 230 63
rect 247 46 254 63
rect 216 42 254 46
rect 224 34 254 42
<< ndiffc >>
rect 67 80 84 97
rect 67 46 84 63
rect 117 80 134 97
rect 117 46 134 63
rect 173 80 190 97
rect 173 46 190 63
rect 230 80 247 97
rect 230 46 247 63
<< psubdiff >>
rect 254 97 283 109
rect 254 80 264 97
rect 281 80 283 97
rect 254 63 283 80
rect 254 46 264 63
rect 281 46 283 63
rect 254 34 283 46
<< psubdiffcont >>
rect 264 80 281 97
rect 264 46 281 63
<< poly >>
rect 151 137 216 142
rect 151 120 159 137
rect 176 120 216 137
rect 151 114 216 120
rect 90 101 110 114
rect 196 101 216 114
rect 90 33 110 42
rect 45 23 110 33
rect 196 29 216 42
rect 45 6 53 23
rect 70 6 110 23
rect 45 1 110 6
<< polycont >>
rect 159 120 176 137
rect 53 6 70 23
<< locali >>
rect 119 137 140 139
rect 117 120 121 137
rect 138 120 159 137
rect 176 120 184 137
rect 117 97 142 120
rect 230 97 281 105
rect 58 80 67 97
rect 84 80 92 97
rect 109 80 117 97
rect 134 80 142 97
rect 164 80 173 97
rect 190 80 198 97
rect 247 80 264 97
rect 58 63 92 80
rect 117 63 134 80
rect 173 63 190 80
rect 230 63 247 80
rect 264 63 281 80
rect 58 46 67 63
rect 84 46 92 63
rect 109 46 117 63
rect 134 46 142 63
rect 164 46 173 63
rect 190 46 198 63
rect 247 46 264 63
rect 173 23 190 46
rect 230 38 281 46
rect 44 6 53 23
rect 70 6 190 23
<< viali >>
rect 121 120 138 137
rect 247 63 264 80
<< metal1 >>
rect 118 137 141 143
rect 118 120 121 137
rect 138 120 141 137
rect 118 0 141 120
rect 244 80 267 129
rect 244 63 247 80
rect 264 63 267 80
rect 244 0 267 63
<< metal2 >>
rect 54 74 283 90
rect 0 4 12 25
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628704305
transform 1 0 24 0 1 15
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628704305
transform 1 0 39 0 1 83
box 0 0 34 33
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
