magic
tech sky130A
timestamp 1628707371
<< metal3 >>
rect 0 0 284 286
<< mimcap >>
rect 42 140 242 243
rect 42 127 127 140
rect 141 127 242 140
rect 42 43 242 127
<< mimcapcontact >>
rect 127 127 141 140
<< metal4 >>
rect 112 152 157 153
rect 110 140 162 152
rect 110 127 127 140
rect 141 127 162 140
rect 110 103 162 127
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
