magic
tech sky130A
timestamp 1627255200
<< nwell >>
rect -61 89 67 373
<< pmos >>
rect -40 295 28 325
rect -40 164 28 194
<< pdiff >>
rect -40 349 28 354
rect -40 331 -33 349
rect -15 331 3 349
rect 21 331 28 349
rect -40 325 28 331
rect -40 289 28 295
rect -40 271 -32 289
rect -15 271 4 289
rect 22 271 28 289
rect -40 265 28 271
rect -40 218 28 224
rect -40 201 -32 218
rect -14 201 4 218
rect 22 201 28 218
rect -40 194 28 201
rect -40 157 28 164
rect -40 140 -32 157
rect -14 140 4 157
rect 22 140 28 157
rect -40 131 28 140
<< pdiffc >>
rect -33 331 -15 349
rect 3 331 21 349
rect -32 271 -15 289
rect 4 271 22 289
rect -32 201 -14 218
rect 4 201 22 218
rect -32 140 -14 157
rect 4 140 22 157
<< nsubdiff >>
rect -40 253 28 265
rect -40 236 -32 253
rect -14 236 4 253
rect 22 236 28 253
rect -40 224 28 236
<< nsubdiffcont >>
rect -32 236 -14 253
rect 4 236 22 253
<< poly >>
rect -53 295 -40 325
rect 28 295 53 325
rect 36 194 53 295
rect -53 164 -40 194
rect 28 164 53 194
rect 36 112 53 164
<< locali >>
rect -41 331 -33 349
rect -15 331 3 349
rect 21 331 29 349
rect -40 271 -32 289
rect -15 271 4 289
rect 22 271 30 289
rect -40 253 30 271
rect -40 236 -32 253
rect -14 236 4 253
rect 22 236 30 253
rect -40 218 30 236
rect -40 201 -32 218
rect -14 201 4 218
rect 22 201 30 218
rect -40 140 -32 157
rect -14 140 4 157
rect 22 140 31 157
rect -5 112 31 140
rect -5 95 28 112
use sky130_hilas_poly2li  sky130_hilas_poly2li_0
timestamp 1627255200
transform 0 1 34 -1 0 108
box -9 -14 18 19
<< end >>
