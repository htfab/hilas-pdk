magic
tech sky130A
timestamp 1634057757
<< metal3 >>
rect 0 580 282 583
rect 0 2 720 580
rect 279 0 720 2
<< mimcap >>
rect 39 143 677 542
rect 39 142 155 143
rect 39 129 127 142
rect 141 129 155 142
rect 169 129 183 143
rect 197 129 211 143
rect 225 129 239 143
rect 253 129 267 143
rect 281 129 294 143
rect 308 129 322 143
rect 336 129 350 143
rect 364 129 677 143
rect 39 42 677 129
<< mimcapcontact >>
rect 127 129 141 142
rect 155 129 169 143
rect 183 129 197 143
rect 211 129 225 143
rect 239 129 253 143
rect 267 129 281 143
rect 294 129 308 143
rect 322 129 336 143
rect 350 129 364 143
<< metal4 >>
rect 89 143 393 157
rect 89 142 155 143
rect 89 129 127 142
rect 141 129 155 142
rect 169 129 183 143
rect 197 129 211 143
rect 225 129 239 143
rect 253 129 267 143
rect 281 129 294 143
rect 308 129 322 143
rect 336 129 350 143
rect 364 129 393 143
rect 89 110 393 129
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
