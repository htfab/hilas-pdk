VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_dac5bit01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_dac5bit01 ;
  ORIGIN -3.820 -5.240 ;
  SIZE 16.580 BY 5.970 ;
  OBS
      LAYER nwell ;
        RECT 6.190 10.200 17.620 10.270 ;
      LAYER li1 ;
        RECT 7.800 10.270 7.970 10.280 ;
        RECT 16.770 10.270 16.980 11.050 ;
        RECT 17.440 10.270 17.610 10.950 ;
        RECT 6.190 10.040 17.620 10.270 ;
        RECT 6.190 6.480 6.360 10.040 ;
        RECT 6.850 5.250 7.020 9.710 ;
        RECT 7.800 6.480 7.970 10.040 ;
        RECT 8.480 5.250 8.650 9.670 ;
        RECT 9.390 6.480 9.560 10.040 ;
        RECT 10.080 5.250 10.250 9.750 ;
        RECT 11.010 6.480 11.180 10.040 ;
        RECT 11.700 5.250 11.870 9.700 ;
        RECT 12.630 6.500 12.800 10.040 ;
        RECT 13.300 5.250 13.470 9.750 ;
        RECT 14.230 6.510 14.400 10.040 ;
        RECT 14.920 5.250 15.090 9.750 ;
        RECT 15.840 6.500 16.010 10.040 ;
        RECT 16.520 5.250 16.690 9.730 ;
        RECT 17.450 6.470 17.620 10.040 ;
        RECT 18.130 5.250 18.300 9.910 ;
      LAYER met1 ;
        RECT 10.560 8.800 14.010 8.970 ;
        RECT 12.110 6.270 12.290 7.810 ;
        RECT 13.810 6.960 14.010 8.800 ;
        RECT 6.860 5.250 20.300 5.480 ;
      LAYER met2 ;
        RECT 3.820 11.020 10.870 11.210 ;
        RECT 3.820 10.200 5.880 10.260 ;
        RECT 7.300 10.200 7.520 10.660 ;
        RECT 12.220 10.210 12.470 10.970 ;
        RECT 12.220 10.200 12.500 10.210 ;
        RECT 3.820 10.050 12.500 10.200 ;
        RECT 4.080 9.810 4.280 10.050 ;
        RECT 5.720 9.900 12.500 10.050 ;
        RECT 13.930 8.330 14.130 10.890 ;
        RECT 3.820 8.120 14.130 8.330 ;
        RECT 15.530 7.350 15.680 11.090 ;
        RECT 16.530 10.930 17.690 11.210 ;
        RECT 17.280 10.920 17.690 10.930 ;
        RECT 3.820 7.150 15.690 7.350 ;
        RECT 3.820 6.030 12.360 6.230 ;
  END
END sky130_hilas_dac5bit01
END LIBRARY

