magic
tech sky130A
timestamp 1628698522
<< error_p >>
rect -540 172 -533 173
rect -601 -66 -516 -60
rect -602 -94 -516 -66
rect -573 -97 -572 -94
rect -560 -97 -554 -94
rect -573 -100 -551 -97
rect -550 -100 -516 -94
rect -498 -95 -495 -92
rect -575 -103 -516 -100
rect -575 -106 -566 -103
rect -573 -122 -572 -106
rect -569 -114 -566 -106
rect -560 -106 -516 -103
rect -560 -114 -551 -106
rect -569 -117 -551 -114
rect -560 -120 -551 -117
rect -560 -122 -554 -120
rect -550 -122 -516 -106
rect -495 -96 -492 -95
rect -495 -121 -494 -96
rect -573 -123 -516 -122
<< nwell >>
rect -572 -43 -425 226
rect -601 -67 -425 -43
rect -602 -150 -425 -67
rect -572 -441 -425 -150
<< mvpmos >>
rect -521 116 -491 166
rect -521 -21 -491 30
rect -521 -94 -491 -42
rect -521 -175 -491 -123
rect -521 -246 -491 -196
rect -521 -381 -491 -331
<< mvndiff >>
rect -573 -123 -550 -94
<< mvpdiff >>
rect -521 189 -491 193
rect -521 172 -515 189
rect -498 172 -491 189
rect -521 166 -491 172
rect -521 110 -491 116
rect -521 93 -515 110
rect -497 93 -491 110
rect -521 88 -491 93
rect -521 53 -491 58
rect -521 36 -515 53
rect -497 36 -491 53
rect -521 30 -491 36
rect -521 -42 -491 -21
rect -521 -100 -491 -94
rect -521 -117 -515 -100
rect -497 -117 -491 -100
rect -521 -123 -491 -117
rect -521 -196 -491 -175
rect -521 -252 -491 -246
rect -521 -269 -515 -252
rect -497 -269 -491 -252
rect -521 -273 -491 -269
rect -521 -308 -491 -304
rect -521 -325 -515 -308
rect -497 -325 -491 -308
rect -521 -331 -491 -325
rect -521 -387 -491 -381
rect -521 -404 -515 -387
rect -497 -404 -491 -387
rect -521 -408 -491 -404
<< mvpdiffc >>
rect -515 172 -498 189
rect -515 93 -497 110
rect -515 36 -497 53
rect -515 -117 -497 -100
rect -515 -269 -497 -252
rect -515 -325 -497 -308
rect -515 -404 -497 -387
<< poly >>
rect -555 116 -521 166
rect -491 116 -478 166
rect -555 30 -534 116
rect -555 -21 -521 30
rect -491 -21 -476 30
rect -534 -94 -521 -42
rect -491 -94 -465 -42
rect -488 -123 -465 -94
rect -534 -175 -521 -123
rect -491 -175 -465 -123
rect -550 -246 -521 -196
rect -491 -246 -478 -196
rect -550 -331 -534 -246
rect -550 -381 -521 -331
rect -491 -381 -478 -331
rect -550 -382 -534 -381
<< locali >>
rect -522 172 -515 189
rect -498 172 -490 189
rect -523 93 -515 110
rect -497 93 -489 110
rect -523 36 -515 53
rect -497 36 -489 53
rect -554 -117 -540 -100
rect -522 -117 -515 -100
rect -497 -117 -489 -100
rect -523 -269 -515 -252
rect -497 -269 -489 -252
rect -523 -325 -515 -308
rect -497 -325 -489 -308
rect -523 -404 -515 -387
rect -497 -404 -489 -387
<< viali >>
rect -540 172 -522 189
rect -569 -117 -554 -100
rect -540 -117 -522 -100
<< metal1 >>
rect -536 196 -502 200
rect -536 195 -532 196
rect -546 189 -532 195
rect -506 195 -502 196
rect -546 172 -540 189
rect -546 170 -532 172
rect -506 170 -490 195
rect -536 167 -502 170
rect -546 -100 -520 -96
rect -546 -117 -540 -100
rect -522 -117 -520 -100
rect -546 -121 -520 -117
rect -495 -121 -492 -96
<< via1 >>
rect -532 189 -506 196
rect -532 172 -522 189
rect -522 172 -506 189
rect -532 170 -506 172
rect -520 -121 -495 -95
<< metal2 >>
rect -536 196 -502 200
rect -572 170 -532 196
rect -506 170 -453 196
rect -536 167 -502 170
rect -522 -94 -492 -93
rect -522 -95 -491 -94
rect -542 -121 -520 -95
rect -495 -121 -489 -95
rect -542 -122 -489 -121
rect -522 -124 -492 -122
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
