magic
tech sky130A
timestamp 1625668104
<< error_s >>
rect 2481 3932 2487 3938
rect 2598 3932 2604 3938
rect 3498 3932 3504 3938
rect 3615 3932 3621 3938
rect 2487 3681 2493 3687
rect 2592 3681 2598 3687
rect 3504 3681 3510 3687
rect 3609 3681 3615 3687
rect 2481 3631 2487 3637
rect 2598 3631 2604 3637
rect 2915 3627 2921 3633
rect 2968 3627 2974 3633
rect 3081 3627 3087 3633
rect 3134 3627 3140 3633
rect 3498 3631 3504 3637
rect 3615 3631 3621 3637
rect 2909 3577 2915 3583
rect 2974 3577 2980 3583
rect 3075 3577 3081 3583
rect 3140 3577 3146 3583
rect 3548 3258 3554 3264
rect 3653 3258 3659 3264
rect 4519 3258 4525 3264
rect 4624 3258 4630 3264
rect 3974 3248 3980 3254
rect 4027 3248 4033 3254
rect 4145 3248 4151 3254
rect 4198 3248 4204 3254
rect 3542 3194 3548 3200
rect 3659 3194 3665 3200
rect 3968 3198 3974 3204
rect 4033 3198 4039 3204
rect 4139 3198 4145 3204
rect 4204 3198 4210 3204
rect 4513 3194 4519 3200
rect 4630 3194 4636 3200
rect 3548 3141 3554 3147
rect 3653 3141 3659 3147
rect 3974 3139 3980 3145
rect 4027 3139 4033 3145
rect 4145 3139 4151 3145
rect 4198 3139 4204 3145
rect 4519 3141 4525 3147
rect 4624 3141 4630 3147
rect 6348 3132 6354 3138
rect 6453 3132 6459 3138
rect 3968 3089 3974 3095
rect 4033 3089 4039 3095
rect 4139 3089 4145 3095
rect 4204 3089 4210 3095
rect 3542 3077 3548 3083
rect 3659 3077 3665 3083
rect 4513 3077 4519 3083
rect 4630 3077 4636 3083
rect 6342 3082 6348 3088
rect 6459 3082 6465 3088
rect 3548 2956 3554 2962
rect 3653 2956 3659 2962
rect 4519 2956 4525 2962
rect 4624 2956 4630 2962
rect 3974 2950 3980 2956
rect 4027 2950 4033 2956
rect 4145 2950 4151 2956
rect 4198 2950 4204 2956
rect 6654 2913 6655 2926
rect 3968 2900 3974 2906
rect 4033 2900 4039 2906
rect 4139 2900 4145 2906
rect 4204 2900 4210 2906
rect 3542 2892 3548 2898
rect 3659 2892 3665 2898
rect 4513 2892 4519 2898
rect 4630 2892 4636 2898
rect 3548 2840 3554 2846
rect 3653 2840 3659 2846
rect 4519 2840 4525 2846
rect 4624 2840 4630 2846
rect 3974 2833 3980 2839
rect 4027 2833 4033 2839
rect 4145 2833 4151 2839
rect 4198 2833 4204 2839
rect 6348 2831 6354 2837
rect 6453 2831 6459 2837
rect 3968 2783 3974 2789
rect 4033 2783 4039 2789
rect 4139 2783 4145 2789
rect 4204 2783 4210 2789
rect 3542 2776 3548 2782
rect 3659 2776 3665 2782
rect 4513 2776 4519 2782
rect 4630 2776 4636 2782
rect 6342 2781 6348 2787
rect 6459 2781 6465 2787
rect 649 2645 678 2661
rect 728 2645 757 2661
rect 807 2645 836 2661
rect 886 2645 915 2661
rect 1196 2621 1202 2627
rect 2046 2621 2053 2627
rect 649 2611 650 2612
rect 677 2611 678 2612
rect 728 2611 729 2612
rect 756 2611 757 2612
rect 807 2611 808 2612
rect 835 2611 836 2612
rect 886 2611 887 2612
rect 914 2611 915 2612
rect 648 2610 679 2611
rect 727 2610 758 2611
rect 806 2610 837 2611
rect 885 2610 916 2611
rect 649 2603 678 2610
rect 728 2603 757 2610
rect 807 2603 836 2610
rect 886 2603 915 2610
rect 649 2589 659 2603
rect 906 2589 915 2603
rect 649 2583 678 2589
rect 728 2583 757 2589
rect 807 2583 836 2589
rect 886 2583 915 2589
rect 648 2582 679 2583
rect 727 2582 758 2583
rect 806 2582 837 2583
rect 885 2582 916 2583
rect 948 2582 965 2611
rect 649 2581 650 2582
rect 677 2581 678 2582
rect 728 2581 729 2582
rect 756 2581 757 2582
rect 807 2581 808 2582
rect 835 2581 836 2582
rect 886 2581 887 2582
rect 914 2581 915 2582
rect 649 2532 678 2547
rect 728 2532 757 2547
rect 807 2532 836 2547
rect 886 2532 915 2547
rect 649 2365 678 2381
rect 728 2365 757 2381
rect 807 2365 836 2381
rect 886 2365 915 2381
rect 2356 2362 2361 2363
rect 649 2331 650 2332
rect 677 2331 678 2332
rect 728 2331 729 2332
rect 756 2331 757 2332
rect 807 2331 808 2332
rect 835 2331 836 2332
rect 886 2331 887 2332
rect 914 2331 915 2332
rect 648 2330 679 2331
rect 727 2330 758 2331
rect 806 2330 837 2331
rect 885 2330 916 2331
rect 649 2323 678 2330
rect 728 2323 757 2330
rect 807 2323 836 2330
rect 886 2323 915 2330
rect 649 2309 659 2323
rect 906 2309 915 2323
rect 649 2303 678 2309
rect 728 2303 757 2309
rect 807 2303 836 2309
rect 886 2303 915 2309
rect 648 2302 679 2303
rect 727 2302 758 2303
rect 806 2302 837 2303
rect 885 2302 916 2303
rect 948 2302 965 2331
rect 649 2301 650 2302
rect 677 2301 678 2302
rect 728 2301 729 2302
rect 756 2301 757 2302
rect 807 2301 808 2302
rect 835 2301 836 2302
rect 886 2301 887 2302
rect 914 2301 915 2302
rect 649 2252 678 2267
rect 728 2252 757 2267
rect 807 2252 836 2267
rect 886 2252 915 2267
rect -210 2251 -209 2252
rect -182 2251 -181 2252
rect -260 2222 -242 2251
rect -211 2250 -180 2251
rect -210 2241 -181 2250
rect -210 2232 -200 2241
rect -191 2232 -181 2241
rect -210 2223 -181 2232
rect -211 2222 -180 2223
rect -149 2222 -131 2251
rect -210 2221 -209 2222
rect -182 2221 -181 2222
rect 259 2221 265 2227
rect 364 2221 370 2227
rect 649 2210 678 2226
rect 728 2210 757 2226
rect 807 2210 836 2226
rect 886 2210 915 2226
rect 2648 2195 2649 2250
rect -210 2172 -181 2190
rect 253 2171 259 2177
rect 370 2171 376 2177
rect 649 2176 650 2177
rect 677 2176 678 2177
rect 728 2176 729 2177
rect 756 2176 757 2177
rect 807 2176 808 2177
rect 835 2176 836 2177
rect 886 2176 887 2177
rect 914 2176 915 2177
rect 599 2147 617 2176
rect 648 2175 679 2176
rect 727 2175 758 2176
rect 806 2175 837 2176
rect 885 2175 916 2176
rect 649 2168 678 2175
rect 728 2168 757 2175
rect 807 2168 836 2175
rect 886 2168 915 2175
rect 649 2154 659 2168
rect 906 2154 915 2168
rect 649 2148 678 2154
rect 728 2148 757 2154
rect 807 2148 836 2154
rect 886 2148 915 2154
rect 648 2147 679 2148
rect 727 2147 758 2148
rect 806 2147 837 2148
rect 885 2147 916 2148
rect 948 2147 965 2176
rect 1190 2155 1196 2161
rect 2052 2155 2058 2161
rect 649 2146 650 2147
rect 677 2146 678 2147
rect 728 2146 729 2147
rect 756 2146 757 2147
rect 807 2146 808 2147
rect 835 2146 836 2147
rect 886 2146 887 2147
rect 914 2146 915 2147
rect 4358 2125 4364 2131
rect 4463 2125 4469 2131
rect 4784 2115 4790 2121
rect 4837 2115 4843 2121
rect 649 2097 678 2112
rect 728 2097 757 2112
rect 807 2097 836 2112
rect 886 2097 915 2112
rect 4352 2061 4358 2067
rect 4469 2061 4475 2067
rect 4778 2065 4784 2071
rect 4843 2065 4849 2071
rect 4358 2008 4364 2014
rect 4463 2008 4469 2014
rect 4784 2006 4790 2012
rect 4837 2006 4843 2012
rect 4778 1956 4784 1962
rect 4843 1956 4849 1962
rect 4352 1944 4358 1950
rect 4469 1944 4475 1950
rect 4358 1823 4364 1829
rect 4463 1823 4469 1829
rect 4621 1818 4638 1822
rect 4784 1817 4790 1823
rect 4837 1817 4843 1823
rect 4778 1767 4784 1773
rect 4843 1767 4849 1773
rect 4352 1759 4358 1765
rect 4469 1759 4475 1765
rect 4358 1707 4364 1713
rect 4463 1707 4469 1713
rect 4784 1700 4790 1706
rect 4837 1700 4843 1706
rect 4778 1650 4784 1656
rect 4843 1650 4849 1656
rect 4352 1643 4358 1649
rect 4469 1643 4475 1649
rect 6228 1325 6230 1326
rect 519 1156 536 1159
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_0
timestamp 1625405207
transform 1 0 -1050 0 1 -5
box 1050 5 1614 610
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_0
timestamp 1624113741
transform 1 0 714 0 1 211
box -30 -102 850 522
use sky130_hilas_Trans4small  sky130_hilas_Trans4small_0
timestamp 1608234847
transform 1 0 -729 0 1 934
box 191 -150 471 438
use sky130_hilas_Trans2med  sky130_hilas_Trans2med_0
timestamp 1625425852
transform 1 0 587 0 1 1190
box -380 -143 -27 452
use sky130_hilas_nFETLarge  sky130_hilas_nFETLarge_0
timestamp 1625426387
transform 1 0 789 0 1 586
box 64 420 501 1003
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_0
timestamp 1608245216
transform 1 0 1645 0 1 508
box 64 419 528 1018
use sky130_hilas_WTA4Stage01  sky130_hilas_WTA4Stage01_0
timestamp 1625404155
transform 1 0 4954 0 1 1626
box -1121 -43 296 562
use sky130_hilas_FGcharacterization01  sky130_hilas_FGcharacterization01_0
timestamp 1625074044
transform 1 0 597 0 1 1820
box -912 259 2083 864
use sky130_hilas_swc4x2cell  sky130_hilas_swc4x2cell_0
timestamp 1625491916
transform 1 0 4087 0 1 2720
box -1004 -4 1009 601
use sky130_hilas_TA2Cell_1FG_Strong  sky130_hilas_TA2Cell_1FG_Strong_0
timestamp 1625491312
transform 1 0 4496 0 1 3369
box -2617 140 193 745
use sky130_hilas_DAC5bit01  sky130_hilas_DAC5bit01_0
timestamp 1625056879
transform 1 0 5165 0 1 436
box 382 524 2040 1121
use sky130_hilas_Tgate4Single01  sky130_hilas_Tgate4Single01_0
timestamp 1608226321
transform 1 0 5682 0 1 3791
box -36 -141 440 464
use sky130_hilas_TA2Cell_1FG  sky130_hilas_TA2Cell_1FG_0
timestamp 1625491133
transform 1 0 8403 0 1 2519
box -2616 140 193 745
<< end >>
