magic
tech sky130A
timestamp 1628704370
<< error_s >>
rect 65 135 115 141
rect 388 136 438 142
rect 545 135 573 142
rect 687 136 715 142
rect 65 93 115 99
rect 388 94 438 100
rect 545 93 573 100
rect 687 94 715 100
rect 136 69 186 75
rect 316 64 367 70
rect 496 64 524 70
rect 736 64 764 70
rect 136 27 186 33
rect 316 22 367 28
rect 496 22 524 28
rect 736 22 764 28
<< nwell >>
rect 0 0 250 175
rect 637 168 814 175
rect 637 0 814 9
<< mvpmos >>
rect 65 99 115 135
rect 136 33 186 69
<< mvpdiff >>
rect 34 123 65 135
rect 34 106 42 123
rect 59 106 65 123
rect 34 99 65 106
rect 115 124 149 135
rect 115 107 121 124
rect 138 107 149 124
rect 115 99 149 107
rect 105 60 136 69
rect 105 43 111 60
rect 129 43 136 60
rect 105 33 136 43
rect 186 62 217 69
rect 186 45 192 62
rect 210 45 217 62
rect 186 33 217 45
<< mvpdiffc >>
rect 42 106 59 123
rect 121 107 138 124
rect 111 43 129 60
rect 192 45 210 62
<< mvnsubdiff >>
rect 35 60 105 69
rect 35 43 61 60
rect 78 43 105 60
rect 35 33 105 43
<< mvnsubdiffcont >>
rect 61 43 78 60
<< poly >>
rect 65 143 215 158
rect 65 135 115 143
rect 188 131 215 143
rect 188 114 193 131
rect 210 114 215 131
rect 188 104 215 114
rect 242 129 276 134
rect 242 112 251 129
rect 268 112 276 129
rect 242 104 276 112
rect 65 84 115 99
rect 136 69 186 83
rect 242 70 258 104
rect 226 46 258 70
rect 136 25 186 33
rect 226 25 242 46
rect 136 10 242 25
<< polycont >>
rect 193 114 210 131
rect 251 112 268 129
<< locali >>
rect 128 131 173 139
rect 128 124 145 131
rect 34 106 42 123
rect 59 106 67 123
rect 113 107 121 124
rect 138 114 145 124
rect 162 114 173 131
rect 138 107 173 114
rect 193 131 210 139
rect 41 97 59 106
rect 58 80 59 97
rect 41 61 59 80
rect 193 63 210 114
rect 243 129 272 132
rect 243 127 251 129
rect 243 110 249 127
rect 268 112 276 129
rect 266 110 272 112
rect 243 108 272 110
rect 193 62 231 63
rect 58 60 59 61
rect 58 44 61 60
rect 41 43 61 44
rect 78 43 111 60
rect 129 43 137 60
rect 184 45 192 62
rect 210 56 231 62
rect 210 51 265 56
rect 210 45 266 51
rect 192 39 266 45
rect 192 34 231 39
<< viali >>
rect 145 114 162 131
rect 41 80 58 97
rect 249 112 251 127
rect 251 112 266 127
rect 249 110 266 112
rect 41 44 58 61
<< metal1 >>
rect 34 97 63 175
rect 465 169 496 175
rect 766 168 790 175
rect 138 136 170 139
rect 138 110 141 136
rect 167 110 170 136
rect 243 132 274 133
rect 138 109 170 110
rect 242 106 245 132
rect 271 106 274 132
rect 242 105 274 106
rect 243 104 272 105
rect 34 80 41 97
rect 58 80 63 97
rect 34 61 63 80
rect 34 44 41 61
rect 58 44 63 61
rect 34 0 63 44
<< via1 >>
rect 141 131 167 136
rect 141 114 145 131
rect 145 114 162 131
rect 162 114 167 131
rect 141 110 167 114
rect 245 127 271 132
rect 245 110 249 127
rect 249 110 266 127
rect 266 110 271 127
rect 245 106 271 110
<< metal2 >>
rect 138 131 141 136
rect 7 111 141 131
rect 138 110 141 111
rect 167 131 170 136
rect 241 132 273 133
rect 241 131 245 132
rect 167 111 245 131
rect 167 110 170 111
rect 241 106 245 111
rect 271 106 274 132
rect 241 104 273 106
use sky130_hilas_StepUpDigitalPart1  StepUpDigitalPart1_0
timestamp 1628704340
transform 1 0 -22 0 1 49
box 0 0 614 169
<< labels >>
rlabel metal2 7 111 14 131 0 Output
rlabel metal1 34 155 63 163 0 Vinj
rlabel metal1 34 4 63 12 0 Vinj
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
