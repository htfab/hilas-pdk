magic
tech sky130A
timestamp 1632575814
<< nwell >>
rect 633 -163 861 0
rect 633 -415 803 -163
rect 632 -617 803 -415
<< nmos >>
rect -437 -281 -422 -18
rect -437 -612 -422 -349
rect -335 -614 -315 -18
rect -282 -614 -262 -18
rect -231 -614 -211 -18
rect -180 -614 -160 -18
rect -129 -614 -109 -18
rect -78 -614 -58 -18
rect -27 -614 -7 -18
rect 24 -614 44 -18
rect 75 -614 95 -18
rect 126 -614 146 -18
rect 177 -614 197 -18
rect 228 -614 248 -18
rect 279 -614 299 -18
rect 330 -614 350 -18
rect 381 -614 401 -18
rect 432 -614 452 -18
rect 541 -218 561 -18
<< pmos >>
rect 683 -599 703 -18
rect 735 -599 755 -18
<< ndiff >>
rect -465 -30 -437 -18
rect -465 -273 -461 -30
rect -444 -273 -437 -30
rect -465 -281 -437 -273
rect -422 -32 -394 -18
rect -422 -275 -416 -32
rect -399 -275 -394 -32
rect -422 -281 -394 -275
rect -414 -349 -394 -281
rect -466 -360 -437 -349
rect -466 -605 -461 -360
rect -444 -605 -437 -360
rect -466 -612 -437 -605
rect -422 -361 -394 -349
rect -422 -606 -416 -361
rect -399 -606 -394 -361
rect -422 -612 -394 -606
rect -364 -26 -335 -18
rect -364 -610 -358 -26
rect -341 -610 -335 -26
rect -364 -614 -335 -610
rect -315 -26 -282 -18
rect -315 -610 -307 -26
rect -290 -610 -282 -26
rect -315 -614 -282 -610
rect -262 -26 -231 -18
rect -262 -610 -256 -26
rect -239 -610 -231 -26
rect -262 -614 -231 -610
rect -211 -26 -180 -18
rect -211 -610 -204 -26
rect -187 -610 -180 -26
rect -211 -614 -180 -610
rect -160 -26 -129 -18
rect -160 -610 -154 -26
rect -137 -610 -129 -26
rect -160 -614 -129 -610
rect -109 -26 -78 -18
rect -109 -610 -103 -26
rect -86 -610 -78 -26
rect -109 -614 -78 -610
rect -58 -26 -27 -18
rect -58 -610 -51 -26
rect -34 -610 -27 -26
rect -58 -614 -27 -610
rect -7 -26 24 -18
rect -7 -610 0 -26
rect 17 -610 24 -26
rect -7 -614 24 -610
rect 44 -26 75 -18
rect 44 -610 51 -26
rect 68 -610 75 -26
rect 44 -614 75 -610
rect 95 -26 126 -18
rect 95 -610 102 -26
rect 119 -610 126 -26
rect 95 -614 126 -610
rect 146 -26 177 -18
rect 146 -610 153 -26
rect 170 -610 177 -26
rect 146 -614 177 -610
rect 197 -26 228 -18
rect 197 -610 203 -26
rect 220 -610 228 -26
rect 197 -614 228 -610
rect 248 -26 279 -18
rect 248 -610 255 -26
rect 272 -610 279 -26
rect 248 -614 279 -610
rect 299 -26 330 -18
rect 299 -610 305 -26
rect 322 -610 330 -26
rect 299 -614 330 -610
rect 350 -26 381 -18
rect 350 -610 356 -26
rect 373 -610 381 -26
rect 350 -614 381 -610
rect 401 -26 432 -18
rect 401 -610 408 -26
rect 425 -610 432 -26
rect 401 -614 432 -610
rect 452 -26 483 -18
rect 452 -610 458 -26
rect 475 -610 483 -26
rect 510 -27 541 -18
rect 510 -210 517 -27
rect 534 -210 541 -27
rect 510 -218 541 -210
rect 561 -27 592 -18
rect 561 -210 568 -27
rect 585 -210 592 -27
rect 561 -218 592 -210
rect 452 -614 483 -610
<< pdiff >>
rect 653 -39 683 -18
rect 653 -589 660 -39
rect 677 -589 683 -39
rect 653 -599 683 -589
rect 703 -39 735 -18
rect 703 -588 710 -39
rect 727 -588 735 -39
rect 703 -599 735 -588
rect 755 -40 784 -18
rect 755 -588 761 -40
rect 778 -588 784 -40
rect 755 -599 784 -588
<< ndiffc >>
rect -461 -273 -444 -30
rect -416 -275 -399 -32
rect -461 -605 -444 -360
rect -416 -606 -399 -361
rect -358 -610 -341 -26
rect -307 -610 -290 -26
rect -256 -610 -239 -26
rect -204 -610 -187 -26
rect -154 -610 -137 -26
rect -103 -610 -86 -26
rect -51 -610 -34 -26
rect 0 -610 17 -26
rect 51 -610 68 -26
rect 102 -610 119 -26
rect 153 -610 170 -26
rect 203 -610 220 -26
rect 255 -610 272 -26
rect 305 -610 322 -26
rect 356 -610 373 -26
rect 408 -610 425 -26
rect 458 -610 475 -26
rect 517 -210 534 -27
rect 568 -210 585 -27
<< pdiffc >>
rect 660 -589 677 -39
rect 710 -588 727 -39
rect 761 -588 778 -40
<< psubdiff >>
rect 511 -258 587 -246
rect 511 -603 522 -258
rect 578 -603 587 -258
rect 511 -615 587 -603
<< nsubdiff >>
rect 811 -39 843 -19
rect 811 -119 818 -39
rect 835 -119 843 -39
rect 811 -132 843 -119
<< psubdiffcont >>
rect 522 -603 578 -258
<< nsubdiffcont >>
rect 818 -119 835 -39
<< poly >>
rect -437 -10 633 5
rect -437 -18 -422 -10
rect -335 -18 -315 -10
rect -282 -18 -262 -10
rect -231 -18 -211 -10
rect -180 -18 -160 -10
rect -129 -18 -109 -10
rect -78 -18 -58 -10
rect -27 -18 -7 -10
rect 24 -18 44 -10
rect 75 -18 95 -10
rect 126 -18 146 -10
rect 177 -18 197 -10
rect 228 -18 248 -10
rect 279 -18 299 -10
rect 330 -18 350 -10
rect 381 -18 401 -10
rect 432 -18 452 -10
rect 541 -18 561 -10
rect -940 -35 -889 -20
rect -940 -541 -925 -35
rect -958 -546 -925 -541
rect -958 -563 -950 -546
rect -933 -563 -925 -546
rect -958 -568 -925 -563
rect -904 -579 -889 -35
rect -868 -35 -817 -20
rect -868 -579 -853 -35
rect -904 -595 -853 -579
rect -832 -579 -817 -35
rect -796 -35 -745 -20
rect -796 -579 -781 -35
rect -832 -595 -781 -579
rect -760 -579 -745 -35
rect -724 -35 -673 -20
rect -724 -579 -709 -35
rect -760 -595 -709 -579
rect -688 -579 -673 -35
rect -652 -35 -601 -20
rect -652 -579 -637 -35
rect -688 -595 -637 -579
rect -616 -579 -601 -35
rect -580 -35 -529 -20
rect -580 -579 -565 -35
rect -616 -595 -565 -579
rect -544 -579 -529 -35
rect -437 -294 -422 -281
rect -492 -313 -458 -308
rect -492 -330 -484 -313
rect -467 -326 -458 -313
rect -467 -330 -422 -326
rect -492 -341 -422 -330
rect -437 -349 -422 -341
rect -508 -443 -477 -434
rect -508 -460 -503 -443
rect -486 -460 -477 -443
rect -508 -469 -477 -460
rect -506 -579 -491 -469
rect -544 -595 -491 -579
rect -437 -625 -422 -612
rect 602 -26 633 -10
rect 683 -18 703 -5
rect 735 -18 755 -5
rect 602 -209 611 -26
rect 628 -209 633 -26
rect 602 -217 633 -209
rect 541 -231 561 -218
rect -335 -627 -315 -614
rect -282 -627 -262 -614
rect -231 -627 -211 -614
rect -180 -627 -160 -614
rect -129 -627 -109 -614
rect -78 -627 -58 -614
rect -27 -627 -7 -614
rect 24 -627 44 -614
rect 75 -627 95 -614
rect 126 -627 146 -614
rect 177 -627 197 -614
rect 228 -627 248 -614
rect 279 -627 299 -614
rect 330 -627 350 -614
rect 381 -627 401 -614
rect 432 -627 452 -614
rect 607 -364 643 -353
rect 607 -589 612 -364
rect 629 -589 643 -364
rect 607 -607 643 -589
rect 683 -607 703 -599
rect 735 -607 755 -599
rect 607 -622 755 -607
<< polycont >>
rect -950 -563 -933 -546
rect -484 -330 -467 -313
rect -503 -460 -486 -443
rect 611 -209 628 -26
rect 612 -589 629 -364
<< locali >>
rect -461 -30 -444 -22
rect -468 -149 -461 -143
rect -468 -159 -462 -149
rect -484 -166 -462 -159
rect -484 -185 -461 -166
rect -484 -202 -462 -185
rect -484 -221 -461 -202
rect -484 -238 -462 -221
rect -484 -253 -461 -238
rect -503 -257 -461 -253
rect -503 -274 -500 -257
rect -483 -274 -463 -257
rect -446 -274 -444 -273
rect -503 -280 -444 -274
rect -416 -32 -399 -16
rect -503 -293 -442 -280
rect -503 -296 -500 -293
rect -502 -310 -500 -296
rect -483 -310 -462 -293
rect -445 -310 -442 -293
rect -502 -311 -442 -310
rect -492 -313 -442 -311
rect -492 -330 -484 -313
rect -467 -316 -442 -313
rect -467 -330 -459 -316
rect -461 -360 -444 -352
rect -503 -442 -486 -435
rect -503 -443 -501 -442
rect -503 -468 -486 -460
rect -416 -361 -399 -275
rect -960 -546 -924 -543
rect -960 -547 -950 -546
rect -960 -564 -951 -547
rect -933 -563 -924 -546
rect -934 -564 -924 -563
rect -960 -566 -924 -564
rect -461 -613 -444 -605
rect -417 -606 -416 -468
rect -360 -26 -339 -18
rect -360 -442 -358 -26
rect -360 -459 -359 -442
rect -417 -608 -415 -606
rect -417 -617 -399 -608
rect -360 -610 -358 -459
rect -341 -610 -339 -26
rect -360 -618 -339 -610
rect -309 -26 -288 -18
rect -309 -610 -307 -26
rect -290 -544 -288 -26
rect -289 -561 -288 -544
rect -290 -610 -288 -561
rect -309 -618 -288 -610
rect -258 -26 -237 -18
rect -258 -441 -256 -26
rect -258 -458 -257 -441
rect -258 -610 -256 -458
rect -239 -610 -237 -26
rect -258 -618 -237 -610
rect -206 -26 -185 -18
rect -206 -610 -204 -26
rect -187 -544 -185 -26
rect -186 -561 -185 -544
rect -187 -610 -185 -561
rect -206 -618 -185 -610
rect -156 -26 -135 -18
rect -156 -441 -154 -26
rect -156 -458 -155 -441
rect -156 -610 -154 -458
rect -137 -610 -135 -26
rect -156 -618 -135 -610
rect -105 -26 -84 -16
rect -105 -610 -103 -26
rect -86 -544 -84 -26
rect -85 -561 -84 -544
rect -86 -610 -84 -561
rect -105 -618 -84 -610
rect -53 -26 -32 -16
rect -53 -441 -51 -26
rect -53 -458 -52 -441
rect -53 -610 -51 -458
rect -34 -610 -32 -26
rect -53 -618 -32 -610
rect -2 -26 19 -16
rect -2 -610 0 -26
rect 17 -34 19 -26
rect 49 -26 70 -16
rect 17 -544 18 -34
rect 17 -610 18 -561
rect -2 -618 18 -610
rect 49 -441 51 -26
rect 68 -34 70 -26
rect 100 -26 121 -16
rect 49 -458 50 -441
rect 49 -610 51 -458
rect 68 -610 69 -34
rect 49 -618 69 -610
rect 100 -610 102 -26
rect 119 -34 121 -26
rect 151 -26 172 -16
rect 119 -544 120 -34
rect 119 -610 120 -561
rect 100 -618 120 -610
rect 151 -441 153 -26
rect 151 -458 152 -441
rect 151 -610 153 -458
rect 170 -610 172 -26
rect 151 -618 172 -610
rect 201 -26 222 -16
rect 201 -610 203 -26
rect 220 -544 222 -26
rect 221 -561 222 -544
rect 220 -610 222 -561
rect 201 -618 222 -610
rect 253 -26 274 -16
rect 253 -441 255 -26
rect 253 -458 254 -441
rect 253 -610 255 -458
rect 272 -610 274 -26
rect 253 -618 274 -610
rect 303 -26 324 -16
rect 303 -610 305 -26
rect 322 -544 324 -26
rect 323 -561 324 -544
rect 322 -610 324 -561
rect 303 -618 324 -610
rect 354 -26 375 -16
rect 354 -441 356 -26
rect 354 -458 355 -441
rect 354 -610 356 -458
rect 373 -610 375 -26
rect 354 -618 375 -610
rect 406 -26 427 -16
rect 406 -610 408 -26
rect 425 -543 427 -26
rect 426 -560 427 -543
rect 425 -610 427 -560
rect 406 -618 427 -610
rect 456 -26 477 -16
rect 456 -441 458 -26
rect 456 -458 457 -441
rect 456 -610 458 -458
rect 475 -610 477 -26
rect 514 -27 538 -16
rect 514 -210 517 -27
rect 534 -210 538 -27
rect 514 -245 538 -210
rect 566 -26 632 -17
rect 566 -27 611 -26
rect 566 -210 568 -27
rect 585 -118 611 -27
rect 587 -135 611 -118
rect 628 -119 632 -26
rect 585 -155 611 -135
rect 630 -136 632 -119
rect 628 -155 632 -136
rect 587 -172 611 -155
rect 630 -172 632 -155
rect 585 -193 611 -172
rect 628 -192 632 -172
rect 586 -209 611 -193
rect 629 -209 632 -192
rect 586 -210 632 -209
rect 566 -221 632 -210
rect 658 -39 679 -31
rect 456 -618 477 -610
rect 512 -251 579 -245
rect 512 -258 540 -251
rect 557 -258 579 -251
rect 512 -603 522 -258
rect 578 -603 579 -258
rect 658 -354 660 -39
rect 610 -364 660 -354
rect 610 -589 612 -364
rect 629 -540 660 -364
rect 629 -557 639 -540
rect 656 -557 660 -540
rect 629 -589 660 -557
rect 677 -589 679 -39
rect 610 -597 679 -589
rect 708 -39 729 -31
rect 708 -41 710 -39
rect 708 -58 709 -41
rect 708 -78 710 -58
rect 708 -95 709 -78
rect 708 -588 710 -95
rect 727 -588 729 -39
rect 708 -597 729 -588
rect 759 -40 780 -31
rect 818 -38 835 -31
rect 759 -118 761 -40
rect 759 -135 760 -118
rect 759 -155 761 -135
rect 759 -172 760 -155
rect 759 -191 761 -172
rect 759 -208 760 -191
rect 759 -588 761 -208
rect 778 -588 780 -40
rect 834 -39 835 -38
rect 818 -132 835 -119
rect 759 -597 780 -588
rect 512 -612 579 -603
<< viali >>
rect -462 -166 -461 -149
rect -461 -166 -445 -149
rect -462 -202 -461 -185
rect -461 -202 -445 -185
rect -462 -238 -461 -221
rect -461 -238 -445 -221
rect -500 -274 -483 -257
rect -463 -273 -461 -257
rect -461 -273 -446 -257
rect -463 -274 -446 -273
rect -500 -310 -483 -293
rect -462 -310 -445 -293
rect -501 -443 -484 -442
rect -501 -459 -486 -443
rect -486 -459 -484 -443
rect -462 -538 -461 -521
rect -461 -538 -445 -521
rect -951 -563 -950 -547
rect -950 -563 -934 -547
rect -951 -564 -934 -563
rect -462 -575 -461 -558
rect -461 -575 -445 -558
rect -359 -459 -358 -442
rect -358 -459 -342 -442
rect -414 -536 -399 -519
rect -399 -536 -397 -519
rect -415 -572 -399 -555
rect -399 -572 -398 -555
rect -415 -606 -399 -591
rect -399 -606 -398 -591
rect -415 -608 -398 -606
rect -306 -561 -290 -544
rect -290 -561 -289 -544
rect -257 -458 -256 -441
rect -256 -458 -240 -441
rect -203 -561 -187 -544
rect -187 -561 -186 -544
rect -155 -458 -154 -441
rect -154 -458 -138 -441
rect -102 -561 -86 -544
rect -86 -561 -85 -544
rect -52 -458 -51 -441
rect -51 -458 -35 -441
rect 1 -561 17 -544
rect 17 -561 18 -544
rect 50 -458 51 -441
rect 51 -458 67 -441
rect 103 -561 119 -544
rect 119 -561 120 -544
rect 152 -458 153 -441
rect 153 -458 169 -441
rect 204 -561 220 -544
rect 220 -561 221 -544
rect 254 -458 255 -441
rect 255 -458 271 -441
rect 306 -561 322 -544
rect 322 -561 323 -544
rect 355 -458 356 -441
rect 356 -458 372 -441
rect 409 -560 425 -543
rect 425 -560 426 -543
rect 457 -458 458 -441
rect 458 -458 474 -441
rect 569 -135 585 -118
rect 585 -135 587 -118
rect 612 -136 628 -119
rect 628 -136 630 -119
rect 569 -172 585 -155
rect 585 -172 587 -155
rect 612 -172 628 -155
rect 628 -172 630 -155
rect 569 -210 585 -193
rect 585 -210 586 -193
rect 612 -209 628 -192
rect 628 -209 629 -192
rect 540 -258 557 -251
rect 540 -268 557 -258
rect 540 -304 557 -287
rect 540 -340 557 -323
rect 540 -376 557 -359
rect 540 -412 557 -395
rect 540 -448 557 -431
rect 540 -484 557 -467
rect 540 -520 557 -503
rect 540 -556 557 -539
rect 540 -592 557 -575
rect 639 -557 656 -540
rect 709 -58 710 -41
rect 710 -58 726 -41
rect 709 -95 710 -78
rect 710 -95 726 -78
rect 760 -135 761 -118
rect 761 -135 778 -118
rect 760 -172 761 -155
rect 761 -172 778 -155
rect 760 -208 761 -191
rect 761 -208 778 -191
rect 817 -39 834 -38
rect 817 -55 818 -39
rect 818 -55 834 -39
rect 817 -94 818 -77
rect 818 -94 834 -77
<< metal1 >>
rect 702 13 734 14
rect 702 -13 705 13
rect 731 -13 734 13
rect 702 -18 734 -13
rect 810 13 843 14
rect 810 -13 813 13
rect 839 -13 843 13
rect 706 -41 729 -18
rect 810 -19 843 -13
rect 706 -58 709 -41
rect 726 -58 729 -41
rect 706 -78 729 -58
rect 706 -95 709 -78
rect 726 -95 729 -78
rect 706 -101 729 -95
rect 814 -38 837 -19
rect 814 -55 817 -38
rect 834 -55 837 -38
rect 814 -77 837 -55
rect 814 -94 817 -77
rect 834 -94 837 -77
rect 814 -100 837 -94
rect 564 -116 595 -112
rect 749 -116 782 -112
rect 564 -118 782 -116
rect 564 -135 569 -118
rect 587 -119 760 -118
rect 587 -135 612 -119
rect 564 -136 612 -135
rect 630 -135 760 -119
rect 778 -135 782 -118
rect 630 -136 782 -135
rect -466 -149 -442 -143
rect -466 -166 -462 -149
rect -445 -166 -442 -149
rect -466 -185 -442 -166
rect -466 -202 -462 -185
rect -445 -202 -442 -185
rect -466 -221 -442 -202
rect 564 -155 781 -136
rect 564 -172 569 -155
rect 587 -172 612 -155
rect 630 -172 760 -155
rect 778 -172 781 -155
rect 564 -173 781 -172
rect 564 -193 584 -173
rect 610 -183 781 -173
rect 610 -191 782 -183
rect 610 -192 760 -191
rect 564 -210 569 -193
rect 610 -199 612 -192
rect 586 -209 612 -199
rect 629 -208 760 -192
rect 778 -208 782 -191
rect 629 -209 782 -208
rect 586 -210 782 -209
rect 564 -216 782 -210
rect -466 -238 -462 -221
rect -445 -238 -442 -221
rect -492 -251 -442 -238
rect -503 -257 -442 -251
rect -503 -274 -500 -257
rect -483 -274 -463 -257
rect -446 -274 -442 -257
rect -503 -281 -442 -274
rect -503 -293 -489 -281
rect -463 -293 -442 -281
rect -503 -310 -500 -293
rect -463 -307 -462 -293
rect -483 -310 -462 -307
rect -445 -310 -442 -293
rect -503 -313 -442 -310
rect -503 -316 -480 -313
rect -466 -316 -442 -313
rect 523 -251 571 -244
rect 523 -268 540 -251
rect 557 -268 571 -251
rect 523 -287 571 -268
rect 523 -304 540 -287
rect 557 -304 571 -287
rect 523 -323 571 -304
rect 523 -340 540 -323
rect 557 -340 571 -323
rect 523 -359 571 -340
rect 523 -376 540 -359
rect 557 -376 571 -359
rect 523 -395 571 -376
rect 523 -412 540 -395
rect 557 -412 571 -395
rect 523 -431 571 -412
rect -506 -437 487 -434
rect -506 -438 -158 -437
rect -506 -442 -260 -438
rect -506 -459 -501 -442
rect -484 -459 -359 -442
rect -342 -459 -260 -442
rect -506 -464 -260 -459
rect -234 -463 -158 -438
rect -132 -463 -56 -437
rect -30 -463 46 -437
rect 72 -463 149 -437
rect 175 -463 250 -437
rect 276 -463 352 -437
rect 378 -463 454 -437
rect 480 -463 487 -437
rect -234 -464 487 -463
rect -506 -468 487 -464
rect 523 -448 540 -431
rect 557 -448 571 -431
rect 523 -467 571 -448
rect 523 -484 540 -467
rect 557 -484 571 -467
rect 523 -503 571 -484
rect -465 -521 -440 -515
rect -465 -536 -462 -521
rect -469 -538 -462 -536
rect -445 -536 -440 -521
rect -417 -519 -390 -512
rect -417 -536 -414 -519
rect -397 -536 -390 -519
rect 523 -520 540 -503
rect 557 -520 571 -503
rect -179 -536 432 -535
rect -445 -538 -439 -536
rect -469 -539 -439 -538
rect -962 -541 -924 -539
rect -962 -567 -956 -541
rect -930 -567 -924 -541
rect -962 -570 -924 -567
rect -469 -565 -466 -539
rect -440 -565 -439 -539
rect -417 -547 -390 -536
rect -469 -568 -462 -565
rect -465 -575 -462 -568
rect -445 -568 -439 -565
rect -423 -555 -390 -547
rect -445 -575 -440 -568
rect -465 -581 -440 -575
rect -423 -572 -415 -555
rect -398 -572 -390 -555
rect -315 -538 432 -536
rect -315 -539 -107 -538
rect -315 -565 -312 -539
rect -286 -565 -208 -539
rect -182 -564 -107 -539
rect -81 -564 -5 -538
rect 21 -564 98 -538
rect 124 -564 200 -538
rect 226 -564 302 -538
rect 328 -564 404 -538
rect 430 -564 432 -538
rect -182 -565 432 -564
rect -315 -568 432 -565
rect 523 -539 571 -520
rect 523 -556 540 -539
rect 557 -556 571 -539
rect 523 -561 571 -556
rect 627 -535 669 -526
rect 627 -561 635 -535
rect 661 -561 669 -535
rect -315 -569 -282 -568
rect -423 -591 -390 -572
rect -423 -596 -415 -591
rect -398 -596 -390 -591
rect -423 -622 -419 -596
rect -393 -622 -390 -596
rect -423 -626 -390 -622
rect 523 -575 577 -561
rect 627 -568 669 -561
rect 523 -592 540 -575
rect 557 -592 577 -575
rect 523 -599 577 -592
rect 523 -625 535 -599
rect 561 -625 577 -599
rect 523 -628 577 -625
<< via1 >>
rect 705 -13 731 13
rect 813 -13 839 13
rect 584 -193 610 -173
rect 584 -199 586 -193
rect 586 -199 610 -193
rect -489 -293 -463 -281
rect -489 -307 -483 -293
rect -483 -307 -463 -293
rect -260 -441 -234 -438
rect -260 -458 -257 -441
rect -257 -458 -240 -441
rect -240 -458 -234 -441
rect -260 -464 -234 -458
rect -158 -441 -132 -437
rect -158 -458 -155 -441
rect -155 -458 -138 -441
rect -138 -458 -132 -441
rect -158 -463 -132 -458
rect -56 -441 -30 -437
rect -56 -458 -52 -441
rect -52 -458 -35 -441
rect -35 -458 -30 -441
rect -56 -463 -30 -458
rect 46 -441 72 -437
rect 46 -458 50 -441
rect 50 -458 67 -441
rect 67 -458 72 -441
rect 46 -463 72 -458
rect 149 -441 175 -437
rect 149 -458 152 -441
rect 152 -458 169 -441
rect 169 -458 175 -441
rect 149 -463 175 -458
rect 250 -441 276 -437
rect 250 -458 254 -441
rect 254 -458 271 -441
rect 271 -458 276 -441
rect 250 -463 276 -458
rect 352 -441 378 -437
rect 352 -458 355 -441
rect 355 -458 372 -441
rect 372 -458 378 -441
rect 352 -463 378 -458
rect 454 -441 480 -437
rect 454 -458 457 -441
rect 457 -458 474 -441
rect 474 -458 480 -441
rect 454 -463 480 -458
rect -956 -547 -930 -541
rect -956 -564 -951 -547
rect -951 -564 -934 -547
rect -934 -564 -930 -547
rect -956 -567 -930 -564
rect -466 -558 -440 -539
rect -466 -565 -462 -558
rect -462 -565 -445 -558
rect -445 -565 -440 -558
rect -312 -544 -286 -539
rect -312 -561 -306 -544
rect -306 -561 -289 -544
rect -289 -561 -286 -544
rect -312 -565 -286 -561
rect -208 -544 -182 -539
rect -208 -561 -203 -544
rect -203 -561 -186 -544
rect -186 -561 -182 -544
rect -208 -565 -182 -561
rect -107 -544 -81 -538
rect -107 -561 -102 -544
rect -102 -561 -85 -544
rect -85 -561 -81 -544
rect -107 -564 -81 -561
rect -5 -544 21 -538
rect -5 -561 1 -544
rect 1 -561 18 -544
rect 18 -561 21 -544
rect -5 -564 21 -561
rect 98 -544 124 -538
rect 98 -561 103 -544
rect 103 -561 120 -544
rect 120 -561 124 -544
rect 98 -564 124 -561
rect 200 -544 226 -538
rect 200 -561 204 -544
rect 204 -561 221 -544
rect 221 -561 226 -544
rect 200 -564 226 -561
rect 302 -544 328 -538
rect 302 -561 306 -544
rect 306 -561 323 -544
rect 323 -561 328 -544
rect 302 -564 328 -561
rect 404 -543 430 -538
rect 404 -560 409 -543
rect 409 -560 426 -543
rect 426 -560 430 -543
rect 404 -564 430 -560
rect 635 -540 661 -535
rect 635 -557 639 -540
rect 639 -557 656 -540
rect 656 -557 661 -540
rect 635 -561 661 -557
rect -419 -608 -415 -596
rect -415 -608 -398 -596
rect -398 -608 -393 -596
rect -419 -622 -393 -608
rect 535 -625 561 -599
<< metal2 >>
rect -984 13 924 17
rect -984 9 705 13
rect -984 -20 -915 9
rect -812 -13 705 9
rect 731 -13 813 13
rect 839 -13 924 13
rect -812 -20 924 -13
rect -984 -21 924 -20
rect -920 -23 -807 -21
rect 864 -75 924 -49
rect 864 -139 924 -113
rect 570 -173 624 -166
rect 570 -199 584 -173
rect 610 -199 924 -173
rect 570 -206 624 -199
rect 864 -253 924 -227
rect -501 -279 -442 -277
rect -501 -309 -493 -279
rect -458 -281 -442 -279
rect -458 -307 -434 -281
rect 861 -307 924 -281
rect -458 -309 -442 -307
rect -501 -312 -442 -309
rect 864 -359 924 -333
rect 864 -411 924 -385
rect -162 -437 -128 -433
rect -59 -437 -25 -433
rect 42 -437 76 -433
rect 145 -437 179 -433
rect 247 -437 281 -433
rect 348 -437 382 -433
rect 449 -437 483 -433
rect -375 -438 -158 -437
rect -375 -463 -260 -438
rect -263 -464 -260 -463
rect -234 -463 -158 -438
rect -132 -463 -56 -437
rect -30 -463 46 -437
rect 72 -463 149 -437
rect 175 -463 250 -437
rect 276 -463 352 -437
rect 378 -463 454 -437
rect 480 -463 483 -437
rect 861 -463 924 -437
rect -234 -464 -232 -463
rect -263 -467 -232 -464
rect -162 -469 -128 -463
rect -59 -469 -25 -463
rect 42 -469 76 -463
rect 145 -469 179 -463
rect 247 -469 281 -463
rect 348 -469 382 -463
rect 449 -469 483 -463
rect 864 -515 924 -489
rect 629 -535 667 -527
rect -470 -539 -438 -536
rect -961 -541 -925 -540
rect -470 -541 -466 -539
rect -984 -567 -956 -541
rect -930 -567 -925 -541
rect -472 -565 -466 -541
rect -440 -541 -438 -539
rect -315 -539 -283 -536
rect -315 -541 -312 -539
rect -440 -565 -312 -541
rect -286 -541 -283 -539
rect -211 -539 -179 -536
rect -211 -541 -208 -539
rect -286 -565 -208 -541
rect -182 -541 -179 -539
rect -109 -538 -78 -535
rect -109 -541 -107 -538
rect -182 -564 -107 -541
rect -81 -541 -78 -538
rect -7 -538 24 -535
rect -7 -541 -5 -538
rect -81 -564 -5 -541
rect 21 -541 24 -538
rect 95 -538 126 -535
rect 95 -541 98 -538
rect 21 -564 98 -541
rect 124 -541 126 -538
rect 197 -538 229 -535
rect 197 -541 200 -538
rect 124 -564 200 -541
rect 226 -541 229 -538
rect 299 -538 330 -535
rect 299 -541 302 -538
rect 226 -564 302 -541
rect 328 -541 330 -538
rect 401 -538 432 -535
rect 401 -541 404 -538
rect 328 -564 404 -541
rect 430 -541 432 -538
rect 629 -541 635 -535
rect 430 -561 635 -541
rect 661 -541 667 -535
rect 661 -561 924 -541
rect 430 -564 924 -561
rect -182 -565 924 -564
rect -472 -567 924 -565
rect -961 -568 -925 -567
rect -470 -569 -438 -567
rect -315 -568 -283 -567
rect -211 -568 -179 -567
rect -109 -568 -78 -567
rect 401 -568 432 -567
rect -984 -596 924 -593
rect -984 -622 -419 -596
rect -393 -599 924 -596
rect -393 -622 535 -599
rect -984 -625 535 -622
rect 561 -625 924 -599
rect -984 -633 924 -625
<< via2 >>
rect -915 -20 -812 9
rect -493 -281 -458 -279
rect -493 -307 -489 -281
rect -489 -307 -463 -281
rect -463 -307 -458 -281
rect -493 -309 -458 -307
<< metal3 >>
rect -920 9 -807 12
rect -920 -20 -915 9
rect -812 -20 -807 9
rect -920 -24 -914 -20
rect -813 -24 -807 -20
rect -920 -25 -807 -24
rect -961 -276 -512 -68
rect -961 -279 -455 -276
rect -961 -309 -493 -279
rect -458 -309 -455 -279
rect -961 -312 -455 -309
rect -961 -585 -512 -312
<< via3 >>
rect -914 -20 -813 8
rect -914 -24 -813 -20
<< mimcap >>
rect -929 -111 -544 -95
rect -929 -144 -913 -111
rect -808 -144 -544 -111
rect -929 -563 -544 -144
<< mimcapcontact >>
rect -913 -144 -808 -111
<< metal4 >>
rect -916 8 -804 10
rect -916 -24 -914 8
rect -813 -24 -804 8
rect -916 -111 -804 -24
rect -916 -144 -913 -111
rect -808 -144 -804 -111
rect -916 -149 -804 -144
<< labels >>
rlabel metal2 912 -21 924 17 0 VPWR
port 2 nsew
rlabel metal2 914 -633 924 -593 0 VGND
port 3 nsew
rlabel metal2 916 -567 924 -541 0 PBIAS
port 4 nsew
rlabel metal2 915 -199 924 -173 0 NBIAS
port 5 nsew
rlabel metal2 -984 -21 -975 17 0 VPWR
port 2 nsew
rlabel metal2 -984 -633 -972 -593 0 VGND
port 3 nsew
rlabel metal2 -984 -567 -972 -541 0 RESIST
port 6 nsew
<< end >>
