VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_wta4stage01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_wta4stage01 ;
  ORIGIN 11.210 0.430 ;
  SIZE 14.170 BY 6.050 ;
  OBS
      LAYER nwell ;
        RECT -11.010 5.610 -8.050 5.620 ;
        RECT -11.010 5.460 -10.600 5.610 ;
        RECT -11.010 5.450 -10.420 5.460 ;
        RECT -11.010 3.690 -10.600 5.450 ;
        RECT -11.120 2.540 -10.600 3.690 ;
        RECT -11.010 -0.420 -10.600 2.540 ;
      LAYER li1 ;
        RECT -11.150 -0.220 -10.970 0.670 ;
      LAYER met1 ;
        RECT -10.250 5.610 -10.090 5.620 ;
        RECT -9.440 5.610 -9.280 5.620 ;
        RECT -7.620 3.990 -7.400 5.370 ;
        RECT 1.310 5.160 1.540 5.620 ;
        RECT 2.570 5.160 2.800 5.620 ;
        RECT -11.120 2.540 -10.910 3.690 ;
        RECT -7.720 1.220 -7.450 2.120 ;
        RECT 1.310 -0.430 1.540 -0.180 ;
        RECT 2.570 -0.430 2.800 -0.180 ;
      LAYER met2 ;
        RECT -7.380 5.300 0.070 5.310 ;
        RECT -7.510 5.120 0.070 5.300 ;
        RECT -11.000 4.940 -10.610 5.120 ;
        RECT -7.510 5.100 0.240 5.120 ;
        RECT -0.140 4.910 0.240 5.100 ;
        RECT -11.120 4.180 -10.970 4.690 ;
        RECT -0.540 4.570 -0.500 4.660 ;
        RECT -0.650 4.370 0.560 4.570 ;
        RECT 1.700 4.260 2.960 4.420 ;
        RECT -11.120 4.020 -7.690 4.180 ;
        RECT -11.070 3.510 -10.900 3.690 ;
        RECT -0.550 3.510 0.660 3.710 ;
        RECT 1.700 3.330 2.960 3.490 ;
        RECT -11.000 3.080 -10.610 3.260 ;
        RECT -7.910 3.040 -7.680 3.050 ;
        RECT -7.910 3.010 -0.340 3.040 ;
        RECT -7.910 2.840 -0.280 3.010 ;
        RECT -7.910 2.740 -7.670 2.840 ;
        RECT -11.120 2.560 -7.670 2.740 ;
        RECT -0.470 2.640 0.240 2.840 ;
        RECT -11.120 2.540 -7.750 2.560 ;
        RECT -7.670 2.340 -0.320 2.360 ;
        RECT -7.670 2.140 0.240 2.340 ;
        RECT -11.000 1.930 -10.610 2.110 ;
        RECT -11.180 1.180 -10.980 1.680 ;
        RECT -0.560 1.520 0.440 1.680 ;
        RECT 1.700 1.490 2.960 1.650 ;
        RECT -11.180 0.980 -7.630 1.180 ;
        RECT -0.550 0.540 0.450 0.710 ;
        RECT 1.720 0.560 2.960 0.720 ;
        RECT -0.550 0.530 0.390 0.540 ;
        RECT -11.000 0.080 -10.610 0.260 ;
        RECT -0.320 0.080 0.230 0.090 ;
        RECT -7.900 -0.140 0.230 0.080 ;
        RECT -7.900 -0.150 -0.310 -0.140 ;
        RECT -7.900 -0.160 -7.130 -0.150 ;
        RECT -7.900 -0.200 -7.660 -0.160 ;
        RECT -11.140 -0.400 -7.660 -0.200 ;
        RECT -11.140 -0.410 -8.470 -0.400 ;
  END
END sky130_hilas_wta4stage01
END LIBRARY

