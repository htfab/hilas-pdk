magic
tech sky130A
timestamp 1628704331
<< checkpaint >>
rect -1026 1640 407 2027
rect -1026 1553 803 1640
rect 985 1553 3870 1640
rect -1026 1257 3870 1553
rect -1026 163 4083 1257
rect -630 -224 4083 163
rect 689 -343 4083 -224
rect 985 -584 4083 -343
rect 985 -610 3911 -584
rect 985 -630 3870 -610
<< error_s >>
rect 539 582 589 588
rect 611 582 661 588
rect 2579 582 2629 588
rect 2651 582 2701 588
rect 3039 586 3066 592
rect 539 540 589 546
rect 611 540 661 546
rect 2579 540 2629 546
rect 2651 540 2701 546
rect 3039 544 3066 550
rect 3039 519 3066 525
rect 3039 477 3066 483
rect 3039 436 3066 442
rect 3039 394 3066 400
rect 3039 369 3066 375
rect 3039 327 3066 333
rect 3039 286 3066 292
rect 3039 244 3066 250
rect 3039 219 3066 225
rect 3039 177 3066 183
rect 3039 136 3066 142
rect 3039 94 3066 100
rect 539 69 589 75
rect 611 69 661 75
rect 2579 69 2629 75
rect 2651 69 2701 75
rect 3039 69 3066 75
rect 539 27 589 33
rect 611 27 661 33
rect 2579 27 2629 33
rect 2651 27 2701 33
rect 3039 27 3066 33
<< nwell >>
rect 472 609 670 610
rect 2768 609 2915 610
rect 3153 592 3281 610
rect 472 542 479 560
rect 472 55 480 73
rect 3153 5 3281 24
<< locali >>
rect 1321 346 1341 353
rect 1321 329 1322 346
rect 1339 329 1341 346
rect 1321 274 1341 329
rect 1321 257 1323 274
rect 1340 257 1341 274
rect 1321 252 1341 257
rect 1896 346 1925 353
rect 1896 329 1901 346
rect 1918 329 1925 346
rect 1896 274 1925 329
rect 1896 257 1901 274
rect 1918 257 1925 274
rect 1896 252 1925 257
<< viali >>
rect 1322 329 1339 346
rect 1323 257 1340 274
rect 1901 329 1918 346
rect 1901 257 1918 274
<< metal1 >>
rect 496 605 524 610
rect 496 604 528 605
rect 549 604 568 610
rect 496 578 499 604
rect 525 578 528 604
rect 1197 601 1220 609
rect 1319 601 1342 609
rect 1548 594 1692 610
rect 1898 601 1921 610
rect 2020 602 2043 610
rect 2672 602 2691 610
rect 2716 605 2744 610
rect 2716 603 2748 605
rect 496 577 528 578
rect 2716 577 2719 603
rect 2745 577 2748 603
rect 3085 596 3119 610
rect 3151 595 3179 610
rect 2716 575 2748 577
rect 1322 328 1339 329
rect 1901 328 1918 329
rect 1320 297 1352 299
rect 1320 258 1323 297
rect 1349 271 1352 297
rect 1340 269 1352 271
rect 1890 291 1922 294
rect 1340 258 1344 269
rect 1890 265 1893 291
rect 1919 265 1922 291
rect 1890 262 1901 265
rect 1342 252 1344 258
rect 1918 262 1922 265
rect 2934 52 2967 54
rect 1890 39 1922 41
rect 1890 13 1893 39
rect 1919 13 1922 39
rect 2934 26 2937 52
rect 2964 26 2967 52
rect 2934 25 2967 26
rect 1890 11 1922 13
rect 2933 22 2975 25
rect 3035 24 3085 25
rect 3035 22 3119 24
rect 2933 11 3119 22
rect 2672 5 2691 10
rect 2716 5 2744 10
rect 2961 8 3051 11
rect 3085 5 3119 11
rect 3152 5 3179 26
<< via1 >>
rect 499 578 525 604
rect 2719 577 2745 603
rect 1323 274 1349 297
rect 1323 271 1340 274
rect 1340 271 1349 274
rect 1893 274 1919 291
rect 1893 265 1901 274
rect 1901 265 1918 274
rect 1918 265 1919 274
rect 1893 13 1919 39
rect 2937 26 2964 52
<< metal2 >>
rect 496 604 528 605
rect 496 578 499 604
rect 525 593 528 604
rect 2716 603 2748 605
rect 2716 593 2719 603
rect 525 578 2719 593
rect 496 577 2719 578
rect 2745 577 2748 603
rect 2828 583 2859 607
rect 496 575 2748 577
rect 472 542 479 560
rect 2939 520 2961 522
rect 1362 482 1446 502
rect 2934 486 2961 520
rect 1407 435 2421 457
rect 2760 436 2795 458
rect 1402 338 2303 360
rect 1320 297 1352 299
rect 1320 271 1323 297
rect 1349 294 1352 297
rect 1349 291 1922 294
rect 1349 271 1893 291
rect 1320 269 1893 271
rect 1890 265 1893 269
rect 1919 265 1922 291
rect 1890 262 1922 265
rect 1407 160 1973 182
rect 1357 130 1405 131
rect 1357 106 1446 130
rect 1951 127 1973 160
rect 2281 177 2303 338
rect 2399 315 2421 435
rect 2941 429 2961 430
rect 2941 396 2963 429
rect 2943 395 2963 396
rect 2836 316 2868 340
rect 3270 339 3281 362
rect 2396 311 2421 315
rect 2396 247 2422 311
rect 3270 257 3281 279
rect 2396 226 2809 247
rect 2788 212 2809 226
rect 2788 191 2990 212
rect 2281 155 2566 177
rect 2388 127 2990 132
rect 1951 111 2990 127
rect 1951 105 2427 111
rect 472 55 480 73
rect 2934 52 2967 54
rect 1890 40 1922 41
rect 2934 40 2937 52
rect 1890 39 2937 40
rect 1890 13 1893 39
rect 1919 26 2937 39
rect 2964 26 2967 52
rect 1919 24 2967 26
rect 1919 23 1959 24
rect 1919 13 1922 23
rect 1890 11 1922 13
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1628704305
transform 1 0 3126 0 1 46
box 0 0 327 581
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1628704305
transform 1 0 2634 0 -1 170
box 133 -454 320 165
use sky130_hilas_FGBias2x1cell  sky130_hilas_FGBias2x1cell_0
timestamp 1628704315
transform 1 0 2011 0 1 387
box 0 0 1625 1010
use sky130_hilas_FGBiasWeakGate2x1cell  sky130_hilas_FGBiasWeakGate2x1cell_0
timestamp 1628704305
transform -1 0 1229 0 1 387
box 0 0 1625 1010
<< labels >>
rlabel metal2 1362 482 1398 501 0 VIN11
port 2 nsew analog default
rlabel metal2 1357 106 1393 131 0 VIN12
port 1 nsew analog default
rlabel metal1 3085 604 3119 610 0 VGND
port 7 nsew analog default
rlabel metal1 3151 604 3179 610 0 VPWR
port 6 nsew analog default
rlabel metal1 3152 5 3179 11 0 VPWR
port 6 nsew power default
rlabel metal1 3085 5 3119 11 0 VGND
port 7 nsew ground default
rlabel metal2 2836 316 2868 340 0 VIN21
port 3 nsew analog default
rlabel metal2 2828 583 2859 607 1 VIN22
port 4 n analog default
rlabel metal1 2716 602 2744 610 0 VINJ
port 8 nsew power default
rlabel metal1 2716 5 2744 10 0 VINJ
port 8 nsew power default
rlabel metal2 3270 339 3281 362 0 OUTPUT1
port 9 nsew analog default
rlabel metal2 3270 257 3281 279 0 OUTPUT2
port 10 nsew analog default
rlabel metal2 472 542 479 560 0 DRAIN1
port 11 nsew
rlabel metal2 472 55 480 73 0 DRAIN2
port 12 nsew
rlabel metal1 496 603 524 610 0 VINJ
port 8 nsew
rlabel metal1 549 604 568 610 0 COLSEL2
port 13 nsew
rlabel metal1 1197 601 1220 609 0 GATE2
port 14 nsew
rlabel metal1 1319 601 1342 609 0 VGND
port 7 nsew
rlabel metal1 2020 602 2043 610 0 GATE1
port 15 nsew
rlabel metal1 1898 602 1921 610 0 VGND
port 7 nsew
rlabel metal1 2672 602 2691 610 0 COLSEL1
port 16 nsew
rlabel metal1 2672 5 2691 10 0 COLSEL1
port 16 nsew
rlabel metal1 1590 598 1650 610 0 VTUN
port 17 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
