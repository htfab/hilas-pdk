magic
tech sky130A
timestamp 1628698463
<< checkpaint >>
rect -517 676 990 816
rect -517 -473 1002 676
rect -502 -611 1002 -473
rect -502 -721 997 -611
<< nwell >>
rect 68 52 472 189
<< mvnmos >>
rect 130 -56 341 5
<< mvpmos >>
rect 130 86 340 148
<< mvndiff >>
rect 101 1 130 5
rect 101 -16 107 1
rect 124 -16 130 1
rect 101 -33 130 -16
rect 101 -50 107 -33
rect 124 -50 130 -33
rect 101 -56 130 -50
rect 341 1 370 5
rect 341 -16 347 1
rect 364 -16 370 1
rect 341 -33 370 -16
rect 341 -50 347 -33
rect 364 -50 370 -33
rect 341 -56 370 -50
<< mvpdiff >>
rect 101 143 130 148
rect 101 126 107 143
rect 124 126 130 143
rect 101 109 130 126
rect 101 92 107 109
rect 124 92 130 109
rect 101 86 130 92
rect 340 143 370 148
rect 340 126 346 143
rect 363 126 370 143
rect 340 109 370 126
rect 340 92 346 109
rect 363 92 370 109
rect 340 86 370 92
<< mvndiffc >>
rect 107 -16 124 1
rect 107 -50 124 -33
rect 347 -16 364 1
rect 347 -50 364 -33
<< mvpdiffc >>
rect 107 126 124 143
rect 107 92 124 109
rect 346 126 363 143
rect 346 92 363 109
<< psubdiff >>
rect 389 -2 458 10
rect 389 -19 399 -2
rect 416 -19 433 -2
rect 450 -19 458 -2
rect 389 -36 458 -19
rect 389 -53 399 -36
rect 416 -53 433 -36
rect 450 -53 458 -36
rect 389 -70 458 -53
rect 382 -87 399 -70
rect 416 -87 433 -70
rect 450 -87 458 -70
rect 389 -99 458 -87
<< mvnsubdiff >>
rect 397 144 439 156
rect 397 127 409 144
rect 426 127 439 144
rect 397 110 439 127
rect 397 93 409 110
rect 426 93 439 110
rect 397 86 439 93
<< psubdiffcont >>
rect 399 -19 416 -2
rect 433 -19 450 -2
rect 399 -53 416 -36
rect 433 -53 450 -36
rect 399 -87 416 -70
rect 433 -87 450 -70
<< mvnsubdiffcont >>
rect 409 127 426 144
rect 409 93 426 110
<< poly >>
rect 130 148 341 163
rect 130 85 340 86
rect 130 68 341 85
rect 130 67 231 68
rect 163 40 164 67
rect 197 40 198 67
rect 304 20 305 46
rect 338 20 339 46
rect 271 19 341 20
rect 130 5 341 19
rect 130 -69 341 -56
<< locali >>
rect 99 183 429 189
rect 99 182 158 183
rect 166 182 265 183
rect 275 182 429 183
rect 99 179 429 182
rect 99 162 377 179
rect 394 162 412 179
rect 99 144 429 162
rect 99 143 409 144
rect 99 126 107 143
rect 124 126 346 143
rect 363 127 409 143
rect 426 127 429 144
rect 363 126 429 127
rect 99 110 428 126
rect 99 109 409 110
rect 99 92 107 109
rect 124 92 346 109
rect 363 93 409 109
rect 426 93 428 110
rect 363 92 428 93
rect 99 85 428 92
rect 99 1 231 67
rect 271 24 428 85
rect 367 4 450 6
rect 361 1 450 4
rect 99 -16 107 1
rect 124 -16 347 1
rect 364 -2 450 1
rect 364 -16 399 -2
rect 99 -19 399 -16
rect 416 -19 433 -2
rect 99 -33 450 -19
rect 99 -50 107 -33
rect 124 -50 347 -33
rect 364 -36 450 -33
rect 364 -50 399 -36
rect 99 -53 399 -50
rect 416 -53 433 -36
rect 99 -70 450 -53
rect 99 -87 382 -70
rect 99 -88 450 -87
rect 375 -95 450 -88
<< viali >>
rect 377 162 394 179
rect 412 162 429 179
rect 382 -87 399 -70
rect 416 -87 433 -70
<< metal1 >>
rect 68 179 473 189
rect 68 162 377 179
rect 394 162 412 179
rect 429 162 473 179
rect 68 142 473 162
rect 99 141 473 142
rect 68 -64 373 -50
rect 68 -70 473 -64
rect 68 -87 382 -70
rect 399 -87 416 -70
rect 433 -87 473 -70
rect 68 -113 473 -87
use sky130_hilas_poly2li  sky130_hilas_poly2li_4
timestamp 1628285143
transform 0 1 285 -1 0 37
box -9 -14 18 19
use sky130_hilas_poly2li  sky130_hilas_poly2li_3
timestamp 1628285143
transform 0 1 353 -1 0 37
box -9 -14 18 19
use sky130_hilas_poly2li  sky130_hilas_poly2li_0
timestamp 1628285143
transform 0 1 319 -1 0 37
box -9 -14 18 19
use sky130_hilas_poly2li  sky130_hilas_poly2li_1
timestamp 1628285143
transform 0 1 144 -1 0 58
box -9 -14 18 19
use sky130_hilas_poly2li  sky130_hilas_poly2li_2
timestamp 1628285143
transform 0 1 178 -1 0 58
box -9 -14 18 19
use sky130_hilas_poly2li  sky130_hilas_poly2li_5
timestamp 1628285143
transform 0 1 212 -1 0 58
box -9 -14 18 19
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1628285143
transform 1 0 174 0 1 -83
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1628285143
transform 1 0 138 0 1 -83
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_3
timestamp 1628285143
transform 1 0 210 0 1 -83
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_2
timestamp 1628285143
transform 1 0 282 0 1 -83
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_5
timestamp 1628285143
transform 1 0 246 0 1 -83
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_7
timestamp 1628285143
transform 1 0 354 0 1 -83
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_4
timestamp 1628285143
transform 1 0 318 0 1 -83
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_10
timestamp 1628285143
transform 1 0 159 0 1 165
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_9
timestamp 1628285143
transform 1 0 123 0 1 165
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_12
timestamp 1628285143
transform 1 0 231 0 1 165
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_11
timestamp 1628285143
transform 1 0 195 0 1 165
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_13
timestamp 1628285143
transform 1 0 267 0 1 165
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_15
timestamp 1628285143
transform 1 0 347 0 1 165
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_14
timestamp 1628285143
transform 1 0 303 0 1 165
box -10 -8 13 21
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
