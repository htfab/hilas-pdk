magic
tech sky130A
magscale 1 2
timestamp 1628276330
<< error_s >>
rect 70 1108 170 1120
rect 716 1110 816 1122
rect 1030 1108 1086 1122
rect 1314 1110 1370 1122
rect 70 1024 170 1036
rect 716 1026 816 1038
rect 1030 1024 1086 1038
rect 1314 1026 1370 1038
rect 212 976 312 988
rect 572 966 674 978
rect 932 966 988 978
rect 1412 966 1468 978
rect 212 892 312 904
rect 572 882 674 894
rect 932 882 988 894
rect 1412 882 1468 894
rect 70 758 170 770
rect 716 760 816 772
rect 1030 758 1086 772
rect 1314 760 1370 772
rect 70 674 170 686
rect 716 676 816 688
rect 1030 674 1086 688
rect 1314 676 1370 688
rect 212 626 312 638
rect 572 616 674 628
rect 932 616 988 628
rect 1412 616 1468 628
rect 212 542 312 554
rect 572 532 674 544
rect 932 532 988 544
rect 1412 532 1468 544
rect 70 408 170 420
rect 716 410 816 422
rect 1030 408 1086 422
rect 1314 410 1370 422
rect 70 324 170 336
rect 716 326 816 338
rect 1030 324 1086 338
rect 1314 326 1370 338
rect 212 276 312 288
rect 572 266 674 278
rect 932 266 988 278
rect 1412 266 1468 278
rect 212 192 312 204
rect 572 182 674 194
rect 932 182 988 194
rect 1412 182 1468 194
rect 70 58 170 70
rect 716 60 816 72
rect 1030 58 1086 72
rect 1314 60 1370 72
rect 70 -26 170 -14
rect 716 -24 816 -12
rect 1030 -26 1086 -12
rect 1314 -24 1370 -12
rect 212 -74 312 -62
rect 572 -84 674 -72
rect 932 -84 988 -72
rect 1412 -84 1468 -72
rect 212 -158 312 -146
rect 572 -168 674 -156
rect 932 -168 988 -156
rect 1412 -168 1468 -156
<< metal2 >>
rect 1676 874 1730 938
rect 1676 524 1784 588
rect 1674 174 1800 238
rect 1674 -114 1708 -112
rect 1646 -176 1871 -114
use sky130_hilas_StepUpDigital  StepUpDigital_0
timestamp 1628276300
transform 1 0 -98 0 1 226
box -148 -88 1778 262
use sky130_hilas_StepUpDigital  StepUpDigital_3
timestamp 1628276300
transform 1 0 -98 0 1 -124
box -148 -88 1778 262
use sky130_hilas_StepUpDigital  StepUpDigital_1
timestamp 1628276300
transform 1 0 -98 0 1 576
box -148 -88 1778 262
use sky130_hilas_StepUpDigital  StepUpDigital_2
timestamp 1628276300
transform 1 0 -98 0 1 926
box -148 -88 1778 262
<< labels >>
rlabel space 1492 1034 1540 1044 0 VPWR
port 5 nsew
rlabel metal1 1492 -204 1540 -194 0 VPWR
port 5 nsew
rlabel space 8 1034 66 1044 0 VINJ
port 6 nsew
rlabel metal1 8 -204 66 -194 0 VINJ
port 6 nsew
rlabel space 890 1030 952 1044 0 VGND
port 11 nsew
rlabel metal1 890 -204 952 -192 0 VGND
port 11 nsew
rlabel metal2 1808 -176 1870 -114 1 INPUT4
port 12 n
rlabel metal2 1784 174 1800 238 1 INPUT3
port 13 n
rlabel metal2 1762 524 1784 588 1 INPUT2
port 14 n
rlabel metal2 1712 874 1728 938 1 INPUT1
port 15 n
rlabel space -140 1060 -124 1100 1 OUTPUT1
port 16 n
rlabel space -140 710 -124 750 1 OUTPUT2
port 8 n
rlabel space -140 360 -110 400 1 OUTPUT3
port 9 n
rlabel space -140 10 -126 50 1 OUTPUT4
port 17 n
<< end >>
