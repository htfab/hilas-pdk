magic
tech sky130A
timestamp 1632251355
<< nwell >>
rect 0 1 173 185
<< mvnsubdiff >>
rect 54 81 113 110
rect 54 54 69 81
rect 97 54 113 81
rect 54 36 113 54
<< mvnsubdiffcont >>
rect 69 54 97 81
<< locali >>
rect 42 81 97 89
rect 42 46 97 54
<< viali >>
rect 42 54 69 81
<< metal1 >>
rect 36 81 75 186
rect 36 54 42 81
rect 69 54 75 81
rect 36 0 75 54
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
