* Copyright 2020 The Hilas PDK Authors
* 
* This file is part of HILAS.
* 
* HILAS is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published by
* the Free Software Foundation, version 3 of the License.
* 
* HILAS is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
* 
* You should have received a copy of the GNU Lesser General Public License
* along with HILAS.  If not, see <https://www.gnu.org/licenses/>.
* 
* Licensed under the Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
* https://www.gnu.org/licenses/lgpl-3.0.en.html
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
* SPDX-License-Identifier: LGPL-3.0
* 
* 

* NGSPICE file created from sky130_hilas_swc4x1BiasCell.ext - technology: sky130A

.subckt sky130_hilas_TunCap01 SUB a_n2872_n666# w_n2902_n800#
X0 a_n2872_n666# w_n2902_n800# w_n2902_n800# sky130_fd_pr__cap_var w=590000u l=500000u
.ends

.subckt sky130_hilas_horizPcell01 a_n502_286# a_n508_162# SUB w_n578_94# a_n578_238#
+ m1_n258_94# a_n300_94# a_n344_286#
X0 w_n578_94# a_n300_94# a_n344_162# w_n578_94# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
X1 a_n344_286# a_n578_238# a_n502_286# w_n578_94# sky130_fd_pr__pfet_g5v0d10v5 w=300000u l=500000u
X2 a_n344_162# a_n578_238# a_n508_162# w_n578_94# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
.ends

.subckt sky130_hilas_FGVaractorCapacitor SUB m1_n1784_n790# a_n1882_n672# w_n1914_n790#
X0 a_n1882_n672# w_n1914_n790# w_n1914_n790# sky130_fd_pr__cap_var w=1.11e+06u l=640000u
.ends

.subckt sky130_hilas_swc4x1BiasCell BIAS1 BIAS2 BIAS3 BIAS4 VTUN GATE VINJ VPWR GATESELECT
+ DRAIN1 DRAIN2 DRAIN3 DRAIN4
Xsky130_hilas_TunCap01_0 SUB a_640_n334# VTUN sky130_hilas_TunCap01
Xsky130_hilas_TunCap01_1 SUB a_640_n618# VTUN sky130_hilas_TunCap01
Xsky130_hilas_TunCap01_2 SUB a_n214_10# VTUN sky130_hilas_TunCap01
Xsky130_hilas_TunCap01_3 SUB a_638_270# VTUN sky130_hilas_TunCap01
Xsky130_hilas_horizPcell01_0 BIAS2 DRAIN2 SUB VINJ a_n214_10# GATESELECT GATESELECT
+ VPWR sky130_hilas_horizPcell01
Xsky130_hilas_horizPcell01_1 BIAS4 DRAIN4 SUB VINJ a_640_n618# GATESELECT GATESELECT
+ VPWR sky130_hilas_horizPcell01
Xsky130_hilas_horizPcell01_2 BIAS3 DRAIN3 SUB VINJ a_640_n334# GATESELECT GATESELECT
+ VPWR sky130_hilas_horizPcell01
Xsky130_hilas_horizPcell01_3 BIAS1 DRAIN1 SUB VINJ a_638_270# GATESELECT GATESELECT
+ VPWR sky130_hilas_horizPcell01
Xsky130_hilas_FGVaractorCapacitor_0 SUB GATE a_640_n618# GATE sky130_hilas_FGVaractorCapacitor
Xsky130_hilas_FGVaractorCapacitor_2 SUB GATE a_n214_10# GATE sky130_hilas_FGVaractorCapacitor
Xsky130_hilas_FGVaractorCapacitor_1 SUB GATE a_640_n334# GATE sky130_hilas_FGVaractorCapacitor
Xsky130_hilas_FGVaractorCapacitor_3 SUB GATE a_638_270# GATE sky130_hilas_FGVaractorCapacitor
.ends

