magic
tech sky130A
timestamp 1628698459
<< metal2 >>
rect 1414 480 2211 498
rect 1414 437 2211 455
rect 1417 337 2211 355
rect 1417 294 2211 312
rect 1416 232 1443 260
rect 2180 234 2211 262
rect 1417 179 2211 196
rect 1417 137 2211 154
rect 1417 39 2211 56
rect 1417 -5 2211 12
<< metal3 >>
rect 1982 222 2180 283
rect 1982 221 2178 222
rect 2179 221 2180 222
rect 1982 208 2180 221
<< metal4 >>
rect 1530 272 1631 273
rect 1459 222 1794 272
rect 1459 221 1566 222
rect 1730 110 1793 222
rect 1730 80 1945 110
rect 1763 79 1945 80
use sky130_hilas_m22m4  sky130_hilas_m22m4_0
timestamp 1607701799
transform 1 0 1452 0 1 242
box -36 -36 43 39
use sky130_hilas_CapModule03  sky130_hilas_CapModule03_0
timestamp 1607813757
transform 1 0 1952 0 1 199
box -392 -247 31 336
use sky130_hilas_m22m4  sky130_hilas_m22m4_1
timestamp 1607701799
transform 1 0 2164 0 1 244
box -36 -36 43 39
<< labels >>
rlabel metal2 1416 232 1423 260 0 CAPTERM01
port 2 nsew analog default
rlabel metal2 2196 234 2211 262 0 CAPTERM02
port 1 nsew analog default
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
