magic
tech sky130A
timestamp 1628617061
<< checkpaint >>
rect -611 1175 821 1253
rect -691 897 821 1175
rect -691 -414 836 897
rect -691 -608 810 -414
rect -691 -650 730 -608
<< error_s >>
rect 1 522 40 525
rect 1 480 40 483
rect 0 426 39 429
rect 0 384 39 387
rect 0 330 39 333
rect 0 288 39 291
rect 0 234 39 237
rect 0 192 39 195
rect 0 138 39 141
rect 0 96 39 99
rect 1 42 40 45
rect 1 0 40 3
use sky130_hilas_pFETdevice01a  sky130_hilas_pFETdevice01a_0
timestamp 1628617045
transform 1 0 19 0 1 22
box 0 0 161 85
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_0
timestamp 1628617059
transform 1 0 18 0 1 118
box 0 0 161 121
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_3
timestamp 1628617059
transform 1 0 18 0 1 310
box 0 0 161 121
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_6
timestamp 1628617059
transform 1 0 18 0 1 406
box 0 0 161 121
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_0
timestamp 1628616950
transform 1 0 19 0 1 502
box 0 0 172 121
use sky130_hilas_pFETdevice01b  sky130_hilas_pFETdevice01b_1
timestamp 1628617034
transform 1 0 18 0 1 214
box 0 0 188 133
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
