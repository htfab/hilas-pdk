magic
tech sky130A
timestamp 1628704290
<< checkpaint >>
rect -1025 1640 408 2027
rect -1025 1598 803 1640
rect -1025 1553 983 1598
rect 986 1553 3871 1640
rect -1025 1242 3871 1553
rect -1025 1020 4051 1242
rect -1025 163 4056 1020
rect -630 -224 4056 163
rect 105 -273 4056 -224
rect 105 -285 4055 -273
rect 106 -345 4055 -285
rect 106 -392 4047 -345
rect 108 -570 4047 -392
rect 108 -583 3912 -570
rect 986 -610 3912 -583
rect 986 -630 3871 -610
<< error_s >>
rect 539 582 589 588
rect 611 582 661 588
rect 2580 582 2630 588
rect 2652 582 2702 588
rect 3040 586 3067 592
rect 539 540 589 546
rect 611 540 661 546
rect 2580 540 2630 546
rect 2652 540 2702 546
rect 3040 544 3067 550
rect 3040 519 3067 525
rect 724 438 727 488
rect 766 438 769 488
rect 860 438 862 488
rect 902 438 904 488
rect 3040 477 3067 483
rect 3040 436 3067 442
rect 724 359 727 409
rect 766 359 769 409
rect 860 359 862 409
rect 902 359 904 409
rect 3040 394 3067 400
rect 3040 369 3067 375
rect 3040 327 3067 333
rect 3040 286 3067 292
rect 724 206 727 256
rect 766 206 769 256
rect 860 206 862 256
rect 902 206 904 256
rect 3040 244 3067 250
rect 3040 219 3067 225
rect 3040 177 3067 183
rect 724 127 727 177
rect 766 127 769 177
rect 860 127 862 177
rect 902 127 904 177
rect 3040 136 3067 142
rect 3040 94 3067 100
rect 539 69 589 75
rect 611 69 661 75
rect 2580 69 2630 75
rect 2652 69 2702 75
rect 3040 69 3067 75
rect 539 27 589 33
rect 611 27 661 33
rect 2580 27 2630 33
rect 2652 27 2702 33
rect 3040 27 3067 33
<< nwell >>
rect 472 609 803 610
rect 2769 609 2903 610
rect 492 578 524 608
rect 2719 578 2751 608
rect 3154 592 3282 610
rect 3154 5 3282 24
<< metal1 >>
rect 508 608 524 610
rect 492 606 524 608
rect 492 580 495 606
rect 521 580 524 606
rect 549 604 568 610
rect 736 599 757 610
rect 783 602 802 610
rect 824 604 845 610
rect 932 603 950 610
rect 1548 595 1590 610
rect 1651 595 1693 610
rect 2021 602 2044 610
rect 2673 602 2692 610
rect 2717 608 2745 610
rect 2717 606 2751 608
rect 2717 602 2722 606
rect 1548 581 1693 595
rect 492 578 524 580
rect 2719 580 2722 602
rect 2748 580 2751 606
rect 3086 596 3120 610
rect 3152 595 3180 610
rect 2719 578 2751 580
rect 2933 53 2965 55
rect 1314 38 1346 40
rect 737 6 760 18
rect 1314 12 1317 38
rect 1343 12 1346 38
rect 1314 10 1346 12
rect 1894 38 1926 40
rect 1894 12 1897 38
rect 1923 12 1926 38
rect 2933 27 2936 53
rect 2962 27 2965 53
rect 2933 25 2965 27
rect 2933 22 2976 25
rect 3036 24 3087 25
rect 3036 22 3120 24
rect 2933 19 3120 22
rect 2948 14 3120 19
rect 1894 10 1926 12
rect 2951 11 3120 14
rect 2673 5 2692 10
rect 2717 5 2745 10
rect 2954 9 3120 11
rect 2961 8 3057 9
rect 3086 5 3120 9
rect 3153 5 3180 26
<< via1 >>
rect 495 580 521 606
rect 2722 580 2748 606
rect 1317 12 1343 38
rect 1897 12 1923 38
rect 2936 27 2962 53
<< metal2 >>
rect 492 606 524 608
rect 492 580 495 606
rect 521 596 524 606
rect 2719 606 2751 608
rect 2719 596 2722 606
rect 521 580 2722 596
rect 2748 580 2751 606
rect 2829 583 2860 607
rect 492 578 2751 580
rect 472 542 480 560
rect 2940 520 2962 522
rect 2935 486 2962 520
rect 2761 436 2796 458
rect 2942 429 2962 430
rect 1623 387 2422 407
rect 2942 396 2964 429
rect 2944 395 2964 396
rect 2282 319 2304 320
rect 1624 294 2307 319
rect 2400 315 2422 387
rect 2837 316 2869 340
rect 3271 339 3282 362
rect 1624 202 1975 221
rect 1952 142 1975 202
rect 2278 177 2307 294
rect 2397 311 2422 315
rect 2397 247 2423 311
rect 3271 257 3282 279
rect 2397 226 2810 247
rect 2789 212 2810 226
rect 2789 191 2990 212
rect 2278 155 2567 177
rect 2278 154 2307 155
rect 1952 127 1974 142
rect 2389 127 2989 132
rect 1952 112 2989 127
rect 1952 111 2976 112
rect 1952 105 2428 111
rect 472 55 480 73
rect 2933 53 2965 55
rect 2933 40 2936 53
rect 1314 38 2936 40
rect 1314 12 1317 38
rect 1343 25 1897 38
rect 1343 12 1346 25
rect 1314 10 1346 12
rect 1894 12 1897 25
rect 1923 27 2936 38
rect 2962 27 2965 53
rect 1923 25 2965 27
rect 1923 12 1926 25
rect 1894 10 1926 12
use sky130_hilas_FGBias2x1cell  sky130_hilas_FGBias2x1cell_0
timestamp 1628704264
transform 1 0 2012 0 1 387
box -396 -387 1229 623
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1628704264
transform 1 0 2635 0 -1 170
box 133 -440 320 165
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1628704272
transform 1 0 3127 0 1 46
box 0 0 327 579
use sky130_hilas_FGtrans2x1cell  sky130_hilas_FGtrans2x1cell_0
timestamp 1628704264
transform -1 0 1229 0 1 387
box 0 0 1624 1010
<< labels >>
rlabel metal1 3086 604 3120 610 0 VGND
port 11 nsew
rlabel metal1 3152 604 3180 610 0 VPWR
port 10 nsew
rlabel metal1 3153 5 3180 11 0 VPWR
port 10 nsew
rlabel metal1 3086 5 3120 11 0 VGND
port 11 nsew
rlabel metal2 2837 316 2869 340 0 VIN21
port 9 nsew
rlabel metal2 2829 583 2860 607 1 VIN22
port 8 n
rlabel metal1 737 6 760 18 0 VIN12
port 18 nsew
rlabel metal1 736 599 757 610 0 VIN11
port 5 nsew
rlabel metal1 1651 603 1693 610 0 VTUN
port 1 nsew
rlabel metal1 1548 603 1590 610 0 VTUN
rlabel metal1 824 604 845 610 0 PROG
port 3 nsew
rlabel metal1 508 604 524 610 0 VINJ
port 6 nsew
rlabel metal1 2717 602 2745 610 0 VINJ
port 6 nsew
rlabel metal2 3271 339 3282 362 0 OUTPUT1
port 13 nsew
rlabel metal2 3271 257 3282 279 0 OUTPUT2
port 12 nsew
rlabel metal1 549 604 568 610 0 GATESEL1
port 14 nsew
rlabel metal1 2673 5 2692 10 0 GATESEL2
port 15 nsew
rlabel metal1 2717 5 2745 10 0 VINJ
port 6 nsew
rlabel metal1 2673 602 2692 610 0 GATESEL2
port 15 nsew
rlabel metal2 472 542 480 560 0 DRAIN1
port 16 nsew
rlabel metal2 472 55 480 73 0 DRAIN2
port 17 nsew
rlabel metal1 2021 602 2044 610 0 GATE1
port 4 nsew
rlabel metal1 783 602 802 610 0 GATE2
port 19 nsew
rlabel metal1 932 603 950 610 0 RUN
port 20 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
