magic
tech sky130A
timestamp 1628694524
<< checkpaint >>
rect -692 1334 1426 1377
rect -692 1284 1460 1334
rect -692 -626 1479 1284
rect -395 -670 1479 -626
<< error_s >>
rect 44 620 94 626
rect 367 621 417 627
rect 524 620 552 627
rect 666 621 694 627
rect 44 578 94 584
rect 367 579 417 585
rect 524 578 552 585
rect 666 579 694 585
rect 115 554 165 560
rect 295 549 346 555
rect 475 549 503 555
rect 715 549 743 555
rect 115 512 165 518
rect 295 507 346 513
rect 475 507 503 513
rect 715 507 743 513
rect 44 445 94 451
rect 367 446 417 452
rect 524 445 552 452
rect 666 446 694 452
rect 44 403 94 409
rect 367 404 417 410
rect 524 403 552 410
rect 666 404 694 410
rect 115 379 165 385
rect 295 374 346 380
rect 475 374 503 380
rect 715 374 743 380
rect 115 337 165 343
rect 295 332 346 338
rect 475 332 503 338
rect 715 332 743 338
rect 44 270 94 276
rect 367 271 417 277
rect 524 270 552 277
rect 666 271 694 277
rect 44 228 94 234
rect 367 229 417 235
rect 524 228 552 235
rect 666 229 694 235
rect 115 204 165 210
rect 295 199 346 205
rect 475 199 503 205
rect 715 199 743 205
rect 115 162 165 168
rect 295 157 346 163
rect 475 157 503 163
rect 715 157 743 163
rect 44 95 94 101
rect 367 96 417 102
rect 524 95 552 102
rect 666 96 694 102
rect 44 53 94 59
rect 367 54 417 60
rect 524 53 552 60
rect 666 54 694 60
rect 115 29 165 35
rect 295 24 346 30
rect 475 24 503 30
rect 715 24 743 30
rect 115 -13 165 -7
rect 295 -18 346 -12
rect 475 -18 503 -12
rect 715 -18 743 -12
<< nwell >>
rect -21 536 -10 556
<< metal1 >>
rect 13 651 42 660
rect 444 654 475 660
rect 745 655 769 660
rect 13 -40 42 -28
rect 444 -40 475 -34
rect 745 -40 769 -35
<< metal2 >>
rect -21 596 -5 616
rect 839 503 849 535
rect -21 421 -4 441
rect 839 328 849 360
rect -21 246 -2 266
rect 839 153 849 185
rect -21 71 -5 91
rect 839 -22 849 10
use sky130_hilas_StepUpDigital  StepUpDigital_2
timestamp 1628617025
transform 1 0 -40 0 1 529
box 0 0 836 218
use sky130_hilas_StepUpDigital  StepUpDigital_1
timestamp 1628617025
transform 1 0 -40 0 1 354
box 0 0 836 218
use sky130_hilas_StepUpDigital  StepUpDigital_3
timestamp 1628617025
transform 1 0 -40 0 1 4
box 0 0 836 218
use sky130_hilas_StepUpDigital  StepUpDigital_0
timestamp 1628617025
transform 1 0 -40 0 1 179
box 0 0 836 218
<< labels >>
rlabel metal1 13 -36 42 -31 0 VINJ
port 6 nsew
rlabel metal2 -21 71 -10 91 0 OUTPUT4
port 10 nsew
rlabel metal2 839 503 849 535 0 INPUT1
port 12 nsew
rlabel metal2 839 328 849 360 0 INPUT2
port 13 nsew
rlabel metal2 839 153 849 185 0 INPUT3
port 14 nsew
rlabel metal2 839 -22 849 10 0 INPUT4
port 15 nsew
rlabel metal2 -21 246 -13 266 0 OUTPUT3
port 9 nsew
rlabel metal2 -21 421 -14 441 0 OUTPUT2
port 8 nsew
rlabel metal2 -21 596 -14 616 0 OUTPUT1
port 7 nsew
rlabel metal1 444 -40 475 -34 0 VGND
port 11 nsew
rlabel metal1 444 654 475 660 0 VGND
port 11 nsew
rlabel metal1 13 651 42 660 0 VINJ
port 6 nsew
rlabel metal1 745 655 769 660 0 VPWR
port 5 nsew
rlabel metal1 745 -40 769 -35 0 VPWR
port 5 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
