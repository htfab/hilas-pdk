magic
tech sky130A
timestamp 1626543161
<< nwell >>
rect 742 -38 1947 556
<< mvndiff >>
rect -558 543 599 548
rect -558 526 -552 543
rect 593 526 599 543
rect -558 517 599 526
rect -558 486 -527 517
rect -558 479 599 486
rect -558 462 -552 479
rect 593 462 599 479
rect -558 455 599 462
rect -558 424 -527 455
rect -558 417 599 424
rect -558 400 -552 417
rect 592 400 599 417
rect -558 394 599 400
rect -558 364 -527 394
rect -558 357 599 364
rect -558 340 -552 357
rect 593 340 599 357
rect -558 334 599 340
rect -558 304 -527 334
rect -558 298 599 304
rect -558 281 -552 298
rect 593 281 599 298
rect -558 275 599 281
rect -558 245 -527 275
rect -558 239 599 245
rect -558 222 -552 239
rect 593 222 599 239
rect -558 216 599 222
rect -558 186 -527 216
rect -558 180 599 186
rect -558 163 -552 180
rect 592 163 599 180
rect -558 156 599 163
rect -558 125 -527 156
rect 568 155 599 156
rect -558 119 599 125
rect -558 102 -552 119
rect 593 102 599 119
rect -558 95 599 102
rect -558 64 -527 95
rect -558 57 599 64
rect -558 40 -551 57
rect 593 40 599 57
rect -558 34 599 40
rect -558 4 -527 34
rect -559 -4 599 4
rect -559 -21 -552 -4
rect 592 -21 599 -4
rect -559 -26 599 -21
<< mvpdiff >>
rect 832 463 1850 472
rect 832 446 839 463
rect 1819 446 1850 463
rect 832 441 1850 446
rect 1819 404 1850 441
rect 836 396 1850 404
rect 836 379 844 396
rect 1813 379 1850 396
rect 836 372 1850 379
rect 1819 330 1850 372
rect 841 323 1850 330
rect 841 306 849 323
rect 1824 306 1850 323
rect 841 298 1850 306
rect 1819 261 1850 298
rect 841 255 1850 261
rect 841 238 848 255
rect 1816 238 1850 255
rect 841 229 1850 238
rect 1819 196 1850 229
rect 837 188 1850 196
rect 837 171 844 188
rect 1818 171 1850 188
rect 837 163 1850 171
rect 1819 132 1850 163
rect 837 124 1850 132
rect 837 107 843 124
rect 1816 107 1850 124
rect 837 99 1850 107
rect 1819 69 1850 99
rect 837 62 1850 69
rect 837 45 845 62
rect 1816 45 1850 62
rect 837 38 1850 45
<< mvndiffc >>
rect -552 526 593 543
rect -552 462 593 479
rect -552 400 592 417
rect -552 340 593 357
rect -552 281 593 298
rect -552 222 593 239
rect -552 163 592 180
rect -552 102 593 119
rect -551 40 593 57
rect -552 -21 592 -4
<< mvpdiffc >>
rect 839 446 1819 463
rect 844 379 1813 396
rect 849 306 1824 323
rect 848 238 1816 255
rect 844 171 1818 188
rect 843 107 1816 124
rect 845 45 1816 62
<< psubdiff >>
rect -698 648 -664 649
rect -698 646 -646 648
rect 646 646 2054 648
rect -698 640 2054 646
rect -698 623 -621 640
rect 1966 623 2054 640
rect -698 606 2054 623
rect -698 589 -621 606
rect 1966 589 2054 606
rect -698 583 2054 589
rect -698 -55 -690 583
rect -673 570 -631 583
rect -673 -39 -656 570
rect -639 -39 -631 570
rect 646 579 2056 583
rect 646 570 709 579
rect -673 -55 -631 -39
rect -698 -56 -631 -55
rect 646 -44 651 570
rect 668 568 709 570
rect 668 -44 685 568
rect 646 -45 685 -44
rect 702 -45 709 568
rect 1988 577 2056 579
rect 646 -52 709 -45
rect 1988 -45 1993 577
rect 2010 573 2056 577
rect 2010 -45 2031 573
rect 1988 -46 2031 -45
rect 2048 -46 2056 573
rect 1988 -52 2056 -46
rect 646 -56 2056 -52
rect -698 -62 2056 -56
rect -698 -79 -624 -62
rect 1977 -79 2056 -62
rect -698 -96 2056 -79
rect -698 -107 -624 -96
rect -697 -113 -624 -107
rect 1977 -113 2056 -96
rect -697 -119 2056 -113
rect -697 -123 -631 -119
rect 535 -121 2056 -119
rect -697 -124 -646 -123
<< nsubdiff >>
rect 773 517 1909 523
rect 773 500 802 517
rect 1869 500 1909 517
rect 773 495 1909 500
rect 773 482 801 495
rect 773 23 778 482
rect 795 23 801 482
rect 1881 492 1909 495
rect 773 11 801 23
rect 1881 23 1886 492
rect 1903 23 1909 492
rect 1881 11 1909 23
rect 767 6 1909 11
rect 767 -11 808 6
rect 1875 -11 1909 6
rect 767 -17 1909 -11
<< psubdiffcont >>
rect -621 623 1966 640
rect -621 589 1966 606
rect -690 -55 -673 583
rect -656 -39 -639 570
rect 651 -44 668 570
rect 685 -45 702 568
rect 1993 -45 2010 577
rect 2031 -46 2048 573
rect -624 -79 1977 -62
rect -624 -113 1977 -96
<< nsubdiffcont >>
rect 802 500 1869 517
rect 778 23 795 482
rect 1886 23 1903 492
rect 808 -11 1875 6
<< poly >>
rect 32 796 49 807
rect 700 796 717 805
rect 23 790 73 796
rect 23 773 32 790
rect 49 773 73 790
rect 23 756 73 773
rect 23 739 32 756
rect 49 739 73 756
rect 23 722 73 739
rect 23 705 32 722
rect 49 705 73 722
rect 23 688 73 705
rect 23 671 32 688
rect 49 671 73 688
rect 23 664 73 671
rect 654 788 726 796
rect 654 771 700 788
rect 717 771 726 788
rect 654 754 726 771
rect 654 737 700 754
rect 717 737 726 754
rect 654 720 726 737
rect 654 703 700 720
rect 717 703 726 720
rect 654 686 726 703
rect 654 669 700 686
rect 717 669 726 686
rect 654 664 726 669
<< polycont >>
rect 32 773 49 790
rect 32 739 49 756
rect 32 705 49 722
rect 32 671 49 688
rect 700 771 717 788
rect 700 737 717 754
rect 700 703 717 720
rect 700 669 717 686
<< npolyres >>
rect 73 664 654 796
<< locali >>
rect 28 807 53 810
rect 28 671 32 807
rect 49 671 53 807
rect 28 664 53 671
rect 696 805 721 808
rect 696 669 700 805
rect 717 669 721 805
rect 32 663 49 664
rect 696 661 721 669
rect -690 624 -621 640
rect -690 606 -682 624
rect 1966 623 2048 640
rect -495 606 1654 623
rect -690 589 -621 606
rect 1970 605 2048 623
rect 1966 600 2048 605
rect 1966 589 2011 600
rect -690 583 -674 589
rect -656 588 -610 589
rect -656 570 -638 588
rect -673 -39 -656 397
rect -639 396 -638 570
rect -620 396 -610 588
rect 651 570 702 589
rect -552 544 -535 552
rect 572 544 595 553
rect -552 543 595 544
rect -553 526 -552 543
rect 593 526 595 543
rect -553 510 595 526
rect -553 493 -519 510
rect 579 493 595 510
rect -553 479 595 493
rect -553 462 -552 479
rect 593 462 595 479
rect -553 448 595 462
rect -553 431 -519 448
rect 579 431 595 448
rect -553 417 595 431
rect -553 400 -552 417
rect 592 400 595 417
rect -553 386 595 400
rect -553 369 -518 386
rect 580 369 595 386
rect -553 357 595 369
rect -553 340 -552 357
rect 593 340 595 357
rect -553 328 595 340
rect -553 311 -516 328
rect 582 311 595 328
rect -553 298 595 311
rect -553 281 -552 298
rect 593 281 595 298
rect -553 269 595 281
rect -553 252 -515 269
rect 583 252 595 269
rect -553 239 595 252
rect -553 222 -552 239
rect 593 222 595 239
rect -553 209 595 222
rect -553 192 -515 209
rect 583 192 595 209
rect -553 180 595 192
rect -553 163 -552 180
rect 592 163 595 180
rect -553 149 595 163
rect -553 132 -520 149
rect 578 132 595 149
rect -553 119 595 132
rect -553 102 -552 119
rect 593 102 595 119
rect -553 88 595 102
rect -553 71 -519 88
rect 579 71 595 88
rect -553 57 595 71
rect -553 40 -551 57
rect 593 40 595 57
rect -553 28 595 40
rect -553 11 -520 28
rect 578 11 595 28
rect -553 -4 595 11
rect -560 -21 -552 -4
rect 592 -21 595 -4
rect -553 -27 -534 -21
rect -673 -55 -639 -39
rect 572 -45 595 -21
rect 668 568 702 570
rect 668 -44 685 568
rect 651 -45 685 -44
rect 1993 577 2011 589
rect 778 500 802 517
rect 1869 500 1903 517
rect 778 482 795 500
rect 1886 492 1903 500
rect 834 467 1845 469
rect 834 463 1847 467
rect 829 446 839 463
rect 1819 446 1847 463
rect 834 434 1847 446
rect 834 417 854 434
rect 1799 417 1847 434
rect 834 396 1847 417
rect 834 379 844 396
rect 1813 379 1847 396
rect 834 359 1847 379
rect 834 342 853 359
rect 1792 342 1847 359
rect 834 323 1847 342
rect 834 306 849 323
rect 1824 306 1847 323
rect 834 287 1847 306
rect 834 270 856 287
rect 1796 270 1847 287
rect 834 255 1847 270
rect 834 238 848 255
rect 1816 238 1847 255
rect 834 221 1847 238
rect 834 204 857 221
rect 1794 204 1847 221
rect 834 188 1847 204
rect 834 171 844 188
rect 1818 171 1847 188
rect 834 156 1847 171
rect 834 139 856 156
rect 1801 139 1847 156
rect 834 124 1847 139
rect 834 107 843 124
rect 1816 107 1847 124
rect 834 92 1847 107
rect 834 75 857 92
rect 1796 75 1847 92
rect 834 62 1847 75
rect 834 45 845 62
rect 1816 45 1847 62
rect 834 44 1847 45
rect 834 36 1845 44
rect 778 13 795 23
rect 777 6 795 13
rect 1903 313 1947 324
rect 1903 23 1904 313
rect 1886 6 1904 23
rect 777 -11 808 6
rect 1875 -11 1904 6
rect 1893 -17 1904 -11
rect 1939 -17 1947 313
rect 1893 -22 1947 -17
rect -690 -62 -639 -55
rect -565 -62 -385 -61
rect 651 -62 702 -45
rect 2010 507 2011 577
rect 2031 573 2048 600
rect 2010 -45 2031 507
rect 1993 -46 2031 -45
rect 1992 -62 2048 -46
rect -690 -79 -624 -62
rect 1977 -79 2048 -62
rect -690 -96 2048 -79
rect -687 -113 -624 -96
rect 1977 -113 2048 -96
rect -687 -115 -618 -113
rect -567 -114 -387 -113
<< viali >>
rect 32 790 49 807
rect 32 756 49 773
rect 32 722 49 739
rect 32 688 49 705
rect 700 788 717 805
rect 700 754 717 771
rect 700 720 717 737
rect 700 686 717 703
rect -682 623 -621 624
rect -621 623 -496 624
rect -682 606 -495 623
rect 1654 606 1970 623
rect 1654 605 1966 606
rect 1966 605 1970 606
rect -674 583 -656 589
rect -674 510 -673 583
rect -673 397 -656 583
rect -638 396 -620 588
rect -519 493 579 510
rect -519 431 579 448
rect -518 369 580 386
rect -516 311 582 328
rect -515 252 583 269
rect -515 192 583 209
rect -520 132 578 149
rect -519 71 579 88
rect -520 11 578 28
rect 854 417 1799 434
rect 853 342 1792 359
rect 856 270 1796 287
rect 857 204 1794 221
rect 856 139 1801 156
rect 857 75 1796 92
rect 1904 -17 1939 313
rect 2011 507 2031 600
<< metal1 >>
rect 26 807 416 858
rect 26 790 32 807
rect 49 799 416 807
rect 690 805 725 811
rect 49 790 55 799
rect 690 796 700 805
rect 26 773 55 790
rect 26 756 32 773
rect 49 756 55 773
rect 26 739 55 756
rect 26 722 32 739
rect 49 722 55 739
rect 26 705 55 722
rect 26 688 32 705
rect 49 688 55 705
rect 689 788 700 796
rect 717 796 725 805
rect 717 788 726 796
rect 689 771 726 788
rect 689 754 700 771
rect 717 754 726 771
rect 689 737 726 754
rect 689 720 700 737
rect 717 720 726 737
rect 689 703 726 720
rect 689 701 700 703
rect 644 700 700 701
rect 26 664 55 688
rect 511 686 700 700
rect 717 701 726 703
rect 717 686 901 701
rect 511 664 901 686
rect -701 632 -464 647
rect -701 624 -679 632
rect -701 606 -682 624
rect -701 599 -679 606
rect -476 599 -464 632
rect -701 589 -464 599
rect -701 584 -674 589
rect -698 575 -674 584
rect -656 588 -464 589
rect -656 575 -638 588
rect -620 584 -464 588
rect -620 575 -603 584
rect -528 582 -470 584
rect -698 513 -685 575
rect -615 513 -603 575
rect 510 518 901 664
rect 1633 634 2046 639
rect 1633 623 1660 634
rect 1959 623 2046 634
rect 1633 605 1654 623
rect 1970 605 2046 623
rect 1633 599 1660 605
rect 1959 600 2046 605
rect 1959 599 2011 600
rect 1633 595 2011 599
rect 2031 599 2046 600
rect 2031 595 2047 599
rect 1633 590 2003 595
rect -461 517 901 518
rect -698 510 -674 513
rect -698 397 -673 510
rect -656 397 -638 513
rect -698 396 -638 397
rect -620 396 -603 513
rect -698 388 -603 396
rect -675 -179 -603 388
rect -528 510 901 517
rect -528 493 -519 510
rect 579 493 901 510
rect 1994 519 2003 590
rect 2038 519 2047 595
rect 1994 507 2011 519
rect 2031 507 2047 519
rect 1994 500 2047 507
rect -528 461 901 493
rect -528 448 1807 461
rect -528 431 -519 448
rect 579 434 1807 448
rect 579 431 854 434
rect -528 417 854 431
rect 1799 417 1807 434
rect -528 386 1807 417
rect -528 369 -518 386
rect 580 369 1807 386
rect -528 359 1807 369
rect -528 342 853 359
rect 1792 342 1807 359
rect -528 328 1807 342
rect -528 311 -516 328
rect 582 311 1807 328
rect -528 287 1807 311
rect -528 270 856 287
rect 1796 270 1807 287
rect -528 269 1807 270
rect -528 252 -515 269
rect 583 252 1807 269
rect -528 221 1807 252
rect -528 209 857 221
rect -528 192 -515 209
rect 583 204 857 209
rect 1794 204 1807 221
rect 583 192 1807 204
rect -528 156 1807 192
rect -528 149 856 156
rect -528 132 -520 149
rect 578 139 856 149
rect 1801 139 1807 156
rect 578 132 1807 139
rect -528 92 1807 132
rect -528 88 857 92
rect -528 71 -519 88
rect 579 75 857 88
rect 1796 75 1807 92
rect 579 71 1807 75
rect -528 31 1807 71
rect 1884 319 1941 320
rect 1884 313 1946 319
rect 1884 307 1904 313
rect 1939 307 1946 313
rect -528 28 901 31
rect -528 11 -520 28
rect 578 11 901 28
rect -528 3 901 11
rect 510 -152 901 3
rect 1884 -10 1900 307
rect 1942 -10 1946 307
rect 1884 -17 1904 -10
rect 1939 -17 1946 -10
rect 1884 -23 1946 -17
rect 1884 -24 1941 -23
rect 1801 -140 1857 -137
rect 508 -229 903 -152
rect 1801 -187 1803 -140
rect 1802 -192 1803 -187
rect 1855 -192 1857 -140
rect 1802 -209 1857 -192
<< via1 >>
rect -679 624 -476 632
rect -679 623 -496 624
rect -496 623 -476 624
rect -679 606 -495 623
rect -495 606 -476 623
rect -679 599 -476 606
rect -685 513 -674 575
rect -674 513 -656 575
rect -656 513 -638 575
rect -638 513 -620 575
rect -620 513 -615 575
rect 1660 623 1959 634
rect 1660 605 1959 623
rect 1660 599 1959 605
rect 2003 519 2011 595
rect 2011 519 2031 595
rect 2031 519 2038 595
rect 1900 -10 1904 307
rect 1904 -10 1939 307
rect 1939 -10 1942 307
rect 1803 -192 1855 -140
<< metal2 >>
rect -745 634 2114 649
rect -745 632 1660 634
rect -745 599 -679 632
rect -476 599 1660 632
rect 1959 599 2114 634
rect -745 595 2114 599
rect -745 575 2003 595
rect -745 513 -685 575
rect -615 519 2003 575
rect 2038 519 2114 595
rect -615 513 2114 519
rect -745 509 2114 513
rect -698 508 -605 509
rect -673 397 -656 508
rect 1889 307 1953 320
rect 1889 19 1900 307
rect -745 -10 1900 19
rect 1942 19 1953 307
rect 1942 -10 2114 19
rect -745 -121 2114 -10
rect 1799 -134 2062 -121
rect 1799 -140 2054 -134
rect 1799 -192 1803 -140
rect 1855 -185 2054 -140
rect 1855 -192 1861 -185
<< labels >>
rlabel metal1 508 -229 903 -152 0 OUTPUT 
port 2 nsew
rlabel space -744 508 -721 649 0 VGND
port 3 nsew
rlabel metal2 2078 509 2114 649 0 VGND
port 3 nsew
rlabel metal2 -744 -121 -723 19 0 VINJ
port 4 nsew
rlabel metal2 2084 -121 2114 19 0 VINJ
port 4 nsew
rlabel metal1 26 811 415 858 0 INPUT
port 5 nsew
rlabel metal2 1875 -185 2054 -160 0 VINJ
port 4 nsew
rlabel metal1 -675 -179 -603 -145 0 VGND
port 3 nsew
<< end >>
