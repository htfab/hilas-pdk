* NGSPICE file created from /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_capacitorSize04.ext - technology: sky130A

.subckt sky130_hilas_CapModule01a VSUBS m3_n832_n432# c1_n802_n404#
X0 c1_n802_n404# m3_n832_n432# sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
.ends

.subckt home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_capacitorSize04
+ Cap1Term02 Cap2Term02 Cap2Term01 Cap1Term01
Xsky130_hilas_CapModule01a_0 VSUBS Cap2Term02 Cap2Term01 sky130_hilas_CapModule01a
Xsky130_hilas_CapModule01a_1 VSUBS Cap1Term02 Cap1Term01 sky130_hilas_CapModule01a
.ends

