magic
tech sky130A
timestamp 1628707346
<< nwell >>
rect 1 0 345 164
<< mvnmos >>
rect 513 95 563 127
rect 442 34 492 65
rect 584 34 634 65
<< mvpmos >>
rect 159 97 211 131
rect 85 33 138 66
rect 232 34 284 66
<< mvndiff >>
rect 482 119 513 127
rect 482 102 489 119
rect 506 102 513 119
rect 482 95 513 102
rect 563 119 590 127
rect 563 102 569 119
rect 586 102 590 119
rect 563 95 590 102
rect 413 58 442 65
rect 413 41 418 58
rect 435 41 442 58
rect 413 34 442 41
rect 492 58 520 65
rect 492 41 498 58
rect 515 41 520 58
rect 492 34 520 41
rect 556 58 584 65
rect 556 41 561 58
rect 578 41 584 58
rect 556 34 584 41
rect 634 58 663 65
rect 634 41 640 58
rect 657 41 663 58
rect 634 34 663 41
<< mvpdiff >>
rect 131 123 159 131
rect 131 106 136 123
rect 153 106 159 123
rect 131 97 159 106
rect 211 123 239 131
rect 211 106 217 123
rect 234 106 239 123
rect 211 97 239 106
rect 58 58 85 66
rect 58 41 62 58
rect 79 41 85 58
rect 58 33 85 41
rect 138 58 166 66
rect 138 41 144 58
rect 161 41 166 58
rect 138 33 166 41
rect 205 58 232 66
rect 205 41 209 58
rect 226 41 232 58
rect 205 34 232 41
rect 284 58 311 66
rect 284 41 290 58
rect 307 41 311 58
rect 284 34 311 41
<< mvndiffc >>
rect 489 102 506 119
rect 569 102 586 119
rect 418 41 435 58
rect 498 41 515 58
rect 561 41 578 58
rect 640 41 657 58
<< mvpdiffc >>
rect 136 106 153 123
rect 217 106 234 123
rect 62 41 79 58
rect 144 41 161 58
rect 209 41 226 58
rect 290 41 307 58
<< psubdiff >>
rect 629 120 670 127
rect 629 103 641 120
rect 658 103 670 120
rect 629 95 670 103
<< mvnsubdiff >>
rect 51 123 92 131
rect 51 106 63 123
rect 80 106 92 123
rect 51 97 92 106
<< psubdiffcont >>
rect 641 103 658 120
<< mvnsubdiffcont >>
rect 63 106 80 123
<< poly >>
rect 194 145 531 151
rect 159 140 531 145
rect 159 134 563 140
rect 159 131 211 134
rect 362 131 397 134
rect 362 114 371 131
rect 388 114 397 131
rect 513 127 563 134
rect 263 107 298 113
rect 362 107 397 114
rect 15 82 101 83
rect 15 68 138 82
rect 159 81 211 97
rect 263 90 273 107
rect 290 90 298 107
rect 263 86 298 90
rect 263 81 460 86
rect 513 81 563 95
rect 15 58 42 68
rect 85 66 138 68
rect 232 79 460 81
rect 232 69 492 79
rect 232 66 284 69
rect 15 41 20 58
rect 37 41 42 58
rect 15 33 42 41
rect 442 65 492 69
rect 584 65 634 79
rect 85 20 138 33
rect 232 21 284 34
rect 442 21 492 34
rect 584 21 634 34
<< polycont >>
rect 371 114 388 131
rect 273 90 290 107
rect 20 41 37 58
<< locali >>
rect 63 123 80 135
rect 371 131 388 139
rect 136 123 153 131
rect 217 123 234 131
rect 63 104 65 106
rect 153 106 157 123
rect 63 94 80 104
rect 136 66 157 106
rect 213 106 217 123
rect 213 98 234 106
rect 273 107 290 115
rect 560 120 586 127
rect 640 120 658 133
rect 560 119 641 120
rect 384 110 388 114
rect 371 106 388 110
rect 213 66 230 98
rect 287 88 290 90
rect 273 78 290 88
rect 427 102 489 119
rect 506 102 514 119
rect 560 102 569 119
rect 586 103 641 119
rect 586 102 658 103
rect 20 58 37 66
rect 35 39 37 41
rect 20 33 37 39
rect 62 60 79 66
rect 62 58 87 60
rect 79 53 87 58
rect 62 36 66 41
rect 83 36 87 53
rect 136 58 161 66
rect 136 41 144 58
rect 62 33 87 36
rect 63 31 87 33
rect 144 32 161 41
rect 209 58 230 66
rect 427 58 444 102
rect 560 88 586 102
rect 640 91 658 102
rect 560 70 563 88
rect 581 70 586 88
rect 560 58 586 70
rect 226 41 230 58
rect 281 41 290 58
rect 307 54 418 58
rect 307 41 358 54
rect 209 33 226 41
rect 375 41 418 54
rect 435 41 444 58
rect 489 41 498 58
rect 515 41 561 58
rect 578 41 586 58
rect 631 41 640 58
rect 657 41 665 58
<< viali >>
rect 65 106 80 121
rect 80 106 82 121
rect 65 104 82 106
rect 367 114 371 127
rect 371 114 384 127
rect 367 110 384 114
rect 270 90 273 105
rect 273 90 287 105
rect 270 88 287 90
rect 18 41 20 56
rect 20 41 35 56
rect 18 39 35 41
rect 66 41 79 53
rect 79 41 83 53
rect 66 36 83 41
rect 563 70 581 88
rect 358 37 375 54
<< metal1 >>
rect 62 126 84 160
rect 62 121 85 126
rect 62 104 65 121
rect 82 104 85 121
rect 62 100 85 104
rect 9 61 40 67
rect 9 35 12 61
rect 38 35 40 61
rect 9 32 40 35
rect 62 60 84 100
rect 264 84 268 110
rect 294 84 297 110
rect 361 109 367 135
rect 393 109 404 135
rect 361 106 404 109
rect 559 88 586 161
rect 559 70 563 88
rect 581 70 586 88
rect 62 53 87 60
rect 62 36 66 53
rect 83 36 87 53
rect 62 29 87 36
rect 348 57 387 58
rect 348 31 354 57
rect 380 31 387 57
rect 62 9 84 29
rect 559 9 586 70
rect 641 61 672 64
rect 641 35 644 61
rect 670 35 672 61
rect 641 32 672 35
<< via1 >>
rect 12 56 38 61
rect 12 39 18 56
rect 18 39 35 56
rect 35 39 38 56
rect 12 35 38 39
rect 268 105 294 110
rect 268 88 270 105
rect 270 88 287 105
rect 287 88 294 105
rect 268 84 294 88
rect 367 127 393 135
rect 367 110 384 127
rect 384 110 393 127
rect 367 109 393 110
rect 354 54 380 57
rect 354 37 358 54
rect 358 37 375 54
rect 375 37 380 54
rect 354 31 380 37
rect 644 35 670 61
<< metal2 >>
rect 0 135 404 145
rect 0 129 367 135
rect 264 102 268 110
rect 237 100 268 102
rect 1 84 268 100
rect 294 84 297 110
rect 362 109 367 129
rect 393 109 404 135
rect 362 106 404 109
rect 641 61 672 64
rect 9 51 12 61
rect 1 35 12 51
rect 38 35 41 61
rect 350 31 354 57
rect 380 49 387 57
rect 380 48 453 49
rect 641 48 644 61
rect 380 35 644 48
rect 670 48 672 61
rect 670 35 688 48
rect 380 31 688 35
<< labels >>
rlabel metal2 682 31 688 48 0 Output
rlabel metal2 0 129 6 145 0 Input1
rlabel space 0 84 6 100 0 Input2
rlabel space 0 35 6 51 0 Input3
rlabel metal1 559 155 586 161 0 GND
rlabel metal1 559 9 586 14 0 GND
rlabel metal1 62 9 84 15 0 Vinj
rlabel metal1 62 153 84 160 0 Vinj
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
