magic
tech sky130A
timestamp 1628704213
<< nwell >>
rect 0 0 203 99
<< pmos >>
rect 103 36 142 78
<< pdiff >>
rect 75 64 103 78
rect 75 47 80 64
rect 97 47 103 64
rect 75 36 103 47
rect 142 64 169 78
rect 142 47 148 64
rect 165 47 169 64
rect 142 36 169 47
<< pdiffc >>
rect 80 47 97 64
rect 148 47 165 64
<< poly >>
rect 103 78 142 91
rect 41 28 67 36
rect 103 28 142 36
rect 41 13 142 28
<< locali >>
rect 66 64 97 72
rect 66 54 80 64
rect 64 52 80 54
rect 80 39 97 47
rect 148 64 165 72
rect 148 39 165 47
<< metal2 >>
rect 0 52 37 71
rect 0 10 38 29
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628285143
transform 1 0 178 0 1 54
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628285143
transform 1 0 48 0 1 64
box -14 -15 20 18
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_0
timestamp 1628285143
transform 0 1 34 -1 0 27
box -9 -26 24 29
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
