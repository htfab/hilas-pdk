VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_Tgate4Single01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_Tgate4Single01 ;
  ORIGIN 0.360 1.410 ;
  SIZE 4.760 BY 6.050 ;
  PIN Input1_4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -0.360 -1.300 1.310 -1.100 ;
    END
  END Input1_4
  PIN Vdd
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 0.380 -1.410 0.580 -0.480 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.380 3.710 0.580 4.640 ;
    END
  END Vdd
  PIN Select4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -0.360 -0.320 -0.040 -0.120 ;
    END
  END Select4
  PIN Select3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -0.360 0.330 -0.040 0.530 ;
    END
  END Select3
  PIN Input1_3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -0.360 1.310 1.310 1.510 ;
    END
  END Input1_3
  PIN Input1_2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -0.360 1.720 1.310 1.920 ;
    END
  END Input1_2
  PIN Select2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -0.360 2.700 -0.040 2.900 ;
    END
  END Select2
  PIN Select1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -0.360 3.350 -0.040 3.550 ;
    END
  END Select1
  PIN Input1_1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -0.360 4.330 1.310 4.530 ;
    END
  END Input1_1
  PIN GND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 3.890 3.710 4.080 4.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.890 -1.410 4.080 -0.480 ;
    END
  END GND
  PIN Output1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 3.500 3.350 4.400 3.550 ;
    END
  END Output1
  PIN Output2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 3.500 2.700 4.400 2.900 ;
    END
  END Output2
  PIN Output3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 3.500 0.330 4.400 0.530 ;
    END
  END Output3
  PIN Output4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 3.500 -0.320 4.400 -0.120 ;
    END
  END Output4
  OBS
      LAYER li1 ;
        RECT -0.120 -1.270 4.320 4.500 ;
      LAYER met1 ;
        RECT -0.130 3.430 0.100 4.530 ;
        RECT 0.860 3.430 3.610 4.530 ;
        RECT -0.130 -0.200 4.100 3.430 ;
        RECT -0.130 -1.300 0.100 -0.200 ;
        RECT 0.860 -1.300 3.610 -0.200 ;
      LAYER met2 ;
        RECT 1.590 4.050 3.530 4.540 ;
        RECT -0.070 3.830 3.530 4.050 ;
        RECT 0.240 2.420 3.220 3.830 ;
        RECT -0.070 2.200 3.530 2.420 ;
        RECT 1.590 1.030 3.530 2.200 ;
        RECT -0.070 0.810 3.530 1.030 ;
        RECT 0.240 -0.600 3.220 0.810 ;
        RECT -0.070 -0.820 3.530 -0.600 ;
        RECT 1.590 -1.310 3.530 -0.820 ;
  END
END sky130_hilas_Tgate4Single01
END LIBRARY

