magic
tech sky130A
timestamp 1627061166
<< error_s >>
rect 432 542 438 548
rect 537 542 543 548
rect 58 532 64 538
rect 111 532 117 538
rect 52 482 58 488
rect 117 482 123 488
rect 426 478 432 484
rect 543 478 549 484
rect 58 423 64 429
rect 111 423 117 429
rect 432 425 438 431
rect 537 425 543 431
rect 52 373 58 379
rect 117 373 123 379
rect 426 361 432 367
rect 543 361 549 367
rect 432 240 438 246
rect 537 240 543 246
rect 58 234 64 240
rect 111 234 117 240
rect 52 184 58 190
rect 117 184 123 190
rect 426 176 432 182
rect 543 176 549 182
rect 432 124 438 130
rect 537 124 543 130
rect 58 117 64 123
rect 111 117 117 123
rect 52 67 58 73
rect 117 67 123 73
rect 426 60 432 66
rect 543 60 549 66
<< nwell >>
rect 376 604 599 605
rect 1 494 8 512
rect 896 310 931 311
rect 896 294 913 310
rect 930 294 931 310
rect 441 1 479 9
rect 376 0 599 1
<< psubdiff >>
rect 279 464 305 487
rect 279 447 283 464
rect 300 447 305 464
rect 279 421 305 447
rect 671 463 698 489
rect 671 446 677 463
rect 694 446 698 463
rect 671 423 698 446
rect 280 352 305 379
rect 280 335 284 352
rect 301 335 305 352
rect 280 318 305 335
rect 280 301 284 318
rect 301 301 305 318
rect 280 284 305 301
rect 280 267 284 284
rect 301 267 305 284
rect 280 239 305 267
rect 673 338 698 365
rect 673 321 677 338
rect 694 321 698 338
rect 673 304 698 321
rect 673 287 677 304
rect 694 287 698 304
rect 673 270 698 287
rect 673 253 677 270
rect 694 253 698 270
rect 673 240 698 253
<< psubdiffcont >>
rect 283 447 300 464
rect 677 446 694 463
rect 284 335 301 352
rect 284 301 301 318
rect 284 267 301 284
rect 677 321 694 338
rect 677 287 694 304
rect 677 253 694 270
<< poly >>
rect 583 529 753 533
rect 157 496 394 520
rect 583 517 752 529
rect 157 387 392 411
rect 583 373 752 390
rect 913 310 931 311
rect 929 294 931 310
rect 157 207 394 231
rect 584 215 752 232
rect 159 87 396 111
rect 584 73 752 90
<< polycont >>
rect 896 294 913 311
<< locali >>
rect 284 352 301 360
rect 284 259 301 267
rect 677 338 694 346
rect 887 294 896 311
rect 677 245 694 253
<< viali >>
rect 283 464 300 481
rect 283 430 300 447
rect 677 463 694 480
rect 677 429 694 446
rect 284 318 301 335
rect 284 284 301 301
rect 677 304 694 321
rect 913 294 931 311
rect 677 270 694 287
<< metal1 >>
rect 36 0 76 605
rect 280 487 304 605
rect 441 595 479 605
rect 673 489 697 605
rect 875 601 891 605
rect 912 600 931 605
rect 956 600 972 605
rect 279 481 305 487
rect 279 464 283 481
rect 300 464 305 481
rect 279 447 305 464
rect 279 430 283 447
rect 300 430 305 447
rect 279 421 305 430
rect 671 480 698 489
rect 671 463 677 480
rect 694 463 698 480
rect 671 446 698 463
rect 671 429 677 446
rect 694 429 698 446
rect 671 423 698 429
rect 280 335 304 421
rect 280 318 284 335
rect 301 318 304 335
rect 280 301 304 318
rect 280 284 284 301
rect 301 284 304 301
rect 280 160 304 284
rect 673 321 697 423
rect 673 304 677 321
rect 694 304 697 321
rect 918 314 931 316
rect 673 287 697 304
rect 910 311 934 314
rect 910 294 913 311
rect 931 294 934 311
rect 910 291 934 294
rect 920 287 931 291
rect 673 270 677 287
rect 694 270 697 287
rect 673 164 697 270
rect 672 161 698 164
rect 279 157 305 160
rect 672 132 698 135
rect 279 128 305 131
rect 280 0 304 128
rect 441 0 479 9
rect 673 0 697 132
<< via1 >>
rect 279 131 305 157
rect 672 135 698 161
<< metal2 >>
rect 1 548 761 555
rect 1 537 764 548
rect 1 494 974 512
rect 0 406 761 412
rect 0 394 764 406
rect 0 351 764 369
rect 2 236 764 253
rect 2 194 764 211
rect 669 161 701 164
rect 276 131 279 157
rect 305 156 308 157
rect 669 156 672 161
rect 305 138 672 156
rect 305 131 308 138
rect 669 135 672 138
rect 698 135 701 161
rect 669 132 701 135
rect 2 96 764 113
rect 80 87 234 96
rect 2 52 764 69
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_0
timestamp 1608066871
transform 1 0 1452 0 1 517
box -1451 -400 -1278 -210
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_1
timestamp 1608066871
transform 1 0 1452 0 1 400
box -1451 -400 -1278 -210
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_0
timestamp 1606741561
transform 1 0 1333 0 1 396
box -957 -395 -734 -209
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_1
timestamp 1606741561
transform 1 0 1333 0 1 512
box -957 -395 -734 -209
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_1
timestamp 1607386385
transform 1 0 1041 0 1 -46
box -289 47 -33 232
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_2
timestamp 1607386385
transform 1 0 1041 0 -1 351
box -289 47 -33 232
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_2
timestamp 1608066871
transform 1 0 1452 0 1 706
box -1451 -400 -1278 -210
use sky130_hilas_wellContact  sky130_hilas_wellContact_1
timestamp 1606753443
transform 1 0 1449 0 1 675
box -1449 -441 -1275 -255
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_2
timestamp 1606741561
transform 1 0 1333 0 1 697
box -957 -395 -734 -209
use sky130_hilas_wellContact  sky130_hilas_wellContact_0
timestamp 1606753443
transform 1 0 1852 0 1 668
box -1449 -441 -1275 -255
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_0
timestamp 1607386385
transform 1 0 1041 0 1 254
box -289 47 -33 232
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_3
timestamp 1608066871
transform 1 0 1452 0 1 815
box -1451 -400 -1278 -210
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_3
timestamp 1606741561
transform 1 0 1333 0 1 814
box -957 -395 -734 -209
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_3
timestamp 1607386385
transform 1 0 1041 0 -1 652
box -289 47 -33 232
<< labels >>
rlabel metal1 36 593 76 605 0 VTUN
port 1 nsew
rlabel metal1 956 600 972 605 0 VINJ
port 2 nsew
rlabel metal1 912 600 931 605 0 COLSEL1
port 3 nsew
rlabel metal1 875 601 891 605 0 COL1
port 4 nsew
rlabel metal1 441 595 479 605 0 GATE1
port 5 nsew
rlabel poly 647 518 658 531 0 FG1
rlabel poly 636 373 653 388 0 FG2
rlabel poly 643 216 660 231 0 FG3
rlabel poly 653 75 670 90 0 FG4
rlabel metal2 1 537 8 555 0 DRAIN1
port 6 nsew
rlabel metal2 0 394 7 412 0 ROW2
port 9 nsew
rlabel metal2 0 351 7 369 0 DRAIN2
port 8 nsew
rlabel metal2 2 236 8 253 0 DRAIN3
port 10 nsew
rlabel metal2 2 194 8 211 0 ROW3
port 7 nsew
rlabel metal2 2 96 8 113 0 ROW4
port 11 nsew
rlabel metal2 2 52 8 69 0 DRAIN4
port 12 nsew
rlabel metal2 1 494 8 512 0 ROW1
port 13 nsew
rlabel metal1 280 600 304 605 0 VGND
port 14 nsew
rlabel metal1 673 600 697 605 0 VGND
port 14 nsew
rlabel metal1 673 0 697 6 0 VGND
port 14 nsew
rlabel metal1 280 0 304 6 0 VGND
port 14 nsew
rlabel metal1 441 0 479 9 0 GATE1
port 5 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
