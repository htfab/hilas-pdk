magic
tech sky130A
timestamp 1606663783
<< error_p >>
rect -1466 227 -1381 259
rect -1393 135 -1387 141
rect -1341 135 -1335 141
rect -1399 77 -1393 83
rect -1335 77 -1329 83
rect -869 77 -863 83
rect -820 77 -814 83
rect -772 54 -769 77
rect -1393 25 -1387 31
rect -1341 25 -1335 31
rect -875 4 -869 10
rect -814 4 -808 10
rect -772 4 -769 27
rect -324 16 -298 238
rect -1399 -32 -1393 -26
rect -1335 -32 -1329 -26
rect -873 -51 -872 -47
rect -873 -72 -867 -66
rect -820 -72 -814 -66
rect -1393 -83 -1387 -77
rect -1341 -83 -1335 -77
rect -1400 -133 -1393 -127
rect -1335 -133 -1329 -127
rect -879 -147 -873 -141
rect -814 -147 -808 -141
rect -471 -175 -451 -167
rect -1394 -183 -1388 -177
rect -1341 -183 -1335 -177
rect -1400 -233 -1394 -227
rect -1335 -233 -1329 -227
rect -900 -244 -875 -223
rect -900 -248 -869 -244
rect -806 -248 -800 -242
rect -900 -275 -875 -248
rect -1394 -283 -1388 -277
rect -1341 -283 -1335 -277
rect -1400 -333 -1394 -327
rect -1335 -333 -1329 -327
rect -884 -362 -875 -344
rect -866 -362 -865 -361
rect -800 -362 -794 -356
rect -778 -362 -775 -250
rect -916 -364 -875 -362
rect -867 -363 -775 -362
rect -866 -364 -775 -363
rect -891 -387 -875 -364
rect -521 -408 -491 -407
rect -554 -441 -507 -440
rect -425 -442 -423 -356
<< nwell >>
rect -1466 175 -1275 227
rect -1465 -440 -1275 175
rect -992 26 -713 224
rect -994 -253 -712 26
rect -990 -440 -712 -253
rect -572 -440 -425 226
rect -324 17 2 238
rect -324 16 -2 17
rect -507 -442 -425 -440
<< mvpmos >>
rect -521 116 -491 166
rect -222 143 -172 173
rect -222 81 -172 112
rect -150 81 -100 112
rect -521 -21 -491 30
rect -521 -94 -491 -42
rect -521 -175 -491 -123
rect -521 -246 -491 -196
rect -521 -381 -491 -331
<< mvvaractor >>
rect -1393 77 -1335 135
rect -1393 -32 -1335 25
rect -869 4 -814 77
rect -1393 -133 -1335 -83
rect -873 -147 -814 -72
rect -1394 -233 -1335 -183
rect -1394 -333 -1335 -283
rect -875 -362 -800 -248
rect -875 -364 -866 -362
<< mvpdiff >>
rect -521 189 -491 193
rect -521 172 -515 189
rect -497 172 -491 189
rect -521 166 -491 172
rect -256 167 -222 173
rect -256 150 -247 167
rect -229 150 -222 167
rect -256 143 -222 150
rect -172 166 -141 173
rect -172 149 -165 166
rect -146 149 -141 166
rect -172 143 -141 149
rect -521 110 -491 116
rect -521 93 -515 110
rect -497 93 -491 110
rect -521 88 -491 93
rect -256 105 -222 112
rect -256 88 -247 105
rect -229 88 -222 105
rect -256 81 -222 88
rect -172 81 -150 112
rect -100 105 -66 112
rect -100 88 -93 105
rect -73 88 -66 105
rect -100 81 -66 88
rect -521 53 -491 58
rect -521 36 -515 53
rect -497 36 -491 53
rect -521 30 -491 36
rect -521 -42 -491 -21
rect -521 -100 -491 -94
rect -521 -117 -515 -100
rect -497 -117 -491 -100
rect -521 -123 -491 -117
rect -521 -196 -491 -175
rect -521 -252 -491 -246
rect -521 -269 -515 -252
rect -497 -269 -491 -252
rect -521 -273 -491 -269
rect -521 -308 -491 -304
rect -521 -325 -515 -308
rect -497 -325 -491 -308
rect -521 -331 -491 -325
rect -521 -387 -491 -381
rect -521 -404 -515 -387
rect -497 -404 -491 -387
rect -521 -408 -491 -404
<< mvpdiffc >>
rect -515 172 -497 189
rect -247 150 -229 167
rect -165 149 -146 166
rect -515 93 -497 110
rect -247 88 -229 105
rect -93 88 -73 105
rect -515 36 -497 53
rect -515 -117 -497 -100
rect -515 -269 -497 -252
rect -515 -325 -497 -308
rect -515 -404 -497 -387
<< psubdiff >>
rect -656 -361 -630 -349
rect -656 -378 -652 -361
rect -634 -378 -630 -361
rect -656 -390 -630 -378
<< mvnsubdiff >>
rect -1393 135 -1335 182
rect -869 77 -814 191
rect -1393 25 -1335 77
rect -100 183 -67 187
rect -100 169 -66 183
rect -100 151 -93 169
rect -73 151 -66 169
rect -100 139 -66 151
rect -1393 -83 -1335 -32
rect -869 -43 -814 4
rect -872 -51 -814 -43
rect -873 -72 -814 -51
rect -1394 -183 -1335 -133
rect -873 -190 -814 -147
rect -1394 -283 -1335 -233
rect -875 -248 -800 -190
rect -1394 -360 -1335 -333
rect -1394 -387 -1379 -360
rect -1351 -387 -1335 -360
rect -866 -364 -800 -362
rect -1394 -397 -1335 -387
rect -875 -403 -800 -364
<< psubdiffcont >>
rect -652 -378 -634 -361
<< mvnsubdiffcont >>
rect -93 151 -73 169
rect -1379 -387 -1351 -360
<< poly >>
rect -1436 77 -1393 135
rect -1335 77 -1292 135
rect -222 173 -172 187
rect -555 166 -534 168
rect -555 116 -521 166
rect -491 116 -478 166
rect -915 54 -869 77
rect -951 27 -869 54
rect -1435 -32 -1393 25
rect -1335 -32 -1292 25
rect -915 4 -869 27
rect -814 54 -772 77
rect -814 27 -743 54
rect -555 30 -534 116
rect -222 112 -172 143
rect -137 127 -117 187
rect -150 112 -100 127
rect -222 66 -172 81
rect -150 67 -100 81
rect -814 4 -772 27
rect -555 -21 -521 30
rect -491 -21 -476 30
rect -1435 -133 -1393 -83
rect -1335 -133 -1291 -83
rect -915 -147 -873 -72
rect -814 -147 -771 -72
rect -535 -94 -521 -42
rect -491 -94 -447 -42
rect -471 -123 -447 -94
rect -1436 -233 -1394 -183
rect -1335 -233 -1292 -183
rect -534 -175 -521 -123
rect -491 -167 -447 -123
rect -491 -175 -472 -167
rect -471 -175 -447 -167
rect -534 -246 -521 -196
rect -491 -246 -472 -196
rect -1436 -333 -1394 -283
rect -1335 -333 -1292 -283
rect -927 -364 -875 -250
rect -800 -362 -778 -248
rect -537 -381 -521 -331
rect -491 -381 -475 -331
<< locali >>
rect -523 172 -515 189
rect -497 172 -489 189
rect -256 150 -247 167
rect -229 150 -221 167
rect -166 166 -146 175
rect -166 149 -165 166
rect -166 141 -146 149
rect -93 169 -73 180
rect -523 93 -515 110
rect -497 93 -489 110
rect -93 105 -73 151
rect -256 88 -247 105
rect -229 88 -221 105
rect -93 80 -73 88
rect -523 36 -515 53
rect -497 36 -489 53
rect -524 -117 -515 -100
rect -497 -117 -489 -100
rect -523 -269 -515 -252
rect -497 -269 -489 -252
rect -523 -325 -515 -308
rect -497 -325 -489 -308
rect -1379 -360 -1351 -352
rect -660 -378 -652 -361
rect -634 -378 -626 -361
rect -1379 -395 -1351 -387
rect -523 -404 -515 -387
rect -497 -404 -489 -387
<< end >>
