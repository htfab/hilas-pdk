magic
tech sky130A
timestamp 1627737364
<< error_s >>
rect -2549 711 -2499 722
rect -2477 711 -2427 722
rect -509 711 -459 722
rect -437 711 -387 722
rect -49 717 -22 724
rect 154 704 171 709
rect -2427 680 -2393 681
rect -543 680 -509 681
rect -2549 669 -2499 680
rect -2477 669 -2427 680
rect -509 669 -459 680
rect -437 669 -387 680
rect -49 675 -22 682
rect -49 651 -22 658
rect -2485 648 -2476 650
rect -2425 648 -2393 650
rect -2361 648 -2322 650
rect -2226 648 -2186 650
rect -750 648 -710 650
rect -614 648 -575 650
rect -543 648 -511 650
rect -460 648 -451 650
rect -2188 640 -2186 648
rect -2504 544 -2499 585
rect -2364 573 -2361 623
rect -2322 573 -2319 623
rect -2228 573 -2226 623
rect -2186 573 -2184 623
rect -752 573 -750 623
rect -710 573 -708 623
rect -617 573 -614 623
rect -575 573 -572 623
rect -49 609 -22 616
rect -437 561 -432 585
rect -49 569 -22 576
rect -413 544 -408 561
rect -2364 494 -2361 544
rect -2322 494 -2319 544
rect -2228 494 -2226 544
rect -2186 494 -2184 544
rect -752 494 -750 544
rect -710 494 -708 544
rect -617 494 -614 544
rect -575 494 -572 544
rect -49 527 -22 534
rect -49 503 -22 510
rect -1766 463 -1749 464
rect -1187 463 -1170 464
rect -49 461 -22 468
rect -1766 444 -1749 445
rect -1187 444 -1170 445
rect -1766 428 -1749 430
rect -1187 428 -1170 430
rect -49 421 -22 428
rect -1765 409 -1748 411
rect -1187 409 -1170 411
rect -2504 324 -2499 365
rect -2364 341 -2361 391
rect -2322 341 -2319 391
rect -2228 341 -2226 391
rect -2186 341 -2184 391
rect -752 341 -750 391
rect -710 341 -708 391
rect -617 341 -614 391
rect -575 341 -572 391
rect -49 379 -22 386
rect -437 341 -432 365
rect -49 355 -22 362
rect -413 324 -408 341
rect -49 313 -22 320
rect -2364 262 -2361 312
rect -2322 262 -2319 312
rect -2228 262 -2226 312
rect -2186 262 -2184 312
rect -752 262 -750 312
rect -710 262 -708 312
rect -617 262 -614 312
rect -575 262 -572 312
rect -49 273 -22 280
rect -2485 235 -2476 237
rect -2425 235 -2393 237
rect -2361 235 -2322 237
rect -2226 235 -2186 237
rect -750 235 -710 237
rect -614 235 -575 237
rect -543 235 -511 237
rect -460 235 -451 237
rect -49 231 -22 238
rect -2549 205 -2499 216
rect -2477 205 -2427 216
rect -509 205 -459 216
rect -437 205 -387 216
rect -49 207 -22 214
rect -2427 204 -2393 205
rect -543 204 -509 205
rect 130 201 154 206
rect -2549 163 -2499 174
rect -2477 163 -2427 174
rect -509 163 -459 174
rect -437 163 -387 174
rect -49 165 -22 172
<< nwell >>
rect -2616 744 -2418 745
rect -320 744 -173 745
rect 65 727 193 745
rect -2616 677 -2609 695
rect -2616 190 -2608 208
rect 65 140 193 159
<< locali >>
rect -1767 480 -1747 488
rect -1767 463 -1766 480
rect -1749 463 -1747 480
rect -1767 411 -1747 463
rect -1767 394 -1765 411
rect -1748 394 -1747 411
rect -1767 387 -1747 394
rect -1192 480 -1163 488
rect -1192 463 -1187 480
rect -1170 463 -1163 480
rect -1192 411 -1163 463
rect -1192 394 -1187 411
rect -1170 394 -1163 411
rect -1192 387 -1163 394
<< viali >>
rect -1766 463 -1749 480
rect -1765 394 -1748 411
rect -1187 463 -1170 480
rect -1187 394 -1170 411
<< metal1 >>
rect -2592 740 -2564 745
rect -2592 739 -2560 740
rect -2539 739 -2520 745
rect -2592 713 -2589 739
rect -2563 713 -2560 739
rect -1891 736 -1868 744
rect -1769 736 -1746 744
rect -1540 729 -1396 745
rect -1190 736 -1167 745
rect -1068 737 -1045 745
rect -416 737 -397 745
rect -372 740 -344 745
rect -372 738 -340 740
rect -2592 712 -2560 713
rect -372 712 -369 738
rect -343 712 -340 738
rect -3 731 31 745
rect 63 730 91 745
rect -372 710 -340 712
rect -1768 432 -1736 434
rect -1768 394 -1765 432
rect -1739 406 -1736 432
rect -1748 404 -1736 406
rect -1198 426 -1166 429
rect -1748 394 -1744 404
rect -1198 400 -1195 426
rect -1169 400 -1166 426
rect -1198 397 -1187 400
rect -1170 397 -1166 400
rect -1768 393 -1744 394
rect -1746 391 -1744 393
rect -154 187 -121 189
rect -1198 174 -1166 176
rect -1198 148 -1195 174
rect -1169 148 -1166 174
rect -154 161 -151 187
rect -124 161 -121 187
rect -154 160 -121 161
rect -1198 146 -1166 148
rect -155 159 -3 160
rect -155 146 31 159
rect -416 140 -397 145
rect -372 140 -344 145
rect -3 140 31 146
rect 64 140 91 161
<< via1 >>
rect -2589 713 -2563 739
rect -369 712 -343 738
rect -1765 411 -1739 432
rect -1765 406 -1748 411
rect -1748 406 -1739 411
rect -1195 411 -1169 426
rect -1195 400 -1187 411
rect -1187 400 -1170 411
rect -1170 400 -1169 411
rect -1195 148 -1169 174
rect -151 161 -124 187
<< metal2 >>
rect -2592 739 -2560 740
rect -2592 713 -2589 739
rect -2563 728 -2560 739
rect -372 738 -340 740
rect -372 728 -369 738
rect -2563 713 -369 728
rect -2592 712 -369 713
rect -343 712 -340 738
rect -260 718 -229 742
rect -2592 710 -340 712
rect -2616 677 -2609 695
rect -149 655 -127 657
rect -1726 617 -1642 637
rect -154 621 -127 655
rect -1681 570 -667 592
rect -328 571 -293 593
rect -1686 473 -785 495
rect -1768 432 -1736 434
rect -1768 406 -1765 432
rect -1739 429 -1736 432
rect -1739 426 -1166 429
rect -1739 406 -1195 426
rect -1768 404 -1195 406
rect -1198 400 -1195 404
rect -1169 400 -1166 426
rect -1198 397 -1166 400
rect -1681 295 -1115 317
rect -1731 265 -1683 266
rect -1731 241 -1642 265
rect -1137 262 -1115 295
rect -807 312 -785 473
rect -689 450 -667 570
rect -147 564 -127 565
rect -147 531 -125 564
rect -145 530 -125 531
rect -252 451 -220 475
rect 182 474 193 497
rect -692 446 -667 450
rect -692 382 -666 446
rect 182 392 193 414
rect -692 361 -279 382
rect -300 347 -279 361
rect -300 326 -113 347
rect -807 290 -522 312
rect -700 262 -113 267
rect -1137 246 -113 262
rect -1137 240 -661 246
rect -2616 190 -2608 208
rect -154 187 -121 189
rect -1198 175 -1166 176
rect -154 175 -151 187
rect -1198 174 -151 175
rect -1198 148 -1195 174
rect -1169 161 -151 174
rect -124 161 -121 187
rect -1169 159 -121 161
rect -1169 158 -1129 159
rect -1169 148 -1166 158
rect -1198 146 -1166 148
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1627737364
transform 1 0 38 0 1 181
box -172 -22 155 550
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1627737364
transform 1 0 -454 0 -1 305
box 133 -440 320 165
use sky130_hilas_FGBiasWeakGate2x1cell  sky130_hilas_FGBiasWeakGate2x1cell_0
timestamp 1627737364
transform -1 0 -1859 0 1 522
box -396 -382 757 223
use sky130_hilas_FGBias2x1cell  sky130_hilas_FGBias2x1cell_0
timestamp 1627737364
transform 1 0 -1077 0 1 522
box -396 -382 757 223
<< labels >>
rlabel metal2 -1726 617 -1690 636 0 VIN11
port 2 nsew analog default
rlabel metal2 -1731 241 -1695 266 0 VIN12
port 1 nsew analog default
rlabel metal1 -3 739 31 745 0 VGND
port 7 nsew analog default
rlabel metal1 63 739 91 745 0 VPWR
port 6 nsew analog default
rlabel metal1 64 140 91 146 0 VPWR
port 6 nsew power default
rlabel metal1 -3 140 31 146 0 VGND
port 7 nsew ground default
rlabel metal2 -252 451 -220 475 0 VIN21
port 3 nsew analog default
rlabel metal2 -260 718 -229 742 1 VIN22
port 4 n analog default
rlabel metal1 -372 737 -344 745 0 VINJ
port 8 nsew power default
rlabel metal1 -372 140 -344 145 0 VINJ
port 8 nsew power default
rlabel metal2 182 474 193 497 0 OUTPUT1
port 9 nsew analog default
rlabel metal2 182 392 193 414 0 OUTPUT2
port 10 nsew analog default
rlabel metal2 -2616 677 -2609 695 0 DRAIN1
port 11 nsew
rlabel metal2 -2616 190 -2608 208 0 DRAIN2
port 12 nsew
rlabel metal1 -2592 738 -2564 745 0 VINJ
port 8 nsew
rlabel metal1 -2539 739 -2520 745 0 COLSEL2
port 13 nsew
rlabel metal1 -1891 736 -1868 744 0 GATE2
port 14 nsew
rlabel metal1 -1769 736 -1746 744 0 VGND
port 7 nsew
rlabel metal1 -1068 737 -1045 745 0 GATE1
port 15 nsew
rlabel metal1 -1190 737 -1167 745 0 VGND
port 7 nsew
rlabel metal1 -416 737 -397 745 0 COLSEL1
port 16 nsew
rlabel metal1 -416 140 -397 145 0 COLSEL1
port 16 nsew
rlabel metal1 -1498 733 -1438 745 0 VTUN
port 17 nsew
<< end >>
