magic
tech sky130A
timestamp 1628698461
<< metal3 >>
rect -416 -216 -186 12
<< mimcap >>
rect -401 -105 -201 -2
rect -401 -118 -316 -105
rect -302 -118 -201 -105
rect -401 -202 -201 -118
<< mimcapcontact >>
rect -316 -118 -302 -105
<< metal4 >>
rect -331 -93 -286 -92
rect -333 -105 -281 -93
rect -333 -118 -316 -105
rect -302 -118 -281 -105
rect -333 -142 -281 -118
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
