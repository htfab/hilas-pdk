magic
tech sky130A
timestamp 1625668354
use sky130_hilas_RightProtection  sky130_hilas_RightProtection_0
timestamp 1625582648
transform 1 0 22518 0 1 -15744
box -2054 8715 -826 28728
use sky130_hilas_LeftProtection  sky130_hilas_LeftProtection_0
timestamp 1625577583
transform 1 0 -13278 0 1 -15672
box -2065 -8439 -833 28728
use sky130_hilas_TopProtection  sky130_hilas_TopProtection_0
timestamp 1625575869
transform 1 0 -13875 0 1 13286
box -2 -76 34131 1170
use sky130_hilas_TopLevelTextStructure  sky130_hilas_TopLevelTextStructure_0
timestamp 1625668104
transform 1 0 510 0 1 -11
box -538 0 8596 4255
<< end >>
