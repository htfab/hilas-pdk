magic
tech sky130A
timestamp 1637975350
<< error_p >>
rect 1430 1276 1480 1281
rect 1610 1276 1660 1282
rect 766 1267 818 1273
rect 818 1266 846 1267
rect 1120 1266 1170 1271
rect 1724 1246 1725 1263
rect 1430 1234 1480 1239
rect 1610 1234 1660 1240
rect 766 1225 818 1231
rect 1120 1224 1170 1229
rect 1430 1209 1480 1215
rect 1750 1209 1800 1215
rect 692 1200 745 1205
rect 839 1200 891 1205
rect 1049 1199 1099 1205
rect 1191 1199 1241 1205
rect 1430 1167 1480 1173
rect 1750 1167 1800 1173
rect 692 1158 745 1163
rect 839 1158 891 1163
rect 1049 1157 1099 1163
rect 1191 1157 1241 1163
rect 766 1107 818 1113
rect 818 1106 846 1107
rect 1120 1106 1170 1111
rect 1430 1106 1480 1112
rect 1750 1106 1800 1112
rect 766 1065 818 1071
rect 1120 1064 1170 1069
rect 1430 1064 1480 1070
rect 1750 1064 1800 1070
rect 692 1040 745 1045
rect 839 1040 891 1045
rect 1049 1039 1099 1045
rect 1191 1039 1241 1045
rect 1430 1040 1480 1045
rect 1610 1039 1660 1045
rect 1724 1016 1725 1033
rect 692 998 745 1003
rect 839 998 891 1003
rect 1049 997 1099 1003
rect 1191 997 1241 1003
rect 1430 998 1480 1003
rect 1610 997 1660 1003
rect 1430 956 1480 961
rect 1610 956 1660 962
rect 766 947 818 953
rect 818 946 846 947
rect 1120 946 1170 951
rect 1724 926 1725 943
rect 1430 914 1480 919
rect 1610 914 1660 920
rect 766 905 818 911
rect 1120 904 1170 909
rect 1430 889 1480 895
rect 1750 889 1800 895
rect 692 880 745 885
rect 839 880 891 885
rect 1049 879 1099 885
rect 1191 879 1241 885
rect 1430 847 1480 853
rect 1750 847 1800 853
rect 692 838 745 843
rect 839 838 891 843
rect 1049 837 1099 843
rect 1191 837 1241 843
rect 766 787 818 793
rect 818 786 846 787
rect 1120 786 1170 791
rect 1430 786 1480 792
rect 1750 786 1800 792
rect 766 745 818 751
rect 1120 744 1170 749
rect 1430 744 1480 750
rect 1750 744 1800 750
rect 692 720 745 725
rect 839 720 891 725
rect 1049 719 1099 725
rect 1191 719 1241 725
rect 1430 720 1480 725
rect 1610 719 1660 725
rect 1724 696 1725 713
rect 692 678 745 683
rect 839 678 891 683
rect 1049 677 1099 683
rect 1191 677 1241 683
rect 1430 678 1480 683
rect 1610 677 1660 683
rect 3022 659 3023 667
rect 1430 626 1480 631
rect 1610 626 1660 632
rect 766 617 818 623
rect 818 616 846 617
rect 1120 616 1170 621
rect 1724 596 1725 613
rect 1430 584 1480 589
rect 1610 584 1660 590
rect 766 575 818 581
rect 1120 574 1170 579
rect 1430 559 1480 565
rect 1750 559 1800 565
rect 692 550 745 555
rect 839 550 891 555
rect 1049 549 1099 555
rect 1191 549 1241 555
rect 1430 517 1480 523
rect 1750 517 1800 523
rect 692 508 745 513
rect 839 508 891 513
rect 1049 507 1099 513
rect 1191 507 1241 513
rect 766 457 818 463
rect 818 456 846 457
rect 1120 456 1170 461
rect 1430 456 1480 462
rect 1750 456 1800 462
rect 766 415 818 421
rect 1120 414 1170 419
rect 1430 414 1480 420
rect 1750 414 1800 420
rect 692 390 745 395
rect 839 390 891 395
rect 1049 389 1099 395
rect 1191 389 1241 395
rect 1430 390 1480 395
rect 1610 389 1660 395
rect 1724 366 1725 383
rect 692 348 745 353
rect 839 348 891 353
rect 1049 347 1099 353
rect 1191 347 1241 353
rect 1430 348 1480 353
rect 1610 347 1660 353
rect 1430 306 1480 311
rect 1610 306 1660 312
rect 766 297 818 303
rect 818 296 846 297
rect 1120 296 1170 301
rect 1724 276 1725 293
rect 1430 264 1480 269
rect 1610 264 1660 270
rect 766 255 818 261
rect 1120 254 1170 259
rect 1430 239 1480 245
rect 1750 239 1800 245
rect 692 230 745 235
rect 839 230 891 235
rect 1049 229 1099 235
rect 1191 229 1241 235
rect 1430 197 1480 203
rect 1750 197 1800 203
rect 692 188 745 193
rect 839 188 891 193
rect 1049 187 1099 193
rect 1191 187 1241 193
rect 766 137 818 143
rect 818 136 846 137
rect 1120 136 1170 141
rect 1430 136 1480 142
rect 1750 136 1800 142
rect 766 95 818 101
rect 1120 94 1170 99
rect 1430 94 1480 100
rect 1750 94 1800 100
rect 692 70 745 75
rect 839 70 891 75
rect 1049 69 1099 75
rect 1191 69 1241 75
rect 1430 70 1480 75
rect 1610 69 1660 75
rect 1724 46 1725 63
rect 692 28 745 33
rect 839 28 891 33
rect 1049 27 1099 33
rect 1191 27 1241 33
rect 1430 28 1480 33
rect 1610 27 1660 33
<< error_s >>
rect 84 10292 137 10299
rect 263 10291 315 10299
rect 84 10250 137 10257
rect 263 10249 315 10257
rect 84 10141 137 10148
rect 263 10140 315 10148
rect 84 10099 137 10106
rect 263 10098 315 10106
rect 84 9990 137 9997
rect 263 9989 315 9997
rect 84 9948 137 9955
rect 263 9947 315 9955
rect 84 9642 137 9649
rect 263 9641 315 9649
rect 84 9600 137 9607
rect 263 9599 315 9607
rect 84 9491 137 9498
rect 263 9490 315 9498
rect 84 9449 137 9456
rect 263 9448 315 9456
rect -688 9375 -636 9381
rect -636 9374 -608 9375
rect -334 9374 -284 9379
rect 84 9340 137 9347
rect 263 9339 315 9347
rect -688 9333 -636 9339
rect -334 9332 -284 9337
rect -762 9308 -709 9313
rect -615 9308 -563 9313
rect -405 9307 -355 9313
rect -263 9307 -213 9313
rect -1370 9300 -1317 9307
rect -1191 9299 -1139 9307
rect 84 9298 137 9305
rect 263 9297 315 9305
rect -762 9266 -709 9271
rect -615 9266 -563 9271
rect -405 9265 -355 9271
rect -263 9265 -213 9271
rect -1370 9258 -1317 9265
rect -1191 9257 -1139 9265
rect -688 9215 -636 9221
rect -636 9214 -608 9215
rect -334 9214 -284 9219
rect -688 9173 -636 9179
rect -334 9172 -284 9177
rect -1370 9149 -1317 9156
rect -1191 9148 -1139 9156
rect -762 9148 -709 9153
rect -615 9148 -563 9153
rect -405 9147 -355 9153
rect -263 9147 -213 9153
rect -1370 9107 -1317 9114
rect -1191 9106 -1139 9114
rect -762 9106 -709 9111
rect -615 9106 -563 9111
rect -405 9105 -355 9111
rect -263 9105 -213 9111
rect -688 9055 -636 9061
rect -636 9054 -608 9055
rect -334 9054 -284 9059
rect -688 9013 -636 9019
rect -334 9012 -284 9017
rect -1370 8998 -1317 9005
rect -1191 8997 -1139 9005
rect -762 8988 -709 8993
rect -615 8988 -563 8993
rect -405 8987 -355 8993
rect -263 8987 -213 8993
rect 84 8992 137 8999
rect 263 8991 315 8999
rect -1370 8956 -1317 8963
rect -1191 8955 -1139 8963
rect -762 8946 -709 8951
rect -615 8946 -563 8951
rect -405 8945 -355 8951
rect -263 8945 -213 8951
rect 84 8950 137 8957
rect 263 8949 315 8957
rect -688 8895 -636 8901
rect -636 8894 -608 8895
rect -334 8894 -284 8899
rect -688 8853 -636 8859
rect -334 8852 -284 8857
rect 84 8841 137 8848
rect 263 8840 315 8848
rect -762 8828 -709 8833
rect -615 8828 -563 8833
rect -405 8827 -355 8833
rect -263 8827 -213 8833
rect 84 8799 137 8806
rect 263 8798 315 8806
rect -762 8786 -709 8791
rect -615 8786 -563 8791
rect -405 8785 -355 8791
rect -263 8785 -213 8791
rect 84 8690 137 8697
rect 263 8689 315 8697
rect 84 8648 137 8655
rect 263 8647 315 8655
rect 84 8342 137 8349
rect 263 8341 315 8349
rect 84 8300 137 8307
rect 263 8299 315 8307
rect 84 8191 137 8198
rect 263 8190 315 8198
rect 84 8149 137 8156
rect 263 8148 315 8156
rect 84 8040 137 8047
rect 263 8039 315 8047
rect 84 7998 137 8005
rect 263 7997 315 8005
rect 84 7692 137 7699
rect 263 7691 315 7699
rect 84 7650 137 7657
rect 263 7649 315 7657
rect 84 7541 137 7548
rect 263 7540 315 7548
rect 84 7499 137 7506
rect 263 7498 315 7506
rect 84 7390 137 7397
rect 263 7389 315 7397
rect 84 7348 137 7355
rect 263 7347 315 7355
rect 84 7042 137 7049
rect 263 7041 315 7049
rect 84 7000 137 7007
rect 263 6999 315 7007
rect 84 6891 137 6898
rect 263 6890 315 6898
rect 84 6849 137 6856
rect 263 6848 315 6856
rect -688 6775 -636 6781
rect -636 6774 -608 6775
rect -334 6774 -284 6779
rect 84 6740 137 6747
rect 263 6739 315 6747
rect -688 6733 -636 6739
rect -334 6732 -284 6737
rect -762 6708 -709 6713
rect -615 6708 -563 6713
rect -405 6707 -355 6713
rect -263 6707 -213 6713
rect -1370 6700 -1317 6707
rect -1191 6699 -1139 6707
rect 84 6698 137 6705
rect 263 6697 315 6705
rect -762 6666 -709 6671
rect -615 6666 -563 6671
rect -405 6665 -355 6671
rect -263 6665 -213 6671
rect -1370 6658 -1317 6665
rect -1191 6657 -1139 6665
rect -688 6615 -636 6621
rect -636 6614 -608 6615
rect -334 6614 -284 6619
rect -688 6573 -636 6579
rect -334 6572 -284 6577
rect -1370 6549 -1317 6556
rect -1191 6548 -1139 6556
rect -762 6548 -709 6553
rect -615 6548 -563 6553
rect -405 6547 -355 6553
rect -263 6547 -213 6553
rect -1370 6507 -1317 6514
rect -1191 6506 -1139 6514
rect -762 6506 -709 6511
rect -615 6506 -563 6511
rect -405 6505 -355 6511
rect -263 6505 -213 6511
rect -688 6455 -636 6461
rect -636 6454 -608 6455
rect -334 6454 -284 6459
rect -688 6413 -636 6419
rect -334 6412 -284 6417
rect -1370 6398 -1317 6405
rect -1191 6397 -1139 6405
rect -762 6388 -709 6393
rect -615 6388 -563 6393
rect -405 6387 -355 6393
rect -263 6387 -213 6393
rect 84 6392 137 6399
rect 263 6391 315 6399
rect -1370 6356 -1317 6363
rect -1191 6355 -1139 6363
rect -762 6346 -709 6351
rect -615 6346 -563 6351
rect -405 6345 -355 6351
rect -263 6345 -213 6351
rect 84 6350 137 6357
rect 263 6349 315 6357
rect -688 6295 -636 6301
rect -636 6294 -608 6295
rect -334 6294 -284 6299
rect -688 6253 -636 6259
rect -334 6252 -284 6257
rect 84 6241 137 6248
rect 263 6240 315 6248
rect -762 6228 -709 6233
rect -615 6228 -563 6233
rect -405 6227 -355 6233
rect -263 6227 -213 6233
rect 84 6199 137 6206
rect 263 6198 315 6206
rect -762 6186 -709 6191
rect -615 6186 -563 6191
rect -405 6185 -355 6191
rect -263 6185 -213 6191
rect 84 6090 137 6097
rect 263 6089 315 6097
rect 84 6048 137 6055
rect 263 6047 315 6055
rect 84 5742 137 5749
rect 263 5741 315 5749
rect 84 5700 137 5707
rect 263 5699 315 5707
rect 84 5591 137 5598
rect 263 5590 315 5598
rect 84 5549 137 5556
rect 263 5548 315 5556
rect -2273 5501 -2221 5507
rect -2221 5500 -2193 5501
rect -1919 5500 -1869 5505
rect -2273 5459 -2221 5465
rect -1919 5458 -1869 5463
rect 84 5440 137 5447
rect 263 5439 315 5447
rect -2347 5434 -2294 5439
rect -2200 5434 -2148 5439
rect -1990 5433 -1940 5439
rect -1848 5433 -1798 5439
rect -2955 5426 -2902 5433
rect -2776 5425 -2724 5433
rect 84 5398 137 5405
rect 263 5397 315 5405
rect -2347 5392 -2294 5397
rect -2200 5392 -2148 5397
rect -1990 5391 -1940 5397
rect -1848 5391 -1798 5397
rect -2955 5384 -2902 5391
rect -2776 5383 -2724 5391
rect -2273 5341 -2221 5347
rect -2221 5340 -2193 5341
rect -1919 5340 -1869 5345
rect -2273 5299 -2221 5305
rect -1919 5298 -1869 5303
rect -2955 5275 -2902 5282
rect -2776 5274 -2724 5282
rect -2347 5274 -2294 5279
rect -2200 5274 -2148 5279
rect -1990 5273 -1940 5279
rect -1848 5273 -1798 5279
rect -2955 5233 -2902 5240
rect -2776 5232 -2724 5240
rect -2347 5232 -2294 5237
rect -2200 5232 -2148 5237
rect -1990 5231 -1940 5237
rect -1848 5231 -1798 5237
rect -2273 5181 -2221 5187
rect -2221 5180 -2193 5181
rect -1919 5180 -1869 5185
rect -2273 5139 -2221 5145
rect -1919 5138 -1869 5143
rect -2955 5124 -2902 5131
rect -2776 5123 -2724 5131
rect -2347 5114 -2294 5119
rect -2200 5114 -2148 5119
rect -1990 5113 -1940 5119
rect -1848 5113 -1798 5119
rect 84 5092 137 5099
rect 263 5091 315 5099
rect -2955 5082 -2902 5089
rect -2776 5081 -2724 5089
rect -2347 5072 -2294 5077
rect -2200 5072 -2148 5077
rect -1990 5071 -1940 5077
rect -1848 5071 -1798 5077
rect 84 5050 137 5057
rect 263 5049 315 5057
rect -2273 5021 -2221 5027
rect -2221 5020 -2193 5021
rect -1919 5020 -1869 5025
rect -2273 4979 -2221 4985
rect -1919 4978 -1869 4983
rect -2347 4954 -2294 4959
rect -2200 4954 -2148 4959
rect -1990 4953 -1940 4959
rect -1848 4953 -1798 4959
rect 84 4941 137 4948
rect 263 4940 315 4948
rect -2347 4912 -2294 4917
rect -2200 4912 -2148 4917
rect -1990 4911 -1940 4917
rect -1848 4911 -1798 4917
rect 84 4899 137 4906
rect 263 4898 315 4906
rect 84 4790 137 4797
rect 263 4789 315 4797
rect 84 4748 137 4755
rect 263 4747 315 4755
rect 84 4442 137 4449
rect 263 4441 315 4449
rect 84 4400 137 4407
rect 263 4399 315 4407
rect 84 4291 137 4298
rect 263 4290 315 4298
rect 84 4249 137 4256
rect 263 4248 315 4256
rect -688 4175 -636 4181
rect -636 4174 -608 4175
rect -334 4174 -284 4179
rect 84 4140 137 4147
rect 263 4139 315 4147
rect -688 4133 -636 4139
rect -334 4132 -284 4137
rect -762 4108 -709 4113
rect -615 4108 -563 4113
rect -405 4107 -355 4113
rect -263 4107 -213 4113
rect -1370 4100 -1317 4107
rect -1191 4099 -1139 4107
rect 84 4098 137 4105
rect 263 4097 315 4105
rect -762 4066 -709 4071
rect -615 4066 -563 4071
rect -405 4065 -355 4071
rect -263 4065 -213 4071
rect -1370 4058 -1317 4065
rect -1191 4057 -1139 4065
rect -688 4015 -636 4021
rect -636 4014 -608 4015
rect -334 4014 -284 4019
rect -688 3973 -636 3979
rect -334 3972 -284 3977
rect -1370 3949 -1317 3956
rect -1191 3948 -1139 3956
rect -762 3948 -709 3953
rect -615 3948 -563 3953
rect -405 3947 -355 3953
rect -263 3947 -213 3953
rect -1370 3907 -1317 3914
rect -1191 3906 -1139 3914
rect -762 3906 -709 3911
rect -615 3906 -563 3911
rect -405 3905 -355 3911
rect -263 3905 -213 3911
rect -688 3855 -636 3861
rect -636 3854 -608 3855
rect -334 3854 -284 3859
rect -688 3813 -636 3819
rect -334 3812 -284 3817
rect -1370 3798 -1317 3805
rect -1191 3797 -1139 3805
rect -762 3788 -709 3793
rect -615 3788 -563 3793
rect -405 3787 -355 3793
rect -263 3787 -213 3793
rect 84 3792 137 3799
rect 263 3791 315 3799
rect -1370 3756 -1317 3763
rect -1191 3755 -1139 3763
rect -762 3746 -709 3751
rect -615 3746 -563 3751
rect -405 3745 -355 3751
rect -263 3745 -213 3751
rect 84 3750 137 3757
rect 263 3749 315 3757
rect -688 3695 -636 3701
rect -636 3694 -608 3695
rect -334 3694 -284 3699
rect -688 3653 -636 3659
rect -334 3652 -284 3657
rect 84 3641 137 3648
rect 263 3640 315 3648
rect -762 3628 -709 3633
rect -615 3628 -563 3633
rect -405 3627 -355 3633
rect -263 3627 -213 3633
rect 84 3599 137 3606
rect 263 3598 315 3606
rect -762 3586 -709 3591
rect -615 3586 -563 3591
rect -405 3585 -355 3591
rect -263 3585 -213 3591
rect 84 3490 137 3497
rect 263 3489 315 3497
rect 84 3448 137 3455
rect 263 3447 315 3455
rect 84 3142 137 3149
rect 263 3141 315 3149
rect 84 3100 137 3107
rect 263 3099 315 3107
rect 84 2991 137 2998
rect 263 2990 315 2998
rect 84 2949 137 2956
rect 263 2948 315 2956
rect 84 2840 137 2847
rect 263 2839 315 2847
rect 84 2798 137 2805
rect 263 2797 315 2805
rect 84 2492 137 2499
rect 263 2491 315 2499
rect 84 2450 137 2457
rect 263 2449 315 2457
rect 84 2341 137 2348
rect 263 2340 315 2348
rect 84 2299 137 2306
rect 263 2298 315 2306
rect 84 2190 137 2197
rect 263 2189 315 2197
rect 84 2148 137 2155
rect 263 2147 315 2155
rect 84 1842 137 1849
rect 263 1841 315 1849
rect 84 1800 137 1807
rect 263 1799 315 1807
rect 84 1691 137 1698
rect 263 1690 315 1698
rect 84 1649 137 1656
rect 263 1648 315 1656
rect -688 1575 -636 1581
rect -636 1574 -608 1575
rect -334 1574 -284 1579
rect 84 1540 137 1547
rect 263 1539 315 1547
rect -688 1533 -636 1539
rect -334 1532 -284 1537
rect -762 1508 -709 1513
rect -615 1508 -563 1513
rect -405 1507 -355 1513
rect -263 1507 -213 1513
rect -1370 1500 -1317 1507
rect -1191 1499 -1139 1507
rect 84 1498 137 1505
rect 263 1497 315 1505
rect -762 1466 -709 1471
rect -615 1466 -563 1471
rect -405 1465 -355 1471
rect -263 1465 -213 1471
rect -1370 1458 -1317 1465
rect -1191 1457 -1139 1465
rect -688 1415 -636 1421
rect -636 1414 -608 1415
rect -334 1414 -284 1419
rect -688 1373 -636 1379
rect -334 1372 -284 1377
rect -1370 1349 -1317 1356
rect -1191 1348 -1139 1356
rect -762 1348 -709 1353
rect -615 1348 -563 1353
rect -405 1347 -355 1353
rect -263 1347 -213 1353
rect -1370 1307 -1317 1314
rect -1191 1306 -1139 1314
rect -762 1306 -709 1311
rect -615 1306 -563 1311
rect -405 1305 -355 1311
rect -263 1305 -213 1311
rect -688 1255 -636 1261
rect -636 1254 -608 1255
rect -334 1254 -284 1259
rect -688 1213 -636 1219
rect -334 1212 -284 1217
rect -1370 1198 -1317 1205
rect -1191 1197 -1139 1205
rect -762 1188 -709 1193
rect -615 1188 -563 1193
rect -405 1187 -355 1193
rect -263 1187 -213 1193
rect 84 1192 137 1199
rect 263 1191 315 1199
rect -1370 1156 -1317 1163
rect -1191 1155 -1139 1163
rect -762 1146 -709 1151
rect -615 1146 -563 1151
rect -405 1145 -355 1151
rect -263 1145 -213 1151
rect 84 1150 137 1157
rect 263 1149 315 1157
rect -688 1095 -636 1101
rect -636 1094 -608 1095
rect -334 1094 -284 1099
rect -688 1053 -636 1059
rect -334 1052 -284 1057
rect 84 1041 137 1048
rect 263 1040 315 1048
rect -762 1028 -709 1033
rect -615 1028 -563 1033
rect -405 1027 -355 1033
rect -263 1027 -213 1033
rect 84 999 137 1006
rect 263 998 315 1006
rect -762 986 -709 991
rect -615 986 -563 991
rect -405 985 -355 991
rect -263 985 -213 991
rect 84 890 137 897
rect 263 889 315 897
rect 84 848 137 855
rect 263 847 315 855
rect 84 542 137 549
rect 263 541 315 549
rect 84 500 137 507
rect 263 499 315 507
rect 84 391 137 398
rect 263 390 315 398
rect 84 349 137 356
rect 263 348 315 356
rect 84 240 137 247
rect 263 239 315 247
rect 84 198 137 205
rect 263 197 315 205
<< metal1 >>
rect -1629 9056 -1594 9059
rect -1629 9030 -1625 9056
rect -1599 9030 -1594 9056
rect -1629 9027 -1594 9030
rect -1623 5423 -1600 9027
rect -1574 6459 -1551 6466
rect -1574 6457 -1548 6459
rect -1576 6456 -1547 6457
rect -1576 6430 -1574 6456
rect -1548 6430 -1547 6456
rect -1576 6429 -1547 6430
rect -1627 5421 -1600 5423
rect -1628 5420 -1600 5421
rect -1628 5394 -1627 5420
rect -1601 5394 -1600 5420
rect -1628 5393 -1600 5394
rect -1574 6427 -1548 6429
rect -1627 5391 -1601 5393
rect -1574 5263 -1551 6427
rect -1575 5261 -1549 5263
rect -1576 5260 -1548 5261
rect -1576 5234 -1575 5260
rect -1549 5234 -1548 5260
rect -1576 5233 -1548 5234
rect -1575 5231 -1549 5233
rect -1576 5104 -1550 5106
rect -1577 5103 -1549 5104
rect -1577 5077 -1576 5103
rect -1550 5077 -1549 5103
rect -1577 5076 -1549 5077
rect -1576 5074 -1550 5076
rect -1630 4940 -1604 4942
rect -1631 4939 -1601 4940
rect -2978 4853 -2956 4914
rect -1631 4913 -1630 4939
rect -1604 4938 -1601 4939
rect -1604 4913 -1600 4938
rect -1631 4912 -1600 4913
rect -1630 4910 -1600 4912
rect -2980 4851 -2954 4853
rect -2981 4850 -2953 4851
rect -2981 4824 -2980 4850
rect -2954 4824 -2953 4850
rect -2981 4823 -2953 4824
rect -2980 4821 -2954 4823
rect -2721 4763 -2698 4910
rect -2735 4762 -2698 4763
rect -2737 4736 -2734 4762
rect -2708 4737 -2698 4762
rect -2708 4736 -2705 4737
rect -2735 4735 -2707 4736
rect -1623 1259 -1600 4910
rect -1574 3859 -1551 5074
rect -787 4854 -761 4856
rect -788 4853 -760 4854
rect -788 4827 -787 4853
rect -761 4827 -760 4853
rect -788 4826 -760 4827
rect -787 4824 -761 4826
rect -291 4766 -264 4768
rect -292 4765 -263 4766
rect -292 4738 -291 4765
rect -264 4738 -263 4765
rect -292 4737 -263 4738
rect -291 4735 -264 4737
rect -1574 3857 -1548 3859
rect -1575 3856 -1547 3857
rect -1575 3830 -1574 3856
rect -1548 3830 -1547 3856
rect -1575 3829 -1547 3830
rect -1574 3827 -1548 3829
rect -1624 1257 -1598 1259
rect -1625 1256 -1597 1257
rect -1625 1230 -1624 1256
rect -1598 1230 -1597 1256
rect -1625 1229 -1597 1230
rect -1624 1227 -1598 1229
<< via1 >>
rect -1625 9030 -1599 9056
rect -1574 6430 -1548 6456
rect -1627 5394 -1601 5420
rect -1575 5234 -1549 5260
rect -1576 5077 -1550 5103
rect -1630 4913 -1604 4939
rect -2980 4824 -2954 4850
rect -2734 4736 -2708 4762
rect -787 4827 -761 4853
rect -291 4738 -264 4765
rect -1574 3830 -1548 3856
rect -1624 1230 -1598 1256
<< metal2 >>
rect -1628 9056 -1596 9058
rect -1628 9030 -1625 9056
rect -1599 9052 -1596 9056
rect -1599 9034 -1522 9052
rect -1599 9030 -1596 9034
rect -1628 9028 -1596 9030
rect -1578 6456 -1545 6458
rect -1578 6430 -1574 6456
rect -1548 6452 -1545 6456
rect -1548 6434 -1522 6452
rect -1548 6430 -1545 6434
rect -1578 6428 -1545 6430
rect -1629 5420 -1599 5422
rect -1630 5414 -1627 5420
rect -1722 5400 -1627 5414
rect -1630 5394 -1627 5400
rect -1601 5394 -1598 5420
rect -1629 5392 -1599 5394
rect -1577 5260 -1547 5262
rect -1578 5254 -1575 5260
rect -1722 5240 -1575 5254
rect -1578 5234 -1575 5240
rect -1549 5234 -1546 5260
rect -1577 5232 -1547 5234
rect -1579 5103 -1547 5105
rect -1579 5097 -1576 5103
rect -1722 5083 -1576 5097
rect -1579 5077 -1576 5083
rect -1550 5077 -1547 5103
rect -1579 5075 -1547 5077
rect -1633 4939 -1601 4941
rect -1633 4933 -1630 4939
rect -1722 4919 -1630 4933
rect -1633 4913 -1630 4919
rect -1604 4913 -1601 4939
rect -1633 4911 -1601 4913
rect -789 4853 -759 4855
rect -2980 4852 -787 4853
rect -2982 4850 -787 4852
rect -2983 4824 -2980 4850
rect -2954 4827 -787 4850
rect -761 4827 -758 4853
rect -2954 4824 -2951 4827
rect -789 4825 -759 4827
rect -2982 4822 -2952 4824
rect -293 4765 -263 4766
rect -2734 4764 -2708 4765
rect -294 4764 -291 4765
rect -2736 4762 -291 4764
rect -2736 4736 -2734 4762
rect -2708 4738 -291 4762
rect -264 4738 -261 4765
rect -2708 4736 -2707 4738
rect -293 4736 -263 4738
rect -2736 4734 -2707 4736
rect -2734 4733 -2708 4734
rect -1576 3856 -1546 3858
rect -1577 3830 -1574 3856
rect -1548 3852 -1545 3856
rect -1548 3834 -1522 3852
rect -1548 3830 -1545 3834
rect -1576 3828 -1546 3830
rect -1626 1256 -1596 1258
rect -1627 1230 -1624 1256
rect -1598 1252 -1595 1256
rect -1598 1234 -1522 1252
rect -1598 1230 -1595 1234
rect -1626 1228 -1596 1230
use sky130_hilas_VinjDecode2to4_Spaced01  sky130_hilas_VinjDecode2to4_Spaced01_0
array 1 1 1548 1 4 2600
timestamp 1637974713
transform 1 0 -1454 0 1 958
box -86 -963 1462 1642
use sky130_hilas_CellVoltageDAC01  sky130_hilas_CellVoltageDAC01_0
array 1 1 3111 1 16 650
timestamp 1637956455
transform 1 0 18 0 1 14
box -92 -14 3093 645
use sky130_hilas_VinjDecode2to4  sky130_hilas_VinjDecode2to4_1
timestamp 1637953024
transform 1 0 -2402 0 1 4853
box -637 31 694 681
<< end >>
