magic
tech sky130A
timestamp 1607954820
<< metal1 >>
rect 38 460 58 464
rect 621 460 640 464
rect 38 -141 58 -137
rect 621 -141 640 -137
<< metal2 >>
rect -36 433 -31 453
rect -36 385 -31 405
rect -36 335 -30 355
rect 665 335 672 355
rect -36 270 -30 290
rect 666 270 672 290
rect -36 220 -31 240
rect -36 172 -31 192
rect -36 131 -31 151
rect -36 83 -31 103
rect -36 33 -30 53
rect 666 33 672 53
rect -36 -32 -30 -12
rect 666 -32 672 -12
rect -36 -82 -31 -62
rect -36 -130 -31 -110
use sky130_hilas_TgateDouble01  sky130_hilas_TgateDouble01_1
timestamp 1607953977
transform 1 0 227 0 1 40
box -263 -181 445 -29
use sky130_hilas_TgateDouble01  sky130_hilas_TgateDouble01_0
timestamp 1607953977
transform 1 0 227 0 -1 283
box -263 -181 445 -29
use sky130_hilas_TgateDouble01  sky130_hilas_TgateDouble01_3
timestamp 1607953977
transform 1 0 227 0 1 342
box -263 -181 445 -29
use sky130_hilas_TgateDouble01  sky130_hilas_TgateDouble01_2
timestamp 1607953977
transform 1 0 227 0 -1 -19
box -263 -181 445 -29
<< labels >>
rlabel metal1 621 460 640 464 0 Vdd
rlabel metal1 38 460 58 464 0 GND
rlabel metal2 665 335 672 355 0 Output1
rlabel metal2 666 33 672 53 0 Output3
rlabel metal2 666 270 672 290 0 Output2
rlabel metal2 666 -32 672 -12 0 Output4
rlabel metal2 -36 335 -30 355 0 Select1
rlabel metal2 -36 270 -30 290 0 Select2
rlabel metal2 -36 33 -30 53 0 Select3
rlabel metal2 -36 -32 -30 -12 0 Select4
rlabel metal1 621 -141 640 -137 0 GND
rlabel metal1 38 -141 58 -137 0 Vdd
rlabel metal2 -36 433 -31 453 0 Input1_1
rlabel metal2 -36 385 -31 405 0 Input2_1
rlabel metal2 -36 172 -31 192 0 Input1_2
rlabel metal2 -36 220 -31 240 0 Input2_2
rlabel metal2 -36 131 -31 151 0 Input1_3
rlabel metal2 -36 83 -31 103 0 Input2_3
rlabel metal2 -36 -82 -31 -62 0 Input2_4
rlabel metal2 -36 -130 -31 -110 0 Input1_4
<< end >>
