VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_horizpcell01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_horizpcell01 ;
  ORIGIN 2.890 -0.470 ;
  SIZE 2.560 BY 1.850 ;
  OBS
      LAYER nwell ;
        RECT -2.890 0.480 -0.330 2.320 ;
        RECT -2.890 0.470 -0.340 0.480 ;
      LAYER li1 ;
        RECT -2.550 1.500 -2.210 1.670 ;
        RECT -1.660 1.170 -1.460 1.740 ;
        RECT -0.940 1.180 -0.720 1.770 ;
        RECT -0.930 1.150 -0.720 1.180 ;
        RECT -2.550 0.880 -2.210 1.050 ;
        RECT -0.930 0.800 -0.730 1.150 ;
      LAYER mcon ;
        RECT -1.650 1.210 -1.480 1.380 ;
        RECT -0.920 1.180 -0.750 1.350 ;
      LAYER met1 ;
        RECT -1.660 1.630 -1.500 2.320 ;
        RECT -1.660 1.410 -1.460 1.630 ;
        RECT -1.260 1.580 -1.100 2.320 ;
        RECT -0.850 1.810 -0.690 2.320 ;
        RECT -0.850 1.720 -0.680 1.810 ;
        RECT -1.270 1.460 -1.100 1.580 ;
        RECT -1.680 1.170 -1.450 1.410 ;
        RECT -1.660 1.150 -1.460 1.170 ;
        RECT -1.660 0.470 -1.500 1.150 ;
        RECT -1.290 0.470 -1.100 1.460 ;
        RECT -0.960 1.670 -0.680 1.720 ;
        RECT -0.960 1.120 -0.690 1.670 ;
        RECT -0.850 0.470 -0.690 1.120 ;
      LAYER met2 ;
        RECT -2.890 1.400 -2.800 1.580 ;
        RECT -2.500 1.400 -0.330 1.580 ;
        RECT -2.510 0.970 -0.330 1.150 ;
  END
END sky130_hilas_horizpcell01
END LIBRARY

