magic
tech sky130A
timestamp 1627737364
<< poly >>
rect -9 17 24 25
rect -9 0 -1 17
rect 16 0 24 17
rect -9 -8 24 0
<< polycont >>
rect -1 0 16 17
<< locali >>
rect -3 17 18 25
rect -3 0 -1 17
rect 16 0 18 17
rect -3 -3 18 0
rect -3 -18 -1 -3
rect 16 -18 18 -3
<< viali >>
rect -1 -20 16 -3
<< metal1 >>
rect -8 26 24 29
rect -8 0 -5 26
rect 21 0 24 26
rect -8 -3 24 0
rect -4 -20 -1 -3
rect 16 -20 19 -3
rect -4 -26 19 -20
<< via1 >>
rect -5 0 21 26
<< metal2 >>
rect -8 26 24 29
rect -8 0 -5 26
rect 21 0 24 26
rect -8 -3 24 0
<< end >>
