magic
tech sky130A
timestamp 1627742263
<< error_s >>
rect 165 440 205 451
rect 315 440 355 451
rect 165 398 205 409
rect 315 398 355 409
rect 89 379 129 389
rect 315 377 355 389
rect 89 337 129 347
rect 315 335 355 347
rect 89 278 129 288
rect 315 278 355 290
rect 89 236 129 246
rect 315 236 355 248
rect 165 216 205 227
rect 315 216 355 227
rect 165 174 205 185
rect 315 174 355 185
rect 165 138 205 149
rect 315 138 355 149
rect 165 96 205 107
rect 315 96 355 107
rect 89 77 129 87
rect 315 75 355 87
rect 89 35 129 45
rect 315 33 355 45
rect 89 -24 129 -14
rect 315 -24 355 -12
rect 89 -66 129 -56
rect 315 -66 355 -54
rect 165 -86 205 -75
rect 315 -86 355 -75
rect 165 -128 205 -117
rect 315 -128 355 -117
<< metal1 >>
rect 38 460 58 464
rect 389 458 408 464
rect 38 -141 58 -137
rect 389 -141 408 -135
<< metal2 >>
rect -36 433 -31 453
rect -36 335 -30 355
rect 433 335 440 355
rect -36 270 -30 290
rect 433 270 440 290
rect -36 172 -31 192
rect -36 131 -31 151
rect -36 33 -30 53
rect 433 33 440 53
rect -36 -32 -30 -12
rect 433 -32 440 -12
rect -36 -130 -31 -110
use sky130_hilas_TgateSingle01  sky130_hilas_TgateSingle01_1
timestamp 1627742263
transform 1 0 227 0 1 40
box -263 -181 213 -29
use sky130_hilas_TgateSingle01  sky130_hilas_TgateSingle01_0
timestamp 1627742263
transform 1 0 227 0 -1 283
box -263 -181 213 -29
use sky130_hilas_TgateSingle01  sky130_hilas_TgateSingle01_3
timestamp 1627742263
transform 1 0 227 0 1 342
box -263 -181 213 -29
use sky130_hilas_TgateSingle01  sky130_hilas_TgateSingle01_2
timestamp 1627742263
transform 1 0 227 0 -1 -19
box -263 -181 213 -29
<< labels >>
rlabel metal2 -36 335 -30 355 0 SELECT1
port 8 nsew analog default
rlabel metal2 -36 270 -30 290 0 SELECT2
port 7 nsew analog default
rlabel metal2 -36 33 -30 53 0 SELECT3
port 4 nsew analog default
rlabel metal2 -36 -32 -30 -12 0 SELECT4
port 3 nsew analog default
rlabel metal1 38 -141 58 -137 0 VPWR
port 2 nsew analog default
rlabel metal2 -36 433 -31 453 0 INPUT1_1
port 9 nsew analog default
rlabel metal2 -36 172 -31 192 0 INPUT1_2
port 6 nsew analog default
rlabel metal2 -36 131 -31 151 0 INPUT1_3
port 5 nsew analog default
rlabel metal2 -36 -130 -31 -110 0 INPUT1_4
port 1 nsew analog default
rlabel metal1 389 458 408 464 0 VGND
port 10 nsew ground default
rlabel metal1 389 -141 408 -135 0 VGND
port 10 nsew ground default
rlabel metal2 433 335 440 355 0 OUTPUT1
port 11 nsew analog default
rlabel metal2 433 270 440 290 0 OUTPUT2
port 12 nsew analog default
rlabel metal2 433 33 440 53 0 OUTPUT3
port 13 nsew analog default
rlabel metal2 433 -32 440 -12 0 OUTPUT4
port 14 nsew analog default
rlabel metal1 38 460 58 464 0 VPWR
port 2 nsew power default
<< end >>
