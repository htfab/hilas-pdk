magic
tech sky130A
timestamp 1637956479
<< error_p >>
rect 1430 1276 1480 1281
rect 1610 1276 1660 1282
rect 766 1267 818 1273
rect 818 1266 846 1267
rect 1120 1266 1170 1271
rect 1724 1246 1725 1263
rect 1430 1234 1480 1239
rect 1610 1234 1660 1240
rect 766 1225 818 1231
rect 1120 1224 1170 1229
rect 1430 1209 1480 1215
rect 1750 1209 1800 1215
rect 692 1200 745 1205
rect 839 1200 891 1205
rect 1049 1199 1099 1205
rect 1191 1199 1241 1205
rect 84 1192 137 1199
rect 263 1191 315 1199
rect 1430 1167 1480 1173
rect 1750 1167 1800 1173
rect 692 1158 745 1163
rect 839 1158 891 1163
rect 1049 1157 1099 1163
rect 1191 1157 1241 1163
rect 84 1150 137 1157
rect 263 1149 315 1157
rect 766 1107 818 1113
rect 818 1106 846 1107
rect 1120 1106 1170 1111
rect 1430 1106 1480 1112
rect 1750 1106 1800 1112
rect 766 1065 818 1071
rect 1120 1064 1170 1069
rect 1430 1064 1480 1070
rect 1750 1064 1800 1070
rect 84 1041 137 1048
rect 263 1040 315 1048
rect 692 1040 745 1045
rect 839 1040 891 1045
rect 1049 1039 1099 1045
rect 1191 1039 1241 1045
rect 1430 1040 1480 1045
rect 1610 1039 1660 1045
rect 1724 1016 1725 1033
rect 84 999 137 1006
rect 263 998 315 1006
rect 692 998 745 1003
rect 839 998 891 1003
rect 1049 997 1099 1003
rect 1191 997 1241 1003
rect 1430 998 1480 1003
rect 1610 997 1660 1003
rect 1430 956 1480 961
rect 1610 956 1660 962
rect 766 947 818 953
rect 818 946 846 947
rect 1120 946 1170 951
rect 1724 926 1725 943
rect 1430 914 1480 919
rect 1610 914 1660 920
rect 766 905 818 911
rect 1120 904 1170 909
rect 84 890 137 897
rect 263 889 315 897
rect 1430 889 1480 895
rect 1750 889 1800 895
rect 692 880 745 885
rect 839 880 891 885
rect 1049 879 1099 885
rect 1191 879 1241 885
rect 84 848 137 855
rect 263 847 315 855
rect 1430 847 1480 853
rect 1750 847 1800 853
rect 692 838 745 843
rect 839 838 891 843
rect 1049 837 1099 843
rect 1191 837 1241 843
rect 766 787 818 793
rect 818 786 846 787
rect 1120 786 1170 791
rect 1430 786 1480 792
rect 1750 786 1800 792
rect 766 745 818 751
rect 1120 744 1170 749
rect 1430 744 1480 750
rect 1750 744 1800 750
rect 692 720 745 725
rect 839 720 891 725
rect 1049 719 1099 725
rect 1191 719 1241 725
rect 1430 720 1480 725
rect 1610 719 1660 725
rect 1724 696 1725 713
rect 692 678 745 683
rect 839 678 891 683
rect 1049 677 1099 683
rect 1191 677 1241 683
rect 1430 678 1480 683
rect 1610 677 1660 683
rect 3022 659 3023 667
rect 1430 626 1480 631
rect 1610 626 1660 632
rect 766 617 818 623
rect 818 616 846 617
rect 1120 616 1170 621
rect 1724 596 1725 613
rect 1430 584 1480 589
rect 1610 584 1660 590
rect 766 575 818 581
rect 1120 574 1170 579
rect 1430 559 1480 565
rect 1750 559 1800 565
rect 692 550 745 555
rect 839 550 891 555
rect 1049 549 1099 555
rect 1191 549 1241 555
rect 84 542 137 549
rect 263 541 315 549
rect 1430 517 1480 523
rect 1750 517 1800 523
rect 692 508 745 513
rect 839 508 891 513
rect 1049 507 1099 513
rect 1191 507 1241 513
rect 84 500 137 507
rect 263 499 315 507
rect 766 457 818 463
rect 818 456 846 457
rect 1120 456 1170 461
rect 1430 456 1480 462
rect 1750 456 1800 462
rect 766 415 818 421
rect 1120 414 1170 419
rect 1430 414 1480 420
rect 1750 414 1800 420
rect 84 391 137 398
rect 263 390 315 398
rect 692 390 745 395
rect 839 390 891 395
rect 1049 389 1099 395
rect 1191 389 1241 395
rect 1430 390 1480 395
rect 1610 389 1660 395
rect 1724 366 1725 383
rect 84 349 137 356
rect 263 348 315 356
rect 692 348 745 353
rect 839 348 891 353
rect 1049 347 1099 353
rect 1191 347 1241 353
rect 1430 348 1480 353
rect 1610 347 1660 353
rect 1430 306 1480 311
rect 1610 306 1660 312
rect 766 297 818 303
rect 818 296 846 297
rect 1120 296 1170 301
rect 1724 276 1725 293
rect 1430 264 1480 269
rect 1610 264 1660 270
rect 766 255 818 261
rect 1120 254 1170 259
rect 84 240 137 247
rect 263 239 315 247
rect 1430 239 1480 245
rect 1750 239 1800 245
rect 692 230 745 235
rect 839 230 891 235
rect 1049 229 1099 235
rect 1191 229 1241 235
rect 84 198 137 205
rect 263 197 315 205
rect 1430 197 1480 203
rect 1750 197 1800 203
rect 692 188 745 193
rect 839 188 891 193
rect 1049 187 1099 193
rect 1191 187 1241 193
rect 766 137 818 143
rect 818 136 846 137
rect 1120 136 1170 141
rect 1430 136 1480 142
rect 1750 136 1800 142
rect 766 95 818 101
rect 1120 94 1170 99
rect 1430 94 1480 100
rect 1750 94 1800 100
rect 692 70 745 75
rect 839 70 891 75
rect 1049 69 1099 75
rect 1191 69 1241 75
rect 1430 70 1480 75
rect 1610 69 1660 75
rect 1724 46 1725 63
rect 692 28 745 33
rect 839 28 891 33
rect 1049 27 1099 33
rect 1191 27 1241 33
rect 1430 28 1480 33
rect 1610 27 1660 33
use sky130_hilas_CellVoltageDAC01  sky130_hilas_CellVoltageDAC01_0
array 1 1 3111 1 16 650
timestamp 1637956455
transform 1 0 18 0 1 14
box -92 -14 3093 645
<< end >>
