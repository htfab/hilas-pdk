magic
tech sky130A
timestamp 1634057736
<< checkpaint >>
rect -543 753 1180 772
rect -556 686 1180 753
rect -584 685 1180 686
rect -607 -608 1180 685
rect -543 -618 1180 -608
<< error_s >>
rect 87 110 486 116
rect 87 68 486 74
rect 87 42 486 48
rect 87 0 486 6
<< psubdiff >>
rect 519 99 562 110
rect 519 82 533 99
rect 550 82 562 99
rect 519 74 562 82
rect 519 33 562 42
rect 519 16 533 33
rect 550 16 562 33
rect 519 6 562 16
<< psubdiffcont >>
rect 533 82 550 99
rect 533 16 550 33
<< poly >>
rect 14 50 487 65
rect 14 41 41 50
<< locali >>
rect 512 103 551 108
rect 512 86 518 103
rect 535 99 551 103
rect 512 82 533 86
rect 550 82 551 99
rect 512 75 551 82
rect 492 33 551 75
rect 492 29 533 33
rect 492 12 518 29
rect 550 16 551 33
rect 535 12 551 16
rect 492 7 551 12
<< viali >>
rect 518 99 535 103
rect 518 86 533 99
rect 533 86 535 99
rect 518 16 533 29
rect 533 16 535 29
rect 518 12 535 16
<< metal1 >>
rect 513 103 540 116
rect 513 86 518 103
rect 535 86 540 103
rect 513 29 540 86
rect 513 12 518 29
rect 535 12 540 29
rect 513 1 540 12
<< metal2 >>
rect 90 80 562 102
rect 0 13 66 34
use sky130_hilas_poly2li  sky130_hilas_poly2li_0
timestamp 1634057707
transform 1 0 23 0 1 22
box 0 0 27 33
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1634057708
transform 1 0 525 0 1 51
box 0 0 23 29
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1634057699
transform 1 0 74 0 1 90
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1634057699
transform 1 0 46 0 1 23
box 0 0 34 33
use sky130_hilas_nFET03_LongL  sky130_hilas_nFET03_LongL_0
timestamp 1634057710
transform 1 0 87 0 1 12
box 0 0 463 62
use sky130_hilas_nFET03_LongL  sky130_hilas_nFET03_LongL_1
timestamp 1634057710
transform 1 0 87 0 1 80
box 0 0 463 62
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
