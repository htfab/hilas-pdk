magic
tech sky130A
timestamp 1632411078
<< error_s >>
rect -350 111 49 117
rect -350 69 49 75
rect -350 43 49 49
rect -350 1 49 7
<< psubdiff >>
rect 82 100 125 111
rect 82 83 96 100
rect 113 83 125 100
rect 82 75 125 83
rect 82 34 125 43
rect 82 17 96 34
rect 113 17 125 34
rect 82 7 125 17
<< psubdiffcont >>
rect 96 83 113 100
rect 96 17 113 34
<< poly >>
rect -423 51 50 66
rect -423 42 -396 51
<< locali >>
rect 75 104 114 109
rect 75 87 81 104
rect 98 100 114 104
rect 75 83 96 87
rect 113 83 114 100
rect 75 76 114 83
rect 55 34 114 76
rect 55 30 96 34
rect 55 13 81 30
rect 113 17 114 34
rect 98 13 114 17
rect 55 8 114 13
<< viali >>
rect 81 100 98 104
rect 81 87 96 100
rect 96 87 98 100
rect 81 17 96 30
rect 96 17 98 30
rect 81 13 98 17
<< metal1 >>
rect 78 104 101 111
rect 78 87 81 104
rect 98 87 101 104
rect 78 30 101 87
rect 78 13 81 30
rect 98 13 101 30
rect 78 7 101 13
<< metal2 >>
rect -437 81 -392 102
rect -437 14 -371 35
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1632409009
transform 1 0 -391 0 1 24
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1632409009
transform 1 0 -381 0 1 91
box -14 -15 20 18
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1629420194
transform 1 0 88 0 1 52
box -10 -8 13 21
use sky130_hilas_nFET03_LongL  sky130_hilas_nFET03_LongL_1
timestamp 1632408239
transform 1 0 -350 0 1 81
box -31 -19 432 43
use sky130_hilas_nFET03_LongL  sky130_hilas_nFET03_LongL_0
timestamp 1632408239
transform 1 0 -350 0 1 13
box -31 -19 432 43
use sky130_hilas_poly2li  sky130_hilas_poly2li_0
timestamp 1629420194
transform 1 0 -414 0 1 23
box -9 -14 18 19
<< end >>
