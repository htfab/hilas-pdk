magic
tech sky130A
timestamp 1627062736
<< psubdiff >>
rect 13 222 53 476
rect 13 205 24 222
rect 41 205 53 222
rect 13 188 53 205
rect 13 171 24 188
rect 41 171 53 188
rect 13 154 53 171
rect 13 137 24 154
rect 41 137 53 154
rect 13 115 53 137
<< psubdiffcont >>
rect 24 205 41 222
rect 24 171 41 188
rect 24 137 41 154
<< poly >>
rect 62 568 364 583
rect 62 305 81 568
rect 62 290 365 305
rect 62 103 82 290
rect 14 93 82 103
rect 14 76 19 93
rect 36 76 53 93
rect 70 76 82 93
rect 14 59 82 76
rect 14 42 20 59
rect 37 42 54 59
rect 71 42 82 59
rect 14 27 82 42
rect 14 25 364 27
rect 14 8 20 25
rect 37 8 54 25
rect 71 10 364 25
rect 71 8 97 10
rect 14 3 97 8
rect 14 0 83 3
<< polycont >>
rect 19 76 36 93
rect 53 76 70 93
rect 20 42 37 59
rect 54 42 71 59
rect 20 8 37 25
rect 54 8 71 25
<< locali >>
rect 95 280 112 318
rect 150 280 167 318
rect 205 280 222 318
rect 260 280 277 318
rect 315 280 332 318
rect 370 280 387 318
rect 19 93 70 101
rect 36 76 53 93
rect 19 75 70 76
rect 19 68 71 75
rect 20 59 71 68
rect 37 42 54 59
rect 20 25 71 42
rect 37 8 54 25
rect 20 0 71 8
<< viali >>
rect 24 222 41 239
rect 24 188 41 205
rect 24 154 41 171
rect 24 120 41 137
<< metal1 >>
rect 18 239 46 245
rect 18 222 24 239
rect 41 222 46 239
rect 18 205 46 222
rect 18 192 24 205
rect 0 188 24 192
rect 41 188 46 205
rect 0 171 46 188
rect 0 160 24 171
rect 18 154 24 160
rect 41 162 46 171
rect 41 154 47 162
rect 18 137 47 154
rect 18 120 24 137
rect 41 120 47 137
rect 18 117 47 120
<< metal2 >>
rect 33 559 339 560
rect 24 526 339 559
rect 24 281 56 526
rect 143 458 437 488
rect 362 454 437 458
rect 399 441 437 454
rect 402 354 437 441
rect 142 321 437 354
rect 24 248 340 281
rect 24 144 56 248
rect 24 112 340 144
rect 0 0 60 82
rect 402 77 437 321
rect 143 45 437 77
rect 143 44 414 45
use sky130_hilas_li2m2  sky130_hilas_li2m2_10
timestamp 1607089160
transform 1 0 210 0 1 126
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_6
timestamp 1607089160
transform 1 0 320 0 1 126
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_15
timestamp 1607089160
transform 1 0 156 0 1 58
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_17
timestamp 1607089160
transform 1 0 265 0 1 58
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_19
timestamp 1607089160
transform 1 0 375 0 1 59
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_9
timestamp 1607089160
transform 1 0 100 0 1 126
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_7
timestamp 1607089160
transform 1 0 44 0 1 15
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_8
timestamp 1607089160
transform 1 0 43 0 1 62
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1607089160
transform 1 0 210 0 1 263
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1607089160
transform 1 0 320 0 1 263
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1607089160
transform 1 0 100 0 1 263
box -14 -15 20 18
use sky130_hilas_nFETLargePart1  sky130_hilas_nFETLargePart1_1
timestamp 1607983547
transform 1 0 255 0 1 53
box -165 -31 137 241
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1607089160
transform 1 0 265 0 1 336
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_4
timestamp 1607089160
transform 1 0 156 0 1 336
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_5
timestamp 1607089160
transform 1 0 375 0 1 336
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_14
timestamp 1607089160
transform 1 0 210 0 1 541
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_18
timestamp 1607089160
transform 1 0 320 0 1 540
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_11
timestamp 1607089160
transform 1 0 101 0 1 541
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_16
timestamp 1607089160
transform 1 0 156 0 1 473
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_12
timestamp 1607089160
transform 1 0 265 0 1 471
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_13
timestamp 1607089160
transform 1 0 376 0 1 470
box -14 -15 20 18
use sky130_hilas_nFETLargePart1  sky130_hilas_nFETLargePart1_0
timestamp 1607983547
transform 1 0 255 0 1 331
box -165 -31 137 241
<< labels >>
rlabel metal2 422 414 436 488 0 DRAIN
port 3 nsew analog default
rlabel metal2 24 485 38 559 0 SOURCE
port 2 nsew analog default
rlabel metal2 0 0 10 82 0 GATE
port 1 nsew analog default
rlabel metal1 0 160 7 192 0 VGND
port 4 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
