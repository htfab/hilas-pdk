magic
tech sky130A
magscale 1 2
timestamp 1632256348
<< error_s >>
rect 714 2034 794 2048
rect 842 1978 862 2012
rect 882 1986 896 2032
rect 920 2010 932 2012
rect 842 1964 856 1978
rect 714 1950 794 1964
rect 1008 1958 1236 1994
rect 766 1912 774 1934
rect 804 1914 814 1924
rect 714 1900 794 1912
rect 652 1852 668 1868
rect 674 1852 682 1870
rect 738 1868 746 1900
rect 766 1896 774 1900
rect 790 1852 800 1862
rect 668 1836 684 1842
rect 806 1836 822 1852
rect 714 1816 794 1828
rect 910 1790 1236 1958
rect 780 1740 1102 1754
rect 24 1656 26 1672
rect 0 1616 28 1656
rect 148 1654 188 1682
rect 646 1666 660 1730
rect 674 1648 688 1740
rect 1376 1732 1414 1760
rect 674 1638 696 1648
rect 680 1624 696 1638
rect 24 1580 26 1616
rect 754 1586 1102 1690
rect 1464 1646 1492 1686
rect 26 1504 192 1580
rect 754 1572 1176 1586
rect 656 1570 1176 1572
rect 0 1420 28 1460
rect 550 1436 1176 1570
rect 550 1428 1200 1436
rect 550 1418 1008 1428
rect 1376 1418 1414 1446
rect 730 1408 742 1418
rect 714 1394 794 1408
rect 730 1390 742 1394
rect 910 1392 964 1408
rect 656 1372 856 1384
rect 656 1338 862 1372
rect 882 1346 896 1392
rect 920 1370 932 1372
rect 656 1324 856 1338
rect 714 1316 794 1324
rect 1008 1318 1236 1402
rect 0 1274 28 1314
rect 662 1294 922 1316
rect 948 1314 1236 1318
rect 938 1294 1236 1314
rect 1376 1306 1414 1334
rect 662 1268 1236 1294
rect 662 1260 924 1268
rect 634 1204 646 1260
rect 656 1228 662 1260
rect 668 1238 680 1260
rect 668 1230 688 1238
rect 668 1228 692 1230
rect 738 1228 746 1260
rect 766 1256 774 1260
rect 854 1246 924 1260
rect 652 1226 692 1228
rect 652 1222 696 1226
rect 652 1214 702 1222
rect 652 1212 714 1214
rect 790 1212 800 1222
rect 634 1196 654 1204
rect 656 1196 662 1212
rect 668 1208 744 1212
rect 668 1202 702 1208
rect 668 1196 684 1202
rect 806 1196 822 1212
rect 634 1192 662 1196
rect 854 1195 922 1246
rect 634 1190 664 1192
rect 794 1191 922 1195
rect 948 1191 1236 1268
rect 794 1190 1236 1191
rect 634 1188 1236 1190
rect 634 1178 680 1188
rect 714 1186 794 1188
rect 908 1186 1236 1188
rect 714 1180 806 1186
rect 634 1168 710 1178
rect 714 1176 794 1180
rect 620 1154 668 1156
rect 646 1144 668 1154
rect 948 1150 1236 1186
rect 592 1120 634 1122
rect 714 1120 730 1144
rect 776 1136 856 1146
rect 0 1078 28 1118
rect 612 1110 634 1120
rect 646 1088 660 1090
rect 580 1078 660 1088
rect 674 1078 688 1116
rect 718 1078 733 1093
rect 776 1078 856 1086
rect 897 1078 912 1093
rect 948 1078 1102 1148
rect 1376 1092 1414 1120
rect 580 1074 1102 1078
rect 526 1052 1102 1074
rect 526 1048 776 1052
rect 596 1046 660 1048
rect 526 1028 660 1046
rect 526 1020 602 1028
rect 0 976 28 1016
rect 608 1010 660 1028
rect 646 1004 660 1010
rect 674 1008 688 1048
rect 726 1042 776 1048
rect 856 1048 1102 1052
rect 1464 1048 1492 1088
rect 856 1042 906 1048
rect 726 1038 906 1042
rect 948 1038 1102 1048
rect 726 1036 1102 1038
rect 714 1032 1102 1036
rect 714 1030 776 1032
rect 718 1016 776 1030
rect 856 1016 1102 1032
rect 674 984 696 1008
rect 718 1001 733 1016
rect 897 1001 912 1016
rect 612 974 634 984
rect 674 978 688 984
rect 592 972 634 974
rect 662 950 922 974
rect 646 940 922 950
rect 948 946 1102 1016
rect 1376 994 1414 1022
rect 1464 1006 1492 1046
rect 620 938 922 940
rect 662 934 922 938
rect 662 930 980 934
rect 550 882 1008 930
rect 1062 906 1142 918
rect 1016 892 1032 898
rect 550 866 1016 882
rect 1214 870 1246 880
rect 0 780 28 820
rect 550 796 1008 866
rect 1062 822 1142 834
rect 550 778 1202 796
rect 1376 778 1414 806
rect 714 770 1202 778
rect 778 762 1202 770
rect 778 744 1236 762
rect 656 700 1236 744
rect 714 686 1236 700
rect 0 634 28 674
rect 702 646 714 676
rect 730 674 742 686
rect 778 676 1236 686
rect 946 674 1236 676
rect 744 660 808 674
rect 938 666 1236 674
rect 1376 666 1414 694
rect 716 632 836 646
rect 910 606 924 646
rect 938 634 966 666
rect 1008 658 1236 666
rect 656 542 946 558
rect 656 522 948 542
rect 0 438 28 478
rect 148 452 188 480
rect 656 428 1102 522
rect 646 364 1102 428
rect 1464 408 1492 448
rect 656 354 1102 364
rect 1376 354 1414 382
rect 910 294 922 304
rect 668 252 684 258
rect 702 252 710 270
rect 714 266 794 278
rect 910 268 980 294
rect 806 242 822 258
rect 652 226 668 242
rect 790 232 800 242
rect 738 194 746 226
rect 776 198 786 208
rect 910 198 922 268
rect 950 266 980 268
rect 1062 266 1142 278
rect 766 194 774 198
rect 714 182 794 194
rect 910 187 924 198
rect 954 187 980 266
rect 1004 242 1008 266
rect 1016 252 1032 258
rect 1000 226 1016 242
rect 1214 230 1246 240
rect 1004 194 1008 226
rect 910 186 980 187
rect 766 160 774 182
rect 714 130 794 144
rect 910 136 924 186
rect 1062 182 1142 194
rect 848 82 862 116
rect 886 108 898 116
rect 882 62 896 108
rect 714 46 794 60
<< nwell >>
rect 24 1504 26 1580
<< metal1 >>
rect 148 1654 188 1662
rect 850 1650 888 1662
rect 148 452 188 460
rect 850 452 888 464
<< metal2 >>
rect 0 1616 10 1656
rect 0 1420 12 1460
rect 938 1420 952 1460
rect 0 1274 12 1314
rect 938 1274 952 1314
rect 0 1078 10 1118
rect 0 976 10 1016
rect 0 780 12 820
rect 938 780 952 820
rect 0 634 12 674
rect 938 634 952 674
rect 0 438 10 478
use sky130_hilas_TgateSingle01  sky130_hilas_TgateSingle01_1
timestamp 1632255311
transform 1 0 526 0 1 778
box 0 0 966 676
use sky130_hilas_TgateSingle01  sky130_hilas_TgateSingle01_2
timestamp 1632255311
transform 1 0 526 0 -1 676
box 0 0 966 676
use sky130_hilas_TgateSingle01  sky130_hilas_TgateSingle01_0
timestamp 1632255311
transform 1 0 526 0 -1 1316
box 0 0 966 676
use sky130_hilas_TgateSingle01  sky130_hilas_TgateSingle01_3
timestamp 1632255311
transform 1 0 526 0 1 1418
box 0 0 966 676
<< labels >>
rlabel metal2 0 1274 12 1314 0 SELECT2
port 7 nsew analog default
rlabel metal1 148 452 188 460 0 VPWR
port 2 nsew analog default
rlabel metal2 0 1078 10 1118 0 INPUT1_2
port 6 nsew analog default
rlabel metal1 850 1650 888 1662 0 VGND
port 10 nsew ground default
rlabel metal1 850 452 888 464 0 VGND
port 10 nsew ground default
rlabel metal2 938 1274 952 1314 0 OUTPUT2
port 12 nsew analog default
rlabel metal1 148 1654 188 1662 0 VPWR
port 2 nsew power default
rlabel metal2 938 634 952 674 0 OUTPUT4
port 14 nsew
rlabel metal2 938 780 952 820 0 OUTPUT3
port 15 nsew
rlabel metal2 938 1420 952 1460 0 OUTPUT1
port 16 nsew
rlabel metal2 0 438 10 478 0 INPUT1_4
port 17 nsew
rlabel metal2 0 634 12 674 0 SELECT4
port 18 nsew
rlabel metal2 0 780 12 820 0 SELECT3
port 19 nsew
rlabel metal2 0 976 10 1016 0 INPUT1_3
port 20 nsew
rlabel metal2 0 1420 12 1460 0 SELECT1
port 21 nsew
rlabel metal2 0 1616 10 1656 0 INPUT1_1
port 22 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
