magic
tech sky130A
timestamp 1627063351
<< error_s >>
rect 100 574 129 592
rect 346 572 375 588
rect 425 572 454 588
rect 504 572 533 588
rect 583 572 612 588
rect 100 542 101 543
rect 128 542 129 543
rect 50 513 68 542
rect 99 541 130 542
rect 100 532 129 541
rect 100 523 110 532
rect 119 523 129 532
rect 100 514 129 523
rect 99 513 130 514
rect 161 513 179 542
rect 346 538 347 539
rect 374 538 375 539
rect 425 538 426 539
rect 453 538 454 539
rect 504 538 505 539
rect 532 538 533 539
rect 583 538 584 539
rect 611 538 612 539
rect 100 512 101 513
rect 128 512 129 513
rect 296 509 314 538
rect 345 537 376 538
rect 424 537 455 538
rect 503 537 534 538
rect 582 537 613 538
rect 346 530 375 537
rect 425 530 454 537
rect 504 530 533 537
rect 583 530 612 537
rect 346 516 356 530
rect 603 516 612 530
rect 346 510 375 516
rect 425 510 454 516
rect 504 510 533 516
rect 583 510 612 516
rect 345 509 376 510
rect 424 509 455 510
rect 503 509 534 510
rect 582 509 613 510
rect 645 509 662 538
rect 679 516 681 517
rect 346 508 347 509
rect 374 508 375 509
rect 425 508 426 509
rect 453 508 454 509
rect 504 508 505 509
rect 532 508 533 509
rect 583 508 584 509
rect 611 508 612 509
rect 100 463 129 481
rect 346 459 375 474
rect 425 459 454 474
rect 504 459 533 474
rect 583 459 612 474
rect 100 422 129 440
rect 346 425 375 441
rect 425 425 454 441
rect 504 425 533 441
rect 583 425 612 441
rect 346 391 347 392
rect 374 391 375 392
rect 425 391 426 392
rect 453 391 454 392
rect 504 391 505 392
rect 532 391 533 392
rect 583 391 584 392
rect 611 391 612 392
rect 100 390 101 391
rect 128 390 129 391
rect 50 361 68 390
rect 99 389 130 390
rect 100 380 129 389
rect 100 371 110 380
rect 119 371 129 380
rect 100 362 129 371
rect 99 361 130 362
rect 161 361 179 390
rect 296 362 314 391
rect 345 390 376 391
rect 424 390 455 391
rect 503 390 534 391
rect 582 390 613 391
rect 346 383 375 390
rect 425 383 454 390
rect 504 383 533 390
rect 583 383 612 390
rect 346 369 356 383
rect 603 369 612 383
rect 346 363 375 369
rect 425 363 454 369
rect 504 363 533 369
rect 583 363 612 369
rect 345 362 376 363
rect 424 362 455 363
rect 503 362 534 363
rect 582 362 613 363
rect 645 362 662 391
rect 674 365 687 369
rect 688 365 701 370
rect 674 362 701 365
rect 346 361 347 362
rect 374 361 375 362
rect 425 361 426 362
rect 453 361 454 362
rect 504 361 505 362
rect 532 361 533 362
rect 583 361 584 362
rect 611 361 612 362
rect 100 360 101 361
rect 128 360 129 361
rect 100 311 129 329
rect 346 312 375 327
rect 425 312 454 327
rect 504 312 533 327
rect 583 312 612 327
rect 100 277 129 295
rect 346 278 375 294
rect 425 278 454 294
rect 504 278 533 294
rect 583 278 612 294
rect 100 245 101 246
rect 128 245 129 246
rect 50 216 68 245
rect 99 244 130 245
rect 100 235 129 244
rect 100 226 110 235
rect 119 226 129 235
rect 100 217 129 226
rect 99 216 130 217
rect 161 216 179 245
rect 346 244 347 245
rect 374 244 375 245
rect 425 244 426 245
rect 453 244 454 245
rect 504 244 505 245
rect 532 244 533 245
rect 583 244 584 245
rect 611 244 612 245
rect 100 215 101 216
rect 128 215 129 216
rect 296 215 314 244
rect 345 243 376 244
rect 424 243 455 244
rect 503 243 534 244
rect 582 243 613 244
rect 346 236 375 243
rect 425 236 454 243
rect 504 236 533 243
rect 583 236 612 243
rect 346 222 356 236
rect 603 222 612 236
rect 346 216 375 222
rect 425 216 454 222
rect 504 216 533 222
rect 583 216 612 222
rect 345 215 376 216
rect 424 215 455 216
rect 503 215 534 216
rect 582 215 613 216
rect 645 215 662 244
rect 346 214 347 215
rect 374 214 375 215
rect 425 214 426 215
rect 453 214 454 215
rect 504 214 505 215
rect 532 214 533 215
rect 583 214 584 215
rect 611 214 612 215
rect 100 166 129 184
rect 346 165 375 180
rect 425 165 454 180
rect 504 165 533 180
rect 583 165 612 180
rect 100 123 129 141
rect 346 131 375 147
rect 425 131 454 147
rect 504 131 533 147
rect 583 131 612 147
rect 346 97 347 98
rect 374 97 375 98
rect 425 97 426 98
rect 453 97 454 98
rect 504 97 505 98
rect 532 97 533 98
rect 583 97 584 98
rect 611 97 612 98
rect 100 91 101 92
rect 128 91 129 92
rect 50 62 68 91
rect 99 90 130 91
rect 100 81 129 90
rect 100 72 110 81
rect 119 72 129 81
rect 100 63 129 72
rect 99 62 130 63
rect 161 62 179 91
rect 296 68 314 97
rect 345 96 376 97
rect 424 96 455 97
rect 503 96 534 97
rect 582 96 613 97
rect 346 89 375 96
rect 425 89 454 96
rect 504 89 533 96
rect 583 89 612 96
rect 346 75 356 89
rect 603 75 612 89
rect 346 69 375 75
rect 425 69 454 75
rect 504 69 533 75
rect 583 69 612 75
rect 345 68 376 69
rect 424 68 455 69
rect 503 68 534 69
rect 582 68 613 69
rect 645 68 662 97
rect 346 67 347 68
rect 374 67 375 68
rect 425 67 426 68
rect 453 67 454 68
rect 504 67 505 68
rect 532 67 533 68
rect 583 67 584 68
rect 611 67 612 68
rect 100 61 101 62
rect 128 61 129 62
rect 100 12 129 30
rect 346 18 375 33
rect 425 18 454 33
rect 504 18 533 33
rect 583 18 612 33
<< nwell >>
rect 823 310 858 311
rect 823 294 840 310
rect 857 294 858 310
<< poly >>
rect 660 529 680 533
rect 172 496 321 520
rect 660 517 679 529
rect 172 387 319 411
rect 660 373 679 390
rect 840 310 858 311
rect 856 294 858 310
rect 172 207 321 231
rect 660 215 679 232
rect 172 87 323 111
rect 660 73 679 90
<< polycont >>
rect 823 294 840 311
<< locali >>
rect 814 294 823 311
<< viali >>
rect 840 294 858 311
<< metal1 >>
rect 101 0 128 605
rect 845 314 858 316
rect 837 311 861 314
rect 837 294 840 311
rect 858 294 861 311
rect 837 291 861 294
rect 847 287 858 291
<< metal2 >>
rect 0 548 688 555
rect 0 537 691 548
rect 0 494 901 512
rect 0 406 688 412
rect 0 394 691 406
rect 0 362 687 369
rect 0 351 691 362
rect 0 236 691 253
rect 0 194 691 211
rect 0 96 691 113
rect 0 52 691 69
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_3
timestamp 1607262215
transform 1 0 112 0 1 55
box -62 -43 67 86
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_2
timestamp 1607262215
transform 1 0 112 0 1 209
box -62 -43 67 86
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_3
timestamp 1607261501
transform 1 0 800 0 1 54
box -521 -54 -121 110
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_2
timestamp 1607261501
transform 1 0 800 0 1 201
box -521 -54 -121 110
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_1
timestamp 1607386385
transform 1 0 968 0 1 -46
box -289 47 -33 232
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_2
timestamp 1607386385
transform 1 0 968 0 -1 351
box -289 47 -33 232
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_1
timestamp 1607262215
transform 1 0 112 0 1 354
box -62 -43 67 86
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_1
timestamp 1607261501
transform 1 0 800 0 1 348
box -521 -54 -121 110
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_0
timestamp 1607386385
transform 1 0 968 0 1 254
box -289 47 -33 232
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_0
timestamp 1607262215
transform 1 0 112 0 1 506
box -62 -43 67 86
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_0
timestamp 1607261501
transform 1 0 800 0 1 495
box -521 -54 -121 110
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_3
timestamp 1607386385
transform 1 0 968 0 -1 652
box -289 47 -33 232
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
