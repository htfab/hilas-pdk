magic
tech sky130A
timestamp 1632256322
<< error_s >>
rect 62 578 101 581
rect 62 536 101 539
rect 62 482 101 485
rect 62 440 101 443
rect 62 386 101 389
rect 62 344 101 347
rect 62 290 101 293
rect 62 248 101 251
rect 0 96 161 212
rect 62 62 101 65
rect 62 20 101 23
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_3
timestamp 1632251308
transform 1 0 0 0 1 480
box 0 0 172 121
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_2
timestamp 1632251308
transform 1 0 0 0 1 384
box 0 0 172 121
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_4
timestamp 1632251308
transform 1 0 0 0 1 288
box 0 0 172 121
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_1
timestamp 1632251308
transform 1 0 0 0 1 192
box 0 0 172 121
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_0
timestamp 1632251308
transform 1 0 0 0 1 96
box 0 0 172 121
use sky130_hilas_pFETdevice01a  sky130_hilas_pFETdevice01a_0
timestamp 1632251417
transform 1 0 0 0 1 0
box 0 0 161 85
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
