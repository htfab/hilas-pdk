magic
tech sky130A
timestamp 1628168646
<< error_s >>
rect 568 195 618 201
rect 640 195 690 201
rect 568 153 618 159
rect 640 153 690 159
rect 568 -318 618 -312
rect 640 -318 690 -312
rect 568 -360 618 -354
rect 640 -360 690 -354
<< nwell >>
rect -337 -242 -281 0
<< psubdiff >>
rect -95 -42 -70 101
rect -95 -59 -92 -42
rect -73 -59 -70 -42
rect -95 -72 -70 -59
rect -95 -75 267 -72
rect -95 -76 146 -75
rect -95 -93 -71 -76
rect -52 -93 -28 -76
rect -9 -93 16 -76
rect 35 -93 56 -76
rect 75 -93 100 -76
rect 119 -92 146 -76
rect 165 -76 267 -75
rect 165 -92 190 -76
rect 119 -93 190 -92
rect 209 -93 236 -76
rect 255 -93 267 -76
rect -95 -97 267 -93
rect -95 -110 -70 -97
rect -95 -127 -92 -110
rect -73 -127 -70 -110
rect -95 -281 -70 -127
<< mvnsubdiff >>
rect -337 -242 -281 0
<< psubdiffcont >>
rect -92 -59 -73 -42
rect -71 -93 -52 -76
rect -28 -93 -9 -76
rect 16 -93 35 -76
rect 56 -93 75 -76
rect 100 -93 119 -76
rect 146 -92 165 -75
rect 190 -93 209 -76
rect 236 -93 255 -76
rect -92 -127 -73 -110
<< poly >>
rect -206 151 293 201
rect -237 134 332 151
rect -237 126 321 134
rect 45 91 64 126
rect 220 90 237 126
rect 46 -293 63 -260
rect 220 -293 237 -260
rect -280 -310 331 -293
rect -202 -367 298 -310
<< locali >>
rect -209 122 297 205
rect -202 114 -154 122
rect -169 89 -154 114
rect -92 -42 -73 -34
rect -92 -75 -73 -59
rect -92 -76 146 -75
rect -92 -93 -71 -76
rect -52 -93 -28 -76
rect -9 -93 16 -76
rect 35 -93 56 -76
rect 75 -93 100 -76
rect 119 -92 146 -76
rect 165 -76 263 -75
rect 165 -92 190 -76
rect 119 -93 190 -92
rect 209 -93 236 -76
rect 255 -93 263 -76
rect -92 -110 -73 -93
rect -92 -135 -73 -127
rect 11 -197 34 -193
rect -172 -279 -170 -254
rect -205 -287 -170 -279
rect -205 -372 300 -287
<< metal1 >>
rect -361 -381 -319 223
rect -113 126 -90 223
rect -113 101 -89 126
rect -113 -382 -90 101
rect 9 -382 32 223
rect 661 217 680 223
rect 661 -382 680 -376
rect 705 -382 733 223
<< metal2 >>
rect -396 155 516 173
rect -217 113 -171 114
rect -396 97 -171 113
rect -396 95 -202 97
rect 554 70 757 71
rect -396 49 757 70
rect -396 48 626 49
rect -396 -49 650 -27
rect 622 -98 648 -63
rect -396 -226 757 -205
rect -396 -227 626 -226
rect -396 -279 -201 -258
rect 510 -315 526 -313
rect -396 -320 526 -315
rect -396 -330 514 -320
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_0
timestamp 1627744303
transform 1 0 986 0 1 62
box -1005 -380 -733 -211
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_2
timestamp 1627744303
transform 1 0 986 0 -1 -231
box -1005 -380 -733 -211
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1628166556
transform 1 0 -103 0 1 -92
box -10 -8 13 21
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_3
timestamp 1628079880
transform 1 0 1056 0 1 433
box -1451 -400 -1278 -210
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_1
timestamp 1628079880
transform 1 0 1056 0 1 19
box -1451 -400 -1278 -210
use sky130_hilas_wellContact  sky130_hilas_wellContact_1
timestamp 1628104465
transform 1 0 1054 0 1 404
box -1448 -441 -1275 -255
use sky130_hilas_wellContact  sky130_hilas_wellContact_0
timestamp 1628104465
transform 1 0 1054 0 1 231
box -1448 -441 -1275 -255
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1628166556
transform 1 0 -191 0 1 -268
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1628166556
transform 1 0 -188 0 1 101
box -14 -15 20 18
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1628164971
transform 1 0 627 0 1 -56
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1628164971
transform 1 0 627 0 1 -116
box -9 -10 23 22
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628166556
transform 1 0 538 0 1 -216
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628166556
transform 1 0 538 0 1 60
box -14 -15 20 18
use sky130_hilas_horizTransCell01  sky130_hilas_horizTransCell01_0
timestamp 1628168286
transform 1 0 790 0 1 -429
box -476 42 -33 359
use sky130_hilas_horizTransCell01  sky130_hilas_horizTransCell01_1
timestamp 1628168286
transform 1 0 790 0 -1 270
box -476 42 -33 359
<< labels >>
rlabel metal1 -361 216 -319 223 0 VTUN
port 9 nsew analog default
rlabel metal1 -113 216 -90 223 0 VGND
port 7 nsew ground default
rlabel metal1 9 215 32 223 0 GATE1
port 8 nsew analog default
rlabel metal1 705 216 733 223 0 VINJ
port 5 nsew power default
rlabel metal2 749 49 757 71 0 ROW1
port 3 nsew analog default
rlabel metal2 750 -226 757 -205 0 ROW2
port 4 nsew analog default
rlabel metal2 -396 155 -389 173 0 DRAIN1
port 1 nsew analog default
rlabel metal2 -396 95 -391 113 0 VIN11
port 2 nsew
rlabel metal1 661 217 680 222 0 COLSEL1
port 6 nsew analog default
rlabel metal1 661 -382 680 -376 0 COLSEL1
port 6 nsew analog default
rlabel metal1 705 -382 733 -375 0 VINJ
port 5 nsew power default
rlabel metal1 -113 -382 -90 -372 0 VGND
port 7 nsew ground default
rlabel metal1 9 -382 32 -374 0 GATE1
port 10 nsew analog default
rlabel metal2 -396 -330 -391 -315 0 DRAIN2
port 11 nsew analog default
rlabel metal2 -396 -279 -390 -258 0 VIN12
port 12 nsew analog default
rlabel metal2 -396 -49 -390 -27 0 COMMONSOURCE
port 13 nsew analog default
<< end >>
