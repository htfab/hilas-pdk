magic
tech sky130A
timestamp 1629137264
<< checkpaint >>
rect -997 2475 436 2508
rect -997 2079 438 2475
rect -997 2046 832 2079
rect -997 2019 834 2046
rect 1014 2019 3928 2079
rect -997 1861 3928 2019
rect -997 644 4178 1861
rect -630 -145 4178 644
rect -630 -204 4006 -145
rect -605 -233 4006 -204
rect 2166 -256 4006 -233
rect 2166 -630 3975 -256
<< error_s >>
rect 568 1021 618 1027
rect 640 1021 690 1027
rect 2608 1021 2658 1027
rect 2680 1021 2730 1027
rect 3068 1025 3095 1031
rect 568 979 618 985
rect 640 979 690 985
rect 2608 979 2658 985
rect 2680 979 2730 985
rect 3068 983 3095 989
rect 3068 958 3095 964
rect 3068 916 3095 922
rect 3068 875 3095 881
rect 3068 833 3095 839
rect 3068 808 3095 814
rect 3068 766 3095 772
rect 3068 725 3095 731
rect 3068 683 3095 689
rect 3068 658 3095 664
rect 3068 616 3095 622
rect 3068 575 3095 581
rect 3068 533 3095 539
rect 568 508 618 514
rect 640 508 690 514
rect 2608 508 2658 514
rect 2680 508 2730 514
rect 3068 508 3095 514
rect 568 466 618 472
rect 640 466 690 472
rect 2608 466 2658 472
rect 2680 466 2730 472
rect 3068 466 3095 472
<< nwell >>
rect 501 1048 699 1049
rect 2797 1048 2944 1049
rect 3182 1031 3310 1049
rect 501 981 508 999
rect 501 494 509 512
rect 3182 444 3310 463
<< locali >>
rect 1350 785 1370 792
rect 1350 768 1351 785
rect 1368 768 1370 785
rect 1350 713 1370 768
rect 1350 696 1352 713
rect 1369 696 1370 713
rect 1350 691 1370 696
rect 1925 785 1954 792
rect 1925 768 1930 785
rect 1947 768 1954 785
rect 1925 713 1954 768
rect 1925 696 1930 713
rect 1947 696 1954 713
rect 1925 691 1954 696
<< viali >>
rect 1351 768 1368 785
rect 1352 696 1369 713
rect 1930 768 1947 785
rect 1930 696 1947 713
<< metal1 >>
rect 525 1044 553 1049
rect 525 1043 557 1044
rect 578 1043 597 1049
rect 525 1017 528 1043
rect 554 1017 557 1043
rect 1226 1040 1249 1048
rect 1348 1040 1371 1048
rect 1577 1033 1721 1049
rect 1927 1040 1950 1049
rect 2049 1041 2072 1049
rect 2701 1041 2720 1049
rect 2745 1044 2773 1049
rect 2745 1042 2777 1044
rect 525 1016 557 1017
rect 2745 1016 2748 1042
rect 2774 1016 2777 1042
rect 3114 1035 3148 1049
rect 3180 1034 3208 1049
rect 2745 1014 2777 1016
rect 1351 767 1368 768
rect 1930 767 1947 768
rect 1349 736 1381 738
rect 1349 697 1352 736
rect 1378 710 1381 736
rect 1369 708 1381 710
rect 1919 730 1951 733
rect 1369 697 1373 708
rect 1919 704 1922 730
rect 1948 704 1951 730
rect 1919 701 1930 704
rect 1371 691 1373 697
rect 1947 701 1951 704
rect 2963 491 2996 493
rect 1919 478 1951 480
rect 1919 452 1922 478
rect 1948 452 1951 478
rect 2963 465 2966 491
rect 2993 465 2996 491
rect 2963 464 2996 465
rect 1919 450 1951 452
rect 2962 461 3004 464
rect 3064 463 3114 464
rect 3064 461 3148 463
rect 2962 450 3148 461
rect 2701 444 2720 449
rect 2745 444 2773 449
rect 2990 447 3080 450
rect 3114 444 3148 450
rect 3181 444 3208 465
<< via1 >>
rect 528 1017 554 1043
rect 2748 1016 2774 1042
rect 1352 713 1378 736
rect 1352 710 1369 713
rect 1369 710 1378 713
rect 1922 713 1948 730
rect 1922 704 1930 713
rect 1930 704 1947 713
rect 1947 704 1948 713
rect 1922 452 1948 478
rect 2966 465 2993 491
<< metal2 >>
rect 525 1043 557 1044
rect 525 1017 528 1043
rect 554 1032 557 1043
rect 2745 1042 2777 1044
rect 2745 1032 2748 1042
rect 554 1017 2748 1032
rect 525 1016 2748 1017
rect 2774 1016 2777 1042
rect 2857 1022 2888 1046
rect 525 1014 2777 1016
rect 501 981 508 999
rect 2968 959 2990 961
rect 1391 921 1475 941
rect 2963 925 2990 959
rect 1436 874 2450 896
rect 2789 875 2824 897
rect 1431 777 2332 799
rect 1349 736 1381 738
rect 1349 710 1352 736
rect 1378 733 1381 736
rect 1378 730 1951 733
rect 1378 710 1922 730
rect 1349 708 1922 710
rect 1919 704 1922 708
rect 1948 704 1951 730
rect 1919 701 1951 704
rect 1436 599 2002 621
rect 1386 569 1434 570
rect 1386 545 1475 569
rect 1980 566 2002 599
rect 2310 616 2332 777
rect 2428 754 2450 874
rect 2970 868 2990 869
rect 2970 835 2992 868
rect 2972 834 2992 835
rect 2865 755 2897 779
rect 3299 778 3310 801
rect 2425 750 2450 754
rect 2425 686 2451 750
rect 3299 696 3310 718
rect 2425 665 2838 686
rect 2817 651 2838 665
rect 2817 630 3019 651
rect 2310 594 2595 616
rect 2417 566 3019 571
rect 1980 550 3019 566
rect 1980 544 2456 550
rect 501 494 509 512
rect 2963 491 2996 493
rect 1919 479 1951 480
rect 2963 479 2966 491
rect 1919 478 2966 479
rect 1919 452 1922 478
rect 1948 465 2966 478
rect 2993 465 2996 491
rect 1948 463 2996 465
rect 1948 462 1988 463
rect 1948 452 1951 462
rect 1919 450 1951 452
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1629137248
transform 1 0 3155 0 1 485
box 0 0 393 746
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1628285143
transform 1 0 2663 0 -1 609
box 133 -454 682 609
use sky130_hilas_FGBias2x1cell  sky130_hilas_FGBias2x1cell_0
timestamp 1629137259
transform 1 0 2040 0 1 826
box 0 0 1654 1052
use sky130_hilas_FGBiasWeakGate2x1cell  sky130_hilas_FGBiasWeakGate2x1cell_0
timestamp 1629137239
transform -1 0 1258 0 1 826
box 0 0 1654 1052
<< labels >>
rlabel metal2 1391 921 1427 940 0 VIN11
port 2 nsew analog default
rlabel metal2 1386 545 1422 570 0 VIN12
port 1 nsew analog default
rlabel metal1 3114 1043 3148 1049 0 VGND
port 7 nsew analog default
rlabel metal1 3180 1043 3208 1049 0 VPWR
port 6 nsew analog default
rlabel metal1 3181 444 3208 450 0 VPWR
port 6 nsew power default
rlabel metal1 3114 444 3148 450 0 VGND
port 7 nsew ground default
rlabel metal2 2865 755 2897 779 0 VIN21
port 3 nsew analog default
rlabel metal2 2857 1022 2888 1046 1 VIN22
port 4 n analog default
rlabel metal1 2745 1041 2773 1049 0 VINJ
port 8 nsew power default
rlabel metal1 2745 444 2773 449 0 VINJ
port 8 nsew power default
rlabel metal2 3299 778 3310 801 0 OUTPUT1
port 9 nsew analog default
rlabel metal2 3299 696 3310 718 0 OUTPUT2
port 10 nsew analog default
rlabel metal2 501 981 508 999 0 DRAIN1
port 11 nsew
rlabel metal2 501 494 509 512 0 DRAIN2
port 12 nsew
rlabel metal1 525 1042 553 1049 0 VINJ
port 8 nsew
rlabel metal1 578 1043 597 1049 0 COLSEL2
port 13 nsew
rlabel metal1 1226 1040 1249 1048 0 GATE2
port 14 nsew
rlabel metal1 1348 1040 1371 1048 0 VGND
port 7 nsew
rlabel metal1 2049 1041 2072 1049 0 GATE1
port 15 nsew
rlabel metal1 1927 1041 1950 1049 0 VGND
port 7 nsew
rlabel metal1 2701 1041 2720 1049 0 COLSEL1
port 16 nsew
rlabel metal1 2701 444 2720 449 0 COLSEL1
port 16 nsew
rlabel metal1 1619 1037 1679 1049 0 VTUN
port 17 nsew
<< end >>
