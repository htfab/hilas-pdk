magic
tech sky130A
timestamp 1628694563
<< error_p >>
rect 146 173 163 174
rect 170 162 171 203
rect 134 150 138 162
rect 170 150 175 162
rect 170 134 171 150
rect 170 102 171 133
rect 170 44 171 73
<< nwell >>
rect 0 304 219 477
<< nmos >>
rect 53 203 86 232
rect 138 203 171 232
rect 53 73 86 102
rect 138 73 171 102
<< pmos >>
rect 21 356 89 386
rect 125 356 193 386
<< ndiff >>
rect 53 256 86 260
rect 53 239 61 256
rect 78 239 86 256
rect 53 232 86 239
rect 138 256 171 260
rect 138 239 146 256
rect 163 239 171 256
rect 138 232 171 239
rect 53 196 86 203
rect 53 179 61 196
rect 78 179 86 196
rect 53 173 86 179
rect 53 125 86 132
rect 53 108 61 125
rect 78 108 86 125
rect 53 102 86 108
rect 138 196 171 203
rect 138 179 146 196
rect 163 179 171 196
rect 138 173 171 179
rect 138 126 171 133
rect 138 109 146 126
rect 163 109 171 126
rect 138 102 171 109
rect 53 66 86 73
rect 53 49 60 66
rect 78 49 86 66
rect 53 45 86 49
rect 138 67 171 73
rect 138 50 145 67
rect 164 50 171 67
rect 138 44 171 50
<< pdiff >>
rect 21 410 89 416
rect 21 393 29 410
rect 47 393 65 410
rect 83 393 89 410
rect 21 386 89 393
rect 125 410 193 416
rect 125 393 133 410
rect 151 393 170 410
rect 189 393 193 410
rect 125 386 193 393
rect 21 349 89 356
rect 21 332 29 349
rect 47 332 65 349
rect 83 332 89 349
rect 21 323 89 332
rect 125 349 193 356
rect 125 332 131 349
rect 149 332 167 349
rect 185 332 193 349
rect 125 328 193 332
rect 132 323 193 328
<< ndiffc >>
rect 61 239 78 256
rect 146 239 163 256
rect 61 179 78 196
rect 61 108 78 125
rect 146 179 163 196
rect 146 109 163 126
rect 60 49 78 66
rect 145 50 164 67
<< pdiffc >>
rect 29 393 47 410
rect 65 393 83 410
rect 133 393 151 410
rect 170 393 189 410
rect 29 332 47 349
rect 65 332 83 349
rect 131 332 149 349
rect 167 332 185 349
<< psubdiff >>
rect 53 161 86 173
rect 53 144 61 161
rect 78 144 86 161
rect 53 132 86 144
rect 138 162 171 173
rect 138 145 146 162
rect 163 145 171 162
rect 138 134 171 145
rect 138 133 170 134
<< nsubdiff >>
rect 21 445 89 457
rect 21 428 29 445
rect 47 428 65 445
rect 83 428 89 445
rect 21 416 89 428
rect 125 445 193 457
rect 125 428 133 445
rect 151 428 170 445
rect 189 428 193 445
rect 125 416 193 428
<< psubdiffcont >>
rect 61 144 78 161
rect 146 145 163 162
<< nsubdiffcont >>
rect 29 428 47 445
rect 65 428 83 445
rect 133 428 151 445
rect 170 428 189 445
<< poly >>
rect 8 356 21 386
rect 89 356 125 386
rect 193 356 206 386
rect 97 312 114 356
rect 91 304 118 312
rect 91 287 96 304
rect 113 287 118 304
rect 91 279 118 287
rect 28 203 53 232
rect 86 203 99 232
rect 124 203 138 232
rect 171 203 194 232
rect 28 102 44 203
rect 178 102 194 203
rect 28 73 53 102
rect 86 73 99 102
rect 123 73 138 102
rect 171 73 194 102
rect 28 34 44 73
rect 28 26 87 34
rect 178 33 194 73
rect 28 9 60 26
rect 78 9 87 26
rect 28 3 87 9
rect 138 25 194 33
rect 138 8 147 25
rect 164 8 194 25
rect 138 3 194 8
<< polycont >>
rect 96 287 113 304
rect 60 9 78 26
rect 147 8 164 25
<< locali >>
rect 21 428 29 445
rect 47 428 65 445
rect 83 428 133 445
rect 151 428 170 445
rect 189 428 197 445
rect 21 410 197 428
rect 21 393 29 410
rect 47 393 65 410
rect 83 393 133 410
rect 151 393 170 410
rect 189 393 197 410
rect 21 332 29 349
rect 47 332 65 349
rect 83 332 92 349
rect 123 332 131 349
rect 149 332 167 349
rect 185 332 193 349
rect 56 315 92 332
rect 56 304 121 315
rect 56 287 96 304
rect 113 287 121 304
rect 56 279 121 287
rect 56 256 83 279
rect 146 257 171 332
rect 138 256 171 257
rect 53 239 61 256
rect 78 239 86 256
rect 138 239 146 256
rect 163 239 171 256
rect 49 179 61 196
rect 78 179 90 196
rect 49 172 90 179
rect 134 179 146 196
rect 163 179 175 196
rect 134 172 175 179
rect 49 162 175 172
rect 49 161 146 162
rect 49 144 61 161
rect 78 145 146 161
rect 163 145 175 162
rect 78 144 175 145
rect 49 134 175 144
rect 49 125 90 134
rect 49 108 61 125
rect 78 108 90 125
rect 134 126 175 134
rect 134 109 146 126
rect 163 109 175 126
rect 52 49 60 66
rect 78 49 86 66
rect 137 50 145 67
rect 164 50 173 67
rect 137 49 173 50
rect 60 26 78 49
rect 60 0 78 9
rect 145 25 164 49
rect 145 8 147 25
rect 145 0 164 8
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
