magic
tech sky130A
timestamp 1634057729
<< checkpaint >>
rect -545 759 804 777
rect -581 694 804 759
rect -586 693 804 694
rect -608 -600 804 693
rect -545 -610 804 -600
<< error_s >>
rect 85 116 112 122
rect 85 74 112 80
rect 137 73 160 79
rect 137 56 140 73
rect 85 49 112 55
rect 137 50 160 56
rect 85 7 112 13
<< nmos >>
rect 85 115 112 116
rect 85 13 112 14
<< ndiff >>
rect 54 115 85 116
rect 112 115 143 116
rect 54 13 85 14
rect 112 13 143 14
<< psubdiff >>
rect 143 106 184 116
rect 143 89 155 106
rect 172 89 184 106
rect 143 80 184 89
rect 143 40 184 49
rect 143 23 155 40
rect 172 23 184 40
rect 143 13 184 23
<< psubdiffcont >>
rect 155 89 172 106
rect 155 23 172 40
<< poly >>
rect 85 128 112 129
rect 13 62 112 72
rect 13 57 85 62
rect 13 49 40 57
rect 85 0 112 1
<< locali >>
rect 138 106 173 114
rect 138 89 155 106
rect 172 89 173 106
rect 118 81 137 82
rect 138 81 173 89
rect 118 48 173 81
rect 138 40 173 48
rect 138 23 155 40
rect 172 23 173 40
rect 138 15 173 23
<< metal2 >>
rect 0 20 33 41
use sky130_hilas_poly2li  sky130_hilas_poly2li_0
timestamp 1634057707
transform 1 0 22 0 1 30
box 0 0 27 33
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1634057708
transform 1 0 147 0 1 58
box 0 0 23 29
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1634057699
transform 1 0 44 0 1 31
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1634057699
transform 1 0 49 0 1 96
box 0 0 34 33
use sky130_hilas_nFET03  sky130_hilas_nFET03_1
timestamp 1634057709
transform 1 0 85 0 1 86
box 0 0 89 61
use sky130_hilas_nFET03  sky130_hilas_nFET03_0
timestamp 1634057709
transform 1 0 85 0 1 20
box 0 0 89 61
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
