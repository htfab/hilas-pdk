magic
tech sky130A
timestamp 1632257806
<< checkpaint >>
rect -630 -248 3387 1717
rect -150 -630 2907 -248
rect -150 -635 1366 -630
rect 1391 -635 2907 -630
<< error_s >>
rect 803 572 832 588
rect 882 572 911 588
rect 961 572 990 588
rect 1040 572 1069 588
rect 1286 574 1315 592
rect 1442 574 1471 592
rect 1688 572 1717 588
rect 1767 572 1796 588
rect 1846 572 1875 588
rect 1925 572 1954 588
rect 1286 542 1287 543
rect 1314 542 1315 543
rect 1442 542 1443 543
rect 1470 542 1471 543
rect 803 538 804 539
rect 831 538 832 539
rect 882 538 883 539
rect 910 538 911 539
rect 961 538 962 539
rect 989 538 990 539
rect 1040 538 1041 539
rect 1068 538 1069 539
rect 753 509 770 538
rect 802 537 833 538
rect 881 537 912 538
rect 960 537 991 538
rect 1039 537 1070 538
rect 803 530 832 537
rect 882 530 911 537
rect 961 530 990 537
rect 1040 530 1069 537
rect 803 516 812 530
rect 1059 516 1069 530
rect 803 510 832 516
rect 882 510 911 516
rect 961 510 990 516
rect 1040 510 1069 516
rect 802 509 833 510
rect 881 509 912 510
rect 960 509 991 510
rect 1039 509 1070 510
rect 1101 509 1119 538
rect 1236 513 1254 542
rect 1285 541 1316 542
rect 1286 532 1315 541
rect 1286 523 1296 532
rect 1305 523 1315 532
rect 1286 514 1315 523
rect 1285 513 1316 514
rect 1347 513 1365 542
rect 1392 513 1410 542
rect 1441 541 1472 542
rect 1442 532 1471 541
rect 1442 523 1452 532
rect 1461 523 1471 532
rect 1442 514 1471 523
rect 1441 513 1472 514
rect 1503 513 1521 542
rect 1688 538 1689 539
rect 1716 538 1717 539
rect 1767 538 1768 539
rect 1795 538 1796 539
rect 1846 538 1847 539
rect 1874 538 1875 539
rect 1925 538 1926 539
rect 1953 538 1954 539
rect 1286 512 1287 513
rect 1314 512 1315 513
rect 1442 512 1443 513
rect 1470 512 1471 513
rect 1638 509 1656 538
rect 1687 537 1718 538
rect 1766 537 1797 538
rect 1845 537 1876 538
rect 1924 537 1955 538
rect 1688 530 1717 537
rect 1767 530 1796 537
rect 1846 530 1875 537
rect 1925 530 1954 537
rect 1688 516 1698 530
rect 1945 516 1954 530
rect 1688 510 1717 516
rect 1767 510 1796 516
rect 1846 510 1875 516
rect 1925 510 1954 516
rect 1687 509 1718 510
rect 1766 509 1797 510
rect 1845 509 1876 510
rect 1924 509 1955 510
rect 1987 509 2004 538
rect 2021 516 2023 517
rect 803 508 804 509
rect 831 508 832 509
rect 882 508 883 509
rect 910 508 911 509
rect 961 508 962 509
rect 989 508 990 509
rect 1040 508 1041 509
rect 1068 508 1069 509
rect 1688 508 1689 509
rect 1716 508 1717 509
rect 1767 508 1768 509
rect 1795 508 1796 509
rect 1846 508 1847 509
rect 1874 508 1875 509
rect 1925 508 1926 509
rect 1953 508 1954 509
rect 803 459 832 474
rect 882 459 911 474
rect 961 459 990 474
rect 1040 459 1069 474
rect 1286 463 1315 481
rect 1442 463 1471 481
rect 1688 459 1717 474
rect 1767 459 1796 474
rect 1846 459 1875 474
rect 1925 459 1954 474
rect 803 425 832 441
rect 882 425 911 441
rect 961 425 990 441
rect 1040 425 1069 441
rect 1286 422 1315 440
rect 1442 422 1471 440
rect 1688 425 1717 441
rect 1767 425 1796 441
rect 1846 425 1875 441
rect 1925 425 1954 441
rect 803 391 804 392
rect 831 391 832 392
rect 882 391 883 392
rect 910 391 911 392
rect 961 391 962 392
rect 989 391 990 392
rect 1040 391 1041 392
rect 1068 391 1069 392
rect 1688 391 1689 392
rect 1716 391 1717 392
rect 1767 391 1768 392
rect 1795 391 1796 392
rect 1846 391 1847 392
rect 1874 391 1875 392
rect 1925 391 1926 392
rect 1953 391 1954 392
rect 753 362 770 391
rect 802 390 833 391
rect 881 390 912 391
rect 960 390 991 391
rect 1039 390 1070 391
rect 803 383 832 390
rect 882 383 911 390
rect 961 383 990 390
rect 1040 383 1069 390
rect 803 369 812 383
rect 1059 369 1069 383
rect 803 363 832 369
rect 882 363 911 369
rect 961 363 990 369
rect 1040 363 1069 369
rect 802 362 833 363
rect 881 362 912 363
rect 960 362 991 363
rect 1039 362 1070 363
rect 1101 362 1119 391
rect 1286 390 1287 391
rect 1314 390 1315 391
rect 1442 390 1443 391
rect 1470 390 1471 391
rect 803 361 804 362
rect 831 361 832 362
rect 882 361 883 362
rect 910 361 911 362
rect 961 361 962 362
rect 989 361 990 362
rect 1040 361 1041 362
rect 1068 361 1069 362
rect 1236 361 1254 390
rect 1285 389 1316 390
rect 1286 380 1315 389
rect 1286 371 1296 380
rect 1305 371 1315 380
rect 1286 362 1315 371
rect 1285 361 1316 362
rect 1347 361 1365 390
rect 1392 361 1410 390
rect 1441 389 1472 390
rect 1442 380 1471 389
rect 1442 371 1452 380
rect 1461 371 1471 380
rect 1442 362 1471 371
rect 1441 361 1472 362
rect 1503 361 1521 390
rect 1638 362 1656 391
rect 1687 390 1718 391
rect 1766 390 1797 391
rect 1845 390 1876 391
rect 1924 390 1955 391
rect 1688 383 1717 390
rect 1767 383 1796 390
rect 1846 383 1875 390
rect 1925 383 1954 390
rect 1688 369 1698 383
rect 1945 369 1954 383
rect 1688 363 1717 369
rect 1767 363 1796 369
rect 1846 363 1875 369
rect 1925 363 1954 369
rect 1687 362 1718 363
rect 1766 362 1797 363
rect 1845 362 1876 363
rect 1924 362 1955 363
rect 1987 362 2004 391
rect 1688 361 1689 362
rect 1716 361 1717 362
rect 1767 361 1768 362
rect 1795 361 1796 362
rect 1846 361 1847 362
rect 1874 361 1875 362
rect 1925 361 1926 362
rect 1953 361 1954 362
rect 1286 360 1287 361
rect 1314 360 1315 361
rect 1442 360 1443 361
rect 1470 360 1471 361
rect 803 312 832 327
rect 882 312 911 327
rect 961 312 990 327
rect 1040 312 1069 327
rect 1286 311 1315 329
rect 1442 311 1471 329
rect 1688 312 1717 327
rect 1767 312 1796 327
rect 1846 312 1875 327
rect 1925 312 1954 327
rect 803 278 832 294
rect 882 278 911 294
rect 961 278 990 294
rect 1040 278 1069 294
rect 1286 277 1315 295
rect 1442 277 1471 295
rect 1688 278 1717 294
rect 1767 278 1796 294
rect 1846 278 1875 294
rect 1925 278 1954 294
rect 1286 245 1287 246
rect 1314 245 1315 246
rect 1442 245 1443 246
rect 1470 245 1471 246
rect 803 244 804 245
rect 831 244 832 245
rect 882 244 883 245
rect 910 244 911 245
rect 961 244 962 245
rect 989 244 990 245
rect 1040 244 1041 245
rect 1068 244 1069 245
rect 753 215 770 244
rect 802 243 833 244
rect 881 243 912 244
rect 960 243 991 244
rect 1039 243 1070 244
rect 803 236 832 243
rect 882 236 911 243
rect 961 236 990 243
rect 1040 236 1069 243
rect 803 222 812 236
rect 1059 222 1069 236
rect 803 216 832 222
rect 882 216 911 222
rect 961 216 990 222
rect 1040 216 1069 222
rect 802 215 833 216
rect 881 215 912 216
rect 960 215 991 216
rect 1039 215 1070 216
rect 1101 215 1119 244
rect 1236 216 1254 245
rect 1285 244 1316 245
rect 1286 235 1315 244
rect 1286 226 1296 235
rect 1305 226 1315 235
rect 1286 217 1315 226
rect 1285 216 1316 217
rect 1347 216 1365 245
rect 1392 216 1410 245
rect 1441 244 1472 245
rect 1442 235 1471 244
rect 1442 226 1452 235
rect 1461 226 1471 235
rect 1442 217 1471 226
rect 1441 216 1472 217
rect 1503 216 1521 245
rect 1688 244 1689 245
rect 1716 244 1717 245
rect 1767 244 1768 245
rect 1795 244 1796 245
rect 1846 244 1847 245
rect 1874 244 1875 245
rect 1925 244 1926 245
rect 1953 244 1954 245
rect 1286 215 1287 216
rect 1314 215 1315 216
rect 1442 215 1443 216
rect 1470 215 1471 216
rect 1638 215 1656 244
rect 1687 243 1718 244
rect 1766 243 1797 244
rect 1845 243 1876 244
rect 1924 243 1955 244
rect 1688 236 1717 243
rect 1767 236 1796 243
rect 1846 236 1875 243
rect 1925 236 1954 243
rect 1688 222 1698 236
rect 1945 222 1954 236
rect 1688 216 1717 222
rect 1767 216 1796 222
rect 1846 216 1875 222
rect 1925 216 1954 222
rect 1687 215 1718 216
rect 1766 215 1797 216
rect 1845 215 1876 216
rect 1924 215 1955 216
rect 1987 215 2004 244
rect 803 214 804 215
rect 831 214 832 215
rect 882 214 883 215
rect 910 214 911 215
rect 961 214 962 215
rect 989 214 990 215
rect 1040 214 1041 215
rect 1068 214 1069 215
rect 1688 214 1689 215
rect 1716 214 1717 215
rect 1767 214 1768 215
rect 1795 214 1796 215
rect 1846 214 1847 215
rect 1874 214 1875 215
rect 1925 214 1926 215
rect 1953 214 1954 215
rect 803 165 832 180
rect 882 165 911 180
rect 961 165 990 180
rect 1040 165 1069 180
rect 1286 166 1315 184
rect 1442 166 1471 184
rect 1688 165 1717 180
rect 1767 165 1796 180
rect 1846 165 1875 180
rect 1925 165 1954 180
rect 803 131 832 147
rect 882 131 911 147
rect 961 131 990 147
rect 1040 131 1069 147
rect 1286 123 1315 141
rect 1442 123 1471 141
rect 1688 131 1717 147
rect 1767 131 1796 147
rect 1846 131 1875 147
rect 1925 131 1954 147
rect 803 97 804 98
rect 831 97 832 98
rect 882 97 883 98
rect 910 97 911 98
rect 961 97 962 98
rect 989 97 990 98
rect 1040 97 1041 98
rect 1068 97 1069 98
rect 1688 97 1689 98
rect 1716 97 1717 98
rect 1767 97 1768 98
rect 1795 97 1796 98
rect 1846 97 1847 98
rect 1874 97 1875 98
rect 1925 97 1926 98
rect 1953 97 1954 98
rect 753 68 770 97
rect 802 96 833 97
rect 881 96 912 97
rect 960 96 991 97
rect 1039 96 1070 97
rect 803 89 832 96
rect 882 89 911 96
rect 961 89 990 96
rect 1040 89 1069 96
rect 803 75 812 89
rect 1059 75 1069 89
rect 803 69 832 75
rect 882 69 911 75
rect 961 69 990 75
rect 1040 69 1069 75
rect 802 68 833 69
rect 881 68 912 69
rect 960 68 991 69
rect 1039 68 1070 69
rect 1101 68 1119 97
rect 1286 91 1287 92
rect 1314 91 1315 92
rect 1442 91 1443 92
rect 1470 91 1471 92
rect 803 67 804 68
rect 831 67 832 68
rect 882 67 883 68
rect 910 67 911 68
rect 961 67 962 68
rect 989 67 990 68
rect 1040 67 1041 68
rect 1068 67 1069 68
rect 1236 62 1254 91
rect 1285 90 1316 91
rect 1286 81 1315 90
rect 1286 72 1296 81
rect 1305 72 1315 81
rect 1286 63 1315 72
rect 1285 62 1316 63
rect 1347 62 1365 91
rect 1392 62 1410 91
rect 1441 90 1472 91
rect 1442 81 1471 90
rect 1442 72 1452 81
rect 1461 72 1471 81
rect 1442 63 1471 72
rect 1441 62 1472 63
rect 1503 62 1521 91
rect 1638 68 1656 97
rect 1687 96 1718 97
rect 1766 96 1797 97
rect 1845 96 1876 97
rect 1924 96 1955 97
rect 1688 89 1717 96
rect 1767 89 1796 96
rect 1846 89 1875 96
rect 1925 89 1954 96
rect 1688 75 1698 89
rect 1945 75 1954 89
rect 1688 69 1717 75
rect 1767 69 1796 75
rect 1846 69 1875 75
rect 1925 69 1954 75
rect 1687 68 1718 69
rect 1766 68 1797 69
rect 1845 68 1876 69
rect 1924 68 1955 69
rect 1987 68 2004 97
rect 1688 67 1689 68
rect 1716 67 1717 68
rect 1767 67 1768 68
rect 1795 67 1796 68
rect 1846 67 1847 68
rect 1874 67 1875 68
rect 1925 67 1926 68
rect 1953 67 1954 68
rect 1286 61 1287 62
rect 1314 61 1315 62
rect 1442 61 1443 62
rect 1470 61 1471 62
rect 803 18 832 33
rect 882 18 911 33
rect 961 18 990 33
rect 1040 18 1069 33
rect 1286 12 1315 30
rect 1442 12 1471 30
rect 1688 18 1717 33
rect 1767 18 1796 33
rect 1846 18 1875 33
rect 1925 18 1954 33
<< metal1 >>
rect 516 599 532 605
rect 557 599 576 605
rect 597 599 613 605
rect 516 1 532 8
rect 557 1 576 8
rect 597 1 613 8
rect 924 0 949 605
rect 1285 0 1315 605
rect 1443 0 1473 605
rect 1809 0 1833 605
rect 2144 598 2160 605
rect 2181 598 2200 605
rect 2225 598 2241 605
rect 2144 1 2160 8
rect 2181 1 2200 8
rect 2225 1 2241 8
<< metal2 >>
rect 480 537 488 555
rect 2266 537 2277 555
rect 480 494 488 512
rect 2267 494 2278 512
rect 480 394 488 412
rect 2267 394 2278 412
rect 480 351 488 369
rect 720 361 732 369
rect 2029 355 2041 369
rect 2267 351 2278 369
rect 480 236 487 254
rect 2266 236 2277 254
rect 480 193 487 211
rect 2266 193 2277 211
rect 480 94 487 112
rect 2266 94 2277 112
rect 480 51 487 69
rect 2266 51 2277 69
use sky130_hilas_swc4x1cellOverlap2  sky130_hilas_swc4x1cellOverlap2_1
timestamp 1632256376
transform -1 0 1224 0 1 382
box 0 0 1224 705
use sky130_hilas_swc4x1cellOverlap2  sky130_hilas_swc4x1cellOverlap2_0
timestamp 1632256376
transform 1 0 1533 0 1 382
box 0 0 1224 705
<< labels >>
rlabel metal1 597 599 613 605 0 VERT1
port 1 nsew analog default
rlabel metal1 516 599 532 605 0 VINJ
port 10 nsew
rlabel metal1 557 599 576 605 0 GATESELECT1
port 11 nsew analog default
rlabel metal2 480 537 488 555 0 DRAIN1
port 3 nsew analog default
rlabel metal2 480 494 488 512 0 HORIZ1
port 2 nsew analog default
rlabel metal2 480 394 488 412 0 HORIZ2
port 4 nsew analog default
rlabel metal2 480 351 488 369 0 DRAIN2
port 5 nsew analog default
rlabel metal2 480 236 487 254 0 DRAIN3
port 6 nsew analog default
rlabel metal2 480 193 487 211 0 HORIZ3
port 7 nsew analog default
rlabel metal2 480 94 487 112 0 HORIZ4
port 8 nsew analog default
rlabel metal2 480 51 487 69 0 DRAIN4
port 9 nsew analog default
rlabel metal1 516 1 532 8 0 VINJ
port 10 nsew power default
rlabel metal1 597 1 613 8 0 VERT1
port 1 nsew analog default
rlabel metal1 557 1 576 8 0 GATESELECT1
port 11 nsew analog default
rlabel metal1 2225 1 2241 8 0 VINJ
port 10 nsew power default
rlabel metal1 2144 598 2160 605 0 VERT2
port 12 nsew analog default
rlabel metal1 2181 598 2200 605 0 GATESELECT2
port 13 nsew analog default
rlabel metal1 2225 598 2241 605 0 VINJ
port 10 nsew power default
rlabel metal1 2144 1 2160 8 0 VERT2
port 12 nsew analog default
rlabel metal1 2181 1 2200 8 0 GATESELECT2
port 13 nsew analog default
rlabel metal2 2266 537 2277 555 0 DRAIN1
port 3 nsew analog default
rlabel metal2 2267 494 2278 512 0 HORIZ1
port 2 nsew analog default
rlabel metal2 2267 394 2278 412 0 HORIZ2
port 4 nsew analog default
rlabel metal2 2267 351 2278 369 0 DRAIN2
port 5 nsew analog default
rlabel metal2 2266 236 2277 254 0 DRAIN3
port 6 nsew analog default
rlabel metal2 2266 193 2277 211 0 HORIZ3
port 7 nsew analog default
rlabel metal2 2266 94 2277 112 0 HORIZ4
port 8 nsew analog default
rlabel metal2 2266 51 2277 69 0 DRAIN
port 14 nsew analog default
rlabel metal1 1809 600 1833 605 0 GATE2
port 15 nsew analog default
rlabel metal1 1809 0 1833 6 0 GATE2
port 15 nsew analog default
rlabel metal1 924 599 949 605 0 GATE1
port 16 nsew analog default
rlabel metal1 924 0 949 6 0 GATE1
port 16 nsew analog default
rlabel metal1 1285 597 1315 605 0 VTUN
port 17 nsew analog default
rlabel metal1 1443 597 1473 605 0 VTUN
rlabel metal1 1285 0 1315 8 0 VTUN
port 17 nsew analog default
rlabel metal1 1443 0 1473 8 0 VTUN
port 17 nsew analog default
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
