magic
tech sky130A
timestamp 1628616748
<< checkpaint >>
rect -132 761 1151 769
rect -142 -520 1151 761
rect -142 -528 1141 -520
<< error_s >>
rect 85 136 135 142
rect 405 136 455 142
rect 85 94 135 100
rect 405 94 455 100
rect 85 70 135 75
rect 225 69 275 75
rect 405 70 455 75
rect 85 28 135 33
rect 225 27 275 33
rect 405 28 455 33
<< nwell >>
rect 0 0 342 169
<< mvnmos >>
rect 405 100 455 136
rect 405 33 455 70
<< mvpmos >>
rect 85 100 135 136
rect 85 33 135 70
rect 225 33 275 69
<< mvndiff >>
rect 377 124 405 136
rect 377 107 382 124
rect 399 107 405 124
rect 377 100 405 107
rect 455 124 483 136
rect 455 107 461 124
rect 478 107 483 124
rect 455 100 483 107
rect 377 62 405 70
rect 377 45 382 62
rect 399 45 405 62
rect 377 33 405 45
rect 455 62 483 70
rect 455 45 461 62
rect 478 45 483 62
rect 455 33 483 45
<< mvpdiff >>
rect 55 123 85 136
rect 55 106 62 123
rect 79 106 85 123
rect 55 100 85 106
rect 135 124 165 136
rect 135 107 141 124
rect 158 107 165 124
rect 135 100 165 107
rect 55 63 85 70
rect 55 46 62 63
rect 79 46 85 63
rect 55 33 85 46
rect 135 62 165 70
rect 135 45 141 62
rect 159 45 165 62
rect 135 33 165 45
rect 195 62 225 69
rect 195 45 202 62
rect 219 45 225 62
rect 195 33 225 45
rect 275 62 305 69
rect 275 45 281 62
rect 298 45 305 62
rect 275 33 305 45
<< mvndiffc >>
rect 382 107 399 124
rect 461 107 478 124
rect 382 45 399 62
rect 461 45 478 62
<< mvpdiffc >>
rect 62 106 79 123
rect 141 107 158 124
rect 62 46 79 63
rect 141 45 159 62
rect 202 45 219 62
rect 281 45 298 62
<< psubdiff >>
rect 515 67 546 79
rect 515 50 519 67
rect 536 50 546 67
rect 515 38 546 50
<< nsubdiff >>
rect 18 101 43 131
rect 18 84 22 101
rect 39 84 43 101
rect 18 67 43 84
rect 18 50 22 67
rect 39 50 43 67
rect 18 38 43 50
<< psubdiffcont >>
rect 519 50 536 67
<< nsubdiffcont >>
rect 22 84 39 101
rect 22 50 39 67
<< poly >>
rect 85 144 551 159
rect 85 136 135 144
rect 405 136 455 144
rect 515 141 551 144
rect 181 112 221 116
rect 181 110 275 112
rect 85 70 135 100
rect 181 93 189 110
rect 206 93 275 110
rect 515 124 526 141
rect 543 124 551 141
rect 515 119 551 124
rect 181 88 275 93
rect 225 69 275 88
rect 405 70 455 100
rect 85 20 135 33
rect 225 20 275 33
rect 405 20 455 33
<< polycont >>
rect 189 93 206 110
rect 526 124 543 141
<< locali >>
rect 526 141 543 149
rect 62 123 79 131
rect 22 101 39 105
rect 22 67 39 69
rect 132 107 141 124
rect 158 110 382 124
rect 158 107 189 110
rect 62 95 79 106
rect 180 93 189 107
rect 206 107 382 110
rect 399 107 407 124
rect 453 107 461 124
rect 478 107 490 124
rect 526 114 543 124
rect 206 93 214 107
rect 526 97 532 114
rect 526 93 543 97
rect 180 89 214 93
rect 62 63 79 78
rect 519 67 536 75
rect 62 38 79 46
rect 132 45 141 62
rect 159 46 160 62
rect 431 62 455 66
rect 177 46 202 62
rect 159 45 202 46
rect 219 45 228 62
rect 273 45 281 62
rect 298 45 360 62
rect 377 45 382 62
rect 399 45 407 62
rect 431 45 435 62
rect 452 45 461 62
rect 478 45 488 62
rect 431 42 455 45
<< viali >>
rect 22 105 39 122
rect 22 84 39 86
rect 22 69 39 84
rect 22 33 39 50
rect 62 78 79 95
rect 532 97 549 114
rect 160 46 177 63
rect 360 45 377 62
rect 435 45 452 62
rect 519 33 536 50
<< metal1 >>
rect 58 134 83 169
rect 19 122 83 134
rect 19 105 22 122
rect 39 105 83 122
rect 19 95 83 105
rect 19 86 62 95
rect 19 69 22 86
rect 39 78 62 86
rect 79 78 83 95
rect 39 69 83 78
rect 19 50 83 69
rect 173 67 207 70
rect 173 66 178 67
rect 19 33 22 50
rect 39 33 83 50
rect 151 63 178 66
rect 151 46 160 63
rect 177 46 178 63
rect 151 43 178 46
rect 173 41 178 43
rect 204 62 207 67
rect 357 62 380 170
rect 492 76 511 170
rect 525 119 557 120
rect 525 93 528 119
rect 554 93 557 119
rect 525 92 557 93
rect 204 45 219 62
rect 357 45 360 62
rect 377 45 380 62
rect 204 41 207 45
rect 173 38 207 41
rect 19 27 83 33
rect 58 5 83 27
rect 357 5 380 45
rect 416 67 453 68
rect 416 41 419 67
rect 445 62 458 67
rect 452 45 458 62
rect 445 41 458 45
rect 492 50 539 76
rect 416 39 453 41
rect 492 33 519 50
rect 536 33 539 50
rect 492 27 539 33
rect 492 5 511 27
<< via1 >>
rect 178 41 204 67
rect 528 114 554 119
rect 528 97 532 114
rect 532 97 549 114
rect 549 97 554 114
rect 528 93 554 97
rect 419 62 445 67
rect 419 45 435 62
rect 435 45 445 62
rect 419 41 445 45
<< metal2 >>
rect 524 119 558 121
rect 524 93 528 119
rect 554 114 558 119
rect 554 93 568 114
rect 524 91 568 93
rect 416 67 448 70
rect 175 41 178 67
rect 204 62 207 67
rect 416 62 419 67
rect 204 43 419 62
rect 204 41 207 43
rect 416 41 419 43
rect 445 41 448 67
rect 416 38 448 41
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1628616665
transform 1 0 498 0 1 110
box 0 0 23 29
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
