magic
tech sky130A
timestamp 1637953024
<< error_s >>
rect 129 648 181 654
rect 181 647 209 648
rect 483 647 533 652
rect 129 606 181 612
rect 483 605 533 610
rect 55 581 108 586
rect 202 581 254 586
rect 412 580 462 586
rect 554 580 604 586
rect -553 573 -500 580
rect -374 572 -322 580
rect 55 539 108 544
rect 202 539 254 544
rect 412 538 462 544
rect 554 538 604 544
rect -553 531 -500 538
rect -374 530 -322 538
rect 129 488 181 494
rect 181 487 209 488
rect 483 487 533 492
rect 129 446 181 452
rect 483 445 533 450
rect -553 422 -500 429
rect -374 421 -322 429
rect 55 421 108 426
rect 202 421 254 426
rect 412 420 462 426
rect 554 420 604 426
rect -553 380 -500 387
rect -374 379 -322 387
rect 55 379 108 384
rect 202 379 254 384
rect 412 378 462 384
rect 554 378 604 384
rect 129 328 181 334
rect 181 327 209 328
rect 483 327 533 332
rect 129 286 181 292
rect 483 285 533 290
rect -553 271 -500 278
rect -374 270 -322 278
rect 55 261 108 266
rect 202 261 254 266
rect 412 260 462 266
rect 554 260 604 266
rect -553 229 -500 236
rect -374 228 -322 236
rect 55 219 108 224
rect 202 219 254 224
rect 412 218 462 224
rect 554 218 604 224
rect 129 168 181 174
rect 181 167 209 168
rect 483 167 533 172
rect 129 126 181 132
rect 483 125 533 130
rect 55 101 108 106
rect 202 101 254 106
rect 412 100 462 106
rect 554 100 604 106
rect 55 59 108 64
rect 202 59 254 64
rect 412 58 462 64
rect 554 58 604 64
<< nwell >>
rect -29 679 315 681
rect 32 659 54 665
rect 32 64 54 69
rect -29 31 315 35
<< metal1 >>
rect -576 658 -554 681
rect -319 657 -296 681
rect -270 631 -243 660
rect 32 659 54 665
rect 529 661 556 666
rect -274 604 -271 631
rect -244 604 -241 631
rect -178 612 -151 617
rect -270 526 -243 604
rect -271 523 -243 526
rect -244 496 -243 523
rect -271 493 -243 496
rect -270 490 -243 493
rect -224 563 -197 570
rect -224 358 -197 536
rect -178 471 -151 585
rect -83 567 -54 572
rect -85 564 -54 567
rect -56 535 -54 564
rect -85 532 -54 535
rect -183 444 -180 471
rect -153 444 -150 471
rect -225 355 -197 358
rect -198 328 -197 355
rect -225 325 -197 328
rect -576 31 -554 235
rect -319 31 -296 236
rect -224 189 -197 325
rect -178 313 -151 444
rect -180 310 -151 313
rect -153 283 -151 310
rect -180 280 -151 283
rect -178 278 -151 280
rect -131 417 -104 423
rect -131 414 -103 417
rect -131 387 -130 414
rect -131 384 -103 387
rect -83 410 -54 532
rect -83 384 -81 410
rect -55 384 -54 410
rect -228 186 -193 189
rect -228 159 -224 186
rect -197 159 -193 186
rect -228 156 -193 159
rect -131 143 -104 384
rect -83 267 -54 384
rect -83 264 -53 267
rect -83 235 -82 264
rect -83 232 -53 235
rect -135 141 -100 143
rect -135 114 -131 141
rect -104 114 -100 141
rect -135 111 -100 114
rect -83 95 -54 232
rect -87 93 -50 95
rect -87 64 -83 93
rect -54 64 -50 93
rect 32 64 54 69
rect 529 64 556 69
rect -87 61 -50 64
rect 32 31 54 39
rect 529 31 556 39
<< via1 >>
rect -271 604 -244 631
rect -178 585 -151 612
rect -271 496 -244 523
rect -224 536 -197 563
rect -85 535 -56 564
rect -180 444 -153 471
rect -225 328 -198 355
rect -180 283 -153 310
rect -130 387 -103 414
rect -81 384 -55 410
rect -224 159 -197 186
rect -82 235 -53 264
rect -131 114 -104 141
rect -83 64 -54 93
<< metal2 >>
rect -268 644 -13 660
rect -268 634 -242 644
rect -271 631 -242 634
rect -637 609 -626 627
rect -294 609 -271 627
rect -244 629 -242 631
rect -244 609 -241 629
rect -162 612 -29 615
rect -271 601 -244 604
rect -181 585 -178 612
rect -151 599 -29 612
rect -151 585 -148 599
rect -54 564 -29 566
rect -227 560 -224 563
rect -294 542 -224 560
rect -227 536 -224 542
rect -197 560 -194 563
rect -197 541 -192 560
rect -197 536 -194 541
rect -88 535 -85 564
rect -56 550 -29 564
rect -56 535 -53 550
rect 681 546 694 563
rect -274 496 -271 523
rect -244 517 -241 523
rect -244 501 -110 517
rect -244 496 -241 501
rect -126 500 -110 501
rect -126 484 -30 500
rect -637 458 -626 476
rect -294 474 -158 476
rect -294 471 -153 474
rect -294 458 -180 471
rect -153 444 -152 455
rect -180 441 -152 444
rect -175 439 -152 441
rect -125 439 -29 455
rect -125 414 -109 439
rect -133 409 -130 414
rect -294 391 -130 409
rect -133 387 -130 391
rect -103 387 -100 414
rect -84 384 -81 410
rect -55 406 -52 410
rect -55 390 -29 406
rect -55 384 -52 390
rect 681 386 694 403
rect -228 328 -225 355
rect -198 340 -195 355
rect -198 328 -14 340
rect -637 307 -626 325
rect -228 324 -14 328
rect -183 283 -180 310
rect -153 295 -150 310
rect -153 283 -14 295
rect -182 279 -14 283
rect -85 258 -82 264
rect -294 240 -82 258
rect -85 235 -82 240
rect -53 249 -50 264
rect -53 246 -23 249
rect -53 230 -29 246
rect 681 226 694 243
rect -227 186 -194 188
rect -227 159 -224 186
rect -197 180 -194 186
rect -197 164 -14 180
rect -197 159 -194 164
rect -227 157 -194 159
rect -134 141 -101 142
rect -134 114 -131 141
rect -104 135 -101 141
rect -104 119 -14 135
rect -104 114 -101 119
rect -134 112 -101 114
rect -86 93 -51 94
rect -86 64 -83 93
rect -54 86 -51 93
rect -54 70 -20 86
rect -54 64 -51 70
rect 681 66 694 83
rect -86 63 -51 64
use sky130_hilas_VinjInv2  VinjInv2_2
timestamp 1637952898
transform 1 0 -301 0 1 60
box -336 143 25 308
use sky130_hilas_VinjInv2  VinjInv2_1
timestamp 1637952898
transform 1 0 -301 0 1 211
box -336 143 25 308
use sky130_hilas_VinjInv2  VinjInv2_0
timestamp 1637952898
transform 1 0 -301 0 1 362
box -336 143 25 308
use sky130_hilas_VinjNOR3  VinjNOR3_2
timestamp 1637951121
transform 1 0 307 0 1 211
box -337 140 387 310
use sky130_hilas_VinjNOR3  VinjNOR3_3
timestamp 1637951121
transform 1 0 307 0 1 371
box -337 140 387 310
use sky130_hilas_VinjNOR3  VinjNOR3_1
timestamp 1637951121
transform 1 0 307 0 1 51
box -337 140 387 310
use sky130_hilas_VinjNOR3  VinjNOR3_0
timestamp 1637951121
transform 1 0 307 0 1 -109
box -337 140 387 310
<< labels >>
rlabel metal1 529 661 556 666 0 VGND
port 5 nsew
rlabel metal1 529 64 556 69 0 VGND
port 5 nsew
rlabel metal1 32 64 54 69 0 VINJ
port 6 nsew
rlabel metal1 32 659 54 665 0 VINJ
port 6 nsew
rlabel metal2 -637 609 -626 627 0 IN1
port 8 nsew
rlabel metal2 -637 458 -626 476 0 IN2
port 7 nsew
rlabel metal2 -637 307 -626 325 0 ENABLE
port 9 nsew
rlabel metal1 -576 658 -554 666 0 VINJ
port 6 nsew
rlabel metal1 -319 657 -296 666 0 VGND
port 5 nsew
rlabel metal2 681 546 694 563 0 OUTPUT00
port 1 nsew
rlabel metal2 681 386 694 403 0 OUTPUT01
port 2 nsew
rlabel metal2 681 226 694 243 0 OUTPUT10
port 3 nsew
rlabel metal2 681 66 694 83 0 OUTPUT11
port 4 nsew
<< end >>
