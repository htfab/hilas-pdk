VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_hilas_TA2Cell_1FG_Strong
  CLASS CORE ;
  FOREIGN sky130_hilas_TA2Cell_1FG_Strong ;
  ORIGIN 0.000 0.000 ;
  SIZE 32.050 BY 9.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 14.710 5.900 15.130 6.050 ;
        RECT 15.740 5.900 16.160 6.050 ;
        RECT 14.710 5.760 16.160 5.900 ;
    END
  END VTUN
  PIN PROG
    PORT
      LAYER met1 ;
        RECT 7.470 5.990 7.680 6.050 ;
    END
  END PROG
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT 19.440 5.970 19.670 6.050 ;
    END
  END GATE1
  PIN VIN11
    PORT
      LAYER met1 ;
        RECT 6.590 5.940 6.800 6.050 ;
    END
  END VIN11
  PIN VINJ
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 1.770 5.970 2.080 6.160 ;
        RECT 4.150 5.970 4.470 6.030 ;
        RECT 1.770 5.910 11.520 5.970 ;
        RECT 26.420 5.910 26.740 6.030 ;
        RECT 1.770 5.830 26.740 5.910 ;
        RECT 1.800 5.780 26.740 5.830 ;
        RECT 4.150 5.730 26.740 5.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 26.400 6.030 26.680 6.050 ;
        RECT 26.400 5.970 26.740 6.030 ;
        RECT 26.420 5.730 26.740 5.970 ;
      LAYER via ;
        RECT 26.450 5.750 26.710 6.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 26.400 0.000 26.680 0.050 ;
    END
  END VINJ
  PIN VIN22
    ANTENNAGATEAREA 4.153100 ;
    ANTENNADIFFAREA 8.050300 ;
    PORT
      LAYER nwell ;
        RECT 27.570 6.050 30.880 9.870 ;
        RECT 26.920 6.040 32.050 6.050 ;
        RECT 26.910 3.830 32.050 6.040 ;
        RECT 26.910 0.000 28.770 3.830 ;
        RECT 30.770 0.000 32.050 3.830 ;
      LAYER met2 ;
        RECT 29.490 7.010 29.810 7.270 ;
        RECT 29.530 6.990 30.710 7.010 ;
        RECT 29.530 6.730 30.750 6.990 ;
        RECT 29.530 6.670 30.710 6.730 ;
        RECT 29.490 6.660 30.710 6.670 ;
        RECT 29.490 6.410 29.810 6.660 ;
        RECT 28.160 6.030 28.470 6.040 ;
        RECT 27.590 6.020 28.470 6.030 ;
        RECT 27.520 5.780 28.470 6.020 ;
        RECT 28.160 5.710 28.470 5.780 ;
        RECT 29.130 5.710 29.440 5.760 ;
        RECT 31.380 5.710 31.690 5.810 ;
        RECT 28.550 5.590 28.860 5.660 ;
        RECT 29.130 5.590 31.690 5.710 ;
        RECT 28.550 5.480 31.690 5.590 ;
        RECT 28.550 5.380 30.880 5.480 ;
        RECT 28.550 5.330 28.860 5.380 ;
        RECT 28.310 5.170 28.620 5.210 ;
        RECT 28.130 5.030 28.850 5.170 ;
        RECT 29.080 5.030 29.390 5.110 ;
        RECT 28.130 4.920 29.390 5.030 ;
        RECT 28.310 4.880 29.390 4.920 ;
        RECT 28.580 4.820 29.390 4.880 ;
        RECT 28.580 4.810 28.850 4.820 ;
        RECT 29.080 4.780 29.390 4.820 ;
        RECT 27.190 4.530 27.500 4.670 ;
        RECT 26.840 4.490 27.500 4.530 ;
        RECT 28.400 4.500 28.710 4.640 ;
        RECT 28.400 4.490 30.880 4.500 ;
        RECT 19.350 4.340 30.880 4.490 ;
        RECT 26.840 4.310 27.190 4.340 ;
        RECT 28.400 4.320 30.880 4.340 ;
        RECT 28.400 4.310 28.710 4.320 ;
        RECT 28.650 4.240 28.850 4.250 ;
        RECT 28.650 4.230 28.870 4.240 ;
        RECT 29.080 4.230 29.390 4.270 ;
        RECT 28.650 4.160 29.390 4.230 ;
        RECT 28.360 4.140 29.390 4.160 ;
        RECT 28.310 4.020 29.390 4.140 ;
        RECT 28.310 3.900 28.870 4.020 ;
        RECT 29.080 3.940 29.390 4.020 ;
        RECT 28.310 3.890 28.780 3.900 ;
        RECT 28.560 0.350 28.880 0.500 ;
        RECT 12.370 0.200 28.880 0.350 ;
        RECT 12.370 0.050 12.690 0.200 ;
        RECT 18.170 0.050 18.490 0.200 ;
    END
  END VIN22
  PIN VIN21
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT 27.920 3.350 28.230 3.390 ;
        RECT 27.600 3.340 28.260 3.350 ;
        RECT 27.600 3.110 28.700 3.340 ;
        RECT 27.920 3.060 28.230 3.110 ;
    END
  END VIN21
  PIN VPWR
    ANTENNADIFFAREA 1.373600 ;
    PORT
      LAYER met1 ;
        RECT 30.750 5.900 31.030 6.050 ;
        RECT 30.760 4.470 31.030 5.900 ;
        RECT 30.760 4.180 31.040 4.470 ;
        RECT 30.760 1.880 31.030 4.180 ;
        RECT 30.760 1.590 31.040 1.880 ;
        RECT 30.760 0.000 31.030 1.590 ;
    END
  END VPWR
  PIN VGND
    ANTENNAGATEAREA 3.745100 ;
    ANTENNADIFFAREA 3.678400 ;
    PORT
      LAYER met1 ;
        RECT 29.920 8.410 30.110 9.870 ;
        RECT 30.360 9.220 30.640 9.870 ;
        RECT 30.250 8.620 30.640 9.220 ;
        RECT 29.920 8.380 30.140 8.410 ;
        RECT 29.900 8.110 30.150 8.380 ;
        RECT 29.910 8.100 30.150 8.110 ;
        RECT 29.910 7.860 30.140 8.100 ;
        RECT 29.520 6.380 29.780 6.700 ;
        RECT 29.520 6.260 29.760 6.380 ;
        RECT 29.950 6.050 30.110 7.860 ;
        RECT 30.360 7.020 30.640 8.620 ;
        RECT 30.360 6.700 30.720 7.020 ;
        RECT 30.360 6.050 30.640 6.700 ;
        RECT 28.150 5.710 28.470 6.030 ;
        RECT 29.950 5.830 30.640 6.050 ;
        RECT 29.130 5.430 29.450 5.750 ;
        RECT 29.910 5.580 30.640 5.830 ;
        RECT 29.900 5.310 30.640 5.580 ;
        RECT 29.080 4.780 29.400 5.100 ;
        RECT 28.400 4.200 28.710 4.640 ;
        RECT 28.410 4.190 28.620 4.200 ;
        RECT 28.390 3.870 28.650 4.190 ;
        RECT 29.080 3.950 29.400 4.270 ;
        RECT 28.410 2.580 28.620 3.870 ;
        RECT 29.920 3.820 30.640 5.310 ;
        RECT 28.390 2.290 28.620 2.580 ;
        RECT 28.560 0.200 28.880 0.500 ;
        RECT 30.090 0.200 30.430 3.820 ;
        RECT 28.560 0.140 30.430 0.200 ;
        RECT 28.610 0.060 30.430 0.140 ;
        RECT 30.090 0.000 30.430 0.060 ;
      LAYER via ;
        RECT 29.520 6.410 29.780 6.670 ;
        RECT 30.460 6.730 30.720 6.990 ;
        RECT 28.180 5.740 28.440 6.000 ;
        RECT 29.160 5.460 29.420 5.720 ;
        RECT 29.110 4.810 29.370 5.070 ;
        RECT 28.430 4.350 28.690 4.610 ;
        RECT 28.390 3.900 28.650 4.160 ;
        RECT 29.110 3.980 29.370 4.240 ;
        RECT 28.590 0.220 28.850 0.480 ;
    END
  END VGND
  PIN OUTPUT2
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER met2 ;
        RECT 29.130 2.740 29.440 2.800 ;
        RECT 31.420 2.740 31.730 2.870 ;
        RECT 29.130 2.520 32.050 2.740 ;
        RECT 29.130 2.470 29.440 2.520 ;
    END
  END OUTPUT2
  PIN OUTPUT1
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER met2 ;
        RECT 29.130 3.570 29.440 3.620 ;
        RECT 31.430 3.570 31.740 3.590 ;
        RECT 29.130 3.340 32.050 3.570 ;
        RECT 29.130 3.290 29.440 3.340 ;
        RECT 31.430 3.260 31.740 3.340 ;
    END
  END OUTPUT1
  PIN GATESEL1
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER met1 ;
        RECT 4.600 6.050 4.780 9.870 ;
        RECT 4.600 5.990 4.910 6.050 ;
        RECT 4.600 5.340 4.780 5.990 ;
        RECT 4.540 5.000 4.830 5.340 ;
        RECT 4.600 3.820 4.780 5.000 ;
    END
  END GATESEL1
  PIN GATESEL2
    PORT
      LAYER met1 ;
        RECT 25.960 0.000 26.150 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.960 5.970 26.150 6.050 ;
    END
  END GATESEL2
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 3.950 5.370 4.030 5.550 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 3.950 0.500 4.030 0.680 ;
    END
  END DRAIN2
  PIN VIN12
    PORT
      LAYER met1 ;
        RECT 6.600 0.010 6.830 0.130 ;
    END
  END VIN12
  PIN GATE2
    PORT
      LAYER met1 ;
        RECT 7.060 5.970 7.250 6.050 ;
    END
  END GATE2
  PIN RUN
    ANTENNADIFFAREA 1.850000 ;
    PORT
      LAYER met1 ;
        RECT 8.470 6.050 8.700 9.870 ;
        RECT 8.470 5.980 8.730 6.050 ;
        RECT 8.470 3.820 8.700 5.980 ;
    END
  END RUN
  OBS
      LAYER nwell ;
        RECT 0.000 3.830 3.310 9.860 ;
        RECT 5.040 7.480 7.760 9.130 ;
        RECT 9.790 9.120 11.520 9.870 ;
        RECT 5.040 7.440 7.750 7.480 ;
        RECT 5.040 6.110 7.750 6.150 ;
        RECT 5.040 6.050 7.760 6.110 ;
        RECT 3.950 6.040 7.760 6.050 ;
        RECT 4.150 5.730 4.470 6.030 ;
        RECT 5.040 4.460 7.760 6.040 ;
        RECT 9.780 5.550 11.520 9.120 ;
        RECT 9.790 3.830 11.520 5.550 ;
        RECT 19.360 9.120 21.090 9.870 ;
        RECT 19.360 5.550 21.100 9.120 ;
        RECT 23.120 7.480 25.840 9.130 ;
        RECT 23.120 7.440 25.830 7.480 ;
        RECT 23.120 6.110 25.830 6.150 ;
        RECT 19.360 3.830 21.090 5.550 ;
        RECT 23.120 4.460 25.840 6.110 ;
        RECT 26.420 5.730 26.740 6.030 ;
      LAYER li1 ;
        RECT 0.400 9.190 0.600 9.540 ;
        RECT 1.880 9.290 2.410 9.460 ;
        RECT 2.650 9.440 2.840 9.470 ;
        RECT 2.650 9.270 3.710 9.440 ;
        RECT 28.470 9.290 29.000 9.460 ;
        RECT 2.650 9.240 2.840 9.270 ;
        RECT 0.390 9.160 0.600 9.190 ;
        RECT 0.390 8.580 0.610 9.160 ;
        RECT 0.390 8.570 0.600 8.580 ;
        RECT 0.770 8.400 0.960 8.410 ;
        RECT 0.760 8.110 0.960 8.400 ;
        RECT 0.730 7.780 0.970 8.110 ;
        RECT 1.160 7.300 1.330 8.910 ;
        RECT 1.990 7.810 2.160 8.900 ;
        RECT 3.120 8.880 3.310 8.910 ;
        RECT 2.580 8.710 3.310 8.880 ;
        RECT 3.540 8.880 3.710 9.270 ;
        RECT 30.280 9.190 30.480 9.540 ;
        RECT 30.280 9.160 30.490 9.190 ;
        RECT 3.540 8.710 4.280 8.880 ;
        RECT 26.600 8.710 26.950 8.880 ;
        RECT 27.970 8.710 28.300 8.880 ;
        RECT 3.120 8.680 3.310 8.710 ;
        RECT 5.340 8.090 5.570 8.610 ;
        RECT 2.580 7.920 5.570 8.090 ;
        RECT 1.760 7.770 2.160 7.810 ;
        RECT 1.750 7.580 2.160 7.770 ;
        RECT 10.540 7.730 11.090 8.160 ;
        RECT 19.790 7.730 20.340 8.160 ;
        RECT 23.420 7.920 23.650 8.610 ;
        RECT 28.720 8.380 28.890 8.900 ;
        RECT 28.560 8.120 28.890 8.380 ;
        RECT 26.600 7.920 26.950 8.090 ;
        RECT 27.970 7.920 28.300 8.090 ;
        RECT 1.760 7.550 2.160 7.580 ;
        RECT 1.150 7.110 1.330 7.300 ;
        RECT 1.990 7.210 2.160 7.550 ;
        RECT 2.650 7.300 2.840 7.480 ;
        RECT 2.580 7.130 2.930 7.300 ;
        RECT 3.500 6.720 3.710 7.150 ;
        RECT 3.930 7.130 4.270 7.300 ;
        RECT 3.520 6.700 3.690 6.720 ;
        RECT 1.150 6.390 1.330 6.580 ;
        RECT 0.730 5.580 0.970 5.910 ;
        RECT 0.760 5.290 0.960 5.580 ;
        RECT 0.770 5.280 0.960 5.290 ;
        RECT 0.390 5.110 0.600 5.120 ;
        RECT 0.390 4.530 0.610 5.110 ;
        RECT 1.160 4.780 1.330 6.390 ;
        RECT 1.990 6.120 2.160 6.480 ;
        RECT 2.580 6.390 2.930 6.560 ;
        RECT 3.120 6.540 3.310 6.590 ;
        RECT 4.020 6.560 4.190 7.130 ;
        RECT 8.300 6.900 8.490 7.300 ;
        RECT 22.390 6.900 22.580 7.300 ;
        RECT 26.610 7.130 26.950 7.300 ;
        RECT 27.970 7.130 28.300 7.300 ;
        RECT 28.720 7.210 28.890 8.120 ;
        RECT 29.550 7.300 29.720 8.910 ;
        RECT 30.270 8.580 30.490 9.160 ;
        RECT 30.280 8.570 30.490 8.580 ;
        RECT 29.920 8.400 30.110 8.410 ;
        RECT 29.920 8.110 30.120 8.400 ;
        RECT 29.910 7.780 30.150 8.110 ;
        RECT 8.300 6.890 8.680 6.900 ;
        RECT 4.940 6.710 8.680 6.890 ;
        RECT 8.300 6.670 8.680 6.710 ;
        RECT 22.200 6.890 22.580 6.900 ;
        RECT 22.200 6.710 25.940 6.890 ;
        RECT 22.200 6.670 22.580 6.710 ;
        RECT 3.120 6.530 3.350 6.540 ;
        RECT 3.930 6.530 4.270 6.560 ;
        RECT 3.120 6.390 4.270 6.530 ;
        RECT 2.660 6.180 2.850 6.390 ;
        RECT 3.120 6.360 4.100 6.390 ;
        RECT 3.260 6.330 4.100 6.360 ;
        RECT 8.300 6.290 8.490 6.670 ;
        RECT 1.750 6.080 2.160 6.120 ;
        RECT 1.740 5.890 2.160 6.080 ;
        RECT 10.540 6.000 11.090 6.430 ;
        RECT 19.790 6.000 20.340 6.430 ;
        RECT 22.390 6.290 22.580 6.670 ;
        RECT 28.050 6.560 28.220 7.130 ;
        RECT 29.550 7.110 29.730 7.300 ;
        RECT 26.610 6.390 26.950 6.560 ;
        RECT 27.970 6.390 28.300 6.560 ;
        RECT 27.900 6.000 28.070 6.050 ;
        RECT 1.750 5.860 2.160 5.890 ;
        RECT 1.990 4.790 2.160 5.860 ;
        RECT 2.580 5.670 5.510 5.770 ;
        RECT 2.580 5.600 5.570 5.670 ;
        RECT 4.600 5.280 4.770 5.340 ;
        RECT 4.580 5.070 4.790 5.280 ;
        RECT 3.110 4.980 3.300 5.010 ;
        RECT 4.600 5.000 4.770 5.070 ;
        RECT 5.340 4.980 5.570 5.600 ;
        RECT 23.420 4.980 23.650 5.710 ;
        RECT 26.600 5.600 26.950 5.770 ;
        RECT 27.900 5.740 28.460 6.000 ;
        RECT 27.900 5.720 28.300 5.740 ;
        RECT 27.970 5.600 28.300 5.720 ;
        RECT 28.720 5.620 28.890 6.480 ;
        RECT 29.550 6.390 29.730 6.580 ;
        RECT 29.550 5.760 29.720 6.390 ;
        RECT 29.370 5.720 29.720 5.760 ;
        RECT 2.580 4.810 3.300 4.980 ;
        RECT 3.110 4.780 3.300 4.810 ;
        RECT 3.470 4.810 4.280 4.980 ;
        RECT 26.600 4.810 26.950 4.980 ;
        RECT 0.390 4.500 0.600 4.530 ;
        RECT 0.400 4.150 0.600 4.500 ;
        RECT 2.680 4.470 2.870 4.500 ;
        RECT 3.470 4.470 3.660 4.810 ;
        RECT 27.320 4.640 27.500 5.570 ;
        RECT 28.050 5.310 28.380 5.480 ;
        RECT 28.560 5.360 28.890 5.620 ;
        RECT 29.140 5.460 29.720 5.720 ;
        RECT 29.910 5.760 30.150 5.910 ;
        RECT 29.910 5.580 30.510 5.760 ;
        RECT 29.370 5.430 29.720 5.460 ;
        RECT 28.130 5.170 28.380 5.310 ;
        RECT 28.130 4.980 28.610 5.170 ;
        RECT 27.970 4.910 28.610 4.980 ;
        RECT 27.970 4.810 28.300 4.910 ;
        RECT 1.880 4.230 2.410 4.400 ;
        RECT 2.680 4.290 3.660 4.470 ;
        RECT 27.200 4.610 27.520 4.640 ;
        RECT 27.200 4.420 27.530 4.610 ;
        RECT 27.200 4.380 27.520 4.420 ;
        RECT 2.680 4.270 2.870 4.290 ;
        RECT 27.320 0.470 27.500 4.380 ;
        RECT 28.130 3.530 28.300 4.810 ;
        RECT 28.720 4.790 28.890 5.360 ;
        RECT 28.960 5.070 29.130 5.110 ;
        RECT 29.550 5.100 29.720 5.430 ;
        RECT 29.920 5.280 30.510 5.580 ;
        RECT 31.330 5.640 31.910 5.810 ;
        RECT 31.330 5.540 31.720 5.640 ;
        RECT 31.330 5.510 31.710 5.540 ;
        RECT 31.330 5.360 31.690 5.510 ;
        RECT 29.370 5.070 29.720 5.100 ;
        RECT 28.960 4.810 29.720 5.070 ;
        RECT 28.960 4.780 29.130 4.810 ;
        RECT 29.370 4.780 29.720 4.810 ;
        RECT 29.370 4.770 29.570 4.780 ;
        RECT 29.960 4.770 30.510 5.280 ;
        RECT 30.980 5.190 31.690 5.360 ;
        RECT 30.270 4.530 30.490 4.770 ;
        RECT 30.280 4.500 30.490 4.530 ;
        RECT 28.470 4.270 29.000 4.400 ;
        RECT 30.280 4.280 30.480 4.500 ;
        RECT 30.980 4.440 31.680 4.750 ;
        RECT 28.470 4.240 29.130 4.270 ;
        RECT 29.370 4.240 29.570 4.280 ;
        RECT 28.470 4.230 29.570 4.240 ;
        RECT 28.960 3.980 29.570 4.230 ;
        RECT 28.960 3.940 29.130 3.980 ;
        RECT 29.370 3.950 29.570 3.980 ;
        RECT 29.370 3.590 29.570 3.620 ;
        RECT 27.930 3.330 28.250 3.360 ;
        RECT 29.140 3.330 29.570 3.590 ;
        RECT 27.930 3.140 28.260 3.330 ;
        RECT 29.370 3.290 29.570 3.330 ;
        RECT 29.960 3.290 30.510 4.280 ;
        RECT 30.830 4.210 31.680 4.440 ;
        RECT 30.980 3.870 31.680 4.210 ;
        RECT 31.440 3.510 31.760 3.550 ;
        RECT 31.440 3.450 31.770 3.510 ;
        RECT 30.970 3.320 31.770 3.450 ;
        RECT 30.970 3.290 31.760 3.320 ;
        RECT 30.970 3.270 31.670 3.290 ;
        RECT 27.930 3.100 28.250 3.140 ;
        RECT 27.930 3.020 28.100 3.100 ;
        RECT 27.880 2.850 28.100 3.020 ;
        RECT 27.880 2.690 28.050 2.850 ;
        RECT 29.370 2.760 29.570 2.800 ;
        RECT 28.410 2.430 28.600 2.550 ;
        RECT 29.140 2.500 29.570 2.760 ;
        RECT 29.370 2.470 29.570 2.500 ;
        RECT 28.050 2.320 28.600 2.430 ;
        RECT 28.050 2.260 28.590 2.320 ;
        RECT 28.130 0.480 28.300 2.260 ;
        RECT 28.960 2.110 29.130 2.150 ;
        RECT 29.370 2.110 29.570 2.140 ;
        RECT 28.960 1.850 29.570 2.110 ;
        RECT 28.960 1.820 29.130 1.850 ;
        RECT 29.370 1.810 29.570 1.850 ;
        RECT 29.960 1.810 30.510 2.800 ;
        RECT 31.430 2.790 31.750 2.830 ;
        RECT 30.970 2.610 31.760 2.790 ;
        RECT 31.430 2.600 31.760 2.610 ;
        RECT 31.430 2.570 31.750 2.600 ;
        RECT 30.980 1.850 31.680 2.190 ;
        RECT 30.830 1.620 31.680 1.850 ;
        RECT 28.960 1.280 29.130 1.310 ;
        RECT 29.370 1.280 29.570 1.320 ;
        RECT 28.960 1.020 29.570 1.280 ;
        RECT 28.960 0.980 29.130 1.020 ;
        RECT 29.370 0.990 29.570 1.020 ;
        RECT 29.370 0.630 29.570 0.660 ;
        RECT 29.140 0.370 29.570 0.630 ;
        RECT 29.370 0.330 29.570 0.370 ;
        RECT 29.960 0.330 30.510 1.320 ;
        RECT 30.980 1.310 31.680 1.620 ;
        RECT 30.980 0.700 31.690 0.870 ;
        RECT 31.330 0.420 31.690 0.700 ;
        RECT 31.330 0.250 31.910 0.420 ;
      LAYER mcon ;
        RECT 2.230 9.290 2.410 9.460 ;
        RECT 2.660 9.270 2.830 9.440 ;
        RECT 0.420 8.990 0.590 9.160 ;
        RECT 0.770 8.150 0.950 8.340 ;
        RECT 3.130 8.710 3.300 8.880 ;
        RECT 30.290 8.990 30.460 9.160 ;
        RECT 5.370 8.410 5.540 8.580 ;
        RECT 23.450 8.410 23.620 8.580 ;
        RECT 5.370 7.960 5.540 8.130 ;
        RECT 1.850 7.590 2.020 7.760 ;
        RECT 10.820 7.810 11.090 8.080 ;
        RECT 19.790 7.810 20.060 8.080 ;
        RECT 23.450 7.960 23.620 8.130 ;
        RECT 28.620 8.160 28.790 8.330 ;
        RECT 2.660 7.280 2.830 7.450 ;
        RECT 29.930 8.150 30.110 8.340 ;
        RECT 8.500 6.700 8.670 6.870 ;
        RECT 22.210 6.700 22.380 6.870 ;
        RECT 0.770 5.350 0.950 5.540 ;
        RECT 3.130 6.390 3.300 6.560 ;
        RECT 2.670 6.210 2.840 6.380 ;
        RECT 1.840 5.900 2.010 6.070 ;
        RECT 10.820 6.080 11.090 6.350 ;
        RECT 19.790 6.080 20.060 6.350 ;
        RECT 28.230 5.780 28.400 5.950 ;
        RECT 5.370 5.460 5.540 5.630 ;
        RECT 5.370 5.010 5.540 5.180 ;
        RECT 23.450 5.460 23.620 5.630 ;
        RECT 23.450 5.010 23.620 5.180 ;
        RECT 3.120 4.810 3.290 4.980 ;
        RECT 0.420 4.530 0.590 4.700 ;
        RECT 28.620 5.400 28.790 5.570 ;
        RECT 29.200 5.500 29.370 5.670 ;
        RECT 28.380 4.950 28.550 5.120 ;
        RECT 2.230 4.230 2.410 4.400 ;
        RECT 2.690 4.300 2.860 4.470 ;
        RECT 27.260 4.430 27.430 4.600 ;
        RECT 29.930 5.350 30.110 5.540 ;
        RECT 31.450 5.550 31.620 5.720 ;
        RECT 29.150 4.850 29.320 5.020 ;
        RECT 30.180 5.180 30.350 5.350 ;
        RECT 30.290 4.530 30.460 4.700 ;
        RECT 29.150 4.030 29.320 4.200 ;
        RECT 30.840 4.240 31.010 4.410 ;
        RECT 30.180 3.700 30.350 3.870 ;
        RECT 29.200 3.380 29.370 3.550 ;
        RECT 27.990 3.150 28.160 3.320 ;
        RECT 31.500 3.330 31.670 3.500 ;
        RECT 28.420 2.350 28.590 2.520 ;
        RECT 29.200 2.540 29.370 2.710 ;
        RECT 31.490 2.610 31.660 2.780 ;
        RECT 30.180 2.220 30.350 2.390 ;
        RECT 29.150 1.890 29.320 2.060 ;
        RECT 30.840 1.650 31.010 1.820 ;
        RECT 29.150 1.070 29.320 1.240 ;
        RECT 30.180 0.740 30.350 0.910 ;
        RECT 29.200 0.420 29.370 0.590 ;
        RECT 31.410 0.360 31.580 0.530 ;
      LAYER met1 ;
        RECT 0.360 9.220 0.520 9.870 ;
        RECT 0.360 8.670 0.630 9.220 ;
        RECT 0.350 8.620 0.630 8.670 ;
        RECT 0.350 8.530 0.520 8.620 ;
        RECT 0.360 5.160 0.520 8.530 ;
        RECT 0.770 8.410 0.960 9.870 ;
        RECT 2.640 9.500 2.850 9.870 ;
        RECT 2.170 9.050 2.480 9.490 ;
        RECT 2.630 9.210 2.860 9.500 ;
        RECT 0.740 8.380 0.960 8.410 ;
        RECT 0.730 8.110 0.980 8.380 ;
        RECT 0.730 8.100 0.970 8.110 ;
        RECT 0.740 7.860 0.970 8.100 ;
        RECT 0.770 5.830 0.930 7.860 ;
        RECT 1.770 7.520 2.090 7.840 ;
        RECT 2.640 7.510 2.850 9.210 ;
        RECT 3.110 8.940 3.300 9.870 ;
        RECT 3.100 8.650 3.330 8.940 ;
        RECT 1.120 7.010 1.360 7.430 ;
        RECT 2.630 7.220 2.860 7.510 ;
        RECT 2.640 7.080 2.850 7.220 ;
        RECT 1.090 6.690 1.360 7.010 ;
        RECT 1.120 6.260 1.360 6.690 ;
        RECT 3.110 6.620 3.300 8.650 ;
        RECT 3.520 7.150 3.730 9.870 ;
        RECT 5.320 7.870 5.580 8.660 ;
        RECT 3.490 6.640 3.730 7.150 ;
        RECT 2.660 6.440 2.850 6.570 ;
        RECT 2.640 6.150 2.870 6.440 ;
        RECT 3.100 6.330 3.330 6.620 ;
        RECT 1.760 5.830 2.080 6.150 ;
        RECT 0.740 5.590 0.970 5.830 ;
        RECT 0.730 5.580 0.970 5.590 ;
        RECT 0.730 5.310 0.980 5.580 ;
        RECT 0.740 5.280 0.960 5.310 ;
        RECT 0.350 5.070 0.520 5.160 ;
        RECT 0.350 5.020 0.630 5.070 ;
        RECT 0.360 4.470 0.630 5.020 ;
        RECT 0.360 3.820 0.520 4.470 ;
        RECT 0.770 3.820 0.960 5.280 ;
        RECT 2.170 4.200 2.480 4.640 ;
        RECT 2.660 4.530 2.850 6.150 ;
        RECT 3.110 5.040 3.300 6.330 ;
        RECT 3.090 4.750 3.320 5.040 ;
        RECT 2.660 4.320 2.890 4.530 ;
        RECT 2.650 4.240 2.890 4.320 ;
        RECT 2.650 3.820 2.880 4.240 ;
        RECT 3.110 3.820 3.300 4.750 ;
        RECT 3.520 3.820 3.730 6.640 ;
        RECT 4.310 6.030 4.470 6.050 ;
        RECT 4.150 5.730 4.470 6.030 ;
        RECT 5.320 4.930 5.580 5.720 ;
        RECT 10.760 3.820 11.180 9.870 ;
        RECT 19.700 3.820 20.120 9.870 ;
        RECT 22.180 3.820 22.410 9.870 ;
        RECT 23.400 8.660 23.630 9.870 ;
        RECT 28.400 9.050 28.710 9.490 ;
        RECT 23.400 7.870 23.660 8.660 ;
        RECT 28.550 8.090 28.870 8.410 ;
        RECT 23.400 5.720 23.630 7.870 ;
        RECT 29.520 7.300 29.760 7.430 ;
        RECT 29.520 6.980 29.780 7.300 ;
        RECT 23.400 4.930 23.660 5.720 ;
        RECT 28.550 5.330 28.870 5.650 ;
        RECT 31.380 5.480 31.700 5.800 ;
        RECT 23.400 3.820 23.630 4.930 ;
        RECT 28.300 4.880 28.620 5.200 ;
        RECT 27.190 4.350 27.510 4.670 ;
        RECT 27.920 3.070 28.240 3.390 ;
        RECT 29.130 3.300 29.450 3.620 ;
        RECT 31.430 3.260 31.750 3.580 ;
        RECT 29.130 2.470 29.450 2.790 ;
        RECT 31.420 2.540 31.740 2.860 ;
        RECT 29.080 1.820 29.400 2.140 ;
        RECT 29.080 0.990 29.400 1.310 ;
        RECT 12.370 0.050 12.690 0.350 ;
        RECT 18.170 0.050 18.490 0.350 ;
        RECT 29.130 0.340 29.450 0.660 ;
        RECT 31.340 0.290 31.660 0.610 ;
      LAYER via ;
        RECT 2.190 9.080 2.450 9.340 ;
        RECT 1.800 7.550 2.060 7.810 ;
        RECT 1.090 6.720 1.350 6.980 ;
        RECT 1.790 5.860 2.050 6.120 ;
        RECT 2.190 4.350 2.450 4.610 ;
        RECT 4.180 5.750 4.440 6.010 ;
        RECT 28.430 9.080 28.690 9.340 ;
        RECT 28.580 8.120 28.840 8.380 ;
        RECT 29.520 7.010 29.780 7.270 ;
        RECT 28.580 5.360 28.840 5.620 ;
        RECT 31.410 5.510 31.670 5.770 ;
        RECT 28.330 4.910 28.590 5.170 ;
        RECT 27.220 4.380 27.480 4.640 ;
        RECT 27.950 3.100 28.210 3.360 ;
        RECT 29.160 3.330 29.420 3.590 ;
        RECT 31.460 3.290 31.720 3.550 ;
        RECT 29.160 2.500 29.420 2.760 ;
        RECT 31.450 2.570 31.710 2.830 ;
        RECT 29.110 1.850 29.370 2.110 ;
        RECT 29.110 1.020 29.370 1.280 ;
        RECT 29.160 0.370 29.420 0.630 ;
        RECT 12.400 0.070 12.660 0.330 ;
        RECT 18.200 0.070 18.460 0.330 ;
        RECT 31.370 0.320 31.630 0.580 ;
      LAYER met2 ;
        RECT 2.410 9.380 2.730 9.390 ;
        RECT 2.170 9.370 2.730 9.380 ;
        RECT 28.400 9.370 28.710 9.380 ;
        RECT 0.000 9.190 11.520 9.370 ;
        RECT 19.350 9.190 30.880 9.370 ;
        RECT 2.170 9.050 2.480 9.190 ;
        RECT 28.400 9.050 28.710 9.190 ;
        RECT 28.550 8.350 28.860 8.420 ;
        RECT 28.550 8.130 30.880 8.350 ;
        RECT 28.550 8.090 28.860 8.130 ;
        RECT 1.780 7.830 2.090 7.850 ;
        RECT 1.780 7.640 11.520 7.830 ;
        RECT 1.780 7.520 2.090 7.640 ;
        RECT 1.060 6.950 1.380 6.980 ;
        RECT 1.060 6.720 11.520 6.950 ;
        RECT 2.170 4.500 2.480 4.640 ;
        RECT 0.000 4.490 2.480 4.500 ;
        RECT 0.000 4.340 11.520 4.490 ;
        RECT 0.000 4.320 2.480 4.340 ;
        RECT 2.170 4.310 2.480 4.320 ;
        RECT 15.460 3.820 23.450 4.020 ;
        RECT 22.050 3.140 22.270 3.150 ;
        RECT 15.470 2.890 22.300 3.140 ;
        RECT 23.230 3.100 23.450 3.820 ;
        RECT 15.470 1.970 18.980 2.160 ;
        RECT 18.750 1.370 18.980 1.970 ;
        RECT 22.010 1.720 22.300 2.890 ;
        RECT 23.200 3.060 23.450 3.100 ;
        RECT 23.200 2.420 23.460 3.060 ;
        RECT 23.200 2.210 27.330 2.420 ;
        RECT 27.120 2.070 27.330 2.210 ;
        RECT 29.080 2.070 29.390 2.150 ;
        RECT 27.120 1.860 29.390 2.070 ;
        RECT 29.080 1.820 29.390 1.860 ;
        RECT 22.010 1.500 24.900 1.720 ;
        RECT 22.010 1.490 22.300 1.500 ;
        RECT 18.750 1.220 18.970 1.370 ;
        RECT 29.080 1.270 29.390 1.310 ;
        RECT 23.120 1.220 29.390 1.270 ;
        RECT 18.750 1.060 29.390 1.220 ;
        RECT 18.750 1.000 23.510 1.060 ;
        RECT 29.080 0.980 29.390 1.060 ;
        RECT 29.130 0.580 29.440 0.660 ;
        RECT 31.340 0.580 31.650 0.620 ;
        RECT 29.130 0.350 31.840 0.580 ;
        RECT 29.130 0.330 29.440 0.350 ;
        RECT 31.340 0.290 31.650 0.350 ;
  END
END sky130_hilas_TA2Cell_1FG_Strong

MACRO sky130_hilas_TA2Cell_NoFG
  CLASS CORE ;
  FOREIGN sky130_hilas_TA2Cell_NoFG ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 9.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN COLSEL1
    PORT
      LAYER met1 ;
        RECT 10.570 5.970 10.760 6.050 ;
    END
  END COLSEL1
  PIN VIN12
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT 12.470 0.270 12.780 0.340 ;
        RECT 11.870 0.020 12.780 0.270 ;
        RECT 12.470 0.010 12.780 0.020 ;
    END
  END VIN12
  PIN VIN21
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT 13.790 3.350 14.100 3.390 ;
        RECT 13.700 3.340 14.130 3.350 ;
        RECT 13.470 3.110 14.570 3.340 ;
        RECT 13.790 3.060 14.100 3.110 ;
    END
  END VIN21
  PIN VIN22
    ANTENNAGATEAREA 4.299400 ;
    ANTENNADIFFAREA 6.715500 ;
    PORT
      LAYER nwell ;
        RECT 12.180 6.050 15.490 9.870 ;
        RECT 11.220 3.830 15.490 6.050 ;
        RECT 11.220 0.010 14.640 3.830 ;
        RECT 12.780 0.000 14.640 0.010 ;
      LAYER met2 ;
        RECT 14.100 7.010 14.420 7.270 ;
        RECT 14.140 6.990 15.320 7.010 ;
        RECT 14.140 6.730 15.360 6.990 ;
        RECT 14.140 6.670 15.320 6.730 ;
        RECT 14.100 6.660 15.320 6.670 ;
        RECT 14.100 6.410 14.420 6.660 ;
        RECT 13.430 6.030 13.680 6.040 ;
        RECT 14.030 6.030 14.340 6.040 ;
        RECT 13.430 5.780 14.340 6.030 ;
        RECT 14.030 5.710 14.340 5.780 ;
        RECT 15.000 5.710 15.310 5.760 ;
        RECT 17.250 5.710 17.560 5.810 ;
        RECT 13.160 5.590 13.470 5.660 ;
        RECT 15.000 5.590 17.560 5.710 ;
        RECT 13.160 5.480 17.560 5.590 ;
        RECT 13.160 5.380 15.490 5.480 ;
        RECT 13.160 5.330 13.470 5.380 ;
        RECT 14.180 5.170 14.490 5.210 ;
        RECT 14.000 5.030 14.740 5.170 ;
        RECT 14.950 5.030 15.260 5.110 ;
        RECT 14.000 4.920 15.260 5.030 ;
        RECT 14.180 4.880 15.260 4.920 ;
        RECT 14.490 4.820 15.260 4.880 ;
        RECT 14.490 4.800 14.740 4.820 ;
        RECT 14.950 4.780 15.260 4.820 ;
        RECT 13.060 4.640 13.370 4.670 ;
        RECT 13.010 4.530 13.370 4.640 ;
        RECT 15.960 4.600 16.300 4.690 ;
        RECT 11.450 4.500 13.370 4.530 ;
        RECT 13.610 4.500 16.300 4.600 ;
        RECT 11.450 4.490 16.300 4.500 ;
        RECT 3.960 4.410 16.300 4.490 ;
        RECT 3.960 4.340 15.490 4.410 ;
        RECT 15.960 4.360 16.300 4.410 ;
        RECT 11.450 4.320 15.490 4.340 ;
        RECT 11.450 4.310 13.320 4.320 ;
        RECT 13.610 3.840 13.800 4.320 ;
        RECT 14.520 4.230 14.730 4.240 ;
        RECT 14.950 4.230 15.260 4.270 ;
        RECT 14.520 4.160 15.260 4.230 ;
        RECT 14.230 4.140 15.260 4.160 ;
        RECT 14.180 4.020 15.260 4.140 ;
        RECT 14.180 3.950 14.730 4.020 ;
        RECT 14.180 3.890 14.650 3.950 ;
        RECT 14.950 3.940 15.260 4.020 ;
        RECT 2.820 3.650 13.800 3.840 ;
        RECT 2.820 3.470 3.010 3.650 ;
        RECT 2.800 2.480 3.150 3.470 ;
        RECT 12.230 2.940 12.540 2.990 ;
        RECT 11.910 2.710 13.010 2.940 ;
        RECT 11.910 2.700 12.570 2.710 ;
        RECT 12.230 2.660 12.540 2.700 ;
    END
  END VIN22
  PIN OUTPUT1
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER met2 ;
        RECT 15.000 2.740 15.310 2.800 ;
        RECT 17.290 2.740 17.600 2.870 ;
        RECT 15.000 2.520 17.920 2.740 ;
        RECT 15.000 2.470 15.310 2.520 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER met2 ;
        RECT 15.000 3.570 15.310 3.620 ;
        RECT 17.300 3.570 17.610 3.590 ;
        RECT 15.000 3.340 17.920 3.570 ;
        RECT 15.000 3.290 15.310 3.340 ;
        RECT 17.300 3.260 17.610 3.340 ;
    END
  END OUTPUT2
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 15.960 0.000 16.300 6.050 ;
      LAYER via ;
        RECT 16.000 4.390 16.260 4.650 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 16.650 5.870 17.920 6.050 ;
        RECT 16.640 0.000 17.920 5.870 ;
      LAYER met1 ;
        RECT 16.630 4.470 16.900 6.050 ;
        RECT 16.630 4.180 16.910 4.470 ;
        RECT 16.630 1.880 16.900 4.180 ;
        RECT 16.630 1.590 16.910 1.880 ;
        RECT 16.630 0.000 16.900 1.590 ;
    END
  END VPWR
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 0.000 5.370 0.070 5.550 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 0.000 0.520 0.080 0.670 ;
    END
  END DRAIN2
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 0.350 5.980 0.770 6.050 ;
    END
  END VTUN
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT 4.050 5.970 4.280 6.050 ;
    END
  END GATE1
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 11.010 5.970 11.290 6.050 ;
    END
  END VINJ
  OBS
      LAYER nwell ;
        RECT 3.970 9.120 5.700 9.870 ;
        RECT 3.970 5.550 5.710 9.120 ;
        RECT 7.730 7.480 10.450 9.130 ;
        RECT 7.730 7.440 10.440 7.480 ;
        RECT 7.730 6.110 10.440 6.150 ;
        RECT 3.970 3.830 5.700 5.550 ;
        RECT 7.730 4.460 10.450 6.110 ;
      LAYER li1 ;
        RECT 13.080 9.290 13.610 9.460 ;
        RECT 14.890 9.190 15.090 9.540 ;
        RECT 14.890 9.160 15.100 9.190 ;
        RECT 11.210 8.710 11.560 8.880 ;
        RECT 12.580 8.710 12.910 8.880 ;
        RECT 4.400 7.730 4.950 8.160 ;
        RECT 8.030 7.920 8.260 8.610 ;
        RECT 13.330 8.380 13.500 8.900 ;
        RECT 13.170 8.120 13.500 8.380 ;
        RECT 11.210 7.920 11.560 8.090 ;
        RECT 12.580 7.920 12.910 8.090 ;
        RECT 7.000 6.900 7.190 7.300 ;
        RECT 11.220 7.130 11.560 7.300 ;
        RECT 12.580 7.130 12.910 7.300 ;
        RECT 13.330 7.210 13.500 8.120 ;
        RECT 14.160 7.300 14.330 8.910 ;
        RECT 14.880 8.580 15.100 9.160 ;
        RECT 14.890 8.570 15.100 8.580 ;
        RECT 14.530 8.400 14.720 8.410 ;
        RECT 14.530 8.110 14.730 8.400 ;
        RECT 14.520 7.780 14.760 8.110 ;
        RECT 6.810 6.890 7.190 6.900 ;
        RECT 6.810 6.710 10.550 6.890 ;
        RECT 6.810 6.670 7.190 6.710 ;
        RECT 4.400 6.000 4.950 6.430 ;
        RECT 7.000 6.290 7.190 6.670 ;
        RECT 12.660 6.560 12.830 7.130 ;
        RECT 14.160 7.110 14.340 7.300 ;
        RECT 11.220 6.390 11.560 6.560 ;
        RECT 12.580 6.390 12.910 6.560 ;
        RECT 8.030 4.980 8.260 5.710 ;
        RECT 11.210 5.600 11.560 5.770 ;
        RECT 12.580 5.600 12.910 5.770 ;
        RECT 13.330 5.620 13.500 6.480 ;
        RECT 14.160 6.390 14.340 6.580 ;
        RECT 13.770 6.000 13.940 6.050 ;
        RECT 14.160 6.000 14.330 6.390 ;
        RECT 13.770 5.740 14.330 6.000 ;
        RECT 13.770 5.720 13.940 5.740 ;
        RECT 11.210 4.810 11.560 4.980 ;
        RECT 2.830 2.470 3.290 3.480 ;
        RECT 11.630 1.670 11.810 5.580 ;
        RECT 12.440 4.980 12.610 5.570 ;
        RECT 13.170 5.360 13.500 5.620 ;
        RECT 14.160 5.480 14.330 5.740 ;
        RECT 14.520 5.580 14.760 5.910 ;
        RECT 15.240 5.720 15.440 5.760 ;
        RECT 12.440 4.810 12.910 4.980 ;
        RECT 12.440 3.790 12.610 4.810 ;
        RECT 13.190 4.790 13.500 5.360 ;
        RECT 13.920 5.310 14.330 5.480 ;
        RECT 14.000 5.170 14.330 5.310 ;
        RECT 14.530 5.290 14.730 5.580 ;
        RECT 15.010 5.460 15.440 5.720 ;
        RECT 15.240 5.430 15.440 5.460 ;
        RECT 14.530 5.280 14.720 5.290 ;
        RECT 14.000 4.910 14.480 5.170 ;
        RECT 14.890 5.110 15.100 5.120 ;
        RECT 14.830 5.070 15.100 5.110 ;
        RECT 15.240 5.070 15.440 5.100 ;
        RECT 13.190 4.640 13.370 4.790 ;
        RECT 14.000 4.780 14.330 4.910 ;
        RECT 14.830 4.810 15.440 5.070 ;
        RECT 14.830 4.780 15.100 4.810 ;
        RECT 13.070 4.610 13.390 4.640 ;
        RECT 13.070 4.420 13.400 4.610 ;
        RECT 13.070 4.400 13.390 4.420 ;
        RECT 13.070 4.380 13.610 4.400 ;
        RECT 13.080 4.230 13.610 4.380 ;
        RECT 12.360 3.730 12.900 3.790 ;
        RECT 12.360 3.620 12.910 3.730 ;
        RECT 12.720 3.500 12.910 3.620 ;
        RECT 12.190 3.200 12.360 3.360 ;
        RECT 12.190 3.030 12.410 3.200 ;
        RECT 12.240 2.950 12.410 3.030 ;
        RECT 12.240 2.910 12.560 2.950 ;
        RECT 12.240 2.720 12.570 2.910 ;
        RECT 12.240 2.690 12.560 2.720 ;
        RECT 11.510 1.630 11.830 1.670 ;
        RECT 11.510 1.440 11.840 1.630 ;
        RECT 11.510 1.410 11.830 1.440 ;
        RECT 11.630 0.480 11.810 1.410 ;
        RECT 12.440 1.140 12.610 2.520 ;
        RECT 12.440 0.880 12.920 1.140 ;
        RECT 12.440 0.740 12.690 0.880 ;
        RECT 12.360 0.570 12.690 0.740 ;
        RECT 13.190 0.470 13.370 4.230 ;
        RECT 14.000 3.530 14.170 4.780 ;
        RECT 14.880 4.530 15.100 4.780 ;
        RECT 15.240 4.770 15.440 4.810 ;
        RECT 15.830 4.770 16.380 5.760 ;
        RECT 17.200 5.640 17.780 5.810 ;
        RECT 17.200 5.540 17.590 5.640 ;
        RECT 17.200 5.510 17.580 5.540 ;
        RECT 17.200 5.360 17.560 5.510 ;
        RECT 16.850 5.190 17.560 5.360 ;
        RECT 14.890 4.500 15.100 4.530 ;
        RECT 14.890 4.270 15.090 4.500 ;
        RECT 16.850 4.440 17.550 4.750 ;
        RECT 14.830 4.240 15.090 4.270 ;
        RECT 15.240 4.240 15.440 4.280 ;
        RECT 14.830 3.980 15.440 4.240 ;
        RECT 14.830 3.940 15.000 3.980 ;
        RECT 15.240 3.950 15.440 3.980 ;
        RECT 15.240 3.590 15.440 3.620 ;
        RECT 13.800 3.330 14.120 3.360 ;
        RECT 15.010 3.330 15.440 3.590 ;
        RECT 13.800 3.140 14.130 3.330 ;
        RECT 15.240 3.290 15.440 3.330 ;
        RECT 15.830 3.290 16.380 4.280 ;
        RECT 16.700 4.210 17.550 4.440 ;
        RECT 16.850 3.870 17.550 4.210 ;
        RECT 17.310 3.510 17.630 3.550 ;
        RECT 17.310 3.450 17.640 3.510 ;
        RECT 16.840 3.320 17.640 3.450 ;
        RECT 16.840 3.290 17.630 3.320 ;
        RECT 16.840 3.270 17.540 3.290 ;
        RECT 13.800 3.100 14.120 3.140 ;
        RECT 13.800 3.020 13.970 3.100 ;
        RECT 13.750 2.850 13.970 3.020 ;
        RECT 13.750 2.690 13.920 2.850 ;
        RECT 15.240 2.760 15.440 2.800 ;
        RECT 14.280 2.430 14.470 2.550 ;
        RECT 15.010 2.500 15.440 2.760 ;
        RECT 15.240 2.470 15.440 2.500 ;
        RECT 13.920 2.320 14.470 2.430 ;
        RECT 13.920 2.260 14.460 2.320 ;
        RECT 14.000 0.480 14.170 2.260 ;
        RECT 14.830 2.110 15.000 2.150 ;
        RECT 15.240 2.110 15.440 2.140 ;
        RECT 14.830 1.850 15.440 2.110 ;
        RECT 14.830 1.820 15.000 1.850 ;
        RECT 15.240 1.810 15.440 1.850 ;
        RECT 15.830 1.810 16.380 2.800 ;
        RECT 17.300 2.790 17.620 2.830 ;
        RECT 16.840 2.610 17.630 2.790 ;
        RECT 17.300 2.600 17.630 2.610 ;
        RECT 17.300 2.570 17.620 2.600 ;
        RECT 16.850 1.850 17.550 2.190 ;
        RECT 16.700 1.620 17.550 1.850 ;
        RECT 14.830 1.280 15.000 1.310 ;
        RECT 15.240 1.280 15.440 1.320 ;
        RECT 14.830 1.020 15.440 1.280 ;
        RECT 14.830 0.980 15.000 1.020 ;
        RECT 15.240 0.990 15.440 1.020 ;
        RECT 15.240 0.630 15.440 0.660 ;
        RECT 15.010 0.370 15.440 0.630 ;
        RECT 15.240 0.330 15.440 0.370 ;
        RECT 15.830 0.330 16.380 1.320 ;
        RECT 16.850 1.310 17.550 1.620 ;
        RECT 16.850 0.700 17.560 0.870 ;
        RECT 17.200 0.420 17.560 0.700 ;
        RECT 12.210 0.310 12.380 0.330 ;
        RECT 12.210 0.050 12.770 0.310 ;
        RECT 17.200 0.250 17.780 0.420 ;
        RECT 12.210 0.000 12.380 0.050 ;
      LAYER mcon ;
        RECT 14.900 8.990 15.070 9.160 ;
        RECT 8.060 8.410 8.230 8.580 ;
        RECT 4.400 7.810 4.670 8.080 ;
        RECT 8.060 7.960 8.230 8.130 ;
        RECT 13.230 8.160 13.400 8.330 ;
        RECT 14.540 8.150 14.720 8.340 ;
        RECT 6.820 6.700 6.990 6.870 ;
        RECT 4.400 6.080 4.670 6.350 ;
        RECT 8.060 5.460 8.230 5.630 ;
        RECT 14.100 5.780 14.270 5.950 ;
        RECT 8.060 5.010 8.230 5.180 ;
        RECT 2.860 3.220 3.030 3.390 ;
        RECT 2.860 2.530 3.030 2.700 ;
        RECT 13.230 5.400 13.400 5.570 ;
        RECT 14.540 5.350 14.720 5.540 ;
        RECT 15.070 5.500 15.240 5.670 ;
        RECT 17.320 5.550 17.490 5.720 ;
        RECT 16.050 5.180 16.220 5.350 ;
        RECT 14.250 4.950 14.420 5.120 ;
        RECT 15.020 4.850 15.190 5.020 ;
        RECT 13.130 4.430 13.300 4.600 ;
        RECT 12.730 3.530 12.900 3.700 ;
        RECT 12.300 2.730 12.470 2.900 ;
        RECT 11.570 1.450 11.740 1.620 ;
        RECT 12.690 0.930 12.860 1.100 ;
        RECT 14.900 4.530 15.070 4.700 ;
        RECT 15.020 4.030 15.190 4.200 ;
        RECT 16.710 4.240 16.880 4.410 ;
        RECT 16.050 3.700 16.220 3.870 ;
        RECT 15.070 3.380 15.240 3.550 ;
        RECT 13.860 3.150 14.030 3.320 ;
        RECT 17.370 3.330 17.540 3.500 ;
        RECT 14.290 2.350 14.460 2.520 ;
        RECT 15.070 2.540 15.240 2.710 ;
        RECT 17.360 2.610 17.530 2.780 ;
        RECT 16.050 2.220 16.220 2.390 ;
        RECT 15.020 1.890 15.190 2.060 ;
        RECT 16.710 1.650 16.880 1.820 ;
        RECT 15.020 1.070 15.190 1.240 ;
        RECT 16.050 0.740 16.220 0.910 ;
        RECT 15.070 0.420 15.240 0.590 ;
        RECT 17.280 0.360 17.450 0.530 ;
        RECT 12.540 0.100 12.710 0.270 ;
      LAYER met1 ;
        RECT 4.310 3.820 4.730 9.870 ;
        RECT 6.790 3.820 7.020 9.870 ;
        RECT 8.010 8.660 8.240 9.870 ;
        RECT 13.010 9.050 13.320 9.490 ;
        RECT 8.010 7.870 8.270 8.660 ;
        RECT 14.530 8.410 14.720 9.870 ;
        RECT 14.970 9.220 15.250 9.870 ;
        RECT 14.860 8.620 15.250 9.220 ;
        RECT 13.160 8.090 13.480 8.410 ;
        RECT 14.530 8.380 14.750 8.410 ;
        RECT 14.510 8.110 14.760 8.380 ;
        RECT 14.520 8.100 14.760 8.110 ;
        RECT 8.010 5.720 8.240 7.870 ;
        RECT 14.520 7.860 14.750 8.100 ;
        RECT 14.130 7.300 14.370 7.430 ;
        RECT 14.130 6.980 14.390 7.300 ;
        RECT 14.130 6.380 14.390 6.700 ;
        RECT 14.130 6.260 14.370 6.380 ;
        RECT 8.010 4.930 8.270 5.720 ;
        RECT 14.020 5.710 14.340 6.030 ;
        RECT 14.560 5.830 14.720 7.860 ;
        RECT 14.970 7.020 15.250 8.620 ;
        RECT 14.970 6.700 15.330 7.020 ;
        RECT 13.160 5.330 13.480 5.650 ;
        RECT 14.520 5.590 14.750 5.830 ;
        RECT 14.970 5.750 15.250 6.700 ;
        RECT 14.520 5.580 14.760 5.590 ;
        RECT 14.510 5.310 14.760 5.580 ;
        RECT 14.970 5.430 15.320 5.750 ;
        RECT 17.250 5.480 17.570 5.800 ;
        RECT 14.530 5.280 14.750 5.310 ;
        RECT 8.010 3.820 8.240 4.930 ;
        RECT 14.170 4.880 14.490 5.200 ;
        RECT 13.060 4.640 13.380 4.670 ;
        RECT 13.010 4.350 13.380 4.640 ;
        RECT 13.010 4.200 13.320 4.350 ;
        RECT 14.280 4.190 14.490 4.300 ;
        RECT 14.260 3.870 14.520 4.190 ;
        RECT 2.790 2.470 3.170 3.480 ;
        RECT 12.700 3.470 12.930 3.760 ;
        RECT 12.230 2.660 12.550 2.980 ;
        RECT 12.720 2.180 12.930 3.470 ;
        RECT 13.790 3.070 14.110 3.390 ;
        RECT 14.280 2.580 14.490 3.870 ;
        RECT 14.530 3.820 14.720 5.280 ;
        RECT 14.970 5.100 15.250 5.430 ;
        RECT 14.950 5.070 15.270 5.100 ;
        RECT 14.860 4.780 15.270 5.070 ;
        RECT 14.860 4.470 15.250 4.780 ;
        RECT 14.970 4.270 15.250 4.470 ;
        RECT 14.950 3.950 15.270 4.270 ;
        RECT 14.970 3.820 15.250 3.950 ;
        RECT 15.000 3.300 15.320 3.620 ;
        RECT 17.300 3.260 17.620 3.580 ;
        RECT 14.260 2.290 14.490 2.580 ;
        RECT 15.000 2.470 15.320 2.790 ;
        RECT 17.290 2.540 17.610 2.860 ;
        RECT 12.700 1.860 12.960 2.180 ;
        RECT 12.720 1.750 12.930 1.860 ;
        RECT 14.950 1.820 15.270 2.140 ;
        RECT 11.500 1.380 11.820 1.700 ;
        RECT 12.610 0.850 12.930 1.170 ;
        RECT 14.950 0.990 15.270 1.310 ;
        RECT 15.000 0.340 15.320 0.660 ;
        RECT 12.460 0.020 12.780 0.340 ;
        RECT 17.210 0.290 17.530 0.610 ;
      LAYER via ;
        RECT 13.040 9.080 13.300 9.340 ;
        RECT 13.190 8.120 13.450 8.380 ;
        RECT 14.130 7.010 14.390 7.270 ;
        RECT 14.130 6.410 14.390 6.670 ;
        RECT 14.050 5.740 14.310 6.000 ;
        RECT 15.070 6.730 15.330 6.990 ;
        RECT 13.190 5.360 13.450 5.620 ;
        RECT 15.030 5.460 15.290 5.720 ;
        RECT 17.280 5.510 17.540 5.770 ;
        RECT 14.200 4.910 14.460 5.170 ;
        RECT 13.090 4.610 13.350 4.640 ;
        RECT 13.040 4.380 13.350 4.610 ;
        RECT 13.040 4.350 13.300 4.380 ;
        RECT 14.260 3.900 14.520 4.160 ;
        RECT 2.830 2.510 3.120 3.440 ;
        RECT 12.260 2.690 12.520 2.950 ;
        RECT 13.820 3.100 14.080 3.360 ;
        RECT 14.980 4.810 15.240 5.070 ;
        RECT 14.980 3.980 15.240 4.240 ;
        RECT 15.030 3.330 15.290 3.590 ;
        RECT 17.330 3.290 17.590 3.550 ;
        RECT 15.030 2.500 15.290 2.760 ;
        RECT 17.320 2.570 17.580 2.830 ;
        RECT 12.700 1.890 12.960 2.150 ;
        RECT 14.980 1.850 15.240 2.110 ;
        RECT 11.530 1.410 11.790 1.670 ;
        RECT 12.640 0.880 12.900 1.140 ;
        RECT 14.980 1.020 15.240 1.280 ;
        RECT 15.030 0.370 15.290 0.630 ;
        RECT 12.490 0.050 12.750 0.310 ;
        RECT 17.240 0.320 17.500 0.580 ;
      LAYER met2 ;
        RECT 13.010 9.370 13.320 9.380 ;
        RECT 3.960 9.190 15.490 9.370 ;
        RECT 13.010 9.050 13.320 9.190 ;
        RECT 13.160 8.350 13.470 8.420 ;
        RECT 13.160 8.130 15.490 8.350 ;
        RECT 13.160 8.090 13.470 8.130 ;
        RECT 12.620 2.070 13.090 2.160 ;
        RECT 14.950 2.070 15.260 2.150 ;
        RECT 12.620 1.910 15.260 2.070 ;
        RECT 12.670 1.890 15.260 1.910 ;
        RECT 12.960 1.870 15.260 1.890 ;
        RECT 14.650 1.860 15.260 1.870 ;
        RECT 14.950 1.820 15.260 1.860 ;
        RECT 11.390 1.710 11.550 1.780 ;
        RECT 11.390 1.380 11.810 1.710 ;
        RECT 14.950 1.270 15.260 1.310 ;
        RECT 12.670 1.170 15.260 1.270 ;
        RECT 12.620 1.130 15.260 1.170 ;
        RECT 12.440 1.060 15.260 1.130 ;
        RECT 12.440 0.880 12.990 1.060 ;
        RECT 14.950 0.980 15.260 1.060 ;
        RECT 12.620 0.840 12.930 0.880 ;
        RECT 15.000 0.580 15.310 0.660 ;
        RECT 17.210 0.580 17.520 0.620 ;
        RECT 15.000 0.350 17.710 0.580 ;
        RECT 15.000 0.330 15.310 0.350 ;
        RECT 17.210 0.290 17.520 0.350 ;
  END
END sky130_hilas_TA2Cell_NoFG

MACRO sky130_hilas_TopLevelTextStructure
  CLASS CORE ;
  FOREIGN sky130_hilas_TopLevelTextStructure ;
  ORIGIN 0.000 0.000 ;
  SIZE 130.250 BY 78.160 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DIG24 
    ANTENNAGATEAREA 0.236000 ;
    ANTENNADIFFAREA 4.378700 ;
    PORT
      LAYER nwell ;
        RECT 66.090 38.200 68.640 38.210 ;
        RECT 66.080 34.390 68.640 38.200 ;
        RECT 70.170 34.390 72.400 38.210 ;
        RECT 66.080 34.380 72.400 34.390 ;
        RECT 66.080 34.230 68.750 34.380 ;
        RECT 66.080 34.220 68.930 34.230 ;
        RECT 66.080 32.180 68.750 34.220 ;
        RECT 66.090 32.170 68.750 32.180 ;
        RECT 68.230 31.310 68.750 32.170 ;
        RECT 70.170 32.160 72.400 34.380 ;
        RECT 68.340 28.350 68.750 31.310 ;
      LAYER met2 ;
        RECT 68.240 34.270 68.550 34.290 ;
        RECT 66.080 34.110 76.150 34.270 ;
        RECT 66.080 34.100 76.140 34.110 ;
        RECT 66.080 34.090 68.640 34.100 ;
        RECT 68.240 33.960 68.550 34.090 ;
        RECT 71.500 34.080 71.820 34.100 ;
        RECT 71.500 33.890 79.420 34.080 ;
        RECT 79.580 33.890 79.890 33.930 ;
        RECT 71.500 33.870 79.890 33.890 ;
        RECT 71.500 33.840 71.820 33.870 ;
        RECT 79.210 33.680 79.890 33.870 ;
        RECT 79.580 33.600 79.890 33.680 ;
        RECT 68.230 33.410 68.380 33.460 ;
        RECT 68.230 33.290 68.550 33.410 ;
        RECT 68.230 33.280 76.150 33.290 ;
        RECT 66.080 33.120 76.150 33.280 ;
        RECT 66.080 33.100 68.640 33.120 ;
        RECT 68.230 33.080 68.550 33.100 ;
        RECT 68.230 32.950 68.380 33.080 ;
        RECT 71.480 32.950 71.800 33.050 ;
        RECT 73.820 33.030 75.360 33.120 ;
        RECT 68.230 32.850 71.800 32.950 ;
        RECT 66.080 32.790 71.800 32.850 ;
        RECT 66.080 32.760 68.650 32.790 ;
        RECT 73.730 32.760 74.050 32.810 ;
        RECT 66.080 32.670 74.050 32.760 ;
        RECT 67.660 32.600 74.050 32.670 ;
        RECT 68.240 32.550 68.550 32.600 ;
        RECT 73.730 32.550 74.050 32.600 ;
        RECT 68.210 32.530 68.550 32.550 ;
        RECT 68.210 32.290 68.530 32.530 ;
        RECT 68.280 32.280 68.450 32.290 ;
        RECT 73.210 31.830 73.530 31.880 ;
        RECT 67.670 31.810 73.530 31.830 ;
        RECT 67.670 31.780 79.010 31.810 ;
        RECT 67.670 31.670 79.070 31.780 ;
        RECT 71.440 31.610 79.070 31.670 ;
        RECT 79.580 31.610 79.890 31.690 ;
        RECT 68.190 31.510 68.510 31.540 ;
        RECT 71.440 31.510 71.680 31.610 ;
        RECT 68.190 31.330 71.680 31.510 ;
        RECT 78.880 31.410 79.890 31.610 ;
        RECT 79.480 31.400 79.890 31.410 ;
        RECT 79.580 31.360 79.890 31.400 ;
        RECT 68.190 31.310 71.600 31.330 ;
        RECT 68.190 31.280 68.510 31.310 ;
        RECT 73.710 23.600 129.540 23.640 ;
        RECT 73.710 23.140 130.250 23.600 ;
        RECT 124.150 22.740 126.160 22.760 ;
        RECT 73.170 22.240 126.160 22.740 ;
        RECT 124.150 3.120 126.160 22.240 ;
        RECT 128.240 3.140 130.250 23.140 ;
        RECT 124.150 2.470 126.190 3.120 ;
        RECT 128.210 2.560 130.250 3.140 ;
        RECT 128.210 2.490 130.240 2.560 ;
        RECT 124.150 2.390 126.160 2.470 ;
    END
  END DIG24 
  PIN DIG22
    ANTENNAGATEAREA 0.118000 ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 71.480 31.130 71.800 31.170 ;
        RECT 71.480 31.110 79.030 31.130 ;
        RECT 79.580 31.120 79.890 31.160 ;
        RECT 79.480 31.110 79.890 31.120 ;
        RECT 71.480 30.910 79.890 31.110 ;
        RECT 71.580 30.900 71.900 30.910 ;
        RECT 79.580 30.830 79.890 30.910 ;
        RECT 68.170 29.990 68.370 30.450 ;
        RECT 72.740 29.990 73.060 30.040 ;
        RECT 67.660 29.830 73.060 29.990 ;
        RECT 68.170 29.750 71.720 29.830 ;
        RECT 72.740 29.780 73.060 29.830 ;
        RECT 71.320 29.730 71.640 29.750 ;
        RECT 72.700 21.820 121.970 21.840 ;
        RECT 72.700 21.340 122.080 21.820 ;
        RECT 120.070 3.140 122.080 21.340 ;
        RECT 120.070 2.490 122.140 3.140 ;
        RECT 120.070 2.450 122.080 2.490 ;
    END
  END DIG22
  PIN DIG21
    ANTENNAGATEAREA 0.118000 ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 68.140 29.210 68.450 29.540 ;
        RECT 72.240 29.060 72.560 29.110 ;
        RECT 67.720 28.900 72.560 29.060 ;
        RECT 68.210 28.850 68.740 28.900 ;
        RECT 72.240 28.850 72.560 28.900 ;
        RECT 79.580 28.860 79.890 28.920 ;
        RECT 79.030 28.850 79.890 28.860 ;
        RECT 68.190 28.570 68.500 28.690 ;
        RECT 71.450 28.630 79.890 28.850 ;
        RECT 71.450 28.620 79.040 28.630 ;
        RECT 71.450 28.610 72.220 28.620 ;
        RECT 71.450 28.570 71.690 28.610 ;
        RECT 79.580 28.590 79.890 28.630 ;
        RECT 68.190 28.370 71.690 28.570 ;
        RECT 68.190 28.360 70.880 28.370 ;
        RECT 72.220 20.930 118.010 20.940 ;
        RECT 72.220 20.440 118.220 20.930 ;
        RECT 116.210 3.140 118.220 20.440 ;
        RECT 116.150 2.620 118.220 3.140 ;
        RECT 116.150 2.490 118.180 2.620 ;
    END
  END DIG21
  PIN DIG29
    PORT
      LAYER met2 ;
        RECT 107.960 3.840 108.150 4.010 ;
        RECT 107.960 3.650 112.960 3.840 ;
        RECT 112.770 3.120 112.960 3.650 ;
        RECT 113.610 3.120 113.800 3.190 ;
        RECT 112.100 2.470 114.130 3.120 ;
    END
  END DIG29
  PIN DIG28
    PORT
      LAYER met2 ;
        RECT 106.990 3.050 107.200 4.030 ;
        RECT 108.120 3.050 110.150 3.140 ;
        RECT 106.990 2.840 110.150 3.050 ;
        RECT 108.120 2.490 110.150 2.840 ;
    END
  END DIG28
  PIN DIG27
    PORT
      LAYER met2 ;
        RECT 105.060 3.140 105.270 4.030 ;
        RECT 103.940 2.490 105.970 3.140 ;
    END
  END DIG27
  PIN DIG26
    ANTENNAGATEAREA 30.021599 ;
    ANTENNADIFFAREA 288.843079 ;
    PORT
      LAYER nwell ;
        RECT 26.350 71.970 29.060 72.010 ;
        RECT 26.340 70.320 29.060 71.970 ;
        RECT 26.350 68.980 29.060 69.020 ;
        RECT 26.340 66.320 29.060 68.980 ;
        RECT 60.410 47.710 63.830 53.760 ;
        RECT 80.180 47.470 83.490 59.530 ;
        RECT 89.970 58.790 91.700 59.540 ;
        RECT 89.960 55.220 91.700 58.790 ;
        RECT 85.220 51.120 87.940 52.770 ;
        RECT 89.970 52.760 91.700 55.220 ;
        RECT 85.230 51.080 87.940 51.120 ;
        RECT 85.230 49.750 87.940 49.790 ;
        RECT 85.220 49.690 87.940 49.750 ;
        RECT 84.140 49.680 87.940 49.690 ;
        RECT 85.220 48.100 87.940 49.680 ;
        RECT 89.960 49.190 91.700 52.760 ;
        RECT 89.970 47.600 91.700 49.190 ;
        RECT 88.340 47.470 91.700 47.600 ;
        RECT 99.540 58.790 101.270 59.540 ;
        RECT 99.540 55.220 101.280 58.790 ;
        RECT 103.300 57.150 106.020 58.800 ;
        RECT 103.300 57.110 106.010 57.150 ;
        RECT 107.750 55.830 111.060 59.540 ;
        RECT 105.740 55.820 111.060 55.830 ;
        RECT 103.300 55.720 111.060 55.820 ;
        RECT 99.540 52.760 101.270 55.220 ;
        RECT 103.300 54.130 112.230 55.720 ;
        RECT 105.740 52.770 112.230 54.130 ;
        RECT 99.540 49.190 101.280 52.760 ;
        RECT 103.300 51.080 112.230 52.770 ;
        RECT 105.740 49.790 112.230 51.080 ;
        RECT 103.300 49.780 112.230 49.790 ;
        RECT 103.300 49.750 106.010 49.780 ;
        RECT 99.540 47.470 101.270 49.190 ;
        RECT 103.300 48.100 106.020 49.750 ;
        RECT 107.090 47.470 112.230 49.780 ;
        RECT 80.830 45.740 82.560 47.470 ;
        RECT 80.820 43.900 82.560 45.740 ;
        RECT 80.830 41.550 82.560 43.900 ;
        RECT 88.340 41.570 90.900 47.470 ;
        RECT 107.090 43.640 108.950 47.470 ;
        RECT 110.950 43.640 112.230 47.470 ;
        RECT 88.340 41.560 90.890 41.570 ;
        RECT 17.720 29.600 18.280 31.570 ;
        RECT 44.580 26.700 47.090 32.940 ;
        RECT 12.550 15.240 13.170 20.940 ;
        RECT 50.830 16.550 51.850 22.250 ;
        RECT 60.640 16.580 61.660 22.280 ;
        RECT 107.860 4.650 109.210 20.120 ;
        RECT 107.850 4.180 109.210 4.650 ;
      LAYER met3 ;
        RECT 77.230 57.250 77.680 58.000 ;
        RECT 77.230 51.090 77.600 57.250 ;
        RECT 78.270 57.240 78.720 57.990 ;
        RECT 78.350 54.600 78.720 57.240 ;
        RECT 78.350 54.000 78.790 54.600 ;
        RECT 77.230 50.760 77.720 51.090 ;
        RECT 77.280 50.600 77.720 50.760 ;
        RECT 78.350 48.890 78.720 54.000 ;
        RECT 78.340 48.020 78.810 48.890 ;
    END
  END DIG26
  PIN DIG25
    ANTENNAGATEAREA 30.021599 ;
    ANTENNADIFFAREA 277.819702 ;
    PORT
      LAYER met2 ;
        RECT 0.770 72.770 1.450 73.990 ;
        RECT 2.000 72.770 2.450 72.870 ;
        RECT 0.770 72.540 2.450 72.770 ;
        RECT 0.770 71.670 1.450 72.540 ;
        RECT 2.000 72.440 2.450 72.540 ;
        RECT 84.620 72.200 85.080 72.220 ;
        RECT 115.490 72.200 116.350 73.550 ;
        RECT 84.620 71.830 116.350 72.200 ;
        RECT 84.620 71.810 85.080 71.830 ;
        RECT 115.490 71.450 116.350 71.830 ;
        RECT 6.970 70.020 7.290 70.340 ;
        RECT 2.100 68.970 2.530 69.440 ;
        RECT 6.990 68.980 7.260 70.020 ;
        RECT 4.470 68.970 7.260 68.980 ;
        RECT 2.100 68.960 7.260 68.970 ;
        RECT 2.190 68.750 7.260 68.960 ;
        RECT 2.190 68.740 6.740 68.750 ;
        RECT 42.240 66.920 42.740 66.940 ;
        RECT 47.980 66.920 48.420 66.970 ;
        RECT 62.350 66.920 62.850 66.940 ;
        RECT 42.240 66.500 68.750 66.920 ;
        RECT 42.390 66.480 68.750 66.500 ;
        RECT 47.980 66.470 48.420 66.480 ;
        RECT 68.150 66.460 68.650 66.480 ;
        RECT 39.490 63.710 39.790 63.770 ;
        RECT 80.810 63.710 81.110 63.740 ;
        RECT 39.490 63.480 81.180 63.710 ;
        RECT 39.490 63.450 39.790 63.480 ;
        RECT 80.810 63.400 81.110 63.480 ;
        RECT 32.410 63.050 32.720 63.070 ;
        RECT 22.620 62.970 22.940 62.980 ;
        RECT 32.410 62.970 32.730 63.050 ;
        RECT 56.590 62.980 56.910 63.000 ;
        RECT 56.590 62.970 56.920 62.980 ;
        RECT 63.360 62.970 63.680 63.000 ;
        RECT 78.130 62.970 78.450 62.990 ;
        RECT 92.790 62.970 93.350 63.110 ;
        RECT 22.620 62.740 93.350 62.970 ;
        RECT 22.620 62.660 22.940 62.740 ;
        RECT 32.410 62.730 32.720 62.740 ;
        RECT 56.590 62.720 56.920 62.740 ;
        RECT 63.360 62.720 63.680 62.740 ;
        RECT 78.130 62.730 78.450 62.740 ;
        RECT 92.790 62.600 93.350 62.740 ;
        RECT 28.410 62.520 28.780 62.580 ;
        RECT 91.610 62.520 92.150 62.540 ;
        RECT 28.410 62.290 92.150 62.520 ;
        RECT 28.410 62.230 28.780 62.290 ;
        RECT 60.210 62.070 60.490 62.080 ;
        RECT 31.240 62.060 31.550 62.070 ;
        RECT 60.190 62.060 60.510 62.070 ;
        RECT 62.920 62.060 63.240 62.090 ;
        RECT 77.240 62.060 77.560 62.120 ;
        RECT 90.530 62.060 91.070 62.070 ;
        RECT 31.240 61.830 91.070 62.060 ;
        RECT 91.610 61.980 92.150 62.290 ;
        RECT 31.240 61.800 31.570 61.830 ;
        RECT 60.190 61.810 60.510 61.830 ;
        RECT 62.920 61.810 63.240 61.830 ;
        RECT 60.210 61.800 60.490 61.810 ;
        RECT 31.240 61.780 31.550 61.800 ;
        RECT 90.530 61.510 91.070 61.830 ;
        RECT 0.280 61.370 0.790 61.390 ;
        RECT 19.920 61.370 20.320 61.380 ;
        RECT 0.280 61.020 20.320 61.370 ;
        RECT 0.280 60.980 0.790 61.020 ;
        RECT 19.920 60.990 20.320 61.020 ;
        RECT 40.560 60.060 40.820 60.860 ;
        RECT 69.480 60.440 69.760 60.460 ;
        RECT 69.460 60.410 69.780 60.440 ;
        RECT 101.600 60.410 102.940 60.950 ;
        RECT 69.460 60.200 102.940 60.410 ;
        RECT 69.460 60.180 69.780 60.200 ;
        RECT 69.480 60.160 69.760 60.180 ;
        RECT 42.560 60.060 42.900 60.120 ;
        RECT 40.460 59.840 42.900 60.060 ;
        RECT 101.600 59.670 102.940 60.200 ;
        RECT 82.590 59.050 82.910 59.060 ;
        RECT 82.350 59.040 82.910 59.050 ;
        RECT 108.580 59.040 108.890 59.050 ;
        RECT 80.180 58.960 91.700 59.040 ;
        RECT 99.530 58.960 111.060 59.040 ;
        RECT 115.460 58.960 116.320 60.940 ;
        RECT 80.180 58.860 116.320 58.960 ;
        RECT 82.350 58.720 82.660 58.860 ;
        RECT 87.110 58.840 116.320 58.860 ;
        RECT 15.800 58.550 16.110 58.640 ;
        RECT 15.200 58.380 16.110 58.550 ;
        RECT 15.800 58.360 16.110 58.380 ;
        RECT 16.890 58.560 17.200 58.650 ;
        RECT 87.110 58.590 116.210 58.840 ;
        RECT 87.110 58.560 87.520 58.590 ;
        RECT 16.890 58.390 18.000 58.560 ;
        RECT 16.890 58.360 17.200 58.390 ;
        RECT 20.300 58.360 20.590 58.380 ;
        RECT 7.850 57.960 20.610 58.360 ;
        RECT 0.290 55.270 1.560 56.140 ;
        RECT 7.850 55.270 8.250 57.960 ;
        RECT 15.330 57.900 15.650 57.960 ;
        RECT 20.300 57.950 20.590 57.960 ;
        RECT 77.180 57.650 77.760 58.090 ;
        RECT 77.180 57.460 77.820 57.650 ;
        RECT 11.650 57.280 12.020 57.290 ;
        RECT 9.860 57.050 12.020 57.280 ;
        RECT 15.330 57.220 15.650 57.300 ;
        RECT 15.200 57.050 15.650 57.220 ;
        RECT 20.310 57.060 20.630 57.110 ;
        RECT 9.860 56.920 17.280 57.050 ;
        RECT 9.860 56.220 10.480 56.920 ;
        RECT 11.650 56.880 17.280 56.920 ;
        RECT 19.740 56.890 20.690 57.060 ;
        RECT 20.310 56.850 20.630 56.890 ;
        RECT 77.580 56.850 77.820 57.460 ;
        RECT 78.200 57.450 78.780 58.080 ;
        RECT 108.730 58.020 109.040 58.090 ;
        RECT 81.020 57.940 81.490 58.000 ;
        RECT 105.920 57.950 106.210 57.960 ;
        RECT 105.920 57.940 106.220 57.950 ;
        RECT 108.730 57.940 111.060 58.020 ;
        RECT 116.450 57.940 116.900 57.960 ;
        RECT 81.020 57.510 116.910 57.940 ;
        RECT 81.960 57.500 82.270 57.510 ;
        RECT 105.920 57.500 106.220 57.510 ;
        RECT 81.960 57.310 91.700 57.500 ;
        RECT 105.920 57.480 106.210 57.500 ;
        RECT 81.960 57.190 82.270 57.310 ;
        RECT 15.800 56.710 16.110 56.800 ;
        RECT 15.200 56.540 16.110 56.710 ;
        RECT 16.890 56.720 17.200 56.810 ;
        RECT 15.800 56.470 16.110 56.540 ;
        RECT 16.540 56.640 16.860 56.690 ;
        RECT 16.890 56.640 18.000 56.720 ;
        RECT 109.670 56.680 109.990 56.940 ;
        RECT 115.950 56.830 116.310 56.840 ;
        RECT 102.100 56.650 102.400 56.670 ;
        RECT 109.710 56.660 110.890 56.680 ;
        RECT 109.710 56.650 110.930 56.660 ;
        RECT 115.390 56.650 116.310 56.830 ;
        RECT 16.540 56.550 18.000 56.640 ;
        RECT 81.240 56.620 81.560 56.650 ;
        RECT 16.540 56.470 17.280 56.550 ;
        RECT 16.540 56.430 16.860 56.470 ;
        RECT 81.240 56.390 91.700 56.620 ;
        RECT 102.090 56.550 116.310 56.650 ;
        RECT 15.330 56.300 15.650 56.380 ;
        RECT 11.650 56.220 12.020 56.260 ;
        RECT 0.290 54.870 8.250 55.270 ;
        RECT 9.330 56.130 12.020 56.220 ;
        RECT 15.200 56.130 15.650 56.300 ;
        RECT 102.090 56.230 116.350 56.550 ;
        RECT 102.100 56.210 102.400 56.230 ;
        RECT 20.310 56.140 20.630 56.190 ;
        RECT 9.330 55.960 17.280 56.130 ;
        RECT 19.740 55.970 20.690 56.140 ;
        RECT 109.670 56.080 109.990 56.230 ;
        RECT 9.330 55.850 12.020 55.960 ;
        RECT 20.310 55.930 20.630 55.970 ;
        RECT 115.390 55.890 116.350 56.230 ;
        RECT 9.330 55.740 10.480 55.850 ;
        RECT 9.330 55.290 10.440 55.740 ;
        RECT 15.610 55.710 15.920 55.820 ;
        RECT 15.200 55.520 15.920 55.710 ;
        RECT 15.610 55.490 15.920 55.520 ;
        RECT 16.510 55.720 16.830 55.770 ;
        RECT 16.510 55.650 17.280 55.720 ;
        RECT 16.510 55.550 18.000 55.650 ;
        RECT 16.510 55.510 16.830 55.550 ;
        RECT 16.910 55.450 18.000 55.550 ;
        RECT 81.950 55.640 82.260 55.830 ;
        RECT 106.490 55.720 107.610 55.730 ;
        RECT 84.330 55.640 84.650 55.700 ;
        RECT 81.950 55.580 91.700 55.640 ;
        RECT 105.620 55.580 109.140 55.720 ;
        RECT 81.950 55.520 109.140 55.580 ;
        RECT 81.950 55.510 107.610 55.520 ;
        RECT 81.950 55.500 106.920 55.510 ;
        RECT 81.980 55.450 106.920 55.500 ;
        RECT 16.910 55.390 17.220 55.450 ;
        RECT 84.330 55.400 106.920 55.450 ;
        RECT 107.260 55.390 107.570 55.510 ;
        RECT 107.700 55.450 108.650 55.520 ;
        RECT 108.340 55.380 108.650 55.450 ;
        RECT 108.830 55.390 109.140 55.520 ;
        RECT 109.310 55.380 109.620 55.430 ;
        RECT 111.560 55.380 111.870 55.480 ;
        RECT 11.650 55.290 12.020 55.330 ;
        RECT 15.610 55.290 15.930 55.350 ;
        RECT 9.330 55.210 12.020 55.290 ;
        RECT 15.200 55.210 15.930 55.290 ;
        RECT 20.280 55.220 20.600 55.270 ;
        RECT 108.730 55.260 109.040 55.330 ;
        RECT 109.310 55.260 111.870 55.380 ;
        RECT 9.330 55.040 17.280 55.210 ;
        RECT 19.740 55.050 20.690 55.220 ;
        RECT 108.730 55.150 111.870 55.260 ;
        RECT 108.730 55.050 111.060 55.150 ;
        RECT 9.330 54.920 12.020 55.040 ;
        RECT 15.610 55.030 15.930 55.040 ;
        RECT 20.280 55.010 20.600 55.050 ;
        RECT 108.730 55.000 109.040 55.050 ;
        RECT 9.330 54.880 10.230 54.920 ;
        RECT 0.290 54.260 1.560 54.870 ;
        RECT 0.720 50.330 1.990 51.210 ;
        RECT 9.330 50.330 9.700 54.880 ;
        RECT 15.610 54.750 15.920 54.860 ;
        RECT 15.200 54.560 15.920 54.750 ;
        RECT 16.520 54.800 16.840 54.850 ;
        RECT 108.490 54.840 108.800 54.880 ;
        RECT 16.520 54.690 17.280 54.800 ;
        RECT 108.310 54.780 109.030 54.840 ;
        RECT 108.180 54.740 109.030 54.780 ;
        RECT 109.260 54.770 109.570 54.780 ;
        RECT 109.190 54.740 109.570 54.770 ;
        RECT 16.520 54.630 18.000 54.690 ;
        RECT 16.520 54.590 16.840 54.630 ;
        RECT 15.610 54.530 15.920 54.560 ;
        RECT 16.910 54.490 18.000 54.630 ;
        RECT 16.910 54.430 17.220 54.490 ;
        RECT 87.480 54.410 96.630 54.640 ;
        RECT 105.620 54.540 106.230 54.740 ;
        RECT 108.130 54.540 110.380 54.740 ;
        RECT 105.910 54.450 106.230 54.540 ;
        RECT 108.180 54.520 108.500 54.540 ;
        RECT 108.760 54.490 109.570 54.540 ;
        RECT 108.760 54.480 109.030 54.490 ;
        RECT 109.260 54.450 109.570 54.490 ;
        RECT 115.450 54.460 116.350 55.890 ;
        RECT 15.610 54.330 15.930 54.390 ;
        RECT 15.200 54.210 15.930 54.330 ;
        RECT 96.340 54.310 96.630 54.410 ;
        RECT 10.810 54.190 17.300 54.210 ;
        RECT 0.720 49.960 9.700 50.330 ;
        RECT 10.520 54.020 17.300 54.190 ;
        RECT 96.340 54.160 105.460 54.310 ;
        RECT 107.370 54.200 107.680 54.340 ;
        RECT 105.910 54.160 106.230 54.180 ;
        RECT 107.020 54.160 107.680 54.200 ;
        RECT 108.580 54.170 108.890 54.310 ;
        RECT 108.580 54.160 111.060 54.170 ;
        RECT 96.340 54.110 111.060 54.160 ;
        RECT 96.340 54.100 96.630 54.110 ;
        RECT 10.520 53.840 12.020 54.020 ;
        RECT 99.530 54.010 111.060 54.110 ;
        RECT 10.520 53.250 11.180 53.840 ;
        RECT 11.650 53.800 12.020 53.840 ;
        RECT 15.610 53.830 15.920 53.900 ;
        RECT 105.620 53.890 106.230 54.010 ;
        RECT 107.020 53.980 107.370 54.010 ;
        RECT 108.130 53.990 111.060 54.010 ;
        RECT 108.130 53.890 110.380 53.990 ;
        RECT 108.180 53.850 108.500 53.890 ;
        RECT 108.830 53.830 109.570 53.890 ;
        RECT 15.610 53.790 16.190 53.830 ;
        RECT 108.540 53.810 109.570 53.830 ;
        RECT 16.910 53.790 17.220 53.800 ;
        RECT 15.200 53.730 17.300 53.790 ;
        RECT 15.200 53.600 18.000 53.730 ;
        RECT 15.610 53.570 16.190 53.600 ;
        RECT 16.910 53.530 18.000 53.600 ;
        RECT 87.480 53.690 95.690 53.810 ;
        RECT 108.490 53.690 109.570 53.810 ;
        RECT 87.480 53.590 103.630 53.690 ;
        RECT 16.910 53.470 17.220 53.530 ;
        RECT 95.470 53.490 103.630 53.590 ;
        RECT 108.490 53.570 109.050 53.690 ;
        RECT 109.260 53.610 109.570 53.690 ;
        RECT 108.490 53.560 108.960 53.570 ;
        RECT 15.610 53.370 15.930 53.430 ;
        RECT 15.200 53.250 15.930 53.370 ;
        RECT 10.520 53.060 17.300 53.250 ;
        RECT 10.520 52.880 12.020 53.060 ;
        RECT 10.520 52.870 11.190 52.880 ;
        RECT 10.520 52.830 11.180 52.870 ;
        RECT 11.650 52.840 12.020 52.880 ;
        RECT 15.830 52.830 16.150 52.870 ;
        RECT 0.720 49.330 1.990 49.960 ;
        RECT 0.660 45.570 1.930 46.460 ;
        RECT 10.520 45.570 10.890 52.830 ;
        RECT 15.830 52.640 17.300 52.830 ;
        RECT 95.470 52.810 95.690 53.490 ;
        RECT 98.090 53.330 98.550 53.460 ;
        RECT 103.410 53.330 103.630 53.490 ;
        RECT 98.090 53.130 105.460 53.330 ;
        RECT 109.310 53.240 109.620 53.290 ;
        RECT 109.820 53.240 111.530 53.330 ;
        RECT 111.610 53.240 111.920 53.260 ;
        RECT 98.090 53.010 98.550 53.130 ;
        RECT 103.410 53.010 103.630 53.130 ;
        RECT 107.260 53.120 107.570 53.240 ;
        RECT 106.490 53.110 107.610 53.120 ;
        RECT 108.830 53.110 109.140 53.240 ;
        RECT 105.620 53.010 109.140 53.110 ;
        RECT 109.310 53.010 112.230 53.240 ;
        RECT 99.530 52.830 111.060 53.010 ;
        RECT 102.230 52.810 102.450 52.820 ;
        RECT 95.470 52.680 102.480 52.810 ;
        RECT 103.410 52.770 103.630 52.830 ;
        RECT 107.780 52.780 108.890 52.830 ;
        RECT 103.380 52.730 103.630 52.770 ;
        RECT 108.100 52.730 108.410 52.780 ;
        RECT 103.380 52.680 103.640 52.730 ;
        RECT 106.490 52.700 107.610 52.710 ;
        RECT 108.580 52.700 108.890 52.780 ;
        RECT 15.830 52.610 16.150 52.640 ;
        RECT 95.470 52.560 105.460 52.680 ;
        RECT 15.870 51.870 16.190 51.910 ;
        RECT 15.870 51.680 17.300 51.870 ;
        RECT 95.470 51.830 95.690 52.560 ;
        RECT 99.100 52.480 105.460 52.560 ;
        RECT 105.620 52.500 109.140 52.700 ;
        RECT 111.330 52.680 111.530 53.010 ;
        RECT 111.610 52.930 111.920 53.010 ;
        RECT 106.490 52.490 107.610 52.500 ;
        RECT 99.100 52.360 99.460 52.480 ;
        RECT 95.470 51.700 99.160 51.830 ;
        RECT 102.190 51.700 102.480 52.480 ;
        RECT 103.380 52.090 103.640 52.480 ;
        RECT 107.260 52.370 107.570 52.490 ;
        RECT 108.830 52.370 109.140 52.500 ;
        RECT 109.820 52.480 111.530 52.680 ;
        RECT 109.310 52.410 109.620 52.470 ;
        RECT 111.330 52.410 111.530 52.480 ;
        RECT 111.600 52.410 111.910 52.540 ;
        RECT 109.310 52.190 112.230 52.410 ;
        RECT 109.310 52.140 109.620 52.190 ;
        RECT 103.380 51.880 107.510 52.090 ;
        RECT 107.300 51.740 107.510 51.880 ;
        RECT 108.730 51.990 109.040 52.060 ;
        RECT 108.730 51.770 111.060 51.990 ;
        RECT 108.180 51.740 108.500 51.760 ;
        RECT 108.730 51.740 109.040 51.770 ;
        RECT 109.260 51.750 109.570 51.770 ;
        RECT 109.190 51.740 109.570 51.750 ;
        RECT 107.300 51.720 109.570 51.740 ;
        RECT 15.870 51.650 16.190 51.680 ;
        RECT 95.470 51.500 105.460 51.700 ;
        RECT 105.620 51.520 106.230 51.720 ;
        RECT 107.300 51.530 110.380 51.720 ;
        RECT 108.130 51.520 110.380 51.530 ;
        RECT 95.470 51.490 97.070 51.500 ;
        RECT 60.190 51.400 60.500 51.410 ;
        RECT 60.180 51.340 60.510 51.400 ;
        RECT 59.830 51.290 60.510 51.340 ;
        RECT 56.600 51.210 60.510 51.290 ;
        RECT 61.830 51.260 63.780 51.400 ;
        RECT 98.930 51.290 99.160 51.500 ;
        RECT 102.190 51.390 102.480 51.500 ;
        RECT 105.910 51.430 106.230 51.520 ;
        RECT 108.180 51.500 108.500 51.520 ;
        RECT 109.190 51.490 109.570 51.520 ;
        RECT 111.330 51.430 111.530 52.190 ;
        RECT 115.420 51.430 116.320 52.100 ;
        RECT 102.190 51.290 105.080 51.390 ;
        RECT 61.760 51.240 63.780 51.260 ;
        RECT 61.760 51.210 62.080 51.240 ;
        RECT 62.560 51.230 63.780 51.240 ;
        RECT 63.260 51.220 63.780 51.230 ;
        RECT 56.600 51.070 62.080 51.210 ;
        RECT 87.480 51.090 105.460 51.290 ;
        RECT 59.350 51.020 62.080 51.070 ;
        RECT 59.350 50.970 59.670 51.020 ;
        RECT 61.760 51.000 62.080 51.020 ;
        RECT 98.930 51.040 99.160 51.090 ;
        RECT 105.910 51.070 106.230 51.160 ;
        RECT 108.180 51.070 108.500 51.090 ;
        RECT 109.190 51.070 109.510 51.100 ;
        RECT 98.930 50.890 99.150 51.040 ;
        RECT 105.620 50.940 106.230 51.070 ;
        RECT 108.130 50.940 110.380 51.070 ;
        RECT 103.300 50.890 110.380 50.940 ;
        RECT 98.930 50.870 110.380 50.890 ;
        RECT 111.330 51.000 116.320 51.430 ;
        RECT 98.930 50.730 109.570 50.870 ;
        RECT 98.930 50.670 103.690 50.730 ;
        RECT 109.260 50.650 109.570 50.730 ;
        RECT 109.670 50.650 109.990 50.870 ;
        RECT 109.710 50.630 110.890 50.650 ;
        RECT 100.020 50.420 100.410 50.440 ;
        RECT 100.010 50.310 100.420 50.420 ;
        RECT 109.710 50.370 110.930 50.630 ;
        RECT 100.010 50.110 105.460 50.310 ;
        RECT 109.310 50.250 109.620 50.330 ;
        RECT 109.710 50.310 110.890 50.370 ;
        RECT 111.330 50.310 111.530 51.000 ;
        RECT 109.670 50.290 111.530 50.310 ;
        RECT 109.670 50.250 111.830 50.290 ;
        RECT 100.010 50.020 100.420 50.110 ;
        RECT 107.260 50.100 107.570 50.220 ;
        RECT 108.830 50.170 109.140 50.220 ;
        RECT 106.490 50.090 107.610 50.100 ;
        RECT 108.740 50.090 109.140 50.170 ;
        RECT 105.620 50.020 109.140 50.090 ;
        RECT 92.550 49.890 109.140 50.020 ;
        RECT 109.310 50.020 112.020 50.250 ;
        RECT 109.310 50.000 109.620 50.020 ;
        RECT 111.330 49.960 111.830 50.020 ;
        RECT 115.420 50.010 116.320 51.000 ;
        RECT 92.550 49.870 109.060 49.890 ;
        RECT 92.550 49.720 92.870 49.870 ;
        RECT 98.350 49.720 98.670 49.870 ;
        RECT 100.840 49.720 101.240 49.730 ;
        RECT 100.820 49.660 101.260 49.720 ;
        RECT 108.340 49.670 108.650 49.680 ;
        RECT 107.770 49.660 108.650 49.670 ;
        RECT 111.330 49.660 111.530 49.960 ;
        RECT 84.380 49.520 84.700 49.640 ;
        RECT 100.820 49.520 105.460 49.660 ;
        RECT 106.580 49.520 106.900 49.640 ;
        RECT 84.380 49.340 106.900 49.520 ;
        RECT 107.700 49.420 108.650 49.660 ;
        RECT 109.820 49.540 111.530 49.660 ;
        RECT 109.820 49.460 111.500 49.540 ;
        RECT 108.340 49.350 108.650 49.420 ;
        RECT 109.310 49.350 109.620 49.400 ;
        RECT 111.560 49.350 111.870 49.450 ;
        RECT 108.730 49.230 109.040 49.300 ;
        RECT 109.310 49.230 111.870 49.350 ;
        RECT 108.730 49.120 111.870 49.230 ;
        RECT 108.730 49.020 111.060 49.120 ;
        RECT 108.730 48.970 109.040 49.020 ;
        RECT 108.490 48.810 108.800 48.850 ;
        RECT 108.310 48.670 109.030 48.810 ;
        RECT 109.260 48.670 109.570 48.750 ;
        RECT 108.310 48.560 109.570 48.670 ;
        RECT 108.490 48.520 109.570 48.560 ;
        RECT 108.760 48.460 109.570 48.520 ;
        RECT 108.760 48.450 109.030 48.460 ;
        RECT 109.260 48.420 109.570 48.460 ;
        RECT 107.370 48.170 107.680 48.310 ;
        RECT 93.490 48.130 103.630 48.160 ;
        RECT 107.020 48.130 107.680 48.170 ;
        RECT 108.580 48.140 108.890 48.280 ;
        RECT 108.580 48.130 111.060 48.140 ;
        RECT 93.490 47.980 111.060 48.130 ;
        RECT 93.490 47.940 103.630 47.980 ;
        RECT 107.020 47.950 107.370 47.980 ;
        RECT 108.580 47.960 111.060 47.980 ;
        RECT 108.580 47.950 108.890 47.960 ;
        RECT 103.410 46.740 103.630 47.940 ;
        RECT 108.830 47.880 109.030 47.890 ;
        RECT 108.830 47.870 109.050 47.880 ;
        RECT 109.260 47.870 109.570 47.910 ;
        RECT 108.830 47.800 109.570 47.870 ;
        RECT 108.540 47.780 109.570 47.800 ;
        RECT 108.490 47.660 109.570 47.780 ;
        RECT 108.490 47.540 109.050 47.660 ;
        RECT 109.260 47.580 109.570 47.660 ;
        RECT 108.490 47.530 108.960 47.540 ;
        RECT 103.380 46.700 103.630 46.740 ;
        RECT 92.620 46.530 92.940 46.580 ;
        RECT 92.620 46.280 98.640 46.530 ;
        RECT 98.320 46.210 98.640 46.280 ;
        RECT 103.380 46.060 103.640 46.700 ;
        RECT 103.380 45.850 107.510 46.060 ;
        RECT 0.660 45.200 10.890 45.570 ;
        RECT 107.300 45.710 107.510 45.850 ;
        RECT 109.260 45.710 109.570 45.790 ;
        RECT 107.300 45.500 109.570 45.710 ;
        RECT 109.260 45.460 109.570 45.500 ;
        RECT 0.660 44.580 1.930 45.200 ;
        RECT 56.830 44.780 57.150 44.790 ;
        RECT 84.640 44.780 85.100 44.850 ;
        RECT 56.830 44.500 85.100 44.780 ;
        RECT 56.830 44.450 57.150 44.500 ;
        RECT 84.640 44.440 85.100 44.500 ;
        RECT 98.320 43.990 98.640 44.000 ;
        RECT 108.760 43.990 109.090 44.130 ;
        RECT 98.320 43.830 109.090 43.990 ;
        RECT 98.320 43.820 99.010 43.830 ;
        RECT 67.660 43.660 67.970 43.680 ;
        RECT 68.340 43.660 71.190 43.740 ;
        RECT 85.230 43.660 88.060 43.740 ;
        RECT 98.320 43.700 98.640 43.820 ;
        RECT 88.430 43.660 88.740 43.680 ;
        RECT 65.500 43.640 75.560 43.660 ;
        RECT 80.840 43.640 90.900 43.660 ;
        RECT 65.500 43.490 90.900 43.640 ;
        RECT 65.500 43.480 68.060 43.490 ;
        RECT 67.660 43.350 67.970 43.480 ;
        RECT 68.340 43.440 68.760 43.490 ;
        RECT 70.750 43.460 85.430 43.490 ;
        RECT 87.740 43.440 88.060 43.490 ;
        RECT 88.340 43.480 90.900 43.490 ;
        RECT 88.430 43.350 88.740 43.480 ;
        RECT 68.570 43.110 68.890 43.190 ;
        RECT 72.500 43.110 72.820 43.120 ;
        RECT 68.570 42.930 72.820 43.110 ;
        RECT 68.570 42.870 68.890 42.930 ;
        RECT 72.500 42.860 72.820 42.930 ;
        RECT 83.580 43.110 83.900 43.120 ;
        RECT 87.510 43.110 87.830 43.190 ;
        RECT 83.580 42.930 87.830 43.110 ;
        RECT 83.580 42.860 83.900 42.930 ;
        RECT 87.510 42.870 87.830 42.930 ;
        RECT 92.700 40.810 93.300 40.870 ;
        RECT 115.420 40.810 116.320 41.840 ;
        RECT 92.700 40.340 116.320 40.810 ;
        RECT 92.700 40.290 93.300 40.340 ;
        RECT 115.420 39.750 116.320 40.340 ;
        RECT 68.240 37.710 68.550 37.850 ;
        RECT 66.080 37.530 68.650 37.710 ;
        RECT 68.240 37.520 68.550 37.530 ;
        RECT 68.240 37.280 68.550 37.300 ;
        RECT 66.080 37.100 76.160 37.280 ;
        RECT 68.240 36.970 68.550 37.100 ;
        RECT 76.010 37.090 76.160 37.100 ;
        RECT 15.830 36.840 16.140 36.860 ;
        RECT 16.490 36.840 16.800 36.860 ;
        RECT 15.830 36.370 23.150 36.840 ;
        RECT 15.830 36.350 16.140 36.370 ;
        RECT 16.490 36.350 16.800 36.370 ;
        RECT 22.680 35.690 23.150 36.370 ;
        RECT 49.450 36.700 49.760 36.720 ;
        RECT 87.090 36.700 87.540 36.730 ;
        RECT 49.450 36.290 87.540 36.700 ;
        RECT 49.450 36.270 49.760 36.290 ;
        RECT 68.240 36.280 68.550 36.290 ;
        RECT 76.040 36.280 76.180 36.290 ;
        RECT 66.070 36.100 76.180 36.280 ;
        RECT 87.090 36.270 87.540 36.290 ;
        RECT 68.240 36.080 68.550 36.100 ;
        RECT 68.240 35.850 68.550 35.860 ;
        RECT 66.080 35.810 68.550 35.850 ;
        RECT 66.080 35.690 68.640 35.810 ;
        RECT 115.450 35.690 116.350 36.660 ;
        RECT 14.500 35.560 14.760 35.630 ;
        RECT 16.550 35.560 16.870 35.580 ;
        RECT 18.310 35.560 18.640 35.600 ;
        RECT 14.500 35.370 18.640 35.560 ;
        RECT 14.500 35.310 14.760 35.370 ;
        RECT 16.550 35.320 16.870 35.370 ;
        RECT 18.310 35.330 18.640 35.370 ;
        RECT 22.680 35.220 116.350 35.690 ;
        RECT 13.950 35.160 14.270 35.200 ;
        RECT 15.890 35.160 16.210 35.220 ;
        RECT 18.810 35.160 19.130 35.200 ;
        RECT 13.950 34.970 19.130 35.160 ;
        RECT 91.610 35.100 92.180 35.220 ;
        RECT 13.950 34.940 14.270 34.970 ;
        RECT 15.890 34.960 16.210 34.970 ;
        RECT 18.810 34.940 19.130 34.970 ;
        RECT 17.290 34.580 17.600 34.650 ;
        RECT 20.290 34.600 20.590 34.620 ;
        RECT 20.280 34.580 20.600 34.600 ;
        RECT 17.290 34.370 20.600 34.580 ;
        RECT 115.450 34.570 116.350 35.220 ;
        RECT 17.290 34.320 17.600 34.370 ;
        RECT 18.060 34.360 20.600 34.370 ;
        RECT 16.120 34.140 16.430 34.210 ;
        RECT 18.060 34.140 18.280 34.360 ;
        RECT 20.280 34.340 20.600 34.360 ;
        RECT 20.290 34.320 20.590 34.340 ;
        RECT 16.120 33.920 18.280 34.140 ;
        RECT 16.120 33.880 16.430 33.920 ;
        RECT 17.800 33.420 18.120 33.480 ;
        RECT 19.670 33.450 19.960 33.470 ;
        RECT 17.800 33.410 18.280 33.420 ;
        RECT 19.660 33.410 19.980 33.450 ;
        RECT 17.800 33.220 19.980 33.410 ;
        RECT 17.800 33.210 18.280 33.220 ;
        RECT 17.800 33.160 18.120 33.210 ;
        RECT 19.660 33.190 19.980 33.220 ;
        RECT 19.670 33.170 19.960 33.190 ;
        RECT 14.970 32.810 15.290 32.830 ;
        RECT 14.750 32.590 15.290 32.810 ;
        RECT 14.970 32.570 15.290 32.590 ;
        RECT 17.720 32.230 18.040 32.350 ;
        RECT 14.750 32.030 18.040 32.230 ;
        RECT 14.750 32.020 17.730 32.030 ;
        RECT 14.750 31.810 17.730 31.830 ;
        RECT 14.750 31.620 18.050 31.810 ;
        RECT 17.730 31.490 18.050 31.620 ;
        RECT 13.980 31.290 14.270 31.300 ;
        RECT 13.970 31.270 14.290 31.290 ;
        RECT 14.970 31.270 15.290 31.280 ;
        RECT 13.970 31.050 15.290 31.270 ;
        RECT 13.970 31.030 14.290 31.050 ;
        RECT 13.980 31.010 14.270 31.030 ;
        RECT 14.970 31.020 15.290 31.050 ;
        RECT 17.780 30.810 18.100 30.860 ;
        RECT 19.240 30.810 19.560 30.860 ;
        RECT 17.780 30.600 19.560 30.810 ;
        RECT 17.780 30.540 18.100 30.600 ;
        RECT 19.240 30.560 19.560 30.600 ;
        RECT 90.490 30.450 91.040 30.460 ;
        RECT 90.490 30.430 91.050 30.450 ;
        RECT 115.420 30.430 116.320 31.580 ;
        RECT 90.490 29.960 116.320 30.430 ;
        RECT 90.490 29.950 91.050 29.960 ;
        RECT 90.490 29.930 91.040 29.950 ;
        RECT 115.420 29.490 116.320 29.960 ;
        RECT 15.080 28.230 15.390 28.240 ;
        RECT 16.170 28.230 16.480 28.240 ;
        RECT 13.760 28.220 16.480 28.230 ;
        RECT 13.530 27.910 16.480 28.220 ;
        RECT 13.530 27.900 16.470 27.910 ;
        RECT 13.530 26.280 13.880 27.900 ;
        RECT 40.460 27.840 42.900 28.060 ;
        RECT 14.530 27.550 14.840 27.560 ;
        RECT 15.630 27.550 15.940 27.560 ;
        RECT 16.730 27.550 17.040 27.560 ;
        RECT 14.500 27.230 17.660 27.550 ;
        RECT 17.340 26.280 17.660 27.230 ;
        RECT 40.560 27.040 40.820 27.840 ;
        RECT 42.560 27.780 42.900 27.840 ;
        RECT 95.680 27.620 96.240 27.690 ;
        RECT 108.400 27.620 109.080 27.680 ;
        RECT 115.930 27.620 116.590 28.260 ;
        RECT 46.740 27.360 47.070 27.380 ;
        RECT 46.730 27.280 47.080 27.360 ;
        RECT 52.480 27.280 52.800 27.340 ;
        RECT 45.390 27.220 45.710 27.230 ;
        RECT 46.730 27.220 52.800 27.280 ;
        RECT 45.390 27.120 52.800 27.220 ;
        RECT 95.680 27.210 116.590 27.620 ;
        RECT 95.680 27.160 96.240 27.210 ;
        RECT 108.400 27.150 109.080 27.210 ;
        RECT 45.390 27.050 47.080 27.120 ;
        RECT 52.480 27.070 52.800 27.120 ;
        RECT 115.930 27.110 116.590 27.210 ;
        RECT 45.390 27.020 47.020 27.050 ;
        RECT 45.390 26.970 45.710 27.020 ;
        RECT 42.310 26.660 42.640 26.900 ;
        RECT 46.790 26.660 46.900 26.820 ;
        RECT 48.170 26.790 48.470 26.800 ;
        RECT 48.160 26.660 48.480 26.790 ;
        RECT 58.700 26.660 58.980 26.960 ;
        RECT 62.730 26.660 63.030 26.940 ;
        RECT 42.310 26.640 63.030 26.660 ;
        RECT 42.310 26.610 63.020 26.640 ;
        RECT 42.310 26.500 62.960 26.610 ;
        RECT 46.120 26.280 46.560 26.290 ;
        RECT 0.800 26.270 46.560 26.280 ;
        RECT 0.800 25.860 46.580 26.270 ;
        RECT 13.530 25.460 13.880 25.860 ;
        RECT 13.530 25.310 16.480 25.460 ;
        RECT 17.340 25.310 17.660 25.860 ;
        RECT 39.270 25.850 39.750 25.860 ;
        RECT 46.100 25.850 46.580 25.860 ;
        RECT 46.120 25.840 46.560 25.850 ;
        RECT 0.780 24.890 42.760 25.310 ;
        RECT 13.530 24.260 13.880 24.890 ;
        RECT 13.530 24.130 13.910 24.260 ;
        RECT 13.530 24.090 14.280 24.130 ;
        RECT 15.080 24.090 15.390 24.110 ;
        RECT 13.530 23.790 16.480 24.090 ;
        RECT 15.080 23.780 15.390 23.790 ;
        RECT 16.170 23.760 16.480 23.790 ;
        RECT 14.530 23.410 14.840 23.420 ;
        RECT 17.340 23.410 17.660 24.890 ;
        RECT 23.830 24.390 24.660 24.890 ;
        RECT 14.510 23.080 17.660 23.410 ;
        RECT 14.510 23.070 17.570 23.080 ;
        RECT 17.420 22.870 17.710 22.890 ;
        RECT 19.650 22.870 19.960 22.890 ;
        RECT 17.410 22.510 19.960 22.870 ;
        RECT 17.420 22.490 17.710 22.510 ;
        RECT 19.650 22.490 19.960 22.510 ;
        RECT 56.950 22.000 60.010 22.010 ;
        RECT 47.140 21.970 50.200 21.980 ;
        RECT 47.050 21.640 50.200 21.970 ;
        RECT 52.480 21.970 55.540 21.980 ;
        RECT 52.480 21.640 55.630 21.970 ;
        RECT 14.370 20.670 14.680 20.680 ;
        RECT 15.460 20.670 15.770 20.680 ;
        RECT 13.050 20.660 15.770 20.670 ;
        RECT 12.820 20.350 15.770 20.660 ;
        RECT 12.820 20.340 15.760 20.350 ;
        RECT 11.610 19.910 11.980 19.920 ;
        RECT 12.820 19.910 13.170 20.340 ;
        RECT 13.820 19.990 14.130 20.000 ;
        RECT 14.920 19.990 15.230 20.000 ;
        RECT 16.020 19.990 16.330 20.000 ;
        RECT 0.720 19.090 1.990 19.790 ;
        RECT 10.290 19.530 13.170 19.910 ;
        RECT 13.790 19.670 16.950 19.990 ;
        RECT 10.290 19.090 10.670 19.530 ;
        RECT 11.610 19.510 11.980 19.530 ;
        RECT 0.720 18.710 10.670 19.090 ;
        RECT 0.720 17.910 1.990 18.710 ;
        RECT 12.820 17.900 13.170 19.530 ;
        RECT 16.630 19.210 16.950 19.670 ;
        RECT 47.050 19.550 47.370 21.640 ;
        RECT 49.870 21.630 50.180 21.640 ;
        RECT 52.500 21.630 52.810 21.640 ;
        RECT 48.230 21.260 48.540 21.290 ;
        RECT 49.320 21.260 49.630 21.270 ;
        RECT 53.050 21.260 53.360 21.270 ;
        RECT 54.140 21.260 54.450 21.290 ;
        RECT 48.230 20.960 51.180 21.260 ;
        RECT 49.320 20.940 49.630 20.960 ;
        RECT 50.430 20.920 51.180 20.960 ;
        RECT 50.800 20.790 51.180 20.920 ;
        RECT 50.830 20.360 51.180 20.790 ;
        RECT 51.500 20.960 54.450 21.260 ;
        RECT 51.500 20.920 52.250 20.960 ;
        RECT 53.050 20.940 53.360 20.960 ;
        RECT 51.500 20.790 51.880 20.920 ;
        RECT 51.500 20.360 51.850 20.790 ;
        RECT 55.310 20.360 55.630 21.640 ;
        RECT 56.860 21.670 60.010 22.000 ;
        RECT 62.290 22.000 65.350 22.010 ;
        RECT 62.290 21.670 65.440 22.000 ;
        RECT 56.860 20.360 57.180 21.670 ;
        RECT 59.680 21.660 59.990 21.670 ;
        RECT 62.310 21.660 62.620 21.670 ;
        RECT 58.040 21.290 58.350 21.320 ;
        RECT 59.130 21.290 59.440 21.300 ;
        RECT 62.860 21.290 63.170 21.300 ;
        RECT 63.950 21.290 64.260 21.320 ;
        RECT 58.040 20.990 60.990 21.290 ;
        RECT 59.130 20.970 59.440 20.990 ;
        RECT 60.240 20.950 60.990 20.990 ;
        RECT 60.610 20.820 60.990 20.950 ;
        RECT 60.640 20.360 60.990 20.820 ;
        RECT 61.310 20.990 64.260 21.290 ;
        RECT 61.310 20.950 62.060 20.990 ;
        RECT 62.860 20.970 63.170 20.990 ;
        RECT 61.310 20.820 61.690 20.950 ;
        RECT 61.310 20.360 61.660 20.820 ;
        RECT 50.810 20.330 61.710 20.360 ;
        RECT 50.800 20.080 61.710 20.330 ;
        RECT 50.800 20.050 51.180 20.080 ;
        RECT 50.830 19.920 51.180 20.050 ;
        RECT 48.230 19.590 51.180 19.920 ;
        RECT 46.880 19.540 47.380 19.550 ;
        RECT 50.830 19.540 51.180 19.590 ;
        RECT 51.500 20.070 51.880 20.080 ;
        RECT 51.500 19.920 51.850 20.070 ;
        RECT 51.500 19.590 54.450 19.920 ;
        RECT 51.500 19.540 51.850 19.590 ;
        RECT 55.310 19.540 55.630 20.080 ;
        RECT 56.860 19.540 57.180 20.080 ;
        RECT 60.610 20.050 60.990 20.080 ;
        RECT 60.640 19.950 60.990 20.050 ;
        RECT 58.040 19.620 60.990 19.950 ;
        RECT 60.640 19.540 60.990 19.620 ;
        RECT 61.310 19.950 61.660 20.080 ;
        RECT 61.310 19.620 64.260 19.950 ;
        RECT 61.310 19.540 61.660 19.620 ;
        RECT 65.120 19.540 65.440 21.670 ;
        RECT 68.780 21.980 71.840 21.990 ;
        RECT 68.780 21.650 71.930 21.980 ;
        RECT 68.800 21.640 69.110 21.650 ;
        RECT 69.350 21.270 69.660 21.280 ;
        RECT 70.440 21.270 70.750 21.300 ;
        RECT 67.800 20.970 70.750 21.270 ;
        RECT 67.800 20.930 68.550 20.970 ;
        RECT 69.350 20.950 69.660 20.970 ;
        RECT 67.800 20.800 68.180 20.930 ;
        RECT 67.800 19.930 68.150 20.800 ;
        RECT 67.800 19.600 70.750 19.930 ;
        RECT 67.800 19.540 68.150 19.600 ;
        RECT 71.610 19.540 71.930 21.650 ;
        RECT 92.810 19.540 93.370 19.560 ;
        RECT 20.280 19.210 20.560 19.220 ;
        RECT 16.630 18.880 20.580 19.210 ;
        RECT 46.880 19.080 93.370 19.540 ;
        RECT 46.880 19.000 50.210 19.080 ;
        RECT 16.630 18.630 16.950 18.880 ;
        RECT 20.280 18.860 20.560 18.880 ;
        RECT 47.050 18.860 50.210 19.000 ;
        RECT 13.790 18.300 16.950 18.630 ;
        RECT 12.820 17.570 15.770 17.900 ;
        RECT 12.820 17.560 13.170 17.570 ;
        RECT 12.820 17.530 13.210 17.560 ;
        RECT 16.630 17.530 16.950 18.300 ;
        RECT 47.050 17.820 47.370 18.860 ;
        RECT 19.240 17.550 19.570 17.590 ;
        RECT 19.230 17.530 19.580 17.550 ;
        RECT 12.820 17.240 22.890 17.530 ;
        RECT 47.050 17.500 50.210 17.820 ;
        RECT 47.670 17.490 47.980 17.500 ;
        RECT 48.770 17.490 49.080 17.500 ;
        RECT 49.870 17.490 50.180 17.500 ;
        RECT 12.820 16.700 13.170 17.240 ;
        RECT 16.630 16.900 16.950 17.240 ;
        RECT 19.240 17.220 19.570 17.240 ;
        RECT 12.820 16.570 13.200 16.700 ;
        RECT 12.820 16.530 13.570 16.570 ;
        RECT 16.630 16.560 19.040 16.900 ;
        RECT 14.370 16.530 14.680 16.550 ;
        RECT 12.820 16.230 15.770 16.530 ;
        RECT 14.370 16.220 14.680 16.230 ;
        RECT 15.460 16.200 15.770 16.230 ;
        RECT 16.630 16.320 19.080 16.560 ;
        RECT 16.630 16.300 19.040 16.320 ;
        RECT 13.820 15.850 14.130 15.860 ;
        RECT 16.630 15.850 16.950 16.300 ;
        RECT 18.070 16.230 18.730 16.300 ;
        RECT 18.100 16.220 18.700 16.230 ;
        RECT 13.800 15.520 16.950 15.850 ;
        RECT 13.800 15.510 16.860 15.520 ;
        RECT 22.590 15.160 22.880 17.240 ;
        RECT 50.830 17.150 51.180 19.080 ;
        RECT 48.240 17.140 51.180 17.150 ;
        RECT 48.230 16.830 51.180 17.140 ;
        RECT 51.500 17.150 51.850 19.080 ;
        RECT 52.470 18.860 55.630 19.080 ;
        RECT 55.310 18.630 55.630 18.860 ;
        RECT 56.860 18.890 60.020 19.080 ;
        RECT 56.860 18.630 57.180 18.890 ;
        RECT 60.640 18.630 60.990 19.080 ;
        RECT 61.310 18.630 61.660 19.080 ;
        RECT 62.280 18.890 65.440 19.080 ;
        RECT 65.120 18.630 65.440 18.890 ;
        RECT 67.800 18.630 68.150 19.080 ;
        RECT 68.770 18.870 71.930 19.080 ;
        RECT 92.810 19.060 93.370 19.080 ;
        RECT 71.610 18.630 71.930 18.870 ;
        RECT 55.190 18.170 92.270 18.630 ;
        RECT 55.260 18.070 55.780 18.170 ;
        RECT 55.310 17.820 55.630 18.070 ;
        RECT 52.470 17.500 55.630 17.820 ;
        RECT 56.860 17.850 57.180 18.170 ;
        RECT 56.860 17.720 60.020 17.850 ;
        RECT 60.640 17.720 60.990 18.170 ;
        RECT 61.310 17.720 61.660 18.170 ;
        RECT 65.120 17.850 65.440 18.170 ;
        RECT 62.280 17.720 65.440 17.850 ;
        RECT 67.800 17.720 68.150 18.170 ;
        RECT 71.610 17.830 71.930 18.170 ;
        RECT 91.620 18.110 92.180 18.170 ;
        RECT 68.770 17.720 71.930 17.830 ;
        RECT 56.630 17.650 91.180 17.720 ;
        RECT 52.500 17.490 52.810 17.500 ;
        RECT 53.600 17.490 53.910 17.500 ;
        RECT 54.700 17.490 55.010 17.500 ;
        RECT 56.620 17.260 91.180 17.650 ;
        RECT 51.500 17.140 54.440 17.150 ;
        RECT 51.500 16.830 54.450 17.140 ;
        RECT 48.230 16.820 50.950 16.830 ;
        RECT 51.730 16.820 54.450 16.830 ;
        RECT 48.230 16.810 48.540 16.820 ;
        RECT 49.320 16.810 49.630 16.820 ;
        RECT 53.050 16.810 53.360 16.820 ;
        RECT 54.140 16.810 54.450 16.820 ;
        RECT 56.620 17.130 57.270 17.260 ;
        RECT 60.640 17.180 60.990 17.260 ;
        RECT 58.050 17.170 60.990 17.180 ;
        RECT 56.620 16.740 57.220 17.130 ;
        RECT 58.040 16.860 60.990 17.170 ;
        RECT 61.310 17.180 61.660 17.260 ;
        RECT 61.310 17.170 64.250 17.180 ;
        RECT 61.310 16.860 64.260 17.170 ;
        RECT 58.040 16.850 60.760 16.860 ;
        RECT 61.540 16.850 64.260 16.860 ;
        RECT 58.040 16.840 58.350 16.850 ;
        RECT 59.130 16.840 59.440 16.850 ;
        RECT 62.860 16.840 63.170 16.850 ;
        RECT 63.950 16.840 64.260 16.850 ;
        RECT 67.800 17.160 68.150 17.260 ;
        RECT 90.490 17.240 91.050 17.260 ;
        RECT 67.800 17.150 70.740 17.160 ;
        RECT 67.800 16.840 70.750 17.150 ;
        RECT 68.030 16.830 70.750 16.840 ;
        RECT 69.350 16.820 69.660 16.830 ;
        RECT 70.440 16.820 70.750 16.830 ;
        RECT 56.620 16.410 57.230 16.740 ;
        RECT 39.010 15.160 39.330 15.180 ;
        RECT 95.010 15.160 96.170 15.190 ;
        RECT 22.400 14.040 96.170 15.160 ;
        RECT 39.010 14.020 39.330 14.040 ;
        RECT 50.380 13.960 52.300 14.040 ;
        RECT 60.190 13.930 62.120 14.040 ;
        RECT 95.010 14.010 96.170 14.040 ;
        RECT 98.850 11.860 99.050 11.870 ;
        RECT 102.570 11.860 102.890 11.910 ;
        RECT 98.850 11.710 102.890 11.860 ;
        RECT 1.930 10.710 2.430 10.820 ;
        RECT 70.900 10.740 71.290 10.750 ;
        RECT 70.890 10.710 71.290 10.740 ;
        RECT 1.930 10.430 71.290 10.710 ;
        RECT 1.930 10.350 2.430 10.430 ;
        RECT 70.890 10.410 71.290 10.430 ;
        RECT 70.900 10.400 71.290 10.410 ;
        RECT 98.170 9.620 98.600 9.640 ;
        RECT 79.670 9.590 81.630 9.620 ;
        RECT 98.150 9.590 98.610 9.620 ;
        RECT 79.670 9.240 98.610 9.590 ;
        RECT 79.670 3.140 81.630 9.240 ;
        RECT 98.150 9.220 98.610 9.240 ;
        RECT 98.170 9.210 98.600 9.220 ;
        RECT 98.850 8.800 99.050 11.710 ;
        RECT 102.570 11.590 102.890 11.710 ;
        RECT 99.820 10.300 102.590 10.310 ;
        RECT 99.820 10.110 102.890 10.300 ;
        RECT 99.070 8.810 99.500 8.830 ;
        RECT 99.060 8.800 99.510 8.810 ;
        RECT 83.600 8.420 99.510 8.800 ;
        RECT 79.640 2.490 81.670 3.140 ;
        RECT 83.600 3.120 85.560 8.420 ;
        RECT 97.700 8.260 97.960 8.420 ;
        RECT 97.730 7.980 97.930 8.260 ;
        RECT 98.850 7.980 99.050 8.420 ;
        RECT 99.070 8.400 99.500 8.420 ;
        RECT 99.820 7.990 100.030 10.110 ;
        RECT 102.570 9.980 102.890 10.110 ;
        RECT 101.600 8.650 101.910 8.680 ;
        RECT 102.560 8.650 102.880 8.690 ;
        RECT 101.600 8.400 102.880 8.650 ;
        RECT 99.820 7.980 100.440 7.990 ;
        RECT 87.750 7.600 100.440 7.980 ;
        RECT 87.750 3.140 89.730 7.600 ;
        RECT 97.730 7.190 97.930 7.600 ;
        RECT 98.850 7.190 99.050 7.600 ;
        RECT 99.820 7.190 100.030 7.600 ;
        RECT 100.830 7.190 101.250 7.220 ;
        RECT 91.860 6.810 101.250 7.190 ;
        RECT 83.590 2.470 85.620 3.120 ;
        RECT 87.710 2.490 89.740 3.140 ;
        RECT 91.860 3.110 93.840 6.810 ;
        RECT 97.730 4.020 97.930 6.810 ;
        RECT 98.850 4.020 99.050 6.810 ;
        RECT 99.820 4.020 100.030 6.810 ;
        RECT 100.830 6.780 101.250 6.810 ;
        RECT 101.600 4.020 101.900 8.400 ;
        RECT 102.560 8.370 102.880 8.400 ;
        RECT 102.560 7.050 102.880 7.070 ;
        RECT 102.560 6.750 102.910 7.050 ;
        RECT 102.720 5.460 102.910 6.750 ;
        RECT 102.560 5.140 102.910 5.460 ;
        RECT 102.720 4.020 102.910 5.140 ;
        RECT 96.930 3.820 103.170 4.020 ;
        RECT 96.930 3.140 97.130 3.820 ;
        RECT 97.730 3.140 97.930 3.820 ;
        RECT 91.850 2.460 93.880 3.110 ;
        RECT 95.840 2.490 97.930 3.140 ;
        RECT 97.730 0.000 97.930 2.490 ;
        RECT 98.850 0.140 99.050 3.820 ;
        RECT 98.840 0.000 99.050 0.140 ;
        RECT 99.820 3.140 100.030 3.820 ;
        RECT 101.600 3.700 101.900 3.820 ;
        RECT 102.190 3.700 102.510 3.820 ;
        RECT 101.600 3.610 102.510 3.700 ;
        RECT 102.720 3.610 102.910 3.820 ;
        RECT 104.090 3.610 104.290 4.020 ;
        RECT 101.600 3.410 104.290 3.610 ;
        RECT 101.600 3.140 102.060 3.410 ;
        RECT 99.820 2.840 102.060 3.140 ;
        RECT 99.820 2.490 101.900 2.840 ;
        RECT 99.820 0.000 100.030 2.490 ;
        RECT 101.600 2.060 101.900 2.490 ;
        RECT 102.720 2.260 102.910 3.410 ;
        RECT 101.600 1.900 101.960 2.060 ;
        RECT 102.570 1.940 102.910 2.260 ;
        RECT 101.250 0.460 101.570 0.530 ;
        RECT 101.750 0.460 101.960 1.900 ;
        RECT 102.720 0.670 102.910 1.940 ;
        RECT 101.250 0.260 101.960 0.460 ;
        RECT 102.560 0.350 102.910 0.670 ;
        RECT 101.250 0.210 101.570 0.260 ;
        RECT 101.750 0.000 101.960 0.260 ;
        RECT 102.720 0.150 102.910 0.350 ;
        RECT 102.700 0.000 102.910 0.150 ;
      LAYER via2 ;
        RECT 77.300 57.620 77.620 57.940 ;
        RECT 78.330 57.610 78.650 57.930 ;
    END
  END DIG25
  PIN DIG16
    PORT
      LAYER met2 ;
        RECT 37.330 58.960 37.720 59.050 ;
        RECT 37.330 58.790 39.060 58.960 ;
        RECT 38.100 58.550 38.190 58.790 ;
        RECT 37.310 10.080 37.730 10.090 ;
        RECT 37.310 9.830 77.580 10.080 ;
        RECT 37.310 9.750 77.590 9.830 ;
        RECT 37.310 9.740 37.730 9.750 ;
        RECT 71.550 9.730 77.590 9.750 ;
        RECT 75.650 9.230 77.590 9.730 ;
        RECT 75.650 3.160 77.580 9.230 ;
        RECT 75.560 2.380 77.590 3.160 ;
    END
  END DIG16
  PIN DIG15
    PORT
      LAYER met2 ;
        RECT 36.730 57.420 37.060 57.430 ;
        RECT 36.710 57.320 37.080 57.420 ;
        RECT 36.710 57.150 39.060 57.320 ;
        RECT 36.710 57.040 37.080 57.150 ;
        RECT 38.100 57.000 38.190 57.150 ;
        RECT 36.710 9.460 37.090 9.470 ;
        RECT 36.710 9.130 73.510 9.460 ;
        RECT 36.710 9.120 37.090 9.130 ;
        RECT 67.440 9.120 73.510 9.130 ;
        RECT 71.550 8.800 73.510 9.120 ;
        RECT 71.550 3.140 73.500 8.800 ;
        RECT 71.490 2.490 73.520 3.140 ;
    END
  END DIG15
  PIN DIG14
    PORT
      LAYER met2 ;
        RECT 36.130 55.840 36.520 55.940 ;
        RECT 36.130 55.670 39.060 55.840 ;
        RECT 36.130 55.570 36.520 55.670 ;
        RECT 38.100 55.450 38.190 55.670 ;
        RECT 36.070 8.830 36.490 8.840 ;
        RECT 36.070 8.500 69.430 8.830 ;
        RECT 36.070 8.490 36.490 8.500 ;
        RECT 67.440 3.140 69.430 8.500 ;
        RECT 67.440 2.490 69.470 3.140 ;
    END
  END DIG14
  PIN DIG13
    PORT
      LAYER met2 ;
        RECT 35.490 54.240 35.880 54.330 ;
        RECT 35.490 54.070 39.060 54.240 ;
        RECT 35.490 53.980 35.880 54.070 ;
        RECT 35.480 8.190 35.880 8.210 ;
        RECT 35.480 7.860 65.420 8.190 ;
        RECT 35.480 7.850 35.880 7.860 ;
        RECT 63.460 3.140 65.410 7.860 ;
        RECT 63.410 2.490 65.440 3.140 ;
    END
  END DIG13
  PIN DIG12
    PORT
      LAYER met2 ;
        RECT 34.850 53.670 35.240 53.780 ;
        RECT 34.850 53.500 39.060 53.670 ;
        RECT 34.850 53.400 35.240 53.500 ;
        RECT 34.820 7.520 35.230 7.530 ;
        RECT 34.810 7.190 61.330 7.520 ;
        RECT 34.820 7.170 35.230 7.190 ;
        RECT 59.420 3.120 61.330 7.190 ;
        RECT 59.340 2.470 61.370 3.120 ;
    END
  END DIG12
  PIN DIG11
    PORT
      LAYER met2 ;
        RECT 34.240 52.100 34.630 52.200 ;
        RECT 38.100 52.100 38.190 52.350 ;
        RECT 34.240 51.930 39.060 52.100 ;
        RECT 34.240 51.830 34.630 51.930 ;
        RECT 34.240 6.900 34.650 6.910 ;
        RECT 34.240 6.880 57.310 6.900 ;
        RECT 34.240 6.570 57.320 6.880 ;
        RECT 34.240 6.560 34.650 6.570 ;
        RECT 55.320 3.190 57.320 6.570 ;
        RECT 55.290 2.490 57.320 3.190 ;
    END
  END DIG11
  PIN DIG10
    PORT
      LAYER met2 ;
        RECT 33.610 50.570 34.030 50.660 ;
        RECT 38.100 50.570 38.190 50.800 ;
        RECT 33.610 50.400 39.060 50.570 ;
        RECT 33.610 50.310 34.030 50.400 ;
        RECT 33.640 6.250 34.030 6.260 ;
        RECT 33.640 5.930 53.330 6.250 ;
        RECT 33.740 5.920 53.330 5.930 ;
        RECT 51.340 3.210 53.330 5.920 ;
        RECT 51.330 2.460 53.360 3.210 ;
    END
  END DIG10
  PIN DIG09
    PORT
      LAYER met2 ;
        RECT 33.050 49.000 33.440 49.090 ;
        RECT 38.100 49.000 38.190 49.250 ;
        RECT 33.050 48.830 39.060 49.000 ;
        RECT 33.050 48.740 33.440 48.830 ;
        RECT 33.060 5.640 33.450 5.690 ;
        RECT 33.060 5.360 49.420 5.640 ;
        RECT 33.320 5.310 49.420 5.360 ;
        RECT 47.350 2.490 49.380 5.310 ;
    END
  END DIG09
  PIN DIG08
    PORT
      LAYER met2 ;
        RECT 32.440 43.530 32.810 43.650 ;
        RECT 32.440 43.360 38.760 43.530 ;
        RECT 32.440 43.250 32.810 43.360 ;
        RECT 32.480 4.670 45.220 5.000 ;
        RECT 43.170 3.140 45.200 4.670 ;
        RECT 43.170 3.130 45.190 3.140 ;
        RECT 43.170 3.080 45.210 3.130 ;
        RECT 43.180 2.470 45.210 3.080 ;
    END
  END DIG08
  PIN DIG07
    PORT
      LAYER met2 ;
        RECT 31.800 41.940 32.190 42.030 ;
        RECT 38.100 41.940 38.190 42.220 ;
        RECT 31.800 41.770 38.760 41.940 ;
        RECT 31.800 41.680 32.190 41.770 ;
        RECT 39.090 4.370 41.110 4.390 ;
        RECT 31.930 4.360 41.110 4.370 ;
        RECT 31.830 4.040 41.110 4.360 ;
        RECT 31.830 4.030 32.220 4.040 ;
        RECT 39.070 3.160 41.110 4.040 ;
        RECT 39.070 3.150 41.090 3.160 ;
        RECT 39.070 3.080 41.120 3.150 ;
        RECT 39.090 2.490 41.120 3.080 ;
    END
  END DIG07
  PIN DIG06
    PORT
      LAYER met2 ;
        RECT 31.180 40.390 31.570 40.470 ;
        RECT 38.100 40.390 38.190 40.670 ;
        RECT 31.180 40.220 38.760 40.390 ;
        RECT 31.180 40.140 31.570 40.220 ;
        RECT 31.190 3.380 37.170 3.720 ;
        RECT 35.160 3.130 37.170 3.380 ;
        RECT 36.830 3.120 37.170 3.130 ;
        RECT 35.130 2.940 37.170 3.120 ;
        RECT 35.130 2.460 37.160 2.940 ;
    END
  END DIG06
  PIN DIG05
    PORT
      LAYER met2 ;
        RECT 30.570 38.910 30.990 39.000 ;
        RECT 38.100 38.910 38.190 39.120 ;
        RECT 30.570 38.740 38.760 38.910 ;
        RECT 30.570 38.640 30.990 38.740 ;
        RECT 30.580 3.130 31.130 3.150 ;
        RECT 30.580 2.700 33.130 3.130 ;
        RECT 31.100 2.470 33.130 2.700 ;
    END
  END DIG05
  PIN DIG04
    PORT
      LAYER met2 ;
        RECT 29.930 33.740 30.340 33.840 ;
        RECT 29.930 33.570 38.760 33.740 ;
        RECT 29.930 33.480 30.340 33.570 ;
        RECT 29.080 3.150 29.730 3.160 ;
        RECT 27.050 2.520 29.730 3.150 ;
        RECT 27.050 2.490 29.080 2.520 ;
    END
  END DIG04
  PIN DIG03
    PORT
      LAYER met2 ;
        RECT 29.270 32.170 29.660 32.280 ;
        RECT 38.100 32.170 38.190 32.450 ;
        RECT 29.270 32.000 38.760 32.170 ;
        RECT 29.270 31.900 29.660 32.000 ;
        RECT 29.250 3.780 29.740 3.980 ;
        RECT 23.640 3.760 29.740 3.780 ;
        RECT 23.070 3.480 29.740 3.760 ;
        RECT 23.070 3.380 29.650 3.480 ;
        RECT 23.070 3.150 25.050 3.380 ;
        RECT 23.050 2.490 25.080 3.150 ;
    END
  END DIG03
  PIN DIG02
    PORT
      LAYER met2 ;
        RECT 28.660 30.630 29.030 30.640 ;
        RECT 38.100 30.630 38.190 30.900 ;
        RECT 28.660 30.460 38.760 30.630 ;
        RECT 28.660 30.250 29.030 30.460 ;
        RECT 28.570 4.590 29.110 4.660 ;
        RECT 19.140 4.160 29.110 4.590 ;
        RECT 19.140 3.150 21.120 4.160 ;
        RECT 19.090 2.490 21.120 3.150 ;
    END
  END DIG02
  PIN DIG01
    PORT
      LAYER met2 ;
        RECT 27.970 29.090 28.360 29.190 ;
        RECT 38.100 29.090 38.190 29.350 ;
        RECT 27.970 28.920 38.760 29.090 ;
        RECT 27.970 28.820 28.360 28.920 ;
        RECT 27.920 5.430 28.460 5.470 ;
        RECT 15.090 5.390 28.460 5.430 ;
        RECT 15.040 5.000 28.460 5.390 ;
        RECT 15.040 3.120 17.050 5.000 ;
        RECT 27.920 4.970 28.460 5.000 ;
        RECT 15.020 2.460 17.050 3.120 ;
    END
  END DIG01
  PIN CAP2    
    ANTENNAGATEAREA 12.473400 ;
    ANTENNADIFFAREA 1.787900 ;
    PORT
      LAYER met2 ;
        RECT 25.160 61.600 25.480 61.610 ;
        RECT 89.590 61.600 90.120 61.630 ;
        RECT 25.160 61.370 90.120 61.600 ;
        RECT 25.160 61.310 25.480 61.370 ;
        RECT 89.590 61.020 90.120 61.370 ;
        RECT 89.460 52.420 89.770 52.470 ;
        RECT 89.460 52.410 89.920 52.420 ;
        RECT 89.460 52.230 91.710 52.410 ;
        RECT 89.460 52.140 89.770 52.230 ;
        RECT 89.490 48.700 89.800 48.780 ;
        RECT 89.490 48.680 91.710 48.700 ;
        RECT 87.480 48.480 105.460 48.680 ;
        RECT 89.490 48.450 89.800 48.480 ;
        RECT 93.040 48.410 93.880 48.480 ;
        RECT 89.440 25.130 90.040 25.180 ;
        RECT 115.850 25.130 117.950 26.070 ;
        RECT 89.440 24.660 117.950 25.130 ;
        RECT 89.440 24.620 90.040 24.660 ;
        RECT 115.850 23.990 117.950 24.660 ;
        RECT 115.870 23.980 116.640 23.990 ;
        RECT 65.080 16.800 65.680 17.230 ;
        RECT 65.070 16.780 65.680 16.800 ;
        RECT 71.570 16.780 72.170 17.210 ;
        RECT 89.560 16.780 90.120 16.790 ;
        RECT 65.070 16.320 90.210 16.780 ;
        RECT 65.070 16.270 65.600 16.320 ;
        RECT 65.070 16.220 65.590 16.270 ;
    END
  END CAP2    
  PIN OUTPUTTA1    
    ANTENNAGATEAREA 0.477400 ;
    PORT
      LAYER met2 ;
        RECT 6.550 68.100 6.860 68.330 ;
        RECT 3.460 68.000 6.860 68.100 ;
        RECT 3.460 67.870 6.840 68.000 ;
        RECT 3.460 67.840 3.780 67.870 ;
        RECT 112.870 65.560 113.640 65.710 ;
        RECT 3.380 65.140 113.640 65.560 ;
        RECT 112.870 65.000 113.640 65.140 ;
        RECT 112.680 45.800 113.460 45.950 ;
        RECT 115.420 45.800 116.320 46.720 ;
        RECT 112.680 45.330 116.320 45.800 ;
        RECT 112.680 45.180 113.460 45.330 ;
        RECT 115.420 44.630 116.320 45.330 ;
    END
  END OUTPUTTA1    
  PIN ROWTERM2
    PORT
      LAYER met2 ;
        RECT 86.230 64.030 86.650 64.050 ;
        RECT 115.460 64.030 116.320 65.330 ;
        RECT 86.230 63.660 116.320 64.030 ;
        RECT 86.230 63.640 86.650 63.660 ;
        RECT 115.460 63.230 116.320 63.660 ;
        RECT 86.170 41.810 86.610 41.930 ;
        RECT 75.410 41.630 86.610 41.810 ;
        RECT 86.170 41.530 86.610 41.630 ;
    END
  END ROWTERM2
  PIN COLUMN2
    ANTENNADIFFAREA 5.542100 ;
    PORT
      LAYER nwell ;
        RECT 85.220 57.150 87.940 58.800 ;
        RECT 85.220 57.110 87.930 57.150 ;
        RECT 85.220 55.780 87.930 55.820 ;
        RECT 85.220 55.720 87.940 55.780 ;
        RECT 84.130 55.710 87.940 55.720 ;
        RECT 85.220 54.130 87.940 55.710 ;
        RECT 84.580 41.550 86.810 47.600 ;
      LAYER met2 ;
        RECT 85.450 68.740 85.890 68.760 ;
        RECT 115.490 68.740 116.350 69.420 ;
        RECT 85.450 68.370 116.350 68.740 ;
        RECT 85.450 68.350 85.890 68.370 ;
        RECT 115.490 67.320 116.350 68.370 ;
        RECT 67.660 44.090 67.970 44.230 ;
        RECT 84.140 44.180 84.220 44.320 ;
        RECT 85.430 44.180 85.860 44.260 ;
        RECT 65.500 44.080 67.970 44.090 ;
        RECT 74.170 44.080 85.860 44.180 ;
        RECT 88.430 44.090 88.740 44.230 ;
        RECT 88.430 44.080 90.900 44.090 ;
        RECT 65.500 43.920 90.900 44.080 ;
        RECT 65.500 43.910 75.560 43.920 ;
        RECT 80.840 43.910 90.900 43.920 ;
        RECT 67.660 43.900 67.970 43.910 ;
        RECT 85.430 43.850 85.860 43.910 ;
        RECT 88.430 43.900 88.740 43.910 ;
    END
  END COLUMN2
  PIN GATE2
    ANTENNADIFFAREA 4.566800 ;
    PORT
      LAYER met1 ;
        RECT 100.550 73.180 103.740 74.300 ;
        RECT 101.640 60.980 102.920 73.180 ;
        RECT 101.630 59.640 102.920 60.980 ;
        RECT 101.640 59.150 102.920 59.640 ;
        RECT 102.360 56.680 102.590 59.150 ;
        RECT 102.090 56.200 102.590 56.680 ;
        RECT 102.190 47.460 102.590 56.200 ;
        RECT 106.360 54.960 106.560 55.830 ;
        RECT 106.350 54.670 106.580 54.960 ;
        RECT 106.360 53.960 106.560 54.670 ;
        RECT 106.350 53.670 106.580 53.960 ;
        RECT 106.360 51.940 106.560 53.670 ;
        RECT 106.350 51.650 106.580 51.940 ;
        RECT 106.360 50.940 106.560 51.650 ;
        RECT 106.350 50.650 106.580 50.940 ;
        RECT 106.360 49.780 106.560 50.650 ;
        RECT 102.190 26.210 102.420 47.460 ;
        RECT 102.190 25.980 102.430 26.210 ;
        RECT 102.190 20.170 102.420 25.980 ;
      LAYER via ;
        RECT 101.630 59.670 102.910 60.950 ;
        RECT 102.120 56.230 102.380 56.650 ;
    END
  END GATE2
  PIN DRAININJECT
    ANTENNADIFFAREA 0.105300 ;
    PORT
      LAYER met2 ;
        RECT 45.000 70.310 45.450 70.330 ;
        RECT 44.990 70.250 45.470 70.310 ;
        RECT 22.600 70.110 45.470 70.250 ;
        RECT 22.580 69.950 45.470 70.110 ;
        RECT 22.580 69.790 22.900 69.950 ;
        RECT 44.990 69.890 45.470 69.950 ;
        RECT 45.000 69.870 45.450 69.890 ;
        RECT 22.580 69.780 22.890 69.790 ;
    END
  END DRAININJECT
  PIN VTUN
    ANTENNADIFFAREA 0.604400 ;
    PORT
      LAYER nwell ;
        RECT 31.540 70.270 33.760 71.960 ;
      LAYER met2 ;
        RECT 41.150 69.550 41.600 69.570 ;
        RECT 41.140 69.540 41.620 69.550 ;
        RECT 64.760 69.540 66.180 69.580 ;
        RECT 41.140 69.140 66.230 69.540 ;
        RECT 41.140 69.130 41.620 69.140 ;
        RECT 41.150 69.110 41.600 69.130 ;
        RECT 64.760 69.100 66.180 69.140 ;
    END
  END VTUN
  PIN CHAROUTPUT
    ANTENNADIFFAREA 0.359600 ;
    PORT
      LAYER met2 ;
        RECT 0.770 68.580 1.450 69.460 ;
        RECT 0.770 68.550 4.430 68.580 ;
        RECT 0.770 68.290 4.730 68.550 ;
        RECT 0.770 68.260 4.430 68.290 ;
        RECT 0.770 67.140 1.450 68.260 ;
    END
  END CHAROUTPUT
  PIN LARGECAPACITOR
    ANTENNADIFFAREA 6.082200 ;
    PORT
      LAYER nwell ;
        RECT 9.520 67.390 19.210 71.990 ;
        RECT 8.920 66.000 19.210 67.390 ;
      LAYER met2 ;
        RECT 0.320 64.320 1.000 64.990 ;
        RECT 9.240 64.320 9.710 64.340 ;
        RECT 0.320 63.740 9.710 64.320 ;
        RECT 0.320 63.500 1.040 63.740 ;
        RECT 9.240 63.720 9.710 63.740 ;
        RECT 0.320 62.670 1.000 63.500 ;
    END
  END LARGECAPACITOR
  PIN DRAIN6P
    PORT
      LAYER met2 ;
        RECT 0.720 13.860 1.990 14.770 ;
        RECT 0.720 13.480 10.690 13.860 ;
        RECT 0.720 12.890 1.990 13.480 ;
        RECT 10.310 12.630 10.690 13.480 ;
        RECT 11.610 12.630 11.980 12.640 ;
        RECT 10.310 12.250 13.030 12.630 ;
        RECT 11.610 12.230 11.980 12.250 ;
    END
  END DRAIN6P
  PIN DRAIN5P
    PORT
      LAYER met2 ;
        RECT 9.880 29.540 10.290 29.560 ;
        RECT 11.650 29.540 13.640 29.560 ;
        RECT 9.880 29.500 13.640 29.540 ;
        RECT 16.620 29.500 16.930 29.550 ;
        RECT 9.880 29.280 16.930 29.500 ;
        RECT 9.880 29.170 12.030 29.280 ;
        RECT 16.620 29.220 16.930 29.280 ;
        RECT 9.880 29.150 10.290 29.170 ;
        RECT 11.650 29.150 12.020 29.170 ;
        RECT 0.660 23.300 1.930 24.080 ;
        RECT 9.890 23.300 10.300 23.320 ;
        RECT 0.660 22.930 10.300 23.300 ;
        RECT 0.660 22.200 1.930 22.930 ;
        RECT 9.890 22.910 10.300 22.930 ;
    END
  END DRAIN5P
  PIN DARIN4P
    ANTENNADIFFAREA 0.727900 ;
    PORT
      LAYER met2 ;
        RECT 0.720 32.550 1.990 33.320 ;
        RECT 0.720 32.180 6.710 32.550 ;
        RECT 0.720 31.440 1.990 32.180 ;
        RECT 6.340 30.520 6.710 32.180 ;
        RECT 6.340 30.340 12.290 30.520 ;
        RECT 6.340 30.270 12.360 30.340 ;
        RECT 13.750 30.270 15.020 30.280 ;
        RECT 15.450 30.270 15.760 30.330 ;
        RECT 6.340 30.150 15.760 30.270 ;
        RECT 11.650 30.110 15.760 30.150 ;
        RECT 12.010 30.060 15.760 30.110 ;
        RECT 15.450 30.000 15.760 30.060 ;
    END
  END DARIN4P
  PIN DRAIN5N
    ANTENNADIFFAREA 0.688800 ;
    PORT
      LAYER met2 ;
        RECT 4.650 34.200 5.420 34.390 ;
        RECT 11.650 34.200 12.040 34.220 ;
        RECT 4.650 34.160 12.040 34.200 ;
        RECT 15.420 34.160 15.730 34.210 ;
        RECT 4.650 33.950 15.730 34.160 ;
        RECT 4.650 33.830 12.030 33.950 ;
        RECT 15.420 33.880 15.730 33.950 ;
        RECT 4.650 33.650 5.420 33.830 ;
        RECT 11.650 33.810 12.020 33.830 ;
        RECT 0.720 28.410 1.990 29.230 ;
        RECT 4.650 28.410 5.450 28.550 ;
        RECT 0.720 27.910 5.450 28.410 ;
        RECT 0.720 27.350 1.990 27.910 ;
        RECT 4.650 27.780 5.450 27.910 ;
    END
  END DRAIN5N
  PIN DRAIN4N
    ANTENNADIFFAREA 0.688800 ;
    PORT
      LAYER met2 ;
        RECT 0.660 36.580 1.930 37.420 ;
        RECT 0.660 36.210 10.360 36.580 ;
        RECT 0.660 35.540 1.930 36.210 ;
        RECT 9.990 34.860 10.360 36.210 ;
        RECT 9.990 34.850 12.020 34.860 ;
        RECT 9.990 34.670 12.240 34.850 ;
        RECT 9.990 34.610 13.640 34.670 ;
        RECT 16.640 34.610 16.950 34.650 ;
        RECT 9.990 34.490 16.950 34.610 ;
        RECT 11.650 34.450 16.950 34.490 ;
        RECT 12.020 34.390 16.950 34.450 ;
        RECT 16.640 34.320 16.950 34.390 ;
    END
  END DRAIN4N
  PIN DRAIN3P
    PORT
      LAYER met2 ;
        RECT 11.650 52.100 17.300 52.290 ;
        RECT 0.720 40.730 1.990 41.640 ;
        RECT 11.650 40.730 12.020 52.100 ;
        RECT 0.720 40.360 12.020 40.730 ;
        RECT 0.720 39.760 1.990 40.360 ;
    END
  END DRAIN3P
  PIN SOURCEP
    PORT
      LAYER met2 ;
        RECT 0.000 59.170 1.270 60.630 ;
        RECT 11.350 59.170 11.650 59.180 ;
        RECT 20.940 59.170 21.230 59.190 ;
        RECT 0.000 58.780 21.260 59.170 ;
        RECT 0.000 58.750 1.270 58.780 ;
        RECT 20.940 58.760 21.230 58.780 ;
        RECT 20.920 54.150 21.240 54.180 ;
        RECT 19.710 53.950 21.340 54.150 ;
        RECT 20.920 53.920 21.240 53.950 ;
        RECT 20.930 53.190 21.250 53.220 ;
        RECT 19.710 52.990 21.340 53.190 ;
        RECT 20.930 52.960 21.250 52.990 ;
        RECT 20.920 52.230 21.240 52.260 ;
        RECT 19.710 52.030 21.340 52.230 ;
        RECT 20.920 52.000 21.240 52.030 ;
        RECT 16.140 30.250 16.450 30.320 ;
        RECT 20.930 30.270 21.220 30.290 ;
        RECT 16.140 30.240 18.280 30.250 ;
        RECT 20.920 30.240 21.240 30.270 ;
        RECT 16.140 30.040 21.240 30.240 ;
        RECT 16.140 29.990 16.450 30.040 ;
        RECT 18.070 30.030 21.240 30.040 ;
        RECT 17.330 29.420 17.640 29.490 ;
        RECT 18.070 29.420 18.280 30.030 ;
        RECT 20.920 30.010 21.240 30.030 ;
        RECT 20.930 29.990 21.220 30.010 ;
        RECT 17.330 29.210 18.280 29.420 ;
        RECT 17.330 29.160 17.640 29.210 ;
        RECT 20.860 11.660 21.170 11.680 ;
        RECT 16.630 11.320 21.170 11.660 ;
        RECT 20.860 11.300 21.170 11.320 ;
    END
  END SOURCEP
  PIN GATE1
    PORT
      LAYER met2 ;
        RECT 57.060 61.020 57.380 61.060 ;
        RECT 72.710 61.020 73.990 61.120 ;
        RECT 57.060 60.810 73.990 61.020 ;
        RECT 57.060 60.780 57.380 60.810 ;
    END
  END GATE1
  PIN VINJ
    ANTENNADIFFAREA 1.921700 ;
    PORT
      LAYER nwell ;
        RECT 3.910 68.480 6.650 71.980 ;
        RECT 20.790 65.980 24.790 71.970 ;
      LAYER met2 ;
        RECT 0.620 70.570 3.100 70.580 ;
        RECT 4.410 70.570 4.730 70.770 ;
        RECT 5.140 70.570 5.450 70.780 ;
        RECT 5.820 70.570 6.140 70.780 ;
        RECT 6.480 70.570 21.130 70.700 ;
        RECT 0.620 70.490 21.130 70.570 ;
        RECT 0.620 70.320 6.620 70.490 ;
        RECT 20.550 70.480 21.300 70.490 ;
        RECT 0.620 70.180 6.480 70.320 ;
        RECT 2.890 69.810 6.480 70.180 ;
        RECT 20.550 70.180 22.170 70.480 ;
        RECT 20.550 70.040 20.790 70.180 ;
        RECT 21.870 70.120 22.170 70.180 ;
        RECT 4.410 69.640 4.730 69.810 ;
        RECT 5.140 69.610 5.450 69.810 ;
        RECT 5.840 69.660 6.160 69.810 ;
        RECT 20.530 69.710 20.840 70.040 ;
        RECT 21.870 69.800 22.200 70.120 ;
        RECT 21.890 69.790 22.200 69.800 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.320 62.170 0.830 62.290 ;
        RECT 0.320 61.880 3.420 62.170 ;
        RECT 0.830 61.870 3.420 61.880 ;
    END
    PORT
      LAYER met2 ;
        RECT 46.660 67.930 47.160 67.960 ;
        RECT 52.380 67.930 52.880 67.960 ;
        RECT 46.660 67.520 76.820 67.930 ;
        RECT 46.810 67.490 76.820 67.520 ;
    END
  END VINJ
  PIN VGND
    ANTENNADIFFAREA 5.176000 ;
    PORT
      LAYER met2 ;
        RECT 5.120 66.930 5.430 67.140 ;
        RECT 6.550 66.930 6.860 67.160 ;
        RECT 2.770 66.770 7.690 66.930 ;
        RECT 0.960 66.600 7.690 66.770 ;
        RECT 0.960 66.550 7.700 66.600 ;
        RECT 0.960 66.440 7.720 66.550 ;
        RECT 0.960 66.370 3.230 66.440 ;
        RECT 0.960 66.170 1.360 66.370 ;
        RECT 4.330 66.230 4.640 66.440 ;
        RECT 5.260 66.230 5.570 66.440 ;
        RECT 5.960 66.230 6.270 66.440 ;
        RECT 6.700 66.260 7.720 66.440 ;
        RECT 19.810 66.260 20.120 66.380 ;
        RECT 29.670 66.260 29.980 66.400 ;
        RECT 6.700 66.230 29.980 66.260 ;
        RECT 0.610 65.770 1.360 66.170 ;
        RECT 6.720 66.070 29.980 66.230 ;
        RECT 6.720 66.050 29.950 66.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.350 74.170 60.330 74.320 ;
        RECT 59.360 66.920 60.330 74.170 ;
        RECT 59.340 66.450 60.350 66.920 ;
      LAYER via ;
        RECT 59.370 66.490 60.320 66.900 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 0.426400 ;
    PORT
      LAYER met1 ;
        RECT 50.950 22.160 51.210 22.360 ;
        RECT 51.470 22.160 51.730 22.360 ;
        RECT 50.950 21.350 51.260 22.160 ;
        RECT 51.420 21.350 51.730 22.160 ;
        RECT 50.950 20.820 51.210 21.350 ;
        RECT 50.840 20.360 51.210 20.820 ;
        RECT 50.830 20.020 51.210 20.360 ;
        RECT 50.840 18.610 51.210 20.020 ;
        RECT 51.470 20.820 51.730 21.350 ;
        RECT 51.470 20.380 51.840 20.820 ;
        RECT 51.470 20.040 51.850 20.380 ;
        RECT 51.470 18.610 51.840 20.040 ;
        RECT 50.840 15.180 51.840 18.610 ;
        RECT 50.360 15.140 52.290 15.180 ;
        RECT 49.820 13.950 52.290 15.140 ;
        RECT 49.820 2.460 50.760 13.950 ;
      LAYER via ;
        RECT 50.830 20.050 51.110 20.330 ;
        RECT 51.570 20.070 51.850 20.350 ;
        RECT 51.150 15.100 52.270 15.120 ;
        RECT 50.410 14.000 52.270 15.100 ;
        RECT 50.410 13.980 51.530 14.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 60.760 22.190 61.020 22.390 ;
        RECT 61.280 22.190 61.540 22.390 ;
        RECT 60.760 21.380 61.070 22.190 ;
        RECT 61.230 21.380 61.540 22.190 ;
        RECT 60.760 20.850 61.020 21.380 ;
        RECT 60.650 20.360 61.020 20.850 ;
        RECT 60.640 20.020 61.020 20.360 ;
        RECT 60.650 18.840 61.020 20.020 ;
        RECT 61.280 20.850 61.540 21.380 ;
        RECT 61.280 18.840 61.650 20.850 ;
        RECT 60.650 15.200 61.650 18.840 ;
        RECT 61.780 15.200 62.670 15.240 ;
        RECT 60.170 13.920 62.670 15.200 ;
        RECT 61.780 3.920 62.670 13.920 ;
        RECT 61.780 3.190 62.700 3.920 ;
        RECT 61.750 2.460 62.670 3.190 ;
      LAYER via ;
        RECT 60.640 20.050 60.920 20.330 ;
        RECT 60.220 13.950 62.080 15.140 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 15.270 52.900 17.840 55.990 ;
        RECT 38.850 54.960 40.620 61.200 ;
        RECT 44.580 54.960 47.090 61.200 ;
        RECT 84.330 55.400 84.650 55.700 ;
        RECT 39.690 53.950 39.930 54.000 ;
        RECT 39.450 53.940 40.920 53.950 ;
        RECT 39.150 53.860 40.920 53.940 ;
        RECT 45.180 53.860 47.390 53.950 ;
        RECT 53.330 53.700 54.010 53.710 ;
        RECT 38.850 46.600 40.620 52.840 ;
        RECT 44.580 46.600 47.090 52.840 ;
        RECT 53.320 47.650 54.020 53.700 ;
        RECT 77.220 50.550 77.780 51.090 ;
        RECT 84.140 49.010 84.210 49.190 ;
        RECT 65.510 47.590 68.060 47.600 ;
        RECT 38.850 36.470 40.620 42.710 ;
        RECT 44.580 36.470 47.090 42.710 ;
        RECT 60.410 37.640 63.830 43.690 ;
        RECT 65.500 41.570 68.060 47.590 ;
        RECT 65.510 41.560 68.060 41.570 ;
        RECT 69.590 41.550 71.820 47.600 ;
        RECT 73.840 45.740 75.570 47.600 ;
        RECT 73.840 43.900 75.580 45.740 ;
        RECT 84.140 44.140 84.220 44.320 ;
        RECT 73.840 41.550 75.570 43.900 ;
        RECT 74.420 37.580 76.150 38.210 ;
        RECT 74.420 34.510 76.160 37.580 ;
        RECT 74.030 34.290 74.410 34.390 ;
        RECT 13.880 28.680 16.250 31.550 ;
        RECT 38.850 26.700 40.620 32.940 ;
        RECT 53.320 27.900 55.070 33.900 ;
        RECT 60.410 27.880 63.830 33.930 ;
        RECT 74.420 32.160 76.150 34.510 ;
        RECT 78.060 34.250 78.460 34.390 ;
        RECT 55.220 22.500 57.240 26.460 ;
        RECT 55.220 22.470 59.260 22.500 ;
        RECT 13.540 18.020 13.550 18.060 ;
        RECT 14.550 15.020 17.940 20.720 ;
        RECT 46.060 16.770 49.450 22.470 ;
        RECT 50.450 19.430 50.460 19.470 ;
        RECT 52.220 19.430 52.230 19.470 ;
        RECT 53.230 16.800 59.260 22.470 ;
        RECT 60.260 19.460 60.270 19.500 ;
        RECT 62.030 19.460 62.040 19.500 ;
        RECT 63.040 16.800 66.430 22.500 ;
        RECT 53.230 16.770 56.620 16.800 ;
        RECT 96.970 0.370 102.620 16.470 ;
      LAYER li1 ;
        RECT 3.910 71.560 4.080 71.860 ;
        RECT 3.910 71.380 4.910 71.560 ;
        RECT 5.310 71.550 5.480 71.860 ;
        RECT 7.110 71.590 7.780 71.760 ;
        RECT 5.310 71.380 6.320 71.550 ;
        RECT 7.110 70.800 7.780 70.970 ;
        RECT 5.120 70.700 5.440 70.740 ;
        RECT 4.240 70.530 6.320 70.700 ;
        RECT 21.130 70.660 24.440 71.640 ;
        RECT 28.530 70.840 28.760 71.530 ;
        RECT 33.230 70.790 33.460 71.480 ;
        RECT 5.110 70.510 5.440 70.530 ;
        RECT 5.120 70.480 5.440 70.510 ;
        RECT 4.420 70.120 6.240 70.290 ;
        RECT 5.120 69.880 5.440 69.900 ;
        RECT 4.240 69.710 6.320 69.880 ;
        RECT 7.030 69.870 7.240 70.300 ;
        RECT 21.240 70.000 21.410 70.350 ;
        RECT 21.960 70.080 22.130 70.110 ;
        RECT 21.870 70.040 22.190 70.080 ;
        RECT 22.640 70.070 22.810 70.110 ;
        RECT 20.510 69.960 21.410 70.000 ;
        RECT 7.050 69.850 7.220 69.870 ;
        RECT 20.500 69.770 21.410 69.960 ;
        RECT 21.860 69.850 22.190 70.040 ;
        RECT 22.560 70.030 22.880 70.070 ;
        RECT 21.870 69.820 22.190 69.850 ;
        RECT 22.550 69.840 22.880 70.030 ;
        RECT 21.960 69.780 22.130 69.820 ;
        RECT 22.560 69.810 22.880 69.840 ;
        RECT 22.640 69.780 22.810 69.810 ;
        RECT 20.510 69.740 21.410 69.770 ;
        RECT 29.740 69.760 29.910 69.780 ;
        RECT 5.110 69.670 5.440 69.710 ;
        RECT 5.120 69.640 5.440 69.670 ;
        RECT 7.110 69.370 7.780 69.540 ;
        RECT 4.240 68.870 4.910 69.040 ;
        RECT 5.640 68.870 6.320 69.040 ;
        RECT 6.620 68.750 6.810 68.810 ;
        RECT 6.620 68.580 7.790 68.750 ;
        RECT 6.550 68.300 6.720 68.330 ;
        RECT 6.550 68.270 6.880 68.300 ;
        RECT 6.550 68.080 6.890 68.270 ;
        RECT 6.550 68.040 6.880 68.080 ;
        RECT 6.550 68.000 6.720 68.040 ;
        RECT 5.300 67.920 5.470 67.980 ;
        RECT 7.120 67.970 7.790 68.140 ;
        RECT 4.240 67.750 4.910 67.920 ;
        RECT 5.300 67.750 6.320 67.920 ;
        RECT 5.300 67.650 5.470 67.750 ;
        RECT 5.100 67.080 5.420 67.100 ;
        RECT 6.530 67.080 6.850 67.120 ;
        RECT 4.230 66.910 7.810 67.080 ;
        RECT 5.090 66.870 5.420 66.910 ;
        RECT 6.520 66.890 6.850 66.910 ;
        RECT 5.100 66.840 5.420 66.870 ;
        RECT 6.530 66.860 6.850 66.890 ;
        RECT 4.310 66.480 4.630 66.520 ;
        RECT 5.240 66.480 5.560 66.520 ;
        RECT 5.940 66.480 6.260 66.520 ;
        RECT 6.680 66.480 7.000 66.520 ;
        RECT 4.300 66.410 4.630 66.480 ;
        RECT 5.230 66.410 5.560 66.480 ;
        RECT 5.930 66.410 6.260 66.480 ;
        RECT 6.670 66.460 7.000 66.480 ;
        RECT 7.390 66.470 7.710 66.510 ;
        RECT 7.380 66.460 7.710 66.470 ;
        RECT 6.670 66.410 7.710 66.460 ;
        RECT 4.280 66.240 7.710 66.410 ;
        RECT 9.380 66.300 9.550 66.970 ;
        RECT 19.870 66.880 20.040 69.530 ;
        RECT 21.240 69.340 21.410 69.740 ;
        RECT 26.850 69.590 29.910 69.760 ;
        RECT 29.740 68.940 29.910 69.590 ;
        RECT 21.130 67.860 24.440 68.840 ;
        RECT 29.740 68.770 31.010 68.940 ;
        RECT 28.530 67.850 28.760 68.540 ;
        RECT 19.870 66.340 20.050 66.880 ;
        RECT 19.790 66.300 20.110 66.340 ;
        RECT 21.130 66.310 24.440 67.290 ;
        RECT 28.530 66.840 28.760 67.530 ;
        RECT 29.740 66.360 29.910 68.770 ;
        RECT 32.480 67.120 32.650 68.010 ;
        RECT 29.650 66.320 29.970 66.360 ;
        RECT 6.860 66.230 7.710 66.240 ;
        RECT 19.780 66.110 20.110 66.300 ;
        RECT 29.640 66.130 29.970 66.320 ;
        RECT 19.790 66.080 20.110 66.110 ;
        RECT 29.650 66.100 29.970 66.130 ;
        RECT 19.820 62.520 21.340 62.530 ;
        RECT 19.820 61.730 21.370 62.520 ;
        RECT 40.510 60.730 40.860 60.830 ;
        RECT 43.580 60.810 45.810 60.960 ;
        RECT 43.580 60.790 45.960 60.810 ;
        RECT 43.580 60.780 43.760 60.790 ;
        RECT 43.120 60.760 43.760 60.780 ;
        RECT 42.170 60.730 42.630 60.760 ;
        RECT 39.100 60.560 39.860 60.730 ;
        RECT 40.110 60.560 41.280 60.730 ;
        RECT 41.520 60.590 42.630 60.730 ;
        RECT 43.080 60.590 43.760 60.760 ;
        RECT 45.360 60.640 45.960 60.790 ;
        RECT 46.420 60.630 46.750 60.800 ;
        RECT 41.520 60.560 42.340 60.590 ;
        RECT 39.100 60.550 39.330 60.560 ;
        RECT 39.060 60.110 39.330 60.550 ;
        RECT 42.080 60.420 42.340 60.560 ;
        RECT 43.580 60.530 43.760 60.590 ;
        RECT 44.700 60.440 45.030 60.610 ;
        RECT 40.540 60.110 40.870 60.370 ;
        RECT 42.080 60.250 43.260 60.420 ;
        RECT 42.080 60.110 42.340 60.250 ;
        RECT 38.510 59.970 38.680 60.030 ;
        RECT 38.480 59.750 38.700 59.970 ;
        RECT 39.030 59.930 39.360 60.110 ;
        RECT 39.610 59.940 41.770 60.110 ;
        RECT 42.010 59.940 42.340 60.110 ;
        RECT 42.170 59.890 42.340 59.940 ;
        RECT 42.630 59.750 42.840 60.080 ;
        RECT 43.080 59.810 43.260 60.250 ;
        RECT 44.780 60.190 45.030 60.440 ;
        RECT 44.780 60.090 45.250 60.190 ;
        RECT 46.500 60.170 46.680 60.630 ;
        RECT 44.610 60.080 45.250 60.090 ;
        RECT 43.810 60.020 45.250 60.080 ;
        RECT 43.810 59.910 45.170 60.020 ;
        RECT 45.720 60.000 46.680 60.170 ;
        RECT 38.510 59.700 38.680 59.750 ;
        RECT 40.510 59.180 40.860 59.280 ;
        RECT 43.580 59.260 45.810 59.410 ;
        RECT 43.580 59.240 45.960 59.260 ;
        RECT 43.580 59.230 43.760 59.240 ;
        RECT 43.120 59.210 43.760 59.230 ;
        RECT 42.170 59.180 42.630 59.210 ;
        RECT 39.100 59.010 39.860 59.180 ;
        RECT 40.110 59.010 41.280 59.180 ;
        RECT 41.520 59.040 42.630 59.180 ;
        RECT 43.080 59.040 43.760 59.210 ;
        RECT 45.360 59.090 45.960 59.240 ;
        RECT 46.420 59.080 46.750 59.250 ;
        RECT 41.520 59.010 42.340 59.040 ;
        RECT 39.100 59.000 39.330 59.010 ;
        RECT 16.120 58.600 16.320 58.640 ;
        RECT 15.810 58.340 16.320 58.600 ;
        RECT 16.120 58.310 16.320 58.340 ;
        RECT 16.710 58.610 16.910 58.640 ;
        RECT 16.710 58.570 17.220 58.610 ;
        RECT 16.710 58.380 17.230 58.570 ;
        RECT 39.060 58.560 39.330 59.000 ;
        RECT 42.080 58.870 42.340 59.010 ;
        RECT 43.580 58.980 43.760 59.040 ;
        RECT 44.700 58.890 45.030 59.060 ;
        RECT 40.540 58.560 40.870 58.820 ;
        RECT 42.080 58.700 43.260 58.870 ;
        RECT 42.080 58.560 42.340 58.700 ;
        RECT 38.510 58.420 38.680 58.480 ;
        RECT 16.710 58.350 17.220 58.380 ;
        RECT 16.710 58.310 16.910 58.350 ;
        RECT 17.400 58.160 17.570 58.210 ;
        RECT 38.480 58.200 38.700 58.420 ;
        RECT 39.030 58.380 39.360 58.560 ;
        RECT 39.610 58.390 41.770 58.560 ;
        RECT 42.010 58.390 42.340 58.560 ;
        RECT 42.170 58.340 42.340 58.390 ;
        RECT 42.630 58.200 42.840 58.530 ;
        RECT 43.080 58.260 43.260 58.700 ;
        RECT 44.780 58.640 45.030 58.890 ;
        RECT 44.780 58.540 45.250 58.640 ;
        RECT 46.500 58.620 46.680 59.080 ;
        RECT 44.610 58.530 45.250 58.540 ;
        RECT 43.810 58.470 45.250 58.530 ;
        RECT 43.810 58.360 45.170 58.470 ;
        RECT 45.720 58.450 46.680 58.620 ;
        RECT 67.790 58.570 68.460 59.440 ;
        RECT 80.070 59.130 82.170 59.440 ;
        RECT 80.070 58.960 82.590 59.130 ;
        RECT 82.830 59.110 83.020 59.140 ;
        RECT 80.070 58.590 82.170 58.960 ;
        RECT 82.830 58.940 83.890 59.110 ;
        RECT 108.650 58.960 109.180 59.130 ;
        RECT 82.830 58.910 83.020 58.940 ;
        RECT 80.570 58.250 80.790 58.590 ;
        RECT 80.570 58.240 80.780 58.250 ;
        RECT 15.370 58.140 15.800 58.160 ;
        RECT 15.370 57.970 15.820 58.140 ;
        RECT 17.390 58.130 17.570 58.160 ;
        RECT 38.510 58.150 38.680 58.200 ;
        RECT 17.390 58.120 17.820 58.130 ;
        RECT 15.370 57.950 15.800 57.970 ;
        RECT 17.390 57.890 17.980 58.120 ;
        RECT 80.950 58.070 81.140 58.080 ;
        RECT 17.390 57.880 17.820 57.890 ;
        RECT 17.390 57.820 17.560 57.880 ;
        RECT 16.120 57.680 16.320 57.720 ;
        RECT 15.810 57.420 16.320 57.680 ;
        RECT 16.120 57.390 16.320 57.420 ;
        RECT 16.710 57.690 16.910 57.720 ;
        RECT 16.710 57.650 17.220 57.690 ;
        RECT 16.710 57.460 17.230 57.650 ;
        RECT 40.510 57.630 40.860 57.730 ;
        RECT 43.580 57.710 45.810 57.860 ;
        RECT 80.940 57.780 81.140 58.070 ;
        RECT 43.580 57.690 45.960 57.710 ;
        RECT 43.580 57.680 43.760 57.690 ;
        RECT 43.120 57.660 43.760 57.680 ;
        RECT 42.170 57.630 42.630 57.660 ;
        RECT 39.100 57.460 39.860 57.630 ;
        RECT 40.110 57.460 41.280 57.630 ;
        RECT 41.520 57.490 42.630 57.630 ;
        RECT 43.080 57.490 43.760 57.660 ;
        RECT 45.360 57.540 45.960 57.690 ;
        RECT 46.420 57.530 46.750 57.700 ;
        RECT 41.520 57.460 42.340 57.490 ;
        RECT 16.710 57.430 17.220 57.460 ;
        RECT 39.100 57.450 39.330 57.460 ;
        RECT 16.710 57.390 16.910 57.430 ;
        RECT 15.370 57.220 15.800 57.240 ;
        RECT 15.370 57.050 15.820 57.220 ;
        RECT 15.370 57.030 15.800 57.050 ;
        RECT 39.060 57.010 39.330 57.450 ;
        RECT 42.080 57.320 42.340 57.460 ;
        RECT 43.580 57.430 43.760 57.490 ;
        RECT 44.700 57.340 45.030 57.510 ;
        RECT 40.540 57.010 40.870 57.270 ;
        RECT 42.080 57.150 43.260 57.320 ;
        RECT 42.080 57.010 42.340 57.150 ;
        RECT 38.510 56.870 38.680 56.930 ;
        RECT 16.120 56.760 16.320 56.800 ;
        RECT 15.810 56.500 16.320 56.760 ;
        RECT 16.120 56.470 16.320 56.500 ;
        RECT 16.710 56.770 16.910 56.800 ;
        RECT 16.710 56.730 17.220 56.770 ;
        RECT 16.710 56.540 17.230 56.730 ;
        RECT 38.480 56.650 38.700 56.870 ;
        RECT 39.030 56.830 39.360 57.010 ;
        RECT 39.610 56.840 41.770 57.010 ;
        RECT 42.010 56.840 42.340 57.010 ;
        RECT 42.170 56.790 42.340 56.840 ;
        RECT 42.630 56.650 42.840 56.980 ;
        RECT 43.080 56.710 43.260 57.150 ;
        RECT 44.780 57.090 45.030 57.340 ;
        RECT 44.780 56.990 45.250 57.090 ;
        RECT 46.500 57.070 46.680 57.530 ;
        RECT 80.910 57.450 81.150 57.780 ;
        RECT 44.610 56.980 45.250 56.990 ;
        RECT 43.810 56.920 45.250 56.980 ;
        RECT 43.810 56.810 45.170 56.920 ;
        RECT 45.720 56.900 46.680 57.070 ;
        RECT 81.340 56.970 81.510 58.580 ;
        RECT 82.170 57.480 82.340 58.570 ;
        RECT 83.300 58.550 83.490 58.580 ;
        RECT 82.760 58.380 83.490 58.550 ;
        RECT 83.720 58.550 83.890 58.940 ;
        RECT 110.460 58.860 110.660 59.210 ;
        RECT 110.460 58.830 110.670 58.860 ;
        RECT 83.720 58.380 84.460 58.550 ;
        RECT 106.780 58.380 107.130 58.550 ;
        RECT 108.150 58.380 108.480 58.550 ;
        RECT 83.300 58.350 83.490 58.380 ;
        RECT 85.520 57.760 85.750 58.280 ;
        RECT 82.760 57.590 85.750 57.760 ;
        RECT 81.940 57.440 82.340 57.480 ;
        RECT 81.930 57.250 82.340 57.440 ;
        RECT 90.720 57.400 91.270 57.830 ;
        RECT 99.970 57.400 100.520 57.830 ;
        RECT 103.600 57.590 103.830 58.280 ;
        RECT 108.900 58.050 109.070 58.570 ;
        RECT 108.740 57.790 109.070 58.050 ;
        RECT 106.780 57.590 107.130 57.760 ;
        RECT 108.150 57.590 108.480 57.760 ;
        RECT 81.940 57.220 82.340 57.250 ;
        RECT 81.330 56.780 81.510 56.970 ;
        RECT 82.170 56.880 82.340 57.220 ;
        RECT 82.830 56.970 83.020 57.150 ;
        RECT 82.760 56.800 83.110 56.970 ;
        RECT 38.510 56.600 38.680 56.650 ;
        RECT 16.710 56.510 17.220 56.540 ;
        RECT 16.710 56.470 16.910 56.510 ;
        RECT 83.680 56.390 83.890 56.820 ;
        RECT 84.110 56.800 84.450 56.970 ;
        RECT 83.700 56.370 83.870 56.390 ;
        RECT 15.370 56.300 15.800 56.320 ;
        RECT 15.370 56.130 15.820 56.300 ;
        RECT 15.370 56.110 15.800 56.130 ;
        RECT 40.510 56.080 40.860 56.180 ;
        RECT 43.580 56.160 45.810 56.310 ;
        RECT 43.580 56.140 45.960 56.160 ;
        RECT 43.580 56.130 43.760 56.140 ;
        RECT 43.120 56.110 43.760 56.130 ;
        RECT 42.170 56.080 42.630 56.110 ;
        RECT 39.100 55.910 39.860 56.080 ;
        RECT 40.110 55.910 41.280 56.080 ;
        RECT 41.520 55.940 42.630 56.080 ;
        RECT 43.080 55.940 43.760 56.110 ;
        RECT 45.360 55.990 45.960 56.140 ;
        RECT 46.420 55.980 46.750 56.150 ;
        RECT 81.330 56.060 81.510 56.250 ;
        RECT 41.520 55.910 42.340 55.940 ;
        RECT 39.100 55.900 39.330 55.910 ;
        RECT 15.620 55.740 15.940 55.780 ;
        RECT 15.620 55.720 15.950 55.740 ;
        RECT 15.620 55.520 16.240 55.720 ;
        RECT 16.070 55.390 16.240 55.520 ;
        RECT 16.750 55.680 16.920 55.720 ;
        RECT 16.750 55.640 17.240 55.680 ;
        RECT 16.750 55.450 17.250 55.640 ;
        RECT 39.060 55.460 39.330 55.900 ;
        RECT 42.080 55.770 42.340 55.910 ;
        RECT 43.580 55.880 43.760 55.940 ;
        RECT 44.700 55.790 45.030 55.960 ;
        RECT 40.540 55.460 40.870 55.720 ;
        RECT 42.080 55.600 43.260 55.770 ;
        RECT 42.080 55.460 42.340 55.600 ;
        RECT 16.750 55.420 17.240 55.450 ;
        RECT 16.750 55.390 16.920 55.420 ;
        RECT 38.510 55.320 38.680 55.380 ;
        RECT 15.460 55.280 15.890 55.300 ;
        RECT 15.440 55.110 15.890 55.280 ;
        RECT 15.460 55.090 15.890 55.110 ;
        RECT 38.480 55.100 38.700 55.320 ;
        RECT 39.030 55.280 39.360 55.460 ;
        RECT 39.610 55.290 41.770 55.460 ;
        RECT 42.010 55.290 42.340 55.460 ;
        RECT 42.170 55.240 42.340 55.290 ;
        RECT 42.630 55.100 42.840 55.430 ;
        RECT 43.080 55.160 43.260 55.600 ;
        RECT 44.780 55.540 45.030 55.790 ;
        RECT 44.780 55.440 45.250 55.540 ;
        RECT 46.500 55.520 46.680 55.980 ;
        RECT 44.610 55.430 45.250 55.440 ;
        RECT 43.810 55.370 45.250 55.430 ;
        RECT 43.810 55.260 45.170 55.370 ;
        RECT 45.720 55.350 46.680 55.520 ;
        RECT 80.910 55.250 81.150 55.580 ;
        RECT 38.510 55.050 38.680 55.100 ;
        RECT 80.940 54.960 81.140 55.250 ;
        RECT 80.950 54.950 81.140 54.960 ;
        RECT 15.620 54.780 15.940 54.820 ;
        RECT 80.570 54.780 80.780 54.790 ;
        RECT 15.620 54.760 15.950 54.780 ;
        RECT 15.620 54.560 16.240 54.760 ;
        RECT 16.070 54.430 16.240 54.560 ;
        RECT 16.750 54.720 16.920 54.760 ;
        RECT 16.750 54.680 17.240 54.720 ;
        RECT 16.750 54.490 17.250 54.680 ;
        RECT 16.750 54.460 17.240 54.490 ;
        RECT 16.750 54.430 16.920 54.460 ;
        RECT 15.460 54.320 15.890 54.340 ;
        RECT 15.440 54.150 15.890 54.320 ;
        RECT 80.570 54.200 80.790 54.780 ;
        RECT 81.340 54.450 81.510 56.060 ;
        RECT 82.170 55.790 82.340 56.150 ;
        RECT 82.760 56.060 83.110 56.230 ;
        RECT 83.300 56.210 83.490 56.260 ;
        RECT 84.200 56.230 84.370 56.800 ;
        RECT 88.480 56.570 88.670 56.970 ;
        RECT 102.570 56.570 102.760 56.970 ;
        RECT 106.790 56.800 107.130 56.970 ;
        RECT 108.150 56.800 108.480 56.970 ;
        RECT 108.900 56.880 109.070 57.790 ;
        RECT 109.730 56.970 109.900 58.580 ;
        RECT 110.450 58.250 110.670 58.830 ;
        RECT 110.460 58.240 110.670 58.250 ;
        RECT 110.100 58.070 110.290 58.080 ;
        RECT 110.100 57.780 110.300 58.070 ;
        RECT 110.090 57.450 110.330 57.780 ;
        RECT 88.480 56.560 88.860 56.570 ;
        RECT 85.120 56.380 88.860 56.560 ;
        RECT 88.480 56.340 88.860 56.380 ;
        RECT 102.380 56.560 102.760 56.570 ;
        RECT 102.380 56.380 106.120 56.560 ;
        RECT 102.380 56.340 102.760 56.380 ;
        RECT 83.300 56.200 83.530 56.210 ;
        RECT 84.110 56.200 84.450 56.230 ;
        RECT 83.300 56.060 84.450 56.200 ;
        RECT 82.840 55.850 83.030 56.060 ;
        RECT 83.300 56.030 84.280 56.060 ;
        RECT 83.440 56.000 84.280 56.030 ;
        RECT 88.480 55.960 88.670 56.340 ;
        RECT 81.930 55.750 82.340 55.790 ;
        RECT 81.920 55.560 82.340 55.750 ;
        RECT 90.720 55.670 91.270 56.100 ;
        RECT 99.970 55.670 100.520 56.100 ;
        RECT 102.570 55.960 102.760 56.340 ;
        RECT 108.230 56.230 108.400 56.800 ;
        RECT 109.730 56.780 109.910 56.970 ;
        RECT 106.790 56.060 107.130 56.230 ;
        RECT 108.150 56.060 108.480 56.230 ;
        RECT 107.270 55.660 107.590 55.690 ;
        RECT 108.080 55.670 108.250 55.720 ;
        RECT 108.900 55.690 109.070 56.150 ;
        RECT 109.730 56.060 109.910 56.250 ;
        RECT 81.930 55.530 82.340 55.560 ;
        RECT 82.170 54.460 82.340 55.530 ;
        RECT 82.760 55.340 85.690 55.440 ;
        RECT 82.760 55.270 85.750 55.340 ;
        RECT 84.780 54.950 84.950 55.010 ;
        RECT 84.760 54.740 84.970 54.950 ;
        RECT 83.290 54.650 83.480 54.680 ;
        RECT 84.780 54.670 84.950 54.740 ;
        RECT 85.520 54.650 85.750 55.270 ;
        RECT 103.600 54.650 103.830 55.380 ;
        RECT 106.050 55.320 106.220 55.600 ;
        RECT 107.270 55.470 107.600 55.660 ;
        RECT 108.080 55.520 108.640 55.670 ;
        RECT 106.050 55.280 106.260 55.320 ;
        RECT 106.050 55.260 106.280 55.280 ;
        RECT 106.780 55.270 107.130 55.440 ;
        RECT 107.270 55.430 107.590 55.470 ;
        RECT 107.400 55.270 107.570 55.430 ;
        RECT 108.010 55.410 108.640 55.520 ;
        RECT 108.840 55.660 109.160 55.690 ;
        RECT 108.840 55.470 109.170 55.660 ;
        RECT 109.410 55.520 109.600 55.550 ;
        RECT 109.730 55.520 109.900 56.060 ;
        RECT 110.130 55.580 110.300 55.610 ;
        RECT 108.840 55.430 109.160 55.470 ;
        RECT 108.010 55.350 108.480 55.410 ;
        RECT 108.150 55.270 108.480 55.350 ;
        RECT 108.900 55.290 109.070 55.430 ;
        RECT 109.410 55.390 109.900 55.520 ;
        RECT 106.050 55.240 106.310 55.260 ;
        RECT 106.050 55.190 106.390 55.240 ;
        RECT 106.050 55.130 106.540 55.190 ;
        RECT 106.050 55.100 106.560 55.130 ;
        RECT 106.090 55.070 106.560 55.100 ;
        RECT 106.220 55.020 106.560 55.070 ;
        RECT 106.340 55.010 106.560 55.020 ;
        RECT 106.350 54.980 106.560 55.010 ;
        RECT 106.370 54.900 106.560 54.980 ;
        RECT 107.500 54.900 107.680 55.240 ;
        RECT 107.730 54.900 108.060 55.020 ;
        RECT 108.230 54.980 108.560 55.150 ;
        RECT 108.740 55.030 109.070 55.290 ;
        RECT 109.320 55.130 109.900 55.390 ;
        RECT 110.090 55.430 110.330 55.580 ;
        RECT 110.090 55.250 110.690 55.430 ;
        RECT 109.550 55.100 109.900 55.130 ;
        RECT 108.310 54.900 108.560 54.980 ;
        RECT 108.900 54.900 109.070 55.030 ;
        RECT 109.730 54.930 109.900 55.100 ;
        RECT 110.100 54.950 110.690 55.250 ;
        RECT 111.510 55.310 112.090 55.480 ;
        RECT 111.510 55.210 111.900 55.310 ;
        RECT 111.510 55.180 111.890 55.210 ;
        RECT 111.510 55.030 111.870 55.180 ;
        RECT 110.130 54.930 110.690 54.950 ;
        RECT 105.880 54.850 106.050 54.870 ;
        RECT 82.760 54.480 83.480 54.650 ;
        RECT 83.290 54.450 83.480 54.480 ;
        RECT 83.650 54.480 84.460 54.650 ;
        RECT 80.570 54.170 80.780 54.200 ;
        RECT 15.460 54.130 15.890 54.150 ;
        RECT 15.620 53.820 15.940 53.860 ;
        RECT 80.580 53.820 80.780 54.170 ;
        RECT 82.860 54.140 83.050 54.170 ;
        RECT 83.650 54.140 83.840 54.480 ;
        RECT 105.860 54.420 106.070 54.850 ;
        RECT 106.370 54.730 106.890 54.900 ;
        RECT 107.240 54.780 109.140 54.900 ;
        RECT 109.730 54.890 110.690 54.930 ;
        RECT 107.240 54.740 109.310 54.780 ;
        RECT 109.520 54.740 110.690 54.890 ;
        RECT 111.160 54.860 111.870 55.030 ;
        RECT 107.240 54.730 110.690 54.740 ;
        RECT 106.370 54.700 106.560 54.730 ;
        RECT 107.240 54.720 110.060 54.730 ;
        RECT 106.780 54.480 107.130 54.650 ;
        RECT 107.500 54.310 107.680 54.720 ;
        RECT 108.310 54.650 108.790 54.720 ;
        RECT 108.150 54.580 108.790 54.650 ;
        RECT 108.150 54.480 108.480 54.580 ;
        RECT 107.380 54.280 107.700 54.310 ;
        RECT 82.060 53.900 82.590 54.070 ;
        RECT 82.860 53.960 83.840 54.140 ;
        RECT 82.860 53.940 83.050 53.960 ;
        RECT 15.620 53.800 15.950 53.820 ;
        RECT 15.620 53.600 16.240 53.800 ;
        RECT 16.070 53.470 16.240 53.600 ;
        RECT 16.750 53.760 16.920 53.800 ;
        RECT 105.860 53.780 106.070 54.210 ;
        RECT 107.380 54.090 107.710 54.280 ;
        RECT 107.380 54.050 107.700 54.090 ;
        RECT 106.370 53.900 106.560 53.930 ;
        RECT 107.500 53.910 107.680 54.050 ;
        RECT 108.310 53.910 108.480 54.480 ;
        RECT 108.900 54.460 109.070 54.720 ;
        RECT 109.140 54.700 110.060 54.720 ;
        RECT 109.140 54.480 109.900 54.700 ;
        RECT 109.140 54.450 109.310 54.480 ;
        RECT 109.550 54.450 109.900 54.480 ;
        RECT 109.550 54.440 109.750 54.450 ;
        RECT 110.140 54.440 110.690 54.730 ;
        RECT 110.450 54.200 110.670 54.440 ;
        RECT 110.460 54.170 110.670 54.200 ;
        RECT 108.650 53.940 109.180 54.070 ;
        RECT 110.460 53.950 110.660 54.170 ;
        RECT 111.160 54.110 111.860 54.420 ;
        RECT 108.650 53.910 109.310 53.940 ;
        RECT 109.550 53.910 109.750 53.950 ;
        RECT 109.870 53.910 110.060 53.930 ;
        RECT 107.240 53.900 110.060 53.910 ;
        RECT 110.140 53.900 110.690 53.950 ;
        RECT 105.880 53.760 106.050 53.780 ;
        RECT 16.750 53.720 17.240 53.760 ;
        RECT 106.370 53.730 106.890 53.900 ;
        RECT 107.240 53.740 110.690 53.900 ;
        RECT 111.010 53.880 111.860 54.110 ;
        RECT 107.240 53.730 109.750 53.740 ;
        RECT 16.750 53.530 17.250 53.720 ;
        RECT 106.370 53.650 106.560 53.730 ;
        RECT 106.350 53.620 106.560 53.650 ;
        RECT 106.340 53.610 106.560 53.620 ;
        RECT 106.220 53.560 106.560 53.610 ;
        RECT 106.090 53.530 106.560 53.560 ;
        RECT 16.750 53.500 17.240 53.530 ;
        RECT 106.050 53.500 106.560 53.530 ;
        RECT 16.750 53.470 16.920 53.500 ;
        RECT 15.460 53.360 15.890 53.380 ;
        RECT 15.440 53.190 15.890 53.360 ;
        RECT 15.460 53.170 15.890 53.190 ;
        RECT 17.250 53.130 17.670 53.300 ;
        RECT 17.350 53.090 17.580 53.130 ;
        RECT 58.470 53.060 58.640 53.480 ;
        RECT 59.280 53.360 59.520 53.390 ;
        RECT 58.950 53.190 59.520 53.360 ;
        RECT 59.760 53.190 61.100 53.360 ;
        RECT 61.550 53.190 62.510 53.360 ;
        RECT 59.280 53.150 59.520 53.190 ;
        RECT 62.060 53.180 62.230 53.190 ;
        RECT 58.400 52.840 58.570 52.880 ;
        RECT 38.510 52.700 38.680 52.750 ;
        RECT 38.480 52.480 38.700 52.700 ;
        RECT 38.510 52.420 38.680 52.480 ;
        RECT 39.030 52.340 39.360 52.520 ;
        RECT 42.170 52.510 42.340 52.560 ;
        RECT 39.610 52.340 41.770 52.510 ;
        RECT 42.010 52.340 42.340 52.510 ;
        RECT 42.630 52.370 42.840 52.700 ;
        RECT 58.340 52.670 58.570 52.840 ;
        RECT 39.060 51.900 39.330 52.340 ;
        RECT 40.540 52.080 40.870 52.340 ;
        RECT 42.080 52.200 42.340 52.340 ;
        RECT 43.080 52.200 43.260 52.640 ;
        RECT 43.810 52.430 45.170 52.540 ;
        RECT 43.810 52.370 45.250 52.430 ;
        RECT 44.610 52.360 45.250 52.370 ;
        RECT 39.100 51.890 39.330 51.900 ;
        RECT 42.080 52.030 43.260 52.200 ;
        RECT 44.780 52.260 45.250 52.360 ;
        RECT 45.720 52.280 46.680 52.450 ;
        RECT 58.400 52.320 58.570 52.670 ;
        RECT 58.740 52.740 58.930 52.760 ;
        RECT 61.740 52.740 62.070 52.920 ;
        RECT 58.740 52.570 59.300 52.740 ;
        RECT 59.760 52.570 62.510 52.740 ;
        RECT 58.740 52.530 58.930 52.570 ;
        RECT 63.040 52.500 63.210 53.430 ;
        RECT 63.440 52.630 63.610 53.480 ;
        RECT 106.050 53.440 106.540 53.500 ;
        RECT 106.050 53.390 106.390 53.440 ;
        RECT 106.050 53.370 106.310 53.390 ;
        RECT 106.050 53.350 106.280 53.370 ;
        RECT 107.500 53.360 107.680 53.730 ;
        RECT 107.730 53.610 108.060 53.730 ;
        RECT 80.580 52.830 80.780 53.180 ;
        RECT 82.060 52.930 82.590 53.100 ;
        RECT 80.570 52.800 80.780 52.830 ;
        RECT 42.080 51.890 42.340 52.030 ;
        RECT 44.780 52.010 45.030 52.260 ;
        RECT 39.100 51.720 39.860 51.890 ;
        RECT 40.110 51.720 41.280 51.890 ;
        RECT 41.520 51.860 42.340 51.890 ;
        RECT 43.580 51.860 43.760 51.920 ;
        RECT 41.520 51.720 42.630 51.860 ;
        RECT 40.510 51.620 40.860 51.720 ;
        RECT 42.170 51.690 42.630 51.720 ;
        RECT 43.080 51.690 43.760 51.860 ;
        RECT 44.700 51.840 45.030 52.010 ;
        RECT 46.500 51.820 46.680 52.280 ;
        RECT 80.570 52.220 80.790 52.800 ;
        RECT 80.570 52.210 80.780 52.220 ;
        RECT 43.120 51.670 43.760 51.690 ;
        RECT 43.580 51.660 43.760 51.670 ;
        RECT 45.360 51.660 45.960 51.810 ;
        RECT 43.580 51.640 45.960 51.660 ;
        RECT 46.420 51.650 46.750 51.820 ;
        RECT 58.400 51.730 58.570 52.080 ;
        RECT 80.950 52.040 81.140 52.050 ;
        RECT 43.580 51.490 45.810 51.640 ;
        RECT 58.340 51.560 58.570 51.730 ;
        RECT 58.740 51.830 58.930 51.870 ;
        RECT 58.740 51.660 59.300 51.830 ;
        RECT 59.760 51.660 62.510 51.830 ;
        RECT 58.740 51.640 58.930 51.660 ;
        RECT 58.400 51.520 58.570 51.560 ;
        RECT 61.740 51.480 62.070 51.660 ;
        RECT 38.510 51.150 38.680 51.200 ;
        RECT 38.480 50.930 38.700 51.150 ;
        RECT 38.510 50.870 38.680 50.930 ;
        RECT 39.030 50.790 39.360 50.970 ;
        RECT 42.170 50.960 42.340 51.010 ;
        RECT 39.610 50.790 41.770 50.960 ;
        RECT 42.010 50.790 42.340 50.960 ;
        RECT 42.630 50.820 42.840 51.150 ;
        RECT 39.060 50.350 39.330 50.790 ;
        RECT 40.540 50.530 40.870 50.790 ;
        RECT 42.080 50.650 42.340 50.790 ;
        RECT 43.080 50.650 43.260 51.090 ;
        RECT 43.810 50.880 45.170 50.990 ;
        RECT 58.470 50.920 58.640 51.340 ;
        RECT 59.280 51.210 59.520 51.250 ;
        RECT 62.060 51.210 62.230 51.220 ;
        RECT 58.950 51.040 59.520 51.210 ;
        RECT 59.760 51.040 61.100 51.210 ;
        RECT 61.550 51.040 62.510 51.210 ;
        RECT 59.280 51.010 59.520 51.040 ;
        RECT 63.040 50.970 63.210 51.900 ;
        RECT 63.440 50.920 63.610 51.770 ;
        RECT 80.940 51.750 81.140 52.040 ;
        RECT 80.910 51.420 81.150 51.750 ;
        RECT 81.340 50.940 81.510 52.550 ;
        RECT 43.810 50.820 45.250 50.880 ;
        RECT 44.610 50.810 45.250 50.820 ;
        RECT 39.100 50.340 39.330 50.350 ;
        RECT 42.080 50.480 43.260 50.650 ;
        RECT 44.780 50.710 45.250 50.810 ;
        RECT 45.720 50.730 46.680 50.900 ;
        RECT 81.330 50.750 81.510 50.940 ;
        RECT 82.170 52.020 82.340 52.540 ;
        RECT 82.760 52.350 83.090 52.520 ;
        RECT 84.110 52.350 84.460 52.520 ;
        RECT 84.780 52.500 89.840 53.330 ;
        RECT 106.050 53.310 106.260 53.350 ;
        RECT 106.050 53.030 106.220 53.310 ;
        RECT 107.400 53.200 107.680 53.360 ;
        RECT 108.310 53.320 108.480 53.730 ;
        RECT 109.140 53.650 109.750 53.730 ;
        RECT 109.870 53.700 110.690 53.740 ;
        RECT 109.140 53.610 109.310 53.650 ;
        RECT 109.550 53.620 109.750 53.650 ;
        RECT 108.280 53.290 108.480 53.320 ;
        RECT 108.260 53.280 108.480 53.290 ;
        RECT 107.270 52.940 107.680 53.200 ;
        RECT 108.010 53.200 108.480 53.280 ;
        RECT 108.900 53.200 109.070 53.360 ;
        RECT 109.410 53.290 109.600 53.310 ;
        RECT 109.410 53.280 109.750 53.290 ;
        RECT 109.410 53.260 109.850 53.280 ;
        RECT 108.010 53.110 108.470 53.200 ;
        RECT 108.280 53.090 108.470 53.110 ;
        RECT 108.840 53.160 109.160 53.200 ;
        RECT 108.840 53.100 109.170 53.160 ;
        RECT 109.320 53.110 109.850 53.260 ;
        RECT 107.500 52.670 107.680 52.940 ;
        RECT 108.110 53.000 108.430 53.030 ;
        RECT 108.110 52.810 108.440 53.000 ;
        RECT 108.650 52.930 109.180 53.100 ;
        RECT 109.320 53.000 109.750 53.110 ;
        RECT 110.130 53.020 110.690 53.700 ;
        RECT 111.160 53.540 111.860 53.880 ;
        RECT 111.620 53.180 111.940 53.220 ;
        RECT 111.620 53.120 111.950 53.180 ;
        RECT 109.550 52.960 109.750 53.000 ;
        RECT 110.140 52.960 110.690 53.020 ;
        RECT 111.150 52.990 111.950 53.120 ;
        RECT 111.150 52.960 111.940 52.990 ;
        RECT 110.460 52.830 110.660 52.960 ;
        RECT 111.150 52.940 111.850 52.960 ;
        RECT 108.110 52.770 108.430 52.810 ;
        RECT 110.460 52.800 110.670 52.830 ;
        RECT 108.110 52.690 108.280 52.770 ;
        RECT 89.290 52.420 89.770 52.500 ;
        RECT 82.170 51.760 82.500 52.020 ;
        RECT 82.170 50.850 82.340 51.760 ;
        RECT 82.760 51.560 83.090 51.730 ;
        RECT 84.110 51.560 84.460 51.730 ;
        RECT 87.410 51.560 87.640 52.250 ;
        RECT 89.290 52.170 89.760 52.420 ;
        RECT 106.050 52.300 106.220 52.580 ;
        RECT 106.780 52.350 107.130 52.520 ;
        RECT 107.270 52.410 107.680 52.670 ;
        RECT 108.060 52.520 108.280 52.690 ;
        RECT 108.840 52.640 109.160 52.670 ;
        RECT 108.060 52.500 108.480 52.520 ;
        RECT 106.050 52.260 106.260 52.300 ;
        RECT 90.720 51.370 91.270 51.800 ;
        RECT 99.970 51.370 100.520 51.800 ;
        RECT 103.600 51.560 103.830 52.250 ;
        RECT 106.050 52.240 106.280 52.260 ;
        RECT 107.400 52.250 107.680 52.410 ;
        RECT 108.010 52.350 108.480 52.500 ;
        RECT 108.840 52.450 109.170 52.640 ;
        RECT 109.410 52.500 109.600 52.530 ;
        RECT 109.730 52.500 109.900 52.550 ;
        RECT 108.840 52.410 109.160 52.450 ;
        RECT 109.410 52.430 109.900 52.500 ;
        RECT 108.010 52.330 108.470 52.350 ;
        RECT 108.260 52.320 108.470 52.330 ;
        RECT 108.280 52.290 108.470 52.320 ;
        RECT 106.050 52.220 106.310 52.240 ;
        RECT 106.050 52.170 106.390 52.220 ;
        RECT 106.050 52.110 106.540 52.170 ;
        RECT 106.050 52.080 106.560 52.110 ;
        RECT 106.090 52.050 106.560 52.080 ;
        RECT 106.220 52.000 106.560 52.050 ;
        RECT 106.340 51.990 106.560 52.000 ;
        RECT 106.350 51.960 106.560 51.990 ;
        RECT 106.370 51.880 106.560 51.960 ;
        RECT 107.500 51.880 107.680 52.250 ;
        RECT 108.590 52.100 108.780 52.220 ;
        RECT 108.230 52.020 108.780 52.100 ;
        RECT 108.900 52.020 109.070 52.410 ;
        RECT 109.320 52.170 109.900 52.430 ;
        RECT 109.550 52.140 109.900 52.170 ;
        RECT 107.730 51.880 108.060 52.000 ;
        RECT 108.230 51.930 109.070 52.020 ;
        RECT 108.310 51.880 108.480 51.930 ;
        RECT 108.740 51.880 109.070 51.930 ;
        RECT 109.730 51.910 109.900 52.140 ;
        RECT 110.130 52.470 110.300 52.590 ;
        RECT 110.450 52.470 110.670 52.800 ;
        RECT 110.130 52.050 110.690 52.470 ;
        RECT 111.610 52.460 111.930 52.500 ;
        RECT 111.150 52.280 111.940 52.460 ;
        RECT 111.610 52.270 111.940 52.280 ;
        RECT 111.610 52.240 111.930 52.270 ;
        RECT 110.100 51.910 110.690 52.050 ;
        RECT 105.880 51.830 106.050 51.850 ;
        RECT 105.860 51.400 106.070 51.830 ;
        RECT 106.370 51.730 106.890 51.880 ;
        RECT 107.240 51.820 109.140 51.880 ;
        RECT 109.730 51.870 110.690 51.910 ;
        RECT 107.240 51.780 109.310 51.820 ;
        RECT 109.520 51.780 110.690 51.870 ;
        RECT 106.370 51.710 107.130 51.730 ;
        RECT 106.370 51.680 106.560 51.710 ;
        RECT 106.780 51.560 107.130 51.710 ;
        RECT 107.240 51.710 110.690 51.780 ;
        RECT 107.240 51.700 110.060 51.710 ;
        RECT 82.760 50.770 83.090 50.940 ;
        RECT 84.110 50.770 84.450 50.940 ;
        RECT 42.080 50.340 42.340 50.480 ;
        RECT 44.780 50.460 45.030 50.710 ;
        RECT 39.100 50.170 39.860 50.340 ;
        RECT 40.110 50.170 41.280 50.340 ;
        RECT 41.520 50.310 42.340 50.340 ;
        RECT 43.580 50.310 43.760 50.370 ;
        RECT 41.520 50.170 42.630 50.310 ;
        RECT 40.510 50.070 40.860 50.170 ;
        RECT 42.170 50.140 42.630 50.170 ;
        RECT 43.080 50.140 43.760 50.310 ;
        RECT 44.700 50.290 45.030 50.460 ;
        RECT 46.500 50.270 46.680 50.730 ;
        RECT 43.120 50.120 43.760 50.140 ;
        RECT 43.580 50.110 43.760 50.120 ;
        RECT 45.360 50.110 45.960 50.260 ;
        RECT 43.580 50.090 45.960 50.110 ;
        RECT 46.420 50.100 46.750 50.270 ;
        RECT 58.470 50.130 58.640 50.550 ;
        RECT 59.280 50.430 59.520 50.460 ;
        RECT 58.950 50.260 59.520 50.430 ;
        RECT 59.760 50.260 61.100 50.430 ;
        RECT 61.550 50.260 62.510 50.430 ;
        RECT 59.280 50.220 59.520 50.260 ;
        RECT 62.060 50.250 62.230 50.260 ;
        RECT 43.580 49.940 45.810 50.090 ;
        RECT 58.400 49.910 58.570 49.950 ;
        RECT 58.340 49.740 58.570 49.910 ;
        RECT 38.510 49.600 38.680 49.650 ;
        RECT 38.480 49.380 38.700 49.600 ;
        RECT 38.510 49.320 38.680 49.380 ;
        RECT 39.030 49.240 39.360 49.420 ;
        RECT 42.170 49.410 42.340 49.460 ;
        RECT 39.610 49.240 41.770 49.410 ;
        RECT 42.010 49.240 42.340 49.410 ;
        RECT 42.630 49.270 42.840 49.600 ;
        RECT 39.060 48.800 39.330 49.240 ;
        RECT 40.540 48.980 40.870 49.240 ;
        RECT 42.080 49.100 42.340 49.240 ;
        RECT 43.080 49.100 43.260 49.540 ;
        RECT 43.810 49.330 45.170 49.440 ;
        RECT 58.400 49.390 58.570 49.740 ;
        RECT 58.740 49.810 58.930 49.830 ;
        RECT 61.740 49.810 62.070 49.990 ;
        RECT 58.740 49.640 59.300 49.810 ;
        RECT 59.760 49.640 62.510 49.810 ;
        RECT 58.740 49.600 58.930 49.640 ;
        RECT 63.040 49.570 63.210 50.500 ;
        RECT 63.440 49.700 63.610 50.550 ;
        RECT 81.330 50.030 81.510 50.220 ;
        RECT 82.840 50.200 83.010 50.770 ;
        RECT 88.480 50.540 88.670 50.940 ;
        RECT 102.570 50.540 102.760 50.940 ;
        RECT 105.860 50.760 106.070 51.190 ;
        RECT 106.370 50.880 106.560 50.910 ;
        RECT 106.790 50.880 107.130 50.940 ;
        RECT 107.500 50.890 107.680 51.700 ;
        RECT 108.150 51.560 108.480 51.700 ;
        RECT 108.310 50.940 108.480 51.560 ;
        RECT 108.150 50.890 108.480 50.940 ;
        RECT 108.900 50.890 109.070 51.700 ;
        RECT 109.140 51.680 110.060 51.700 ;
        RECT 109.140 51.520 109.900 51.680 ;
        RECT 109.140 51.490 109.310 51.520 ;
        RECT 109.550 51.480 109.900 51.520 ;
        RECT 109.730 50.990 109.900 51.480 ;
        RECT 110.090 51.480 110.690 51.710 ;
        RECT 111.160 51.520 111.860 51.860 ;
        RECT 110.090 51.420 110.330 51.480 ;
        RECT 111.010 51.290 111.860 51.520 ;
        RECT 109.140 50.950 109.310 50.980 ;
        RECT 109.550 50.950 109.900 50.990 ;
        RECT 109.140 50.940 109.900 50.950 ;
        RECT 109.140 50.910 109.910 50.940 ;
        RECT 109.140 50.890 110.060 50.910 ;
        RECT 106.370 50.770 107.130 50.880 ;
        RECT 107.240 50.880 110.060 50.890 ;
        RECT 110.140 50.880 110.690 50.990 ;
        RECT 111.160 50.980 111.860 51.290 ;
        RECT 105.880 50.740 106.050 50.760 ;
        RECT 106.370 50.710 106.890 50.770 ;
        RECT 107.240 50.720 110.690 50.880 ;
        RECT 107.240 50.710 109.750 50.720 ;
        RECT 106.370 50.630 106.560 50.710 ;
        RECT 106.350 50.600 106.560 50.630 ;
        RECT 106.340 50.590 106.560 50.600 ;
        RECT 106.220 50.540 106.560 50.590 ;
        RECT 88.480 50.530 88.860 50.540 ;
        RECT 85.120 50.350 88.860 50.530 ;
        RECT 88.480 50.310 88.860 50.350 ;
        RECT 102.380 50.530 102.760 50.540 ;
        RECT 106.090 50.530 106.560 50.540 ;
        RECT 102.380 50.480 106.560 50.530 ;
        RECT 102.380 50.420 106.540 50.480 ;
        RECT 102.380 50.370 106.390 50.420 ;
        RECT 102.380 50.350 106.310 50.370 ;
        RECT 102.380 50.310 102.760 50.350 ;
        RECT 43.810 49.270 45.250 49.330 ;
        RECT 44.610 49.260 45.250 49.270 ;
        RECT 39.100 48.790 39.330 48.800 ;
        RECT 42.080 48.930 43.260 49.100 ;
        RECT 44.780 49.160 45.250 49.260 ;
        RECT 45.720 49.180 46.680 49.350 ;
        RECT 80.910 49.220 81.150 49.550 ;
        RECT 42.080 48.790 42.340 48.930 ;
        RECT 44.780 48.910 45.030 49.160 ;
        RECT 39.100 48.620 39.860 48.790 ;
        RECT 40.110 48.620 41.280 48.790 ;
        RECT 41.520 48.760 42.340 48.790 ;
        RECT 43.580 48.760 43.760 48.820 ;
        RECT 41.520 48.620 42.630 48.760 ;
        RECT 40.510 48.520 40.860 48.620 ;
        RECT 42.170 48.590 42.630 48.620 ;
        RECT 43.080 48.590 43.760 48.760 ;
        RECT 44.700 48.740 45.030 48.910 ;
        RECT 46.500 48.720 46.680 49.180 ;
        RECT 58.400 48.800 58.570 49.150 ;
        RECT 43.120 48.570 43.760 48.590 ;
        RECT 43.580 48.560 43.760 48.570 ;
        RECT 45.360 48.560 45.960 48.710 ;
        RECT 43.580 48.540 45.960 48.560 ;
        RECT 46.420 48.550 46.750 48.720 ;
        RECT 58.340 48.630 58.570 48.800 ;
        RECT 58.740 48.900 58.930 48.940 ;
        RECT 58.740 48.730 59.300 48.900 ;
        RECT 59.760 48.730 62.510 48.900 ;
        RECT 58.740 48.710 58.930 48.730 ;
        RECT 58.400 48.590 58.570 48.630 ;
        RECT 61.740 48.550 62.070 48.730 ;
        RECT 43.580 48.390 45.810 48.540 ;
        RECT 38.510 48.050 38.680 48.100 ;
        RECT 38.480 47.830 38.700 48.050 ;
        RECT 38.510 47.770 38.680 47.830 ;
        RECT 39.030 47.690 39.360 47.870 ;
        RECT 42.170 47.860 42.340 47.910 ;
        RECT 39.610 47.690 41.770 47.860 ;
        RECT 42.010 47.690 42.340 47.860 ;
        RECT 42.630 47.720 42.840 48.050 ;
        RECT 58.470 47.990 58.640 48.410 ;
        RECT 59.280 48.280 59.520 48.320 ;
        RECT 62.060 48.280 62.230 48.290 ;
        RECT 58.950 48.110 59.520 48.280 ;
        RECT 59.760 48.110 61.100 48.280 ;
        RECT 61.550 48.110 62.510 48.280 ;
        RECT 59.280 48.080 59.520 48.110 ;
        RECT 63.040 48.040 63.210 48.970 ;
        RECT 80.940 48.930 81.140 49.220 ;
        RECT 80.950 48.920 81.140 48.930 ;
        RECT 63.440 47.990 63.610 48.840 ;
        RECT 80.570 48.750 80.780 48.760 ;
        RECT 80.570 48.170 80.790 48.750 ;
        RECT 81.340 48.420 81.510 50.030 ;
        RECT 82.170 49.260 82.340 50.120 ;
        RECT 82.760 50.030 83.090 50.200 ;
        RECT 84.110 50.030 84.450 50.200 ;
        RECT 88.480 49.930 88.670 50.310 ;
        RECT 90.720 49.640 91.270 50.070 ;
        RECT 99.970 49.640 100.520 50.070 ;
        RECT 102.570 49.930 102.760 50.310 ;
        RECT 106.050 50.330 106.280 50.350 ;
        RECT 107.500 50.340 107.680 50.710 ;
        RECT 107.730 50.590 108.060 50.710 ;
        RECT 106.050 50.290 106.260 50.330 ;
        RECT 106.050 50.010 106.220 50.290 ;
        RECT 106.790 50.030 107.130 50.200 ;
        RECT 107.400 50.180 107.680 50.340 ;
        RECT 108.230 50.260 108.480 50.710 ;
        RECT 109.140 50.690 109.750 50.710 ;
        RECT 109.140 50.650 109.310 50.690 ;
        RECT 109.550 50.660 109.750 50.690 ;
        RECT 109.870 50.680 110.690 50.720 ;
        RECT 107.270 50.140 107.680 50.180 ;
        RECT 107.270 49.950 107.600 50.140 ;
        RECT 108.010 50.090 108.480 50.260 ;
        RECT 108.900 50.180 109.070 50.340 ;
        RECT 109.550 50.300 109.750 50.330 ;
        RECT 109.320 50.260 109.750 50.300 ;
        RECT 109.320 50.220 109.850 50.260 ;
        RECT 108.150 50.030 108.480 50.090 ;
        RECT 108.840 50.140 109.160 50.180 ;
        RECT 108.840 49.950 109.170 50.140 ;
        RECT 109.320 50.040 109.910 50.220 ;
        RECT 109.550 50.030 109.910 50.040 ;
        RECT 109.550 50.000 109.900 50.030 ;
        RECT 110.130 50.000 110.690 50.680 ;
        RECT 111.160 50.370 111.870 50.540 ;
        RECT 111.510 50.090 111.870 50.370 ;
        RECT 107.270 49.920 107.590 49.950 ;
        RECT 108.840 49.920 109.160 49.950 ;
        RECT 108.080 49.640 108.250 49.690 ;
        RECT 82.170 49.000 82.500 49.260 ;
        RECT 82.760 49.240 83.090 49.410 ;
        RECT 84.110 49.240 84.460 49.410 ;
        RECT 82.170 48.430 82.340 49.000 ;
        RECT 87.410 48.620 87.640 49.350 ;
        RECT 82.760 48.450 83.090 48.620 ;
        RECT 84.110 48.450 84.460 48.620 ;
        RECT 89.450 48.490 89.790 48.740 ;
        RECT 103.600 48.620 103.830 49.350 ;
        RECT 106.780 49.240 107.130 49.410 ;
        RECT 108.080 49.380 108.640 49.640 ;
        RECT 108.080 49.360 108.480 49.380 ;
        RECT 108.150 49.240 108.480 49.360 ;
        RECT 108.900 49.260 109.070 49.920 ;
        RECT 109.730 49.400 109.900 50.000 ;
        RECT 111.510 49.920 112.090 50.090 ;
        RECT 109.550 49.360 109.900 49.400 ;
        RECT 89.450 48.410 89.800 48.490 ;
        RECT 106.780 48.450 107.130 48.620 ;
        RECT 80.570 48.140 80.780 48.170 ;
        RECT 39.060 47.250 39.330 47.690 ;
        RECT 40.540 47.430 40.870 47.690 ;
        RECT 42.080 47.550 42.340 47.690 ;
        RECT 43.080 47.550 43.260 47.990 ;
        RECT 43.810 47.780 45.170 47.890 ;
        RECT 43.810 47.720 45.250 47.780 ;
        RECT 44.610 47.710 45.250 47.720 ;
        RECT 39.100 47.240 39.330 47.250 ;
        RECT 42.080 47.380 43.260 47.550 ;
        RECT 44.780 47.610 45.250 47.710 ;
        RECT 45.720 47.630 46.680 47.800 ;
        RECT 80.580 47.790 80.780 48.140 ;
        RECT 82.060 47.870 82.590 48.040 ;
        RECT 42.080 47.240 42.340 47.380 ;
        RECT 44.780 47.360 45.030 47.610 ;
        RECT 39.100 47.070 39.860 47.240 ;
        RECT 40.110 47.070 41.280 47.240 ;
        RECT 41.520 47.210 42.340 47.240 ;
        RECT 43.580 47.210 43.760 47.270 ;
        RECT 41.520 47.070 42.630 47.210 ;
        RECT 40.510 46.970 40.860 47.070 ;
        RECT 42.170 47.040 42.630 47.070 ;
        RECT 43.080 47.040 43.760 47.210 ;
        RECT 44.700 47.190 45.030 47.360 ;
        RECT 46.500 47.170 46.680 47.630 ;
        RECT 84.750 47.560 89.800 48.410 ;
        RECT 107.500 48.280 107.680 49.210 ;
        RECT 108.230 48.950 108.560 49.120 ;
        RECT 108.740 49.000 109.070 49.260 ;
        RECT 109.320 49.100 109.900 49.360 ;
        RECT 110.090 49.400 110.330 49.550 ;
        RECT 110.090 49.220 110.690 49.400 ;
        RECT 109.550 49.070 109.900 49.100 ;
        RECT 108.310 48.810 108.560 48.950 ;
        RECT 108.310 48.620 108.790 48.810 ;
        RECT 108.150 48.550 108.790 48.620 ;
        RECT 108.150 48.450 108.480 48.550 ;
        RECT 107.380 48.250 107.700 48.280 ;
        RECT 107.380 48.060 107.710 48.250 ;
        RECT 107.380 48.020 107.700 48.060 ;
        RECT 43.120 47.020 43.760 47.040 ;
        RECT 43.580 47.010 43.760 47.020 ;
        RECT 45.360 47.010 45.960 47.160 ;
        RECT 43.580 46.990 45.960 47.010 ;
        RECT 46.420 47.000 46.750 47.170 ;
        RECT 43.580 46.840 45.810 46.990 ;
        RECT 65.900 46.920 66.100 47.270 ;
        RECT 67.640 47.190 67.960 47.200 ;
        RECT 67.380 47.020 67.960 47.190 ;
        RECT 67.630 46.970 67.960 47.020 ;
        RECT 67.640 46.940 67.960 46.970 ;
        RECT 88.440 47.190 88.760 47.200 ;
        RECT 88.440 47.020 89.020 47.190 ;
        RECT 88.440 46.970 88.770 47.020 ;
        RECT 88.440 46.940 88.760 46.970 ;
        RECT 65.890 46.890 66.100 46.920 ;
        RECT 90.300 46.920 90.500 47.270 ;
        RECT 65.890 46.300 66.110 46.890 ;
        RECT 66.630 46.330 66.830 46.900 ;
        RECT 67.640 46.610 67.960 46.650 ;
        RECT 67.630 46.570 67.960 46.610 ;
        RECT 67.380 46.400 67.960 46.570 ;
        RECT 67.640 46.390 67.960 46.400 ;
        RECT 88.440 46.610 88.760 46.650 ;
        RECT 88.440 46.570 88.770 46.610 ;
        RECT 88.440 46.400 89.020 46.570 ;
        RECT 88.440 46.390 88.760 46.400 ;
        RECT 65.890 45.270 66.110 45.860 ;
        RECT 68.640 45.840 68.810 46.350 ;
        RECT 72.580 45.850 72.750 46.360 ;
        RECT 83.650 45.850 83.820 46.360 ;
        RECT 87.590 45.840 87.760 46.350 ;
        RECT 89.570 46.330 89.770 46.900 ;
        RECT 90.300 46.890 90.510 46.920 ;
        RECT 90.290 46.300 90.510 46.890 ;
        RECT 92.630 46.110 92.830 47.120 ;
        RECT 98.380 46.110 98.670 47.120 ;
        RECT 65.890 45.240 66.100 45.270 ;
        RECT 66.630 45.260 66.830 45.830 ;
        RECT 67.640 45.760 67.960 45.770 ;
        RECT 67.380 45.590 67.960 45.760 ;
        RECT 67.630 45.550 67.960 45.590 ;
        RECT 67.640 45.510 67.960 45.550 ;
        RECT 88.440 45.760 88.760 45.770 ;
        RECT 88.440 45.590 89.020 45.760 ;
        RECT 88.440 45.550 88.770 45.590 ;
        RECT 88.440 45.510 88.760 45.550 ;
        RECT 89.570 45.260 89.770 45.830 ;
        RECT 90.290 45.270 90.510 45.860 ;
        RECT 65.900 44.890 66.100 45.240 ;
        RECT 90.300 45.240 90.510 45.270 ;
        RECT 67.640 45.190 67.960 45.220 ;
        RECT 67.630 45.140 67.960 45.190 ;
        RECT 88.440 45.190 88.760 45.220 ;
        RECT 67.380 44.970 67.960 45.140 ;
        RECT 67.640 44.960 67.960 44.970 ;
        RECT 66.270 44.490 66.710 44.660 ;
        RECT 65.900 43.910 66.100 44.260 ;
        RECT 67.640 44.180 67.960 44.190 ;
        RECT 67.380 44.010 67.960 44.180 ;
        RECT 67.630 43.960 67.960 44.010 ;
        RECT 68.640 44.000 68.810 45.010 ;
        RECT 70.570 44.280 71.120 44.710 ;
        RECT 72.570 44.140 72.740 45.150 ;
        RECT 74.600 44.350 75.150 44.780 ;
        RECT 81.250 44.350 81.800 44.780 ;
        RECT 83.660 44.140 83.830 45.150 ;
        RECT 88.440 45.140 88.770 45.190 ;
        RECT 85.280 44.280 85.830 44.710 ;
        RECT 87.590 44.000 87.760 45.010 ;
        RECT 88.440 44.970 89.020 45.140 ;
        RECT 88.440 44.960 88.760 44.970 ;
        RECT 90.300 44.890 90.500 45.240 ;
        RECT 89.690 44.490 90.130 44.660 ;
        RECT 88.440 44.180 88.760 44.190 ;
        RECT 88.440 44.010 89.020 44.180 ;
        RECT 67.640 43.930 67.960 43.960 ;
        RECT 88.440 43.960 88.770 44.010 ;
        RECT 88.440 43.930 88.760 43.960 ;
        RECT 65.890 43.880 66.100 43.910 ;
        RECT 90.300 43.910 90.500 44.260 ;
        RECT 107.500 44.110 107.680 48.020 ;
        RECT 108.310 47.170 108.480 48.450 ;
        RECT 108.900 48.430 109.070 49.000 ;
        RECT 109.140 48.710 109.310 48.750 ;
        RECT 109.730 48.740 109.900 49.070 ;
        RECT 110.100 48.920 110.690 49.220 ;
        RECT 111.510 49.280 112.090 49.450 ;
        RECT 111.510 49.180 111.900 49.280 ;
        RECT 111.510 49.150 111.890 49.180 ;
        RECT 111.510 49.000 111.870 49.150 ;
        RECT 109.550 48.710 109.900 48.740 ;
        RECT 109.140 48.450 109.900 48.710 ;
        RECT 109.140 48.420 109.310 48.450 ;
        RECT 109.550 48.420 109.900 48.450 ;
        RECT 109.550 48.410 109.750 48.420 ;
        RECT 110.140 48.410 110.690 48.920 ;
        RECT 111.160 48.830 111.870 49.000 ;
        RECT 110.450 48.170 110.670 48.410 ;
        RECT 110.460 48.140 110.670 48.170 ;
        RECT 108.650 47.910 109.180 48.040 ;
        RECT 110.460 47.920 110.660 48.140 ;
        RECT 111.160 48.080 111.860 48.390 ;
        RECT 108.650 47.880 109.310 47.910 ;
        RECT 109.550 47.880 109.750 47.920 ;
        RECT 108.650 47.870 109.750 47.880 ;
        RECT 109.140 47.620 109.750 47.870 ;
        RECT 109.140 47.580 109.310 47.620 ;
        RECT 109.550 47.590 109.750 47.620 ;
        RECT 109.550 47.230 109.750 47.260 ;
        RECT 108.110 46.970 108.430 47.000 ;
        RECT 109.320 46.970 109.750 47.230 ;
        RECT 108.110 46.780 108.440 46.970 ;
        RECT 109.550 46.930 109.750 46.970 ;
        RECT 110.140 46.930 110.690 47.920 ;
        RECT 111.010 47.850 111.860 48.080 ;
        RECT 111.160 47.510 111.860 47.850 ;
        RECT 111.620 47.150 111.940 47.190 ;
        RECT 111.620 47.090 111.950 47.150 ;
        RECT 111.150 46.960 111.950 47.090 ;
        RECT 111.150 46.930 111.940 46.960 ;
        RECT 111.150 46.910 111.850 46.930 ;
        RECT 108.110 46.740 108.430 46.780 ;
        RECT 108.110 46.660 108.280 46.740 ;
        RECT 108.060 46.490 108.280 46.660 ;
        RECT 108.060 46.330 108.230 46.490 ;
        RECT 109.550 46.400 109.750 46.440 ;
        RECT 108.590 46.070 108.780 46.190 ;
        RECT 109.320 46.140 109.750 46.400 ;
        RECT 109.550 46.110 109.750 46.140 ;
        RECT 108.230 45.960 108.780 46.070 ;
        RECT 108.230 45.900 108.770 45.960 ;
        RECT 108.310 44.120 108.480 45.900 ;
        RECT 109.140 45.750 109.310 45.790 ;
        RECT 109.550 45.750 109.750 45.780 ;
        RECT 109.140 45.490 109.750 45.750 ;
        RECT 109.140 45.460 109.310 45.490 ;
        RECT 109.550 45.450 109.750 45.490 ;
        RECT 110.140 45.450 110.690 46.440 ;
        RECT 111.610 46.430 111.930 46.470 ;
        RECT 111.150 46.250 111.940 46.430 ;
        RECT 111.610 46.240 111.940 46.250 ;
        RECT 111.610 46.210 111.930 46.240 ;
        RECT 111.160 45.490 111.860 45.830 ;
        RECT 111.010 45.260 111.860 45.490 ;
        RECT 109.140 44.920 109.310 44.950 ;
        RECT 109.550 44.920 109.750 44.960 ;
        RECT 109.140 44.660 109.750 44.920 ;
        RECT 109.140 44.620 109.310 44.660 ;
        RECT 109.550 44.630 109.750 44.660 ;
        RECT 109.550 44.270 109.750 44.300 ;
        RECT 109.320 44.010 109.750 44.270 ;
        RECT 109.550 43.970 109.750 44.010 ;
        RECT 110.140 43.970 110.690 44.960 ;
        RECT 111.160 44.950 111.860 45.260 ;
        RECT 111.160 44.340 111.870 44.510 ;
        RECT 111.510 44.060 111.870 44.340 ;
        RECT 58.470 42.990 58.640 43.410 ;
        RECT 59.280 43.290 59.520 43.320 ;
        RECT 58.950 43.120 59.520 43.290 ;
        RECT 59.760 43.120 61.100 43.290 ;
        RECT 61.550 43.120 62.510 43.290 ;
        RECT 59.280 43.080 59.520 43.120 ;
        RECT 62.060 43.110 62.230 43.120 ;
        RECT 58.400 42.770 58.570 42.810 ;
        RECT 38.510 42.570 38.680 42.620 ;
        RECT 58.340 42.600 58.570 42.770 ;
        RECT 38.480 42.350 38.700 42.570 ;
        RECT 38.510 42.290 38.680 42.350 ;
        RECT 39.030 42.210 39.360 42.390 ;
        RECT 42.170 42.380 42.340 42.430 ;
        RECT 39.610 42.210 41.770 42.380 ;
        RECT 42.010 42.210 42.340 42.380 ;
        RECT 42.630 42.240 42.840 42.570 ;
        RECT 39.060 41.770 39.330 42.210 ;
        RECT 40.540 41.950 40.870 42.210 ;
        RECT 42.080 42.070 42.340 42.210 ;
        RECT 43.080 42.070 43.260 42.510 ;
        RECT 43.810 42.300 45.170 42.410 ;
        RECT 43.810 42.240 45.250 42.300 ;
        RECT 44.610 42.230 45.250 42.240 ;
        RECT 39.100 41.760 39.330 41.770 ;
        RECT 42.080 41.900 43.260 42.070 ;
        RECT 44.780 42.130 45.250 42.230 ;
        RECT 45.720 42.150 46.680 42.320 ;
        RECT 58.400 42.250 58.570 42.600 ;
        RECT 58.740 42.670 58.930 42.690 ;
        RECT 61.740 42.670 62.070 42.850 ;
        RECT 58.740 42.500 59.300 42.670 ;
        RECT 59.760 42.500 62.510 42.670 ;
        RECT 58.740 42.460 58.930 42.500 ;
        RECT 63.040 42.430 63.210 43.360 ;
        RECT 63.440 42.560 63.610 43.410 ;
        RECT 65.890 43.290 66.110 43.880 ;
        RECT 66.630 43.320 66.830 43.890 ;
        RECT 67.640 43.600 67.960 43.640 ;
        RECT 67.630 43.560 67.960 43.600 ;
        RECT 67.380 43.390 67.960 43.560 ;
        RECT 67.640 43.380 67.960 43.390 ;
        RECT 88.440 43.600 88.760 43.640 ;
        RECT 88.440 43.560 88.770 43.600 ;
        RECT 88.440 43.390 89.020 43.560 ;
        RECT 88.440 43.380 88.760 43.390 ;
        RECT 89.570 43.320 89.770 43.890 ;
        RECT 90.300 43.880 90.510 43.910 ;
        RECT 111.510 43.890 112.090 44.060 ;
        RECT 90.290 43.290 90.510 43.880 ;
        RECT 65.890 42.270 66.110 42.860 ;
        RECT 65.890 42.240 66.100 42.270 ;
        RECT 66.630 42.260 66.830 42.830 ;
        RECT 67.640 42.760 67.960 42.770 ;
        RECT 67.380 42.590 67.960 42.760 ;
        RECT 67.630 42.550 67.960 42.590 ;
        RECT 67.640 42.510 67.960 42.550 ;
        RECT 88.440 42.760 88.760 42.770 ;
        RECT 88.440 42.590 89.020 42.760 ;
        RECT 88.440 42.550 88.770 42.590 ;
        RECT 88.440 42.510 88.760 42.550 ;
        RECT 89.570 42.260 89.770 42.830 ;
        RECT 90.290 42.270 90.510 42.860 ;
        RECT 42.080 41.760 42.340 41.900 ;
        RECT 44.780 41.880 45.030 42.130 ;
        RECT 39.100 41.590 39.860 41.760 ;
        RECT 40.110 41.590 41.280 41.760 ;
        RECT 41.520 41.730 42.340 41.760 ;
        RECT 43.580 41.730 43.760 41.790 ;
        RECT 41.520 41.590 42.630 41.730 ;
        RECT 40.510 41.490 40.860 41.590 ;
        RECT 42.170 41.560 42.630 41.590 ;
        RECT 43.080 41.560 43.760 41.730 ;
        RECT 44.700 41.710 45.030 41.880 ;
        RECT 46.500 41.690 46.680 42.150 ;
        RECT 43.120 41.540 43.760 41.560 ;
        RECT 43.580 41.530 43.760 41.540 ;
        RECT 45.360 41.530 45.960 41.680 ;
        RECT 43.580 41.510 45.960 41.530 ;
        RECT 46.420 41.520 46.750 41.690 ;
        RECT 58.400 41.660 58.570 42.010 ;
        RECT 65.900 41.890 66.100 42.240 ;
        RECT 90.300 42.240 90.510 42.270 ;
        RECT 67.640 42.190 67.960 42.220 ;
        RECT 67.630 42.140 67.960 42.190 ;
        RECT 67.380 41.970 67.960 42.140 ;
        RECT 67.640 41.960 67.960 41.970 ;
        RECT 88.440 42.190 88.760 42.220 ;
        RECT 88.440 42.140 88.770 42.190 ;
        RECT 88.440 41.970 89.020 42.140 ;
        RECT 88.440 41.960 88.760 41.970 ;
        RECT 90.300 41.890 90.500 42.240 ;
        RECT 43.580 41.360 45.810 41.510 ;
        RECT 58.340 41.490 58.570 41.660 ;
        RECT 58.740 41.760 58.930 41.800 ;
        RECT 58.740 41.590 59.300 41.760 ;
        RECT 59.760 41.590 62.510 41.760 ;
        RECT 58.740 41.570 58.930 41.590 ;
        RECT 58.400 41.450 58.570 41.490 ;
        RECT 61.740 41.410 62.070 41.590 ;
        RECT 38.510 41.020 38.680 41.070 ;
        RECT 38.480 40.800 38.700 41.020 ;
        RECT 38.510 40.740 38.680 40.800 ;
        RECT 39.030 40.660 39.360 40.840 ;
        RECT 42.170 40.830 42.340 40.880 ;
        RECT 39.610 40.660 41.770 40.830 ;
        RECT 42.010 40.660 42.340 40.830 ;
        RECT 42.630 40.690 42.840 41.020 ;
        RECT 39.060 40.220 39.330 40.660 ;
        RECT 40.540 40.400 40.870 40.660 ;
        RECT 42.080 40.520 42.340 40.660 ;
        RECT 43.080 40.520 43.260 40.960 ;
        RECT 43.810 40.750 45.170 40.860 ;
        RECT 58.470 40.850 58.640 41.270 ;
        RECT 59.280 41.140 59.520 41.180 ;
        RECT 62.060 41.140 62.230 41.150 ;
        RECT 58.950 40.970 59.520 41.140 ;
        RECT 59.760 40.970 61.100 41.140 ;
        RECT 61.550 40.970 62.510 41.140 ;
        RECT 59.280 40.940 59.520 40.970 ;
        RECT 63.040 40.900 63.210 41.830 ;
        RECT 63.440 40.850 63.610 41.700 ;
        RECT 43.810 40.690 45.250 40.750 ;
        RECT 44.610 40.680 45.250 40.690 ;
        RECT 39.100 40.210 39.330 40.220 ;
        RECT 42.080 40.350 43.260 40.520 ;
        RECT 44.780 40.580 45.250 40.680 ;
        RECT 45.720 40.600 46.680 40.770 ;
        RECT 42.080 40.210 42.340 40.350 ;
        RECT 44.780 40.330 45.030 40.580 ;
        RECT 39.100 40.040 39.860 40.210 ;
        RECT 40.110 40.040 41.280 40.210 ;
        RECT 41.520 40.180 42.340 40.210 ;
        RECT 43.580 40.180 43.760 40.240 ;
        RECT 41.520 40.040 42.630 40.180 ;
        RECT 40.510 39.940 40.860 40.040 ;
        RECT 42.170 40.010 42.630 40.040 ;
        RECT 43.080 40.010 43.760 40.180 ;
        RECT 44.700 40.160 45.030 40.330 ;
        RECT 46.500 40.140 46.680 40.600 ;
        RECT 43.120 39.990 43.760 40.010 ;
        RECT 43.580 39.980 43.760 39.990 ;
        RECT 45.360 39.980 45.960 40.130 ;
        RECT 43.580 39.960 45.960 39.980 ;
        RECT 46.420 39.970 46.750 40.140 ;
        RECT 58.470 40.060 58.640 40.480 ;
        RECT 59.280 40.360 59.520 40.390 ;
        RECT 58.950 40.190 59.520 40.360 ;
        RECT 59.760 40.190 61.100 40.360 ;
        RECT 61.550 40.190 62.510 40.360 ;
        RECT 59.280 40.150 59.520 40.190 ;
        RECT 62.060 40.180 62.230 40.190 ;
        RECT 43.580 39.810 45.810 39.960 ;
        RECT 58.400 39.840 58.570 39.880 ;
        RECT 58.340 39.670 58.570 39.840 ;
        RECT 38.510 39.470 38.680 39.520 ;
        RECT 38.480 39.250 38.700 39.470 ;
        RECT 38.510 39.190 38.680 39.250 ;
        RECT 39.030 39.110 39.360 39.290 ;
        RECT 42.170 39.280 42.340 39.330 ;
        RECT 39.610 39.110 41.770 39.280 ;
        RECT 42.010 39.110 42.340 39.280 ;
        RECT 42.630 39.140 42.840 39.470 ;
        RECT 39.060 38.670 39.330 39.110 ;
        RECT 40.540 38.850 40.870 39.110 ;
        RECT 42.080 38.970 42.340 39.110 ;
        RECT 43.080 38.970 43.260 39.410 ;
        RECT 58.400 39.320 58.570 39.670 ;
        RECT 58.740 39.740 58.930 39.760 ;
        RECT 61.740 39.740 62.070 39.920 ;
        RECT 58.740 39.570 59.300 39.740 ;
        RECT 59.760 39.570 62.510 39.740 ;
        RECT 58.740 39.530 58.930 39.570 ;
        RECT 63.040 39.500 63.210 40.430 ;
        RECT 63.440 39.630 63.610 40.480 ;
        RECT 43.810 39.200 45.170 39.310 ;
        RECT 43.810 39.140 45.250 39.200 ;
        RECT 44.610 39.130 45.250 39.140 ;
        RECT 39.100 38.660 39.330 38.670 ;
        RECT 42.080 38.800 43.260 38.970 ;
        RECT 44.780 39.030 45.250 39.130 ;
        RECT 45.720 39.050 46.680 39.220 ;
        RECT 42.080 38.660 42.340 38.800 ;
        RECT 44.780 38.780 45.030 39.030 ;
        RECT 39.100 38.490 39.860 38.660 ;
        RECT 40.110 38.490 41.280 38.660 ;
        RECT 41.520 38.630 42.340 38.660 ;
        RECT 43.580 38.630 43.760 38.690 ;
        RECT 41.520 38.490 42.630 38.630 ;
        RECT 40.510 38.390 40.860 38.490 ;
        RECT 42.170 38.460 42.630 38.490 ;
        RECT 43.080 38.460 43.760 38.630 ;
        RECT 44.700 38.610 45.030 38.780 ;
        RECT 46.500 38.590 46.680 39.050 ;
        RECT 58.400 38.730 58.570 39.080 ;
        RECT 43.120 38.440 43.760 38.460 ;
        RECT 43.580 38.430 43.760 38.440 ;
        RECT 45.360 38.430 45.960 38.580 ;
        RECT 43.580 38.410 45.960 38.430 ;
        RECT 46.420 38.420 46.750 38.590 ;
        RECT 58.340 38.560 58.570 38.730 ;
        RECT 58.740 38.830 58.930 38.870 ;
        RECT 58.740 38.660 59.300 38.830 ;
        RECT 59.760 38.660 62.510 38.830 ;
        RECT 58.740 38.640 58.930 38.660 ;
        RECT 58.400 38.520 58.570 38.560 ;
        RECT 61.740 38.480 62.070 38.660 ;
        RECT 43.580 38.260 45.810 38.410 ;
        RECT 38.510 37.920 38.680 37.970 ;
        RECT 58.470 37.920 58.640 38.340 ;
        RECT 59.280 38.210 59.520 38.250 ;
        RECT 62.060 38.210 62.230 38.220 ;
        RECT 58.950 38.040 59.520 38.210 ;
        RECT 59.760 38.040 61.100 38.210 ;
        RECT 61.550 38.040 62.510 38.210 ;
        RECT 59.280 38.010 59.520 38.040 ;
        RECT 63.040 37.970 63.210 38.900 ;
        RECT 63.440 37.920 63.610 38.770 ;
        RECT 38.480 37.700 38.700 37.920 ;
        RECT 38.510 37.640 38.680 37.700 ;
        RECT 39.030 37.560 39.360 37.740 ;
        RECT 42.170 37.730 42.340 37.780 ;
        RECT 39.610 37.560 41.770 37.730 ;
        RECT 42.010 37.560 42.340 37.730 ;
        RECT 42.630 37.590 42.840 37.920 ;
        RECT 39.060 37.120 39.330 37.560 ;
        RECT 40.540 37.300 40.870 37.560 ;
        RECT 42.080 37.420 42.340 37.560 ;
        RECT 43.080 37.420 43.260 37.860 ;
        RECT 43.810 37.650 45.170 37.760 ;
        RECT 43.810 37.590 45.250 37.650 ;
        RECT 44.610 37.580 45.250 37.590 ;
        RECT 39.100 37.110 39.330 37.120 ;
        RECT 42.080 37.250 43.260 37.420 ;
        RECT 44.780 37.480 45.250 37.580 ;
        RECT 45.720 37.500 46.680 37.670 ;
        RECT 66.480 37.530 66.680 37.880 ;
        RECT 68.220 37.800 68.540 37.810 ;
        RECT 67.960 37.630 68.540 37.800 ;
        RECT 68.210 37.580 68.540 37.630 ;
        RECT 68.220 37.550 68.540 37.580 ;
        RECT 42.080 37.110 42.340 37.250 ;
        RECT 44.780 37.230 45.030 37.480 ;
        RECT 39.100 36.940 39.860 37.110 ;
        RECT 40.110 36.940 41.280 37.110 ;
        RECT 41.520 37.080 42.340 37.110 ;
        RECT 43.580 37.080 43.760 37.140 ;
        RECT 41.520 36.940 42.630 37.080 ;
        RECT 40.510 36.840 40.860 36.940 ;
        RECT 42.170 36.910 42.630 36.940 ;
        RECT 43.080 36.910 43.760 37.080 ;
        RECT 44.700 37.060 45.030 37.230 ;
        RECT 46.500 37.040 46.680 37.500 ;
        RECT 66.470 37.500 66.680 37.530 ;
        RECT 43.120 36.890 43.760 36.910 ;
        RECT 43.580 36.880 43.760 36.890 ;
        RECT 45.360 36.880 45.960 37.030 ;
        RECT 43.580 36.860 45.960 36.880 ;
        RECT 46.420 36.870 46.750 37.040 ;
        RECT 66.470 36.910 66.690 37.500 ;
        RECT 67.210 36.940 67.410 37.510 ;
        RECT 68.220 37.220 68.540 37.260 ;
        RECT 68.210 37.180 68.540 37.220 ;
        RECT 67.960 37.010 68.540 37.180 ;
        RECT 68.220 37.000 68.540 37.010 ;
        RECT 43.580 36.710 45.810 36.860 ;
        RECT 66.470 35.880 66.690 36.470 ;
        RECT 66.470 35.850 66.680 35.880 ;
        RECT 67.210 35.870 67.410 36.440 ;
        RECT 69.350 36.430 69.520 36.940 ;
        RECT 73.370 36.460 73.540 36.970 ;
        RECT 68.220 36.370 68.540 36.380 ;
        RECT 67.960 36.200 68.540 36.370 ;
        RECT 68.210 36.160 68.540 36.200 ;
        RECT 68.220 36.120 68.540 36.160 ;
        RECT 66.480 35.500 66.680 35.850 ;
        RECT 68.220 35.800 68.540 35.830 ;
        RECT 68.210 35.750 68.540 35.800 ;
        RECT 67.960 35.580 68.540 35.750 ;
        RECT 68.220 35.570 68.540 35.580 ;
        RECT 66.850 35.100 67.290 35.270 ;
        RECT 15.580 34.180 15.750 34.670 ;
        RECT 15.430 34.150 15.750 34.180 ;
        RECT 16.130 34.180 16.300 34.670 ;
        RECT 16.770 34.620 16.940 34.670 ;
        RECT 17.320 34.620 17.490 34.670 ;
        RECT 16.650 34.590 16.970 34.620 ;
        RECT 17.300 34.590 17.620 34.620 ;
        RECT 16.650 34.400 16.980 34.590 ;
        RECT 17.300 34.400 17.630 34.590 ;
        RECT 66.480 34.520 66.680 34.870 ;
        RECT 68.220 34.790 68.540 34.800 ;
        RECT 67.960 34.620 68.540 34.790 ;
        RECT 68.210 34.570 68.540 34.620 ;
        RECT 69.340 34.570 69.510 35.760 ;
        RECT 71.150 34.890 71.700 35.320 ;
        RECT 68.220 34.540 68.540 34.570 ;
        RECT 66.470 34.490 66.680 34.520 ;
        RECT 73.360 34.510 73.530 35.700 ;
        RECT 75.180 34.960 75.730 35.390 ;
        RECT 16.650 34.360 16.970 34.400 ;
        RECT 17.300 34.360 17.620 34.400 ;
        RECT 16.130 34.150 16.450 34.180 ;
        RECT 15.430 33.960 15.760 34.150 ;
        RECT 16.130 33.960 16.460 34.150 ;
        RECT 15.430 33.920 15.750 33.960 ;
        RECT 15.040 32.460 15.210 32.480 ;
        RECT 15.020 32.030 15.230 32.460 ;
        RECT 15.580 32.270 15.750 33.920 ;
        RECT 16.130 33.920 16.450 33.960 ;
        RECT 16.130 32.270 16.300 33.920 ;
        RECT 16.770 32.270 16.940 34.360 ;
        RECT 17.320 32.270 17.490 34.360 ;
        RECT 66.470 33.900 66.690 34.490 ;
        RECT 67.210 33.930 67.410 34.500 ;
        RECT 68.220 34.210 68.540 34.250 ;
        RECT 68.210 34.170 68.540 34.210 ;
        RECT 67.960 34.000 68.540 34.170 ;
        RECT 68.220 33.990 68.540 34.000 ;
        RECT 79.590 33.870 79.910 33.900 ;
        RECT 17.870 32.910 18.040 33.760 ;
        RECT 79.590 33.700 81.380 33.870 ;
        RECT 79.590 33.680 79.920 33.700 ;
        RECT 58.470 33.230 58.640 33.650 ;
        RECT 59.280 33.530 59.520 33.560 ;
        RECT 58.950 33.360 59.520 33.530 ;
        RECT 59.760 33.360 61.100 33.530 ;
        RECT 61.550 33.360 62.510 33.530 ;
        RECT 59.280 33.320 59.520 33.360 ;
        RECT 62.060 33.350 62.230 33.360 ;
        RECT 58.400 33.010 58.570 33.050 ;
        RECT 38.510 32.800 38.680 32.850 ;
        RECT 58.340 32.840 58.570 33.010 ;
        RECT 38.480 32.580 38.700 32.800 ;
        RECT 38.510 32.520 38.680 32.580 ;
        RECT 39.030 32.440 39.360 32.620 ;
        RECT 42.170 32.610 42.340 32.660 ;
        RECT 39.610 32.440 41.770 32.610 ;
        RECT 42.010 32.440 42.340 32.610 ;
        RECT 42.630 32.470 42.840 32.800 ;
        RECT 17.760 32.280 18.190 32.300 ;
        RECT 17.760 32.110 18.210 32.280 ;
        RECT 17.760 32.090 18.190 32.110 ;
        RECT 39.060 32.000 39.330 32.440 ;
        RECT 40.540 32.180 40.870 32.440 ;
        RECT 42.080 32.300 42.340 32.440 ;
        RECT 43.080 32.300 43.260 32.740 ;
        RECT 43.810 32.530 45.170 32.640 ;
        RECT 43.810 32.470 45.250 32.530 ;
        RECT 44.610 32.460 45.250 32.470 ;
        RECT 39.100 31.990 39.330 32.000 ;
        RECT 42.080 32.130 43.260 32.300 ;
        RECT 44.780 32.360 45.250 32.460 ;
        RECT 45.720 32.380 46.680 32.550 ;
        RECT 58.400 32.490 58.570 32.840 ;
        RECT 58.740 32.910 58.930 32.930 ;
        RECT 61.740 32.910 62.070 33.090 ;
        RECT 58.740 32.740 59.300 32.910 ;
        RECT 59.760 32.740 62.510 32.910 ;
        RECT 58.740 32.700 58.930 32.740 ;
        RECT 63.040 32.670 63.210 33.600 ;
        RECT 63.440 32.800 63.610 33.650 ;
        RECT 79.590 33.640 79.910 33.680 ;
        RECT 81.210 33.470 81.380 33.700 ;
        RECT 66.470 32.880 66.690 33.470 ;
        RECT 66.470 32.850 66.680 32.880 ;
        RECT 67.210 32.870 67.410 33.440 ;
        RECT 68.220 33.370 68.540 33.380 ;
        RECT 67.960 33.200 68.540 33.370 ;
        RECT 80.060 33.220 80.400 33.470 ;
        RECT 80.570 33.300 80.900 33.470 ;
        RECT 81.120 33.300 81.460 33.470 ;
        RECT 68.210 33.160 68.540 33.200 ;
        RECT 68.220 33.120 68.540 33.160 ;
        RECT 79.740 32.960 80.400 33.220 ;
        RECT 80.650 33.130 80.820 33.300 ;
        RECT 81.210 33.130 81.380 33.300 ;
        RECT 80.570 32.960 80.900 33.130 ;
        RECT 81.120 32.960 81.460 33.130 ;
        RECT 66.480 32.500 66.680 32.850 ;
        RECT 68.220 32.800 68.540 32.830 ;
        RECT 68.210 32.750 68.540 32.800 ;
        RECT 67.960 32.580 68.540 32.750 ;
        RECT 68.220 32.570 68.540 32.580 ;
        RECT 80.650 32.730 80.900 32.960 ;
        RECT 81.780 32.880 82.290 33.550 ;
        RECT 80.650 32.560 81.320 32.730 ;
        RECT 42.080 31.990 42.340 32.130 ;
        RECT 44.780 32.110 45.030 32.360 ;
        RECT 39.100 31.820 39.860 31.990 ;
        RECT 40.110 31.820 41.280 31.990 ;
        RECT 41.520 31.960 42.340 31.990 ;
        RECT 43.580 31.960 43.760 32.020 ;
        RECT 41.520 31.820 42.630 31.960 ;
        RECT 14.120 28.910 14.290 31.400 ;
        RECT 14.670 28.910 14.840 31.410 ;
        RECT 15.030 31.390 15.240 31.820 ;
        RECT 17.770 31.740 18.200 31.760 ;
        RECT 17.770 31.570 18.220 31.740 ;
        RECT 40.510 31.720 40.860 31.820 ;
        RECT 42.170 31.790 42.630 31.820 ;
        RECT 43.080 31.790 43.760 31.960 ;
        RECT 44.700 31.940 45.030 32.110 ;
        RECT 46.500 31.920 46.680 32.380 ;
        RECT 80.650 32.330 80.900 32.560 ;
        RECT 43.120 31.770 43.760 31.790 ;
        RECT 43.580 31.760 43.760 31.770 ;
        RECT 45.360 31.760 45.960 31.910 ;
        RECT 43.580 31.740 45.960 31.760 ;
        RECT 46.420 31.750 46.750 31.920 ;
        RECT 58.400 31.900 58.570 32.250 ;
        RECT 79.740 32.070 80.400 32.330 ;
        RECT 80.570 32.160 80.900 32.330 ;
        RECT 81.120 32.160 81.460 32.330 ;
        RECT 43.580 31.590 45.810 31.740 ;
        RECT 58.340 31.730 58.570 31.900 ;
        RECT 58.740 32.000 58.930 32.040 ;
        RECT 58.740 31.830 59.300 32.000 ;
        RECT 59.760 31.830 62.510 32.000 ;
        RECT 58.740 31.810 58.930 31.830 ;
        RECT 58.400 31.690 58.570 31.730 ;
        RECT 61.740 31.650 62.070 31.830 ;
        RECT 17.770 31.550 18.200 31.570 ;
        RECT 15.050 31.370 15.220 31.390 ;
        RECT 15.300 30.300 15.470 31.400 ;
        RECT 15.300 30.270 15.780 30.300 ;
        RECT 15.300 30.080 15.790 30.270 ;
        RECT 15.300 30.040 15.780 30.080 ;
        RECT 15.300 28.910 15.470 30.040 ;
        RECT 15.850 28.910 16.020 31.410 ;
        RECT 38.510 31.250 38.680 31.300 ;
        RECT 38.480 31.030 38.700 31.250 ;
        RECT 17.860 30.360 18.030 31.030 ;
        RECT 38.510 30.970 38.680 31.030 ;
        RECT 39.030 30.890 39.360 31.070 ;
        RECT 42.170 31.060 42.340 31.110 ;
        RECT 39.610 30.890 41.770 31.060 ;
        RECT 42.010 30.890 42.340 31.060 ;
        RECT 42.630 30.920 42.840 31.250 ;
        RECT 39.060 30.450 39.330 30.890 ;
        RECT 40.540 30.630 40.870 30.890 ;
        RECT 42.080 30.750 42.340 30.890 ;
        RECT 43.080 30.750 43.260 31.190 ;
        RECT 58.470 31.090 58.640 31.510 ;
        RECT 59.280 31.380 59.520 31.420 ;
        RECT 62.060 31.380 62.230 31.390 ;
        RECT 58.950 31.210 59.520 31.380 ;
        RECT 59.760 31.210 61.100 31.380 ;
        RECT 61.550 31.210 62.510 31.380 ;
        RECT 59.280 31.180 59.520 31.210 ;
        RECT 63.040 31.140 63.210 32.070 ;
        RECT 63.440 31.090 63.610 31.940 ;
        RECT 80.060 31.820 80.400 32.070 ;
        RECT 80.650 31.990 80.820 32.160 ;
        RECT 81.210 31.990 81.380 32.160 ;
        RECT 80.570 31.820 80.900 31.990 ;
        RECT 81.120 31.820 81.460 31.990 ;
        RECT 79.590 31.610 79.910 31.650 ;
        RECT 79.590 31.590 79.920 31.610 ;
        RECT 81.210 31.590 81.380 31.820 ;
        RECT 81.780 31.740 82.290 32.410 ;
        RECT 79.590 31.420 81.380 31.590 ;
        RECT 79.590 31.390 79.910 31.420 ;
        RECT 79.590 31.100 79.910 31.130 ;
        RECT 43.810 30.980 45.170 31.090 ;
        RECT 43.810 30.920 45.250 30.980 ;
        RECT 44.610 30.910 45.250 30.920 ;
        RECT 39.100 30.440 39.330 30.450 ;
        RECT 42.080 30.580 43.260 30.750 ;
        RECT 44.780 30.810 45.250 30.910 ;
        RECT 45.720 30.830 46.680 31.000 ;
        RECT 79.590 30.930 81.380 31.100 ;
        RECT 79.590 30.910 79.920 30.930 ;
        RECT 79.590 30.870 79.910 30.910 ;
        RECT 42.080 30.440 42.340 30.580 ;
        RECT 44.780 30.560 45.030 30.810 ;
        RECT 16.150 30.260 16.470 30.290 ;
        RECT 39.100 30.270 39.860 30.440 ;
        RECT 40.110 30.270 41.280 30.440 ;
        RECT 41.520 30.410 42.340 30.440 ;
        RECT 43.580 30.410 43.760 30.470 ;
        RECT 41.520 30.270 42.630 30.410 ;
        RECT 16.150 30.070 16.480 30.260 ;
        RECT 40.510 30.170 40.860 30.270 ;
        RECT 42.170 30.240 42.630 30.270 ;
        RECT 43.080 30.240 43.760 30.410 ;
        RECT 44.700 30.390 45.030 30.560 ;
        RECT 46.500 30.370 46.680 30.830 ;
        RECT 43.120 30.220 43.760 30.240 ;
        RECT 43.580 30.210 43.760 30.220 ;
        RECT 45.360 30.210 45.960 30.360 ;
        RECT 43.580 30.190 45.960 30.210 ;
        RECT 46.420 30.200 46.750 30.370 ;
        RECT 58.470 30.300 58.640 30.720 ;
        RECT 59.280 30.600 59.520 30.630 ;
        RECT 58.950 30.430 59.520 30.600 ;
        RECT 59.760 30.430 61.100 30.600 ;
        RECT 61.550 30.430 62.510 30.600 ;
        RECT 59.280 30.390 59.520 30.430 ;
        RECT 62.060 30.420 62.230 30.430 ;
        RECT 16.150 30.030 16.470 30.070 ;
        RECT 43.580 30.040 45.810 30.190 ;
        RECT 58.400 30.080 58.570 30.120 ;
        RECT 58.340 29.910 58.570 30.080 ;
        RECT 38.510 29.700 38.680 29.750 ;
        RECT 16.630 29.490 16.950 29.520 ;
        RECT 16.630 29.300 16.960 29.490 ;
        RECT 38.480 29.480 38.700 29.700 ;
        RECT 17.340 29.430 17.660 29.460 ;
        RECT 16.630 29.260 16.950 29.300 ;
        RECT 17.340 29.240 17.670 29.430 ;
        RECT 38.510 29.420 38.680 29.480 ;
        RECT 39.030 29.340 39.360 29.520 ;
        RECT 42.170 29.510 42.340 29.560 ;
        RECT 39.610 29.340 41.770 29.510 ;
        RECT 42.010 29.340 42.340 29.510 ;
        RECT 42.630 29.370 42.840 29.700 ;
        RECT 17.340 29.200 17.660 29.240 ;
        RECT 39.060 28.900 39.330 29.340 ;
        RECT 40.540 29.080 40.870 29.340 ;
        RECT 42.080 29.200 42.340 29.340 ;
        RECT 43.080 29.200 43.260 29.640 ;
        RECT 58.400 29.560 58.570 29.910 ;
        RECT 58.740 29.980 58.930 30.000 ;
        RECT 61.740 29.980 62.070 30.160 ;
        RECT 58.740 29.810 59.300 29.980 ;
        RECT 59.760 29.810 62.510 29.980 ;
        RECT 58.740 29.770 58.930 29.810 ;
        RECT 63.040 29.740 63.210 30.670 ;
        RECT 63.440 29.870 63.610 30.720 ;
        RECT 81.210 30.700 81.380 30.930 ;
        RECT 80.060 30.450 80.400 30.700 ;
        RECT 80.570 30.530 80.900 30.700 ;
        RECT 81.120 30.530 81.460 30.700 ;
        RECT 79.740 30.190 80.400 30.450 ;
        RECT 80.650 30.360 80.820 30.530 ;
        RECT 81.210 30.360 81.380 30.530 ;
        RECT 80.570 30.190 80.900 30.360 ;
        RECT 81.120 30.190 81.460 30.360 ;
        RECT 80.650 29.960 80.900 30.190 ;
        RECT 81.780 30.110 82.290 30.780 ;
        RECT 80.650 29.790 81.320 29.960 ;
        RECT 80.650 29.560 80.900 29.790 ;
        RECT 43.810 29.430 45.170 29.540 ;
        RECT 68.150 29.460 68.470 29.500 ;
        RECT 43.810 29.370 45.250 29.430 ;
        RECT 44.610 29.360 45.250 29.370 ;
        RECT 39.100 28.890 39.330 28.900 ;
        RECT 42.080 29.030 43.260 29.200 ;
        RECT 44.780 29.260 45.250 29.360 ;
        RECT 45.720 29.280 46.680 29.450 ;
        RECT 42.080 28.890 42.340 29.030 ;
        RECT 44.780 29.010 45.030 29.260 ;
        RECT 39.100 28.720 39.860 28.890 ;
        RECT 40.110 28.720 41.280 28.890 ;
        RECT 41.520 28.860 42.340 28.890 ;
        RECT 43.580 28.860 43.760 28.920 ;
        RECT 41.520 28.720 42.630 28.860 ;
        RECT 14.030 28.200 14.200 28.270 ;
        RECT 13.960 28.170 14.280 28.200 ;
        RECT 13.950 27.980 14.280 28.170 ;
        RECT 13.960 27.940 14.280 27.980 ;
        RECT 14.030 25.430 14.200 27.940 ;
        RECT 14.580 27.530 14.750 28.270 ;
        RECT 15.130 28.210 15.300 28.270 ;
        RECT 15.060 28.180 15.380 28.210 ;
        RECT 15.050 27.990 15.380 28.180 ;
        RECT 15.060 27.950 15.380 27.990 ;
        RECT 14.510 27.500 14.830 27.530 ;
        RECT 14.500 27.310 14.830 27.500 ;
        RECT 14.510 27.270 14.830 27.310 ;
        RECT 14.580 26.160 14.750 27.270 ;
        RECT 14.510 26.130 14.830 26.160 ;
        RECT 14.500 25.940 14.830 26.130 ;
        RECT 14.510 25.900 14.830 25.940 ;
        RECT 13.960 25.400 14.280 25.430 ;
        RECT 13.950 25.210 14.280 25.400 ;
        RECT 13.960 25.170 14.280 25.210 ;
        RECT 14.030 24.090 14.200 25.170 ;
        RECT 13.950 24.060 14.270 24.090 ;
        RECT 13.940 23.870 14.270 24.060 ;
        RECT 13.950 23.830 14.270 23.870 ;
        RECT 14.030 23.090 14.200 23.830 ;
        RECT 14.580 23.390 14.750 25.900 ;
        RECT 15.130 25.430 15.300 27.950 ;
        RECT 15.680 27.530 15.850 28.270 ;
        RECT 16.230 28.210 16.400 28.270 ;
        RECT 16.150 28.180 16.470 28.210 ;
        RECT 16.140 27.990 16.470 28.180 ;
        RECT 16.150 27.950 16.470 27.990 ;
        RECT 15.610 27.500 15.930 27.530 ;
        RECT 15.600 27.310 15.930 27.500 ;
        RECT 15.610 27.270 15.930 27.310 ;
        RECT 15.680 26.160 15.850 27.270 ;
        RECT 15.610 26.130 15.930 26.160 ;
        RECT 15.600 25.940 15.930 26.130 ;
        RECT 15.610 25.900 15.930 25.940 ;
        RECT 15.060 25.400 15.380 25.430 ;
        RECT 15.050 25.210 15.380 25.400 ;
        RECT 15.060 25.170 15.380 25.210 ;
        RECT 15.130 24.080 15.300 25.170 ;
        RECT 15.060 24.050 15.380 24.080 ;
        RECT 15.050 23.860 15.380 24.050 ;
        RECT 15.060 23.820 15.380 23.860 ;
        RECT 14.510 23.360 14.830 23.390 ;
        RECT 14.500 23.170 14.830 23.360 ;
        RECT 14.510 23.130 14.830 23.170 ;
        RECT 14.580 23.090 14.750 23.130 ;
        RECT 15.130 23.090 15.300 23.820 ;
        RECT 15.680 23.380 15.850 25.900 ;
        RECT 16.230 25.430 16.400 27.950 ;
        RECT 16.780 27.530 16.950 28.270 ;
        RECT 17.190 27.990 17.700 28.670 ;
        RECT 40.510 28.620 40.860 28.720 ;
        RECT 42.170 28.690 42.630 28.720 ;
        RECT 43.080 28.690 43.760 28.860 ;
        RECT 44.700 28.840 45.030 29.010 ;
        RECT 46.500 28.820 46.680 29.280 ;
        RECT 58.400 28.970 58.570 29.320 ;
        RECT 68.150 29.270 68.480 29.460 ;
        RECT 79.740 29.300 80.400 29.560 ;
        RECT 80.570 29.390 80.900 29.560 ;
        RECT 81.120 29.390 81.460 29.560 ;
        RECT 68.150 29.240 68.470 29.270 ;
        RECT 43.120 28.670 43.760 28.690 ;
        RECT 43.580 28.660 43.760 28.670 ;
        RECT 45.360 28.660 45.960 28.810 ;
        RECT 43.580 28.640 45.960 28.660 ;
        RECT 46.420 28.650 46.750 28.820 ;
        RECT 58.340 28.800 58.570 28.970 ;
        RECT 58.740 29.070 58.930 29.110 ;
        RECT 58.740 28.900 59.300 29.070 ;
        RECT 59.760 28.900 62.510 29.070 ;
        RECT 58.740 28.880 58.930 28.900 ;
        RECT 58.400 28.760 58.570 28.800 ;
        RECT 61.740 28.720 62.070 28.900 ;
        RECT 43.580 28.490 45.810 28.640 ;
        RECT 38.510 28.150 38.680 28.200 ;
        RECT 58.470 28.160 58.640 28.580 ;
        RECT 59.280 28.450 59.520 28.490 ;
        RECT 62.060 28.450 62.230 28.460 ;
        RECT 58.950 28.280 59.520 28.450 ;
        RECT 59.760 28.280 61.100 28.450 ;
        RECT 61.550 28.280 62.510 28.450 ;
        RECT 59.280 28.250 59.520 28.280 ;
        RECT 63.040 28.210 63.210 29.140 ;
        RECT 63.440 28.160 63.610 29.010 ;
        RECT 68.200 28.650 68.380 29.240 ;
        RECT 80.060 29.050 80.400 29.300 ;
        RECT 80.650 29.220 80.820 29.390 ;
        RECT 81.210 29.220 81.380 29.390 ;
        RECT 80.570 29.050 80.900 29.220 ;
        RECT 81.120 29.050 81.460 29.220 ;
        RECT 79.590 28.840 79.910 28.880 ;
        RECT 79.590 28.820 79.920 28.840 ;
        RECT 81.210 28.820 81.380 29.050 ;
        RECT 81.780 28.970 82.290 29.640 ;
        RECT 79.590 28.650 81.380 28.820 ;
        RECT 68.200 28.610 68.520 28.650 ;
        RECT 79.590 28.620 79.910 28.650 ;
        RECT 68.200 28.420 68.530 28.610 ;
        RECT 68.200 28.390 68.520 28.420 ;
        RECT 17.190 27.920 17.710 27.990 ;
        RECT 38.480 27.930 38.700 28.150 ;
        RECT 17.200 27.660 17.710 27.920 ;
        RECT 38.510 27.870 38.680 27.930 ;
        RECT 39.030 27.790 39.360 27.970 ;
        RECT 42.170 27.960 42.340 28.010 ;
        RECT 39.610 27.790 41.770 27.960 ;
        RECT 42.010 27.790 42.340 27.960 ;
        RECT 42.630 27.820 42.840 28.150 ;
        RECT 16.710 27.500 17.030 27.530 ;
        RECT 16.700 27.310 17.030 27.500 ;
        RECT 16.710 27.270 17.030 27.310 ;
        RECT 16.780 26.160 16.950 27.270 ;
        RECT 17.490 26.280 17.660 27.470 ;
        RECT 39.060 27.350 39.330 27.790 ;
        RECT 40.540 27.530 40.870 27.790 ;
        RECT 42.080 27.650 42.340 27.790 ;
        RECT 43.080 27.650 43.260 28.090 ;
        RECT 43.810 27.880 45.170 27.990 ;
        RECT 43.810 27.820 45.250 27.880 ;
        RECT 44.610 27.810 45.250 27.820 ;
        RECT 39.100 27.340 39.330 27.350 ;
        RECT 42.080 27.480 43.260 27.650 ;
        RECT 44.780 27.710 45.250 27.810 ;
        RECT 45.720 27.730 46.680 27.900 ;
        RECT 42.080 27.340 42.340 27.480 ;
        RECT 44.780 27.460 45.030 27.710 ;
        RECT 39.100 27.170 39.860 27.340 ;
        RECT 40.110 27.170 41.280 27.340 ;
        RECT 41.520 27.310 42.340 27.340 ;
        RECT 43.580 27.310 43.760 27.370 ;
        RECT 41.520 27.170 42.630 27.310 ;
        RECT 40.510 27.070 40.860 27.170 ;
        RECT 42.170 27.140 42.630 27.170 ;
        RECT 43.080 27.140 43.760 27.310 ;
        RECT 44.700 27.290 45.030 27.460 ;
        RECT 46.500 27.270 46.680 27.730 ;
        RECT 43.120 27.120 43.760 27.140 ;
        RECT 43.580 27.110 43.760 27.120 ;
        RECT 45.360 27.110 45.960 27.260 ;
        RECT 43.580 27.090 45.960 27.110 ;
        RECT 46.420 27.100 46.750 27.270 ;
        RECT 43.580 26.940 45.810 27.090 ;
        RECT 16.710 26.130 17.030 26.160 ;
        RECT 16.700 25.940 17.030 26.130 ;
        RECT 16.710 25.900 17.030 25.940 ;
        RECT 16.150 25.400 16.470 25.430 ;
        RECT 16.140 25.210 16.470 25.400 ;
        RECT 16.150 25.170 16.470 25.210 ;
        RECT 16.230 24.060 16.400 25.170 ;
        RECT 16.150 24.030 16.470 24.060 ;
        RECT 16.140 23.840 16.470 24.030 ;
        RECT 16.150 23.800 16.470 23.840 ;
        RECT 15.610 23.350 15.930 23.380 ;
        RECT 15.600 23.160 15.930 23.350 ;
        RECT 15.610 23.120 15.930 23.160 ;
        RECT 15.680 23.090 15.850 23.120 ;
        RECT 16.230 23.090 16.400 23.800 ;
        RECT 16.780 23.380 16.950 25.900 ;
        RECT 23.820 23.970 24.580 24.390 ;
        RECT 16.700 23.350 17.020 23.380 ;
        RECT 16.690 23.160 17.020 23.350 ;
        RECT 23.840 23.180 24.580 23.970 ;
        RECT 16.700 23.120 17.020 23.160 ;
        RECT 16.780 23.090 16.950 23.120 ;
        RECT 56.110 22.240 56.280 22.270 ;
        RECT 13.250 20.610 13.570 20.640 ;
        RECT 14.350 20.620 14.670 20.650 ;
        RECT 15.440 20.620 15.760 20.650 ;
        RECT 13.240 20.420 13.570 20.610 ;
        RECT 14.340 20.430 14.670 20.620 ;
        RECT 15.430 20.580 15.760 20.620 ;
        RECT 16.480 20.580 16.990 21.110 ;
        RECT 13.250 20.380 13.570 20.420 ;
        RECT 14.350 20.390 14.670 20.430 ;
        RECT 14.780 19.970 14.950 20.580 ;
        RECT 15.330 20.390 15.760 20.580 ;
        RECT 13.800 19.940 14.120 19.970 ;
        RECT 13.790 19.750 14.120 19.940 ;
        RECT 13.800 19.710 14.120 19.750 ;
        RECT 14.780 19.710 15.220 19.970 ;
        RECT 14.780 18.600 14.950 19.710 ;
        RECT 13.800 18.570 14.120 18.600 ;
        RECT 13.790 18.380 14.120 18.570 ;
        RECT 13.800 18.340 14.120 18.380 ;
        RECT 14.780 18.340 15.220 18.600 ;
        RECT 13.320 18.300 13.480 18.310 ;
        RECT 13.870 18.300 14.030 18.310 ;
        RECT 14.420 18.300 14.580 18.310 ;
        RECT 13.310 17.950 13.480 18.300 ;
        RECT 13.860 17.970 14.030 18.300 ;
        RECT 14.410 17.970 14.580 18.300 ;
        RECT 14.780 18.080 14.950 18.340 ;
        RECT 14.970 18.300 15.130 18.310 ;
        RECT 13.320 17.930 13.480 17.950 ;
        RECT 13.870 17.930 14.030 17.970 ;
        RECT 14.420 17.930 14.580 17.970 ;
        RECT 14.960 17.900 15.130 18.300 ;
        RECT 15.330 18.080 15.500 20.390 ;
        RECT 15.880 19.970 16.050 20.580 ;
        RECT 16.430 20.100 17.150 20.580 ;
        RECT 15.880 19.710 16.320 19.970 ;
        RECT 15.880 18.600 16.050 19.710 ;
        RECT 15.880 18.340 16.320 18.600 ;
        RECT 15.520 18.300 15.680 18.310 ;
        RECT 15.510 17.970 15.680 18.300 ;
        RECT 15.880 18.080 16.050 18.340 ;
        RECT 16.070 18.300 16.230 18.310 ;
        RECT 15.520 17.930 15.680 17.970 ;
        RECT 16.060 17.960 16.230 18.300 ;
        RECT 16.430 18.080 16.600 20.100 ;
        RECT 16.980 18.080 17.150 20.100 ;
        RECT 17.530 18.080 17.700 20.570 ;
        RECT 46.300 19.750 46.470 22.240 ;
        RECT 46.850 19.740 47.020 22.240 ;
        RECT 47.400 19.740 47.570 22.240 ;
        RECT 47.950 21.930 48.120 22.240 ;
        RECT 47.690 21.670 48.120 21.930 ;
        RECT 47.950 19.740 48.120 21.670 ;
        RECT 48.500 21.250 48.670 22.240 ;
        RECT 49.050 21.930 49.220 22.240 ;
        RECT 48.780 21.670 49.220 21.930 ;
        RECT 48.240 20.990 48.670 21.250 ;
        RECT 48.500 19.880 48.670 20.990 ;
        RECT 48.240 19.740 48.670 19.880 ;
        RECT 49.050 19.740 49.220 21.670 ;
        RECT 49.880 21.880 50.200 21.920 ;
        RECT 49.880 21.690 50.210 21.880 ;
        RECT 49.880 21.660 50.200 21.690 ;
        RECT 51.060 21.290 51.230 22.050 ;
        RECT 51.450 21.290 51.620 22.050 ;
        RECT 53.460 21.930 53.630 22.240 ;
        RECT 52.480 21.880 52.800 21.920 ;
        RECT 52.470 21.690 52.800 21.880 ;
        RECT 52.480 21.660 52.800 21.690 ;
        RECT 53.460 21.670 53.900 21.930 ;
        RECT 49.330 21.190 49.650 21.230 ;
        RECT 49.330 21.000 49.660 21.190 ;
        RECT 50.440 21.180 50.760 21.220 ;
        RECT 51.920 21.180 52.240 21.220 ;
        RECT 53.030 21.190 53.350 21.230 ;
        RECT 49.330 20.970 49.650 21.000 ;
        RECT 50.440 20.990 50.770 21.180 ;
        RECT 51.910 20.990 52.240 21.180 ;
        RECT 53.020 21.000 53.350 21.190 ;
        RECT 50.440 20.960 50.760 20.990 ;
        RECT 51.920 20.960 52.240 20.990 ;
        RECT 53.030 20.970 53.350 21.000 ;
        RECT 49.330 19.840 49.650 19.880 ;
        RECT 50.430 19.840 50.750 19.880 ;
        RECT 51.930 19.840 52.250 19.880 ;
        RECT 53.030 19.840 53.350 19.880 ;
        RECT 48.240 19.650 48.570 19.740 ;
        RECT 49.330 19.650 49.660 19.840 ;
        RECT 50.430 19.650 50.760 19.840 ;
        RECT 51.920 19.650 52.250 19.840 ;
        RECT 53.020 19.650 53.350 19.840 ;
        RECT 53.460 19.740 53.630 21.670 ;
        RECT 54.010 21.250 54.180 22.240 ;
        RECT 54.560 21.930 54.730 22.240 ;
        RECT 54.560 21.670 54.990 21.930 ;
        RECT 54.010 20.990 54.440 21.250 ;
        RECT 54.010 19.880 54.180 20.990 ;
        RECT 54.010 19.740 54.440 19.880 ;
        RECT 54.560 19.740 54.730 21.670 ;
        RECT 55.110 19.740 55.280 22.240 ;
        RECT 55.660 19.740 55.830 22.240 ;
        RECT 56.110 19.780 56.380 22.240 ;
        RECT 56.210 19.750 56.380 19.780 ;
        RECT 56.660 19.770 56.830 22.270 ;
        RECT 57.210 19.770 57.380 22.270 ;
        RECT 57.760 21.960 57.930 22.270 ;
        RECT 57.500 21.700 57.930 21.960 ;
        RECT 57.760 19.770 57.930 21.700 ;
        RECT 58.310 21.280 58.480 22.270 ;
        RECT 58.860 21.960 59.030 22.270 ;
        RECT 58.590 21.700 59.030 21.960 ;
        RECT 58.050 21.020 58.480 21.280 ;
        RECT 58.310 19.910 58.480 21.020 ;
        RECT 58.050 19.770 58.480 19.910 ;
        RECT 58.860 19.770 59.030 21.700 ;
        RECT 59.690 21.910 60.010 21.950 ;
        RECT 59.690 21.720 60.020 21.910 ;
        RECT 59.690 21.690 60.010 21.720 ;
        RECT 60.870 21.320 61.040 22.080 ;
        RECT 61.260 21.320 61.430 22.080 ;
        RECT 63.270 21.960 63.440 22.270 ;
        RECT 62.290 21.910 62.610 21.950 ;
        RECT 62.280 21.720 62.610 21.910 ;
        RECT 62.290 21.690 62.610 21.720 ;
        RECT 63.270 21.700 63.710 21.960 ;
        RECT 59.140 21.220 59.460 21.260 ;
        RECT 59.140 21.030 59.470 21.220 ;
        RECT 60.250 21.210 60.570 21.250 ;
        RECT 61.730 21.210 62.050 21.250 ;
        RECT 62.840 21.220 63.160 21.260 ;
        RECT 59.140 21.000 59.460 21.030 ;
        RECT 60.250 21.020 60.580 21.210 ;
        RECT 61.720 21.020 62.050 21.210 ;
        RECT 62.830 21.030 63.160 21.220 ;
        RECT 60.250 20.990 60.570 21.020 ;
        RECT 61.730 20.990 62.050 21.020 ;
        RECT 62.840 21.000 63.160 21.030 ;
        RECT 59.140 19.870 59.460 19.910 ;
        RECT 60.240 19.870 60.560 19.910 ;
        RECT 61.740 19.870 62.060 19.910 ;
        RECT 62.840 19.870 63.160 19.910 ;
        RECT 54.110 19.650 54.440 19.740 ;
        RECT 58.050 19.680 58.380 19.770 ;
        RECT 59.140 19.680 59.470 19.870 ;
        RECT 60.240 19.680 60.570 19.870 ;
        RECT 61.730 19.680 62.060 19.870 ;
        RECT 62.830 19.680 63.160 19.870 ;
        RECT 63.270 19.770 63.440 21.700 ;
        RECT 63.820 21.280 63.990 22.270 ;
        RECT 64.370 21.960 64.540 22.270 ;
        RECT 64.370 21.700 64.800 21.960 ;
        RECT 63.820 21.020 64.250 21.280 ;
        RECT 63.820 19.910 63.990 21.020 ;
        RECT 63.820 19.770 64.250 19.910 ;
        RECT 64.370 19.770 64.540 21.700 ;
        RECT 64.920 19.770 65.090 22.270 ;
        RECT 65.470 19.770 65.640 22.270 ;
        RECT 66.020 19.780 66.190 22.270 ;
        RECT 68.300 21.230 68.470 21.970 ;
        RECT 68.850 21.930 69.020 21.970 ;
        RECT 68.780 21.890 69.100 21.930 ;
        RECT 68.770 21.700 69.100 21.890 ;
        RECT 68.780 21.670 69.100 21.700 ;
        RECT 68.220 21.190 68.540 21.230 ;
        RECT 68.210 21.000 68.540 21.190 ;
        RECT 68.220 20.970 68.540 21.000 ;
        RECT 68.300 19.890 68.470 20.970 ;
        RECT 68.230 19.850 68.550 19.890 ;
        RECT 63.920 19.680 64.250 19.770 ;
        RECT 58.050 19.650 58.370 19.680 ;
        RECT 59.140 19.650 59.460 19.680 ;
        RECT 60.240 19.650 60.560 19.680 ;
        RECT 61.740 19.650 62.060 19.680 ;
        RECT 62.840 19.650 63.160 19.680 ;
        RECT 63.930 19.650 64.250 19.680 ;
        RECT 68.220 19.660 68.550 19.850 ;
        RECT 48.240 19.620 48.560 19.650 ;
        RECT 49.330 19.620 49.650 19.650 ;
        RECT 50.430 19.620 50.750 19.650 ;
        RECT 51.930 19.620 52.250 19.650 ;
        RECT 53.030 19.620 53.350 19.650 ;
        RECT 54.120 19.620 54.440 19.650 ;
        RECT 68.230 19.630 68.550 19.660 ;
        RECT 47.770 19.530 47.930 19.560 ;
        RECT 16.070 17.930 16.230 17.960 ;
        RECT 13.250 17.840 13.570 17.870 ;
        RECT 14.350 17.840 14.670 17.870 ;
        RECT 15.440 17.840 15.760 17.870 ;
        RECT 13.240 17.650 13.570 17.840 ;
        RECT 14.340 17.650 14.670 17.840 ;
        RECT 15.430 17.750 15.760 17.840 ;
        RECT 13.250 17.610 13.570 17.650 ;
        RECT 14.350 17.610 14.670 17.650 ;
        RECT 13.240 16.500 13.560 16.530 ;
        RECT 13.230 16.310 13.560 16.500 ;
        RECT 14.350 16.490 14.670 16.520 ;
        RECT 13.240 16.270 13.560 16.310 ;
        RECT 14.340 16.300 14.670 16.490 ;
        RECT 14.350 16.260 14.670 16.300 ;
        RECT 12.770 15.440 12.940 16.200 ;
        RECT 13.800 15.800 14.120 15.830 ;
        RECT 13.790 15.610 14.120 15.800 ;
        RECT 13.800 15.570 14.120 15.610 ;
        RECT 14.780 15.820 14.950 17.750 ;
        RECT 15.330 17.610 15.760 17.750 ;
        RECT 15.330 16.500 15.500 17.610 ;
        RECT 15.330 16.240 15.760 16.500 ;
        RECT 14.780 15.560 15.220 15.820 ;
        RECT 14.780 15.250 14.950 15.560 ;
        RECT 15.330 15.250 15.500 16.240 ;
        RECT 15.880 15.820 16.050 17.750 ;
        RECT 15.880 15.560 16.310 15.820 ;
        RECT 15.880 15.250 16.050 15.560 ;
        RECT 16.430 15.250 16.600 17.750 ;
        RECT 16.980 15.250 17.150 17.750 ;
        RECT 17.530 15.250 17.700 17.740 ;
        RECT 46.300 16.920 46.470 19.410 ;
        RECT 46.850 17.390 47.020 19.410 ;
        RECT 47.400 17.390 47.570 19.410 ;
        RECT 47.770 19.190 47.940 19.530 ;
        RECT 48.320 19.520 48.480 19.560 ;
        RECT 47.770 19.180 47.930 19.190 ;
        RECT 47.950 19.150 48.120 19.410 ;
        RECT 48.320 19.190 48.490 19.520 ;
        RECT 48.320 19.180 48.480 19.190 ;
        RECT 47.680 18.890 48.120 19.150 ;
        RECT 47.950 17.780 48.120 18.890 ;
        RECT 47.680 17.520 48.120 17.780 ;
        RECT 46.850 16.910 47.570 17.390 ;
        RECT 47.950 16.910 48.120 17.520 ;
        RECT 48.500 17.100 48.670 19.410 ;
        RECT 48.870 19.190 49.040 19.590 ;
        RECT 49.420 19.520 49.580 19.560 ;
        RECT 49.970 19.520 50.130 19.560 ;
        RECT 50.520 19.540 50.680 19.560 ;
        RECT 52.000 19.540 52.160 19.560 ;
        RECT 48.870 19.180 49.030 19.190 ;
        RECT 49.050 19.150 49.220 19.410 ;
        RECT 49.420 19.190 49.590 19.520 ;
        RECT 49.970 19.190 50.140 19.520 ;
        RECT 50.520 19.190 50.690 19.540 ;
        RECT 51.990 19.190 52.160 19.540 ;
        RECT 52.550 19.520 52.710 19.560 ;
        RECT 53.100 19.520 53.260 19.560 ;
        RECT 52.540 19.190 52.710 19.520 ;
        RECT 53.090 19.190 53.260 19.520 ;
        RECT 49.420 19.180 49.580 19.190 ;
        RECT 49.970 19.180 50.130 19.190 ;
        RECT 50.520 19.180 50.680 19.190 ;
        RECT 52.000 19.180 52.160 19.190 ;
        RECT 52.550 19.180 52.710 19.190 ;
        RECT 53.100 19.180 53.260 19.190 ;
        RECT 53.460 19.150 53.630 19.410 ;
        RECT 53.640 19.190 53.810 19.590 ;
        RECT 57.580 19.560 57.740 19.590 ;
        RECT 54.200 19.520 54.360 19.560 ;
        RECT 54.750 19.530 54.910 19.560 ;
        RECT 53.650 19.180 53.810 19.190 ;
        RECT 48.780 18.890 49.220 19.150 ;
        RECT 49.880 19.110 50.200 19.150 ;
        RECT 52.480 19.110 52.800 19.150 ;
        RECT 49.880 18.920 50.210 19.110 ;
        RECT 52.470 18.920 52.800 19.110 ;
        RECT 49.880 18.890 50.200 18.920 ;
        RECT 52.480 18.890 52.800 18.920 ;
        RECT 53.460 18.890 53.900 19.150 ;
        RECT 49.050 17.780 49.220 18.890 ;
        RECT 53.460 17.780 53.630 18.890 ;
        RECT 48.780 17.520 49.220 17.780 ;
        RECT 49.880 17.740 50.200 17.780 ;
        RECT 52.480 17.740 52.800 17.780 ;
        RECT 49.880 17.550 50.210 17.740 ;
        RECT 52.470 17.550 52.800 17.740 ;
        RECT 49.880 17.520 50.200 17.550 ;
        RECT 52.480 17.520 52.800 17.550 ;
        RECT 53.460 17.520 53.900 17.780 ;
        RECT 48.240 16.910 48.670 17.100 ;
        RECT 49.050 16.910 49.220 17.520 ;
        RECT 49.330 17.060 49.650 17.100 ;
        RECT 50.430 17.070 50.750 17.110 ;
        RECT 51.930 17.070 52.250 17.110 ;
        RECT 47.010 16.380 47.520 16.910 ;
        RECT 48.240 16.870 48.570 16.910 ;
        RECT 49.330 16.870 49.660 17.060 ;
        RECT 50.430 16.880 50.760 17.070 ;
        RECT 51.920 16.880 52.250 17.070 ;
        RECT 53.030 17.060 53.350 17.100 ;
        RECT 48.240 16.840 48.560 16.870 ;
        RECT 49.330 16.840 49.650 16.870 ;
        RECT 50.430 16.850 50.750 16.880 ;
        RECT 51.930 16.850 52.250 16.880 ;
        RECT 53.020 16.870 53.350 17.060 ;
        RECT 53.460 16.910 53.630 17.520 ;
        RECT 54.010 17.100 54.180 19.410 ;
        RECT 54.190 19.190 54.360 19.520 ;
        RECT 54.200 19.180 54.360 19.190 ;
        RECT 54.560 19.150 54.730 19.410 ;
        RECT 54.740 19.190 54.910 19.530 ;
        RECT 56.110 19.410 56.280 19.440 ;
        RECT 54.750 19.180 54.910 19.190 ;
        RECT 54.560 18.890 55.000 19.150 ;
        RECT 54.560 17.780 54.730 18.890 ;
        RECT 54.560 17.520 55.000 17.780 ;
        RECT 54.010 16.910 54.440 17.100 ;
        RECT 54.560 16.910 54.730 17.520 ;
        RECT 55.110 17.390 55.280 19.410 ;
        RECT 55.660 17.390 55.830 19.410 ;
        RECT 55.110 16.910 55.830 17.390 ;
        RECT 56.110 16.950 56.380 19.410 ;
        RECT 56.210 16.920 56.380 16.950 ;
        RECT 56.660 17.420 56.830 19.440 ;
        RECT 57.210 17.420 57.380 19.440 ;
        RECT 57.580 19.220 57.750 19.560 ;
        RECT 58.130 19.550 58.290 19.590 ;
        RECT 57.580 19.210 57.740 19.220 ;
        RECT 57.760 19.180 57.930 19.440 ;
        RECT 58.130 19.220 58.300 19.550 ;
        RECT 58.130 19.210 58.290 19.220 ;
        RECT 57.490 18.920 57.930 19.180 ;
        RECT 57.760 17.810 57.930 18.920 ;
        RECT 57.490 17.550 57.930 17.810 ;
        RECT 56.660 16.940 57.380 17.420 ;
        RECT 57.760 16.940 57.930 17.550 ;
        RECT 58.310 17.130 58.480 19.440 ;
        RECT 58.680 19.220 58.850 19.620 ;
        RECT 59.230 19.550 59.390 19.590 ;
        RECT 59.780 19.550 59.940 19.590 ;
        RECT 60.330 19.570 60.490 19.590 ;
        RECT 61.810 19.570 61.970 19.590 ;
        RECT 58.680 19.210 58.840 19.220 ;
        RECT 58.860 19.180 59.030 19.440 ;
        RECT 59.230 19.220 59.400 19.550 ;
        RECT 59.780 19.220 59.950 19.550 ;
        RECT 60.330 19.220 60.500 19.570 ;
        RECT 61.800 19.220 61.970 19.570 ;
        RECT 62.360 19.550 62.520 19.590 ;
        RECT 62.910 19.550 63.070 19.590 ;
        RECT 62.350 19.220 62.520 19.550 ;
        RECT 62.900 19.220 63.070 19.550 ;
        RECT 59.230 19.210 59.390 19.220 ;
        RECT 59.780 19.210 59.940 19.220 ;
        RECT 60.330 19.210 60.490 19.220 ;
        RECT 61.810 19.210 61.970 19.220 ;
        RECT 62.360 19.210 62.520 19.220 ;
        RECT 62.910 19.210 63.070 19.220 ;
        RECT 63.270 19.180 63.440 19.440 ;
        RECT 63.450 19.220 63.620 19.620 ;
        RECT 64.010 19.550 64.170 19.590 ;
        RECT 64.560 19.560 64.720 19.590 ;
        RECT 63.460 19.210 63.620 19.220 ;
        RECT 58.590 18.920 59.030 19.180 ;
        RECT 59.690 19.140 60.010 19.180 ;
        RECT 62.290 19.140 62.610 19.180 ;
        RECT 59.690 18.950 60.020 19.140 ;
        RECT 62.280 18.950 62.610 19.140 ;
        RECT 59.690 18.920 60.010 18.950 ;
        RECT 62.290 18.920 62.610 18.950 ;
        RECT 63.270 18.920 63.710 19.180 ;
        RECT 58.860 17.810 59.030 18.920 ;
        RECT 63.270 17.810 63.440 18.920 ;
        RECT 58.590 17.550 59.030 17.810 ;
        RECT 59.690 17.770 60.010 17.810 ;
        RECT 62.290 17.770 62.610 17.810 ;
        RECT 59.690 17.580 60.020 17.770 ;
        RECT 62.280 17.580 62.610 17.770 ;
        RECT 59.690 17.550 60.010 17.580 ;
        RECT 62.290 17.550 62.610 17.580 ;
        RECT 63.270 17.550 63.710 17.810 ;
        RECT 58.050 16.940 58.480 17.130 ;
        RECT 58.860 16.940 59.030 17.550 ;
        RECT 59.140 17.090 59.460 17.130 ;
        RECT 60.240 17.100 60.560 17.140 ;
        RECT 61.740 17.100 62.060 17.140 ;
        RECT 54.110 16.870 54.440 16.910 ;
        RECT 53.030 16.840 53.350 16.870 ;
        RECT 54.120 16.840 54.440 16.870 ;
        RECT 55.160 16.380 55.670 16.910 ;
        RECT 56.820 16.410 57.330 16.940 ;
        RECT 58.050 16.900 58.380 16.940 ;
        RECT 59.140 16.900 59.470 17.090 ;
        RECT 60.240 16.910 60.570 17.100 ;
        RECT 61.730 16.910 62.060 17.100 ;
        RECT 62.840 17.090 63.160 17.130 ;
        RECT 58.050 16.870 58.370 16.900 ;
        RECT 59.140 16.870 59.460 16.900 ;
        RECT 60.240 16.880 60.560 16.910 ;
        RECT 61.740 16.880 62.060 16.910 ;
        RECT 62.830 16.900 63.160 17.090 ;
        RECT 63.270 16.940 63.440 17.550 ;
        RECT 63.820 17.130 63.990 19.440 ;
        RECT 64.000 19.220 64.170 19.550 ;
        RECT 64.010 19.210 64.170 19.220 ;
        RECT 64.370 19.180 64.540 19.440 ;
        RECT 64.550 19.220 64.720 19.560 ;
        RECT 64.560 19.210 64.720 19.220 ;
        RECT 64.370 18.920 64.810 19.180 ;
        RECT 64.370 17.810 64.540 18.920 ;
        RECT 64.370 17.550 64.810 17.810 ;
        RECT 63.820 16.940 64.250 17.130 ;
        RECT 64.370 16.940 64.540 17.550 ;
        RECT 64.920 17.420 65.090 19.440 ;
        RECT 65.470 17.420 65.640 19.440 ;
        RECT 64.920 16.940 65.640 17.420 ;
        RECT 66.020 16.950 66.190 19.440 ;
        RECT 68.300 17.120 68.470 19.630 ;
        RECT 68.850 19.160 69.020 21.670 ;
        RECT 69.400 21.240 69.570 21.970 ;
        RECT 69.950 21.940 70.120 21.970 ;
        RECT 69.880 21.900 70.200 21.940 ;
        RECT 69.870 21.710 70.200 21.900 ;
        RECT 69.880 21.680 70.200 21.710 ;
        RECT 69.330 21.200 69.650 21.240 ;
        RECT 69.320 21.010 69.650 21.200 ;
        RECT 69.330 20.980 69.650 21.010 ;
        RECT 69.400 19.890 69.570 20.980 ;
        RECT 69.330 19.850 69.650 19.890 ;
        RECT 69.320 19.660 69.650 19.850 ;
        RECT 69.330 19.630 69.650 19.660 ;
        RECT 68.780 19.120 69.100 19.160 ;
        RECT 68.770 18.930 69.100 19.120 ;
        RECT 68.780 18.900 69.100 18.930 ;
        RECT 68.850 17.790 69.020 18.900 ;
        RECT 68.780 17.750 69.100 17.790 ;
        RECT 68.770 17.560 69.100 17.750 ;
        RECT 68.780 17.530 69.100 17.560 ;
        RECT 68.230 17.080 68.550 17.120 ;
        RECT 63.920 16.900 64.250 16.940 ;
        RECT 62.840 16.870 63.160 16.900 ;
        RECT 63.930 16.870 64.250 16.900 ;
        RECT 64.970 16.410 65.480 16.940 ;
        RECT 68.220 16.890 68.550 17.080 ;
        RECT 68.230 16.860 68.550 16.890 ;
        RECT 68.300 16.790 68.470 16.860 ;
        RECT 68.850 16.790 69.020 17.530 ;
        RECT 69.400 17.110 69.570 19.630 ;
        RECT 69.950 19.160 70.120 21.680 ;
        RECT 70.500 21.260 70.670 21.970 ;
        RECT 71.050 21.940 71.220 21.970 ;
        RECT 70.970 21.900 71.290 21.940 ;
        RECT 70.960 21.710 71.290 21.900 ;
        RECT 70.970 21.680 71.290 21.710 ;
        RECT 70.420 21.220 70.740 21.260 ;
        RECT 70.410 21.030 70.740 21.220 ;
        RECT 70.420 21.000 70.740 21.030 ;
        RECT 70.500 19.890 70.670 21.000 ;
        RECT 70.420 19.850 70.740 19.890 ;
        RECT 70.410 19.660 70.740 19.850 ;
        RECT 70.420 19.630 70.740 19.660 ;
        RECT 69.880 19.120 70.200 19.160 ;
        RECT 69.870 18.930 70.200 19.120 ;
        RECT 69.880 18.900 70.200 18.930 ;
        RECT 69.950 17.790 70.120 18.900 ;
        RECT 69.880 17.750 70.200 17.790 ;
        RECT 69.870 17.560 70.200 17.750 ;
        RECT 69.880 17.530 70.200 17.560 ;
        RECT 69.330 17.070 69.650 17.110 ;
        RECT 69.320 16.880 69.650 17.070 ;
        RECT 69.330 16.850 69.650 16.880 ;
        RECT 69.400 16.790 69.570 16.850 ;
        RECT 69.950 16.790 70.120 17.530 ;
        RECT 70.500 17.110 70.670 19.630 ;
        RECT 71.050 19.160 71.220 21.680 ;
        RECT 70.980 19.120 71.300 19.160 ;
        RECT 70.970 18.930 71.300 19.120 ;
        RECT 70.980 18.900 71.300 18.930 ;
        RECT 71.050 17.790 71.220 18.900 ;
        RECT 70.980 17.750 71.300 17.790 ;
        RECT 70.970 17.560 71.300 17.750 ;
        RECT 71.760 17.590 71.930 18.780 ;
        RECT 70.980 17.530 71.300 17.560 ;
        RECT 70.420 17.070 70.740 17.110 ;
        RECT 70.410 16.880 70.740 17.070 ;
        RECT 70.420 16.850 70.740 16.880 ;
        RECT 70.500 16.790 70.670 16.850 ;
        RECT 71.050 16.790 71.220 17.530 ;
        RECT 71.470 17.140 71.980 17.400 ;
        RECT 71.460 17.070 71.980 17.140 ;
        RECT 71.460 16.390 71.970 17.070 ;
        RECT 18.170 15.280 20.560 15.650 ;
        RECT 18.220 12.020 20.560 15.280 ;
        RECT 96.970 14.480 97.200 14.490 ;
        RECT 96.950 14.310 101.610 14.480 ;
        RECT 96.970 14.300 97.200 14.310 ;
        RECT 102.510 13.830 102.700 13.840 ;
        RECT 98.170 13.790 101.970 13.800 ;
        RECT 102.480 13.790 102.740 13.830 ;
        RECT 98.170 13.630 102.740 13.790 ;
        RECT 101.740 13.620 102.740 13.630 ;
        RECT 101.740 13.160 101.970 13.620 ;
        RECT 102.480 13.510 102.740 13.620 ;
        RECT 102.510 13.160 102.700 13.170 ;
        RECT 101.740 12.950 102.750 13.160 ;
        RECT 96.970 12.870 97.200 12.880 ;
        RECT 96.950 12.700 101.430 12.870 ;
        RECT 96.970 12.690 97.200 12.700 ;
        RECT 101.740 12.190 101.970 12.950 ;
        RECT 102.480 12.840 102.740 12.950 ;
        RECT 98.190 12.020 101.970 12.190 ;
        RECT 18.220 12.010 20.550 12.020 ;
        RECT 96.970 11.270 97.200 11.280 ;
        RECT 96.950 11.100 101.450 11.270 ;
        RECT 96.970 11.090 97.200 11.100 ;
        RECT 98.190 11.090 98.520 11.100 ;
        RECT 99.150 11.090 99.480 11.100 ;
        RECT 100.110 11.090 100.440 11.100 ;
        RECT 101.070 11.090 101.400 11.100 ;
        RECT 101.740 10.580 101.970 12.020 ;
        RECT 102.420 11.830 102.850 11.850 ;
        RECT 102.400 11.660 102.850 11.830 ;
        RECT 102.420 11.640 102.850 11.660 ;
        RECT 98.190 10.410 101.970 10.580 ;
        RECT 98.250 10.180 98.680 10.200 ;
        RECT 98.230 10.010 98.680 10.180 ;
        RECT 98.250 9.990 98.680 10.010 ;
        RECT 96.970 9.650 97.200 9.660 ;
        RECT 96.950 9.480 101.450 9.650 ;
        RECT 96.970 9.470 97.200 9.480 ;
        RECT 101.740 8.980 101.970 10.410 ;
        RECT 102.420 10.220 102.850 10.240 ;
        RECT 102.400 10.050 102.850 10.220 ;
        RECT 102.420 10.030 102.850 10.050 ;
        RECT 98.200 8.970 101.970 8.980 ;
        RECT 98.190 8.810 101.970 8.970 ;
        RECT 98.190 8.800 98.520 8.810 ;
        RECT 100.110 8.800 100.440 8.810 ;
        RECT 101.070 8.800 101.400 8.810 ;
        RECT 99.250 8.440 99.680 8.460 ;
        RECT 99.250 8.270 99.700 8.440 ;
        RECT 99.250 8.250 99.680 8.270 ;
        RECT 96.970 8.050 97.200 8.060 ;
        RECT 96.950 7.880 101.400 8.050 ;
        RECT 96.970 7.870 97.200 7.880 ;
        RECT 98.190 7.870 98.520 7.880 ;
        RECT 99.150 7.870 99.480 7.880 ;
        RECT 100.110 7.870 100.440 7.880 ;
        RECT 101.070 7.870 101.400 7.880 ;
        RECT 101.740 7.360 101.970 8.810 ;
        RECT 102.410 8.610 102.840 8.630 ;
        RECT 102.390 8.440 102.840 8.610 ;
        RECT 102.410 8.420 102.840 8.440 ;
        RECT 98.180 7.190 101.970 7.360 ;
        RECT 100.160 6.930 100.590 6.950 ;
        RECT 100.140 6.760 100.590 6.930 ;
        RECT 100.160 6.740 100.590 6.760 ;
        RECT 96.970 6.430 97.200 6.440 ;
        RECT 96.950 6.260 101.450 6.430 ;
        RECT 96.970 6.250 97.200 6.260 ;
        RECT 98.190 5.740 98.520 5.750 ;
        RECT 99.150 5.740 99.480 5.750 ;
        RECT 100.110 5.740 100.440 5.750 ;
        RECT 101.070 5.740 101.400 5.750 ;
        RECT 101.740 5.740 101.970 7.190 ;
        RECT 102.410 6.990 102.840 7.010 ;
        RECT 102.390 6.820 102.840 6.990 ;
        RECT 102.410 6.800 102.840 6.820 ;
        RECT 98.180 5.570 101.970 5.740 ;
        RECT 96.970 4.830 97.200 4.840 ;
        RECT 96.950 4.820 101.370 4.830 ;
        RECT 96.950 4.660 101.400 4.820 ;
        RECT 96.970 4.650 97.200 4.660 ;
        RECT 98.190 4.650 98.520 4.660 ;
        RECT 99.150 4.650 99.480 4.660 ;
        RECT 100.110 4.650 100.440 4.660 ;
        RECT 101.070 4.650 101.400 4.660 ;
        RECT 101.740 4.150 101.970 5.570 ;
        RECT 102.410 5.380 102.840 5.400 ;
        RECT 102.390 5.210 102.840 5.380 ;
        RECT 102.410 5.190 102.840 5.210 ;
        RECT 108.400 5.020 108.770 19.890 ;
        RECT 108.400 4.770 108.780 5.020 ;
        RECT 98.180 3.980 101.980 4.150 ;
        RECT 98.190 3.970 98.520 3.980 ;
        RECT 99.150 3.970 99.480 3.980 ;
        RECT 100.110 3.970 100.440 3.980 ;
        RECT 101.070 3.970 101.400 3.980 ;
        RECT 96.970 3.200 97.200 3.220 ;
        RECT 98.190 3.200 98.520 3.210 ;
        RECT 99.150 3.200 99.480 3.210 ;
        RECT 100.110 3.200 100.440 3.210 ;
        RECT 101.070 3.200 101.400 3.210 ;
        RECT 96.950 3.030 101.410 3.200 ;
        RECT 101.740 2.540 101.970 3.980 ;
        RECT 102.250 3.390 102.460 3.820 ;
        RECT 102.270 3.370 102.440 3.390 ;
        RECT 98.180 2.370 101.970 2.540 ;
        RECT 98.190 2.360 98.520 2.370 ;
        RECT 99.150 2.360 99.480 2.370 ;
        RECT 100.110 2.360 100.440 2.370 ;
        RECT 101.070 2.360 101.400 2.370 ;
        RECT 102.420 2.180 102.850 2.200 ;
        RECT 102.400 2.010 102.850 2.180 ;
        RECT 102.420 1.990 102.850 2.010 ;
        RECT 102.410 0.590 102.840 0.610 ;
        RECT 99.210 0.510 99.640 0.530 ;
        RECT 100.150 0.510 100.580 0.530 ;
        RECT 99.190 0.340 99.640 0.510 ;
        RECT 100.130 0.340 100.580 0.510 ;
        RECT 101.100 0.450 101.530 0.470 ;
        RECT 99.210 0.320 99.640 0.340 ;
        RECT 100.150 0.320 100.580 0.340 ;
        RECT 101.080 0.280 101.530 0.450 ;
        RECT 102.390 0.420 102.840 0.590 ;
        RECT 102.410 0.400 102.840 0.420 ;
        RECT 101.100 0.260 101.530 0.280 ;
      LAYER mcon ;
        RECT 4.490 71.380 4.660 71.550 ;
        RECT 7.360 71.590 7.530 71.760 ;
        RECT 5.900 71.380 6.070 71.550 ;
        RECT 22.700 71.410 22.870 71.580 ;
        RECT 22.700 71.060 22.870 71.230 ;
        RECT 7.360 70.800 7.530 70.970 ;
        RECT 22.700 70.720 22.870 70.890 ;
        RECT 28.560 71.320 28.730 71.490 ;
        RECT 28.560 70.870 28.730 71.040 ;
        RECT 33.260 71.270 33.430 71.440 ;
        RECT 33.260 70.820 33.430 70.990 ;
        RECT 4.490 70.530 4.660 70.700 ;
        RECT 5.210 70.520 5.380 70.690 ;
        RECT 5.900 70.530 6.070 70.700 ;
        RECT 4.670 70.120 4.840 70.290 ;
        RECT 5.730 70.120 5.900 70.290 ;
        RECT 4.490 69.710 4.660 69.880 ;
        RECT 5.210 69.680 5.380 69.850 ;
        RECT 5.900 69.710 6.070 69.880 ;
        RECT 20.600 69.780 20.770 69.950 ;
        RECT 21.960 69.860 22.130 70.030 ;
        RECT 22.650 69.850 22.820 70.020 ;
        RECT 7.360 69.370 7.530 69.540 ;
        RECT 4.490 68.870 4.660 69.040 ;
        RECT 5.900 68.870 6.070 69.040 ;
        RECT 6.630 68.610 6.800 68.780 ;
        RECT 6.620 68.090 6.790 68.260 ;
        RECT 7.370 67.970 7.540 68.140 ;
        RECT 4.490 67.750 4.660 67.920 ;
        RECT 5.900 67.750 6.070 67.920 ;
        RECT 5.190 66.880 5.360 67.050 ;
        RECT 6.620 66.900 6.790 67.070 ;
        RECT 9.380 66.550 9.550 66.720 ;
        RECT 4.400 66.300 4.570 66.470 ;
        RECT 5.330 66.300 5.500 66.470 ;
        RECT 6.030 66.300 6.200 66.470 ;
        RECT 6.770 66.300 6.940 66.470 ;
        RECT 7.480 66.290 7.650 66.460 ;
        RECT 22.700 68.610 22.870 68.780 ;
        RECT 22.700 68.260 22.870 68.430 ;
        RECT 22.700 67.920 22.870 68.090 ;
        RECT 28.560 68.330 28.730 68.500 ;
        RECT 28.560 67.880 28.730 68.050 ;
        RECT 28.560 67.320 28.730 67.490 ;
        RECT 22.700 67.060 22.870 67.230 ;
        RECT 22.700 66.710 22.870 66.880 ;
        RECT 28.560 66.870 28.730 67.040 ;
        RECT 22.700 66.370 22.870 66.540 ;
        RECT 32.480 67.810 32.650 67.980 ;
        RECT 19.880 66.120 20.050 66.290 ;
        RECT 29.740 66.140 29.910 66.310 ;
        RECT 19.890 61.760 20.320 62.500 ;
        RECT 40.590 60.600 40.800 60.810 ;
        RECT 45.470 60.710 45.640 60.880 ;
        RECT 39.120 60.230 39.290 60.400 ;
        RECT 46.510 60.360 46.680 60.530 ;
        RECT 46.510 60.010 46.680 60.180 ;
        RECT 40.590 59.050 40.800 59.260 ;
        RECT 45.470 59.160 45.640 59.330 ;
        RECT 39.120 58.680 39.290 58.850 ;
        RECT 15.870 58.380 16.040 58.550 ;
        RECT 16.960 58.390 17.130 58.560 ;
        RECT 46.510 58.810 46.680 58.980 ;
        RECT 46.510 58.460 46.680 58.630 ;
        RECT 68.180 58.600 68.440 59.420 ;
        RECT 80.130 58.630 80.450 59.420 ;
        RECT 82.410 58.960 82.590 59.130 ;
        RECT 82.840 58.940 83.010 59.110 ;
        RECT 80.600 58.660 80.770 58.830 ;
        RECT 15.650 57.970 15.820 58.140 ;
        RECT 17.800 57.920 17.970 58.090 ;
        RECT 80.950 57.820 81.130 58.010 ;
        RECT 15.870 57.460 16.040 57.630 ;
        RECT 16.960 57.470 17.130 57.640 ;
        RECT 40.590 57.500 40.800 57.710 ;
        RECT 45.470 57.610 45.640 57.780 ;
        RECT 15.650 57.050 15.820 57.220 ;
        RECT 39.120 57.130 39.290 57.300 ;
        RECT 15.870 56.540 16.040 56.710 ;
        RECT 16.960 56.550 17.130 56.720 ;
        RECT 46.510 57.260 46.680 57.430 ;
        RECT 46.510 56.910 46.680 57.080 ;
        RECT 83.310 58.380 83.480 58.550 ;
        RECT 110.470 58.660 110.640 58.830 ;
        RECT 85.550 58.080 85.720 58.250 ;
        RECT 103.630 58.080 103.800 58.250 ;
        RECT 85.550 57.630 85.720 57.800 ;
        RECT 82.030 57.260 82.200 57.430 ;
        RECT 91.000 57.480 91.270 57.750 ;
        RECT 99.970 57.480 100.240 57.750 ;
        RECT 103.630 57.630 103.800 57.800 ;
        RECT 108.800 57.830 108.970 58.000 ;
        RECT 82.840 56.950 83.010 57.120 ;
        RECT 15.650 56.130 15.820 56.300 ;
        RECT 40.590 55.950 40.800 56.160 ;
        RECT 45.470 56.060 45.640 56.230 ;
        RECT 110.110 57.820 110.290 58.010 ;
        RECT 88.680 56.370 88.850 56.540 ;
        RECT 102.390 56.370 102.560 56.540 ;
        RECT 15.680 55.560 15.850 55.730 ;
        RECT 16.980 55.460 17.150 55.630 ;
        RECT 39.120 55.580 39.290 55.750 ;
        RECT 46.510 55.710 46.680 55.880 ;
        RECT 46.510 55.360 46.680 55.530 ;
        RECT 80.950 55.020 81.130 55.210 ;
        RECT 15.680 54.600 15.850 54.770 ;
        RECT 16.980 54.500 17.150 54.670 ;
        RECT 83.310 56.060 83.480 56.230 ;
        RECT 82.850 55.880 83.020 56.050 ;
        RECT 82.020 55.570 82.190 55.740 ;
        RECT 91.000 55.750 91.270 56.020 ;
        RECT 99.970 55.750 100.240 56.020 ;
        RECT 85.550 55.130 85.720 55.300 ;
        RECT 85.550 54.680 85.720 54.850 ;
        RECT 103.630 55.130 103.800 55.300 ;
        RECT 107.330 55.480 107.500 55.650 ;
        RECT 108.410 55.510 108.580 55.620 ;
        RECT 108.290 55.450 108.580 55.510 ;
        RECT 108.290 55.340 108.460 55.450 ;
        RECT 108.900 55.480 109.070 55.650 ;
        RECT 108.800 55.070 108.970 55.240 ;
        RECT 109.420 55.350 109.590 55.520 ;
        RECT 109.380 55.170 109.550 55.340 ;
        RECT 110.110 55.020 110.290 55.210 ;
        RECT 111.630 55.220 111.800 55.390 ;
        RECT 103.630 54.680 103.800 54.850 ;
        RECT 105.880 54.700 106.050 54.870 ;
        RECT 106.380 54.730 106.550 54.900 ;
        RECT 83.300 54.480 83.470 54.650 ;
        RECT 80.600 54.200 80.770 54.370 ;
        RECT 108.560 54.620 108.730 54.790 ;
        RECT 109.880 54.730 110.050 54.900 ;
        RECT 110.360 54.850 110.530 55.020 ;
        RECT 82.410 53.900 82.590 54.070 ;
        RECT 82.870 53.970 83.040 54.140 ;
        RECT 107.440 54.100 107.610 54.270 ;
        RECT 15.680 53.640 15.850 53.810 ;
        RECT 109.330 54.520 109.500 54.690 ;
        RECT 110.470 54.200 110.640 54.370 ;
        RECT 108.650 53.900 108.830 54.070 ;
        RECT 106.380 53.730 106.550 53.900 ;
        RECT 16.980 53.540 17.150 53.710 ;
        RECT 58.470 53.310 58.640 53.480 ;
        RECT 17.380 53.100 17.550 53.270 ;
        RECT 59.310 53.190 59.480 53.360 ;
        RECT 60.060 53.190 60.230 53.360 ;
        RECT 39.120 52.050 39.290 52.220 ;
        RECT 46.510 52.270 46.680 52.440 ;
        RECT 63.040 52.860 63.210 53.030 ;
        RECT 58.750 52.560 58.920 52.730 ;
        RECT 63.440 53.310 63.610 53.480 ;
        RECT 63.440 52.970 63.610 53.140 ;
        RECT 82.410 52.930 82.590 53.100 ;
        RECT 80.600 52.630 80.770 52.800 ;
        RECT 40.590 51.640 40.800 51.850 ;
        RECT 46.510 51.920 46.680 52.090 ;
        RECT 45.470 51.570 45.640 51.740 ;
        RECT 58.750 51.670 58.920 51.840 ;
        RECT 80.950 51.790 81.130 51.980 ;
        RECT 63.040 51.370 63.210 51.540 ;
        RECT 39.120 50.500 39.290 50.670 ;
        RECT 59.310 51.040 59.480 51.210 ;
        RECT 60.060 51.040 60.230 51.210 ;
        RECT 62.060 51.050 62.230 51.220 ;
        RECT 63.440 51.600 63.610 51.770 ;
        RECT 63.440 51.260 63.610 51.430 ;
        RECT 46.510 50.720 46.680 50.890 ;
        RECT 109.330 53.700 109.500 53.870 ;
        RECT 109.880 53.730 110.050 53.900 ;
        RECT 111.020 53.910 111.190 54.080 ;
        RECT 110.360 53.370 110.530 53.540 ;
        RECT 107.330 52.980 107.500 53.150 ;
        RECT 108.290 53.120 108.460 53.290 ;
        RECT 109.420 53.220 109.590 53.280 ;
        RECT 108.170 52.820 108.340 52.990 ;
        RECT 108.900 52.980 109.070 53.150 ;
        RECT 109.380 53.110 109.590 53.220 ;
        RECT 109.380 53.050 109.550 53.110 ;
        RECT 111.680 53.000 111.850 53.170 ;
        RECT 87.440 52.050 87.610 52.220 ;
        RECT 89.530 52.210 89.700 52.380 ;
        RECT 107.330 52.460 107.500 52.630 ;
        RECT 82.270 51.800 82.440 51.970 ;
        RECT 103.630 52.050 103.800 52.220 ;
        RECT 108.290 52.320 108.460 52.490 ;
        RECT 108.900 52.460 109.070 52.630 ;
        RECT 110.470 52.630 110.640 52.800 ;
        RECT 87.440 51.600 87.610 51.770 ;
        RECT 91.000 51.450 91.270 51.720 ;
        RECT 99.970 51.450 100.240 51.720 ;
        RECT 108.600 52.020 108.770 52.190 ;
        RECT 109.420 52.380 109.590 52.500 ;
        RECT 109.380 52.330 109.590 52.380 ;
        RECT 109.380 52.210 109.550 52.330 ;
        RECT 103.630 51.600 103.800 51.770 ;
        RECT 105.880 51.680 106.050 51.850 ;
        RECT 106.380 51.710 106.550 51.880 ;
        RECT 108.800 51.800 108.970 51.970 ;
        RECT 111.670 52.280 111.840 52.450 ;
        RECT 40.590 50.090 40.800 50.300 ;
        RECT 46.510 50.370 46.680 50.540 ;
        RECT 58.470 50.380 58.640 50.550 ;
        RECT 45.470 50.020 45.640 50.190 ;
        RECT 59.310 50.260 59.480 50.430 ;
        RECT 60.060 50.260 60.230 50.430 ;
        RECT 39.120 48.950 39.290 49.120 ;
        RECT 63.040 49.930 63.210 50.100 ;
        RECT 58.750 49.630 58.920 49.800 ;
        RECT 63.440 50.380 63.610 50.550 ;
        RECT 63.440 50.040 63.610 50.210 ;
        RECT 109.330 51.560 109.500 51.730 ;
        RECT 109.880 51.710 110.050 51.880 ;
        RECT 110.110 51.790 110.290 51.980 ;
        RECT 110.360 51.890 110.530 52.060 ;
        RECT 111.020 51.320 111.190 51.490 ;
        RECT 106.380 50.710 106.550 50.880 ;
        RECT 109.330 50.740 109.500 50.910 ;
        RECT 109.730 50.880 109.910 50.940 ;
        RECT 109.730 50.750 110.050 50.880 ;
        RECT 88.680 50.340 88.850 50.510 ;
        RECT 102.390 50.340 102.560 50.510 ;
        RECT 46.510 49.170 46.680 49.340 ;
        RECT 40.590 48.540 40.800 48.750 ;
        RECT 46.510 48.820 46.680 48.990 ;
        RECT 80.950 48.990 81.130 49.180 ;
        RECT 45.470 48.470 45.640 48.640 ;
        RECT 58.750 48.740 58.920 48.910 ;
        RECT 63.040 48.440 63.210 48.610 ;
        RECT 59.310 48.110 59.480 48.280 ;
        RECT 60.060 48.110 60.230 48.280 ;
        RECT 62.060 48.120 62.230 48.290 ;
        RECT 63.440 48.670 63.610 48.840 ;
        RECT 63.440 48.330 63.610 48.500 ;
        RECT 91.000 49.720 91.270 49.990 ;
        RECT 99.970 49.720 100.240 49.990 ;
        RECT 109.880 50.710 110.050 50.750 ;
        RECT 110.360 50.410 110.530 50.580 ;
        RECT 107.330 49.960 107.500 50.130 ;
        RECT 108.290 50.100 108.460 50.270 ;
        RECT 108.900 49.960 109.070 50.130 ;
        RECT 109.380 50.090 109.590 50.260 ;
        RECT 109.730 50.030 109.910 50.220 ;
        RECT 111.590 50.030 111.760 50.200 ;
        RECT 108.410 49.420 108.580 49.590 ;
        RECT 82.270 49.040 82.440 49.210 ;
        RECT 87.440 49.100 87.610 49.270 ;
        RECT 87.440 48.650 87.610 48.820 ;
        RECT 103.630 49.100 103.800 49.270 ;
        RECT 89.560 48.520 89.730 48.690 ;
        RECT 103.630 48.650 103.800 48.820 ;
        RECT 80.600 48.170 80.770 48.340 ;
        RECT 39.120 47.400 39.290 47.570 ;
        RECT 82.410 47.870 82.590 48.040 ;
        RECT 46.510 47.620 46.680 47.790 ;
        RECT 40.590 46.990 40.800 47.200 ;
        RECT 108.800 49.040 108.970 49.210 ;
        RECT 109.380 49.140 109.550 49.310 ;
        RECT 108.560 48.590 108.730 48.760 ;
        RECT 107.440 48.070 107.610 48.240 ;
        RECT 46.510 47.270 46.680 47.440 ;
        RECT 45.470 46.920 45.640 47.090 ;
        RECT 67.730 46.980 67.900 47.150 ;
        RECT 88.500 46.980 88.670 47.150 ;
        RECT 65.920 46.720 66.090 46.890 ;
        RECT 66.650 46.690 66.820 46.860 ;
        RECT 89.580 46.690 89.750 46.860 ;
        RECT 67.730 46.430 67.900 46.600 ;
        RECT 88.500 46.430 88.670 46.600 ;
        RECT 68.640 46.180 68.810 46.350 ;
        RECT 72.580 46.190 72.750 46.360 ;
        RECT 83.650 46.190 83.820 46.360 ;
        RECT 87.590 46.180 87.760 46.350 ;
        RECT 90.310 46.720 90.480 46.890 ;
        RECT 92.640 46.870 92.810 47.040 ;
        RECT 92.650 46.180 92.820 46.350 ;
        RECT 98.430 46.870 98.600 47.040 ;
        RECT 98.430 46.190 98.600 46.360 ;
        RECT 65.920 45.270 66.090 45.440 ;
        RECT 67.730 45.560 67.900 45.730 ;
        RECT 88.500 45.560 88.670 45.730 ;
        RECT 66.650 45.300 66.820 45.470 ;
        RECT 89.580 45.300 89.750 45.470 ;
        RECT 90.310 45.270 90.480 45.440 ;
        RECT 67.730 45.010 67.900 45.180 ;
        RECT 68.640 44.590 68.810 44.760 ;
        RECT 72.570 44.730 72.740 44.900 ;
        RECT 88.500 45.010 88.670 45.180 ;
        RECT 68.640 44.250 68.810 44.420 ;
        RECT 70.850 44.360 71.120 44.630 ;
        RECT 72.570 44.390 72.740 44.560 ;
        RECT 67.730 43.970 67.900 44.140 ;
        RECT 74.880 44.430 75.150 44.700 ;
        RECT 81.250 44.430 81.520 44.700 ;
        RECT 83.660 44.730 83.830 44.900 ;
        RECT 83.660 44.390 83.830 44.560 ;
        RECT 85.280 44.360 85.550 44.630 ;
        RECT 87.590 44.590 87.760 44.760 ;
        RECT 89.950 44.490 90.130 44.660 ;
        RECT 87.590 44.250 87.760 44.420 ;
        RECT 88.500 43.970 88.670 44.140 ;
        RECT 110.110 48.990 110.290 49.180 ;
        RECT 111.630 49.190 111.800 49.360 ;
        RECT 109.330 48.490 109.500 48.660 ;
        RECT 110.360 48.820 110.530 48.990 ;
        RECT 110.470 48.170 110.640 48.340 ;
        RECT 109.330 47.670 109.500 47.840 ;
        RECT 111.020 47.880 111.190 48.050 ;
        RECT 110.360 47.340 110.530 47.510 ;
        RECT 109.380 47.020 109.550 47.190 ;
        RECT 108.170 46.790 108.340 46.960 ;
        RECT 111.680 46.970 111.850 47.140 ;
        RECT 108.600 45.990 108.770 46.160 ;
        RECT 109.380 46.180 109.550 46.350 ;
        RECT 111.670 46.250 111.840 46.420 ;
        RECT 110.360 45.860 110.530 46.030 ;
        RECT 109.330 45.530 109.500 45.700 ;
        RECT 111.020 45.290 111.190 45.460 ;
        RECT 109.330 44.710 109.500 44.880 ;
        RECT 110.360 44.380 110.530 44.550 ;
        RECT 109.380 44.060 109.550 44.230 ;
        RECT 111.590 44.000 111.760 44.170 ;
        RECT 65.920 43.710 66.090 43.880 ;
        RECT 58.470 43.240 58.640 43.410 ;
        RECT 59.310 43.120 59.480 43.290 ;
        RECT 60.060 43.120 60.230 43.290 ;
        RECT 39.120 41.920 39.290 42.090 ;
        RECT 46.510 42.140 46.680 42.310 ;
        RECT 63.040 42.790 63.210 42.960 ;
        RECT 58.750 42.490 58.920 42.660 ;
        RECT 63.440 43.240 63.610 43.410 ;
        RECT 66.650 43.680 66.820 43.850 ;
        RECT 89.580 43.680 89.750 43.850 ;
        RECT 67.730 43.420 67.900 43.590 ;
        RECT 88.500 43.420 88.670 43.590 ;
        RECT 90.310 43.710 90.480 43.880 ;
        RECT 63.440 42.900 63.610 43.070 ;
        RECT 65.920 42.270 66.090 42.440 ;
        RECT 67.730 42.560 67.900 42.730 ;
        RECT 88.500 42.560 88.670 42.730 ;
        RECT 66.650 42.300 66.820 42.470 ;
        RECT 89.580 42.300 89.750 42.470 ;
        RECT 90.310 42.270 90.480 42.440 ;
        RECT 40.590 41.510 40.800 41.720 ;
        RECT 46.510 41.790 46.680 41.960 ;
        RECT 45.470 41.440 45.640 41.610 ;
        RECT 67.730 42.010 67.900 42.180 ;
        RECT 88.500 42.010 88.670 42.180 ;
        RECT 58.750 41.600 58.920 41.770 ;
        RECT 63.040 41.300 63.210 41.470 ;
        RECT 39.120 40.370 39.290 40.540 ;
        RECT 59.310 40.970 59.480 41.140 ;
        RECT 60.060 40.970 60.230 41.140 ;
        RECT 62.060 40.980 62.230 41.150 ;
        RECT 63.440 41.530 63.610 41.700 ;
        RECT 63.440 41.190 63.610 41.360 ;
        RECT 46.510 40.590 46.680 40.760 ;
        RECT 40.590 39.960 40.800 40.170 ;
        RECT 46.510 40.240 46.680 40.410 ;
        RECT 58.470 40.310 58.640 40.480 ;
        RECT 45.470 39.890 45.640 40.060 ;
        RECT 59.310 40.190 59.480 40.360 ;
        RECT 60.060 40.190 60.230 40.360 ;
        RECT 39.120 38.820 39.290 38.990 ;
        RECT 63.040 39.860 63.210 40.030 ;
        RECT 58.750 39.560 58.920 39.730 ;
        RECT 63.440 40.310 63.610 40.480 ;
        RECT 63.440 39.970 63.610 40.140 ;
        RECT 46.510 39.040 46.680 39.210 ;
        RECT 40.590 38.410 40.800 38.620 ;
        RECT 46.510 38.690 46.680 38.860 ;
        RECT 45.470 38.340 45.640 38.510 ;
        RECT 58.750 38.670 58.920 38.840 ;
        RECT 63.040 38.370 63.210 38.540 ;
        RECT 59.310 38.040 59.480 38.210 ;
        RECT 60.060 38.040 60.230 38.210 ;
        RECT 62.060 38.050 62.230 38.220 ;
        RECT 63.440 38.600 63.610 38.770 ;
        RECT 63.440 38.260 63.610 38.430 ;
        RECT 39.120 37.270 39.290 37.440 ;
        RECT 46.510 37.490 46.680 37.660 ;
        RECT 68.310 37.590 68.480 37.760 ;
        RECT 40.590 36.860 40.800 37.070 ;
        RECT 46.510 37.140 46.680 37.310 ;
        RECT 66.500 37.330 66.670 37.500 ;
        RECT 45.470 36.790 45.640 36.960 ;
        RECT 67.230 37.300 67.400 37.470 ;
        RECT 68.310 37.040 68.480 37.210 ;
        RECT 69.350 36.770 69.520 36.940 ;
        RECT 66.500 35.880 66.670 36.050 ;
        RECT 73.370 36.800 73.540 36.970 ;
        RECT 68.310 36.170 68.480 36.340 ;
        RECT 67.230 35.910 67.400 36.080 ;
        RECT 68.310 35.620 68.480 35.790 ;
        RECT 69.340 35.590 69.510 35.760 ;
        RECT 69.340 35.250 69.510 35.420 ;
        RECT 73.360 35.530 73.530 35.700 ;
        RECT 69.340 34.910 69.510 35.080 ;
        RECT 16.710 34.410 16.880 34.580 ;
        RECT 17.360 34.410 17.530 34.580 ;
        RECT 68.310 34.580 68.480 34.750 ;
        RECT 71.430 34.970 71.700 35.240 ;
        RECT 73.360 35.190 73.530 35.360 ;
        RECT 73.360 34.850 73.530 35.020 ;
        RECT 75.460 35.040 75.730 35.310 ;
        RECT 15.490 33.970 15.660 34.140 ;
        RECT 16.190 33.970 16.360 34.140 ;
        RECT 15.040 32.310 15.210 32.480 ;
        RECT 66.500 34.320 66.670 34.490 ;
        RECT 67.230 34.290 67.400 34.460 ;
        RECT 68.310 34.030 68.480 34.200 ;
        RECT 17.870 33.590 18.040 33.760 ;
        RECT 79.650 33.690 79.820 33.860 ;
        RECT 17.870 33.250 18.040 33.420 ;
        RECT 58.470 33.480 58.640 33.650 ;
        RECT 59.310 33.360 59.480 33.530 ;
        RECT 60.060 33.360 60.230 33.530 ;
        RECT 18.040 32.110 18.210 32.280 ;
        RECT 39.120 32.150 39.290 32.320 ;
        RECT 46.510 32.370 46.680 32.540 ;
        RECT 63.040 33.030 63.210 33.200 ;
        RECT 58.750 32.730 58.920 32.900 ;
        RECT 63.440 33.480 63.610 33.650 ;
        RECT 63.440 33.140 63.610 33.310 ;
        RECT 66.500 32.880 66.670 33.050 ;
        RECT 68.310 33.170 68.480 33.340 ;
        RECT 67.230 32.910 67.400 33.080 ;
        RECT 79.800 33.010 79.970 33.180 ;
        RECT 81.950 33.130 82.120 33.300 ;
        RECT 68.310 32.620 68.480 32.790 ;
        RECT 80.690 32.560 80.860 32.730 ;
        RECT 40.590 31.740 40.800 31.950 ;
        RECT 46.510 32.020 46.680 32.190 ;
        RECT 18.050 31.570 18.220 31.740 ;
        RECT 45.470 31.670 45.640 31.840 ;
        RECT 79.800 32.110 79.970 32.280 ;
        RECT 58.750 31.840 58.920 32.010 ;
        RECT 63.040 31.540 63.210 31.710 ;
        RECT 15.520 30.090 15.690 30.260 ;
        RECT 17.860 30.610 18.030 30.780 ;
        RECT 39.120 30.600 39.290 30.770 ;
        RECT 59.310 31.210 59.480 31.380 ;
        RECT 60.060 31.210 60.230 31.380 ;
        RECT 62.060 31.220 62.230 31.390 ;
        RECT 63.440 31.770 63.610 31.940 ;
        RECT 81.950 31.990 82.120 32.160 ;
        RECT 63.440 31.430 63.610 31.600 ;
        RECT 79.650 31.430 79.820 31.600 ;
        RECT 46.510 30.820 46.680 30.990 ;
        RECT 79.650 30.920 79.820 31.090 ;
        RECT 16.210 30.080 16.380 30.250 ;
        RECT 40.590 30.190 40.800 30.400 ;
        RECT 46.510 30.470 46.680 30.640 ;
        RECT 58.470 30.550 58.640 30.720 ;
        RECT 45.470 30.120 45.640 30.290 ;
        RECT 59.310 30.430 59.480 30.600 ;
        RECT 60.060 30.430 60.230 30.600 ;
        RECT 16.690 29.310 16.860 29.480 ;
        RECT 17.400 29.250 17.570 29.420 ;
        RECT 39.120 29.050 39.290 29.220 ;
        RECT 63.040 30.100 63.210 30.270 ;
        RECT 58.750 29.800 58.920 29.970 ;
        RECT 63.440 30.550 63.610 30.720 ;
        RECT 63.440 30.210 63.610 30.380 ;
        RECT 79.800 30.240 79.970 30.410 ;
        RECT 81.950 30.360 82.120 30.530 ;
        RECT 80.690 29.790 80.860 29.960 ;
        RECT 46.510 29.270 46.680 29.440 ;
        RECT 40.590 28.640 40.800 28.850 ;
        RECT 46.510 28.920 46.680 29.090 ;
        RECT 68.210 29.280 68.380 29.450 ;
        RECT 79.800 29.340 79.970 29.510 ;
        RECT 17.360 28.430 17.530 28.600 ;
        RECT 45.470 28.570 45.640 28.740 ;
        RECT 58.750 28.910 58.920 29.080 ;
        RECT 63.040 28.610 63.210 28.780 ;
        RECT 14.050 27.990 14.220 28.160 ;
        RECT 15.150 28.000 15.320 28.170 ;
        RECT 14.600 27.320 14.770 27.490 ;
        RECT 14.600 25.950 14.770 26.120 ;
        RECT 14.050 25.220 14.220 25.390 ;
        RECT 14.040 23.880 14.210 24.050 ;
        RECT 16.240 28.000 16.410 28.170 ;
        RECT 15.700 27.320 15.870 27.490 ;
        RECT 15.700 25.950 15.870 26.120 ;
        RECT 15.150 25.220 15.320 25.390 ;
        RECT 15.150 23.870 15.320 24.040 ;
        RECT 14.600 23.180 14.770 23.350 ;
        RECT 59.310 28.280 59.480 28.450 ;
        RECT 60.060 28.280 60.230 28.450 ;
        RECT 62.060 28.290 62.230 28.460 ;
        RECT 63.440 28.840 63.610 29.010 ;
        RECT 63.440 28.500 63.610 28.670 ;
        RECT 81.950 29.220 82.120 29.390 ;
        RECT 79.650 28.660 79.820 28.830 ;
        RECT 68.260 28.430 68.430 28.600 ;
        RECT 17.370 27.960 17.540 28.130 ;
        RECT 16.800 27.320 16.970 27.490 ;
        RECT 39.120 27.500 39.290 27.670 ;
        RECT 17.490 27.300 17.660 27.470 ;
        RECT 46.510 27.720 46.680 27.890 ;
        RECT 17.490 26.960 17.660 27.130 ;
        RECT 40.590 27.090 40.800 27.300 ;
        RECT 46.510 27.370 46.680 27.540 ;
        RECT 45.470 27.020 45.640 27.190 ;
        RECT 17.490 26.620 17.660 26.790 ;
        RECT 16.800 25.950 16.970 26.120 ;
        RECT 16.240 25.220 16.410 25.390 ;
        RECT 16.240 23.850 16.410 24.020 ;
        RECT 15.700 23.170 15.870 23.340 ;
        RECT 24.070 24.050 24.240 24.390 ;
        RECT 24.410 24.050 24.580 24.390 ;
        RECT 16.790 23.170 16.960 23.340 ;
        RECT 16.650 20.870 16.820 21.040 ;
        RECT 13.340 20.430 13.510 20.600 ;
        RECT 14.440 20.440 14.610 20.610 ;
        RECT 15.530 20.440 15.700 20.610 ;
        RECT 13.890 19.760 14.060 19.930 ;
        RECT 14.990 19.760 15.160 19.930 ;
        RECT 13.890 18.390 14.060 18.560 ;
        RECT 14.990 18.390 15.160 18.560 ;
        RECT 16.660 20.400 16.830 20.570 ;
        RECT 16.090 19.760 16.260 19.930 ;
        RECT 16.090 18.390 16.260 18.560 ;
        RECT 47.750 21.710 47.920 21.880 ;
        RECT 48.840 21.710 49.010 21.880 ;
        RECT 48.300 21.030 48.470 21.200 ;
        RECT 48.300 19.660 48.470 19.830 ;
        RECT 51.060 21.880 51.230 22.050 ;
        RECT 49.940 21.700 50.110 21.870 ;
        RECT 51.060 21.540 51.230 21.710 ;
        RECT 51.450 21.880 51.620 22.050 ;
        RECT 51.450 21.540 51.620 21.710 ;
        RECT 52.570 21.700 52.740 21.870 ;
        RECT 53.670 21.710 53.840 21.880 ;
        RECT 49.390 21.010 49.560 21.180 ;
        RECT 50.500 21.000 50.670 21.170 ;
        RECT 52.010 21.000 52.180 21.170 ;
        RECT 53.120 21.010 53.290 21.180 ;
        RECT 49.390 19.660 49.560 19.830 ;
        RECT 50.490 19.660 50.660 19.830 ;
        RECT 52.020 19.660 52.190 19.830 ;
        RECT 53.120 19.660 53.290 19.830 ;
        RECT 54.760 21.710 54.930 21.880 ;
        RECT 54.210 21.030 54.380 21.200 ;
        RECT 54.210 19.660 54.380 19.830 ;
        RECT 57.560 21.740 57.730 21.910 ;
        RECT 58.650 21.740 58.820 21.910 ;
        RECT 58.110 21.060 58.280 21.230 ;
        RECT 58.110 19.690 58.280 19.860 ;
        RECT 60.870 21.910 61.040 22.080 ;
        RECT 59.750 21.730 59.920 21.900 ;
        RECT 60.870 21.570 61.040 21.740 ;
        RECT 61.260 21.910 61.430 22.080 ;
        RECT 61.260 21.570 61.430 21.740 ;
        RECT 62.380 21.730 62.550 21.900 ;
        RECT 63.480 21.740 63.650 21.910 ;
        RECT 59.200 21.040 59.370 21.210 ;
        RECT 60.310 21.030 60.480 21.200 ;
        RECT 61.820 21.030 61.990 21.200 ;
        RECT 62.930 21.040 63.100 21.210 ;
        RECT 59.200 19.690 59.370 19.860 ;
        RECT 60.300 19.690 60.470 19.860 ;
        RECT 61.830 19.690 62.000 19.860 ;
        RECT 62.930 19.690 63.100 19.860 ;
        RECT 64.570 21.740 64.740 21.910 ;
        RECT 64.020 21.060 64.190 21.230 ;
        RECT 64.020 19.690 64.190 19.860 ;
        RECT 68.870 21.710 69.040 21.880 ;
        RECT 68.310 21.010 68.480 21.180 ;
        RECT 68.320 19.670 68.490 19.840 ;
        RECT 13.340 17.660 13.510 17.830 ;
        RECT 14.440 17.660 14.610 17.830 ;
        RECT 13.330 16.320 13.500 16.490 ;
        RECT 14.440 16.310 14.610 16.480 ;
        RECT 12.770 15.780 12.940 15.950 ;
        RECT 13.890 15.620 14.060 15.790 ;
        RECT 15.530 17.660 15.700 17.830 ;
        RECT 15.530 16.290 15.700 16.460 ;
        RECT 14.990 15.610 15.160 15.780 ;
        RECT 16.080 15.610 16.250 15.780 ;
        RECT 47.740 18.930 47.910 19.100 ;
        RECT 47.740 17.560 47.910 17.730 ;
        RECT 47.170 16.920 47.340 17.090 ;
        RECT 48.840 18.930 49.010 19.100 ;
        RECT 49.940 18.930 50.110 19.100 ;
        RECT 52.570 18.930 52.740 19.100 ;
        RECT 53.670 18.930 53.840 19.100 ;
        RECT 48.840 17.560 49.010 17.730 ;
        RECT 49.940 17.560 50.110 17.730 ;
        RECT 52.570 17.560 52.740 17.730 ;
        RECT 53.670 17.560 53.840 17.730 ;
        RECT 48.300 16.880 48.470 17.050 ;
        RECT 49.390 16.880 49.560 17.050 ;
        RECT 50.490 16.890 50.660 17.060 ;
        RECT 52.020 16.890 52.190 17.060 ;
        RECT 53.120 16.880 53.290 17.050 ;
        RECT 54.770 18.930 54.940 19.100 ;
        RECT 54.770 17.560 54.940 17.730 ;
        RECT 54.210 16.880 54.380 17.050 ;
        RECT 55.340 16.920 55.510 17.090 ;
        RECT 57.550 18.960 57.720 19.130 ;
        RECT 57.550 17.590 57.720 17.760 ;
        RECT 56.980 16.950 57.150 17.120 ;
        RECT 58.650 18.960 58.820 19.130 ;
        RECT 59.750 18.960 59.920 19.130 ;
        RECT 62.380 18.960 62.550 19.130 ;
        RECT 63.480 18.960 63.650 19.130 ;
        RECT 58.650 17.590 58.820 17.760 ;
        RECT 59.750 17.590 59.920 17.760 ;
        RECT 62.380 17.590 62.550 17.760 ;
        RECT 63.480 17.590 63.650 17.760 ;
        RECT 47.180 16.450 47.350 16.620 ;
        RECT 55.330 16.450 55.500 16.620 ;
        RECT 58.110 16.910 58.280 17.080 ;
        RECT 59.200 16.910 59.370 17.080 ;
        RECT 60.300 16.920 60.470 17.090 ;
        RECT 61.830 16.920 62.000 17.090 ;
        RECT 62.930 16.910 63.100 17.080 ;
        RECT 64.580 18.960 64.750 19.130 ;
        RECT 64.580 17.590 64.750 17.760 ;
        RECT 64.020 16.910 64.190 17.080 ;
        RECT 65.150 16.950 65.320 17.120 ;
        RECT 69.970 21.720 70.140 21.890 ;
        RECT 69.420 21.020 69.590 21.190 ;
        RECT 69.420 19.670 69.590 19.840 ;
        RECT 68.870 18.940 69.040 19.110 ;
        RECT 68.870 17.570 69.040 17.740 ;
        RECT 56.990 16.480 57.160 16.650 ;
        RECT 68.320 16.900 68.490 17.070 ;
        RECT 71.060 21.720 71.230 21.890 ;
        RECT 70.510 21.040 70.680 21.210 ;
        RECT 70.510 19.670 70.680 19.840 ;
        RECT 69.970 18.940 70.140 19.110 ;
        RECT 69.970 17.570 70.140 17.740 ;
        RECT 69.420 16.890 69.590 17.060 ;
        RECT 71.070 18.940 71.240 19.110 ;
        RECT 71.760 18.610 71.930 18.780 ;
        RECT 71.760 18.270 71.930 18.440 ;
        RECT 71.760 17.930 71.930 18.100 ;
        RECT 71.070 17.570 71.240 17.740 ;
        RECT 70.510 16.890 70.680 17.060 ;
        RECT 71.640 16.930 71.810 17.100 ;
        RECT 65.140 16.480 65.310 16.650 ;
        RECT 71.630 16.460 71.800 16.630 ;
        RECT 18.230 12.080 18.400 15.600 ;
        RECT 18.600 12.080 18.770 15.600 ;
        RECT 18.950 12.080 19.120 15.600 ;
        RECT 19.290 12.080 19.460 15.600 ;
        RECT 19.640 12.080 19.810 15.600 ;
        RECT 20.000 12.080 20.170 15.600 ;
        RECT 20.360 12.080 20.530 15.600 ;
        RECT 97.000 14.310 97.170 14.480 ;
        RECT 102.520 13.570 102.690 13.740 ;
        RECT 97.000 12.700 97.170 12.870 ;
        RECT 102.520 12.900 102.690 13.070 ;
        RECT 97.000 11.100 97.170 11.270 ;
        RECT 97.000 9.480 97.170 9.650 ;
        RECT 99.530 8.270 99.700 8.440 ;
        RECT 97.000 7.880 97.170 8.050 ;
        RECT 97.000 6.260 97.170 6.430 ;
        RECT 97.000 4.660 97.170 4.830 ;
        RECT 108.600 4.870 108.770 19.820 ;
        RECT 97.000 3.040 97.170 3.210 ;
      LAYER met1 ;
        RECT 80.150 76.420 80.490 76.560 ;
        RECT 88.030 76.420 88.750 78.160 ;
        RECT 80.150 75.700 88.750 76.420 ;
        RECT 28.080 73.250 29.420 73.700 ;
        RECT 1.980 72.410 2.480 72.890 ;
        RECT 28.080 72.830 41.600 73.250 ;
        RECT 43.390 73.160 46.580 74.280 ;
        RECT 28.080 72.690 29.420 72.830 ;
        RECT 2.080 69.450 2.470 72.410 ;
        RECT 22.670 72.090 25.440 72.330 ;
        RECT 4.450 71.630 4.710 71.830 ;
        RECT 7.310 71.790 7.570 71.880 ;
        RECT 4.390 71.320 4.770 71.630 ;
        RECT 5.800 71.320 6.830 71.630 ;
        RECT 7.300 71.560 7.590 71.790 ;
        RECT 4.440 70.530 4.700 70.800 ;
        RECT 5.130 70.530 5.450 70.770 ;
        RECT 5.850 70.530 6.110 70.810 ;
        RECT 4.400 69.870 6.150 70.530 ;
        RECT 4.440 69.610 4.700 69.870 ;
        RECT 5.130 69.610 5.450 69.870 ;
        RECT 5.870 69.630 6.130 69.870 ;
        RECT 2.080 68.960 2.550 69.450 ;
        RECT 2.080 68.950 2.530 68.960 ;
        RECT 2.080 10.840 2.470 68.950 ;
        RECT 4.460 68.580 4.690 69.100 ;
        RECT 4.440 68.260 4.700 68.580 ;
        RECT 3.490 67.810 3.750 68.130 ;
        RECT 3.500 65.590 3.740 67.810 ;
        RECT 4.460 67.690 4.690 68.260 ;
        RECT 5.870 67.690 6.100 69.100 ;
        RECT 6.590 68.550 6.830 71.320 ;
        RECT 22.670 71.000 22.910 72.090 ;
        RECT 7.250 70.870 7.640 71.000 ;
        RECT 7.250 70.580 7.670 70.870 ;
        RECT 22.670 70.740 22.900 71.000 ;
        RECT 6.970 70.020 7.290 70.340 ;
        RECT 7.020 69.790 7.250 70.020 ;
        RECT 7.440 69.640 7.670 70.580 ;
        RECT 22.660 70.520 22.900 70.740 ;
        RECT 20.520 69.710 20.840 70.030 ;
        RECT 21.880 69.790 22.200 70.110 ;
        RECT 22.570 69.780 22.890 70.100 ;
        RECT 7.310 69.570 7.670 69.640 ;
        RECT 7.250 69.460 7.670 69.570 ;
        RECT 7.250 69.340 7.640 69.460 ;
        RECT 6.550 68.010 6.870 68.330 ;
        RECT 7.310 68.170 7.580 69.340 ;
        RECT 22.670 68.200 22.910 68.840 ;
        RECT 7.310 67.940 7.640 68.170 ;
        RECT 22.670 67.940 22.900 68.200 ;
        RECT 22.660 67.290 22.900 67.940 ;
        RECT 5.110 66.810 5.430 67.130 ;
        RECT 6.540 66.830 6.860 67.150 ;
        RECT 4.320 66.230 4.640 66.550 ;
        RECT 5.250 66.230 5.570 66.550 ;
        RECT 5.950 66.230 6.270 66.550 ;
        RECT 6.690 66.230 7.010 66.550 ;
        RECT 7.400 66.220 7.720 66.540 ;
        RECT 3.410 65.110 3.830 65.590 ;
        RECT 9.300 64.350 9.590 67.040 ;
        RECT 22.660 66.650 22.910 67.290 ;
        RECT 19.800 66.050 20.120 66.370 ;
        RECT 9.280 63.680 9.690 64.350 ;
        RECT 22.660 62.990 22.900 66.650 ;
        RECT 22.610 62.650 22.950 62.990 ;
        RECT 19.860 62.550 20.350 62.560 ;
        RECT 15.800 58.310 16.120 58.630 ;
        RECT 16.890 58.320 17.210 58.640 ;
        RECT 15.330 58.170 15.650 58.220 ;
        RECT 15.330 57.940 15.880 58.170 ;
        RECT 15.330 57.900 15.650 57.940 ;
        RECT 15.800 57.390 16.120 57.710 ;
        RECT 16.890 57.400 17.210 57.720 ;
        RECT 15.330 57.250 15.650 57.300 ;
        RECT 15.330 57.020 15.880 57.250 ;
        RECT 15.330 56.980 15.650 57.020 ;
        RECT 15.930 56.790 16.160 57.340 ;
        RECT 15.800 56.470 16.160 56.790 ;
        RECT 16.600 56.720 16.820 57.340 ;
        RECT 15.330 56.330 15.650 56.380 ;
        RECT 15.330 56.100 15.880 56.330 ;
        RECT 15.330 56.060 15.650 56.100 ;
        RECT 15.930 55.810 16.160 56.470 ;
        RECT 16.570 56.400 16.830 56.720 ;
        RECT 16.890 56.480 17.210 56.800 ;
        RECT 15.610 55.490 16.160 55.810 ;
        RECT 16.600 55.800 16.820 56.400 ;
        RECT 15.930 55.350 16.160 55.490 ;
        RECT 16.540 55.480 16.820 55.800 ;
        RECT 15.610 55.310 16.160 55.350 ;
        RECT 15.380 55.080 16.160 55.310 ;
        RECT 15.610 55.030 16.160 55.080 ;
        RECT 15.930 54.850 16.160 55.030 ;
        RECT 16.600 54.880 16.820 55.480 ;
        RECT 16.910 55.390 17.230 55.710 ;
        RECT 15.610 54.530 16.160 54.850 ;
        RECT 16.550 54.560 16.820 54.880 ;
        RECT 15.930 54.390 16.160 54.530 ;
        RECT 15.610 54.350 16.160 54.390 ;
        RECT 15.380 54.120 16.160 54.350 ;
        RECT 15.610 54.070 16.160 54.120 ;
        RECT 15.930 53.890 16.160 54.070 ;
        RECT 15.610 53.570 16.160 53.890 ;
        RECT 15.900 53.540 16.160 53.570 ;
        RECT 15.930 53.430 16.160 53.540 ;
        RECT 15.610 53.390 16.160 53.430 ;
        RECT 15.380 53.160 16.160 53.390 ;
        RECT 15.610 53.110 16.160 53.160 ;
        RECT 15.930 52.900 16.160 53.110 ;
        RECT 15.860 52.580 16.160 52.900 ;
        RECT 15.930 51.940 16.160 52.580 ;
        RECT 15.900 51.620 16.160 51.940 ;
        RECT 15.930 36.870 16.160 51.620 ;
        RECT 16.600 36.870 16.820 54.560 ;
        RECT 16.910 54.430 17.230 54.750 ;
        RECT 16.910 53.470 17.230 53.790 ;
        RECT 17.380 53.300 17.600 58.780 ;
        RECT 17.780 58.150 18.000 58.780 ;
        RECT 17.770 57.860 18.000 58.150 ;
        RECT 17.320 53.070 17.610 53.300 ;
        RECT 17.380 52.900 17.600 53.070 ;
        RECT 17.780 52.900 18.000 57.860 ;
        RECT 19.290 57.060 19.510 61.610 ;
        RECT 19.850 61.400 20.360 62.550 ;
        RECT 25.200 61.620 25.440 72.090 ;
        RECT 28.510 71.760 31.540 72.030 ;
        RECT 28.510 70.780 28.780 71.760 ;
        RECT 28.520 68.570 28.780 68.590 ;
        RECT 28.480 62.590 28.790 68.570 ;
        RECT 29.660 66.070 29.980 66.390 ;
        RECT 28.400 62.220 28.790 62.590 ;
        RECT 31.270 62.080 31.540 71.760 ;
        RECT 33.220 70.740 33.480 72.830 ;
        RECT 41.180 69.580 41.600 72.830 ;
        RECT 44.990 70.340 45.410 73.160 ;
        RECT 44.990 69.860 45.460 70.340 ;
        RECT 41.140 69.100 41.620 69.580 ;
        RECT 32.450 68.030 32.680 68.200 ;
        RECT 32.440 66.160 32.690 68.030 ;
        RECT 46.690 67.490 47.130 67.990 ;
        RECT 52.410 67.490 52.850 67.990 ;
        RECT 42.270 66.470 42.710 66.970 ;
        RECT 32.440 65.980 32.700 66.160 ;
        RECT 32.440 63.080 32.690 65.980 ;
        RECT 39.480 63.730 39.800 63.780 ;
        RECT 39.390 63.440 39.800 63.730 ;
        RECT 32.400 62.720 32.730 63.080 ;
        RECT 31.230 61.770 31.570 62.080 ;
        RECT 19.800 61.300 20.360 61.400 ;
        RECT 25.150 61.300 25.490 61.620 ;
        RECT 38.900 61.550 39.140 61.600 ;
        RECT 19.690 60.900 20.360 61.300 ;
        RECT 19.690 60.870 20.350 60.900 ;
        RECT 19.690 57.060 19.910 60.870 ;
        RECT 38.350 59.700 38.760 60.030 ;
        RECT 20.910 58.750 21.260 59.210 ;
        RECT 37.340 58.770 37.710 59.080 ;
        RECT 20.310 58.390 20.560 58.510 ;
        RECT 20.280 57.930 20.600 58.390 ;
        RECT 20.310 57.140 20.560 57.930 ;
        RECT 20.310 56.820 20.600 57.140 ;
        RECT 20.310 56.220 20.560 56.820 ;
        RECT 20.310 55.900 20.600 56.220 ;
        RECT 20.310 55.300 20.560 55.900 ;
        RECT 20.310 54.980 20.570 55.300 ;
        RECT 15.820 36.340 16.160 36.870 ;
        RECT 16.480 36.340 16.820 36.870 ;
        RECT 14.510 35.600 14.740 35.670 ;
        RECT 14.470 35.340 14.790 35.600 ;
        RECT 14.020 35.230 14.250 35.270 ;
        RECT 13.980 34.910 14.250 35.230 ;
        RECT 4.670 33.670 5.390 34.370 ;
        RECT 4.680 28.520 5.340 33.670 ;
        RECT 14.020 31.390 14.250 34.910 ;
        RECT 14.510 32.870 14.740 35.340 ;
        RECT 15.930 35.250 16.160 36.340 ;
        RECT 16.600 35.610 16.820 36.340 ;
        RECT 18.360 35.630 18.630 35.670 ;
        RECT 16.580 35.290 16.840 35.610 ;
        RECT 18.340 35.300 18.630 35.630 ;
        RECT 15.920 34.930 16.180 35.250 ;
        RECT 16.640 34.330 16.960 34.650 ;
        RECT 17.290 34.330 17.610 34.650 ;
        RECT 15.420 33.890 15.740 34.210 ;
        RECT 16.120 33.890 16.440 34.210 ;
        RECT 17.810 32.880 18.100 33.790 ;
        RECT 14.510 32.860 15.240 32.870 ;
        RECT 14.510 32.540 15.260 32.860 ;
        RECT 14.510 32.500 15.240 32.540 ;
        RECT 14.020 31.320 14.280 31.390 ;
        RECT 14.000 31.310 14.280 31.320 ;
        RECT 13.970 31.000 14.290 31.310 ;
        RECT 9.870 29.140 10.300 29.570 ;
        RECT 4.680 27.800 5.420 28.520 ;
        RECT 9.920 23.330 10.290 29.140 ;
        RECT 13.970 27.910 14.290 28.230 ;
        RECT 14.510 27.560 14.740 32.500 ;
        RECT 15.010 32.250 15.240 32.500 ;
        RECT 17.720 32.310 18.040 32.350 ;
        RECT 18.360 32.330 18.630 35.300 ;
        RECT 18.240 32.310 18.630 32.330 ;
        RECT 15.010 32.030 15.230 32.250 ;
        RECT 17.720 32.080 18.630 32.310 ;
        RECT 18.840 35.230 19.080 35.270 ;
        RECT 18.840 34.910 19.100 35.230 ;
        RECT 17.720 32.030 18.040 32.080 ;
        RECT 15.030 31.600 15.250 31.820 ;
        RECT 15.020 31.310 15.250 31.600 ;
        RECT 17.730 31.770 18.050 31.810 ;
        RECT 18.840 31.770 19.080 34.910 ;
        RECT 17.730 31.540 19.080 31.770 ;
        RECT 17.730 31.490 18.050 31.540 ;
        RECT 15.000 30.990 15.260 31.310 ;
        RECT 17.800 30.860 18.070 31.040 ;
        RECT 17.780 30.540 18.100 30.860 ;
        RECT 17.800 30.370 18.070 30.540 ;
        RECT 15.450 30.010 15.770 30.330 ;
        RECT 16.140 30.000 16.460 30.320 ;
        RECT 16.620 29.230 16.940 29.550 ;
        RECT 17.330 29.170 17.650 29.490 ;
        RECT 17.280 28.350 17.600 28.670 ;
        RECT 15.070 27.920 15.390 28.240 ;
        RECT 16.160 27.920 16.480 28.240 ;
        RECT 17.290 27.880 17.610 28.200 ;
        RECT 14.510 27.240 14.840 27.560 ;
        RECT 15.620 27.240 15.940 27.560 ;
        RECT 16.720 27.240 17.040 27.560 ;
        RECT 14.510 26.190 14.740 27.240 ;
        RECT 17.430 27.070 17.720 27.500 ;
        RECT 17.430 27.050 17.900 27.070 ;
        RECT 17.440 26.750 17.900 27.050 ;
        RECT 17.440 26.220 17.720 26.750 ;
        RECT 14.510 25.870 14.840 26.190 ;
        RECT 15.620 25.870 15.940 26.190 ;
        RECT 16.720 25.870 17.040 26.190 ;
        RECT 13.970 25.140 14.290 25.460 ;
        RECT 14.510 25.000 14.740 25.870 ;
        RECT 15.070 25.140 15.390 25.460 ;
        RECT 16.160 25.140 16.480 25.460 ;
        RECT 14.510 24.770 16.960 25.000 ;
        RECT 16.640 24.440 16.960 24.770 ;
        RECT 13.960 23.800 14.280 24.120 ;
        RECT 15.070 23.790 15.390 24.110 ;
        RECT 16.160 23.770 16.480 24.090 ;
        RECT 9.880 22.900 10.310 23.330 ;
        RECT 14.520 23.100 14.840 23.420 ;
        RECT 15.620 23.090 15.940 23.410 ;
        RECT 16.710 23.090 17.030 23.410 ;
        RECT 17.400 22.870 17.730 22.900 ;
        RECT 17.260 22.790 17.730 22.870 ;
        RECT 17.020 22.550 17.730 22.790 ;
        RECT 17.400 22.480 17.730 22.550 ;
        RECT 12.790 17.590 13.050 21.120 ;
        RECT 16.570 20.790 16.890 21.110 ;
        RECT 13.260 20.350 13.580 20.670 ;
        RECT 14.360 20.360 14.680 20.680 ;
        RECT 15.450 20.360 15.770 20.680 ;
        RECT 16.580 20.320 16.900 20.640 ;
        RECT 13.810 19.680 14.130 20.000 ;
        RECT 14.910 19.680 15.230 20.000 ;
        RECT 16.010 19.680 16.330 20.000 ;
        RECT 13.810 18.310 14.130 18.630 ;
        RECT 14.910 18.310 15.230 18.630 ;
        RECT 16.010 18.310 16.330 18.630 ;
        RECT 12.790 17.240 13.180 17.590 ;
        RECT 13.260 17.580 13.580 17.900 ;
        RECT 14.360 17.580 14.680 17.900 ;
        RECT 15.450 17.580 15.770 17.900 ;
        RECT 12.790 16.670 13.160 17.240 ;
        RECT 18.840 16.880 19.080 31.540 ;
        RECT 19.290 30.870 19.510 51.620 ;
        RECT 19.690 33.480 19.910 51.620 ;
        RECT 20.310 34.630 20.560 54.980 ;
        RECT 20.930 54.210 21.190 58.750 ;
        RECT 36.700 57.050 37.090 57.420 ;
        RECT 36.120 55.560 36.510 55.950 ;
        RECT 20.930 53.890 21.210 54.210 ;
        RECT 35.480 53.970 35.870 54.350 ;
        RECT 35.510 53.960 35.850 53.970 ;
        RECT 20.930 53.250 21.190 53.890 ;
        RECT 34.870 53.770 35.210 53.780 ;
        RECT 34.860 53.380 35.220 53.770 ;
        RECT 20.930 52.930 21.220 53.250 ;
        RECT 20.930 52.290 21.190 52.930 ;
        RECT 20.930 51.970 21.210 52.290 ;
        RECT 20.310 34.610 20.570 34.630 ;
        RECT 20.300 34.330 20.580 34.610 ;
        RECT 20.310 34.310 20.570 34.330 ;
        RECT 19.650 33.160 19.970 33.480 ;
        RECT 19.250 30.550 19.530 30.870 ;
        RECT 19.290 17.580 19.510 30.550 ;
        RECT 19.690 25.340 19.910 33.160 ;
        RECT 19.690 24.860 19.980 25.340 ;
        RECT 19.690 22.900 19.910 24.860 ;
        RECT 19.670 22.480 19.930 22.900 ;
        RECT 19.690 17.860 19.910 22.480 ;
        RECT 20.310 19.240 20.560 34.310 ;
        RECT 20.930 30.300 21.190 51.970 ;
        RECT 34.250 51.820 34.610 52.210 ;
        RECT 33.600 50.280 34.010 50.680 ;
        RECT 33.070 48.720 33.430 49.110 ;
        RECT 32.490 43.660 32.820 43.680 ;
        RECT 32.430 43.240 32.820 43.660 ;
        RECT 31.860 42.050 32.190 42.070 ;
        RECT 31.810 41.660 32.200 42.050 ;
        RECT 31.240 40.500 31.570 40.510 ;
        RECT 31.210 40.110 31.570 40.500 ;
        RECT 30.590 38.630 30.980 39.030 ;
        RECT 29.920 33.460 30.350 33.860 ;
        RECT 29.260 31.890 29.670 32.290 ;
        RECT 20.920 29.980 21.230 30.300 ;
        RECT 28.650 30.250 29.040 30.650 ;
        RECT 20.270 18.840 20.570 19.240 ;
        RECT 19.690 17.720 19.930 17.860 ;
        RECT 19.250 17.230 19.560 17.580 ;
        RECT 19.700 17.090 19.930 17.720 ;
        RECT 12.790 16.140 13.050 16.670 ;
        RECT 13.250 16.240 13.570 16.560 ;
        RECT 14.360 16.230 14.680 16.550 ;
        RECT 15.450 16.210 15.770 16.530 ;
        RECT 18.050 16.320 19.080 16.880 ;
        RECT 19.690 17.060 19.930 17.090 ;
        RECT 18.050 16.210 18.840 16.320 ;
        RECT 12.740 15.330 13.050 16.140 ;
        RECT 13.810 15.540 14.130 15.860 ;
        RECT 14.910 15.530 15.230 15.850 ;
        RECT 16.000 15.530 16.320 15.850 ;
        RECT 19.690 15.670 19.910 17.060 ;
        RECT 12.790 15.130 13.050 15.330 ;
        RECT 18.160 11.990 20.580 15.670 ;
        RECT 20.930 11.700 21.190 29.980 ;
        RECT 27.960 28.810 28.370 29.200 ;
        RECT 23.750 23.660 24.680 25.310 ;
        RECT 23.840 23.180 24.580 23.660 ;
        RECT 20.840 11.290 21.190 11.700 ;
        RECT 1.910 10.320 2.470 10.840 ;
        RECT 28.020 5.470 28.350 28.810 ;
        RECT 27.970 5.460 28.400 5.470 ;
        RECT 27.940 5.000 28.430 5.460 ;
        RECT 27.970 4.980 28.400 5.000 ;
        RECT 28.670 4.680 29.000 30.250 ;
        RECT 28.580 4.190 29.070 4.680 ;
        RECT 29.320 3.970 29.650 31.890 ;
        RECT 29.290 3.510 29.690 3.970 ;
        RECT 29.080 3.020 29.660 3.130 ;
        RECT 29.990 3.020 30.320 33.460 ;
        RECT 30.630 7.600 30.960 38.630 ;
        RECT 30.630 3.140 30.950 7.600 ;
        RECT 31.240 3.750 31.570 40.110 ;
        RECT 31.860 4.000 32.190 41.660 ;
        RECT 32.490 5.030 32.820 43.240 ;
        RECT 33.090 5.330 33.420 48.720 ;
        RECT 33.670 5.900 34.000 50.280 ;
        RECT 34.280 6.930 34.610 51.820 ;
        RECT 34.870 7.540 35.200 53.380 ;
        RECT 35.510 8.210 35.840 53.960 ;
        RECT 36.130 8.860 36.460 55.560 ;
        RECT 36.730 9.490 37.060 57.050 ;
        RECT 37.360 10.100 37.690 58.770 ;
        RECT 38.350 58.150 38.760 58.480 ;
        RECT 38.350 56.600 38.760 56.930 ;
        RECT 39.090 55.410 39.330 61.200 ;
        RECT 39.390 59.940 39.630 63.440 ;
        RECT 41.840 61.530 42.150 61.600 ;
        RECT 42.330 61.200 42.640 66.470 ;
        RECT 46.270 61.550 46.560 61.600 ;
        RECT 40.510 60.560 40.860 60.850 ;
        RECT 40.510 60.540 40.710 60.560 ;
        RECT 42.030 60.140 42.640 61.200 ;
        RECT 45.390 60.660 45.710 60.960 ;
        RECT 42.030 59.870 42.870 60.140 ;
        RECT 40.510 59.010 40.860 59.300 ;
        RECT 40.510 58.990 40.710 59.010 ;
        RECT 40.510 57.460 40.860 57.750 ;
        RECT 40.510 57.440 40.710 57.460 ;
        RECT 40.510 55.910 40.860 56.200 ;
        RECT 40.510 55.890 40.710 55.910 ;
        RECT 42.030 55.420 42.340 59.870 ;
        RECT 42.590 59.810 42.870 59.870 ;
        RECT 45.390 59.110 45.710 59.410 ;
        RECT 42.590 58.260 42.870 58.590 ;
        RECT 45.390 57.560 45.710 57.860 ;
        RECT 42.590 56.710 42.870 57.040 ;
        RECT 45.390 56.010 45.710 56.310 ;
        RECT 38.350 55.050 38.760 55.380 ;
        RECT 38.900 55.360 39.330 55.410 ;
        RECT 41.840 55.360 42.340 55.420 ;
        RECT 39.090 54.960 39.330 55.360 ;
        RECT 42.030 54.960 42.340 55.360 ;
        RECT 42.590 55.160 42.870 55.490 ;
        RECT 46.460 55.410 46.750 61.200 ;
        RECT 46.760 59.890 47.050 67.490 ;
        RECT 47.950 66.500 48.450 66.940 ;
        RECT 46.270 55.360 46.750 55.410 ;
        RECT 46.460 54.960 46.750 55.360 ;
        RECT 42.630 53.940 42.640 53.950 ;
        RECT 39.390 53.860 39.630 53.940 ;
        RECT 42.330 53.860 42.640 53.940 ;
        RECT 46.760 53.860 47.050 53.940 ;
        RECT 48.220 53.500 48.410 66.500 ;
        RECT 52.500 53.460 52.750 67.490 ;
        RECT 54.200 67.450 54.930 74.320 ;
        RECT 71.980 73.150 75.170 74.270 ;
        RECT 64.750 69.080 66.220 69.610 ;
        RECT 54.360 57.060 54.530 67.450 ;
        RECT 62.380 66.470 62.820 66.970 ;
        RECT 56.580 62.720 56.920 63.010 ;
        RECT 56.630 62.690 56.890 62.720 ;
        RECT 54.750 59.160 55.010 59.480 ;
        RECT 54.780 56.930 54.970 59.160 ;
        RECT 56.650 56.910 56.860 62.690 ;
        RECT 60.220 62.090 60.480 62.100 ;
        RECT 60.200 61.790 60.500 62.090 ;
        RECT 60.220 61.780 60.480 61.790 ;
        RECT 57.050 60.760 57.390 61.080 ;
        RECT 57.120 56.930 57.310 60.760 ;
        RECT 57.490 58.670 57.780 58.990 ;
        RECT 57.530 56.910 57.740 58.670 ;
        RECT 58.530 58.190 58.870 58.510 ;
        RECT 58.610 56.940 58.790 58.190 ;
        RECT 60.250 53.760 60.450 61.780 ;
        RECT 62.480 56.890 62.710 66.470 ;
        RECT 63.380 62.700 63.660 63.020 ;
        RECT 62.940 61.790 63.220 62.110 ;
        RECT 58.720 53.540 58.910 53.760 ;
        RECT 58.440 53.050 58.910 53.540 ;
        RECT 59.300 53.400 59.670 53.420 ;
        RECT 59.250 53.140 59.670 53.400 ;
        RECT 59.300 53.130 59.670 53.140 ;
        RECT 38.350 52.420 38.760 52.750 ;
        RECT 39.090 52.440 39.330 52.840 ;
        RECT 42.030 52.440 42.340 52.840 ;
        RECT 38.900 52.390 39.330 52.440 ;
        RECT 38.350 50.870 38.760 51.200 ;
        RECT 38.350 49.320 38.760 49.650 ;
        RECT 38.350 47.770 38.760 48.100 ;
        RECT 39.090 46.600 39.330 52.390 ;
        RECT 41.840 52.380 42.340 52.440 ;
        RECT 40.510 51.890 40.710 51.910 ;
        RECT 40.510 51.600 40.860 51.890 ;
        RECT 40.510 50.340 40.710 50.360 ;
        RECT 40.510 50.050 40.860 50.340 ;
        RECT 40.510 48.790 40.710 48.810 ;
        RECT 40.510 48.500 40.860 48.790 ;
        RECT 42.030 47.930 42.340 52.380 ;
        RECT 42.590 52.310 42.870 52.640 ;
        RECT 46.460 52.440 46.750 52.840 ;
        RECT 58.260 52.610 58.580 52.890 ;
        RECT 58.720 52.790 58.910 53.050 ;
        RECT 46.270 52.390 46.750 52.440 ;
        RECT 45.390 51.490 45.710 51.790 ;
        RECT 42.590 50.760 42.870 51.090 ;
        RECT 45.390 49.940 45.710 50.240 ;
        RECT 42.590 49.210 42.870 49.540 ;
        RECT 45.390 48.390 45.710 48.690 ;
        RECT 42.590 47.930 42.870 47.990 ;
        RECT 38.900 46.200 39.140 46.250 ;
        RECT 39.390 43.490 39.630 47.860 ;
        RECT 42.030 47.660 42.870 47.930 ;
        RECT 40.510 47.240 40.710 47.260 ;
        RECT 40.510 46.950 40.860 47.240 ;
        RECT 42.030 46.600 42.640 47.660 ;
        RECT 45.390 46.840 45.710 47.140 ;
        RECT 46.460 46.600 46.750 52.390 ;
        RECT 58.720 52.500 58.950 52.790 ;
        RECT 58.720 51.900 58.910 52.500 ;
        RECT 58.260 51.510 58.580 51.790 ;
        RECT 58.720 51.610 58.950 51.900 ;
        RECT 58.720 51.350 58.910 51.610 ;
        RECT 58.440 50.860 58.910 51.350 ;
        RECT 60.030 51.420 60.450 53.760 ;
        RECT 62.970 53.760 63.190 61.790 ;
        RECT 62.970 53.540 63.250 53.760 ;
        RECT 63.400 53.540 63.630 62.700 ;
        RECT 64.770 56.700 65.190 69.080 ;
        RECT 65.800 56.700 66.220 69.080 ;
        RECT 68.180 66.430 68.620 66.930 ;
        RECT 68.280 59.450 68.510 66.430 ;
        RECT 72.700 61.180 73.980 73.150 ;
        RECT 76.460 67.960 76.740 68.080 ;
        RECT 76.460 67.460 76.790 67.960 ;
        RECT 72.700 61.100 74.000 61.180 ;
        RECT 72.690 60.800 74.000 61.100 ;
        RECT 69.470 60.150 69.770 60.470 ;
        RECT 68.150 59.440 68.510 59.450 ;
        RECT 68.120 58.590 68.510 59.440 ;
        RECT 68.150 58.580 68.510 58.590 ;
        RECT 68.280 56.890 68.510 58.580 ;
        RECT 69.500 56.890 69.730 60.150 ;
        RECT 75.780 59.600 76.210 59.940 ;
        RECT 76.020 56.930 76.210 59.600 ;
        RECT 76.460 56.840 76.740 67.460 ;
        RECT 78.160 62.700 78.420 63.020 ;
        RECT 77.270 61.830 77.530 62.150 ;
        RECT 77.300 58.110 77.490 61.830 ;
        RECT 78.180 58.110 78.400 62.700 ;
        RECT 80.150 59.480 80.490 75.700 ;
        RECT 84.650 72.240 85.020 72.250 ;
        RECT 84.600 71.790 85.100 72.240 ;
        RECT 80.800 63.380 81.120 63.750 ;
        RECT 80.820 59.540 81.090 63.380 ;
        RECT 80.100 59.400 80.490 59.480 ;
        RECT 80.090 58.630 80.490 59.400 ;
        RECT 80.100 58.560 80.490 58.630 ;
        RECT 77.130 57.420 77.810 58.110 ;
        RECT 78.170 57.420 78.850 58.110 ;
        RECT 80.150 56.780 80.490 58.560 ;
        RECT 80.540 58.890 80.700 59.540 ;
        RECT 80.540 58.340 80.810 58.890 ;
        RECT 80.530 58.290 80.810 58.340 ;
        RECT 80.530 58.200 80.700 58.290 ;
        RECT 80.540 54.830 80.700 58.200 ;
        RECT 80.820 58.050 81.140 59.540 ;
        RECT 82.820 59.170 83.030 59.540 ;
        RECT 82.350 58.720 82.660 59.160 ;
        RECT 82.810 58.880 83.040 59.170 ;
        RECT 80.820 58.000 81.160 58.050 ;
        RECT 80.820 57.500 81.500 58.000 ;
        RECT 80.820 56.850 81.110 57.500 ;
        RECT 81.950 57.190 82.270 57.510 ;
        RECT 82.820 57.180 83.030 58.880 ;
        RECT 83.290 58.610 83.480 59.540 ;
        RECT 83.280 58.320 83.510 58.610 ;
        RECT 80.950 55.500 81.110 56.850 ;
        RECT 81.300 56.680 81.540 57.100 ;
        RECT 82.810 56.890 83.040 57.180 ;
        RECT 82.820 56.750 83.030 56.890 ;
        RECT 81.270 56.360 81.540 56.680 ;
        RECT 81.300 55.930 81.540 56.360 ;
        RECT 83.290 56.290 83.480 58.320 ;
        RECT 83.700 56.820 83.910 59.540 ;
        RECT 83.670 56.310 83.910 56.820 ;
        RECT 82.840 56.110 83.030 56.240 ;
        RECT 82.820 55.820 83.050 56.110 ;
        RECT 83.280 56.000 83.510 56.290 ;
        RECT 81.940 55.500 82.260 55.820 ;
        RECT 80.920 55.260 81.150 55.500 ;
        RECT 80.910 55.250 81.150 55.260 ;
        RECT 80.910 54.980 81.160 55.250 ;
        RECT 80.920 54.950 81.140 54.980 ;
        RECT 80.530 54.740 80.700 54.830 ;
        RECT 80.530 54.690 80.810 54.740 ;
        RECT 80.540 54.140 80.810 54.690 ;
        RECT 61.760 53.380 62.100 53.430 ;
        RECT 61.760 53.360 62.320 53.380 ;
        RECT 61.640 53.190 62.320 53.360 ;
        RECT 61.760 53.150 62.320 53.190 ;
        RECT 61.760 53.110 62.100 53.150 ;
        RECT 62.970 52.470 63.640 53.540 ;
        RECT 80.540 53.510 80.700 54.140 ;
        RECT 80.420 52.860 80.700 53.510 ;
        RECT 62.970 51.930 63.250 52.470 ;
        RECT 63.400 51.930 63.630 52.470 ;
        RECT 80.420 52.260 80.810 52.860 ;
        RECT 59.300 51.260 59.670 51.270 ;
        RECT 59.250 51.000 59.670 51.260 ;
        RECT 59.300 50.980 59.670 51.000 ;
        RECT 60.030 51.090 60.510 51.420 ;
        RECT 61.760 51.250 62.100 51.290 ;
        RECT 61.760 51.210 62.320 51.250 ;
        RECT 58.720 50.610 58.910 50.860 ;
        RECT 58.440 50.120 58.910 50.610 ;
        RECT 59.300 50.470 59.670 50.490 ;
        RECT 59.250 50.210 59.670 50.470 ;
        RECT 59.300 50.200 59.670 50.210 ;
        RECT 58.260 49.680 58.580 49.960 ;
        RECT 58.720 49.860 58.910 50.120 ;
        RECT 58.720 49.570 58.950 49.860 ;
        RECT 58.720 48.970 58.910 49.570 ;
        RECT 58.260 48.580 58.580 48.860 ;
        RECT 58.720 48.680 58.950 48.970 ;
        RECT 58.720 48.420 58.910 48.680 ;
        RECT 58.440 47.930 58.910 48.420 ;
        RECT 59.300 48.330 59.670 48.340 ;
        RECT 59.250 48.070 59.670 48.330 ;
        RECT 59.300 48.050 59.670 48.070 ;
        RECT 41.840 46.200 42.150 46.270 ;
        RECT 42.330 43.420 42.640 46.600 ;
        RECT 46.270 46.200 46.560 46.250 ;
        RECT 46.760 43.440 47.050 47.910 ;
        RECT 48.220 43.450 48.410 47.850 ;
        RECT 49.530 43.640 49.760 47.890 ;
        RECT 52.500 43.640 52.750 47.910 ;
        RECT 58.720 47.710 58.910 47.930 ;
        RECT 60.030 47.710 60.260 51.090 ;
        RECT 61.640 51.040 62.320 51.210 ;
        RECT 61.760 51.020 62.320 51.040 ;
        RECT 61.760 50.970 62.100 51.020 ;
        RECT 62.970 50.860 63.640 51.930 ;
        RECT 62.970 50.610 63.250 50.860 ;
        RECT 63.400 50.610 63.630 50.860 ;
        RECT 61.760 50.450 62.100 50.500 ;
        RECT 61.760 50.430 62.320 50.450 ;
        RECT 61.640 50.260 62.320 50.430 ;
        RECT 61.760 50.220 62.320 50.260 ;
        RECT 62.970 50.250 63.640 50.610 ;
        RECT 61.760 50.180 62.100 50.220 ;
        RECT 62.960 50.180 63.640 50.250 ;
        RECT 62.950 49.580 63.640 50.180 ;
        RECT 62.960 49.550 63.640 49.580 ;
        RECT 62.970 49.540 63.640 49.550 ;
        RECT 62.970 49.000 63.250 49.540 ;
        RECT 61.760 48.320 62.100 48.360 ;
        RECT 61.760 48.280 62.320 48.320 ;
        RECT 61.640 48.110 62.320 48.280 ;
        RECT 61.760 48.090 62.320 48.110 ;
        RECT 61.760 48.040 62.100 48.090 ;
        RECT 62.970 47.930 63.640 49.000 ;
        RECT 80.420 48.710 80.700 52.260 ;
        RECT 80.950 52.050 81.140 54.950 ;
        RECT 82.350 53.870 82.660 54.310 ;
        RECT 82.840 54.200 83.030 55.820 ;
        RECT 83.290 54.710 83.480 56.000 ;
        RECT 83.270 54.420 83.500 54.710 ;
        RECT 82.840 53.990 83.070 54.200 ;
        RECT 82.830 53.910 83.070 53.990 ;
        RECT 82.830 53.490 83.060 53.910 ;
        RECT 83.290 53.490 83.480 54.420 ;
        RECT 83.700 53.490 83.910 56.310 ;
        RECT 84.650 55.720 85.020 71.790 ;
        RECT 85.440 68.340 85.900 68.770 ;
        RECT 84.490 55.700 85.090 55.720 ;
        RECT 84.330 55.660 85.090 55.700 ;
        RECT 84.330 55.400 85.020 55.660 ;
        RECT 82.350 52.690 82.660 53.130 ;
        RECT 80.920 52.020 81.140 52.050 ;
        RECT 80.910 51.750 81.160 52.020 ;
        RECT 80.910 51.740 81.150 51.750 ;
        RECT 80.920 51.500 81.150 51.740 ;
        RECT 82.190 51.730 82.510 52.050 ;
        RECT 80.950 49.470 81.110 51.500 ;
        RECT 81.300 50.940 81.540 51.070 ;
        RECT 81.280 50.620 81.540 50.940 ;
        RECT 81.280 50.020 81.540 50.340 ;
        RECT 81.300 49.900 81.540 50.020 ;
        RECT 84.650 49.690 85.020 55.400 ;
        RECT 84.380 49.630 85.100 49.690 ;
        RECT 80.920 49.230 81.150 49.470 ;
        RECT 84.380 49.360 85.020 49.630 ;
        RECT 80.910 49.220 81.150 49.230 ;
        RECT 80.910 48.950 81.160 49.220 ;
        RECT 82.190 48.970 82.510 49.290 ;
        RECT 80.920 48.920 81.140 48.950 ;
        RECT 80.420 48.110 80.810 48.710 ;
        RECT 62.970 47.710 63.250 47.930 ;
        RECT 62.970 46.350 63.190 47.710 ;
        RECT 65.860 46.950 66.020 47.600 ;
        RECT 65.860 46.400 66.130 46.950 ;
        RECT 65.850 46.350 66.130 46.400 ;
        RECT 66.270 46.610 66.460 47.600 ;
        RECT 66.670 46.920 66.830 47.600 ;
        RECT 66.630 46.900 66.830 46.920 ;
        RECT 67.650 46.910 67.970 47.230 ;
        RECT 66.620 46.660 66.850 46.900 ;
        RECT 66.270 46.490 66.440 46.610 ;
        RECT 62.970 46.260 63.320 46.350 ;
        RECT 65.850 46.260 66.020 46.350 ;
        RECT 62.970 46.040 63.480 46.260 ;
        RECT 65.860 45.900 66.020 46.260 ;
        RECT 65.850 45.810 66.020 45.900 ;
        RECT 65.850 45.760 66.130 45.810 ;
        RECT 65.860 45.460 66.130 45.760 ;
        RECT 66.270 45.670 66.430 46.490 ;
        RECT 66.630 46.440 66.830 46.660 ;
        RECT 66.670 45.720 66.830 46.440 ;
        RECT 67.650 46.360 67.970 46.680 ;
        RECT 68.610 46.440 68.850 47.600 ;
        RECT 66.270 45.550 66.440 45.670 ;
        RECT 54.260 44.210 54.540 45.320 ;
        RECT 54.790 44.630 54.980 45.230 ;
        RECT 56.790 44.790 57.180 44.810 ;
        RECT 56.780 44.700 57.180 44.790 ;
        RECT 54.790 44.440 56.420 44.630 ;
        RECT 54.260 43.930 55.980 44.210 ;
        RECT 55.700 43.700 55.980 43.930 ;
        RECT 56.230 43.660 56.420 44.440 ;
        RECT 56.630 44.450 57.180 44.700 ;
        RECT 56.630 44.430 57.170 44.450 ;
        RECT 56.630 43.580 56.790 44.430 ;
        RECT 60.750 44.360 61.130 44.380 ;
        RECT 61.270 44.360 61.500 45.270 ;
        RECT 60.750 44.130 61.500 44.360 ;
        RECT 62.490 44.270 62.720 45.270 ;
        RECT 65.800 44.280 66.220 45.460 ;
        RECT 66.270 44.690 66.460 45.550 ;
        RECT 66.630 45.500 66.830 45.720 ;
        RECT 66.620 45.260 66.850 45.500 ;
        RECT 67.650 45.480 67.970 45.800 ;
        RECT 68.600 45.780 68.870 46.440 ;
        RECT 66.630 45.240 66.830 45.260 ;
        RECT 66.240 44.460 66.480 44.690 ;
        RECT 58.720 43.470 58.910 43.690 ;
        RECT 58.440 42.980 58.910 43.470 ;
        RECT 59.300 43.330 59.670 43.350 ;
        RECT 59.250 43.070 59.670 43.330 ;
        RECT 59.300 43.060 59.670 43.070 ;
        RECT 38.350 42.290 38.760 42.620 ;
        RECT 39.090 42.310 39.330 42.710 ;
        RECT 42.030 42.310 42.340 42.710 ;
        RECT 38.900 42.260 39.330 42.310 ;
        RECT 38.350 40.740 38.760 41.070 ;
        RECT 38.350 39.190 38.760 39.520 ;
        RECT 38.350 37.640 38.760 37.970 ;
        RECT 39.090 36.470 39.330 42.260 ;
        RECT 41.840 42.250 42.340 42.310 ;
        RECT 40.510 41.760 40.710 41.780 ;
        RECT 40.510 41.470 40.860 41.760 ;
        RECT 40.510 40.210 40.710 40.230 ;
        RECT 40.510 39.920 40.860 40.210 ;
        RECT 40.510 38.660 40.710 38.680 ;
        RECT 40.510 38.370 40.860 38.660 ;
        RECT 42.030 37.800 42.340 42.250 ;
        RECT 42.590 42.180 42.870 42.510 ;
        RECT 46.460 42.310 46.750 42.710 ;
        RECT 58.260 42.540 58.580 42.820 ;
        RECT 58.720 42.720 58.910 42.980 ;
        RECT 46.270 42.260 46.750 42.310 ;
        RECT 45.390 41.360 45.710 41.660 ;
        RECT 42.590 40.630 42.870 40.960 ;
        RECT 45.390 39.810 45.710 40.110 ;
        RECT 42.590 39.080 42.870 39.410 ;
        RECT 45.390 38.260 45.710 38.560 ;
        RECT 42.590 37.800 42.870 37.860 ;
        RECT 38.900 36.070 39.140 36.120 ;
        RECT 39.390 33.960 39.630 37.730 ;
        RECT 42.030 37.530 42.870 37.800 ;
        RECT 40.510 37.110 40.710 37.130 ;
        RECT 40.510 36.820 40.860 37.110 ;
        RECT 42.030 36.470 42.640 37.530 ;
        RECT 45.390 36.710 45.710 37.010 ;
        RECT 46.460 36.470 46.750 42.260 ;
        RECT 58.720 42.430 58.950 42.720 ;
        RECT 58.720 41.830 58.910 42.430 ;
        RECT 58.260 41.440 58.580 41.720 ;
        RECT 58.720 41.540 58.950 41.830 ;
        RECT 58.720 41.280 58.910 41.540 ;
        RECT 58.440 40.790 58.910 41.280 ;
        RECT 59.300 41.190 59.670 41.200 ;
        RECT 59.250 40.930 59.670 41.190 ;
        RECT 59.300 40.910 59.670 40.930 ;
        RECT 58.720 40.540 58.910 40.790 ;
        RECT 58.440 40.050 58.910 40.540 ;
        RECT 59.300 40.400 59.670 40.420 ;
        RECT 59.250 40.140 59.670 40.400 ;
        RECT 59.300 40.130 59.670 40.140 ;
        RECT 58.260 39.610 58.580 39.890 ;
        RECT 58.720 39.790 58.910 40.050 ;
        RECT 58.720 39.500 58.950 39.790 ;
        RECT 58.720 38.900 58.910 39.500 ;
        RECT 58.260 38.510 58.580 38.790 ;
        RECT 58.720 38.610 58.950 38.900 ;
        RECT 58.720 38.350 58.910 38.610 ;
        RECT 58.440 37.860 58.910 38.350 ;
        RECT 59.300 38.260 59.670 38.270 ;
        RECT 59.250 38.000 59.670 38.260 ;
        RECT 59.300 37.980 59.670 38.000 ;
        RECT 41.840 36.070 42.150 36.140 ;
        RECT 42.330 33.960 42.640 36.470 ;
        RECT 46.270 36.070 46.560 36.120 ;
        RECT 46.760 33.960 47.050 37.780 ;
        RECT 48.220 33.690 48.410 37.780 ;
        RECT 49.530 36.740 49.760 37.820 ;
        RECT 49.440 36.260 49.770 36.740 ;
        RECT 49.530 33.650 49.760 36.260 ;
        RECT 52.500 33.860 52.750 37.840 ;
        RECT 55.820 33.800 55.980 37.850 ;
        RECT 58.570 37.640 58.910 37.860 ;
        RECT 60.030 37.640 60.260 43.690 ;
        RECT 60.750 43.360 61.130 44.130 ;
        RECT 62.490 43.970 62.740 44.270 ;
        RECT 62.500 43.500 62.740 43.970 ;
        RECT 65.800 43.890 66.260 44.280 ;
        RECT 63.000 43.470 63.250 43.690 ;
        RECT 61.760 43.310 62.100 43.360 ;
        RECT 61.760 43.290 62.320 43.310 ;
        RECT 61.640 43.120 62.320 43.290 ;
        RECT 61.760 43.080 62.320 43.120 ;
        RECT 61.760 43.040 62.100 43.080 ;
        RECT 63.000 42.400 63.640 43.470 ;
        RECT 65.860 43.390 66.260 43.890 ;
        RECT 65.850 43.340 66.260 43.390 ;
        RECT 66.270 43.600 66.460 44.460 ;
        RECT 66.670 43.910 66.830 45.240 ;
        RECT 67.650 44.930 67.970 45.250 ;
        RECT 68.280 44.290 68.510 45.270 ;
        RECT 66.630 43.890 66.830 43.910 ;
        RECT 67.650 43.900 67.970 44.220 ;
        RECT 68.280 43.940 68.540 44.290 ;
        RECT 66.620 43.650 66.850 43.890 ;
        RECT 68.300 43.780 68.540 43.940 ;
        RECT 68.610 43.780 68.850 45.780 ;
        RECT 70.790 45.680 71.170 47.600 ;
        RECT 72.540 46.420 72.780 47.600 ;
        RECT 72.530 45.760 72.790 46.420 ;
        RECT 69.500 44.380 69.730 45.270 ;
        RECT 69.480 44.000 70.290 44.380 ;
        RECT 66.270 43.480 66.440 43.600 ;
        RECT 65.850 43.250 66.020 43.340 ;
        RECT 65.860 42.900 66.020 43.250 ;
        RECT 65.850 42.810 66.020 42.900 ;
        RECT 65.850 42.760 66.130 42.810 ;
        RECT 63.000 41.860 63.250 42.400 ;
        RECT 65.860 42.210 66.130 42.760 ;
        RECT 66.270 42.670 66.430 43.480 ;
        RECT 66.630 43.430 66.830 43.650 ;
        RECT 66.670 42.720 66.830 43.430 ;
        RECT 67.650 43.350 67.970 43.670 ;
        RECT 68.300 43.500 68.850 43.780 ;
        RECT 68.910 43.730 69.100 43.780 ;
        RECT 69.310 43.730 69.470 43.780 ;
        RECT 68.340 43.440 68.850 43.500 ;
        RECT 68.610 43.190 68.850 43.440 ;
        RECT 69.910 43.360 70.290 44.000 ;
        RECT 70.790 43.820 71.180 45.680 ;
        RECT 68.600 42.870 68.860 43.190 ;
        RECT 66.270 42.550 66.440 42.670 ;
        RECT 61.760 41.180 62.100 41.220 ;
        RECT 61.760 41.140 62.320 41.180 ;
        RECT 61.640 40.970 62.320 41.140 ;
        RECT 61.760 40.950 62.320 40.970 ;
        RECT 61.760 40.900 62.100 40.950 ;
        RECT 63.000 40.790 63.640 41.860 ;
        RECT 65.860 41.560 66.020 42.210 ;
        RECT 66.270 41.560 66.460 42.550 ;
        RECT 66.630 42.500 66.830 42.720 ;
        RECT 66.620 42.260 66.850 42.500 ;
        RECT 67.650 42.480 67.970 42.800 ;
        RECT 66.630 42.240 66.830 42.260 ;
        RECT 66.670 41.560 66.830 42.240 ;
        RECT 67.650 41.930 67.970 42.250 ;
        RECT 68.610 41.550 68.850 42.870 ;
        RECT 70.790 41.550 71.170 43.820 ;
        RECT 71.250 43.690 71.490 43.780 ;
        RECT 72.540 43.150 72.780 45.760 ;
        RECT 74.820 44.250 75.220 47.600 ;
        RECT 80.420 47.460 80.700 48.110 ;
        RECT 80.950 47.460 81.140 48.920 ;
        RECT 82.350 47.840 82.660 48.280 ;
        RECT 76.020 44.250 76.210 45.230 ;
        RECT 74.190 43.880 74.470 44.200 ;
        RECT 74.620 44.060 76.210 44.250 ;
        RECT 73.430 43.680 73.810 43.780 ;
        RECT 74.250 43.580 74.410 43.880 ;
        RECT 74.620 43.710 74.810 44.060 ;
        RECT 74.820 43.870 75.220 44.060 ;
        RECT 76.460 43.870 76.740 45.320 ;
        RECT 74.820 43.590 76.740 43.870 ;
        RECT 81.180 43.780 81.580 47.600 ;
        RECT 83.620 46.420 83.860 47.600 ;
        RECT 83.610 45.760 83.870 46.420 ;
        RECT 77.460 43.650 77.860 43.780 ;
        RECT 78.540 43.680 78.940 43.780 ;
        RECT 80.980 43.730 81.580 43.780 ;
        RECT 72.530 42.830 72.790 43.150 ;
        RECT 72.540 41.550 72.780 42.830 ;
        RECT 74.820 41.550 75.220 43.590 ;
        RECT 77.860 43.420 78.540 43.640 ;
        RECT 81.180 41.550 81.580 43.730 ;
        RECT 82.590 43.680 82.970 43.780 ;
        RECT 83.620 43.150 83.860 45.760 ;
        RECT 84.650 44.880 85.020 49.360 ;
        RECT 85.460 47.600 85.830 68.340 ;
        RECT 86.210 63.630 86.660 64.060 ;
        RECT 85.230 45.680 85.830 47.600 ;
        RECT 84.620 44.420 85.070 44.880 ;
        RECT 84.650 44.380 85.020 44.420 ;
        RECT 85.220 44.290 85.830 45.680 ;
        RECT 85.220 43.830 85.870 44.290 ;
        RECT 85.220 43.820 85.830 43.830 ;
        RECT 85.230 43.780 85.830 43.820 ;
        RECT 84.910 43.710 85.150 43.780 ;
        RECT 83.610 42.830 83.870 43.150 ;
        RECT 83.620 41.550 83.860 42.830 ;
        RECT 85.230 41.550 85.610 43.780 ;
        RECT 86.230 41.940 86.600 63.630 ;
        RECT 92.780 62.580 93.360 63.140 ;
        RECT 89.570 61.010 90.130 61.660 ;
        RECT 90.520 61.500 91.080 62.080 ;
        RECT 91.600 61.960 92.160 62.550 ;
        RECT 87.100 58.550 87.530 58.990 ;
        RECT 86.770 55.610 86.980 55.720 ;
        RECT 87.110 53.510 87.480 58.550 ;
        RECT 88.650 55.720 88.880 59.540 ;
        RECT 87.650 55.660 87.860 55.720 ;
        RECT 88.650 55.650 88.910 55.720 ;
        RECT 86.780 49.680 87.010 49.800 ;
        RECT 87.110 47.600 87.660 53.510 ;
        RECT 88.650 52.540 88.880 55.650 ;
        RECT 88.640 52.290 88.880 52.540 ;
        RECT 89.590 52.460 90.090 61.010 ;
        RECT 87.110 47.460 87.790 47.600 ;
        RECT 88.650 47.460 88.880 52.290 ;
        RECT 89.450 52.140 90.090 52.460 ;
        RECT 89.590 48.770 90.090 52.140 ;
        RECT 89.480 48.450 90.090 48.770 ;
        RECT 89.590 47.600 90.090 48.450 ;
        RECT 90.520 59.540 91.020 61.500 ;
        RECT 90.520 47.600 91.360 59.540 ;
        RECT 91.390 49.600 91.620 49.680 ;
        RECT 87.110 43.780 87.480 47.460 ;
        RECT 87.550 46.440 87.790 47.460 ;
        RECT 88.430 46.910 88.750 47.230 ;
        RECT 89.570 46.900 90.130 47.600 ;
        RECT 90.380 47.470 91.360 47.600 ;
        RECT 90.380 46.950 91.020 47.470 ;
        RECT 87.530 45.780 87.800 46.440 ;
        RECT 88.430 46.360 88.750 46.680 ;
        RECT 89.550 46.660 90.130 46.900 ;
        RECT 87.550 43.780 87.790 45.780 ;
        RECT 88.430 45.480 88.750 45.800 ;
        RECT 89.570 45.500 90.130 46.660 ;
        RECT 90.270 46.350 91.020 46.950 ;
        RECT 90.380 45.810 91.020 46.350 ;
        RECT 89.550 45.260 90.130 45.500 ;
        RECT 88.430 44.930 88.750 45.250 ;
        RECT 89.570 44.690 90.130 45.260 ;
        RECT 90.270 45.210 91.020 45.810 ;
        RECT 89.570 44.460 90.160 44.690 ;
        RECT 88.430 43.900 88.750 44.220 ;
        RECT 89.570 43.890 90.130 44.460 ;
        RECT 90.380 43.940 91.020 45.210 ;
        RECT 86.930 43.730 87.090 43.780 ;
        RECT 87.110 43.730 87.490 43.780 ;
        RECT 87.550 43.740 87.900 43.780 ;
        RECT 86.200 41.930 86.600 41.940 ;
        RECT 86.190 41.510 86.610 41.930 ;
        RECT 86.230 41.500 86.600 41.510 ;
        RECT 63.000 40.540 63.250 40.790 ;
        RECT 61.760 40.380 62.100 40.430 ;
        RECT 61.760 40.360 62.320 40.380 ;
        RECT 61.640 40.190 62.320 40.360 ;
        RECT 61.760 40.150 62.320 40.190 ;
        RECT 61.760 40.110 62.100 40.150 ;
        RECT 63.000 39.470 63.640 40.540 ;
        RECT 63.000 38.930 63.250 39.470 ;
        RECT 61.760 38.250 62.100 38.290 ;
        RECT 61.760 38.210 62.320 38.250 ;
        RECT 58.570 34.210 58.810 37.640 ;
        RECT 58.550 33.960 58.940 34.210 ;
        RECT 58.690 33.710 58.940 33.960 ;
        RECT 58.440 33.220 58.910 33.710 ;
        RECT 59.300 33.570 59.670 33.590 ;
        RECT 59.250 33.310 59.670 33.570 ;
        RECT 59.300 33.300 59.670 33.310 ;
        RECT 38.350 32.520 38.760 32.850 ;
        RECT 39.090 32.540 39.330 32.940 ;
        RECT 42.030 32.540 42.340 32.940 ;
        RECT 38.900 32.490 39.330 32.540 ;
        RECT 38.350 30.970 38.760 31.300 ;
        RECT 38.350 29.420 38.760 29.750 ;
        RECT 38.350 27.870 38.760 28.200 ;
        RECT 39.090 26.700 39.330 32.490 ;
        RECT 41.840 32.480 42.340 32.540 ;
        RECT 40.510 31.990 40.710 32.010 ;
        RECT 40.510 31.700 40.860 31.990 ;
        RECT 40.510 30.440 40.710 30.460 ;
        RECT 40.510 30.150 40.860 30.440 ;
        RECT 40.510 28.890 40.710 28.910 ;
        RECT 40.510 28.600 40.860 28.890 ;
        RECT 42.030 28.030 42.340 32.480 ;
        RECT 42.590 32.410 42.870 32.740 ;
        RECT 46.460 32.540 46.750 32.940 ;
        RECT 46.270 32.490 46.750 32.540 ;
        RECT 53.850 32.530 54.170 32.870 ;
        RECT 58.260 32.780 58.580 33.060 ;
        RECT 58.720 32.960 58.910 33.220 ;
        RECT 58.720 32.670 58.950 32.960 ;
        RECT 45.390 31.590 45.710 31.890 ;
        RECT 42.590 30.860 42.870 31.190 ;
        RECT 45.390 30.040 45.710 30.340 ;
        RECT 42.590 29.310 42.870 29.640 ;
        RECT 45.390 28.490 45.710 28.790 ;
        RECT 42.590 28.030 42.870 28.090 ;
        RECT 38.900 26.300 39.140 26.350 ;
        RECT 39.390 15.330 39.630 27.960 ;
        RECT 42.030 27.760 42.870 28.030 ;
        RECT 40.510 27.340 40.710 27.360 ;
        RECT 40.510 27.050 40.860 27.340 ;
        RECT 42.030 26.880 42.640 27.760 ;
        RECT 46.460 27.390 46.750 32.490 ;
        RECT 46.760 27.390 47.050 28.010 ;
        RECT 47.260 27.410 47.600 27.730 ;
        RECT 45.390 26.940 45.710 27.240 ;
        RECT 46.460 27.040 47.080 27.390 ;
        RECT 42.030 26.700 42.660 26.880 ;
        RECT 46.460 26.700 46.750 27.040 ;
        RECT 42.290 26.550 42.660 26.700 ;
        RECT 46.760 26.580 47.050 27.040 ;
        RECT 47.260 26.800 47.510 27.410 ;
        RECT 48.220 26.820 48.410 28.020 ;
        RECT 52.500 27.350 52.750 28.080 ;
        RECT 53.930 27.770 54.140 32.530 ;
        RECT 58.720 32.070 58.910 32.670 ;
        RECT 58.260 31.680 58.580 31.960 ;
        RECT 58.720 31.780 58.950 32.070 ;
        RECT 58.720 31.520 58.910 31.780 ;
        RECT 55.190 30.840 55.580 31.090 ;
        RECT 58.440 31.030 58.910 31.520 ;
        RECT 59.300 31.430 59.670 31.440 ;
        RECT 59.250 31.170 59.670 31.430 ;
        RECT 59.300 31.150 59.670 31.170 ;
        RECT 54.470 29.740 54.810 30.080 ;
        RECT 54.510 29.720 54.730 29.740 ;
        RECT 53.900 27.450 54.180 27.770 ;
        RECT 54.510 27.440 54.710 29.720 ;
        RECT 54.970 27.760 55.160 28.260 ;
        RECT 52.470 27.060 52.810 27.350 ;
        RECT 54.470 27.120 54.750 27.440 ;
        RECT 54.930 27.430 55.210 27.760 ;
        RECT 41.840 26.300 42.150 26.370 ;
        RECT 42.330 25.340 42.640 26.550 ;
        RECT 46.190 26.300 47.050 26.580 ;
        RECT 46.110 26.290 47.050 26.300 ;
        RECT 47.210 26.690 47.510 26.800 ;
        RECT 46.110 25.820 46.570 26.290 ;
        RECT 42.280 24.860 42.700 25.340 ;
        RECT 47.210 25.180 47.400 26.690 ;
        RECT 48.160 26.500 48.480 26.820 ;
        RECT 50.840 26.290 51.590 26.480 ;
        RECT 51.090 25.450 51.590 26.290 ;
        RECT 55.400 26.210 55.580 30.840 ;
        RECT 58.720 30.780 58.910 31.030 ;
        RECT 58.440 30.290 58.910 30.780 ;
        RECT 59.300 30.640 59.670 30.660 ;
        RECT 59.250 30.380 59.670 30.640 ;
        RECT 59.300 30.370 59.670 30.380 ;
        RECT 58.260 29.850 58.580 30.130 ;
        RECT 58.720 30.030 58.910 30.290 ;
        RECT 58.720 29.740 58.950 30.030 ;
        RECT 58.720 29.140 58.910 29.740 ;
        RECT 58.260 28.750 58.580 29.030 ;
        RECT 58.720 28.850 58.950 29.140 ;
        RECT 58.720 28.590 58.910 28.850 ;
        RECT 58.440 28.160 58.910 28.590 ;
        RECT 59.300 28.500 59.670 28.510 ;
        RECT 59.250 28.240 59.670 28.500 ;
        RECT 59.300 28.220 59.670 28.240 ;
        RECT 58.440 28.100 58.940 28.160 ;
        RECT 56.720 27.370 56.980 27.400 ;
        RECT 56.700 27.070 57.000 27.370 ;
        RECT 56.720 27.060 56.980 27.070 ;
        RECT 55.400 25.910 55.880 26.210 ;
        RECT 56.730 26.140 56.950 27.060 ;
        RECT 58.690 26.930 58.940 28.100 ;
        RECT 60.030 27.880 60.260 33.930 ;
        RECT 60.750 33.580 61.130 38.070 ;
        RECT 61.640 38.040 62.320 38.210 ;
        RECT 61.760 38.020 62.320 38.040 ;
        RECT 61.760 37.970 62.100 38.020 ;
        RECT 62.500 34.190 62.740 37.930 ;
        RECT 63.000 37.860 63.640 38.930 ;
        RECT 63.000 37.640 63.250 37.860 ;
        RECT 62.500 33.920 62.970 34.190 ;
        RECT 62.700 33.690 62.970 33.920 ;
        RECT 63.000 33.710 63.250 33.930 ;
        RECT 61.760 33.550 62.100 33.600 ;
        RECT 61.760 33.530 62.320 33.550 ;
        RECT 61.640 33.360 62.320 33.530 ;
        RECT 61.760 33.320 62.320 33.360 ;
        RECT 61.760 33.280 62.100 33.320 ;
        RECT 63.000 32.640 63.640 33.710 ;
        RECT 64.780 33.560 65.180 38.090 ;
        RECT 66.440 37.560 66.600 38.210 ;
        RECT 66.440 37.010 66.710 37.560 ;
        RECT 66.430 36.960 66.710 37.010 ;
        RECT 66.850 37.220 67.040 38.210 ;
        RECT 67.250 37.530 67.410 38.210 ;
        RECT 68.300 37.840 68.540 37.930 ;
        RECT 67.210 37.510 67.410 37.530 ;
        RECT 68.230 37.790 68.550 37.840 ;
        RECT 68.230 37.730 68.660 37.790 ;
        RECT 68.910 37.740 69.100 37.800 ;
        RECT 68.230 37.520 68.550 37.730 ;
        RECT 67.200 37.270 67.430 37.510 ;
        RECT 68.300 37.290 68.540 37.520 ;
        RECT 66.850 37.100 67.020 37.220 ;
        RECT 66.430 36.870 66.600 36.960 ;
        RECT 66.440 36.510 66.600 36.870 ;
        RECT 66.430 36.420 66.600 36.510 ;
        RECT 66.430 36.370 66.710 36.420 ;
        RECT 66.440 35.820 66.710 36.370 ;
        RECT 66.850 36.280 67.010 37.100 ;
        RECT 67.210 37.050 67.410 37.270 ;
        RECT 67.250 36.330 67.410 37.050 ;
        RECT 68.230 36.970 68.550 37.290 ;
        RECT 68.300 36.410 68.540 36.970 ;
        RECT 66.850 36.160 67.020 36.280 ;
        RECT 66.440 34.550 66.600 35.820 ;
        RECT 66.850 35.300 67.040 36.160 ;
        RECT 67.210 36.110 67.410 36.330 ;
        RECT 67.200 35.870 67.430 36.110 ;
        RECT 68.230 36.090 68.550 36.410 ;
        RECT 67.210 35.850 67.410 35.870 ;
        RECT 68.300 35.860 68.540 36.090 ;
        RECT 66.820 35.070 67.060 35.300 ;
        RECT 66.440 34.000 66.710 34.550 ;
        RECT 66.430 33.950 66.710 34.000 ;
        RECT 66.850 34.210 67.040 35.070 ;
        RECT 67.250 34.520 67.410 35.850 ;
        RECT 68.230 35.540 68.550 35.860 ;
        RECT 68.300 35.420 68.540 35.540 ;
        RECT 68.300 35.180 68.880 35.420 ;
        RECT 67.210 34.500 67.410 34.520 ;
        RECT 68.230 34.510 68.550 34.830 ;
        RECT 67.200 34.260 67.430 34.500 ;
        RECT 66.850 34.090 67.020 34.210 ;
        RECT 66.430 33.860 66.600 33.950 ;
        RECT 66.440 33.510 66.600 33.860 ;
        RECT 66.430 33.420 66.600 33.510 ;
        RECT 66.430 33.370 66.710 33.420 ;
        RECT 66.440 32.820 66.710 33.370 ;
        RECT 66.850 33.280 67.010 34.090 ;
        RECT 67.210 34.040 67.410 34.260 ;
        RECT 67.250 33.330 67.410 34.040 ;
        RECT 68.230 33.960 68.550 34.280 ;
        RECT 68.640 33.840 68.880 35.180 ;
        RECT 69.310 34.390 69.560 38.210 ;
        RECT 71.370 37.810 71.750 38.210 ;
        RECT 71.250 37.730 71.750 37.810 ;
        RECT 71.370 36.290 71.750 37.730 ;
        RECT 73.320 37.820 73.590 38.210 ;
        RECT 73.320 37.730 73.810 37.820 ;
        RECT 75.400 37.800 75.800 38.210 ;
        RECT 75.180 37.730 75.800 37.800 ;
        RECT 77.460 37.730 77.860 37.850 ;
        RECT 78.540 37.730 78.940 37.850 ;
        RECT 80.980 37.730 81.220 37.800 ;
        RECT 82.590 37.730 82.970 37.880 ;
        RECT 87.110 37.800 87.480 43.730 ;
        RECT 87.550 43.440 88.060 43.740 ;
        RECT 87.550 43.190 87.790 43.440 ;
        RECT 88.430 43.350 88.750 43.670 ;
        RECT 89.550 43.650 90.130 43.890 ;
        RECT 87.540 42.870 87.800 43.190 ;
        RECT 87.550 41.550 87.790 42.870 ;
        RECT 88.430 42.480 88.750 42.800 ;
        RECT 89.570 42.500 90.130 43.650 ;
        RECT 90.270 43.340 91.020 43.940 ;
        RECT 90.380 42.810 91.020 43.340 ;
        RECT 89.550 42.260 90.130 42.500 ;
        RECT 88.430 41.930 88.750 42.250 ;
        RECT 89.570 41.560 90.130 42.260 ;
        RECT 90.270 42.210 91.020 42.810 ;
        RECT 90.380 41.560 91.020 42.210 ;
        RECT 84.910 37.730 85.150 37.790 ;
        RECT 86.930 37.740 87.090 37.800 ;
        RECT 87.110 37.740 87.490 37.800 ;
        RECT 87.740 37.740 87.900 37.800 ;
        RECT 71.370 34.430 71.760 36.290 ;
        RECT 69.100 34.320 69.260 34.390 ;
        RECT 69.310 34.320 69.700 34.390 ;
        RECT 69.910 34.320 70.070 34.390 ;
        RECT 69.310 33.770 69.560 34.320 ;
        RECT 71.370 34.130 71.750 34.430 ;
        RECT 71.370 33.810 71.790 34.130 ;
        RECT 69.290 33.740 69.570 33.770 ;
        RECT 69.280 33.460 69.580 33.740 ;
        RECT 69.290 33.440 69.570 33.460 ;
        RECT 66.850 33.160 67.020 33.280 ;
        RECT 63.000 32.100 63.250 32.640 ;
        RECT 66.440 32.170 66.600 32.820 ;
        RECT 66.850 32.170 67.040 33.160 ;
        RECT 67.210 33.110 67.410 33.330 ;
        RECT 67.200 32.870 67.430 33.110 ;
        RECT 68.230 33.090 68.550 33.410 ;
        RECT 67.210 32.850 67.410 32.870 ;
        RECT 67.250 32.170 67.410 32.850 ;
        RECT 68.230 32.540 68.550 32.860 ;
        RECT 68.240 32.460 68.500 32.540 ;
        RECT 68.230 32.260 68.500 32.460 ;
        RECT 61.760 31.420 62.100 31.460 ;
        RECT 61.760 31.380 62.320 31.420 ;
        RECT 61.640 31.210 62.320 31.380 ;
        RECT 61.760 31.190 62.320 31.210 ;
        RECT 61.760 31.140 62.100 31.190 ;
        RECT 63.000 31.030 63.640 32.100 ;
        RECT 68.230 31.570 68.440 32.260 ;
        RECT 69.310 32.160 69.560 33.440 ;
        RECT 71.370 33.080 71.750 33.810 ;
        RECT 73.320 33.740 73.590 37.730 ;
        RECT 74.030 34.290 74.410 34.390 ;
        RECT 73.300 33.430 73.610 33.740 ;
        RECT 71.370 32.760 71.770 33.080 ;
        RECT 71.370 32.160 71.750 32.760 ;
        RECT 73.320 32.160 73.590 33.430 ;
        RECT 73.760 32.780 74.020 32.840 ;
        RECT 73.750 32.520 74.020 32.780 ;
        RECT 73.240 31.590 73.500 31.910 ;
        RECT 68.220 31.250 68.480 31.570 ;
        RECT 63.000 30.780 63.250 31.030 ;
        RECT 71.510 30.880 71.770 31.200 ;
        RECT 61.760 30.620 62.100 30.670 ;
        RECT 61.760 30.600 62.320 30.620 ;
        RECT 61.640 30.430 62.320 30.600 ;
        RECT 61.760 30.390 62.320 30.430 ;
        RECT 61.760 30.350 62.100 30.390 ;
        RECT 63.000 29.710 63.640 30.780 ;
        RECT 71.510 30.020 71.670 30.880 ;
        RECT 63.000 29.170 63.250 29.710 ;
        RECT 71.350 29.700 71.670 30.020 ;
        RECT 72.770 29.750 73.030 30.070 ;
        RECT 68.140 29.210 68.460 29.530 ;
        RECT 61.760 28.490 62.100 28.530 ;
        RECT 61.760 28.450 62.320 28.490 ;
        RECT 61.640 28.280 62.320 28.450 ;
        RECT 61.760 28.260 62.320 28.280 ;
        RECT 61.760 28.210 62.100 28.260 ;
        RECT 62.700 26.950 62.970 28.180 ;
        RECT 63.000 28.100 63.640 29.170 ;
        RECT 72.270 28.820 72.530 29.140 ;
        RECT 68.190 28.360 68.510 28.680 ;
        RECT 63.000 27.880 63.250 28.100 ;
        RECT 65.520 27.380 65.950 27.780 ;
        RECT 58.680 26.670 59.000 26.930 ;
        RECT 62.700 26.640 63.050 26.950 ;
        RECT 55.480 25.800 55.880 25.910 ;
        RECT 56.670 25.740 57.010 26.140 ;
        RECT 56.730 25.660 56.950 25.740 ;
        RECT 60.680 25.470 61.620 26.400 ;
        RECT 65.560 25.590 65.910 27.380 ;
        RECT 67.380 26.820 67.600 28.140 ;
        RECT 68.640 27.420 68.870 28.140 ;
        RECT 68.640 27.190 71.850 27.420 ;
        RECT 68.640 27.180 68.870 27.190 ;
        RECT 67.090 26.580 67.600 26.820 ;
        RECT 46.770 24.860 47.400 25.180 ;
        RECT 50.600 25.130 50.840 25.450 ;
        RECT 51.840 25.130 52.080 25.450 ;
        RECT 60.410 25.150 60.650 25.470 ;
        RECT 61.650 25.150 61.890 25.470 ;
        RECT 67.090 25.330 67.320 26.580 ;
        RECT 71.620 26.220 71.850 27.190 ;
        RECT 71.570 25.820 71.880 26.220 ;
        RECT 66.980 24.890 67.440 25.330 ;
        RECT 46.770 24.760 47.210 24.860 ;
        RECT 50.600 23.790 50.840 24.110 ;
        RECT 51.840 23.780 52.080 24.100 ;
        RECT 60.410 23.810 60.650 24.130 ;
        RECT 61.650 23.800 61.890 24.120 ;
        RECT 71.620 22.650 71.850 25.820 ;
        RECT 71.490 22.430 71.850 22.650 ;
        RECT 71.290 22.200 71.850 22.430 ;
        RECT 71.290 22.190 71.830 22.200 ;
        RECT 47.680 21.640 48.000 21.960 ;
        RECT 48.770 21.640 49.090 21.960 ;
        RECT 49.870 21.630 50.190 21.950 ;
        RECT 52.490 21.630 52.810 21.950 ;
        RECT 53.590 21.640 53.910 21.960 ;
        RECT 54.680 21.640 55.000 21.960 ;
        RECT 57.490 21.670 57.810 21.990 ;
        RECT 58.580 21.670 58.900 21.990 ;
        RECT 59.680 21.660 60.000 21.980 ;
        RECT 62.300 21.660 62.620 21.980 ;
        RECT 63.400 21.670 63.720 21.990 ;
        RECT 64.490 21.670 64.810 21.990 ;
        RECT 68.790 21.640 69.110 21.960 ;
        RECT 69.890 21.650 70.210 21.970 ;
        RECT 70.980 21.650 71.300 21.970 ;
        RECT 46.980 19.580 47.300 21.330 ;
        RECT 48.230 20.960 48.550 21.280 ;
        RECT 49.320 20.940 49.640 21.260 ;
        RECT 50.600 21.250 50.840 21.340 ;
        RECT 50.430 21.020 50.840 21.250 ;
        RECT 51.840 21.250 52.080 21.330 ;
        RECT 50.430 20.930 50.750 21.020 ;
        RECT 51.840 21.010 52.250 21.250 ;
        RECT 51.930 20.930 52.250 21.010 ;
        RECT 53.040 20.940 53.360 21.260 ;
        RECT 54.130 20.960 54.450 21.280 ;
        RECT 48.230 19.590 48.550 19.910 ;
        RECT 49.320 19.590 49.640 19.910 ;
        RECT 50.420 19.590 50.740 19.910 ;
        RECT 51.940 19.590 52.260 19.910 ;
        RECT 53.040 19.590 53.360 19.910 ;
        RECT 54.130 19.590 54.450 19.910 ;
        RECT 46.860 18.980 47.400 19.580 ;
        RECT 47.670 18.860 47.990 19.180 ;
        RECT 48.770 18.860 49.090 19.180 ;
        RECT 49.870 18.860 50.190 19.180 ;
        RECT 52.490 18.860 52.810 19.180 ;
        RECT 53.590 18.860 53.910 19.180 ;
        RECT 54.690 18.860 55.010 19.180 ;
        RECT 55.350 18.560 55.690 21.350 ;
        RECT 55.290 18.040 55.750 18.560 ;
        RECT 47.670 17.490 47.990 17.810 ;
        RECT 48.770 17.490 49.090 17.810 ;
        RECT 49.870 17.490 50.190 17.810 ;
        RECT 52.490 17.490 52.810 17.810 ;
        RECT 53.590 17.490 53.910 17.810 ;
        RECT 54.690 17.490 55.010 17.810 ;
        RECT 56.780 17.670 57.120 21.340 ;
        RECT 58.040 20.990 58.360 21.310 ;
        RECT 59.130 20.970 59.450 21.290 ;
        RECT 60.410 21.280 60.650 21.360 ;
        RECT 60.240 21.040 60.650 21.280 ;
        RECT 61.650 21.280 61.890 21.360 ;
        RECT 61.650 21.040 62.060 21.280 ;
        RECT 60.240 20.960 60.560 21.040 ;
        RECT 61.740 20.960 62.060 21.040 ;
        RECT 62.850 20.970 63.170 21.290 ;
        RECT 63.940 20.990 64.260 21.310 ;
        RECT 58.040 19.620 58.360 19.940 ;
        RECT 59.130 19.620 59.450 19.940 ;
        RECT 60.230 19.620 60.550 19.940 ;
        RECT 61.750 19.620 62.070 19.940 ;
        RECT 62.850 19.620 63.170 19.940 ;
        RECT 63.940 19.620 64.260 19.940 ;
        RECT 57.480 18.890 57.800 19.210 ;
        RECT 58.580 18.890 58.900 19.210 ;
        RECT 59.680 18.890 60.000 19.210 ;
        RECT 62.300 18.890 62.620 19.210 ;
        RECT 63.400 18.890 63.720 19.210 ;
        RECT 64.500 18.890 64.820 19.210 ;
        RECT 56.690 17.200 57.210 17.670 ;
        RECT 57.480 17.520 57.800 17.840 ;
        RECT 58.580 17.520 58.900 17.840 ;
        RECT 59.680 17.520 60.000 17.840 ;
        RECT 62.300 17.520 62.620 17.840 ;
        RECT 63.400 17.520 63.720 17.840 ;
        RECT 64.500 17.520 64.820 17.840 ;
        RECT 65.200 17.200 65.470 21.380 ;
        RECT 68.230 20.940 68.550 21.260 ;
        RECT 69.340 20.950 69.660 21.270 ;
        RECT 70.430 20.970 70.750 21.290 ;
        RECT 72.270 20.980 72.520 28.820 ;
        RECT 72.770 21.880 73.020 29.750 ;
        RECT 73.250 22.790 73.500 31.590 ;
        RECT 73.750 23.680 74.000 32.520 ;
        RECT 75.400 32.160 75.800 37.730 ;
        RECT 87.110 36.760 87.480 37.740 ;
        RECT 87.070 36.250 87.560 36.760 ;
        RECT 87.110 36.220 87.480 36.250 ;
        RECT 78.060 34.250 78.460 34.390 ;
        RECT 79.580 33.610 79.900 33.930 ;
        RECT 79.730 32.930 80.050 33.250 ;
        RECT 79.730 32.040 80.050 32.360 ;
        RECT 79.580 31.360 79.900 31.680 ;
        RECT 79.580 30.840 79.900 31.160 ;
        RECT 79.730 30.160 80.050 30.480 ;
        RECT 79.730 29.270 80.050 29.590 ;
        RECT 79.580 28.590 79.900 28.910 ;
        RECT 74.030 28.340 74.410 28.440 ;
        RECT 80.660 28.340 80.890 34.390 ;
        RECT 81.920 30.040 82.150 34.390 ;
        RECT 81.880 30.030 82.160 30.040 ;
        RECT 81.880 29.710 82.180 30.030 ;
        RECT 81.920 28.340 82.150 29.710 ;
        RECT 89.590 25.180 90.090 41.560 ;
        RECT 90.520 30.460 91.020 41.560 ;
        RECT 91.650 35.690 92.150 61.960 ;
        RECT 92.780 50.020 93.280 62.580 ;
        RECT 94.890 55.570 95.310 55.720 ;
        RECT 95.920 55.570 96.340 55.720 ;
        RECT 99.620 55.640 99.850 55.720 ;
        RECT 94.890 55.430 96.340 55.570 ;
        RECT 98.100 53.000 98.570 53.490 ;
        RECT 92.550 49.720 93.280 50.020 ;
        RECT 92.780 49.680 93.280 49.720 ;
        RECT 98.150 50.020 98.550 53.000 ;
        RECT 99.070 52.390 99.490 52.750 ;
        RECT 98.150 49.720 98.670 50.020 ;
        RECT 98.150 49.690 98.550 49.720 ;
        RECT 92.610 49.600 93.280 49.680 ;
        RECT 92.780 47.040 93.280 49.600 ;
        RECT 94.900 49.530 96.340 49.690 ;
        RECT 98.150 49.600 98.630 49.690 ;
        RECT 92.640 46.870 93.280 47.040 ;
        RECT 92.780 46.580 93.280 46.870 ;
        RECT 92.620 46.280 93.280 46.580 ;
        RECT 92.650 46.180 93.280 46.280 ;
        RECT 92.780 40.860 93.280 46.180 ;
        RECT 92.730 40.300 93.280 40.860 ;
        RECT 91.640 35.130 92.160 35.690 ;
        RECT 90.510 29.940 91.030 30.460 ;
        RECT 89.430 24.610 90.090 25.180 ;
        RECT 73.700 23.100 74.070 23.680 ;
        RECT 73.170 22.210 73.540 22.790 ;
        RECT 72.680 21.300 73.050 21.880 ;
        RECT 68.240 19.600 68.560 19.920 ;
        RECT 69.340 19.600 69.660 19.920 ;
        RECT 70.430 19.600 70.750 19.920 ;
        RECT 70.940 19.190 71.270 20.760 ;
        RECT 72.210 20.410 72.560 20.980 ;
        RECT 68.790 18.870 69.110 19.190 ;
        RECT 69.890 18.870 70.210 19.190 ;
        RECT 70.940 18.870 71.310 19.190 ;
        RECT 70.940 17.820 71.270 18.870 ;
        RECT 71.710 18.310 71.990 18.840 ;
        RECT 71.710 18.010 72.170 18.310 ;
        RECT 71.700 17.990 72.170 18.010 ;
        RECT 68.790 17.500 69.110 17.820 ;
        RECT 69.890 17.500 70.210 17.820 ;
        RECT 70.940 17.500 71.310 17.820 ;
        RECT 71.700 17.560 71.990 17.990 ;
        RECT 47.100 16.850 47.420 17.170 ;
        RECT 48.230 16.810 48.550 17.130 ;
        RECT 49.320 16.810 49.640 17.130 ;
        RECT 50.420 16.820 50.740 17.140 ;
        RECT 51.940 16.820 52.260 17.140 ;
        RECT 53.040 16.810 53.360 17.130 ;
        RECT 54.130 16.810 54.450 17.130 ;
        RECT 55.260 16.850 55.580 17.170 ;
        RECT 56.690 17.150 57.230 17.200 ;
        RECT 56.910 16.880 57.230 17.150 ;
        RECT 58.040 16.840 58.360 17.160 ;
        RECT 59.130 16.840 59.450 17.160 ;
        RECT 60.230 16.850 60.550 17.170 ;
        RECT 61.750 16.850 62.070 17.170 ;
        RECT 62.850 16.840 63.170 17.160 ;
        RECT 63.940 16.840 64.260 17.160 ;
        RECT 65.070 16.880 65.470 17.200 ;
        RECT 65.200 16.790 65.470 16.880 ;
        RECT 68.240 16.830 68.560 17.150 ;
        RECT 69.340 16.820 69.660 17.140 ;
        RECT 70.430 16.820 70.750 17.140 ;
        RECT 65.090 16.730 65.580 16.790 ;
        RECT 47.110 16.380 47.430 16.700 ;
        RECT 55.250 16.380 55.570 16.700 ;
        RECT 56.920 16.410 57.240 16.730 ;
        RECT 65.060 16.410 65.580 16.730 ;
        RECT 65.090 16.230 65.580 16.410 ;
        RECT 38.990 14.010 39.640 15.330 ;
        RECT 70.940 10.770 71.270 17.500 ;
        RECT 71.560 16.860 71.880 17.180 ;
        RECT 71.550 16.390 71.870 16.710 ;
        RECT 89.590 16.300 90.090 24.610 ;
        RECT 90.520 17.210 91.020 29.940 ;
        RECT 91.650 18.080 92.150 35.130 ;
        RECT 92.780 19.590 93.280 40.300 ;
        RECT 98.150 47.040 98.550 49.600 ;
        RECT 98.150 46.870 98.600 47.040 ;
        RECT 98.150 46.530 98.550 46.870 ;
        RECT 98.150 46.210 98.640 46.530 ;
        RECT 98.150 46.190 98.600 46.210 ;
        RECT 98.150 44.000 98.550 46.190 ;
        RECT 98.150 43.700 98.640 44.000 ;
        RECT 95.670 27.150 96.250 27.710 ;
        RECT 95.700 27.140 96.210 27.150 ;
        RECT 92.780 19.030 93.340 19.590 ;
        RECT 92.780 18.900 93.280 19.030 ;
        RECT 95.700 15.270 96.200 27.140 ;
        RECT 95.070 13.990 96.200 15.270 ;
        RECT 96.950 14.510 97.180 16.580 ;
        RECT 96.940 14.280 97.230 14.510 ;
        RECT 96.950 12.900 97.180 14.280 ;
        RECT 96.940 12.670 97.230 12.900 ;
        RECT 96.950 11.300 97.180 12.670 ;
        RECT 96.940 11.070 97.230 11.300 ;
        RECT 70.880 10.380 71.310 10.770 ;
        RECT 37.340 9.720 37.710 10.100 ;
        RECT 96.950 9.680 97.180 11.070 ;
        RECT 98.150 10.210 98.550 43.700 ;
        RECT 98.150 10.190 98.680 10.210 ;
        RECT 99.080 10.190 99.470 52.390 ;
        RECT 99.880 50.430 100.300 59.540 ;
        RECT 103.580 58.330 103.810 59.540 ;
        RECT 108.580 58.720 108.890 59.160 ;
        RECT 103.580 57.540 103.840 58.330 ;
        RECT 106.000 57.970 106.200 58.000 ;
        RECT 103.580 55.390 103.810 57.540 ;
        RECT 105.910 57.470 106.220 57.970 ;
        RECT 108.730 57.760 109.050 58.080 ;
        RECT 106.000 55.720 106.200 57.470 ;
        RECT 109.510 57.100 109.700 74.500 ;
        RECT 112.850 65.650 113.670 65.740 ;
        RECT 112.790 64.960 113.670 65.650 ;
        RECT 110.100 58.080 110.290 59.540 ;
        RECT 110.540 58.890 110.820 59.540 ;
        RECT 110.430 58.290 110.820 58.890 ;
        RECT 110.100 58.050 110.320 58.080 ;
        RECT 110.080 57.780 110.330 58.050 ;
        RECT 110.090 57.770 110.330 57.780 ;
        RECT 110.090 57.530 110.320 57.770 ;
        RECT 109.510 56.970 109.940 57.100 ;
        RECT 109.510 56.650 109.960 56.970 ;
        RECT 109.510 56.370 109.700 56.650 ;
        RECT 109.510 56.050 109.960 56.370 ;
        RECT 109.510 55.930 109.940 56.050 ;
        RECT 106.000 55.640 106.330 55.720 ;
        RECT 106.580 55.700 106.860 55.720 ;
        RECT 106.580 55.640 106.920 55.700 ;
        RECT 103.580 54.600 103.840 55.390 ;
        RECT 106.000 54.930 106.200 55.640 ;
        RECT 106.600 55.400 106.920 55.640 ;
        RECT 107.260 55.400 107.580 55.720 ;
        RECT 108.330 55.570 108.650 55.700 ;
        RECT 108.260 55.380 108.650 55.570 ;
        RECT 108.830 55.400 109.150 55.720 ;
        RECT 109.510 55.580 109.700 55.930 ;
        RECT 109.390 55.420 109.700 55.580 ;
        RECT 108.260 55.280 108.490 55.380 ;
        RECT 105.850 54.640 106.200 54.930 ;
        RECT 108.280 54.810 108.470 55.280 ;
        RECT 108.730 55.000 109.050 55.320 ;
        RECT 109.310 55.100 109.700 55.420 ;
        RECT 103.580 52.300 103.810 54.600 ;
        RECT 105.860 54.420 106.200 54.640 ;
        RECT 108.210 54.490 108.470 54.810 ;
        RECT 108.480 54.550 108.800 54.870 ;
        RECT 109.390 54.800 109.700 55.100 ;
        RECT 109.870 54.960 110.060 55.830 ;
        RECT 110.130 55.720 110.290 57.530 ;
        RECT 110.540 56.690 110.820 58.290 ;
        RECT 110.540 56.370 110.900 56.690 ;
        RECT 110.540 55.720 110.820 56.370 ;
        RECT 110.130 55.500 110.820 55.720 ;
        RECT 110.930 55.570 111.210 55.720 ;
        RECT 110.090 55.250 110.820 55.500 ;
        RECT 110.080 54.980 110.820 55.250 ;
        RECT 109.220 54.480 109.700 54.800 ;
        RECT 109.850 54.670 110.080 54.960 ;
        RECT 109.260 54.450 109.700 54.480 ;
        RECT 106.000 54.220 106.200 54.420 ;
        RECT 105.860 53.990 106.200 54.210 ;
        RECT 107.370 54.020 107.690 54.340 ;
        RECT 105.850 53.890 106.200 53.990 ;
        RECT 105.850 53.700 106.080 53.890 ;
        RECT 108.210 53.820 108.470 54.140 ;
        RECT 108.580 53.870 108.890 54.310 ;
        RECT 109.510 54.230 109.700 54.450 ;
        RECT 109.220 54.080 109.480 54.150 ;
        RECT 108.590 53.860 108.800 53.870 ;
        RECT 108.280 53.350 108.470 53.820 ;
        RECT 108.570 53.540 108.830 53.860 ;
        RECT 109.220 53.830 109.580 54.080 ;
        RECT 109.870 53.960 110.060 54.670 ;
        RECT 109.260 53.620 109.580 53.830 ;
        RECT 109.850 53.670 110.080 53.960 ;
        RECT 107.260 52.910 107.580 53.230 ;
        RECT 108.260 53.060 108.490 53.350 ;
        RECT 108.590 53.130 108.800 53.540 ;
        RECT 109.390 53.340 109.580 53.620 ;
        RECT 109.390 53.290 109.620 53.340 ;
        RECT 108.830 53.130 109.150 53.230 ;
        RECT 108.100 52.740 108.420 53.060 ;
        RECT 108.580 52.910 109.150 53.130 ;
        RECT 109.310 52.970 109.630 53.290 ;
        RECT 108.580 52.700 108.890 52.910 ;
        RECT 107.260 52.380 107.580 52.700 ;
        RECT 108.580 52.690 109.150 52.700 ;
        RECT 103.580 51.510 103.840 52.300 ;
        RECT 108.260 52.260 108.490 52.550 ;
        RECT 105.850 51.720 106.080 51.910 ;
        RECT 108.280 51.790 108.470 52.260 ;
        RECT 108.590 52.250 108.800 52.690 ;
        RECT 108.830 52.380 109.150 52.690 ;
        RECT 109.390 52.460 109.620 52.560 ;
        RECT 108.570 52.050 108.800 52.250 ;
        RECT 109.310 52.140 109.630 52.460 ;
        RECT 108.570 51.960 109.050 52.050 ;
        RECT 105.850 51.620 106.200 51.720 ;
        RECT 99.880 50.000 100.440 50.430 ;
        RECT 99.620 49.610 99.850 49.690 ;
        RECT 99.880 47.460 100.400 50.000 ;
        RECT 100.850 49.740 101.230 49.750 ;
        RECT 100.830 49.440 101.250 49.740 ;
        RECT 100.010 10.190 100.400 47.460 ;
        RECT 98.150 9.990 100.670 10.190 ;
        RECT 36.690 9.100 37.080 9.490 ;
        RECT 96.940 9.450 97.230 9.680 ;
        RECT 98.150 9.650 98.550 9.990 ;
        RECT 36.090 8.470 36.470 8.860 ;
        RECT 35.500 7.840 35.850 8.210 ;
        RECT 96.950 8.080 97.180 9.450 ;
        RECT 98.140 9.190 98.610 9.650 ;
        RECT 99.080 8.850 99.470 9.990 ;
        RECT 97.670 8.470 97.990 8.550 ;
        RECT 99.050 8.470 99.510 8.850 ;
        RECT 97.670 8.290 99.760 8.470 ;
        RECT 99.250 8.250 99.760 8.290 ;
        RECT 99.470 8.240 99.760 8.250 ;
        RECT 96.940 7.850 97.230 8.080 ;
        RECT 100.010 8.030 100.400 9.990 ;
        RECT 34.860 7.160 35.220 7.540 ;
        RECT 34.270 6.920 34.610 6.930 ;
        RECT 34.250 6.550 34.630 6.920 ;
        RECT 34.270 6.540 34.600 6.550 ;
        RECT 96.950 6.460 97.180 7.850 ;
        RECT 99.990 7.570 100.460 8.030 ;
        RECT 100.500 6.960 100.670 9.990 ;
        RECT 100.850 7.230 101.230 49.440 ;
        RECT 103.580 49.360 103.810 51.510 ;
        RECT 105.860 51.400 106.200 51.620 ;
        RECT 108.210 51.470 108.470 51.790 ;
        RECT 108.730 51.730 109.050 51.960 ;
        RECT 109.390 51.810 109.580 52.140 ;
        RECT 109.870 51.940 110.060 53.670 ;
        RECT 110.100 52.020 110.820 54.980 ;
        RECT 110.080 51.940 110.820 52.020 ;
        RECT 109.260 51.780 109.580 51.810 ;
        RECT 109.220 51.490 109.580 51.780 ;
        RECT 109.850 51.750 110.820 51.940 ;
        RECT 109.850 51.650 110.080 51.750 ;
        RECT 109.220 51.460 109.480 51.490 ;
        RECT 105.860 50.970 106.200 51.190 ;
        RECT 105.850 50.870 106.200 50.970 ;
        RECT 105.850 50.680 106.080 50.870 ;
        RECT 108.210 50.800 108.470 51.120 ;
        RECT 109.220 51.060 109.480 51.130 ;
        RECT 109.870 51.070 110.060 51.650 ;
        RECT 110.090 51.500 110.820 51.750 ;
        RECT 109.220 50.810 109.580 51.060 ;
        RECT 108.280 50.330 108.470 50.800 ;
        RECT 109.260 50.660 109.580 50.810 ;
        RECT 109.390 50.330 109.580 50.660 ;
        RECT 109.700 50.940 110.060 51.070 ;
        RECT 109.700 50.650 110.080 50.940 ;
        RECT 110.130 50.660 110.820 51.500 ;
        RECT 110.940 54.140 111.210 55.570 ;
        RECT 111.560 55.150 111.880 55.470 ;
        RECT 110.940 53.850 111.220 54.140 ;
        RECT 110.940 51.550 111.210 53.850 ;
        RECT 111.610 52.930 111.930 53.250 ;
        RECT 111.600 52.210 111.920 52.530 ;
        RECT 110.940 51.260 111.220 51.550 ;
        RECT 109.700 50.620 110.060 50.650 ;
        RECT 109.870 50.340 110.060 50.620 ;
        RECT 107.260 49.890 107.580 50.210 ;
        RECT 108.260 50.040 108.490 50.330 ;
        RECT 108.830 50.170 109.150 50.210 ;
        RECT 108.740 49.890 109.150 50.170 ;
        RECT 109.310 50.010 109.630 50.330 ;
        RECT 109.700 49.900 110.060 50.340 ;
        RECT 108.740 49.870 109.060 49.890 ;
        RECT 109.870 49.870 110.060 49.900 ;
        RECT 110.130 50.340 110.900 50.660 ;
        RECT 110.130 49.870 110.820 50.340 ;
        RECT 108.740 49.810 110.820 49.870 ;
        RECT 108.790 49.730 110.820 49.810 ;
        RECT 106.140 49.610 106.330 49.720 ;
        RECT 106.580 49.640 106.860 49.720 ;
        RECT 103.580 48.570 103.840 49.360 ;
        RECT 106.580 49.340 106.900 49.640 ;
        RECT 108.330 49.350 108.650 49.670 ;
        RECT 110.130 49.470 110.820 49.730 ;
        RECT 110.940 49.690 111.210 51.260 ;
        RECT 111.520 49.960 111.840 50.280 ;
        RECT 110.930 49.540 111.210 49.690 ;
        RECT 108.730 48.970 109.050 49.290 ;
        RECT 109.310 49.070 109.630 49.390 ;
        RECT 110.090 49.220 110.820 49.470 ;
        RECT 110.080 48.950 110.820 49.220 ;
        RECT 103.580 47.460 103.810 48.570 ;
        RECT 108.480 48.520 108.800 48.840 ;
        RECT 109.260 48.420 109.580 48.740 ;
        RECT 107.370 47.990 107.690 48.310 ;
        RECT 108.580 47.840 108.890 48.280 ;
        RECT 108.590 47.830 108.800 47.840 ;
        RECT 108.570 47.510 108.830 47.830 ;
        RECT 109.260 47.590 109.580 47.910 ;
        RECT 108.100 46.710 108.420 47.030 ;
        RECT 108.590 46.220 108.800 47.510 ;
        RECT 110.100 47.460 110.820 48.950 ;
        RECT 110.940 48.110 111.210 49.540 ;
        RECT 111.560 49.120 111.880 49.440 ;
        RECT 110.940 47.820 111.220 48.110 ;
        RECT 109.310 46.940 109.630 47.260 ;
        RECT 108.570 45.930 108.800 46.220 ;
        RECT 109.310 46.110 109.630 46.430 ;
        RECT 109.260 45.460 109.580 45.780 ;
        RECT 109.260 44.630 109.580 44.950 ;
        RECT 108.760 43.840 109.090 44.130 ;
        RECT 109.310 43.980 109.630 44.300 ;
        RECT 110.270 43.840 110.610 47.460 ;
        RECT 108.750 43.700 110.610 43.840 ;
        RECT 106.140 43.640 106.330 43.690 ;
        RECT 106.580 43.640 106.860 43.690 ;
        RECT 110.270 43.640 110.610 43.700 ;
        RECT 110.940 45.520 111.210 47.820 ;
        RECT 111.610 46.900 111.930 47.220 ;
        RECT 111.600 46.180 111.920 46.500 ;
        RECT 112.790 45.960 113.500 64.960 ;
        RECT 110.940 45.230 111.220 45.520 ;
        RECT 110.940 43.640 111.210 45.230 ;
        RECT 112.660 45.170 113.500 45.960 ;
        RECT 111.520 43.930 111.840 44.250 ;
        RECT 108.380 27.130 109.100 27.700 ;
        RECT 108.440 20.120 108.950 27.130 ;
        RECT 108.300 20.070 108.950 20.120 ;
        RECT 108.290 19.890 108.950 20.070 ;
        RECT 108.260 19.880 108.950 19.890 ;
        RECT 108.260 19.510 108.860 19.880 ;
        RECT 108.260 17.640 108.840 19.510 ;
        RECT 107.910 16.650 108.840 17.640 ;
        RECT 108.260 15.870 108.840 16.650 ;
        RECT 108.270 15.260 108.840 15.870 ;
        RECT 108.260 14.260 108.840 15.260 ;
        RECT 102.450 13.500 102.770 13.820 ;
        RECT 108.270 13.660 108.840 14.260 ;
        RECT 102.450 12.830 102.770 13.150 ;
        RECT 102.570 11.860 102.890 11.910 ;
        RECT 102.340 11.630 102.890 11.860 ;
        RECT 102.570 11.590 102.890 11.630 ;
        RECT 102.570 10.250 102.890 10.300 ;
        RECT 102.340 10.020 102.890 10.250 ;
        RECT 102.570 9.980 102.890 10.020 ;
        RECT 102.560 8.640 102.880 8.690 ;
        RECT 102.330 8.410 102.880 8.640 ;
        RECT 102.560 8.370 102.880 8.410 ;
        RECT 100.080 6.740 100.670 6.960 ;
        RECT 100.820 6.770 101.260 7.230 ;
        RECT 102.560 7.020 102.880 7.070 ;
        RECT 102.330 6.790 102.880 7.020 ;
        RECT 102.560 6.750 102.880 6.790 ;
        RECT 100.080 6.730 100.370 6.740 ;
        RECT 96.940 6.230 97.230 6.460 ;
        RECT 32.490 4.700 32.840 5.030 ;
        RECT 96.950 4.860 97.180 6.230 ;
        RECT 108.260 6.220 108.840 13.660 ;
        RECT 108.270 5.620 108.840 6.220 ;
        RECT 102.560 5.410 102.880 5.460 ;
        RECT 102.330 5.180 102.880 5.410 ;
        RECT 102.560 5.140 102.880 5.180 ;
        RECT 32.510 4.640 32.840 4.700 ;
        RECT 96.940 4.630 97.230 4.860 ;
        RECT 108.260 4.800 108.840 5.620 ;
        RECT 108.260 4.790 108.800 4.800 ;
        RECT 31.220 3.420 31.570 3.750 ;
        RECT 31.220 3.350 31.550 3.420 ;
        RECT 96.950 3.240 97.180 4.630 ;
        RECT 102.190 3.540 102.510 3.860 ;
        RECT 102.240 3.310 102.470 3.540 ;
        RECT 29.080 2.690 30.320 3.020 ;
        RECT 30.610 2.720 31.050 3.140 ;
        RECT 96.940 3.010 97.230 3.240 ;
        RECT 29.080 2.580 29.660 2.690 ;
        RECT 102.570 2.210 102.890 2.260 ;
        RECT 102.340 1.980 102.890 2.210 ;
        RECT 102.570 1.940 102.890 1.980 ;
        RECT 102.560 0.620 102.880 0.670 ;
        RECT 99.360 0.540 99.680 0.590 ;
        RECT 100.300 0.540 100.620 0.590 ;
        RECT 99.130 0.310 99.680 0.540 ;
        RECT 100.070 0.310 100.620 0.540 ;
        RECT 101.250 0.480 101.570 0.530 ;
        RECT 99.360 0.270 99.680 0.310 ;
        RECT 100.300 0.270 100.620 0.310 ;
        RECT 101.020 0.250 101.570 0.480 ;
        RECT 102.330 0.390 102.880 0.620 ;
        RECT 102.560 0.350 102.880 0.390 ;
        RECT 101.250 0.210 101.570 0.250 ;
      LAYER via ;
        RECT 2.030 72.460 2.420 72.850 ;
        RECT 4.450 71.540 4.710 71.800 ;
        RECT 7.310 71.590 7.570 71.850 ;
        RECT 4.440 70.510 4.700 70.770 ;
        RECT 5.160 70.480 5.420 70.740 ;
        RECT 5.850 70.520 6.110 70.780 ;
        RECT 4.440 70.060 4.700 70.320 ;
        RECT 5.850 70.080 6.110 70.340 ;
        RECT 4.440 69.640 4.700 69.900 ;
        RECT 5.160 69.640 5.420 69.900 ;
        RECT 5.870 69.660 6.130 69.920 ;
        RECT 2.110 69.010 2.500 69.400 ;
        RECT 4.440 68.290 4.700 68.550 ;
        RECT 3.490 67.840 3.750 68.100 ;
        RECT 7.000 70.050 7.260 70.310 ;
        RECT 20.550 69.740 20.810 70.000 ;
        RECT 21.910 69.820 22.170 70.080 ;
        RECT 22.600 69.810 22.860 70.070 ;
        RECT 6.580 68.040 6.840 68.300 ;
        RECT 5.140 66.840 5.400 67.100 ;
        RECT 6.570 66.860 6.830 67.120 ;
        RECT 4.350 66.260 4.610 66.520 ;
        RECT 5.280 66.260 5.540 66.520 ;
        RECT 5.980 66.260 6.240 66.520 ;
        RECT 6.720 66.260 6.980 66.520 ;
        RECT 7.430 66.250 7.690 66.510 ;
        RECT 3.410 65.140 3.830 65.560 ;
        RECT 19.830 66.080 20.090 66.340 ;
        RECT 9.360 63.740 9.650 64.320 ;
        RECT 22.650 62.680 22.910 62.940 ;
        RECT 15.830 58.340 16.090 58.600 ;
        RECT 16.920 58.350 17.180 58.610 ;
        RECT 15.360 57.930 15.620 58.190 ;
        RECT 15.830 57.420 16.090 57.680 ;
        RECT 16.920 57.430 17.180 57.690 ;
        RECT 15.360 57.010 15.620 57.270 ;
        RECT 15.830 56.500 16.090 56.760 ;
        RECT 15.360 56.090 15.620 56.350 ;
        RECT 16.570 56.430 16.830 56.690 ;
        RECT 16.920 56.510 17.180 56.770 ;
        RECT 15.640 55.520 15.900 55.780 ;
        RECT 16.540 55.510 16.800 55.770 ;
        RECT 15.640 55.060 15.900 55.320 ;
        RECT 16.940 55.420 17.200 55.680 ;
        RECT 15.640 54.560 15.900 54.820 ;
        RECT 16.550 54.590 16.810 54.850 ;
        RECT 15.640 54.100 15.900 54.360 ;
        RECT 15.640 53.830 15.900 53.860 ;
        RECT 15.640 53.600 16.160 53.830 ;
        RECT 15.900 53.570 16.160 53.600 ;
        RECT 15.640 53.140 15.900 53.400 ;
        RECT 15.860 52.610 16.120 52.870 ;
        RECT 15.900 51.650 16.160 51.910 ;
        RECT 16.940 54.460 17.200 54.720 ;
        RECT 16.940 53.500 17.200 53.760 ;
        RECT 29.690 66.100 29.950 66.360 ;
        RECT 28.440 62.250 28.750 62.560 ;
        RECT 45.020 69.890 45.440 70.310 ;
        RECT 41.170 69.130 41.590 69.550 ;
        RECT 46.690 67.520 47.130 67.960 ;
        RECT 52.410 67.520 52.850 67.960 ;
        RECT 64.790 69.130 66.140 69.550 ;
        RECT 54.230 67.490 54.670 67.930 ;
        RECT 42.270 66.500 42.710 66.940 ;
        RECT 39.510 63.480 39.770 63.740 ;
        RECT 32.440 62.790 32.700 63.050 ;
        RECT 31.270 61.800 31.540 62.060 ;
        RECT 19.940 61.020 20.290 61.370 ;
        RECT 25.190 61.330 25.450 61.590 ;
        RECT 38.460 59.730 38.720 59.990 ;
        RECT 20.960 58.780 21.220 59.170 ;
        RECT 37.360 58.790 37.690 59.050 ;
        RECT 20.320 57.960 20.580 58.360 ;
        RECT 20.340 56.850 20.600 57.110 ;
        RECT 20.340 55.930 20.600 56.190 ;
        RECT 20.310 55.010 20.570 55.270 ;
        RECT 15.860 36.370 16.120 36.840 ;
        RECT 16.500 36.370 16.760 36.840 ;
        RECT 14.500 35.340 14.760 35.600 ;
        RECT 13.980 34.940 14.240 35.200 ;
        RECT 4.700 33.690 5.360 34.350 ;
        RECT 16.580 35.320 16.840 35.580 ;
        RECT 18.340 35.330 18.610 35.600 ;
        RECT 15.920 34.960 16.180 35.220 ;
        RECT 16.670 34.360 16.930 34.620 ;
        RECT 17.320 34.360 17.580 34.620 ;
        RECT 15.450 33.920 15.710 34.180 ;
        RECT 16.150 33.920 16.410 34.180 ;
        RECT 17.830 33.190 18.090 33.450 ;
        RECT 15.000 32.570 15.260 32.830 ;
        RECT 14.000 31.030 14.260 31.290 ;
        RECT 9.910 29.170 10.280 29.540 ;
        RECT 4.740 27.830 5.400 28.490 ;
        RECT 14.000 27.940 14.260 28.200 ;
        RECT 17.750 32.060 18.010 32.320 ;
        RECT 18.840 34.940 19.100 35.200 ;
        RECT 17.760 31.520 18.020 31.780 ;
        RECT 15.000 31.020 15.260 31.280 ;
        RECT 17.810 30.570 18.070 30.830 ;
        RECT 15.480 30.040 15.740 30.300 ;
        RECT 16.170 30.030 16.430 30.290 ;
        RECT 16.650 29.260 16.910 29.520 ;
        RECT 17.360 29.200 17.620 29.460 ;
        RECT 17.310 28.380 17.570 28.640 ;
        RECT 15.100 27.950 15.360 28.210 ;
        RECT 16.190 27.950 16.450 28.210 ;
        RECT 17.320 27.910 17.580 28.170 ;
        RECT 14.550 27.270 14.810 27.530 ;
        RECT 15.650 27.270 15.910 27.530 ;
        RECT 16.750 27.270 17.010 27.530 ;
        RECT 14.550 25.900 14.810 26.160 ;
        RECT 15.650 25.900 15.910 26.160 ;
        RECT 16.750 25.900 17.010 26.160 ;
        RECT 14.000 25.170 14.260 25.430 ;
        RECT 15.100 25.170 15.360 25.430 ;
        RECT 16.190 25.170 16.450 25.430 ;
        RECT 13.990 23.830 14.250 24.090 ;
        RECT 15.100 23.820 15.360 24.080 ;
        RECT 16.190 23.800 16.450 24.060 ;
        RECT 9.900 22.930 10.270 23.300 ;
        RECT 14.550 23.130 14.810 23.390 ;
        RECT 15.650 23.120 15.910 23.380 ;
        RECT 16.740 23.120 17.000 23.380 ;
        RECT 17.440 22.510 17.700 22.870 ;
        RECT 16.600 20.820 16.860 21.080 ;
        RECT 13.290 20.380 13.550 20.640 ;
        RECT 14.390 20.390 14.650 20.650 ;
        RECT 15.480 20.390 15.740 20.650 ;
        RECT 16.610 20.350 16.870 20.610 ;
        RECT 13.840 19.710 14.100 19.970 ;
        RECT 14.940 19.710 15.200 19.970 ;
        RECT 16.040 19.710 16.300 19.970 ;
        RECT 13.840 18.340 14.100 18.600 ;
        RECT 14.940 18.340 15.200 18.600 ;
        RECT 16.040 18.340 16.300 18.600 ;
        RECT 13.290 17.610 13.550 17.870 ;
        RECT 14.390 17.610 14.650 17.870 ;
        RECT 15.480 17.610 15.740 17.870 ;
        RECT 12.890 17.270 13.180 17.560 ;
        RECT 36.730 57.070 37.060 57.400 ;
        RECT 36.160 55.590 36.490 55.920 ;
        RECT 20.950 53.920 21.210 54.180 ;
        RECT 35.520 53.990 35.850 54.320 ;
        RECT 34.880 53.420 35.210 53.750 ;
        RECT 20.960 52.960 21.220 53.220 ;
        RECT 20.950 52.000 21.210 52.260 ;
        RECT 20.310 34.340 20.570 34.600 ;
        RECT 19.690 33.190 19.950 33.450 ;
        RECT 19.270 30.580 19.530 30.840 ;
        RECT 19.710 24.890 19.970 25.310 ;
        RECT 19.670 22.510 19.930 22.870 ;
        RECT 34.270 51.850 34.600 52.180 ;
        RECT 33.640 50.320 33.970 50.650 ;
        RECT 33.080 48.750 33.410 49.080 ;
        RECT 32.460 43.280 32.790 43.610 ;
        RECT 31.830 41.690 32.160 42.020 ;
        RECT 31.210 40.140 31.540 40.470 ;
        RECT 30.610 38.660 30.940 38.990 ;
        RECT 29.970 33.490 30.300 33.820 ;
        RECT 29.300 31.920 29.630 32.250 ;
        RECT 20.950 30.010 21.210 30.270 ;
        RECT 28.680 30.280 29.010 30.610 ;
        RECT 20.290 18.880 20.550 19.210 ;
        RECT 19.260 17.260 19.550 17.550 ;
        RECT 13.280 16.270 13.540 16.530 ;
        RECT 14.390 16.260 14.650 16.520 ;
        RECT 15.480 16.240 15.740 16.500 ;
        RECT 18.100 16.250 18.700 16.850 ;
        RECT 13.840 15.570 14.100 15.830 ;
        RECT 14.940 15.560 15.200 15.820 ;
        RECT 16.030 15.560 16.290 15.820 ;
        RECT 28.000 28.840 28.330 29.170 ;
        RECT 23.960 24.480 24.540 25.190 ;
        RECT 20.880 11.320 21.140 11.660 ;
        RECT 1.970 10.380 2.360 10.770 ;
        RECT 27.970 5.010 28.400 5.440 ;
        RECT 28.620 4.220 29.050 4.650 ;
        RECT 29.290 3.540 29.690 3.940 ;
        RECT 29.120 2.600 29.630 3.110 ;
        RECT 38.460 58.180 38.720 58.440 ;
        RECT 38.460 56.630 38.720 56.890 ;
        RECT 40.560 60.570 40.820 60.830 ;
        RECT 45.420 60.670 45.680 60.930 ;
        RECT 40.560 59.020 40.820 59.280 ;
        RECT 40.560 57.470 40.820 57.730 ;
        RECT 40.560 55.920 40.820 56.180 ;
        RECT 42.600 59.850 42.860 60.110 ;
        RECT 45.420 59.120 45.680 59.380 ;
        RECT 42.600 58.300 42.860 58.560 ;
        RECT 45.420 57.570 45.680 57.830 ;
        RECT 42.600 56.750 42.860 57.010 ;
        RECT 45.420 56.020 45.680 56.280 ;
        RECT 38.460 55.080 38.720 55.340 ;
        RECT 42.600 55.200 42.860 55.460 ;
        RECT 47.980 66.500 48.420 66.940 ;
        RECT 62.380 66.500 62.820 66.940 ;
        RECT 56.630 62.720 56.890 62.980 ;
        RECT 54.750 59.190 55.010 59.450 ;
        RECT 60.220 61.810 60.480 62.070 ;
        RECT 57.090 60.790 57.350 61.050 ;
        RECT 57.510 58.700 57.770 58.960 ;
        RECT 58.570 58.220 58.830 58.480 ;
        RECT 63.390 62.730 63.650 62.990 ;
        RECT 62.950 61.820 63.210 62.080 ;
        RECT 59.380 53.140 59.640 53.400 ;
        RECT 38.460 52.460 38.720 52.720 ;
        RECT 38.460 50.910 38.720 51.170 ;
        RECT 38.460 49.360 38.720 49.620 ;
        RECT 38.460 47.810 38.720 48.070 ;
        RECT 40.560 51.620 40.820 51.880 ;
        RECT 40.560 50.070 40.820 50.330 ;
        RECT 40.560 48.520 40.820 48.780 ;
        RECT 42.600 52.340 42.860 52.600 ;
        RECT 58.290 52.620 58.550 52.880 ;
        RECT 45.420 51.520 45.680 51.780 ;
        RECT 42.600 50.790 42.860 51.050 ;
        RECT 45.420 49.970 45.680 50.230 ;
        RECT 42.600 49.240 42.860 49.500 ;
        RECT 45.420 48.420 45.680 48.680 ;
        RECT 42.600 47.690 42.860 47.950 ;
        RECT 40.560 46.970 40.820 47.230 ;
        RECT 45.420 46.870 45.680 47.130 ;
        RECT 58.290 51.520 58.550 51.780 ;
        RECT 68.180 66.460 68.620 66.900 ;
        RECT 76.510 67.490 76.790 67.930 ;
        RECT 72.730 60.830 73.950 61.090 ;
        RECT 69.490 60.180 69.750 60.440 ;
        RECT 75.820 59.640 76.080 59.900 ;
        RECT 78.160 62.730 78.420 62.990 ;
        RECT 77.270 61.860 77.530 62.120 ;
        RECT 84.680 71.830 85.050 72.200 ;
        RECT 80.830 63.440 81.090 63.710 ;
        RECT 77.270 57.650 77.530 57.910 ;
        RECT 78.290 57.660 78.550 57.920 ;
        RECT 82.370 58.750 82.630 59.010 ;
        RECT 81.040 57.540 81.470 57.970 ;
        RECT 81.980 57.220 82.240 57.480 ;
        RECT 81.270 56.390 81.530 56.650 ;
        RECT 81.970 55.530 82.230 55.790 ;
        RECT 61.790 53.140 62.050 53.400 ;
        RECT 59.380 51.000 59.640 51.260 ;
        RECT 60.210 51.120 60.480 51.390 ;
        RECT 59.380 50.210 59.640 50.470 ;
        RECT 58.290 49.690 58.550 49.950 ;
        RECT 58.290 48.590 58.550 48.850 ;
        RECT 59.380 48.070 59.640 48.330 ;
        RECT 61.790 51.000 62.050 51.260 ;
        RECT 61.790 50.210 62.050 50.470 ;
        RECT 61.790 48.070 62.050 48.330 ;
        RECT 82.370 54.020 82.630 54.280 ;
        RECT 85.500 68.370 85.870 68.740 ;
        RECT 84.360 55.420 84.620 55.680 ;
        RECT 82.370 52.720 82.630 52.980 ;
        RECT 82.220 51.760 82.480 52.020 ;
        RECT 81.280 50.650 81.540 50.910 ;
        RECT 81.280 50.050 81.540 50.310 ;
        RECT 84.410 49.370 84.670 49.630 ;
        RECT 82.220 49.000 82.480 49.260 ;
        RECT 67.680 46.940 67.940 47.200 ;
        RECT 67.680 46.390 67.940 46.650 ;
        RECT 56.850 44.480 57.130 44.760 ;
        RECT 67.680 45.510 67.940 45.770 ;
        RECT 59.380 43.070 59.640 43.330 ;
        RECT 38.460 42.330 38.720 42.590 ;
        RECT 38.460 40.780 38.720 41.040 ;
        RECT 38.460 39.230 38.720 39.490 ;
        RECT 38.460 37.680 38.720 37.940 ;
        RECT 40.560 41.490 40.820 41.750 ;
        RECT 40.560 39.940 40.820 40.200 ;
        RECT 40.560 38.390 40.820 38.650 ;
        RECT 42.600 42.210 42.860 42.470 ;
        RECT 58.290 42.550 58.550 42.810 ;
        RECT 45.420 41.390 45.680 41.650 ;
        RECT 42.600 40.660 42.860 40.920 ;
        RECT 45.420 39.840 45.680 40.100 ;
        RECT 42.600 39.110 42.860 39.370 ;
        RECT 45.420 38.290 45.680 38.550 ;
        RECT 42.600 37.560 42.860 37.820 ;
        RECT 40.560 36.840 40.820 37.100 ;
        RECT 45.420 36.740 45.680 37.000 ;
        RECT 58.290 41.450 58.550 41.710 ;
        RECT 59.380 40.930 59.640 41.190 ;
        RECT 59.380 40.140 59.640 40.400 ;
        RECT 58.290 39.620 58.550 39.880 ;
        RECT 58.290 38.520 58.550 38.780 ;
        RECT 59.380 38.000 59.640 38.260 ;
        RECT 49.480 36.290 49.740 36.700 ;
        RECT 61.790 43.070 62.050 43.330 ;
        RECT 67.680 44.960 67.940 45.220 ;
        RECT 67.680 43.930 67.940 44.190 ;
        RECT 67.680 43.380 67.940 43.640 ;
        RECT 68.370 43.460 68.630 43.720 ;
        RECT 68.600 42.900 68.860 43.160 ;
        RECT 61.790 40.930 62.050 41.190 ;
        RECT 67.680 42.510 67.940 42.770 ;
        RECT 67.680 41.960 67.940 42.220 ;
        RECT 82.370 47.990 82.630 48.250 ;
        RECT 74.200 43.910 74.460 44.170 ;
        RECT 72.530 42.860 72.790 43.120 ;
        RECT 86.270 63.660 86.640 64.030 ;
        RECT 84.690 44.460 85.060 44.830 ;
        RECT 85.460 43.870 85.830 44.240 ;
        RECT 83.610 42.860 83.870 43.120 ;
        RECT 92.820 62.610 93.320 63.110 ;
        RECT 89.600 61.050 90.100 61.550 ;
        RECT 90.550 61.540 91.050 62.040 ;
        RECT 91.630 62.010 92.130 62.510 ;
        RECT 87.150 58.590 87.520 58.960 ;
        RECT 89.480 52.170 89.740 52.430 ;
        RECT 89.510 48.480 89.770 48.740 ;
        RECT 88.460 46.940 88.720 47.200 ;
        RECT 88.460 46.390 88.720 46.650 ;
        RECT 88.460 45.510 88.720 45.770 ;
        RECT 88.460 44.960 88.720 45.220 ;
        RECT 88.460 43.930 88.720 44.190 ;
        RECT 86.200 41.540 86.570 41.910 ;
        RECT 61.790 40.140 62.050 40.400 ;
        RECT 59.380 33.310 59.640 33.570 ;
        RECT 38.460 32.560 38.720 32.820 ;
        RECT 38.460 31.010 38.720 31.270 ;
        RECT 38.460 29.460 38.720 29.720 ;
        RECT 38.460 27.910 38.720 28.170 ;
        RECT 40.560 31.720 40.820 31.980 ;
        RECT 40.560 30.170 40.820 30.430 ;
        RECT 40.560 28.620 40.820 28.880 ;
        RECT 42.600 32.440 42.860 32.700 ;
        RECT 53.880 32.570 54.140 32.830 ;
        RECT 58.290 32.790 58.550 33.050 ;
        RECT 45.420 31.620 45.680 31.880 ;
        RECT 42.600 30.890 42.860 31.150 ;
        RECT 45.420 30.070 45.680 30.330 ;
        RECT 42.600 29.340 42.860 29.600 ;
        RECT 45.420 28.520 45.680 28.780 ;
        RECT 42.600 27.790 42.860 28.050 ;
        RECT 40.560 27.070 40.820 27.330 ;
        RECT 47.300 27.440 47.560 27.700 ;
        RECT 45.420 26.970 45.680 27.230 ;
        RECT 46.760 27.070 47.050 27.360 ;
        RECT 42.320 26.560 42.630 26.870 ;
        RECT 58.290 31.690 58.550 31.950 ;
        RECT 59.380 31.170 59.640 31.430 ;
        RECT 54.510 29.790 54.770 30.050 ;
        RECT 53.910 27.480 54.170 27.740 ;
        RECT 54.940 27.470 55.200 27.730 ;
        RECT 52.510 27.070 52.770 27.330 ;
        RECT 54.480 27.150 54.740 27.410 ;
        RECT 46.130 25.850 46.550 26.270 ;
        RECT 42.280 24.890 42.700 25.310 ;
        RECT 48.190 26.530 48.450 26.790 ;
        RECT 59.380 30.380 59.640 30.640 ;
        RECT 58.290 29.860 58.550 30.120 ;
        RECT 58.290 28.760 58.550 29.020 ;
        RECT 59.380 28.240 59.640 28.500 ;
        RECT 56.720 27.090 56.980 27.350 ;
        RECT 55.520 25.840 55.850 26.170 ;
        RECT 61.790 38.000 62.050 38.260 ;
        RECT 61.790 33.310 62.050 33.570 ;
        RECT 68.260 37.550 68.520 37.810 ;
        RECT 68.260 37.000 68.520 37.260 ;
        RECT 68.260 36.120 68.520 36.380 ;
        RECT 68.260 35.570 68.520 35.830 ;
        RECT 68.260 34.540 68.520 34.800 ;
        RECT 68.260 33.990 68.520 34.250 ;
        RECT 87.770 43.460 88.030 43.720 ;
        RECT 88.460 43.380 88.720 43.640 ;
        RECT 87.540 42.900 87.800 43.160 ;
        RECT 88.460 42.510 88.720 42.770 ;
        RECT 88.460 41.960 88.720 42.220 ;
        RECT 71.530 33.840 71.790 34.100 ;
        RECT 69.300 33.470 69.560 33.730 ;
        RECT 68.260 33.120 68.520 33.380 ;
        RECT 68.260 32.570 68.520 32.830 ;
        RECT 68.240 32.290 68.500 32.550 ;
        RECT 61.790 31.170 62.050 31.430 ;
        RECT 73.320 33.450 73.590 33.710 ;
        RECT 71.510 32.790 71.770 33.050 ;
        RECT 73.760 32.550 74.020 32.810 ;
        RECT 73.240 31.620 73.500 31.880 ;
        RECT 68.220 31.280 68.480 31.540 ;
        RECT 71.510 30.910 71.770 31.170 ;
        RECT 61.790 30.380 62.050 30.640 ;
        RECT 71.350 29.730 71.610 29.990 ;
        RECT 72.770 29.780 73.030 30.040 ;
        RECT 68.170 29.240 68.430 29.500 ;
        RECT 61.790 28.240 62.050 28.500 ;
        RECT 72.270 28.850 72.530 29.110 ;
        RECT 68.220 28.390 68.480 28.650 ;
        RECT 65.560 27.400 65.910 27.750 ;
        RECT 58.710 26.670 58.970 26.930 ;
        RECT 62.750 26.640 63.020 26.910 ;
        RECT 56.670 25.770 57.010 26.110 ;
        RECT 65.600 25.630 65.860 25.950 ;
        RECT 71.590 25.850 71.850 26.190 ;
        RECT 46.810 24.800 47.130 25.120 ;
        RECT 67.020 24.920 67.400 25.300 ;
        RECT 47.710 21.670 47.970 21.930 ;
        RECT 48.800 21.670 49.060 21.930 ;
        RECT 49.900 21.660 50.160 21.920 ;
        RECT 52.520 21.660 52.780 21.920 ;
        RECT 53.620 21.670 53.880 21.930 ;
        RECT 54.710 21.670 54.970 21.930 ;
        RECT 57.520 21.700 57.780 21.960 ;
        RECT 58.610 21.700 58.870 21.960 ;
        RECT 59.710 21.690 59.970 21.950 ;
        RECT 62.330 21.690 62.590 21.950 ;
        RECT 63.430 21.700 63.690 21.960 ;
        RECT 64.520 21.700 64.780 21.960 ;
        RECT 68.820 21.670 69.080 21.930 ;
        RECT 69.920 21.680 70.180 21.940 ;
        RECT 71.010 21.680 71.270 21.940 ;
        RECT 48.260 20.990 48.520 21.250 ;
        RECT 49.350 20.970 49.610 21.230 ;
        RECT 50.460 20.960 50.720 21.220 ;
        RECT 51.960 20.960 52.220 21.220 ;
        RECT 53.070 20.970 53.330 21.230 ;
        RECT 54.160 20.990 54.420 21.250 ;
        RECT 48.260 19.620 48.520 19.880 ;
        RECT 49.350 19.620 49.610 19.880 ;
        RECT 50.450 19.620 50.710 19.880 ;
        RECT 51.970 19.620 52.230 19.880 ;
        RECT 53.070 19.620 53.330 19.880 ;
        RECT 54.160 19.620 54.420 19.880 ;
        RECT 46.910 19.020 47.370 19.480 ;
        RECT 47.700 18.890 47.960 19.150 ;
        RECT 48.800 18.890 49.060 19.150 ;
        RECT 49.900 18.890 50.160 19.150 ;
        RECT 52.520 18.890 52.780 19.150 ;
        RECT 53.620 18.890 53.880 19.150 ;
        RECT 54.720 18.890 54.980 19.150 ;
        RECT 55.290 18.070 55.750 18.530 ;
        RECT 47.700 17.520 47.960 17.780 ;
        RECT 48.800 17.520 49.060 17.780 ;
        RECT 49.900 17.520 50.160 17.780 ;
        RECT 52.520 17.520 52.780 17.780 ;
        RECT 53.620 17.520 53.880 17.780 ;
        RECT 54.720 17.520 54.980 17.780 ;
        RECT 58.070 21.020 58.330 21.280 ;
        RECT 59.160 21.000 59.420 21.260 ;
        RECT 60.270 20.990 60.530 21.250 ;
        RECT 61.770 20.990 62.030 21.250 ;
        RECT 62.880 21.000 63.140 21.260 ;
        RECT 63.970 21.020 64.230 21.280 ;
        RECT 58.070 19.650 58.330 19.910 ;
        RECT 59.160 19.650 59.420 19.910 ;
        RECT 60.260 19.650 60.520 19.910 ;
        RECT 61.780 19.650 62.040 19.910 ;
        RECT 62.880 19.650 63.140 19.910 ;
        RECT 63.970 19.650 64.230 19.910 ;
        RECT 57.510 18.920 57.770 19.180 ;
        RECT 58.610 18.920 58.870 19.180 ;
        RECT 59.710 18.920 59.970 19.180 ;
        RECT 62.330 18.920 62.590 19.180 ;
        RECT 63.430 18.920 63.690 19.180 ;
        RECT 64.530 18.920 64.790 19.180 ;
        RECT 56.720 17.180 57.180 17.640 ;
        RECT 57.510 17.550 57.770 17.810 ;
        RECT 58.610 17.550 58.870 17.810 ;
        RECT 59.710 17.550 59.970 17.810 ;
        RECT 62.330 17.550 62.590 17.810 ;
        RECT 63.430 17.550 63.690 17.810 ;
        RECT 64.530 17.550 64.790 17.810 ;
        RECT 68.260 20.970 68.520 21.230 ;
        RECT 69.370 20.980 69.630 21.240 ;
        RECT 70.460 21.000 70.720 21.260 ;
        RECT 87.130 36.290 87.500 36.700 ;
        RECT 79.610 33.640 79.870 33.900 ;
        RECT 79.760 32.960 80.020 33.220 ;
        RECT 79.760 32.070 80.020 32.330 ;
        RECT 79.610 31.390 79.870 31.650 ;
        RECT 79.610 30.870 79.870 31.130 ;
        RECT 79.760 30.190 80.020 30.450 ;
        RECT 79.760 29.300 80.020 29.560 ;
        RECT 79.610 28.620 79.870 28.880 ;
        RECT 81.890 29.740 82.160 30.010 ;
        RECT 98.120 53.030 98.520 53.430 ;
        RECT 92.580 49.740 92.840 50.000 ;
        RECT 99.100 52.390 99.460 52.750 ;
        RECT 98.380 49.740 98.640 50.000 ;
        RECT 92.650 46.300 92.910 46.560 ;
        RECT 92.730 40.330 93.230 40.830 ;
        RECT 91.650 35.140 92.150 35.610 ;
        RECT 90.520 29.950 91.020 30.450 ;
        RECT 89.470 24.650 89.970 25.150 ;
        RECT 73.740 23.140 74.000 23.640 ;
        RECT 73.200 22.240 73.460 22.740 ;
        RECT 72.730 21.340 72.990 21.840 ;
        RECT 68.270 19.630 68.530 19.890 ;
        RECT 69.370 19.630 69.630 19.890 ;
        RECT 70.460 19.630 70.720 19.890 ;
        RECT 72.250 20.440 72.510 20.940 ;
        RECT 68.820 18.900 69.080 19.160 ;
        RECT 69.920 18.900 70.180 19.160 ;
        RECT 71.020 18.900 71.280 19.160 ;
        RECT 68.820 17.530 69.080 17.790 ;
        RECT 69.920 17.530 70.180 17.790 ;
        RECT 71.020 17.530 71.280 17.790 ;
        RECT 47.130 16.880 47.390 17.140 ;
        RECT 48.260 16.840 48.520 17.100 ;
        RECT 49.350 16.840 49.610 17.100 ;
        RECT 50.450 16.850 50.710 17.110 ;
        RECT 51.970 16.850 52.230 17.110 ;
        RECT 53.070 16.840 53.330 17.100 ;
        RECT 54.160 16.840 54.420 17.100 ;
        RECT 55.290 16.880 55.550 17.140 ;
        RECT 56.940 16.910 57.200 17.170 ;
        RECT 58.070 16.870 58.330 17.130 ;
        RECT 59.160 16.870 59.420 17.130 ;
        RECT 60.260 16.880 60.520 17.140 ;
        RECT 61.780 16.880 62.040 17.140 ;
        RECT 62.880 16.870 63.140 17.130 ;
        RECT 63.970 16.870 64.230 17.130 ;
        RECT 65.100 16.910 65.360 17.170 ;
        RECT 68.270 16.860 68.530 17.120 ;
        RECT 69.370 16.850 69.630 17.110 ;
        RECT 70.460 16.850 70.720 17.110 ;
        RECT 47.140 16.410 47.400 16.670 ;
        RECT 55.280 16.410 55.540 16.670 ;
        RECT 56.950 16.440 57.210 16.700 ;
        RECT 65.110 16.700 65.570 16.730 ;
        RECT 65.090 16.440 65.570 16.700 ;
        RECT 65.110 16.270 65.570 16.440 ;
        RECT 39.040 14.040 39.300 15.160 ;
        RECT 71.590 16.890 71.850 17.150 ;
        RECT 98.350 46.240 98.610 46.500 ;
        RECT 98.350 43.720 98.610 43.980 ;
        RECT 95.710 27.170 96.210 27.670 ;
        RECT 92.840 19.060 93.340 19.560 ;
        RECT 91.650 18.110 92.150 18.570 ;
        RECT 90.520 17.240 91.020 17.700 ;
        RECT 71.580 16.420 71.840 16.680 ;
        RECT 89.590 16.330 90.090 16.790 ;
        RECT 95.130 14.040 96.070 15.160 ;
        RECT 70.920 10.410 71.250 10.740 ;
        RECT 37.360 9.750 37.690 10.080 ;
        RECT 108.610 58.750 108.870 59.010 ;
        RECT 105.950 57.510 106.210 57.940 ;
        RECT 108.760 57.790 109.020 58.050 ;
        RECT 112.900 65.000 113.610 65.710 ;
        RECT 109.700 56.680 109.960 56.940 ;
        RECT 109.700 56.080 109.960 56.340 ;
        RECT 106.630 55.420 106.890 55.680 ;
        RECT 107.290 55.430 107.550 55.690 ;
        RECT 108.360 55.410 108.620 55.670 ;
        RECT 108.860 55.430 109.120 55.690 ;
        RECT 108.760 55.030 109.020 55.290 ;
        RECT 109.340 55.130 109.600 55.390 ;
        RECT 105.940 54.450 106.200 54.710 ;
        RECT 108.210 54.520 108.470 54.780 ;
        RECT 108.510 54.580 108.770 54.840 ;
        RECT 110.640 56.400 110.900 56.660 ;
        RECT 109.220 54.740 109.480 54.770 ;
        RECT 109.220 54.510 109.550 54.740 ;
        RECT 109.290 54.480 109.550 54.510 ;
        RECT 105.940 53.920 106.200 54.180 ;
        RECT 107.400 54.050 107.660 54.310 ;
        RECT 108.210 53.850 108.470 54.110 ;
        RECT 108.610 54.020 108.870 54.280 ;
        RECT 109.220 53.910 109.480 54.120 ;
        RECT 109.220 53.860 109.550 53.910 ;
        RECT 108.570 53.570 108.830 53.830 ;
        RECT 109.290 53.650 109.550 53.860 ;
        RECT 107.290 52.940 107.550 53.200 ;
        RECT 108.130 52.770 108.390 53.030 ;
        RECT 108.860 52.980 109.120 53.200 ;
        RECT 108.610 52.940 109.120 52.980 ;
        RECT 109.340 53.000 109.600 53.260 ;
        RECT 108.610 52.720 108.870 52.940 ;
        RECT 107.290 52.410 107.550 52.670 ;
        RECT 108.860 52.410 109.120 52.670 ;
        RECT 109.340 52.170 109.600 52.430 ;
        RECT 100.020 50.020 100.410 50.410 ;
        RECT 100.850 49.460 101.230 49.720 ;
        RECT 36.740 9.130 37.070 9.460 ;
        RECT 36.110 8.500 36.440 8.830 ;
        RECT 35.510 7.870 35.840 8.200 ;
        RECT 98.180 9.220 98.580 9.620 ;
        RECT 97.700 8.290 97.960 8.550 ;
        RECT 99.090 8.420 99.480 8.810 ;
        RECT 34.870 7.190 35.200 7.520 ;
        RECT 34.270 6.570 34.600 6.900 ;
        RECT 100.020 7.600 100.410 7.990 ;
        RECT 105.940 51.430 106.200 51.690 ;
        RECT 108.210 51.500 108.470 51.760 ;
        RECT 108.760 51.760 109.020 52.020 ;
        RECT 109.290 51.750 109.550 51.780 ;
        RECT 109.220 51.520 109.550 51.750 ;
        RECT 105.940 50.900 106.200 51.160 ;
        RECT 108.210 50.830 108.470 51.090 ;
        RECT 109.220 50.950 109.480 51.100 ;
        RECT 109.220 50.840 109.550 50.950 ;
        RECT 109.290 50.690 109.550 50.840 ;
        RECT 111.590 55.180 111.850 55.440 ;
        RECT 111.640 52.960 111.900 53.220 ;
        RECT 111.630 52.240 111.890 52.500 ;
        RECT 107.290 49.920 107.550 50.180 ;
        RECT 108.860 50.150 109.120 50.180 ;
        RECT 108.770 49.920 109.120 50.150 ;
        RECT 109.340 50.040 109.600 50.300 ;
        RECT 109.700 50.050 109.960 50.310 ;
        RECT 108.770 49.890 109.030 49.920 ;
        RECT 110.640 50.370 110.900 50.630 ;
        RECT 106.610 49.360 106.870 49.620 ;
        RECT 108.360 49.380 108.620 49.640 ;
        RECT 111.550 49.990 111.810 50.250 ;
        RECT 108.760 49.000 109.020 49.260 ;
        RECT 109.340 49.100 109.600 49.360 ;
        RECT 108.510 48.550 108.770 48.810 ;
        RECT 109.290 48.450 109.550 48.710 ;
        RECT 107.400 48.020 107.660 48.280 ;
        RECT 108.610 47.990 108.870 48.250 ;
        RECT 108.570 47.540 108.830 47.800 ;
        RECT 109.290 47.620 109.550 47.880 ;
        RECT 108.130 46.740 108.390 47.000 ;
        RECT 111.590 49.150 111.850 49.410 ;
        RECT 109.340 46.970 109.600 47.230 ;
        RECT 109.340 46.140 109.600 46.400 ;
        RECT 109.290 45.490 109.550 45.750 ;
        RECT 109.290 44.660 109.550 44.920 ;
        RECT 108.790 43.850 109.060 44.110 ;
        RECT 109.340 44.010 109.600 44.270 ;
        RECT 111.640 46.930 111.900 47.190 ;
        RECT 111.630 46.210 111.890 46.470 ;
        RECT 112.710 45.210 113.420 45.920 ;
        RECT 111.550 43.960 111.810 44.220 ;
        RECT 108.510 27.160 109.020 27.670 ;
        RECT 102.480 13.530 102.740 13.790 ;
        RECT 102.480 12.860 102.740 13.120 ;
        RECT 102.600 11.620 102.860 11.880 ;
        RECT 102.600 10.010 102.860 10.270 ;
        RECT 102.590 8.400 102.850 8.660 ;
        RECT 100.840 6.810 101.220 7.190 ;
        RECT 102.590 6.780 102.850 7.040 ;
        RECT 33.670 5.930 34.000 6.260 ;
        RECT 33.090 5.360 33.420 5.690 ;
        RECT 32.510 4.670 32.840 5.000 ;
        RECT 102.590 5.170 102.850 5.430 ;
        RECT 31.860 4.030 32.190 4.360 ;
        RECT 31.220 3.380 31.550 3.720 ;
        RECT 102.220 3.570 102.480 3.830 ;
        RECT 30.640 2.740 31.010 3.110 ;
        RECT 102.600 1.970 102.860 2.230 ;
        RECT 99.390 0.300 99.650 0.560 ;
        RECT 100.330 0.300 100.590 0.560 ;
        RECT 101.280 0.240 101.540 0.500 ;
        RECT 102.590 0.380 102.850 0.640 ;
      LAYER met2 ;
        RECT 7.280 71.800 7.600 71.850 ;
        RECT 4.420 71.560 7.600 71.800 ;
        RECT 4.420 71.540 4.740 71.560 ;
        RECT 46.790 61.080 46.900 61.280 ;
        RECT 45.390 60.880 45.710 60.930 ;
        RECT 45.390 60.680 47.020 60.880 ;
        RECT 45.390 60.670 45.710 60.680 ;
        RECT 38.100 60.100 38.190 60.420 ;
        RECT 38.290 59.700 38.750 60.020 ;
        RECT 75.790 59.870 76.100 59.930 ;
        RECT 47.490 59.860 76.100 59.870 ;
        RECT 46.790 59.530 46.900 59.730 ;
        RECT 47.160 59.670 76.100 59.860 ;
        RECT 47.160 59.660 47.740 59.670 ;
        RECT 75.790 59.610 76.100 59.670 ;
        RECT 54.720 59.400 55.040 59.450 ;
        RECT 45.390 59.330 45.710 59.380 ;
        RECT 40.560 58.510 40.820 59.310 ;
        RECT 45.390 59.130 47.020 59.330 ;
        RECT 49.720 59.200 55.090 59.400 ;
        RECT 45.390 59.120 45.710 59.130 ;
        RECT 42.560 58.510 42.900 58.570 ;
        RECT 38.290 58.150 38.750 58.470 ;
        RECT 40.460 58.290 42.900 58.510 ;
        RECT 49.720 58.320 49.920 59.200 ;
        RECT 54.720 59.190 55.040 59.200 ;
        RECT 57.480 58.960 57.790 58.970 ;
        RECT 57.480 58.930 57.800 58.960 ;
        RECT 47.480 58.310 49.920 58.320 ;
        RECT 46.790 57.980 46.900 58.180 ;
        RECT 47.190 58.120 49.920 58.310 ;
        RECT 50.230 58.730 57.800 58.930 ;
        RECT 47.190 58.110 47.680 58.120 ;
        RECT 45.390 57.780 45.710 57.830 ;
        RECT 15.800 57.630 16.110 57.720 ;
        RECT 15.200 57.460 16.110 57.630 ;
        RECT 15.800 57.390 16.110 57.460 ;
        RECT 16.890 57.640 17.200 57.730 ;
        RECT 16.890 57.470 18.000 57.640 ;
        RECT 16.890 57.400 17.200 57.470 ;
        RECT 40.560 56.960 40.820 57.760 ;
        RECT 45.390 57.580 47.020 57.780 ;
        RECT 45.390 57.570 45.710 57.580 ;
        RECT 42.560 56.960 42.900 57.020 ;
        RECT 38.290 56.600 38.750 56.920 ;
        RECT 40.460 56.740 42.900 56.960 ;
        RECT 50.230 56.770 50.430 58.730 ;
        RECT 57.480 58.700 57.800 58.730 ;
        RECT 57.480 58.690 57.790 58.700 ;
        RECT 58.540 58.450 58.860 58.490 ;
        RECT 47.480 56.760 50.430 56.770 ;
        RECT 46.790 56.430 46.900 56.630 ;
        RECT 47.190 56.570 50.430 56.760 ;
        RECT 50.780 58.250 58.940 58.450 ;
        RECT 47.190 56.560 47.690 56.570 ;
        RECT 45.390 56.230 45.710 56.280 ;
        RECT 40.560 55.410 40.820 56.210 ;
        RECT 45.390 56.030 47.020 56.230 ;
        RECT 45.390 56.020 45.710 56.030 ;
        RECT 42.560 55.410 42.900 55.470 ;
        RECT 38.290 55.050 38.750 55.370 ;
        RECT 40.460 55.190 42.900 55.410 ;
        RECT 50.780 55.220 50.980 58.250 ;
        RECT 58.540 58.210 58.860 58.250 ;
        RECT 47.490 55.210 50.980 55.220 ;
        RECT 47.190 55.020 50.980 55.210 ;
        RECT 53.930 56.450 54.220 56.630 ;
        RECT 47.190 55.010 47.650 55.020 ;
        RECT 53.930 53.190 54.110 56.450 ;
        RECT 84.130 55.040 84.210 55.220 ;
        RECT 78.280 54.020 78.880 54.580 ;
        RECT 81.880 54.410 87.110 54.640 ;
        RECT 82.350 54.170 82.660 54.310 ;
        RECT 80.180 54.160 82.660 54.170 ;
        RECT 80.180 54.010 91.700 54.160 ;
        RECT 80.180 53.990 82.660 54.010 ;
        RECT 82.350 53.980 82.660 53.990 ;
        RECT 81.890 53.590 87.110 53.810 ;
        RECT 53.100 53.010 54.110 53.190 ;
        RECT 59.350 53.380 59.670 53.430 ;
        RECT 61.760 53.380 62.080 53.400 ;
        RECT 59.350 53.240 62.080 53.380 ;
        RECT 59.350 53.190 63.780 53.240 ;
        RECT 59.350 53.110 59.670 53.190 ;
        RECT 61.760 53.140 63.780 53.190 ;
        RECT 61.800 53.070 63.780 53.140 ;
        RECT 63.260 53.060 63.780 53.070 ;
        RECT 82.350 53.010 82.660 53.020 ;
        RECT 47.490 52.800 47.790 52.830 ;
        RECT 47.490 52.790 47.880 52.800 ;
        RECT 38.290 52.430 38.750 52.750 ;
        RECT 40.460 52.390 42.900 52.610 ;
        RECT 47.190 52.590 47.880 52.790 ;
        RECT 58.110 52.670 58.590 52.900 ;
        RECT 80.180 52.830 91.710 53.010 ;
        RECT 82.350 52.690 82.660 52.830 ;
        RECT 58.250 52.600 58.590 52.670 ;
        RECT 40.560 51.590 40.820 52.390 ;
        RECT 42.560 52.330 42.900 52.390 ;
        RECT 82.200 51.990 82.510 52.060 ;
        RECT 80.180 51.980 82.510 51.990 ;
        RECT 45.390 51.770 45.710 51.780 ;
        RECT 45.390 51.570 47.020 51.770 ;
        RECT 45.390 51.520 45.710 51.570 ;
        RECT 47.460 51.480 47.790 51.680 ;
        RECT 53.490 51.560 54.220 51.740 ;
        RECT 58.250 51.730 58.590 51.800 ;
        RECT 80.180 51.770 91.710 51.980 ;
        RECT 81.490 51.760 91.710 51.770 ;
        RECT 82.200 51.730 82.510 51.760 ;
        RECT 38.290 50.880 38.750 51.200 ;
        RECT 46.790 51.170 46.900 51.370 ;
        RECT 47.460 51.260 47.640 51.480 ;
        RECT 53.490 51.350 53.670 51.560 ;
        RECT 58.110 51.500 58.590 51.730 ;
        RECT 47.440 51.240 47.640 51.260 ;
        RECT 40.460 50.840 42.900 51.060 ;
        RECT 47.190 51.040 47.640 51.240 ;
        RECT 53.100 51.170 53.670 51.350 ;
        RECT 82.660 51.130 87.110 51.290 ;
        RECT 82.630 51.090 87.110 51.130 ;
        RECT 40.560 50.040 40.820 50.840 ;
        RECT 42.560 50.780 42.900 50.840 ;
        RECT 53.590 50.410 54.140 50.590 ;
        RECT 77.220 50.550 77.780 51.090 ;
        RECT 82.630 51.010 82.860 51.090 ;
        RECT 81.250 50.790 91.710 51.010 ;
        RECT 81.250 50.650 81.570 50.790 ;
        RECT 59.350 50.450 59.670 50.500 ;
        RECT 61.760 50.450 62.080 50.470 ;
        RECT 45.390 50.220 45.710 50.230 ;
        RECT 45.390 50.020 47.020 50.220 ;
        RECT 53.590 50.200 53.770 50.410 ;
        RECT 53.100 50.020 53.770 50.200 ;
        RECT 59.350 50.260 62.080 50.450 ;
        RECT 81.270 50.310 81.530 50.650 ;
        RECT 59.350 50.180 59.670 50.260 ;
        RECT 61.760 50.250 62.080 50.260 ;
        RECT 61.760 50.210 63.780 50.250 ;
        RECT 61.870 50.090 63.780 50.210 ;
        RECT 62.590 50.070 63.780 50.090 ;
        RECT 81.250 50.050 81.570 50.310 ;
        RECT 45.390 49.970 45.710 50.020 ;
        RECT 47.440 49.850 47.790 49.920 ;
        RECT 38.290 49.330 38.750 49.650 ;
        RECT 46.790 49.620 46.900 49.820 ;
        RECT 47.440 49.690 47.830 49.850 ;
        RECT 58.110 49.740 58.590 49.970 ;
        RECT 47.250 49.620 47.830 49.690 ;
        RECT 58.250 49.670 58.590 49.740 ;
        RECT 40.460 49.290 42.900 49.510 ;
        RECT 47.250 49.490 47.640 49.620 ;
        RECT 40.560 48.490 40.820 49.290 ;
        RECT 42.560 49.230 42.900 49.290 ;
        RECT 82.200 49.230 82.510 49.300 ;
        RECT 82.630 49.230 82.860 50.790 ;
        RECT 84.130 50.170 84.210 50.350 ;
        RECT 80.180 49.020 91.710 49.230 ;
        RECT 81.490 49.010 91.710 49.020 ;
        RECT 82.200 48.970 82.510 49.010 ;
        RECT 58.250 48.800 58.590 48.870 ;
        RECT 45.390 48.670 45.710 48.680 ;
        RECT 45.390 48.470 47.020 48.670 ;
        RECT 47.530 48.540 47.790 48.750 ;
        RECT 58.110 48.570 58.590 48.800 ;
        RECT 82.630 48.610 82.860 49.010 ;
        RECT 45.390 48.420 45.710 48.470 ;
        RECT 38.290 47.780 38.750 48.100 ;
        RECT 46.790 48.070 46.900 48.270 ;
        RECT 47.530 48.140 47.730 48.540 ;
        RECT 62.530 48.380 63.780 48.390 ;
        RECT 53.100 48.160 53.870 48.340 ;
        RECT 40.460 47.740 42.900 47.960 ;
        RECT 47.390 47.940 47.730 48.140 ;
        RECT 47.530 47.930 47.730 47.940 ;
        RECT 38.100 47.380 38.190 47.700 ;
        RECT 40.560 46.940 40.820 47.740 ;
        RECT 42.560 47.680 42.900 47.740 ;
        RECT 45.390 47.120 45.710 47.130 ;
        RECT 45.390 46.920 47.020 47.120 ;
        RECT 45.390 46.870 45.710 46.920 ;
        RECT 46.790 46.520 46.900 46.720 ;
        RECT 53.690 45.720 53.870 48.160 ;
        RECT 59.350 48.280 59.670 48.360 ;
        RECT 61.840 48.330 63.780 48.380 ;
        RECT 61.760 48.280 63.780 48.330 ;
        RECT 59.350 48.220 63.780 48.280 ;
        RECT 59.350 48.090 62.080 48.220 ;
        RECT 62.530 48.210 63.780 48.220 ;
        RECT 59.350 48.040 59.670 48.090 ;
        RECT 61.760 48.070 62.080 48.090 ;
        RECT 78.260 48.000 78.880 48.530 ;
        RECT 81.880 48.380 82.860 48.610 ;
        RECT 83.470 48.480 87.110 48.680 ;
        RECT 82.350 48.140 82.660 48.280 ;
        RECT 80.180 48.130 82.660 48.140 ;
        RECT 83.470 48.130 83.670 48.480 ;
        RECT 80.180 47.980 91.710 48.130 ;
        RECT 80.180 47.960 82.660 47.980 ;
        RECT 82.350 47.950 82.660 47.960 ;
        RECT 83.470 47.780 83.670 47.980 ;
        RECT 81.890 47.630 83.670 47.780 ;
        RECT 81.890 47.560 83.640 47.630 ;
        RECT 67.660 47.100 67.970 47.240 ;
        RECT 88.430 47.100 88.740 47.240 ;
        RECT 109.310 47.210 109.620 47.260 ;
        RECT 111.610 47.210 111.920 47.230 ;
        RECT 65.500 46.920 75.570 47.100 ;
        RECT 80.830 46.920 90.900 47.100 ;
        RECT 93.440 46.970 102.450 47.190 ;
        RECT 108.100 46.990 108.410 47.030 ;
        RECT 67.660 46.910 67.970 46.920 ;
        RECT 88.430 46.910 88.740 46.920 ;
        RECT 67.660 46.670 67.970 46.690 ;
        RECT 88.430 46.670 88.740 46.690 ;
        RECT 65.500 46.490 75.570 46.670 ;
        RECT 80.830 46.490 90.900 46.670 ;
        RECT 67.660 46.360 67.970 46.490 ;
        RECT 88.430 46.360 88.740 46.490 ;
        RECT 53.690 45.540 54.230 45.720 ;
        RECT 67.660 45.670 67.970 45.800 ;
        RECT 88.430 45.670 88.740 45.800 ;
        RECT 65.500 45.490 75.580 45.670 ;
        RECT 80.820 45.490 90.900 45.670 ;
        RECT 67.660 45.470 67.970 45.490 ;
        RECT 88.430 45.470 88.740 45.490 ;
        RECT 67.660 45.240 67.970 45.250 ;
        RECT 88.430 45.240 88.740 45.250 ;
        RECT 65.500 45.060 75.580 45.240 ;
        RECT 80.820 45.060 90.900 45.240 ;
        RECT 93.490 45.190 99.150 45.410 ;
        RECT 67.660 44.920 67.970 45.060 ;
        RECT 88.430 44.920 88.740 45.060 ;
        RECT 92.990 44.890 93.470 44.900 ;
        RECT 92.990 44.650 93.880 44.890 ;
        RECT 98.930 44.860 99.150 45.190 ;
        RECT 102.230 45.360 102.450 46.970 ;
        RECT 107.780 46.980 108.440 46.990 ;
        RECT 109.310 46.980 112.230 47.210 ;
        RECT 107.780 46.750 108.880 46.980 ;
        RECT 109.310 46.930 109.620 46.980 ;
        RECT 111.610 46.900 111.920 46.980 ;
        RECT 108.100 46.700 108.410 46.750 ;
        RECT 109.310 46.380 109.620 46.440 ;
        RECT 111.600 46.380 111.910 46.510 ;
        RECT 109.310 46.160 112.230 46.380 ;
        RECT 109.310 46.110 109.620 46.160 ;
        RECT 102.230 45.140 105.080 45.360 ;
        RECT 109.260 44.910 109.570 44.950 ;
        RECT 103.300 44.860 109.570 44.910 ;
        RECT 98.930 44.700 109.570 44.860 ;
        RECT 98.930 44.640 103.690 44.700 ;
        RECT 109.260 44.620 109.570 44.700 ;
        RECT 109.310 44.220 109.620 44.300 ;
        RECT 111.520 44.220 111.830 44.260 ;
        RECT 109.310 43.990 112.020 44.220 ;
        RECT 109.310 43.970 109.620 43.990 ;
        RECT 111.520 43.930 111.830 43.990 ;
        RECT 59.350 43.310 59.670 43.360 ;
        RECT 61.760 43.310 62.080 43.330 ;
        RECT 53.860 43.120 55.640 43.240 ;
        RECT 53.270 43.060 55.640 43.120 ;
        RECT 59.350 43.170 62.080 43.310 ;
        RECT 59.350 43.120 63.780 43.170 ;
        RECT 53.270 42.940 54.110 43.060 ;
        RECT 59.350 43.040 59.670 43.120 ;
        RECT 61.760 43.070 63.780 43.120 ;
        RECT 68.140 43.100 68.280 43.290 ;
        RECT 88.170 43.100 88.260 43.280 ;
        RECT 61.800 43.000 63.780 43.070 ;
        RECT 63.260 42.990 63.780 43.000 ;
        RECT 47.530 42.760 47.780 42.780 ;
        RECT 47.530 42.660 47.790 42.760 ;
        RECT 38.290 42.300 38.750 42.620 ;
        RECT 40.460 42.260 42.900 42.480 ;
        RECT 47.190 42.460 47.790 42.660 ;
        RECT 58.110 42.600 58.590 42.830 ;
        RECT 67.660 42.680 67.970 42.800 ;
        RECT 68.140 42.680 68.280 42.860 ;
        RECT 75.400 42.680 75.960 42.810 ;
        RECT 88.170 42.680 88.260 42.850 ;
        RECT 88.430 42.680 88.740 42.800 ;
        RECT 67.660 42.670 75.960 42.680 ;
        RECT 58.250 42.530 58.590 42.600 ;
        RECT 65.500 42.630 75.960 42.670 ;
        RECT 80.840 42.670 88.740 42.680 ;
        RECT 65.500 42.510 75.560 42.630 ;
        RECT 80.840 42.510 90.900 42.670 ;
        RECT 65.500 42.490 68.060 42.510 ;
        RECT 67.660 42.470 67.970 42.490 ;
        RECT 73.240 42.420 74.780 42.510 ;
        RECT 81.620 42.420 83.160 42.510 ;
        RECT 88.340 42.490 90.900 42.510 ;
        RECT 88.430 42.470 88.740 42.490 ;
        RECT 40.560 41.460 40.820 42.260 ;
        RECT 42.560 42.200 42.900 42.260 ;
        RECT 67.660 42.240 67.970 42.250 ;
        RECT 88.430 42.240 88.740 42.250 ;
        RECT 65.500 42.070 75.560 42.240 ;
        RECT 80.840 42.070 90.900 42.240 ;
        RECT 65.500 42.060 67.970 42.070 ;
        RECT 67.660 41.920 67.970 42.060 ;
        RECT 88.430 42.060 90.900 42.070 ;
        RECT 88.430 41.920 88.740 42.060 ;
        RECT 58.250 41.660 58.590 41.730 ;
        RECT 68.140 41.670 68.290 41.860 ;
        RECT 88.140 41.670 88.270 41.850 ;
        RECT 45.390 41.640 45.710 41.650 ;
        RECT 45.390 41.440 47.020 41.640 ;
        RECT 45.390 41.390 45.710 41.440 ;
        RECT 47.380 41.410 47.760 41.610 ;
        RECT 58.110 41.430 58.590 41.660 ;
        RECT 47.380 41.380 47.750 41.410 ;
        RECT 38.290 40.750 38.750 41.070 ;
        RECT 46.790 41.040 46.900 41.240 ;
        RECT 47.380 41.110 47.580 41.380 ;
        RECT 53.880 41.280 55.640 41.380 ;
        RECT 40.460 40.710 42.900 40.930 ;
        RECT 47.190 40.910 47.580 41.110 ;
        RECT 53.280 41.200 55.640 41.280 ;
        RECT 53.280 41.100 54.160 41.200 ;
        RECT 59.350 41.140 59.670 41.220 ;
        RECT 61.830 41.190 63.780 41.330 ;
        RECT 68.140 41.240 68.270 41.420 ;
        RECT 88.130 41.240 88.270 41.420 ;
        RECT 61.760 41.170 63.780 41.190 ;
        RECT 61.760 41.140 62.080 41.170 ;
        RECT 62.560 41.160 63.780 41.170 ;
        RECT 63.260 41.150 63.780 41.160 ;
        RECT 59.350 40.950 62.080 41.140 ;
        RECT 59.350 40.900 59.670 40.950 ;
        RECT 61.760 40.930 62.080 40.950 ;
        RECT 40.560 39.910 40.820 40.710 ;
        RECT 42.560 40.650 42.900 40.710 ;
        RECT 59.350 40.380 59.670 40.430 ;
        RECT 61.760 40.380 62.080 40.400 ;
        RECT 53.890 40.130 55.640 40.230 ;
        RECT 45.390 40.090 45.710 40.100 ;
        RECT 45.390 39.890 47.020 40.090 ;
        RECT 53.280 40.050 55.640 40.130 ;
        RECT 59.350 40.190 62.080 40.380 ;
        RECT 59.350 40.110 59.670 40.190 ;
        RECT 61.760 40.180 62.080 40.190 ;
        RECT 61.760 40.140 63.780 40.180 ;
        RECT 53.280 39.950 54.160 40.050 ;
        RECT 61.870 40.020 63.780 40.140 ;
        RECT 68.140 40.090 68.210 40.270 ;
        RECT 88.180 40.090 88.270 40.270 ;
        RECT 62.590 40.000 63.780 40.020 ;
        RECT 45.390 39.840 45.710 39.890 ;
        RECT 38.290 39.200 38.750 39.520 ;
        RECT 46.790 39.490 46.900 39.690 ;
        RECT 47.590 39.560 47.790 39.840 ;
        RECT 58.110 39.670 58.590 39.900 ;
        RECT 58.250 39.600 58.590 39.670 ;
        RECT 68.140 39.660 68.210 39.840 ;
        RECT 88.180 39.660 88.270 39.840 ;
        RECT 40.460 39.160 42.900 39.380 ;
        RECT 47.190 39.360 47.790 39.560 ;
        RECT 40.560 38.360 40.820 39.160 ;
        RECT 42.560 39.100 42.900 39.160 ;
        RECT 74.840 39.110 81.600 39.290 ;
        RECT 58.250 38.730 58.590 38.800 ;
        RECT 45.390 38.540 45.710 38.550 ;
        RECT 45.390 38.340 47.020 38.540 ;
        RECT 45.390 38.290 45.710 38.340 ;
        RECT 38.290 37.650 38.750 37.970 ;
        RECT 46.790 37.940 46.900 38.140 ;
        RECT 47.590 38.010 47.790 38.680 ;
        RECT 58.110 38.500 58.590 38.730 ;
        RECT 68.140 38.670 68.210 38.850 ;
        RECT 88.180 38.670 88.270 38.850 ;
        RECT 53.860 38.270 55.640 38.380 ;
        RECT 62.530 38.310 63.780 38.320 ;
        RECT 53.280 38.200 55.640 38.270 ;
        RECT 59.350 38.210 59.670 38.290 ;
        RECT 61.840 38.260 63.780 38.310 ;
        RECT 61.760 38.210 63.780 38.260 ;
        RECT 68.140 38.240 68.210 38.420 ;
        RECT 88.180 38.240 88.270 38.420 ;
        RECT 53.280 38.090 54.160 38.200 ;
        RECT 59.350 38.150 63.780 38.210 ;
        RECT 40.460 37.610 42.900 37.830 ;
        RECT 47.190 37.810 47.790 38.010 ;
        RECT 59.350 38.020 62.080 38.150 ;
        RECT 62.530 38.140 63.780 38.150 ;
        RECT 59.350 37.970 59.670 38.020 ;
        RECT 61.760 38.000 62.080 38.020 ;
        RECT 38.100 37.250 38.190 37.570 ;
        RECT 40.560 36.810 40.820 37.610 ;
        RECT 42.560 37.550 42.900 37.610 ;
        RECT 45.390 36.990 45.710 37.000 ;
        RECT 45.390 36.790 47.020 36.990 ;
        RECT 45.390 36.740 45.710 36.790 ;
        RECT 46.790 36.390 46.900 36.590 ;
        RECT 68.240 34.700 68.550 34.840 ;
        RECT 66.070 34.690 68.550 34.700 ;
        RECT 66.070 34.520 68.670 34.690 ;
        RECT 68.240 34.510 68.550 34.520 ;
        RECT 68.190 33.710 68.740 33.890 ;
        RECT 69.270 33.680 69.590 33.740 ;
        RECT 73.290 33.680 73.620 33.710 ;
        RECT 59.350 33.550 59.670 33.600 ;
        RECT 61.760 33.550 62.080 33.570 ;
        RECT 53.130 33.280 55.090 33.460 ;
        RECT 59.350 33.410 62.080 33.550 ;
        RECT 69.270 33.510 73.620 33.680 ;
        RECT 69.270 33.460 69.590 33.510 ;
        RECT 73.290 33.450 73.620 33.510 ;
        RECT 59.350 33.360 63.780 33.410 ;
        RECT 59.350 33.280 59.670 33.360 ;
        RECT 61.760 33.310 63.780 33.360 ;
        RECT 78.810 33.340 78.850 33.430 ;
        RECT 61.800 33.240 63.780 33.310 ;
        RECT 63.260 33.230 63.780 33.240 ;
        RECT 78.700 33.250 79.910 33.340 ;
        RECT 78.700 33.190 80.040 33.250 ;
        RECT 78.700 33.140 82.310 33.190 ;
        RECT 38.290 32.530 38.750 32.850 ;
        RECT 40.460 32.490 42.900 32.710 ;
        RECT 47.170 32.690 47.820 32.890 ;
        RECT 53.930 32.870 55.100 33.020 ;
        RECT 53.870 32.540 54.150 32.870 ;
        RECT 58.110 32.840 58.590 33.070 ;
        RECT 79.730 33.030 82.310 33.140 ;
        RECT 79.730 32.920 80.040 33.030 ;
        RECT 58.250 32.770 58.590 32.840 ;
        RECT 40.560 31.690 40.820 32.490 ;
        RECT 42.560 32.430 42.900 32.490 ;
        RECT 78.800 32.370 80.010 32.480 ;
        RECT 78.800 32.280 80.040 32.370 ;
        RECT 79.730 32.260 80.040 32.280 ;
        RECT 79.730 32.100 82.310 32.260 ;
        RECT 79.730 32.040 80.040 32.100 ;
        RECT 58.250 31.900 58.590 31.970 ;
        RECT 45.390 31.870 45.710 31.880 ;
        RECT 45.390 31.670 47.020 31.870 ;
        RECT 45.390 31.620 45.710 31.670 ;
        RECT 47.550 31.640 47.800 31.870 ;
        RECT 58.110 31.670 58.590 31.900 ;
        RECT 68.170 31.850 68.740 32.030 ;
        RECT 38.290 30.980 38.750 31.300 ;
        RECT 46.790 31.270 46.900 31.470 ;
        RECT 47.550 31.340 47.750 31.640 ;
        RECT 40.460 30.940 42.900 31.160 ;
        RECT 47.190 31.140 47.750 31.340 ;
        RECT 53.130 31.420 55.470 31.600 ;
        RECT 53.130 31.320 53.310 31.420 ;
        RECT 59.350 31.380 59.670 31.460 ;
        RECT 61.830 31.430 63.780 31.570 ;
        RECT 61.760 31.410 63.780 31.430 ;
        RECT 61.760 31.380 62.080 31.410 ;
        RECT 62.560 31.400 63.780 31.410 ;
        RECT 63.260 31.390 63.780 31.400 ;
        RECT 59.350 31.190 62.080 31.380 ;
        RECT 59.350 31.140 59.670 31.190 ;
        RECT 61.760 31.170 62.080 31.190 ;
        RECT 40.560 30.140 40.820 30.940 ;
        RECT 42.560 30.880 42.900 30.940 ;
        RECT 68.190 30.700 68.740 30.880 ;
        RECT 68.190 30.690 68.350 30.700 ;
        RECT 59.350 30.620 59.670 30.670 ;
        RECT 61.760 30.620 62.080 30.640 ;
        RECT 45.390 30.320 45.710 30.330 ;
        RECT 45.390 30.120 47.020 30.320 ;
        RECT 53.140 30.270 55.100 30.450 ;
        RECT 59.350 30.430 62.080 30.620 ;
        RECT 79.730 30.450 80.040 30.480 ;
        RECT 59.350 30.350 59.670 30.430 ;
        RECT 61.760 30.420 62.080 30.430 ;
        RECT 78.790 30.420 80.040 30.450 ;
        RECT 61.760 30.380 63.780 30.420 ;
        RECT 61.870 30.260 63.780 30.380 ;
        RECT 78.790 30.290 82.310 30.420 ;
        RECT 62.590 30.240 63.780 30.260 ;
        RECT 79.730 30.260 82.310 30.290 ;
        RECT 79.730 30.150 80.040 30.260 ;
        RECT 45.390 30.070 45.710 30.120 ;
        RECT 47.560 30.080 47.760 30.090 ;
        RECT 38.290 29.430 38.750 29.750 ;
        RECT 46.790 29.720 46.900 29.920 ;
        RECT 47.560 29.810 47.850 30.080 ;
        RECT 54.480 30.020 54.800 30.070 ;
        RECT 54.480 29.820 55.090 30.020 ;
        RECT 58.110 29.910 58.590 30.140 ;
        RECT 81.860 29.930 82.190 30.020 ;
        RECT 58.250 29.840 58.590 29.910 ;
        RECT 47.560 29.790 47.760 29.810 ;
        RECT 40.460 29.390 42.900 29.610 ;
        RECT 47.150 29.590 47.760 29.790 ;
        RECT 54.480 29.750 54.940 29.820 ;
        RECT 75.510 29.760 82.190 29.930 ;
        RECT 81.860 29.730 82.190 29.760 ;
        RECT 79.730 29.490 80.040 29.600 ;
        RECT 79.730 29.480 82.310 29.490 ;
        RECT 17.290 28.340 17.900 28.670 ;
        RECT 40.560 28.590 40.820 29.390 ;
        RECT 42.560 29.330 42.900 29.390 ;
        RECT 78.800 29.330 82.310 29.480 ;
        RECT 78.800 29.300 80.040 29.330 ;
        RECT 79.730 29.270 80.040 29.300 ;
        RECT 58.250 28.970 58.590 29.040 ;
        RECT 47.540 28.930 47.840 28.970 ;
        RECT 45.390 28.770 45.710 28.780 ;
        RECT 45.390 28.570 47.020 28.770 ;
        RECT 47.530 28.690 47.840 28.930 ;
        RECT 58.110 28.740 58.590 28.970 ;
        RECT 45.390 28.520 45.710 28.570 ;
        RECT 17.300 27.850 17.900 28.340 ;
        RECT 38.290 27.880 38.750 28.200 ;
        RECT 46.790 28.170 46.900 28.370 ;
        RECT 47.530 28.240 47.730 28.690 ;
        RECT 53.140 28.420 55.430 28.600 ;
        RECT 62.530 28.550 63.780 28.560 ;
        RECT 59.350 28.450 59.670 28.530 ;
        RECT 61.840 28.500 63.780 28.550 ;
        RECT 61.760 28.450 63.780 28.500 ;
        RECT 47.180 28.040 47.730 28.240 ;
        RECT 59.350 28.390 63.780 28.450 ;
        RECT 59.350 28.260 62.080 28.390 ;
        RECT 62.530 28.380 63.780 28.390 ;
        RECT 59.350 28.210 59.670 28.260 ;
        RECT 61.760 28.240 62.080 28.260 ;
        RECT 38.100 27.480 38.190 27.800 ;
        RECT 47.270 27.650 47.590 27.700 ;
        RECT 53.880 27.650 54.200 27.750 ;
        RECT 47.270 27.490 54.200 27.650 ;
        RECT 47.270 27.440 47.590 27.490 ;
        RECT 53.880 27.470 54.200 27.490 ;
        RECT 54.910 27.650 55.230 27.740 ;
        RECT 65.530 27.650 65.940 27.760 ;
        RECT 54.910 27.490 65.940 27.650 ;
        RECT 54.910 27.460 55.230 27.490 ;
        RECT 54.470 27.410 54.750 27.420 ;
        RECT 54.450 27.320 54.770 27.410 ;
        RECT 65.530 27.390 65.940 27.490 ;
        RECT 56.690 27.320 57.010 27.350 ;
        RECT 54.420 27.160 57.010 27.320 ;
        RECT 54.450 27.150 54.770 27.160 ;
        RECT 54.470 27.140 54.750 27.150 ;
        RECT 56.690 27.090 57.010 27.160 ;
        RECT 56.710 27.080 56.990 27.090 ;
        RECT 55.490 25.810 55.870 26.200 ;
        RECT 71.570 26.190 71.870 26.210 ;
        RECT 56.640 25.770 57.040 26.110 ;
        RECT 65.230 25.610 65.890 25.970 ;
        RECT 70.860 25.850 71.880 26.190 ;
        RECT 71.570 25.830 71.880 25.850 ;
        RECT 46.790 24.770 47.170 25.150 ;
        RECT 66.980 24.890 67.430 25.320 ;
        RECT 115.730 21.110 115.740 21.120 ;
        RECT 16.580 20.780 17.190 21.110 ;
        RECT 16.590 20.290 17.190 20.780 ;
        RECT 46.810 16.710 47.410 17.200 ;
        RECT 55.270 16.710 55.870 17.200 ;
        RECT 46.810 16.380 47.420 16.710 ;
        RECT 55.260 16.380 55.870 16.710 ;
        RECT 102.620 13.810 102.910 13.870 ;
        RECT 102.450 13.500 102.910 13.810 ;
        RECT 102.620 13.460 102.910 13.500 ;
        RECT 102.630 13.140 102.910 13.460 ;
        RECT 102.450 12.830 102.910 13.140 ;
        RECT 102.630 12.710 102.910 12.830 ;
        RECT 0.590 7.350 1.860 9.230 ;
        RECT 0.660 2.600 1.930 4.480 ;
        RECT 99.360 0.270 99.680 0.590 ;
        RECT 100.300 0.270 100.620 0.590 ;
      LAYER via2 ;
        RECT 78.410 54.130 78.750 54.470 ;
        RECT 77.340 50.650 77.670 51.000 ;
        RECT 78.430 48.080 78.770 48.440 ;
  END
END sky130_hilas_TopLevelTextStructure

MACRO sky130_hilas_pFETLarge
  CLASS CORE ;
  FOREIGN sky130_hilas_pFETLarge ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.610 BY 6.100 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA 5.457400 ;
    ANTENNADIFFAREA 1.079500 ;
    PORT
      LAYER met2 ;
        RECT 0.750 0.340 1.350 0.830 ;
        RECT 0.750 0.010 1.360 0.340 ;
    END
  END GATE
  PIN SOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 2.724600 ;
    PORT
      LAYER met2 ;
        RECT 1.080 5.600 4.140 5.610 ;
        RECT 0.990 5.270 4.140 5.600 ;
        RECT 0.990 2.820 1.310 5.270 ;
        RECT 3.810 5.260 4.120 5.270 ;
        RECT 0.990 2.490 4.150 2.820 ;
        RECT 0.990 1.450 1.310 2.490 ;
        RECT 0.990 1.130 4.150 1.450 ;
        RECT 1.610 1.120 1.920 1.130 ;
        RECT 2.710 1.120 3.020 1.130 ;
        RECT 3.810 1.120 4.120 1.130 ;
    END
  END SOURCE
  PIN DRAIN
    USE ANALOG ;
    ANTENNADIFFAREA 1.386200 ;
    PORT
      LAYER met2 ;
        RECT 2.170 4.890 2.480 4.920 ;
        RECT 3.260 4.890 3.570 4.900 ;
        RECT 2.170 4.590 5.120 4.890 ;
        RECT 3.260 4.570 3.570 4.590 ;
        RECT 4.370 4.550 5.120 4.590 ;
        RECT 4.740 4.420 5.120 4.550 ;
        RECT 4.770 3.550 5.120 4.420 ;
        RECT 2.170 3.220 5.120 3.550 ;
        RECT 4.770 0.780 5.120 3.220 ;
        RECT 2.180 0.770 5.120 0.780 ;
        RECT 2.170 0.460 5.120 0.770 ;
        RECT 2.170 0.450 4.890 0.460 ;
        RECT 2.170 0.440 2.480 0.450 ;
        RECT 3.260 0.440 3.570 0.450 ;
    END
  END DRAIN
  PIN WELL
    USE ANALOG ;
    ANTENNADIFFAREA 0.213200 ;
    PORT
      LAYER nwell ;
        RECT 4.770 0.180 5.390 5.880 ;
      LAYER met1 ;
        RECT 4.890 5.790 5.150 5.990 ;
        RECT 4.890 4.980 5.200 5.790 ;
        RECT 4.890 0.000 5.150 4.980 ;
    END
  END WELL
  OBS
      LAYER nwell ;
        RECT 0.000 0.400 3.390 6.100 ;
        RECT 4.390 3.060 4.400 3.100 ;
      LAYER li1 ;
        RECT 0.240 3.380 0.410 5.870 ;
        RECT 0.790 3.370 0.960 5.870 ;
        RECT 1.340 3.370 1.510 5.870 ;
        RECT 1.890 5.560 2.060 5.870 ;
        RECT 1.630 5.300 2.060 5.560 ;
        RECT 1.890 3.370 2.060 5.300 ;
        RECT 2.440 4.880 2.610 5.870 ;
        RECT 2.990 5.560 3.160 5.870 ;
        RECT 2.720 5.300 3.160 5.560 ;
        RECT 2.180 4.620 2.610 4.880 ;
        RECT 2.440 3.510 2.610 4.620 ;
        RECT 2.180 3.370 2.610 3.510 ;
        RECT 2.990 3.370 3.160 5.300 ;
        RECT 3.820 5.510 4.140 5.550 ;
        RECT 3.820 5.320 4.150 5.510 ;
        RECT 3.820 5.290 4.140 5.320 ;
        RECT 5.000 4.920 5.170 5.680 ;
        RECT 3.270 4.820 3.590 4.860 ;
        RECT 3.270 4.630 3.600 4.820 ;
        RECT 4.380 4.810 4.700 4.850 ;
        RECT 3.270 4.600 3.590 4.630 ;
        RECT 4.380 4.620 4.710 4.810 ;
        RECT 4.380 4.590 4.700 4.620 ;
        RECT 3.270 3.470 3.590 3.510 ;
        RECT 4.370 3.470 4.690 3.510 ;
        RECT 2.180 3.280 2.510 3.370 ;
        RECT 3.270 3.280 3.600 3.470 ;
        RECT 4.370 3.280 4.700 3.470 ;
        RECT 2.180 3.250 2.500 3.280 ;
        RECT 3.270 3.250 3.590 3.280 ;
        RECT 4.370 3.250 4.690 3.280 ;
        RECT 1.710 3.160 1.870 3.190 ;
        RECT 0.240 0.550 0.410 3.040 ;
        RECT 0.790 1.020 0.960 3.040 ;
        RECT 1.340 1.020 1.510 3.040 ;
        RECT 1.710 2.820 1.880 3.160 ;
        RECT 2.260 3.150 2.420 3.190 ;
        RECT 1.710 2.810 1.870 2.820 ;
        RECT 1.890 2.780 2.060 3.040 ;
        RECT 2.260 2.820 2.430 3.150 ;
        RECT 2.260 2.810 2.420 2.820 ;
        RECT 1.620 2.520 2.060 2.780 ;
        RECT 1.890 1.410 2.060 2.520 ;
        RECT 1.620 1.150 2.060 1.410 ;
        RECT 0.790 0.540 1.510 1.020 ;
        RECT 1.890 0.540 2.060 1.150 ;
        RECT 2.440 0.730 2.610 3.040 ;
        RECT 2.810 2.820 2.980 3.220 ;
        RECT 3.360 3.150 3.520 3.190 ;
        RECT 3.910 3.150 4.070 3.190 ;
        RECT 4.460 3.170 4.620 3.190 ;
        RECT 2.810 2.810 2.970 2.820 ;
        RECT 2.990 2.780 3.160 3.040 ;
        RECT 3.360 2.820 3.530 3.150 ;
        RECT 3.910 2.820 4.080 3.150 ;
        RECT 4.460 2.820 4.630 3.170 ;
        RECT 3.360 2.810 3.520 2.820 ;
        RECT 3.910 2.810 4.070 2.820 ;
        RECT 4.460 2.810 4.620 2.820 ;
        RECT 2.720 2.520 3.160 2.780 ;
        RECT 3.820 2.740 4.140 2.780 ;
        RECT 3.820 2.550 4.150 2.740 ;
        RECT 3.820 2.520 4.140 2.550 ;
        RECT 2.990 1.410 3.160 2.520 ;
        RECT 2.720 1.150 3.160 1.410 ;
        RECT 3.820 1.370 4.140 1.410 ;
        RECT 3.820 1.180 4.150 1.370 ;
        RECT 3.820 1.150 4.140 1.180 ;
        RECT 2.180 0.540 2.610 0.730 ;
        RECT 2.990 0.540 3.160 1.150 ;
        RECT 3.270 0.690 3.590 0.730 ;
        RECT 4.370 0.700 4.690 0.740 ;
        RECT 0.950 0.010 1.460 0.540 ;
        RECT 2.180 0.500 2.510 0.540 ;
        RECT 3.270 0.500 3.600 0.690 ;
        RECT 4.370 0.510 4.700 0.700 ;
        RECT 2.180 0.470 2.500 0.500 ;
        RECT 3.270 0.470 3.590 0.500 ;
        RECT 4.370 0.480 4.690 0.510 ;
      LAYER mcon ;
        RECT 1.690 5.340 1.860 5.510 ;
        RECT 2.780 5.340 2.950 5.510 ;
        RECT 2.240 4.660 2.410 4.830 ;
        RECT 2.240 3.290 2.410 3.460 ;
        RECT 5.000 5.510 5.170 5.680 ;
        RECT 3.880 5.330 4.050 5.500 ;
        RECT 5.000 5.170 5.170 5.340 ;
        RECT 3.330 4.640 3.500 4.810 ;
        RECT 4.440 4.630 4.610 4.800 ;
        RECT 3.330 3.290 3.500 3.460 ;
        RECT 4.430 3.290 4.600 3.460 ;
        RECT 1.680 2.560 1.850 2.730 ;
        RECT 1.680 1.190 1.850 1.360 ;
        RECT 1.110 0.550 1.280 0.720 ;
        RECT 2.780 2.560 2.950 2.730 ;
        RECT 3.880 2.560 4.050 2.730 ;
        RECT 2.780 1.190 2.950 1.360 ;
        RECT 3.880 1.190 4.050 1.360 ;
        RECT 2.240 0.510 2.410 0.680 ;
        RECT 3.330 0.510 3.500 0.680 ;
        RECT 4.430 0.520 4.600 0.690 ;
        RECT 1.120 0.080 1.290 0.250 ;
      LAYER met1 ;
        RECT 1.620 5.270 1.940 5.590 ;
        RECT 2.710 5.270 3.030 5.590 ;
        RECT 3.810 5.260 4.130 5.580 ;
        RECT 2.170 4.590 2.490 4.910 ;
        RECT 3.260 4.570 3.580 4.890 ;
        RECT 4.370 4.560 4.690 4.880 ;
        RECT 2.170 3.220 2.490 3.540 ;
        RECT 3.260 3.220 3.580 3.540 ;
        RECT 4.360 3.220 4.680 3.540 ;
        RECT 1.610 2.490 1.930 2.810 ;
        RECT 2.710 2.490 3.030 2.810 ;
        RECT 3.810 2.490 4.130 2.810 ;
        RECT 1.610 1.120 1.930 1.440 ;
        RECT 2.710 1.120 3.030 1.440 ;
        RECT 3.810 1.120 4.130 1.440 ;
        RECT 1.040 0.480 1.360 0.800 ;
        RECT 2.170 0.440 2.490 0.760 ;
        RECT 3.260 0.440 3.580 0.760 ;
        RECT 4.360 0.450 4.680 0.770 ;
        RECT 1.050 0.010 1.370 0.330 ;
      LAYER via ;
        RECT 1.650 5.300 1.910 5.560 ;
        RECT 2.740 5.300 3.000 5.560 ;
        RECT 3.840 5.290 4.100 5.550 ;
        RECT 2.200 4.620 2.460 4.880 ;
        RECT 3.290 4.600 3.550 4.860 ;
        RECT 4.400 4.590 4.660 4.850 ;
        RECT 2.200 3.250 2.460 3.510 ;
        RECT 3.290 3.250 3.550 3.510 ;
        RECT 4.390 3.250 4.650 3.510 ;
        RECT 1.640 2.520 1.900 2.780 ;
        RECT 2.740 2.520 3.000 2.780 ;
        RECT 3.840 2.520 4.100 2.780 ;
        RECT 1.640 1.150 1.900 1.410 ;
        RECT 2.740 1.150 3.000 1.410 ;
        RECT 3.840 1.150 4.100 1.410 ;
        RECT 1.070 0.510 1.330 0.770 ;
        RECT 2.200 0.470 2.460 0.730 ;
        RECT 3.290 0.470 3.550 0.730 ;
        RECT 4.390 0.480 4.650 0.740 ;
        RECT 1.080 0.040 1.340 0.300 ;
  END
END sky130_hilas_pFETLarge

MACRO sky130_hilas_VinjInv2
  CLASS CORE ;
  FOREIGN sky130_hilas_VinjInv2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.610 BY 1.640 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 0.000 0.000 1.980 1.640 ;
      LAYER li1 ;
        RECT 0.620 1.210 0.790 1.350 ;
        RECT 0.620 1.040 0.810 1.210 ;
        RECT 0.620 0.940 0.790 1.040 ;
        RECT 0.190 0.560 0.360 0.660 ;
        RECT 0.170 0.390 0.360 0.560 ;
        RECT 0.190 0.330 0.360 0.390 ;
        RECT 0.610 0.600 0.780 0.660 ;
        RECT 0.610 0.330 0.860 0.600 ;
        RECT 1.350 0.580 1.600 0.660 ;
        RECT 1.350 0.410 2.650 0.580 ;
        RECT 3.210 0.570 3.380 1.200 ;
        RECT 0.620 0.310 0.860 0.330 ;
        RECT 1.430 0.320 1.600 0.410 ;
        RECT 3.130 0.400 3.460 0.570 ;
      LAYER mcon ;
        RECT 0.640 1.040 0.810 1.210 ;
        RECT 3.210 0.680 3.380 0.850 ;
        RECT 0.650 0.360 0.820 0.530 ;
        RECT 1.990 0.410 2.160 0.580 ;
      LAYER met1 ;
        RECT 0.610 1.260 0.830 1.600 ;
        RECT 0.610 1.000 0.840 1.260 ;
        RECT 0.080 0.320 0.390 0.670 ;
        RECT 0.610 0.600 0.830 1.000 ;
        RECT 0.610 0.290 0.860 0.600 ;
        RECT 1.910 0.360 2.230 0.620 ;
        RECT 0.610 0.090 0.830 0.290 ;
        RECT 3.180 0.090 3.410 1.600 ;
      LAYER via ;
        RECT 0.110 0.350 0.370 0.610 ;
        RECT 1.940 0.360 2.200 0.620 ;
      LAYER met2 ;
        RECT 0.000 1.030 3.610 1.210 ;
        RECT 0.080 0.510 0.400 0.610 ;
        RECT 0.070 0.350 0.400 0.510 ;
        RECT 1.910 0.540 2.230 0.620 ;
        RECT 1.910 0.360 3.610 0.540 ;
  END
END sky130_hilas_VinjInv2

MACRO sky130_hilas_capacitorSize03
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize03 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.790 BY 5.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 4.960 2.630 5.620 3.290 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 2.570 4.530 3.020 4.540 ;
        RECT 2.550 4.040 3.070 4.530 ;
        RECT 0.110 3.190 0.770 3.250 ;
        RECT 2.580 3.200 3.020 4.040 ;
        RECT 1.160 3.190 2.170 3.200 ;
        RECT 2.570 3.190 3.030 3.200 ;
        RECT 0.110 2.690 3.030 3.190 ;
        RECT 0.110 2.680 1.520 2.690 ;
        RECT 0.110 2.590 0.770 2.680 ;
        RECT 2.570 2.030 3.030 2.690 ;
        RECT 2.570 1.520 3.050 2.030 ;
        RECT 2.550 1.030 3.070 1.520 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 0.000 5.270 5.780 5.450 ;
        RECT 0.000 4.840 5.780 5.020 ;
        RECT 0.030 3.840 5.780 4.020 ;
        RECT 0.030 3.410 5.780 3.590 ;
        RECT 0.240 3.070 0.610 3.130 ;
        RECT 0.020 2.790 0.610 3.070 ;
        RECT 0.240 2.730 0.610 2.790 ;
        RECT 5.090 3.110 5.460 3.170 ;
        RECT 5.090 2.830 5.790 3.110 ;
        RECT 5.090 2.770 5.460 2.830 ;
        RECT 0.030 2.260 5.780 2.430 ;
        RECT 0.030 1.840 5.780 2.010 ;
        RECT 0.030 0.860 5.780 1.030 ;
        RECT 0.030 0.420 5.780 0.590 ;
      LAYER via2 ;
        RECT 0.290 2.790 0.570 3.070 ;
        RECT 5.140 2.830 5.420 3.110 ;
      LAYER met3 ;
        RECT 1.450 3.320 4.290 5.870 ;
        RECT 0.020 2.530 0.810 3.280 ;
        RECT 1.450 2.570 5.660 3.320 ;
        RECT 1.450 0.000 4.290 2.570 ;
      LAYER via3 ;
        RECT 0.210 2.680 0.640 3.160 ;
        RECT 5.060 2.720 5.490 3.200 ;
  END
END sky130_hilas_capacitorSize03

MACRO sky130_hilas_swc4x1BiasCell
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x1BiasCell ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.110 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN ROW1
    USE ANALOG ;
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 7.630 5.120 7.940 5.140 ;
        RECT 0.020 4.940 10.100 5.120 ;
        RECT 0.020 4.930 0.170 4.940 ;
        RECT 7.630 4.810 7.940 4.940 ;
    END
  END ROW1
  PIN ROW2
    USE ANALOG ;
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 0.000 4.120 0.140 4.140 ;
        RECT 7.630 4.120 7.940 4.250 ;
        RECT 0.000 3.940 10.110 4.120 ;
        RECT 7.630 3.920 7.940 3.940 ;
    END
  END ROW2
  PIN ROW3
    USE ANALOG ;
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 7.630 2.110 7.940 2.130 ;
        RECT 0.030 1.950 10.100 2.110 ;
        RECT 0.040 1.940 10.100 1.950 ;
        RECT 7.540 1.930 10.100 1.940 ;
        RECT 7.630 1.800 7.940 1.930 ;
    END
  END ROW3
  PIN ROW4
    USE ANALOG ;
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 7.630 1.130 7.940 1.250 ;
        RECT 0.030 1.120 7.940 1.130 ;
        RECT 0.030 0.960 10.100 1.120 ;
        RECT 0.820 0.870 2.360 0.960 ;
        RECT 7.540 0.940 10.100 0.960 ;
        RECT 7.630 0.920 7.940 0.940 ;
    END
  END ROW4
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 1.978000 ;
    PORT
      LAYER nwell ;
        RECT 0.030 5.420 1.760 6.050 ;
        RECT 0.020 2.350 1.760 5.420 ;
        RECT 0.030 0.000 1.760 2.350 ;
      LAYER met1 ;
        RECT 0.380 0.000 0.780 6.050 ;
    END
  END VTUN
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 2.743300 ;
    PORT
      LAYER nwell ;
        RECT 3.780 0.000 6.010 6.050 ;
      LAYER met1 ;
        RECT 4.430 4.130 4.810 6.050 ;
        RECT 4.420 2.270 4.810 4.130 ;
        RECT 4.430 0.000 4.810 2.270 ;
    END
  END GATE1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 7.540 6.040 10.090 6.050 ;
        RECT 7.540 0.020 10.100 6.040 ;
        RECT 7.540 0.010 10.090 0.020 ;
      LAYER met1 ;
        RECT 9.580 5.400 9.740 6.050 ;
        RECT 9.470 4.850 9.740 5.400 ;
        RECT 9.470 4.800 9.750 4.850 ;
        RECT 9.580 4.710 9.750 4.800 ;
        RECT 9.580 4.350 9.740 4.710 ;
        RECT 9.580 4.260 9.750 4.350 ;
        RECT 9.470 4.210 9.750 4.260 ;
        RECT 9.470 3.660 9.740 4.210 ;
        RECT 9.580 2.390 9.740 3.660 ;
        RECT 9.470 1.840 9.740 2.390 ;
        RECT 9.470 1.790 9.750 1.840 ;
        RECT 9.580 1.700 9.750 1.790 ;
        RECT 9.580 1.350 9.740 1.700 ;
        RECT 9.580 1.260 9.750 1.350 ;
        RECT 9.470 1.210 9.750 1.260 ;
        RECT 9.470 0.660 9.740 1.210 ;
        RECT 9.580 0.010 9.740 0.660 ;
    END
  END VINJ
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 8.770 5.370 8.930 6.050 ;
        RECT 8.770 5.350 8.970 5.370 ;
        RECT 8.750 5.110 8.980 5.350 ;
        RECT 8.770 4.890 8.970 5.110 ;
        RECT 8.770 4.170 8.930 4.890 ;
        RECT 8.770 3.950 8.970 4.170 ;
        RECT 8.750 3.710 8.980 3.950 ;
        RECT 8.770 3.690 8.970 3.710 ;
        RECT 8.770 2.360 8.930 3.690 ;
        RECT 8.770 2.340 8.970 2.360 ;
        RECT 8.750 2.100 8.980 2.340 ;
        RECT 8.770 1.880 8.970 2.100 ;
        RECT 8.770 1.170 8.930 1.880 ;
        RECT 8.770 0.950 8.970 1.170 ;
        RECT 8.750 0.710 8.980 0.950 ;
        RECT 8.770 0.690 8.970 0.710 ;
        RECT 8.770 0.010 8.930 0.690 ;
    END
  END VPWR
  PIN COLSEL1
    USE ANALOG ;
    ANTENNAGATEAREA 0.620000 ;
    PORT
      LAYER met1 ;
        RECT 9.140 5.060 9.330 6.050 ;
        RECT 9.160 4.940 9.330 5.060 ;
        RECT 9.170 4.120 9.330 4.940 ;
        RECT 9.160 4.000 9.330 4.120 ;
        RECT 9.140 3.140 9.330 4.000 ;
        RECT 9.120 2.910 9.360 3.140 ;
        RECT 9.140 2.050 9.330 2.910 ;
        RECT 9.160 1.930 9.330 2.050 ;
        RECT 9.170 1.120 9.330 1.930 ;
        RECT 9.160 1.000 9.330 1.120 ;
        RECT 9.140 0.010 9.330 1.000 ;
    END
  END COLSEL1
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER met2 ;
        RECT 7.630 5.550 7.940 5.690 ;
        RECT 7.530 5.370 10.100 5.550 ;
        RECT 7.630 5.360 7.940 5.370 ;
    END
  END DRAIN1
  PIN DRAIN2
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER met2 ;
        RECT 7.630 3.690 7.940 3.700 ;
        RECT 7.630 3.650 10.100 3.690 ;
        RECT 7.540 3.510 10.100 3.650 ;
        RECT 7.630 3.370 7.940 3.510 ;
    END
  END DRAIN2
  PIN DRAIN3
    USE ANALOG ;
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER met2 ;
        RECT 7.630 2.540 7.940 2.680 ;
        RECT 7.630 2.530 10.110 2.540 ;
        RECT 7.510 2.360 10.110 2.530 ;
        RECT 7.630 2.350 7.940 2.360 ;
    END
  END DRAIN3
  PIN DRAIN4
    USE ANALOG ;
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER met2 ;
        RECT 7.630 0.690 7.940 0.700 ;
        RECT 7.530 0.520 10.100 0.690 ;
        RECT 7.630 0.510 10.100 0.520 ;
        RECT 7.630 0.370 7.940 0.510 ;
    END
  END DRAIN4
  PIN VGND
    ANTENNADIFFAREA 1.053100 ;
    PORT
      LAYER met2 ;
        RECT 2.560 1.520 2.890 1.550 ;
        RECT 6.590 1.520 6.910 1.580 ;
        RECT 2.560 1.350 6.910 1.520 ;
        RECT 2.560 1.290 2.890 1.350 ;
        RECT 6.590 1.300 6.910 1.350 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.620 1.610 6.870 6.050 ;
        RECT 6.610 1.580 6.890 1.610 ;
        RECT 6.600 1.300 6.900 1.580 ;
        RECT 6.610 1.280 6.890 1.300 ;
        RECT 6.620 0.000 6.870 1.280 ;
      LAYER via ;
        RECT 6.620 1.310 6.880 1.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.590 1.580 2.860 6.050 ;
        RECT 2.570 1.270 2.880 1.580 ;
        RECT 2.590 0.000 2.860 1.270 ;
      LAYER via ;
        RECT 2.590 1.290 2.860 1.550 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 7.640 5.640 7.960 5.650 ;
        RECT 7.640 5.470 8.220 5.640 ;
        RECT 7.640 5.420 7.970 5.470 ;
        RECT 7.640 5.390 7.960 5.420 ;
        RECT 9.500 5.370 9.700 5.720 ;
        RECT 7.640 5.060 7.960 5.100 ;
        RECT 7.640 5.020 7.970 5.060 ;
        RECT 7.640 4.850 8.220 5.020 ;
        RECT 7.640 4.840 7.960 4.850 ;
        RECT 2.640 4.300 2.810 4.810 ;
        RECT 8.770 4.780 8.970 5.350 ;
        RECT 9.500 5.340 9.710 5.370 ;
        RECT 6.660 4.270 6.830 4.780 ;
        RECT 9.490 4.750 9.710 5.340 ;
        RECT 7.640 4.210 7.960 4.220 ;
        RECT 7.640 4.040 8.220 4.210 ;
        RECT 7.640 4.000 7.970 4.040 ;
        RECT 7.640 3.960 7.960 4.000 ;
        RECT 8.770 3.710 8.970 4.280 ;
        RECT 9.490 3.720 9.710 4.310 ;
        RECT 9.500 3.690 9.710 3.720 ;
        RECT 7.640 3.640 7.960 3.670 ;
        RECT 0.450 2.800 1.000 3.230 ;
        RECT 2.650 2.350 2.820 3.540 ;
        RECT 4.480 2.730 5.030 3.160 ;
        RECT 6.670 2.410 6.840 3.600 ;
        RECT 7.640 3.590 7.970 3.640 ;
        RECT 7.640 3.420 8.220 3.590 ;
        RECT 7.640 3.410 7.960 3.420 ;
        RECT 9.500 3.340 9.700 3.690 ;
        RECT 8.890 2.940 9.330 3.110 ;
        RECT 7.640 2.630 7.960 2.640 ;
        RECT 7.640 2.460 8.220 2.630 ;
        RECT 7.640 2.410 7.970 2.460 ;
        RECT 7.640 2.380 7.960 2.410 ;
        RECT 9.500 2.360 9.700 2.710 ;
        RECT 7.640 2.050 7.960 2.090 ;
        RECT 7.640 2.010 7.970 2.050 ;
        RECT 7.640 1.840 8.220 2.010 ;
        RECT 7.640 1.830 7.960 1.840 ;
        RECT 8.770 1.770 8.970 2.340 ;
        RECT 9.500 2.330 9.710 2.360 ;
        RECT 9.490 1.740 9.710 2.330 ;
        RECT 7.640 1.210 7.960 1.220 ;
        RECT 7.640 1.040 8.220 1.210 ;
        RECT 7.640 1.000 7.970 1.040 ;
        RECT 7.640 0.960 7.960 1.000 ;
        RECT 8.770 0.710 8.970 1.280 ;
        RECT 9.490 0.720 9.710 1.310 ;
        RECT 9.500 0.690 9.710 0.720 ;
        RECT 7.640 0.640 7.960 0.670 ;
        RECT 7.640 0.590 7.970 0.640 ;
        RECT 7.640 0.420 8.220 0.590 ;
        RECT 7.640 0.410 7.960 0.420 ;
        RECT 9.500 0.340 9.700 0.690 ;
      LAYER mcon ;
        RECT 7.700 5.430 7.870 5.600 ;
        RECT 8.780 5.140 8.950 5.310 ;
        RECT 7.700 4.880 7.870 5.050 ;
        RECT 2.640 4.640 2.810 4.810 ;
        RECT 9.510 5.170 9.680 5.340 ;
        RECT 6.660 4.610 6.830 4.780 ;
        RECT 7.700 4.010 7.870 4.180 ;
        RECT 8.780 3.750 8.950 3.920 ;
        RECT 9.510 3.720 9.680 3.890 ;
        RECT 2.650 3.370 2.820 3.540 ;
        RECT 0.450 2.880 0.720 3.150 ;
        RECT 2.650 3.030 2.820 3.200 ;
        RECT 6.670 3.430 6.840 3.600 ;
        RECT 7.700 3.460 7.870 3.630 ;
        RECT 2.650 2.690 2.820 2.860 ;
        RECT 4.480 2.810 4.750 3.080 ;
        RECT 6.670 3.090 6.840 3.260 ;
        RECT 9.150 2.940 9.330 3.110 ;
        RECT 6.670 2.750 6.840 2.920 ;
        RECT 7.700 2.420 7.870 2.590 ;
        RECT 8.780 2.130 8.950 2.300 ;
        RECT 7.700 1.870 7.870 2.040 ;
        RECT 9.510 2.160 9.680 2.330 ;
        RECT 7.700 1.010 7.870 1.180 ;
        RECT 8.780 0.750 8.950 0.920 ;
        RECT 9.510 0.720 9.680 0.890 ;
        RECT 7.700 0.460 7.870 0.630 ;
      LAYER met1 ;
        RECT 7.630 5.360 7.950 5.680 ;
        RECT 7.630 4.810 7.950 5.130 ;
        RECT 7.630 3.930 7.950 4.250 ;
        RECT 7.630 3.380 7.950 3.700 ;
        RECT 7.630 2.350 7.950 2.670 ;
        RECT 7.630 1.800 7.950 2.120 ;
        RECT 7.630 0.930 7.950 1.250 ;
        RECT 7.630 0.380 7.950 0.700 ;
      LAYER via ;
        RECT 7.660 5.390 7.920 5.650 ;
        RECT 7.660 4.840 7.920 5.100 ;
        RECT 7.660 3.960 7.920 4.220 ;
        RECT 7.660 3.410 7.920 3.670 ;
        RECT 7.660 2.380 7.920 2.640 ;
        RECT 7.660 1.830 7.920 2.090 ;
        RECT 7.660 0.960 7.920 1.220 ;
        RECT 7.660 0.410 7.920 0.670 ;
  END
END sky130_hilas_swc4x1BiasCell

MACRO sky130_hilas_FGtrans2x1cell
  CLASS CORE ;
  FOREIGN sky130_hilas_FGtrans2x1cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.520 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN COLSEL1
    USE ANALOG ;
    ANTENNAGATEAREA 0.310000 ;
    PORT
      LAYER met1 ;
        RECT 10.560 4.590 10.750 6.050 ;
        RECT 10.560 4.560 10.780 4.590 ;
        RECT 10.540 4.290 10.790 4.560 ;
        RECT 10.550 4.280 10.790 4.290 ;
        RECT 10.550 4.040 10.780 4.280 ;
        RECT 10.590 2.010 10.750 4.040 ;
        RECT 10.550 1.770 10.780 2.010 ;
        RECT 10.550 1.760 10.790 1.770 ;
        RECT 10.540 1.490 10.790 1.760 ;
        RECT 10.560 1.460 10.780 1.490 ;
        RECT 10.560 0.000 10.750 1.460 ;
    END
  END COLSEL1
  PIN VINJ
    USE ANALOG ;
    ANTENNADIFFAREA 0.510000 ;
    PORT
      LAYER nwell ;
        RECT 8.210 0.010 11.520 6.040 ;
      LAYER met1 ;
        RECT 11.000 5.400 11.160 6.050 ;
        RECT 10.890 4.850 11.160 5.400 ;
        RECT 10.890 4.800 11.170 4.850 ;
        RECT 11.000 4.710 11.170 4.800 ;
        RECT 11.000 1.340 11.160 4.710 ;
        RECT 11.000 1.250 11.170 1.340 ;
        RECT 10.890 1.200 11.170 1.250 ;
        RECT 10.890 0.650 11.160 1.200 ;
        RECT 11.000 0.000 11.160 0.650 ;
    END
  END VINJ
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.105400 ;
    PORT
      LAYER met2 ;
        RECT 8.790 5.560 9.110 5.570 ;
        RECT 8.790 5.550 9.350 5.560 ;
        RECT 0.000 5.370 11.520 5.550 ;
        RECT 9.040 5.230 9.350 5.370 ;
    END
  END DRAIN1
  PIN DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.105400 ;
    PORT
      LAYER met2 ;
        RECT 9.040 0.680 9.350 0.820 ;
        RECT 9.040 0.670 11.520 0.680 ;
        RECT 0.000 0.520 11.520 0.670 ;
        RECT 9.040 0.500 11.520 0.520 ;
        RECT 9.040 0.490 9.350 0.500 ;
    END
  END DRAIN2
  PIN PROG
    USE ANALOG ;
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER met1 ;
        RECT 7.790 3.330 8.000 6.050 ;
        RECT 7.790 2.820 8.030 3.330 ;
        RECT 7.790 0.000 8.000 2.820 ;
    END
  END PROG
  PIN RUN
    USE ANALOG ;
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER met1 ;
        RECT 6.740 1.520 6.920 6.050 ;
        RECT 6.690 1.180 6.980 1.520 ;
        RECT 6.740 0.000 6.920 1.180 ;
    END
  END RUN
  PIN VIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.217200 ;
    PORT
      LAYER met1 ;
        RECT 8.670 2.620 8.860 2.750 ;
        RECT 8.650 2.330 8.880 2.620 ;
        RECT 8.670 0.710 8.860 2.330 ;
        RECT 8.630 0.500 8.860 0.710 ;
        RECT 8.630 0.420 8.870 0.500 ;
        RECT 8.640 0.000 8.870 0.420 ;
    END
  END VIN2
  PIN VIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.217200 ;
    PORT
      LAYER met1 ;
        RECT 8.670 5.680 8.880 6.050 ;
        RECT 8.660 5.390 8.890 5.680 ;
        RECT 8.670 3.690 8.880 5.390 ;
        RECT 8.660 3.400 8.890 3.690 ;
        RECT 8.670 3.260 8.880 3.400 ;
    END
  END VIN1
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 0.434600 ;
    PORT
      LAYER met1 ;
        RECT 8.220 5.120 8.410 6.050 ;
        RECT 8.190 4.830 8.420 5.120 ;
        RECT 8.220 2.800 8.410 4.830 ;
        RECT 8.190 2.510 8.420 2.800 ;
        RECT 8.220 1.220 8.410 2.510 ;
        RECT 8.200 0.930 8.430 1.220 ;
        RECT 8.220 0.000 8.410 0.930 ;
    END
  END GATE1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2.820 0.000 3.050 6.050 ;
    END
  END VGND
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 2.516100 ;
    PORT
      LAYER nwell ;
        RECT 0.000 5.300 1.730 6.050 ;
        RECT 0.000 1.730 1.740 5.300 ;
        RECT 0.000 0.010 1.730 1.730 ;
      LAYER met1 ;
        RECT 0.340 0.000 0.760 6.050 ;
    END
  END VTUN
  PIN COL1
    ANTENNADIFFAREA 1.030400 ;
    PORT
      LAYER met2 ;
        RECT 10.140 3.130 10.460 3.160 ;
        RECT 0.000 2.900 10.460 3.130 ;
    END
  END COL1
  PIN ROW1
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 9.430 4.010 9.740 4.030 ;
        RECT 0.000 3.820 9.740 4.010 ;
        RECT 9.430 3.700 9.740 3.820 ;
    END
  END ROW1
  PIN ROW2
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 9.440 2.150 9.750 2.340 ;
        RECT 0.000 2.010 9.750 2.150 ;
        RECT 0.000 1.960 9.720 2.010 ;
    END
  END ROW2
  OBS
      LAYER nwell ;
        RECT 3.760 3.660 6.480 5.310 ;
        RECT 3.770 3.620 6.480 3.660 ;
        RECT 3.770 2.290 6.480 2.330 ;
        RECT 3.760 0.640 6.480 2.290 ;
      LAYER li1 ;
        RECT 8.680 5.620 8.870 5.650 ;
        RECT 7.810 5.450 8.870 5.620 ;
        RECT 9.110 5.470 9.640 5.640 ;
        RECT 7.810 5.060 7.980 5.450 ;
        RECT 8.680 5.420 8.870 5.450 ;
        RECT 10.920 5.370 11.120 5.720 ;
        RECT 10.920 5.340 11.130 5.370 ;
        RECT 7.240 4.890 7.980 5.060 ;
        RECT 8.210 5.060 8.400 5.090 ;
        RECT 8.210 4.890 8.940 5.060 ;
        RECT 8.210 4.860 8.400 4.890 ;
        RECT 0.430 3.910 0.980 4.340 ;
        RECT 5.950 4.270 6.180 4.790 ;
        RECT 5.950 4.100 8.940 4.270 ;
        RECT 9.360 3.990 9.530 5.080 ;
        RECT 9.360 3.950 9.760 3.990 ;
        RECT 9.360 3.760 9.770 3.950 ;
        RECT 9.360 3.730 9.760 3.760 ;
        RECT 8.680 3.480 8.870 3.660 ;
        RECT 3.030 3.080 3.220 3.480 ;
        RECT 7.250 3.310 7.590 3.480 ;
        RECT 2.840 3.070 3.220 3.080 ;
        RECT 2.840 2.890 6.580 3.070 ;
        RECT 2.840 2.850 3.220 2.890 ;
        RECT 0.430 2.180 0.980 2.610 ;
        RECT 3.030 2.470 3.220 2.850 ;
        RECT 7.330 2.740 7.500 3.310 ;
        RECT 7.810 2.900 8.020 3.330 ;
        RECT 8.590 3.310 8.940 3.480 ;
        RECT 9.360 3.390 9.530 3.730 ;
        RECT 10.190 3.480 10.360 5.090 ;
        RECT 10.910 4.760 11.130 5.340 ;
        RECT 10.920 4.750 11.130 4.760 ;
        RECT 10.560 4.580 10.750 4.590 ;
        RECT 10.560 4.290 10.760 4.580 ;
        RECT 10.550 3.960 10.790 4.290 ;
        RECT 10.190 3.290 10.370 3.480 ;
        RECT 7.830 2.880 8.000 2.900 ;
        RECT 7.250 2.710 7.590 2.740 ;
        RECT 8.210 2.720 8.400 2.770 ;
        RECT 8.170 2.710 8.400 2.720 ;
        RECT 7.250 2.570 8.400 2.710 ;
        RECT 8.590 2.570 8.940 2.740 ;
        RECT 7.420 2.540 8.400 2.570 ;
        RECT 7.420 2.510 8.260 2.540 ;
        RECT 8.670 2.360 8.860 2.570 ;
        RECT 9.360 2.300 9.530 2.660 ;
        RECT 10.190 2.570 10.370 2.760 ;
        RECT 9.360 2.260 9.770 2.300 ;
        RECT 9.360 2.070 9.780 2.260 ;
        RECT 9.360 2.040 9.770 2.070 ;
        RECT 6.010 1.850 8.940 1.950 ;
        RECT 5.950 1.780 8.940 1.850 ;
        RECT 5.950 1.160 6.180 1.780 ;
        RECT 6.750 1.460 6.920 1.520 ;
        RECT 6.730 1.250 6.940 1.460 ;
        RECT 6.750 1.180 6.920 1.250 ;
        RECT 8.220 1.160 8.410 1.190 ;
        RECT 7.240 0.990 8.050 1.160 ;
        RECT 7.860 0.650 8.050 0.990 ;
        RECT 8.220 0.990 8.940 1.160 ;
        RECT 8.220 0.960 8.410 0.990 ;
        RECT 9.360 0.970 9.530 2.040 ;
        RECT 10.190 0.960 10.360 2.570 ;
        RECT 10.550 1.760 10.790 2.090 ;
        RECT 10.560 1.470 10.760 1.760 ;
        RECT 10.560 1.460 10.750 1.470 ;
        RECT 10.920 1.290 11.130 1.300 ;
        RECT 10.910 0.710 11.130 1.290 ;
        RECT 10.920 0.680 11.130 0.710 ;
        RECT 8.650 0.650 8.840 0.680 ;
        RECT 7.860 0.470 8.840 0.650 ;
        RECT 8.650 0.450 8.840 0.470 ;
        RECT 9.110 0.410 9.640 0.580 ;
        RECT 10.920 0.330 11.120 0.680 ;
      LAYER mcon ;
        RECT 8.690 5.450 8.860 5.620 ;
        RECT 10.930 5.170 11.100 5.340 ;
        RECT 8.220 4.890 8.390 5.060 ;
        RECT 5.980 4.590 6.150 4.760 ;
        RECT 0.430 3.990 0.700 4.260 ;
        RECT 5.980 4.140 6.150 4.310 ;
        RECT 9.500 3.770 9.670 3.940 ;
        RECT 8.690 3.460 8.860 3.630 ;
        RECT 2.850 2.880 3.020 3.050 ;
        RECT 0.430 2.260 0.700 2.530 ;
        RECT 10.570 4.330 10.750 4.520 ;
        RECT 8.220 2.570 8.390 2.740 ;
        RECT 8.680 2.390 8.850 2.560 ;
        RECT 9.510 2.080 9.680 2.250 ;
        RECT 5.980 1.640 6.150 1.810 ;
        RECT 5.980 1.190 6.150 1.360 ;
        RECT 8.230 0.990 8.400 1.160 ;
        RECT 10.570 1.530 10.750 1.720 ;
        RECT 10.930 0.710 11.100 0.880 ;
        RECT 8.660 0.480 8.830 0.650 ;
      LAYER met1 ;
        RECT 9.040 5.230 9.350 5.670 ;
        RECT 5.940 4.050 6.200 4.840 ;
        RECT 9.430 3.700 9.750 4.020 ;
        RECT 10.160 3.190 10.400 3.610 ;
        RECT 10.160 2.870 10.430 3.190 ;
        RECT 10.160 2.440 10.400 2.870 ;
        RECT 9.440 2.010 9.760 2.330 ;
        RECT 5.940 1.110 6.200 1.900 ;
        RECT 9.040 0.380 9.350 0.820 ;
      LAYER via ;
        RECT 9.070 5.260 9.330 5.520 ;
        RECT 9.460 3.730 9.720 3.990 ;
        RECT 10.170 2.900 10.430 3.160 ;
        RECT 9.470 2.040 9.730 2.300 ;
        RECT 9.070 0.530 9.330 0.790 ;
  END
END sky130_hilas_FGtrans2x1cell

MACRO sky130_hilas_capacitorSize01
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.420 BY 5.830 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 9.600 2.610 10.260 3.270 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 0.110 3.200 0.770 3.260 ;
        RECT 1.160 3.200 2.170 3.210 ;
        RECT 0.110 2.700 3.800 3.200 ;
        RECT 0.110 2.690 1.520 2.700 ;
        RECT 0.110 2.600 0.770 2.690 ;
        RECT 3.160 1.580 3.790 2.700 ;
        RECT 3.160 1.570 5.310 1.580 ;
        RECT 2.350 1.100 5.390 1.570 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 0.000 5.280 10.420 5.460 ;
        RECT 0.000 4.850 10.420 5.030 ;
        RECT 0.030 3.850 10.420 4.030 ;
        RECT 8.510 3.600 10.420 3.610 ;
        RECT 0.030 3.420 10.420 3.600 ;
        RECT 0.240 3.080 0.610 3.140 ;
        RECT 0.020 2.800 0.610 3.080 ;
        RECT 0.240 2.740 0.610 2.800 ;
        RECT 9.730 3.090 10.100 3.150 ;
        RECT 9.730 2.810 10.420 3.090 ;
        RECT 9.730 2.750 10.100 2.810 ;
        RECT 0.030 2.270 10.420 2.440 ;
        RECT 0.030 1.850 10.420 2.020 ;
        RECT 0.030 0.870 10.420 1.040 ;
        RECT 0.030 0.430 10.420 0.600 ;
      LAYER via2 ;
        RECT 0.290 2.800 0.570 3.080 ;
        RECT 9.780 2.810 10.060 3.090 ;
      LAYER met3 ;
        RECT 1.460 5.800 4.280 5.830 ;
        RECT 1.460 3.300 8.660 5.800 ;
        RECT 0.020 2.540 0.810 3.290 ;
        RECT 1.460 2.550 10.300 3.300 ;
        RECT 1.460 0.020 8.660 2.550 ;
        RECT 4.250 0.000 8.660 0.020 ;
      LAYER via3 ;
        RECT 0.210 2.690 0.640 3.170 ;
        RECT 9.700 2.700 10.130 3.180 ;
  END
END sky130_hilas_capacitorSize01

MACRO sky130_hilas_Tgate4Double01
  CLASS CORE ;
  FOREIGN sky130_hilas_Tgate4Double01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.080 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER nwell ;
        RECT 0.120 0.000 3.590 6.050 ;
      LAYER met1 ;
        RECT 0.740 5.180 0.940 6.050 ;
        RECT 0.730 4.890 0.960 5.180 ;
        RECT 0.740 4.180 0.940 4.890 ;
        RECT 0.730 3.890 0.960 4.180 ;
        RECT 0.740 2.160 0.940 3.890 ;
        RECT 0.730 1.870 0.960 2.160 ;
        RECT 0.740 1.160 0.940 1.870 ;
        RECT 0.730 0.870 0.960 1.160 ;
        RECT 0.740 0.000 0.940 0.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.570 5.180 6.760 6.050 ;
        RECT 6.550 4.890 6.780 5.180 ;
        RECT 6.570 4.180 6.760 4.890 ;
        RECT 6.550 3.890 6.780 4.180 ;
        RECT 6.570 2.160 6.760 3.890 ;
        RECT 6.550 1.870 6.780 2.160 ;
        RECT 6.570 1.160 6.760 1.870 ;
        RECT 6.550 0.870 6.780 1.160 ;
        RECT 6.570 0.000 6.760 0.870 ;
    END
  END VGND
  PIN INPUT1_1
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.450 5.940 2.760 5.950 ;
        RECT 0.000 5.740 5.840 5.940 ;
        RECT 2.450 5.620 2.760 5.740 ;
        RECT 5.530 5.610 5.840 5.740 ;
    END
  END INPUT1_1
  PIN SELECT1
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER met2 ;
        RECT 0.000 4.760 0.610 4.960 ;
        RECT 0.290 4.670 0.610 4.760 ;
    END
  END SELECT1
  PIN SELECT2
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER met2 ;
        RECT 0.290 4.310 0.610 4.400 ;
        RECT 0.000 4.110 0.610 4.310 ;
    END
  END SELECT2
  PIN INPUT2_2
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 1.100 3.810 1.410 3.820 ;
        RECT 4.020 3.810 4.330 3.820 ;
        RECT 0.000 3.610 4.370 3.810 ;
        RECT 1.100 3.490 1.410 3.610 ;
        RECT 4.020 3.490 4.330 3.610 ;
    END
  END INPUT2_2
  PIN INPUT1_2
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.450 3.330 2.760 3.450 ;
        RECT 5.530 3.330 5.840 3.460 ;
        RECT 0.000 3.130 5.840 3.330 ;
        RECT 2.450 3.120 2.760 3.130 ;
    END
  END INPUT1_2
  PIN SELECT3
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER met2 ;
        RECT 0.000 1.740 0.610 1.940 ;
        RECT 0.290 1.650 0.610 1.740 ;
    END
  END SELECT3
  PIN INPUT2_3
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 1.100 2.440 1.410 2.560 ;
        RECT 4.020 2.440 4.330 2.560 ;
        RECT 0.000 2.240 4.370 2.440 ;
        RECT 1.100 2.230 1.410 2.240 ;
        RECT 4.020 2.230 4.330 2.240 ;
    END
  END INPUT2_3
  PIN SELECT4
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER met2 ;
        RECT 0.290 1.290 0.610 1.380 ;
        RECT 0.000 1.090 0.610 1.290 ;
    END
  END SELECT4
  PIN INPUT2_4
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 1.100 0.790 1.410 0.800 ;
        RECT 4.020 0.790 4.330 0.800 ;
        RECT 0.000 0.590 4.370 0.790 ;
        RECT 1.100 0.470 1.410 0.590 ;
        RECT 4.020 0.470 4.330 0.590 ;
    END
  END INPUT2_4
  PIN INPUT1_4
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.450 0.310 2.760 0.430 ;
        RECT 5.530 0.310 5.840 0.440 ;
        RECT 0.000 0.110 5.840 0.310 ;
        RECT 2.450 0.100 2.760 0.110 ;
    END
  END INPUT1_4
  PIN OUTPUT4
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER met2 ;
        RECT 1.680 1.290 2.000 1.300 ;
        RECT 3.100 1.290 3.420 1.310 ;
        RECT 4.850 1.290 5.170 1.330 ;
        RECT 5.890 1.290 6.210 1.320 ;
        RECT 1.680 1.090 7.080 1.290 ;
        RECT 1.680 1.040 2.000 1.090 ;
        RECT 3.100 1.050 3.420 1.090 ;
        RECT 4.850 1.070 5.170 1.090 ;
        RECT 5.890 1.060 6.210 1.090 ;
    END
  END OUTPUT4
  PIN OUTPUT3
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER met2 ;
        RECT 1.680 1.940 2.000 1.990 ;
        RECT 3.100 1.940 3.420 1.980 ;
        RECT 4.850 1.940 5.170 1.960 ;
        RECT 5.890 1.940 6.210 1.970 ;
        RECT 1.680 1.740 7.080 1.940 ;
        RECT 1.680 1.730 2.000 1.740 ;
        RECT 3.100 1.720 3.420 1.740 ;
        RECT 4.850 1.700 5.170 1.740 ;
        RECT 5.890 1.710 6.210 1.740 ;
    END
  END OUTPUT3
  PIN OUTPUT2
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER met2 ;
        RECT 1.680 4.310 2.000 4.320 ;
        RECT 3.100 4.310 3.420 4.330 ;
        RECT 4.850 4.310 5.170 4.350 ;
        RECT 5.890 4.310 6.210 4.340 ;
        RECT 1.680 4.110 7.080 4.310 ;
        RECT 1.680 4.060 2.000 4.110 ;
        RECT 3.100 4.070 3.420 4.110 ;
        RECT 4.850 4.090 5.170 4.110 ;
        RECT 5.890 4.080 6.210 4.110 ;
    END
  END OUTPUT2
  PIN OUTPUT1
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER met2 ;
        RECT 1.680 4.960 2.000 5.010 ;
        RECT 3.100 4.960 3.420 5.000 ;
        RECT 4.850 4.960 5.170 4.980 ;
        RECT 5.890 4.960 6.210 4.990 ;
        RECT 1.680 4.760 7.080 4.960 ;
        RECT 1.680 4.750 2.000 4.760 ;
        RECT 3.100 4.740 3.420 4.760 ;
        RECT 4.850 4.720 5.170 4.760 ;
        RECT 5.890 4.730 6.210 4.760 ;
    END
  END OUTPUT1
  PIN INPUT2_1
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 1.100 5.460 1.410 5.580 ;
        RECT 4.020 5.460 4.330 5.580 ;
        RECT 0.000 5.260 4.370 5.460 ;
        RECT 1.100 5.250 1.410 5.260 ;
        RECT 4.020 5.250 4.330 5.260 ;
    END
  END INPUT2_1
  PIN INPUT1_3
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.450 2.920 2.760 2.930 ;
        RECT 0.000 2.720 5.840 2.920 ;
        RECT 2.450 2.600 2.760 2.720 ;
        RECT 5.530 2.590 5.840 2.720 ;
    END
  END INPUT1_3
  OBS
      LAYER li1 ;
        RECT 2.460 5.890 2.780 5.920 ;
        RECT 0.430 5.540 0.600 5.820 ;
        RECT 0.940 5.580 1.290 5.750 ;
        RECT 1.110 5.550 1.290 5.580 ;
        RECT 1.710 5.560 1.880 5.830 ;
        RECT 2.460 5.700 2.790 5.890 ;
        RECT 5.540 5.880 5.860 5.910 ;
        RECT 2.460 5.660 2.780 5.700 ;
        RECT 0.430 5.500 0.640 5.540 ;
        RECT 1.110 5.520 1.430 5.550 ;
        RECT 0.430 5.480 0.660 5.500 ;
        RECT 0.430 5.460 0.690 5.480 ;
        RECT 0.430 5.410 0.770 5.460 ;
        RECT 0.430 5.350 0.920 5.410 ;
        RECT 0.430 5.320 0.940 5.350 ;
        RECT 0.470 5.290 0.940 5.320 ;
        RECT 1.110 5.330 1.440 5.520 ;
        RECT 1.710 5.340 1.910 5.560 ;
        RECT 2.490 5.490 2.660 5.660 ;
        RECT 3.180 5.540 3.350 5.830 ;
        RECT 4.140 5.550 4.310 5.830 ;
        RECT 4.880 5.550 5.050 5.840 ;
        RECT 5.540 5.690 5.870 5.880 ;
        RECT 6.110 5.740 6.300 5.770 ;
        RECT 5.540 5.650 5.860 5.690 ;
        RECT 1.720 5.330 1.910 5.340 ;
        RECT 1.110 5.290 1.430 5.330 ;
        RECT 3.170 5.310 3.360 5.540 ;
        RECT 4.030 5.520 4.350 5.550 ;
        RECT 4.030 5.330 4.360 5.520 ;
        RECT 4.030 5.290 4.350 5.330 ;
        RECT 4.880 5.320 5.070 5.550 ;
        RECT 5.600 5.490 5.770 5.650 ;
        RECT 6.110 5.570 6.550 5.740 ;
        RECT 6.110 5.540 6.300 5.570 ;
        RECT 0.600 5.240 0.940 5.290 ;
        RECT 0.720 5.230 0.940 5.240 ;
        RECT 0.730 5.200 0.940 5.230 ;
        RECT 0.750 5.120 0.940 5.200 ;
        RECT 2.110 5.120 2.440 5.240 ;
        RECT 6.830 5.150 7.000 5.830 ;
        RECT 0.260 5.070 0.430 5.090 ;
        RECT 0.240 4.640 0.450 5.070 ;
        RECT 0.750 4.950 1.270 5.120 ;
        RECT 0.750 4.920 0.940 4.950 ;
        RECT 1.620 4.940 5.840 5.120 ;
        RECT 6.570 5.110 7.000 5.150 ;
        RECT 6.220 4.950 7.000 5.110 ;
        RECT 6.220 4.940 6.760 4.950 ;
        RECT 6.570 4.920 6.760 4.940 ;
        RECT 0.240 4.000 0.450 4.430 ;
        RECT 0.750 4.120 0.940 4.150 ;
        RECT 6.570 4.130 6.760 4.150 ;
        RECT 0.260 3.980 0.430 4.000 ;
        RECT 0.750 3.950 1.270 4.120 ;
        RECT 1.620 3.950 5.840 4.130 ;
        RECT 6.220 4.120 6.760 4.130 ;
        RECT 6.220 3.960 7.000 4.120 ;
        RECT 0.750 3.870 0.940 3.950 ;
        RECT 0.730 3.840 0.940 3.870 ;
        RECT 0.720 3.830 0.940 3.840 ;
        RECT 2.110 3.830 2.440 3.950 ;
        RECT 6.570 3.920 7.000 3.960 ;
        RECT 0.600 3.780 0.940 3.830 ;
        RECT 0.470 3.750 0.940 3.780 ;
        RECT 0.430 3.720 0.940 3.750 ;
        RECT 1.110 3.740 1.430 3.780 ;
        RECT 0.430 3.660 0.920 3.720 ;
        RECT 0.430 3.610 0.770 3.660 ;
        RECT 0.430 3.590 0.690 3.610 ;
        RECT 0.430 3.570 0.660 3.590 ;
        RECT 0.430 3.530 0.640 3.570 ;
        RECT 1.110 3.550 1.440 3.740 ;
        RECT 1.720 3.730 1.910 3.740 ;
        RECT 0.430 3.250 0.600 3.530 ;
        RECT 1.110 3.520 1.430 3.550 ;
        RECT 1.110 3.490 1.290 3.520 ;
        RECT 0.940 3.320 1.290 3.490 ;
        RECT 1.710 3.510 1.910 3.730 ;
        RECT 1.710 3.240 1.880 3.510 ;
        RECT 2.490 3.410 2.660 3.580 ;
        RECT 3.170 3.530 3.360 3.760 ;
        RECT 4.030 3.740 4.350 3.780 ;
        RECT 4.030 3.550 4.360 3.740 ;
        RECT 2.460 3.370 2.780 3.410 ;
        RECT 2.460 3.180 2.790 3.370 ;
        RECT 3.180 3.240 3.350 3.530 ;
        RECT 4.030 3.520 4.350 3.550 ;
        RECT 4.880 3.520 5.070 3.750 ;
        RECT 4.140 3.240 4.310 3.520 ;
        RECT 4.880 3.230 5.050 3.520 ;
        RECT 5.600 3.420 5.770 3.580 ;
        RECT 6.110 3.500 6.300 3.530 ;
        RECT 5.540 3.380 5.860 3.420 ;
        RECT 5.540 3.190 5.870 3.380 ;
        RECT 6.110 3.330 6.550 3.500 ;
        RECT 6.110 3.300 6.300 3.330 ;
        RECT 6.830 3.240 7.000 3.920 ;
        RECT 2.460 3.150 2.780 3.180 ;
        RECT 5.540 3.160 5.860 3.190 ;
        RECT 2.460 2.870 2.780 2.900 ;
        RECT 0.430 2.520 0.600 2.800 ;
        RECT 0.940 2.560 1.290 2.730 ;
        RECT 1.110 2.530 1.290 2.560 ;
        RECT 1.710 2.540 1.880 2.810 ;
        RECT 2.460 2.680 2.790 2.870 ;
        RECT 5.540 2.860 5.860 2.890 ;
        RECT 2.460 2.640 2.780 2.680 ;
        RECT 0.430 2.480 0.640 2.520 ;
        RECT 1.110 2.500 1.430 2.530 ;
        RECT 0.430 2.460 0.660 2.480 ;
        RECT 0.430 2.440 0.690 2.460 ;
        RECT 0.430 2.390 0.770 2.440 ;
        RECT 0.430 2.330 0.920 2.390 ;
        RECT 0.430 2.300 0.940 2.330 ;
        RECT 0.470 2.270 0.940 2.300 ;
        RECT 1.110 2.310 1.440 2.500 ;
        RECT 1.710 2.320 1.910 2.540 ;
        RECT 2.490 2.470 2.660 2.640 ;
        RECT 3.180 2.520 3.350 2.810 ;
        RECT 4.140 2.530 4.310 2.810 ;
        RECT 4.880 2.530 5.050 2.820 ;
        RECT 5.540 2.670 5.870 2.860 ;
        RECT 6.110 2.720 6.300 2.750 ;
        RECT 5.540 2.630 5.860 2.670 ;
        RECT 1.720 2.310 1.910 2.320 ;
        RECT 1.110 2.270 1.430 2.310 ;
        RECT 3.170 2.290 3.360 2.520 ;
        RECT 4.030 2.500 4.350 2.530 ;
        RECT 4.030 2.310 4.360 2.500 ;
        RECT 4.030 2.270 4.350 2.310 ;
        RECT 4.880 2.300 5.070 2.530 ;
        RECT 5.600 2.470 5.770 2.630 ;
        RECT 6.110 2.550 6.550 2.720 ;
        RECT 6.110 2.520 6.300 2.550 ;
        RECT 0.600 2.220 0.940 2.270 ;
        RECT 0.720 2.210 0.940 2.220 ;
        RECT 0.730 2.180 0.940 2.210 ;
        RECT 0.750 2.100 0.940 2.180 ;
        RECT 2.110 2.100 2.440 2.220 ;
        RECT 6.830 2.130 7.000 2.810 ;
        RECT 0.260 2.050 0.430 2.070 ;
        RECT 0.240 1.620 0.450 2.050 ;
        RECT 0.750 1.930 1.270 2.100 ;
        RECT 0.750 1.900 0.940 1.930 ;
        RECT 1.620 1.920 5.840 2.100 ;
        RECT 6.570 2.090 7.000 2.130 ;
        RECT 6.220 1.930 7.000 2.090 ;
        RECT 6.220 1.920 6.760 1.930 ;
        RECT 6.570 1.900 6.760 1.920 ;
        RECT 0.240 0.980 0.450 1.410 ;
        RECT 0.750 1.100 0.940 1.130 ;
        RECT 6.570 1.110 6.760 1.130 ;
        RECT 0.260 0.960 0.430 0.980 ;
        RECT 0.750 0.930 1.270 1.100 ;
        RECT 1.620 0.930 5.840 1.110 ;
        RECT 6.220 1.100 6.760 1.110 ;
        RECT 6.220 0.940 7.000 1.100 ;
        RECT 0.750 0.850 0.940 0.930 ;
        RECT 0.730 0.820 0.940 0.850 ;
        RECT 0.720 0.810 0.940 0.820 ;
        RECT 2.110 0.810 2.440 0.930 ;
        RECT 6.570 0.900 7.000 0.940 ;
        RECT 0.600 0.760 0.940 0.810 ;
        RECT 0.470 0.730 0.940 0.760 ;
        RECT 0.430 0.700 0.940 0.730 ;
        RECT 1.110 0.720 1.430 0.760 ;
        RECT 0.430 0.640 0.920 0.700 ;
        RECT 0.430 0.590 0.770 0.640 ;
        RECT 0.430 0.570 0.690 0.590 ;
        RECT 0.430 0.550 0.660 0.570 ;
        RECT 0.430 0.510 0.640 0.550 ;
        RECT 1.110 0.530 1.440 0.720 ;
        RECT 1.720 0.710 1.910 0.720 ;
        RECT 0.430 0.230 0.600 0.510 ;
        RECT 1.110 0.500 1.430 0.530 ;
        RECT 1.110 0.470 1.290 0.500 ;
        RECT 0.940 0.300 1.290 0.470 ;
        RECT 1.710 0.490 1.910 0.710 ;
        RECT 1.710 0.220 1.880 0.490 ;
        RECT 2.490 0.390 2.660 0.560 ;
        RECT 3.170 0.510 3.360 0.740 ;
        RECT 4.030 0.720 4.350 0.760 ;
        RECT 4.030 0.530 4.360 0.720 ;
        RECT 2.460 0.350 2.780 0.390 ;
        RECT 2.460 0.160 2.790 0.350 ;
        RECT 3.180 0.220 3.350 0.510 ;
        RECT 4.030 0.500 4.350 0.530 ;
        RECT 4.880 0.500 5.070 0.730 ;
        RECT 4.140 0.220 4.310 0.500 ;
        RECT 4.880 0.210 5.050 0.500 ;
        RECT 5.600 0.400 5.770 0.560 ;
        RECT 6.110 0.480 6.300 0.510 ;
        RECT 5.540 0.360 5.860 0.400 ;
        RECT 5.540 0.170 5.870 0.360 ;
        RECT 6.110 0.310 6.550 0.480 ;
        RECT 6.110 0.280 6.300 0.310 ;
        RECT 6.830 0.220 7.000 0.900 ;
        RECT 2.460 0.130 2.780 0.160 ;
        RECT 5.540 0.140 5.860 0.170 ;
      LAYER mcon ;
        RECT 2.520 5.710 2.690 5.880 ;
        RECT 1.170 5.340 1.340 5.510 ;
        RECT 1.730 5.360 1.900 5.530 ;
        RECT 5.600 5.700 5.770 5.870 ;
        RECT 3.180 5.340 3.350 5.510 ;
        RECT 4.090 5.340 4.260 5.510 ;
        RECT 4.890 5.350 5.060 5.520 ;
        RECT 6.120 5.570 6.290 5.740 ;
        RECT 0.260 4.920 0.430 5.090 ;
        RECT 0.760 4.950 0.930 5.120 ;
        RECT 6.580 4.950 6.750 5.120 ;
        RECT 0.760 3.950 0.930 4.120 ;
        RECT 6.580 3.950 6.750 4.120 ;
        RECT 1.170 3.560 1.340 3.730 ;
        RECT 1.730 3.540 1.900 3.710 ;
        RECT 3.180 3.560 3.350 3.730 ;
        RECT 4.090 3.560 4.260 3.730 ;
        RECT 4.890 3.550 5.060 3.720 ;
        RECT 2.520 3.190 2.690 3.360 ;
        RECT 5.600 3.200 5.770 3.370 ;
        RECT 6.120 3.330 6.290 3.500 ;
        RECT 2.520 2.690 2.690 2.860 ;
        RECT 1.170 2.320 1.340 2.490 ;
        RECT 1.730 2.340 1.900 2.510 ;
        RECT 5.600 2.680 5.770 2.850 ;
        RECT 3.180 2.320 3.350 2.490 ;
        RECT 4.090 2.320 4.260 2.490 ;
        RECT 4.890 2.330 5.060 2.500 ;
        RECT 6.120 2.550 6.290 2.720 ;
        RECT 0.260 1.900 0.430 2.070 ;
        RECT 0.760 1.930 0.930 2.100 ;
        RECT 6.580 1.930 6.750 2.100 ;
        RECT 0.760 0.930 0.930 1.100 ;
        RECT 6.580 0.930 6.750 1.100 ;
        RECT 1.170 0.540 1.340 0.710 ;
        RECT 1.730 0.520 1.900 0.690 ;
        RECT 3.180 0.540 3.350 0.710 ;
        RECT 4.090 0.540 4.260 0.710 ;
        RECT 4.890 0.530 5.060 0.700 ;
        RECT 2.520 0.170 2.690 0.340 ;
        RECT 5.600 0.180 5.770 0.350 ;
        RECT 6.120 0.310 6.290 0.480 ;
      LAYER met1 ;
        RECT 2.450 5.630 2.770 5.950 ;
        RECT 5.530 5.620 5.850 5.940 ;
        RECT 1.100 5.260 1.420 5.580 ;
        RECT 1.700 5.300 1.930 5.590 ;
        RECT 0.230 4.960 0.460 5.150 ;
        RECT 1.720 5.040 1.890 5.300 ;
        RECT 3.150 5.280 3.380 5.570 ;
        RECT 0.230 4.860 0.580 4.960 ;
        RECT 0.240 4.640 0.580 4.860 ;
        RECT 1.710 4.720 1.970 5.040 ;
        RECT 3.170 5.030 3.340 5.280 ;
        RECT 4.020 5.260 4.340 5.580 ;
        RECT 4.860 5.290 5.090 5.580 ;
        RECT 6.090 5.510 6.320 5.800 ;
        RECT 3.130 4.710 3.390 5.030 ;
        RECT 4.890 5.010 5.060 5.290 ;
        RECT 6.090 5.020 6.280 5.510 ;
        RECT 4.880 4.690 5.140 5.010 ;
        RECT 5.920 4.770 6.280 5.020 ;
        RECT 5.920 4.700 6.180 4.770 ;
        RECT 0.240 4.210 0.580 4.430 ;
        RECT 0.230 4.110 0.580 4.210 ;
        RECT 0.230 3.920 0.460 4.110 ;
        RECT 1.710 4.030 1.970 4.350 ;
        RECT 3.130 4.040 3.390 4.360 ;
        RECT 4.880 4.060 5.140 4.380 ;
        RECT 5.920 4.300 6.180 4.370 ;
        RECT 1.100 3.490 1.420 3.810 ;
        RECT 1.720 3.770 1.890 4.030 ;
        RECT 3.170 3.790 3.340 4.040 ;
        RECT 1.700 3.480 1.930 3.770 ;
        RECT 3.150 3.500 3.380 3.790 ;
        RECT 4.020 3.490 4.340 3.810 ;
        RECT 4.890 3.780 5.060 4.060 ;
        RECT 5.920 4.050 6.280 4.300 ;
        RECT 4.860 3.490 5.090 3.780 ;
        RECT 6.090 3.560 6.280 4.050 ;
        RECT 2.450 3.120 2.770 3.440 ;
        RECT 5.530 3.130 5.850 3.450 ;
        RECT 6.090 3.270 6.320 3.560 ;
        RECT 2.450 2.610 2.770 2.930 ;
        RECT 5.530 2.600 5.850 2.920 ;
        RECT 1.100 2.240 1.420 2.560 ;
        RECT 1.700 2.280 1.930 2.570 ;
        RECT 0.230 1.940 0.460 2.130 ;
        RECT 1.720 2.020 1.890 2.280 ;
        RECT 3.150 2.260 3.380 2.550 ;
        RECT 0.230 1.840 0.580 1.940 ;
        RECT 0.240 1.620 0.580 1.840 ;
        RECT 1.710 1.700 1.970 2.020 ;
        RECT 3.170 2.010 3.340 2.260 ;
        RECT 4.020 2.240 4.340 2.560 ;
        RECT 4.860 2.270 5.090 2.560 ;
        RECT 6.090 2.490 6.320 2.780 ;
        RECT 3.130 1.690 3.390 2.010 ;
        RECT 4.890 1.990 5.060 2.270 ;
        RECT 6.090 2.000 6.280 2.490 ;
        RECT 4.880 1.670 5.140 1.990 ;
        RECT 5.920 1.750 6.280 2.000 ;
        RECT 5.920 1.680 6.180 1.750 ;
        RECT 0.240 1.190 0.580 1.410 ;
        RECT 0.230 1.090 0.580 1.190 ;
        RECT 0.230 0.900 0.460 1.090 ;
        RECT 1.710 1.010 1.970 1.330 ;
        RECT 3.130 1.020 3.390 1.340 ;
        RECT 4.880 1.040 5.140 1.360 ;
        RECT 5.920 1.280 6.180 1.350 ;
        RECT 1.100 0.470 1.420 0.790 ;
        RECT 1.720 0.750 1.890 1.010 ;
        RECT 3.170 0.770 3.340 1.020 ;
        RECT 1.700 0.460 1.930 0.750 ;
        RECT 3.150 0.480 3.380 0.770 ;
        RECT 4.020 0.470 4.340 0.790 ;
        RECT 4.890 0.760 5.060 1.040 ;
        RECT 5.920 1.030 6.280 1.280 ;
        RECT 4.860 0.470 5.090 0.760 ;
        RECT 6.090 0.540 6.280 1.030 ;
        RECT 2.450 0.100 2.770 0.420 ;
        RECT 5.530 0.110 5.850 0.430 ;
        RECT 6.090 0.250 6.320 0.540 ;
      LAYER via ;
        RECT 2.480 5.660 2.740 5.920 ;
        RECT 5.560 5.650 5.820 5.910 ;
        RECT 1.130 5.290 1.390 5.550 ;
        RECT 4.050 5.290 4.310 5.550 ;
        RECT 0.320 4.670 0.580 4.930 ;
        RECT 1.710 4.750 1.970 5.010 ;
        RECT 3.130 4.740 3.390 5.000 ;
        RECT 4.880 4.720 5.140 4.980 ;
        RECT 5.920 4.730 6.180 4.990 ;
        RECT 0.320 4.140 0.580 4.400 ;
        RECT 1.710 4.060 1.970 4.320 ;
        RECT 3.130 4.070 3.390 4.330 ;
        RECT 4.880 4.090 5.140 4.350 ;
        RECT 5.920 4.080 6.180 4.340 ;
        RECT 1.130 3.520 1.390 3.780 ;
        RECT 4.050 3.520 4.310 3.780 ;
        RECT 2.480 3.150 2.740 3.410 ;
        RECT 5.560 3.160 5.820 3.420 ;
        RECT 2.480 2.640 2.740 2.900 ;
        RECT 5.560 2.630 5.820 2.890 ;
        RECT 1.130 2.270 1.390 2.530 ;
        RECT 4.050 2.270 4.310 2.530 ;
        RECT 0.320 1.650 0.580 1.910 ;
        RECT 1.710 1.730 1.970 1.990 ;
        RECT 3.130 1.720 3.390 1.980 ;
        RECT 4.880 1.700 5.140 1.960 ;
        RECT 5.920 1.710 6.180 1.970 ;
        RECT 0.320 1.120 0.580 1.380 ;
        RECT 1.710 1.040 1.970 1.300 ;
        RECT 3.130 1.050 3.390 1.310 ;
        RECT 4.880 1.070 5.140 1.330 ;
        RECT 5.920 1.060 6.180 1.320 ;
        RECT 1.130 0.500 1.390 0.760 ;
        RECT 4.050 0.500 4.310 0.760 ;
        RECT 2.480 0.130 2.740 0.390 ;
        RECT 5.560 0.140 5.820 0.400 ;
  END
END sky130_hilas_Tgate4Double01

MACRO sky130_hilas_cellAttempt01
  CLASS CORE ;
  FOREIGN sky130_hilas_cellAttempt01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VTUN
    ANTENNADIFFAREA 1.978000 ;
    PORT
      LAYER nwell ;
        RECT 0.010 4.190 1.740 6.050 ;
        RECT 0.000 2.350 1.740 4.190 ;
        RECT 0.010 0.000 1.740 2.350 ;
      LAYER met1 ;
        RECT 0.360 0.000 0.760 6.050 ;
    END
  END VTUN
  PIN VINJ
    ANTENNADIFFAREA 1.020000 ;
    PORT
      LAYER nwell ;
        RECT 7.520 6.040 10.070 6.050 ;
        RECT 7.520 0.020 10.080 6.040 ;
        RECT 7.520 0.010 10.070 0.020 ;
      LAYER met1 ;
        RECT 9.560 5.400 9.720 6.050 ;
        RECT 9.450 4.850 9.720 5.400 ;
        RECT 9.450 4.800 9.730 4.850 ;
        RECT 9.560 4.710 9.730 4.800 ;
        RECT 9.560 4.350 9.720 4.710 ;
        RECT 9.560 4.260 9.730 4.350 ;
        RECT 9.450 4.210 9.730 4.260 ;
        RECT 9.450 3.660 9.720 4.210 ;
        RECT 9.560 2.390 9.720 3.660 ;
        RECT 9.450 1.840 9.720 2.390 ;
        RECT 9.450 1.790 9.730 1.840 ;
        RECT 9.560 1.700 9.730 1.790 ;
        RECT 9.560 1.350 9.720 1.700 ;
        RECT 9.560 1.260 9.730 1.350 ;
        RECT 9.450 1.210 9.730 1.260 ;
        RECT 9.450 0.660 9.720 1.210 ;
        RECT 9.560 0.010 9.720 0.660 ;
    END
  END VINJ
  PIN COLSEL1
    ANTENNAGATEAREA 0.620000 ;
    PORT
      LAYER met1 ;
        RECT 9.120 5.060 9.310 6.050 ;
        RECT 9.140 4.940 9.310 5.060 ;
        RECT 9.150 4.120 9.310 4.940 ;
        RECT 9.140 4.000 9.310 4.120 ;
        RECT 9.120 3.140 9.310 4.000 ;
        RECT 9.100 2.910 9.340 3.140 ;
        RECT 9.120 2.050 9.310 2.910 ;
        RECT 9.140 1.930 9.310 2.050 ;
        RECT 9.150 1.120 9.310 1.930 ;
        RECT 9.140 1.000 9.310 1.120 ;
        RECT 9.120 0.010 9.310 1.000 ;
    END
  END COLSEL1
  PIN COL1
    ANTENNADIFFAREA 0.372000 ;
    PORT
      LAYER met1 ;
        RECT 8.750 5.370 8.910 6.050 ;
        RECT 8.750 5.350 8.950 5.370 ;
        RECT 8.730 5.110 8.960 5.350 ;
        RECT 8.750 4.890 8.950 5.110 ;
        RECT 8.750 4.170 8.910 4.890 ;
        RECT 8.750 3.950 8.950 4.170 ;
        RECT 8.730 3.710 8.960 3.950 ;
        RECT 8.750 3.690 8.950 3.710 ;
        RECT 8.750 2.360 8.910 3.690 ;
        RECT 8.750 2.340 8.950 2.360 ;
        RECT 8.730 2.100 8.960 2.340 ;
        RECT 8.750 1.880 8.950 2.100 ;
        RECT 8.750 1.170 8.910 1.880 ;
        RECT 8.750 0.950 8.950 1.170 ;
        RECT 8.730 0.710 8.960 0.950 ;
        RECT 8.750 0.690 8.950 0.710 ;
        RECT 8.750 0.010 8.910 0.690 ;
    END
  END COL1
  PIN GATE1
    ANTENNADIFFAREA 2.743300 ;
    PORT
      LAYER nwell ;
        RECT 3.760 0.000 5.990 6.050 ;
      LAYER met1 ;
        RECT 4.410 4.130 4.790 6.050 ;
        RECT 4.400 2.270 4.790 4.130 ;
        RECT 4.410 0.000 4.790 2.270 ;
    END
  END GATE1
  PIN DRAIN1
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER met2 ;
        RECT 7.610 5.550 7.920 5.690 ;
        RECT 0.010 5.370 10.080 5.550 ;
        RECT 7.610 5.360 7.920 5.370 ;
    END
  END DRAIN1
  PIN ROW3
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 7.610 2.110 7.920 2.130 ;
        RECT 0.020 1.940 10.080 2.110 ;
        RECT 7.520 1.930 10.080 1.940 ;
        RECT 7.610 1.800 7.920 1.930 ;
    END
  END ROW3
  PIN DRAIN2
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER met2 ;
        RECT 7.610 3.690 7.920 3.700 ;
        RECT 0.000 3.510 10.080 3.690 ;
        RECT 7.610 3.370 7.920 3.510 ;
    END
  END DRAIN2
  PIN ROW2
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 7.610 4.120 7.920 4.250 ;
        RECT 0.000 3.940 10.080 4.120 ;
        RECT 7.610 3.920 7.920 3.940 ;
    END
  END ROW2
  PIN DRAIN3
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER met2 ;
        RECT 7.610 2.540 7.920 2.680 ;
        RECT 7.610 2.530 10.080 2.540 ;
        RECT 0.020 2.360 10.080 2.530 ;
        RECT 7.610 2.350 7.920 2.360 ;
    END
  END DRAIN3
  PIN ROW4
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 7.610 1.130 7.920 1.250 ;
        RECT 0.020 1.120 7.920 1.130 ;
        RECT 0.020 0.960 10.080 1.120 ;
        RECT 0.800 0.870 2.340 0.960 ;
        RECT 7.520 0.940 10.080 0.960 ;
        RECT 7.610 0.920 7.920 0.940 ;
    END
  END ROW4
  PIN DRAIN4
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER met2 ;
        RECT 7.610 0.690 7.920 0.700 ;
        RECT 0.020 0.520 10.080 0.690 ;
        RECT 7.610 0.510 10.080 0.520 ;
        RECT 7.610 0.370 7.920 0.510 ;
    END
  END DRAIN4
  PIN ROW1
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 7.610 5.120 7.920 5.140 ;
        RECT 0.010 4.940 10.080 5.120 ;
        RECT 7.610 4.810 7.920 4.940 ;
    END
  END ROW1
  PIN VGND
    ANTENNADIFFAREA 1.012300 ;
    PORT
      LAYER met2 ;
        RECT 2.760 1.560 3.080 1.570 ;
        RECT 6.690 1.560 7.010 1.640 ;
        RECT 2.760 1.380 7.010 1.560 ;
        RECT 2.760 1.310 3.080 1.380 ;
        RECT 6.690 1.320 7.010 1.380 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.730 4.890 6.970 6.050 ;
        RECT 6.710 4.230 6.980 4.890 ;
        RECT 6.730 1.640 6.970 4.230 ;
        RECT 6.720 1.320 6.980 1.640 ;
        RECT 6.730 0.000 6.970 1.320 ;
      LAYER via ;
        RECT 6.720 1.350 6.980 1.610 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.800 4.870 3.040 6.050 ;
        RECT 2.790 4.210 3.050 4.870 ;
        RECT 2.800 1.600 3.040 4.210 ;
        RECT 2.790 1.280 3.050 1.600 ;
        RECT 2.800 0.000 3.040 1.280 ;
      LAYER via ;
        RECT 2.790 1.310 3.050 1.570 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 7.620 5.640 7.940 5.650 ;
        RECT 7.620 5.470 8.200 5.640 ;
        RECT 7.620 5.420 7.950 5.470 ;
        RECT 7.620 5.390 7.940 5.420 ;
        RECT 9.480 5.370 9.680 5.720 ;
        RECT 7.620 5.060 7.940 5.100 ;
        RECT 7.620 5.020 7.950 5.060 ;
        RECT 7.620 4.850 8.200 5.020 ;
        RECT 7.620 4.840 7.940 4.850 ;
        RECT 2.830 4.300 3.000 4.810 ;
        RECT 6.770 4.290 6.940 4.800 ;
        RECT 8.750 4.780 8.950 5.350 ;
        RECT 9.480 5.340 9.690 5.370 ;
        RECT 9.470 4.750 9.690 5.340 ;
        RECT 7.620 4.210 7.940 4.220 ;
        RECT 7.620 4.040 8.200 4.210 ;
        RECT 7.620 4.000 7.950 4.040 ;
        RECT 7.620 3.960 7.940 4.000 ;
        RECT 8.750 3.710 8.950 4.280 ;
        RECT 9.470 3.720 9.690 4.310 ;
        RECT 9.480 3.690 9.690 3.720 ;
        RECT 7.620 3.640 7.940 3.670 ;
        RECT 0.430 2.800 0.980 3.230 ;
        RECT 2.840 2.590 3.010 3.600 ;
        RECT 7.620 3.590 7.950 3.640 ;
        RECT 4.460 2.730 5.010 3.160 ;
        RECT 6.770 2.450 6.940 3.460 ;
        RECT 7.620 3.420 8.200 3.590 ;
        RECT 7.620 3.410 7.940 3.420 ;
        RECT 9.480 3.340 9.680 3.690 ;
        RECT 8.870 2.940 9.310 3.110 ;
        RECT 7.620 2.630 7.940 2.640 ;
        RECT 7.620 2.460 8.200 2.630 ;
        RECT 7.620 2.410 7.950 2.460 ;
        RECT 7.620 2.380 7.940 2.410 ;
        RECT 9.480 2.360 9.680 2.710 ;
        RECT 7.620 2.050 7.940 2.090 ;
        RECT 7.620 2.010 7.950 2.050 ;
        RECT 7.620 1.840 8.200 2.010 ;
        RECT 7.620 1.830 7.940 1.840 ;
        RECT 8.750 1.770 8.950 2.340 ;
        RECT 9.480 2.330 9.690 2.360 ;
        RECT 9.470 1.740 9.690 2.330 ;
        RECT 7.620 1.210 7.940 1.220 ;
        RECT 7.620 1.040 8.200 1.210 ;
        RECT 7.620 1.000 7.950 1.040 ;
        RECT 7.620 0.960 7.940 1.000 ;
        RECT 8.750 0.710 8.950 1.280 ;
        RECT 9.470 0.720 9.690 1.310 ;
        RECT 9.480 0.690 9.690 0.720 ;
        RECT 7.620 0.640 7.940 0.670 ;
        RECT 7.620 0.590 7.950 0.640 ;
        RECT 7.620 0.420 8.200 0.590 ;
        RECT 7.620 0.410 7.940 0.420 ;
        RECT 9.480 0.340 9.680 0.690 ;
      LAYER mcon ;
        RECT 7.680 5.430 7.850 5.600 ;
        RECT 8.760 5.140 8.930 5.310 ;
        RECT 7.680 4.880 7.850 5.050 ;
        RECT 2.830 4.640 3.000 4.810 ;
        RECT 6.770 4.630 6.940 4.800 ;
        RECT 9.490 5.170 9.660 5.340 ;
        RECT 7.680 4.010 7.850 4.180 ;
        RECT 8.760 3.750 8.930 3.920 ;
        RECT 9.490 3.720 9.660 3.890 ;
        RECT 7.680 3.460 7.850 3.630 ;
        RECT 0.430 2.880 0.700 3.150 ;
        RECT 2.840 3.180 3.010 3.350 ;
        RECT 2.840 2.840 3.010 3.010 ;
        RECT 4.460 2.810 4.730 3.080 ;
        RECT 6.770 3.040 6.940 3.210 ;
        RECT 9.130 2.940 9.310 3.110 ;
        RECT 6.770 2.700 6.940 2.870 ;
        RECT 7.680 2.420 7.850 2.590 ;
        RECT 8.760 2.130 8.930 2.300 ;
        RECT 7.680 1.870 7.850 2.040 ;
        RECT 9.490 2.160 9.660 2.330 ;
        RECT 7.680 1.010 7.850 1.180 ;
        RECT 8.760 0.750 8.930 0.920 ;
        RECT 9.490 0.720 9.660 0.890 ;
        RECT 7.680 0.460 7.850 0.630 ;
      LAYER met1 ;
        RECT 7.610 5.360 7.930 5.680 ;
        RECT 7.610 4.810 7.930 5.130 ;
        RECT 7.610 3.930 7.930 4.250 ;
        RECT 7.610 3.380 7.930 3.700 ;
        RECT 7.610 2.350 7.930 2.670 ;
        RECT 7.610 1.800 7.930 2.120 ;
        RECT 7.610 0.930 7.930 1.250 ;
        RECT 7.610 0.380 7.930 0.700 ;
      LAYER via ;
        RECT 7.640 5.390 7.900 5.650 ;
        RECT 7.640 4.840 7.900 5.100 ;
        RECT 7.640 3.960 7.900 4.220 ;
        RECT 7.640 3.410 7.900 3.670 ;
        RECT 7.640 2.380 7.900 2.640 ;
        RECT 7.640 1.830 7.900 2.090 ;
        RECT 7.640 0.960 7.900 1.220 ;
        RECT 7.640 0.410 7.900 0.670 ;
  END
END sky130_hilas_cellAttempt01

MACRO sky130_hilas_StepUpDigital
  CLASS CORE ;
  FOREIGN sky130_hilas_StepUpDigital ;
  ORIGIN 0.000 0.800 ;
  SIZE 8.800 BY 1.590 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 0.000 -0.800 2.510 0.790 ;
        RECT 6.470 -0.800 8.240 0.790 ;
      LAYER li1 ;
        RECT 1.280 0.400 3.510 0.550 ;
        RECT 0.340 0.220 0.670 0.390 ;
        RECT 1.130 0.380 3.510 0.400 ;
        RECT 1.130 0.230 1.730 0.380 ;
        RECT 3.330 0.370 3.510 0.380 ;
        RECT 3.330 0.350 3.970 0.370 ;
        RECT 0.410 -0.240 0.590 0.220 ;
        RECT 2.060 0.030 2.390 0.200 ;
        RECT 3.330 0.180 4.010 0.350 ;
        RECT 4.460 0.320 4.920 0.350 ;
        RECT 6.230 0.320 6.580 0.420 ;
        RECT 4.460 0.180 5.570 0.320 ;
        RECT 3.330 0.120 3.510 0.180 ;
        RECT 4.750 0.150 5.570 0.180 ;
        RECT 5.810 0.150 6.980 0.320 ;
        RECT 7.230 0.150 7.990 0.320 ;
        RECT 2.060 -0.220 2.310 0.030 ;
        RECT 4.750 0.010 5.010 0.150 ;
        RECT 0.410 -0.410 1.370 -0.240 ;
        RECT 1.840 -0.320 2.310 -0.220 ;
        RECT 3.830 -0.160 5.010 0.010 ;
        RECT 7.760 0.140 7.990 0.150 ;
        RECT 1.840 -0.330 2.480 -0.320 ;
        RECT 1.840 -0.390 3.280 -0.330 ;
        RECT 1.920 -0.500 3.280 -0.390 ;
        RECT 3.830 -0.600 4.010 -0.160 ;
        RECT 4.750 -0.300 5.010 -0.160 ;
        RECT 6.220 -0.300 6.550 -0.040 ;
        RECT 7.760 -0.300 8.030 0.140 ;
        RECT 4.250 -0.660 4.460 -0.330 ;
        RECT 4.750 -0.470 5.080 -0.300 ;
        RECT 5.320 -0.470 7.480 -0.300 ;
        RECT 4.750 -0.520 4.920 -0.470 ;
        RECT 7.730 -0.480 8.060 -0.300 ;
        RECT 8.410 -0.440 8.580 -0.380 ;
        RECT 8.390 -0.660 8.610 -0.440 ;
        RECT 8.410 -0.710 8.580 -0.660 ;
      LAYER mcon ;
        RECT 1.450 0.300 1.620 0.470 ;
        RECT 0.410 -0.050 0.580 0.120 ;
        RECT 6.290 0.190 6.500 0.400 ;
        RECT 0.410 -0.400 0.580 -0.230 ;
        RECT 7.800 -0.180 7.970 -0.010 ;
      LAYER met1 ;
        RECT 0.340 -0.800 0.630 0.790 ;
        RECT 1.380 0.250 1.700 0.550 ;
        RECT 4.220 -0.600 4.500 -0.270 ;
        RECT 4.750 -0.800 5.060 0.790 ;
        RECT 6.230 0.150 6.580 0.440 ;
        RECT 6.380 0.130 6.580 0.150 ;
        RECT 7.760 -0.800 8.000 0.790 ;
        RECT 8.330 -0.710 8.740 -0.380 ;
      LAYER via ;
        RECT 1.410 0.260 1.670 0.520 ;
        RECT 4.230 -0.560 4.490 -0.300 ;
        RECT 6.270 0.160 6.530 0.420 ;
        RECT 8.370 -0.680 8.630 -0.420 ;
      LAYER met2 ;
        RECT 1.380 0.470 1.700 0.520 ;
        RECT 0.070 0.270 1.700 0.470 ;
        RECT 1.380 0.260 1.700 0.270 ;
        RECT 4.190 -0.350 4.530 -0.290 ;
        RECT 6.270 -0.350 6.530 0.450 ;
        RECT 4.190 -0.570 6.630 -0.350 ;
        RECT 8.340 -0.710 8.800 -0.390 ;
  END
END sky130_hilas_StepUpDigital

MACRO sky130_hilas_VinjNOR3
  CLASS CORE ;
  FOREIGN sky130_hilas_VinjNOR3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.880 BY 1.640 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 0.010 0.000 3.450 1.640 ;
      LAYER li1 ;
        RECT 0.630 1.210 0.800 1.350 ;
        RECT 1.360 1.230 1.530 1.310 ;
        RECT 2.170 1.230 2.340 1.310 ;
        RECT 3.710 1.270 3.880 1.390 ;
        RECT 0.630 1.040 0.820 1.210 ;
        RECT 0.630 0.940 0.800 1.040 ;
        RECT 1.360 0.660 1.570 1.230 ;
        RECT 2.130 0.980 2.340 1.230 ;
        RECT 2.730 1.050 2.900 1.150 ;
        RECT 3.670 1.100 3.880 1.270 ;
        RECT 5.600 1.200 5.860 1.270 ;
        RECT 6.400 1.200 6.580 1.330 ;
        RECT 3.710 1.060 3.880 1.100 ;
        RECT 2.130 0.660 2.300 0.980 ;
        RECT 2.700 0.880 2.900 1.050 ;
        RECT 2.730 0.780 2.900 0.880 ;
        RECT 4.270 1.020 5.140 1.190 ;
        RECT 5.600 1.020 6.580 1.200 ;
        RECT 0.200 0.560 0.370 0.660 ;
        RECT 0.180 0.390 0.370 0.560 ;
        RECT 0.200 0.330 0.370 0.390 ;
        RECT 0.620 0.600 0.790 0.660 ;
        RECT 0.620 0.330 0.870 0.600 ;
        RECT 1.360 0.410 1.610 0.660 ;
        RECT 0.630 0.310 0.870 0.330 ;
        RECT 1.440 0.320 1.610 0.410 ;
        RECT 2.090 0.410 2.300 0.660 ;
        RECT 4.270 0.580 4.440 1.020 ;
        RECT 5.600 0.580 5.860 1.020 ;
        RECT 6.400 0.910 6.580 1.020 ;
        RECT 2.810 0.410 4.440 0.580 ;
        RECT 4.890 0.410 5.860 0.580 ;
        RECT 6.310 0.410 6.650 0.580 ;
        RECT 2.090 0.330 2.260 0.410 ;
        RECT 3.580 0.370 3.750 0.410 ;
      LAYER mcon ;
        RECT 0.650 1.040 0.820 1.210 ;
        RECT 0.660 0.360 0.830 0.530 ;
        RECT 5.630 0.700 5.810 0.880 ;
      LAYER met1 ;
        RECT 0.620 1.260 0.840 1.600 ;
        RECT 0.620 1.000 0.850 1.260 ;
        RECT 0.090 0.320 0.400 0.670 ;
        RECT 0.620 0.600 0.840 1.000 ;
        RECT 2.640 0.840 2.970 1.100 ;
        RECT 3.610 1.060 4.040 1.350 ;
        RECT 0.620 0.290 0.870 0.600 ;
        RECT 3.480 0.310 3.870 0.580 ;
        RECT 0.620 0.090 0.840 0.290 ;
        RECT 5.590 0.090 5.860 1.610 ;
        RECT 6.410 0.320 6.720 0.640 ;
      LAYER via ;
        RECT 0.120 0.350 0.380 0.610 ;
        RECT 2.680 0.840 2.940 1.100 ;
        RECT 3.670 1.090 3.930 1.350 ;
        RECT 3.540 0.310 3.800 0.570 ;
        RECT 6.440 0.350 6.700 0.610 ;
      LAYER met2 ;
        RECT 0.000 1.290 4.040 1.450 ;
        RECT 2.640 1.020 2.970 1.100 ;
        RECT 3.620 1.060 4.040 1.290 ;
        RECT 2.370 1.000 2.970 1.020 ;
        RECT 0.010 0.840 2.970 1.000 ;
        RECT 0.090 0.510 0.410 0.610 ;
        RECT 0.010 0.350 0.410 0.510 ;
        RECT 3.500 0.490 3.870 0.570 ;
        RECT 3.500 0.480 4.530 0.490 ;
        RECT 6.410 0.480 6.720 0.640 ;
        RECT 3.500 0.310 6.880 0.480 ;
  END
END sky130_hilas_VinjNOR3

MACRO sky130_hilas_VinjDiodeProtect01
  CLASS CORE ;
  FOREIGN sky130_hilas_VinjDiodeProtect01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.590 BY 10.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN OUTPUT 
    ANTENNADIFFAREA 58.900799 ;
    PORT
      LAYER met1 ;
        RECT 14.350 10.250 14.700 10.400 ;
        RECT 14.340 9.300 14.710 10.250 ;
        RECT 12.560 8.930 16.460 9.300 ;
        RECT 12.550 7.470 16.460 8.930 ;
        RECT 2.840 7.460 16.460 7.470 ;
        RECT 2.170 6.900 16.460 7.460 ;
        RECT 2.170 2.600 25.520 6.900 ;
        RECT 2.170 2.320 16.460 2.600 ;
        RECT 12.550 0.770 16.460 2.320 ;
        RECT 12.530 0.000 16.480 0.770 ;
    END
  END OUTPUT 
  PIN VGND
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met2 ;
        RECT 0.000 7.380 28.590 8.780 ;
        RECT 0.470 7.370 1.400 7.380 ;
        RECT 0.720 6.260 0.890 7.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.440 8.130 2.810 8.760 ;
        RECT 23.780 8.280 27.910 8.680 ;
        RECT 23.780 8.190 27.920 8.280 ;
        RECT 0.470 6.170 1.420 8.130 ;
        RECT 2.170 8.110 2.750 8.130 ;
        RECT 27.390 7.290 27.920 8.190 ;
        RECT 0.700 0.500 1.420 6.170 ;
      LAYER via ;
        RECT 0.660 8.280 2.690 8.610 ;
        RECT 24.050 8.280 27.040 8.630 ;
        RECT 0.600 7.420 1.300 8.040 ;
        RECT 27.480 7.480 27.830 8.240 ;
    END
  END VGND
  PIN VINJ
    ANTENNADIFFAREA 9.088799 ;
    PORT
      LAYER nwell ;
        RECT 14.870 1.910 26.920 7.850 ;
      LAYER met2 ;
        RECT 26.340 2.480 26.980 5.490 ;
        RECT 0.000 1.080 28.590 2.480 ;
        RECT 25.440 0.950 28.070 1.080 ;
        RECT 25.440 0.440 27.990 0.950 ;
        RECT 25.440 0.370 26.060 0.440 ;
    END
  END VINJ
  PIN INPUT
    PORT
      LAYER met1 ;
        RECT 7.710 10.280 11.610 10.870 ;
        RECT 7.710 8.930 8.000 10.280 ;
    END
  END INPUT
  OBS
      LAYER li1 ;
        RECT 7.730 8.930 7.980 10.390 ;
        RECT 7.770 8.920 7.940 8.930 ;
        RECT 14.410 8.900 14.660 10.370 ;
        RECT 0.550 8.180 27.930 8.690 ;
        RECT 0.550 6.250 1.350 8.180 ;
        RECT 1.930 7.730 2.100 7.810 ;
        RECT 13.170 7.730 13.400 7.820 ;
        RECT 1.930 7.720 13.400 7.730 ;
        RECT 0.550 1.670 1.060 6.250 ;
        RECT 1.920 2.250 13.400 7.720 ;
        RECT 1.850 2.080 13.400 2.250 ;
        RECT 1.920 2.020 2.110 2.080 ;
        RECT 13.170 1.840 13.400 2.080 ;
        RECT 1.800 1.670 3.600 1.680 ;
        RECT 13.960 1.670 14.470 8.180 ;
        RECT 15.230 7.290 26.480 7.460 ;
        RECT 15.230 2.420 15.400 7.290 ;
        RECT 15.790 6.960 25.900 6.980 ;
        RECT 15.790 6.920 25.920 6.960 ;
        RECT 15.740 6.750 25.920 6.920 ;
        RECT 15.790 2.730 25.920 6.750 ;
        RECT 26.310 5.530 26.480 7.290 ;
        RECT 15.790 2.650 25.900 2.730 ;
        RECT 15.220 2.350 15.400 2.420 ;
        RECT 26.310 2.350 26.920 5.530 ;
        RECT 15.220 2.180 26.920 2.350 ;
        RECT 26.380 2.070 26.920 2.180 ;
        RECT 27.380 1.830 27.930 8.180 ;
        RECT 27.370 1.670 27.930 1.830 ;
        RECT 0.550 1.330 27.930 1.670 ;
        RECT 0.580 1.160 27.930 1.330 ;
        RECT 0.580 1.140 1.270 1.160 ;
        RECT 1.780 1.150 3.580 1.160 ;
      LAYER mcon ;
        RECT 7.770 10.190 7.940 10.360 ;
        RECT 7.770 9.850 7.940 10.020 ;
        RECT 7.770 9.510 7.940 9.680 ;
        RECT 7.770 9.170 7.940 9.340 ;
        RECT 14.450 10.170 14.620 10.340 ;
        RECT 14.450 9.830 14.620 10.000 ;
        RECT 14.450 9.490 14.620 9.660 ;
        RECT 14.450 9.150 14.620 9.320 ;
        RECT 0.630 8.520 2.490 8.530 ;
        RECT 0.630 8.350 2.500 8.520 ;
        RECT 23.990 8.340 27.150 8.520 ;
        RECT 0.710 7.390 0.890 8.180 ;
        RECT 0.720 6.260 0.890 7.390 ;
        RECT 1.070 6.250 1.250 8.170 ;
        RECT 2.260 7.220 13.240 7.390 ;
        RECT 2.260 6.600 13.240 6.770 ;
        RECT 2.270 5.980 13.250 6.150 ;
        RECT 2.290 5.400 13.270 5.570 ;
        RECT 2.300 4.810 13.280 4.980 ;
        RECT 2.300 4.210 13.280 4.380 ;
        RECT 2.250 3.610 13.230 3.780 ;
        RECT 2.260 3.000 13.240 3.170 ;
        RECT 2.250 2.400 13.230 2.570 ;
        RECT 15.990 6.460 25.440 6.630 ;
        RECT 15.980 5.710 25.370 5.880 ;
        RECT 16.010 4.990 25.410 5.160 ;
        RECT 16.020 4.330 25.390 4.500 ;
        RECT 16.010 3.680 25.460 3.850 ;
        RECT 16.020 3.040 25.410 3.210 ;
        RECT 27.560 7.360 27.760 8.290 ;
        RECT 26.490 2.120 26.840 5.420 ;
      LAYER met1 ;
        RECT 26.290 5.480 26.860 5.490 ;
        RECT 26.290 2.060 26.910 5.480 ;
        RECT 26.290 2.050 26.860 2.060 ;
        RECT 25.460 0.420 26.020 0.920 ;
        RECT 25.470 0.200 26.020 0.420 ;
      LAYER via ;
        RECT 26.450 2.190 26.870 5.360 ;
        RECT 25.480 0.370 26.000 0.890 ;
  END
END sky130_hilas_VinjDiodeProtect01

MACRO sky130_hilas_LevelShift4InputUp
  CLASS CORE ;
  FOREIGN sky130_hilas_LevelShift4InputUp ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.040 BY 6.730 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN INPUT1
    PORT
      LAYER met2 ;
        RECT 8.900 5.140 8.990 5.460 ;
    END
  END INPUT1
  PIN INPUT2
    PORT
      LAYER met2 ;
        RECT 8.900 3.590 8.990 3.910 ;
    END
  END INPUT2
  PIN INPUT3
    PORT
      LAYER met2 ;
        RECT 8.900 2.040 8.990 2.360 ;
    END
  END INPUT3
  PIN INPUT4
    PORT
      LAYER met2 ;
        RECT 8.900 0.490 8.990 0.810 ;
    END
  END INPUT4
  PIN VPWR
    PORT
      LAYER met1 ;
        RECT 7.950 6.590 8.190 6.640 ;
    END
    PORT
      LAYER nwell ;
        RECT 6.470 0.000 8.240 6.240 ;
      LAYER met1 ;
        RECT 7.760 0.450 8.000 6.240 ;
        RECT 7.760 0.400 8.190 0.450 ;
        RECT 7.760 0.000 8.000 0.400 ;
    END
  END VPWR
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 0.530 6.590 0.820 6.640 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.000 0.000 2.510 6.240 ;
      LAYER met1 ;
        RECT 0.340 0.450 0.630 6.240 ;
        RECT 0.340 0.400 0.820 0.450 ;
        RECT 0.340 0.000 0.630 0.400 ;
    END
  END VINJ
  PIN OUTPUT1
    PORT
      LAYER met2 ;
        RECT 0.190 6.120 0.300 6.320 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    PORT
      LAYER met2 ;
        RECT 0.190 4.570 0.300 4.770 ;
    END
  END OUTPUT2
  PIN OUTPUT3
    PORT
      LAYER met2 ;
        RECT 0.190 3.020 0.300 3.220 ;
    END
  END OUTPUT3
  PIN OUTPUT4
    PORT
      LAYER met2 ;
        RECT 0.190 1.470 0.300 1.670 ;
    END
  END OUTPUT4
  PIN VGND
    PORT
      LAYER met1 ;
        RECT 4.940 6.570 5.250 6.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.750 0.460 5.060 6.240 ;
        RECT 4.750 0.400 5.250 0.460 ;
        RECT 4.750 0.000 5.060 0.400 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.280 5.850 3.510 6.000 ;
        RECT 0.340 5.670 0.670 5.840 ;
        RECT 1.130 5.830 3.510 5.850 ;
        RECT 1.130 5.680 1.730 5.830 ;
        RECT 3.330 5.820 3.510 5.830 ;
        RECT 3.330 5.800 3.970 5.820 ;
        RECT 0.410 5.210 0.590 5.670 ;
        RECT 2.060 5.480 2.390 5.650 ;
        RECT 3.330 5.630 4.010 5.800 ;
        RECT 4.460 5.770 4.920 5.800 ;
        RECT 6.230 5.770 6.580 5.870 ;
        RECT 4.460 5.630 5.570 5.770 ;
        RECT 3.330 5.570 3.510 5.630 ;
        RECT 4.750 5.600 5.570 5.630 ;
        RECT 5.810 5.600 6.980 5.770 ;
        RECT 7.230 5.600 7.990 5.770 ;
        RECT 2.060 5.230 2.310 5.480 ;
        RECT 4.750 5.460 5.010 5.600 ;
        RECT 0.410 5.040 1.370 5.210 ;
        RECT 1.840 5.130 2.310 5.230 ;
        RECT 3.830 5.290 5.010 5.460 ;
        RECT 7.760 5.590 7.990 5.600 ;
        RECT 1.840 5.120 2.480 5.130 ;
        RECT 1.840 5.060 3.280 5.120 ;
        RECT 1.920 4.950 3.280 5.060 ;
        RECT 3.830 4.850 4.010 5.290 ;
        RECT 4.750 5.150 5.010 5.290 ;
        RECT 6.220 5.150 6.550 5.410 ;
        RECT 7.760 5.150 8.030 5.590 ;
        RECT 4.250 4.790 4.460 5.120 ;
        RECT 4.750 4.980 5.080 5.150 ;
        RECT 5.320 4.980 7.480 5.150 ;
        RECT 4.750 4.930 4.920 4.980 ;
        RECT 7.730 4.970 8.060 5.150 ;
        RECT 8.410 5.010 8.580 5.070 ;
        RECT 8.390 4.790 8.610 5.010 ;
        RECT 8.410 4.740 8.580 4.790 ;
        RECT 1.280 4.300 3.510 4.450 ;
        RECT 0.340 4.120 0.670 4.290 ;
        RECT 1.130 4.280 3.510 4.300 ;
        RECT 1.130 4.130 1.730 4.280 ;
        RECT 3.330 4.270 3.510 4.280 ;
        RECT 3.330 4.250 3.970 4.270 ;
        RECT 0.410 3.660 0.590 4.120 ;
        RECT 2.060 3.930 2.390 4.100 ;
        RECT 3.330 4.080 4.010 4.250 ;
        RECT 4.460 4.220 4.920 4.250 ;
        RECT 6.230 4.220 6.580 4.320 ;
        RECT 4.460 4.080 5.570 4.220 ;
        RECT 3.330 4.020 3.510 4.080 ;
        RECT 4.750 4.050 5.570 4.080 ;
        RECT 5.810 4.050 6.980 4.220 ;
        RECT 7.230 4.050 7.990 4.220 ;
        RECT 2.060 3.680 2.310 3.930 ;
        RECT 4.750 3.910 5.010 4.050 ;
        RECT 0.410 3.490 1.370 3.660 ;
        RECT 1.840 3.580 2.310 3.680 ;
        RECT 3.830 3.740 5.010 3.910 ;
        RECT 7.760 4.040 7.990 4.050 ;
        RECT 1.840 3.570 2.480 3.580 ;
        RECT 1.840 3.510 3.280 3.570 ;
        RECT 1.920 3.400 3.280 3.510 ;
        RECT 3.830 3.300 4.010 3.740 ;
        RECT 4.750 3.600 5.010 3.740 ;
        RECT 6.220 3.600 6.550 3.860 ;
        RECT 7.760 3.600 8.030 4.040 ;
        RECT 4.250 3.240 4.460 3.570 ;
        RECT 4.750 3.430 5.080 3.600 ;
        RECT 5.320 3.430 7.480 3.600 ;
        RECT 4.750 3.380 4.920 3.430 ;
        RECT 7.730 3.420 8.060 3.600 ;
        RECT 8.410 3.460 8.580 3.520 ;
        RECT 8.390 3.240 8.610 3.460 ;
        RECT 8.410 3.190 8.580 3.240 ;
        RECT 1.280 2.750 3.510 2.900 ;
        RECT 0.340 2.570 0.670 2.740 ;
        RECT 1.130 2.730 3.510 2.750 ;
        RECT 1.130 2.580 1.730 2.730 ;
        RECT 3.330 2.720 3.510 2.730 ;
        RECT 3.330 2.700 3.970 2.720 ;
        RECT 0.410 2.110 0.590 2.570 ;
        RECT 2.060 2.380 2.390 2.550 ;
        RECT 3.330 2.530 4.010 2.700 ;
        RECT 4.460 2.670 4.920 2.700 ;
        RECT 6.230 2.670 6.580 2.770 ;
        RECT 4.460 2.530 5.570 2.670 ;
        RECT 3.330 2.470 3.510 2.530 ;
        RECT 4.750 2.500 5.570 2.530 ;
        RECT 5.810 2.500 6.980 2.670 ;
        RECT 7.230 2.500 7.990 2.670 ;
        RECT 2.060 2.130 2.310 2.380 ;
        RECT 4.750 2.360 5.010 2.500 ;
        RECT 0.410 1.940 1.370 2.110 ;
        RECT 1.840 2.030 2.310 2.130 ;
        RECT 3.830 2.190 5.010 2.360 ;
        RECT 7.760 2.490 7.990 2.500 ;
        RECT 1.840 2.020 2.480 2.030 ;
        RECT 1.840 1.960 3.280 2.020 ;
        RECT 1.920 1.850 3.280 1.960 ;
        RECT 3.830 1.750 4.010 2.190 ;
        RECT 4.750 2.050 5.010 2.190 ;
        RECT 6.220 2.050 6.550 2.310 ;
        RECT 7.760 2.050 8.030 2.490 ;
        RECT 4.250 1.690 4.460 2.020 ;
        RECT 4.750 1.880 5.080 2.050 ;
        RECT 5.320 1.880 7.480 2.050 ;
        RECT 4.750 1.830 4.920 1.880 ;
        RECT 7.730 1.870 8.060 2.050 ;
        RECT 8.410 1.910 8.580 1.970 ;
        RECT 8.390 1.690 8.610 1.910 ;
        RECT 8.410 1.640 8.580 1.690 ;
        RECT 1.280 1.200 3.510 1.350 ;
        RECT 0.340 1.020 0.670 1.190 ;
        RECT 1.130 1.180 3.510 1.200 ;
        RECT 1.130 1.030 1.730 1.180 ;
        RECT 3.330 1.170 3.510 1.180 ;
        RECT 3.330 1.150 3.970 1.170 ;
        RECT 0.410 0.560 0.590 1.020 ;
        RECT 2.060 0.830 2.390 1.000 ;
        RECT 3.330 0.980 4.010 1.150 ;
        RECT 4.460 1.120 4.920 1.150 ;
        RECT 6.230 1.120 6.580 1.220 ;
        RECT 4.460 0.980 5.570 1.120 ;
        RECT 3.330 0.920 3.510 0.980 ;
        RECT 4.750 0.950 5.570 0.980 ;
        RECT 5.810 0.950 6.980 1.120 ;
        RECT 7.230 0.950 7.990 1.120 ;
        RECT 2.060 0.580 2.310 0.830 ;
        RECT 4.750 0.810 5.010 0.950 ;
        RECT 0.410 0.390 1.370 0.560 ;
        RECT 1.840 0.480 2.310 0.580 ;
        RECT 3.830 0.640 5.010 0.810 ;
        RECT 7.760 0.940 7.990 0.950 ;
        RECT 1.840 0.470 2.480 0.480 ;
        RECT 1.840 0.410 3.280 0.470 ;
        RECT 1.920 0.300 3.280 0.410 ;
        RECT 3.830 0.200 4.010 0.640 ;
        RECT 4.750 0.500 5.010 0.640 ;
        RECT 6.220 0.500 6.550 0.760 ;
        RECT 7.760 0.500 8.030 0.940 ;
        RECT 4.250 0.140 4.460 0.470 ;
        RECT 4.750 0.330 5.080 0.500 ;
        RECT 5.320 0.330 7.480 0.500 ;
        RECT 4.750 0.280 4.920 0.330 ;
        RECT 7.730 0.320 8.060 0.500 ;
        RECT 8.410 0.360 8.580 0.420 ;
        RECT 8.390 0.140 8.610 0.360 ;
        RECT 8.410 0.090 8.580 0.140 ;
      LAYER mcon ;
        RECT 1.450 5.750 1.620 5.920 ;
        RECT 0.410 5.400 0.580 5.570 ;
        RECT 6.290 5.640 6.500 5.850 ;
        RECT 0.410 5.050 0.580 5.220 ;
        RECT 7.800 5.270 7.970 5.440 ;
        RECT 1.450 4.200 1.620 4.370 ;
        RECT 0.410 3.850 0.580 4.020 ;
        RECT 6.290 4.090 6.500 4.300 ;
        RECT 0.410 3.500 0.580 3.670 ;
        RECT 7.800 3.720 7.970 3.890 ;
        RECT 1.450 2.650 1.620 2.820 ;
        RECT 0.410 2.300 0.580 2.470 ;
        RECT 6.290 2.540 6.500 2.750 ;
        RECT 0.410 1.950 0.580 2.120 ;
        RECT 7.800 2.170 7.970 2.340 ;
        RECT 1.450 1.100 1.620 1.270 ;
        RECT 0.410 0.750 0.580 0.920 ;
        RECT 6.290 0.990 6.500 1.200 ;
        RECT 0.410 0.400 0.580 0.570 ;
        RECT 7.800 0.620 7.970 0.790 ;
      LAYER met1 ;
        RECT 1.380 5.700 1.700 6.000 ;
        RECT 6.230 5.600 6.580 5.890 ;
        RECT 6.380 5.580 6.580 5.600 ;
        RECT 4.220 4.850 4.500 5.180 ;
        RECT 8.330 4.740 8.740 5.070 ;
        RECT 1.380 4.150 1.700 4.450 ;
        RECT 6.230 4.050 6.580 4.340 ;
        RECT 6.380 4.030 6.580 4.050 ;
        RECT 4.220 3.300 4.500 3.630 ;
        RECT 8.330 3.190 8.740 3.520 ;
        RECT 1.380 2.600 1.700 2.900 ;
        RECT 6.230 2.500 6.580 2.790 ;
        RECT 6.380 2.480 6.580 2.500 ;
        RECT 4.220 1.750 4.500 2.080 ;
        RECT 8.330 1.640 8.740 1.970 ;
        RECT 1.380 1.050 1.700 1.350 ;
        RECT 6.230 0.950 6.580 1.240 ;
        RECT 6.380 0.930 6.580 0.950 ;
        RECT 4.220 0.200 4.500 0.530 ;
        RECT 8.330 0.090 8.740 0.420 ;
      LAYER via ;
        RECT 1.410 5.710 1.670 5.970 ;
        RECT 6.270 5.610 6.530 5.870 ;
        RECT 4.230 4.890 4.490 5.150 ;
        RECT 8.370 4.770 8.630 5.030 ;
        RECT 1.410 4.160 1.670 4.420 ;
        RECT 6.270 4.060 6.530 4.320 ;
        RECT 4.230 3.340 4.490 3.600 ;
        RECT 8.370 3.220 8.630 3.480 ;
        RECT 1.410 2.610 1.670 2.870 ;
        RECT 6.270 2.510 6.530 2.770 ;
        RECT 4.230 1.790 4.490 2.050 ;
        RECT 8.370 1.670 8.630 1.930 ;
        RECT 1.410 1.060 1.670 1.320 ;
        RECT 6.270 0.960 6.530 1.220 ;
        RECT 4.230 0.240 4.490 0.500 ;
        RECT 8.370 0.120 8.630 0.380 ;
      LAYER met2 ;
        RECT 1.380 5.920 1.700 5.970 ;
        RECT 0.070 5.720 1.700 5.920 ;
        RECT 1.380 5.710 1.700 5.720 ;
        RECT 4.190 5.100 4.530 5.160 ;
        RECT 6.270 5.100 6.530 5.900 ;
        RECT 4.190 4.880 6.630 5.100 ;
        RECT 8.340 4.740 8.800 5.060 ;
        RECT 1.380 4.370 1.700 4.420 ;
        RECT 0.070 4.170 1.700 4.370 ;
        RECT 1.380 4.160 1.700 4.170 ;
        RECT 4.190 3.550 4.530 3.610 ;
        RECT 6.270 3.550 6.530 4.350 ;
        RECT 4.190 3.330 6.630 3.550 ;
        RECT 8.340 3.190 8.800 3.510 ;
        RECT 1.380 2.820 1.700 2.870 ;
        RECT 0.070 2.620 1.700 2.820 ;
        RECT 1.380 2.610 1.700 2.620 ;
        RECT 4.190 2.000 4.530 2.060 ;
        RECT 6.270 2.000 6.530 2.800 ;
        RECT 4.190 1.780 6.630 2.000 ;
        RECT 8.340 1.640 8.800 1.960 ;
        RECT 1.380 1.270 1.700 1.320 ;
        RECT 0.070 1.070 1.700 1.270 ;
        RECT 1.380 1.060 1.700 1.070 ;
        RECT 4.190 0.450 4.530 0.510 ;
        RECT 6.270 0.450 6.530 1.250 ;
        RECT 4.190 0.230 6.630 0.450 ;
        RECT 8.340 0.090 8.800 0.410 ;
  END
END sky130_hilas_LevelShift4InputUp

MACRO sky130_hilas_WTA4Stage01
  CLASS CORE ;
  FOREIGN sky130_hilas_WTA4Stage01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.240 BY 9.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 15.790 1.590 16.120 1.680 ;
        RECT 9.440 1.420 16.120 1.590 ;
        RECT 15.790 1.390 16.120 1.420 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.850 1.700 16.080 6.050 ;
        RECT 15.810 1.690 16.090 1.700 ;
        RECT 15.810 1.370 16.110 1.690 ;
        RECT 15.850 0.000 16.080 1.370 ;
      LAYER via ;
        RECT 15.820 1.400 16.090 1.670 ;
    END
  END VGND
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 12.740 5.000 12.780 5.090 ;
        RECT 12.630 4.910 13.840 5.000 ;
        RECT 12.630 4.850 13.970 4.910 ;
        RECT 12.630 4.800 16.240 4.850 ;
        RECT 13.660 4.690 16.240 4.800 ;
        RECT 13.660 4.580 13.970 4.690 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 12.730 4.030 13.940 4.140 ;
        RECT 12.730 3.940 13.970 4.030 ;
        RECT 13.660 3.920 13.970 3.940 ;
        RECT 13.660 3.760 16.240 3.920 ;
        RECT 13.660 3.700 13.970 3.760 ;
    END
  END OUTPUT2
  PIN OUTPUT3
    USE ANALOG ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 13.660 2.110 13.970 2.140 ;
        RECT 12.720 2.080 13.970 2.110 ;
        RECT 12.720 1.950 16.240 2.080 ;
        RECT 13.660 1.920 16.240 1.950 ;
        RECT 13.660 1.810 13.970 1.920 ;
    END
  END OUTPUT3
  PIN OUTPUT4
    USE ANALOG ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 13.660 1.150 13.970 1.260 ;
        RECT 13.660 1.140 16.240 1.150 ;
        RECT 12.730 0.990 16.240 1.140 ;
        RECT 12.730 0.960 13.970 0.990 ;
        RECT 13.660 0.930 13.970 0.960 ;
    END
  END OUTPUT4
  PIN INPUT1
    USE ANALOG ;
    ANTENNAGATEAREA 0.236000 ;
    ANTENNADIFFAREA 4.378700 ;
    PORT
      LAYER nwell ;
        RECT 0.020 9.860 2.570 9.870 ;
        RECT 0.010 6.050 2.570 9.860 ;
        RECT 4.100 6.050 6.330 9.870 ;
        RECT 0.010 6.040 6.330 6.050 ;
        RECT 0.010 5.890 2.680 6.040 ;
        RECT 0.010 5.880 2.860 5.890 ;
        RECT 0.010 3.840 2.680 5.880 ;
        RECT 0.020 3.830 2.680 3.840 ;
        RECT 2.160 2.970 2.680 3.830 ;
        RECT 4.100 3.820 6.330 6.040 ;
        RECT 2.270 0.010 2.680 2.970 ;
      LAYER met2 ;
        RECT 2.170 5.930 2.480 5.950 ;
        RECT 0.010 5.770 10.080 5.930 ;
        RECT 0.010 5.760 10.070 5.770 ;
        RECT 0.010 5.750 2.570 5.760 ;
        RECT 2.170 5.620 2.480 5.750 ;
        RECT 5.430 5.740 5.750 5.760 ;
        RECT 5.430 5.550 13.350 5.740 ;
        RECT 13.510 5.550 13.820 5.590 ;
        RECT 5.430 5.530 13.820 5.550 ;
        RECT 5.430 5.500 5.750 5.530 ;
        RECT 13.140 5.340 13.820 5.530 ;
        RECT 13.510 5.260 13.820 5.340 ;
        RECT 2.160 5.070 2.310 5.120 ;
        RECT 2.160 4.950 2.480 5.070 ;
        RECT 2.160 4.940 10.080 4.950 ;
        RECT 0.010 4.780 10.080 4.940 ;
        RECT 0.010 4.760 2.570 4.780 ;
        RECT 2.160 4.740 2.480 4.760 ;
        RECT 2.160 4.610 2.310 4.740 ;
        RECT 5.410 4.610 5.730 4.710 ;
        RECT 7.750 4.690 9.290 4.780 ;
        RECT 2.160 4.510 5.730 4.610 ;
        RECT 0.010 4.450 5.730 4.510 ;
        RECT 0.010 4.340 2.580 4.450 ;
        RECT 0.010 4.330 2.480 4.340 ;
        RECT 2.170 4.210 2.480 4.330 ;
        RECT 2.140 4.190 2.480 4.210 ;
        RECT 2.140 3.950 2.460 4.190 ;
        RECT 2.210 3.940 2.380 3.950 ;
        RECT 5.370 3.470 5.600 3.480 ;
        RECT 5.370 3.440 12.940 3.470 ;
        RECT 5.370 3.270 13.000 3.440 ;
        RECT 13.510 3.270 13.820 3.350 ;
        RECT 2.120 3.170 2.440 3.200 ;
        RECT 5.370 3.170 5.610 3.270 ;
        RECT 2.120 2.990 5.610 3.170 ;
        RECT 12.810 3.070 13.820 3.270 ;
        RECT 13.410 3.060 13.820 3.070 ;
        RECT 13.510 3.020 13.820 3.060 ;
        RECT 2.120 2.970 5.530 2.990 ;
        RECT 2.120 2.940 2.440 2.970 ;
    END
  END INPUT1
  PIN INPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.099200 ;
    PORT
      LAYER met1 ;
        RECT 2.160 4.200 2.480 4.520 ;
        RECT 2.170 4.120 2.430 4.200 ;
        RECT 2.160 3.920 2.430 4.120 ;
        RECT 2.160 3.230 2.370 3.920 ;
        RECT 2.150 2.910 2.410 3.230 ;
      LAYER via ;
        RECT 2.190 4.230 2.450 4.490 ;
        RECT 2.170 3.950 2.430 4.210 ;
        RECT 2.150 2.940 2.410 3.200 ;
    END
  END INPUT2
  PIN INPUT3
    USE ANALOG ;
    ANTENNAGATEAREA 0.118000 ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 5.410 2.790 5.730 2.830 ;
        RECT 5.410 2.770 12.960 2.790 ;
        RECT 13.510 2.780 13.820 2.820 ;
        RECT 13.410 2.770 13.820 2.780 ;
        RECT 5.410 2.570 13.820 2.770 ;
        RECT 5.510 2.560 5.830 2.570 ;
        RECT 13.510 2.490 13.820 2.570 ;
        RECT 2.100 1.610 2.300 2.110 ;
        RECT 5.250 1.610 5.570 1.650 ;
        RECT 2.100 1.410 5.650 1.610 ;
        RECT 5.250 1.390 5.570 1.410 ;
    END
  END INPUT3
  PIN INPUT4
    USE ANALOG ;
    ANTENNAGATEAREA 0.118000 ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 2.070 0.870 2.380 1.200 ;
        RECT 13.510 0.520 13.820 0.580 ;
        RECT 12.960 0.510 13.820 0.520 ;
        RECT 2.120 0.230 2.430 0.350 ;
        RECT 5.380 0.290 13.820 0.510 ;
        RECT 5.380 0.280 12.970 0.290 ;
        RECT 5.380 0.270 6.150 0.280 ;
        RECT 5.380 0.230 5.620 0.270 ;
        RECT 13.510 0.250 13.820 0.290 ;
        RECT 2.120 0.030 5.620 0.230 ;
        RECT 2.120 0.020 4.810 0.030 ;
    END
  END INPUT4
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 2.120 5.370 2.670 5.550 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 2.100 3.510 2.670 3.690 ;
    END
  END DRAIN2
  PIN DRAIN3
    PORT
      LAYER met2 ;
        RECT 2.120 2.360 2.670 2.540 ;
        RECT 2.120 2.350 2.280 2.360 ;
    END
  END DRAIN3
  PIN DRAIN4
    PORT
      LAYER met2 ;
        RECT 2.140 0.690 2.300 0.700 ;
        RECT 2.140 0.510 2.670 0.690 ;
    END
  END DRAIN4
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT 7.960 5.950 8.340 6.050 ;
    END
  END GATE1
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 11.990 5.910 12.390 6.050 ;
    END
  END VTUN
  PIN WTAMIDDLENODE
    ANTENNAGATEAREA 0.472000 ;
    ANTENNADIFFAREA 0.708000 ;
    PORT
      LAYER met1 ;
        RECT 14.590 0.000 14.820 6.050 ;
    END
  END WTAMIDDLENODE
  PIN COLSEL1
    ANTENNADIFFAREA 1.053100 ;
    PORT
      LAYER met2 ;
        RECT 3.200 5.340 3.520 5.400 ;
        RECT 7.220 5.340 7.550 5.370 ;
        RECT 3.200 5.170 7.550 5.340 ;
        RECT 3.200 5.120 3.520 5.170 ;
        RECT 7.220 5.110 7.550 5.170 ;
    END
  END COLSEL1
  PIN VPWR
    PORT
      LAYER met1 ;
        RECT 3.840 5.980 4.000 6.050 ;
    END
  END VPWR
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 3.030 5.980 3.190 6.050 ;
    END
  END VINJ
  OBS
      LAYER nwell ;
        RECT 8.350 9.240 10.080 9.870 ;
        RECT 8.350 6.170 10.090 9.240 ;
        RECT 7.960 5.950 8.340 6.050 ;
        RECT 8.350 3.820 10.080 6.170 ;
        RECT 11.990 5.910 12.390 6.050 ;
      LAYER li1 ;
        RECT 0.410 9.190 0.610 9.540 ;
        RECT 2.150 9.460 2.470 9.470 ;
        RECT 1.890 9.290 2.470 9.460 ;
        RECT 2.140 9.240 2.470 9.290 ;
        RECT 2.150 9.210 2.470 9.240 ;
        RECT 0.400 9.160 0.610 9.190 ;
        RECT 0.400 8.570 0.620 9.160 ;
        RECT 1.140 8.600 1.340 9.170 ;
        RECT 2.150 8.880 2.470 8.920 ;
        RECT 2.140 8.840 2.470 8.880 ;
        RECT 1.890 8.670 2.470 8.840 ;
        RECT 2.150 8.660 2.470 8.670 ;
        RECT 0.400 7.540 0.620 8.130 ;
        RECT 0.400 7.510 0.610 7.540 ;
        RECT 1.140 7.530 1.340 8.100 ;
        RECT 3.280 8.090 3.450 8.600 ;
        RECT 7.300 8.120 7.470 8.630 ;
        RECT 2.150 8.030 2.470 8.040 ;
        RECT 1.890 7.860 2.470 8.030 ;
        RECT 2.140 7.820 2.470 7.860 ;
        RECT 2.150 7.780 2.470 7.820 ;
        RECT 0.410 7.160 0.610 7.510 ;
        RECT 2.150 7.460 2.470 7.490 ;
        RECT 2.140 7.410 2.470 7.460 ;
        RECT 1.890 7.240 2.470 7.410 ;
        RECT 2.150 7.230 2.470 7.240 ;
        RECT 0.780 6.760 1.220 6.930 ;
        RECT 0.410 6.180 0.610 6.530 ;
        RECT 2.150 6.450 2.470 6.460 ;
        RECT 1.890 6.280 2.470 6.450 ;
        RECT 2.140 6.230 2.470 6.280 ;
        RECT 3.270 6.230 3.440 7.420 ;
        RECT 5.080 6.550 5.630 6.980 ;
        RECT 2.150 6.200 2.470 6.230 ;
        RECT 0.400 6.150 0.610 6.180 ;
        RECT 7.290 6.170 7.460 7.360 ;
        RECT 9.110 6.620 9.660 7.050 ;
        RECT 0.400 5.560 0.620 6.150 ;
        RECT 1.140 5.590 1.340 6.160 ;
        RECT 2.150 5.870 2.470 5.910 ;
        RECT 2.140 5.830 2.470 5.870 ;
        RECT 1.890 5.660 2.470 5.830 ;
        RECT 2.150 5.650 2.470 5.660 ;
        RECT 13.520 5.530 13.840 5.560 ;
        RECT 13.520 5.360 15.310 5.530 ;
        RECT 13.520 5.340 13.850 5.360 ;
        RECT 13.520 5.300 13.840 5.340 ;
        RECT 15.140 5.130 15.310 5.360 ;
        RECT 0.400 4.540 0.620 5.130 ;
        RECT 0.400 4.510 0.610 4.540 ;
        RECT 1.140 4.530 1.340 5.100 ;
        RECT 2.150 5.030 2.470 5.040 ;
        RECT 1.890 4.860 2.470 5.030 ;
        RECT 13.990 4.880 14.330 5.130 ;
        RECT 14.500 4.960 14.830 5.130 ;
        RECT 15.050 4.960 15.390 5.130 ;
        RECT 2.140 4.820 2.470 4.860 ;
        RECT 2.150 4.780 2.470 4.820 ;
        RECT 13.670 4.620 14.330 4.880 ;
        RECT 14.580 4.790 14.750 4.960 ;
        RECT 15.140 4.790 15.310 4.960 ;
        RECT 14.500 4.620 14.830 4.790 ;
        RECT 15.050 4.620 15.390 4.790 ;
        RECT 0.410 4.160 0.610 4.510 ;
        RECT 2.150 4.460 2.470 4.490 ;
        RECT 2.140 4.410 2.470 4.460 ;
        RECT 1.890 4.240 2.470 4.410 ;
        RECT 2.150 4.230 2.470 4.240 ;
        RECT 14.580 4.390 14.830 4.620 ;
        RECT 15.710 4.540 16.220 5.210 ;
        RECT 14.580 4.220 15.250 4.390 ;
        RECT 14.580 3.990 14.830 4.220 ;
        RECT 13.670 3.730 14.330 3.990 ;
        RECT 14.500 3.820 14.830 3.990 ;
        RECT 15.050 3.820 15.390 3.990 ;
        RECT 13.990 3.480 14.330 3.730 ;
        RECT 14.580 3.650 14.750 3.820 ;
        RECT 15.140 3.650 15.310 3.820 ;
        RECT 14.500 3.480 14.830 3.650 ;
        RECT 15.050 3.480 15.390 3.650 ;
        RECT 13.520 3.270 13.840 3.310 ;
        RECT 13.520 3.250 13.850 3.270 ;
        RECT 15.140 3.250 15.310 3.480 ;
        RECT 15.710 3.400 16.220 4.070 ;
        RECT 13.520 3.080 15.310 3.250 ;
        RECT 13.520 3.050 13.840 3.080 ;
        RECT 13.520 2.760 13.840 2.790 ;
        RECT 13.520 2.590 15.310 2.760 ;
        RECT 13.520 2.570 13.850 2.590 ;
        RECT 13.520 2.530 13.840 2.570 ;
        RECT 15.140 2.360 15.310 2.590 ;
        RECT 13.990 2.110 14.330 2.360 ;
        RECT 14.500 2.190 14.830 2.360 ;
        RECT 15.050 2.190 15.390 2.360 ;
        RECT 13.670 1.850 14.330 2.110 ;
        RECT 14.580 2.020 14.750 2.190 ;
        RECT 15.140 2.020 15.310 2.190 ;
        RECT 14.500 1.850 14.830 2.020 ;
        RECT 15.050 1.850 15.390 2.020 ;
        RECT 14.580 1.620 14.830 1.850 ;
        RECT 15.710 1.770 16.220 2.440 ;
        RECT 14.580 1.450 15.250 1.620 ;
        RECT 14.580 1.220 14.830 1.450 ;
        RECT 2.080 1.120 2.400 1.160 ;
        RECT 2.080 0.930 2.410 1.120 ;
        RECT 13.670 0.960 14.330 1.220 ;
        RECT 14.500 1.050 14.830 1.220 ;
        RECT 15.050 1.050 15.390 1.220 ;
        RECT 2.080 0.900 2.400 0.930 ;
        RECT 2.130 0.310 2.310 0.900 ;
        RECT 13.990 0.710 14.330 0.960 ;
        RECT 14.580 0.880 14.750 1.050 ;
        RECT 15.140 0.880 15.310 1.050 ;
        RECT 14.500 0.710 14.830 0.880 ;
        RECT 15.050 0.710 15.390 0.880 ;
        RECT 13.520 0.500 13.840 0.540 ;
        RECT 13.520 0.480 13.850 0.500 ;
        RECT 15.140 0.480 15.310 0.710 ;
        RECT 15.710 0.630 16.220 1.300 ;
        RECT 13.520 0.310 15.310 0.480 ;
        RECT 2.130 0.270 2.450 0.310 ;
        RECT 13.520 0.280 13.840 0.310 ;
        RECT 2.130 0.080 2.460 0.270 ;
        RECT 2.130 0.050 2.450 0.080 ;
      LAYER mcon ;
        RECT 2.240 9.250 2.410 9.420 ;
        RECT 0.430 8.990 0.600 9.160 ;
        RECT 1.160 8.960 1.330 9.130 ;
        RECT 2.240 8.700 2.410 8.870 ;
        RECT 3.280 8.430 3.450 8.600 ;
        RECT 0.430 7.540 0.600 7.710 ;
        RECT 7.300 8.460 7.470 8.630 ;
        RECT 2.240 7.830 2.410 8.000 ;
        RECT 1.160 7.570 1.330 7.740 ;
        RECT 2.240 7.280 2.410 7.450 ;
        RECT 3.270 7.250 3.440 7.420 ;
        RECT 3.270 6.910 3.440 7.080 ;
        RECT 7.290 7.190 7.460 7.360 ;
        RECT 3.270 6.570 3.440 6.740 ;
        RECT 2.240 6.240 2.410 6.410 ;
        RECT 5.360 6.630 5.630 6.900 ;
        RECT 7.290 6.850 7.460 7.020 ;
        RECT 7.290 6.510 7.460 6.680 ;
        RECT 9.390 6.700 9.660 6.970 ;
        RECT 0.430 5.980 0.600 6.150 ;
        RECT 1.160 5.950 1.330 6.120 ;
        RECT 2.240 5.690 2.410 5.860 ;
        RECT 13.580 5.350 13.750 5.520 ;
        RECT 0.430 4.540 0.600 4.710 ;
        RECT 2.240 4.830 2.410 5.000 ;
        RECT 1.160 4.570 1.330 4.740 ;
        RECT 13.730 4.670 13.900 4.840 ;
        RECT 15.880 4.790 16.050 4.960 ;
        RECT 2.240 4.280 2.410 4.450 ;
        RECT 14.620 4.220 14.790 4.390 ;
        RECT 13.730 3.770 13.900 3.940 ;
        RECT 15.880 3.650 16.050 3.820 ;
        RECT 13.580 3.090 13.750 3.260 ;
        RECT 13.580 2.580 13.750 2.750 ;
        RECT 13.730 1.900 13.900 2.070 ;
        RECT 15.880 2.020 16.050 2.190 ;
        RECT 14.620 1.450 14.790 1.620 ;
        RECT 2.140 0.940 2.310 1.110 ;
        RECT 13.730 1.000 13.900 1.170 ;
        RECT 15.880 0.880 16.050 1.050 ;
        RECT 13.580 0.320 13.750 0.490 ;
        RECT 2.190 0.090 2.360 0.260 ;
      LAYER met1 ;
        RECT 0.370 9.220 0.530 9.870 ;
        RECT 0.370 8.670 0.640 9.220 ;
        RECT 0.360 8.620 0.640 8.670 ;
        RECT 0.780 8.880 0.970 9.870 ;
        RECT 1.180 9.190 1.340 9.870 ;
        RECT 1.140 9.170 1.340 9.190 ;
        RECT 2.160 9.180 2.480 9.500 ;
        RECT 1.130 8.930 1.360 9.170 ;
        RECT 0.780 8.760 0.950 8.880 ;
        RECT 0.360 8.530 0.530 8.620 ;
        RECT 0.370 8.170 0.530 8.530 ;
        RECT 0.360 8.080 0.530 8.170 ;
        RECT 0.360 8.030 0.640 8.080 ;
        RECT 0.370 7.480 0.640 8.030 ;
        RECT 0.780 7.940 0.940 8.760 ;
        RECT 1.140 8.710 1.340 8.930 ;
        RECT 1.180 7.990 1.340 8.710 ;
        RECT 2.160 8.630 2.480 8.950 ;
        RECT 0.780 7.820 0.950 7.940 ;
        RECT 0.370 6.210 0.530 7.480 ;
        RECT 0.780 6.960 0.970 7.820 ;
        RECT 1.140 7.770 1.340 7.990 ;
        RECT 1.130 7.530 1.360 7.770 ;
        RECT 2.160 7.750 2.480 8.070 ;
        RECT 1.140 7.510 1.340 7.530 ;
        RECT 0.750 6.730 0.990 6.960 ;
        RECT 0.370 5.660 0.640 6.210 ;
        RECT 0.360 5.610 0.640 5.660 ;
        RECT 0.780 5.870 0.970 6.730 ;
        RECT 1.180 6.180 1.340 7.510 ;
        RECT 2.160 7.200 2.480 7.520 ;
        RECT 1.140 6.160 1.340 6.180 ;
        RECT 2.160 6.170 2.480 6.490 ;
        RECT 1.130 5.920 1.360 6.160 ;
        RECT 3.240 6.050 3.490 9.870 ;
        RECT 5.300 7.950 5.680 9.870 ;
        RECT 5.300 6.090 5.690 7.950 ;
        RECT 3.240 5.980 3.630 6.050 ;
        RECT 0.780 5.750 0.950 5.870 ;
        RECT 0.360 5.520 0.530 5.610 ;
        RECT 0.370 5.170 0.530 5.520 ;
        RECT 0.360 5.080 0.530 5.170 ;
        RECT 0.360 5.030 0.640 5.080 ;
        RECT 0.370 4.480 0.640 5.030 ;
        RECT 0.780 4.940 0.940 5.750 ;
        RECT 1.140 5.700 1.340 5.920 ;
        RECT 1.180 4.990 1.340 5.700 ;
        RECT 2.160 5.620 2.480 5.940 ;
        RECT 3.240 5.430 3.490 5.980 ;
        RECT 5.300 5.790 5.680 6.090 ;
        RECT 5.300 5.470 5.720 5.790 ;
        RECT 3.220 5.400 3.500 5.430 ;
        RECT 3.210 5.120 3.510 5.400 ;
        RECT 3.220 5.100 3.500 5.120 ;
        RECT 0.780 4.820 0.950 4.940 ;
        RECT 0.370 3.830 0.530 4.480 ;
        RECT 0.780 3.830 0.970 4.820 ;
        RECT 1.140 4.770 1.340 4.990 ;
        RECT 1.130 4.530 1.360 4.770 ;
        RECT 2.160 4.750 2.480 5.070 ;
        RECT 1.140 4.510 1.340 4.530 ;
        RECT 1.180 3.830 1.340 4.510 ;
        RECT 3.240 3.820 3.490 5.100 ;
        RECT 5.300 4.740 5.680 5.470 ;
        RECT 7.250 5.400 7.520 9.870 ;
        RECT 7.230 5.090 7.540 5.400 ;
        RECT 5.300 4.420 5.700 4.740 ;
        RECT 5.300 3.820 5.680 4.420 ;
        RECT 7.250 3.820 7.520 5.090 ;
        RECT 9.330 3.820 9.730 9.870 ;
        RECT 13.510 5.270 13.830 5.590 ;
        RECT 13.660 4.590 13.980 4.910 ;
        RECT 13.660 3.700 13.980 4.020 ;
        RECT 13.510 3.020 13.830 3.340 ;
        RECT 5.440 2.540 5.700 2.860 ;
        RECT 5.440 1.680 5.600 2.540 ;
        RECT 13.510 2.500 13.830 2.820 ;
        RECT 13.660 1.820 13.980 2.140 ;
        RECT 5.280 1.360 5.600 1.680 ;
        RECT 2.070 0.870 2.390 1.190 ;
        RECT 13.660 0.930 13.980 1.250 ;
        RECT 2.120 0.020 2.440 0.340 ;
        RECT 13.510 0.250 13.830 0.570 ;
        RECT 7.960 0.000 8.340 0.100 ;
      LAYER via ;
        RECT 2.190 9.210 2.450 9.470 ;
        RECT 2.190 8.660 2.450 8.920 ;
        RECT 2.190 7.780 2.450 8.040 ;
        RECT 2.190 7.230 2.450 7.490 ;
        RECT 2.190 6.200 2.450 6.460 ;
        RECT 2.190 5.650 2.450 5.910 ;
        RECT 5.460 5.500 5.720 5.760 ;
        RECT 3.230 5.130 3.490 5.390 ;
        RECT 2.190 4.780 2.450 5.040 ;
        RECT 7.250 5.110 7.520 5.370 ;
        RECT 5.440 4.450 5.700 4.710 ;
        RECT 13.540 5.300 13.800 5.560 ;
        RECT 13.690 4.620 13.950 4.880 ;
        RECT 13.690 3.730 13.950 3.990 ;
        RECT 13.540 3.050 13.800 3.310 ;
        RECT 5.440 2.570 5.700 2.830 ;
        RECT 13.540 2.530 13.800 2.790 ;
        RECT 13.690 1.850 13.950 2.110 ;
        RECT 5.280 1.390 5.540 1.650 ;
        RECT 2.100 0.900 2.360 1.160 ;
        RECT 13.690 0.960 13.950 1.220 ;
        RECT 2.150 0.050 2.410 0.310 ;
        RECT 13.540 0.280 13.800 0.540 ;
      LAYER met2 ;
        RECT 2.170 9.370 2.480 9.510 ;
        RECT 0.010 9.190 2.580 9.370 ;
        RECT 2.170 9.180 2.480 9.190 ;
        RECT 2.170 8.940 2.480 8.960 ;
        RECT 0.010 8.760 10.090 8.940 ;
        RECT 2.170 8.630 2.480 8.760 ;
        RECT 9.940 8.750 10.090 8.760 ;
        RECT 2.170 7.940 2.480 8.070 ;
        RECT 9.970 7.940 10.110 7.960 ;
        RECT 0.000 7.760 10.110 7.940 ;
        RECT 2.170 7.740 2.480 7.760 ;
        RECT 2.170 7.510 2.480 7.520 ;
        RECT 0.010 7.470 2.480 7.510 ;
        RECT 0.010 7.330 2.570 7.470 ;
        RECT 2.170 7.190 2.480 7.330 ;
        RECT 2.170 6.360 2.480 6.500 ;
        RECT 0.000 6.350 2.480 6.360 ;
        RECT 0.000 6.180 2.600 6.350 ;
        RECT 2.170 6.170 2.480 6.180 ;
  END
END sky130_hilas_WTA4Stage01

MACRO sky130_hilas_Trans4small
  CLASS CORE ;
  FOREIGN sky130_hilas_Trans4small ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.800 BY 5.880 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN NFET_SOURCE1
    USE ANALOG ;
    ANTENNADIFFAREA 0.108500 ;
    PORT
      LAYER met2 ;
        RECT 0.600 5.650 0.910 5.740 ;
        RECT 0.000 5.480 0.910 5.650 ;
        RECT 0.600 5.410 0.910 5.480 ;
    END
  END NFET_SOURCE1
  PIN NFET_GATE1
    USE ANALOG ;
    ANTENNAGATEAREA 0.094500 ;
    PORT
      LAYER met2 ;
        RECT 0.130 5.240 0.450 5.320 ;
        RECT 0.000 5.070 0.450 5.240 ;
        RECT 0.130 5.000 0.450 5.070 ;
    END
  END NFET_GATE1
  PIN NFET_SOURCE2
    USE ANALOG ;
    ANTENNADIFFAREA 0.108500 ;
    PORT
      LAYER met2 ;
        RECT 0.600 4.730 0.910 4.820 ;
        RECT 0.000 4.560 0.910 4.730 ;
        RECT 0.600 4.490 0.910 4.560 ;
    END
  END NFET_SOURCE2
  PIN NFET_GATE2
    USE ANALOG ;
    ANTENNAGATEAREA 0.094500 ;
    PORT
      LAYER met2 ;
        RECT 0.130 4.320 0.450 4.400 ;
        RECT 0.000 4.150 0.450 4.320 ;
        RECT 0.130 4.080 0.450 4.150 ;
    END
  END NFET_GATE2
  PIN NFET_SOURCE3
    USE ANALOG ;
    ANTENNADIFFAREA 0.108500 ;
    PORT
      LAYER met2 ;
        RECT 0.600 3.810 0.910 3.900 ;
        RECT 0.000 3.640 0.910 3.810 ;
        RECT 0.600 3.570 0.910 3.640 ;
    END
  END NFET_SOURCE3
  PIN NFET_GATE3
    USE ANALOG ;
    ANTENNAGATEAREA 0.094500 ;
    PORT
      LAYER met2 ;
        RECT 0.130 3.400 0.450 3.480 ;
        RECT 0.000 3.230 0.450 3.400 ;
        RECT 0.130 3.160 0.450 3.230 ;
    END
  END NFET_GATE3
  PIN PFET_SOURCE1
    USE ANALOG ;
    ANTENNADIFFAREA 0.109200 ;
    PORT
      LAYER met2 ;
        RECT 0.410 2.810 0.720 2.920 ;
        RECT 0.000 2.620 0.720 2.810 ;
        RECT 0.410 2.590 0.720 2.620 ;
    END
  END PFET_SOURCE1
  PIN PFET_GATE1
    USE ANALOG ;
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER met2 ;
        RECT 0.410 2.390 0.730 2.450 ;
        RECT 0.000 2.200 0.730 2.390 ;
        RECT 0.410 2.130 0.730 2.200 ;
    END
  END PFET_GATE1
  PIN PFET_SOURCE2
    USE ANALOG ;
    ANTENNADIFFAREA 0.109200 ;
    PORT
      LAYER met2 ;
        RECT 0.410 1.850 0.720 1.960 ;
        RECT 0.000 1.660 0.720 1.850 ;
        RECT 0.410 1.630 0.720 1.660 ;
    END
  END PFET_SOURCE2
  PIN PFET_GATE2
    USE ANALOG ;
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER met2 ;
        RECT 0.410 1.430 0.730 1.490 ;
        RECT 0.000 1.240 0.730 1.430 ;
        RECT 0.410 1.170 0.730 1.240 ;
    END
  END PFET_GATE2
  PIN PFET_SOURCE3
    USE ANALOG ;
    ANTENNADIFFAREA 0.109200 ;
    PORT
      LAYER met2 ;
        RECT 0.410 0.890 0.720 1.000 ;
        RECT 0.000 0.700 0.720 0.890 ;
        RECT 0.410 0.670 0.720 0.700 ;
    END
  END PFET_SOURCE3
  PIN PFET_GATE3
    USE ANALOG ;
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER met2 ;
        RECT 0.410 0.470 0.730 0.530 ;
        RECT 0.000 0.280 0.730 0.470 ;
        RECT 0.410 0.210 0.730 0.280 ;
    END
  END PFET_GATE3
  PIN WELL
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.070 0.000 2.640 3.090 ;
      LAYER met1 ;
        RECT 2.180 0.400 2.400 5.880 ;
        RECT 2.120 0.170 2.410 0.400 ;
        RECT 2.180 0.000 2.400 0.170 ;
    END
  END WELL
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2.580 5.250 2.800 5.880 ;
        RECT 2.570 4.960 2.800 5.250 ;
        RECT 2.580 0.000 2.800 4.960 ;
    END
  END VGND
  PIN PFET_DRAIN3
    USE ANALOG ;
    ANTENNADIFFAREA 0.105300 ;
    PORT
      LAYER met2 ;
        RECT 1.710 0.830 2.020 0.900 ;
        RECT 1.710 0.630 2.800 0.830 ;
        RECT 1.710 0.570 2.020 0.630 ;
    END
  END PFET_DRAIN3
  PIN PFET_DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.105300 ;
    PORT
      LAYER met2 ;
        RECT 1.710 1.790 2.020 1.860 ;
        RECT 1.710 1.590 2.800 1.790 ;
        RECT 1.710 1.530 2.020 1.590 ;
    END
  END PFET_DRAIN2
  PIN PFET_DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.105300 ;
    PORT
      LAYER met2 ;
        RECT 1.710 2.750 2.020 2.820 ;
        RECT 1.710 2.550 2.800 2.750 ;
        RECT 1.710 2.490 2.020 2.550 ;
    END
  END PFET_DRAIN1
  PIN NFET_DRAIN3
    USE ANALOG ;
    ANTENNADIFFAREA 0.108500 ;
    PORT
      LAYER met2 ;
        RECT 1.690 3.820 2.000 3.910 ;
        RECT 1.690 3.650 2.800 3.820 ;
        RECT 1.690 3.580 2.000 3.650 ;
    END
  END NFET_DRAIN3
  PIN NFET_DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.108500 ;
    PORT
      LAYER met2 ;
        RECT 1.690 4.740 2.000 4.830 ;
        RECT 1.690 4.570 2.800 4.740 ;
        RECT 1.690 4.500 2.000 4.570 ;
    END
  END NFET_DRAIN2
  PIN NFET_DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.108500 ;
    PORT
      LAYER met2 ;
        RECT 1.690 5.660 2.000 5.750 ;
        RECT 1.690 5.490 2.800 5.660 ;
        RECT 1.690 5.420 2.000 5.490 ;
    END
  END NFET_DRAIN1
  OBS
      LAYER li1 ;
        RECT 0.920 5.700 1.120 5.740 ;
        RECT 0.610 5.440 1.120 5.700 ;
        RECT 0.920 5.410 1.120 5.440 ;
        RECT 1.510 5.710 1.710 5.740 ;
        RECT 1.510 5.670 2.020 5.710 ;
        RECT 1.510 5.480 2.030 5.670 ;
        RECT 1.510 5.450 2.020 5.480 ;
        RECT 1.510 5.410 1.710 5.450 ;
        RECT 2.200 5.260 2.370 5.310 ;
        RECT 0.170 5.240 0.600 5.260 ;
        RECT 0.170 5.070 0.620 5.240 ;
        RECT 2.190 5.230 2.370 5.260 ;
        RECT 2.190 5.220 2.620 5.230 ;
        RECT 0.170 5.050 0.600 5.070 ;
        RECT 2.190 4.990 2.780 5.220 ;
        RECT 2.190 4.980 2.620 4.990 ;
        RECT 2.190 4.920 2.360 4.980 ;
        RECT 0.920 4.780 1.120 4.820 ;
        RECT 0.610 4.520 1.120 4.780 ;
        RECT 0.920 4.490 1.120 4.520 ;
        RECT 1.510 4.790 1.710 4.820 ;
        RECT 1.510 4.750 2.020 4.790 ;
        RECT 1.510 4.560 2.030 4.750 ;
        RECT 1.510 4.530 2.020 4.560 ;
        RECT 1.510 4.490 1.710 4.530 ;
        RECT 0.170 4.320 0.600 4.340 ;
        RECT 0.170 4.150 0.620 4.320 ;
        RECT 0.170 4.130 0.600 4.150 ;
        RECT 0.920 3.860 1.120 3.900 ;
        RECT 0.610 3.600 1.120 3.860 ;
        RECT 0.920 3.570 1.120 3.600 ;
        RECT 1.510 3.870 1.710 3.900 ;
        RECT 1.510 3.830 2.020 3.870 ;
        RECT 1.510 3.640 2.030 3.830 ;
        RECT 1.510 3.610 2.020 3.640 ;
        RECT 1.510 3.570 1.710 3.610 ;
        RECT 0.170 3.400 0.600 3.420 ;
        RECT 0.170 3.230 0.620 3.400 ;
        RECT 0.170 3.210 0.600 3.230 ;
        RECT 0.420 2.840 0.740 2.880 ;
        RECT 0.420 2.820 0.750 2.840 ;
        RECT 0.420 2.620 1.040 2.820 ;
        RECT 0.870 2.490 1.040 2.620 ;
        RECT 1.550 2.780 1.720 2.820 ;
        RECT 1.550 2.740 2.040 2.780 ;
        RECT 1.550 2.550 2.050 2.740 ;
        RECT 1.550 2.520 2.040 2.550 ;
        RECT 1.550 2.490 1.720 2.520 ;
        RECT 0.260 2.380 0.690 2.400 ;
        RECT 0.240 2.210 0.690 2.380 ;
        RECT 0.260 2.190 0.690 2.210 ;
        RECT 0.420 1.880 0.740 1.920 ;
        RECT 0.420 1.860 0.750 1.880 ;
        RECT 0.420 1.660 1.040 1.860 ;
        RECT 0.870 1.530 1.040 1.660 ;
        RECT 1.550 1.820 1.720 1.860 ;
        RECT 1.550 1.780 2.040 1.820 ;
        RECT 1.550 1.590 2.050 1.780 ;
        RECT 1.550 1.560 2.040 1.590 ;
        RECT 1.550 1.530 1.720 1.560 ;
        RECT 0.260 1.420 0.690 1.440 ;
        RECT 0.240 1.250 0.690 1.420 ;
        RECT 0.260 1.230 0.690 1.250 ;
        RECT 0.420 0.920 0.740 0.960 ;
        RECT 0.420 0.900 0.750 0.920 ;
        RECT 0.420 0.700 1.040 0.900 ;
        RECT 0.870 0.570 1.040 0.700 ;
        RECT 1.550 0.860 1.720 0.900 ;
        RECT 1.550 0.820 2.040 0.860 ;
        RECT 1.550 0.630 2.050 0.820 ;
        RECT 1.550 0.600 2.040 0.630 ;
        RECT 1.550 0.570 1.720 0.600 ;
        RECT 0.260 0.460 0.690 0.480 ;
        RECT 0.240 0.290 0.690 0.460 ;
        RECT 0.260 0.270 0.690 0.290 ;
        RECT 2.050 0.230 2.470 0.400 ;
        RECT 2.150 0.190 2.380 0.230 ;
      LAYER mcon ;
        RECT 0.670 5.480 0.840 5.650 ;
        RECT 1.760 5.490 1.930 5.660 ;
        RECT 0.450 5.070 0.620 5.240 ;
        RECT 2.600 5.020 2.770 5.190 ;
        RECT 0.670 4.560 0.840 4.730 ;
        RECT 1.760 4.570 1.930 4.740 ;
        RECT 0.450 4.150 0.620 4.320 ;
        RECT 0.670 3.640 0.840 3.810 ;
        RECT 1.760 3.650 1.930 3.820 ;
        RECT 0.450 3.230 0.620 3.400 ;
        RECT 0.480 2.660 0.650 2.830 ;
        RECT 1.780 2.560 1.950 2.730 ;
        RECT 0.480 1.700 0.650 1.870 ;
        RECT 1.780 1.600 1.950 1.770 ;
        RECT 0.480 0.740 0.650 0.910 ;
        RECT 1.780 0.640 1.950 0.810 ;
        RECT 2.180 0.200 2.350 0.370 ;
      LAYER met1 ;
        RECT 0.600 5.410 0.920 5.730 ;
        RECT 1.690 5.420 2.010 5.740 ;
        RECT 0.130 5.270 0.450 5.320 ;
        RECT 0.130 5.040 0.680 5.270 ;
        RECT 0.130 5.000 0.450 5.040 ;
        RECT 0.600 4.490 0.920 4.810 ;
        RECT 1.690 4.500 2.010 4.820 ;
        RECT 0.130 4.350 0.450 4.400 ;
        RECT 0.130 4.120 0.680 4.350 ;
        RECT 0.130 4.080 0.450 4.120 ;
        RECT 0.600 3.570 0.920 3.890 ;
        RECT 1.690 3.580 2.010 3.900 ;
        RECT 0.130 3.430 0.450 3.480 ;
        RECT 0.130 3.200 0.680 3.430 ;
        RECT 0.130 3.160 0.450 3.200 ;
        RECT 0.410 2.590 0.730 2.910 ;
        RECT 1.710 2.490 2.030 2.810 ;
        RECT 0.410 2.410 0.730 2.450 ;
        RECT 0.180 2.180 0.730 2.410 ;
        RECT 0.410 2.130 0.730 2.180 ;
        RECT 0.410 1.630 0.730 1.950 ;
        RECT 1.710 1.530 2.030 1.850 ;
        RECT 0.410 1.450 0.730 1.490 ;
        RECT 0.180 1.220 0.730 1.450 ;
        RECT 0.410 1.170 0.730 1.220 ;
        RECT 0.410 0.670 0.730 0.990 ;
        RECT 1.710 0.570 2.030 0.890 ;
        RECT 0.410 0.490 0.730 0.530 ;
        RECT 0.180 0.260 0.730 0.490 ;
        RECT 0.410 0.210 0.730 0.260 ;
      LAYER via ;
        RECT 0.630 5.440 0.890 5.700 ;
        RECT 1.720 5.450 1.980 5.710 ;
        RECT 0.160 5.030 0.420 5.290 ;
        RECT 0.630 4.520 0.890 4.780 ;
        RECT 1.720 4.530 1.980 4.790 ;
        RECT 0.160 4.110 0.420 4.370 ;
        RECT 0.630 3.600 0.890 3.860 ;
        RECT 1.720 3.610 1.980 3.870 ;
        RECT 0.160 3.190 0.420 3.450 ;
        RECT 0.440 2.620 0.700 2.880 ;
        RECT 1.740 2.520 2.000 2.780 ;
        RECT 0.440 2.160 0.700 2.420 ;
        RECT 0.440 1.660 0.700 1.920 ;
        RECT 1.740 1.560 2.000 1.820 ;
        RECT 0.440 1.200 0.700 1.460 ;
        RECT 0.440 0.700 0.700 0.960 ;
        RECT 1.740 0.600 2.000 0.860 ;
        RECT 0.440 0.240 0.700 0.500 ;
  END
END sky130_hilas_Trans4small

MACRO sky130_hilas_FGBiasWeakGate2x1cell
  CLASS CORE ;
  FOREIGN sky130_hilas_FGBiasWeakGate2x1cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.530 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.105400 ;
    PORT
      LAYER met2 ;
        RECT 9.050 5.550 9.360 5.560 ;
        RECT 0.000 5.370 11.530 5.550 ;
        RECT 9.050 5.230 9.360 5.370 ;
    END
  END DRAIN1
  PIN VIN11
    PORT
      LAYER met2 ;
        RECT 1.940 4.960 2.250 5.010 ;
        RECT 1.790 4.950 2.250 4.960 ;
        RECT 0.000 4.770 2.250 4.950 ;
        RECT 1.940 4.680 2.250 4.770 ;
    END
  END VIN11
  PIN ROW1
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 9.200 4.530 9.510 4.600 ;
        RECT 9.200 4.520 11.530 4.530 ;
        RECT 0.000 4.310 11.530 4.520 ;
        RECT 0.000 4.300 10.220 4.310 ;
        RECT 9.200 4.270 9.510 4.300 ;
    END
  END ROW1
  PIN ROW2
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 9.200 1.770 9.510 1.840 ;
        RECT 0.000 1.560 11.530 1.770 ;
        RECT 0.000 1.550 10.220 1.560 ;
        RECT 9.200 1.510 9.510 1.550 ;
    END
  END ROW2
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 8.220 0.010 11.530 6.040 ;
      LAYER met1 ;
        RECT 11.010 5.400 11.290 6.050 ;
        RECT 10.900 4.800 11.290 5.400 ;
        RECT 11.010 1.250 11.290 4.800 ;
        RECT 10.900 0.650 11.290 1.250 ;
        RECT 11.010 0.000 11.290 0.650 ;
    END
  END VINJ
  PIN COLSEL1
    USE ANALOG ;
    ANTENNAGATEAREA 0.310000 ;
    PORT
      LAYER met1 ;
        RECT 10.570 4.590 10.760 6.050 ;
        RECT 10.570 4.560 10.790 4.590 ;
        RECT 10.550 4.290 10.800 4.560 ;
        RECT 10.560 4.280 10.800 4.290 ;
        RECT 10.560 4.040 10.790 4.280 ;
        RECT 10.600 2.010 10.760 4.040 ;
        RECT 10.560 1.770 10.790 2.010 ;
        RECT 10.560 1.760 10.800 1.770 ;
        RECT 10.550 1.490 10.800 1.760 ;
        RECT 10.570 1.460 10.790 1.490 ;
        RECT 10.570 0.000 10.760 1.460 ;
    END
  END COLSEL1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2.830 5.080 3.060 6.050 ;
        RECT 2.830 4.830 3.070 5.080 ;
        RECT 2.830 0.000 3.060 4.830 ;
    END
  END VGND
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT 3.770 3.660 6.490 5.310 ;
        RECT 3.770 3.620 6.480 3.660 ;
        RECT 3.770 2.290 6.480 2.330 ;
        RECT 3.770 0.640 6.490 2.290 ;
      LAYER met1 ;
        RECT 4.050 4.840 4.280 6.050 ;
        RECT 4.050 4.050 4.310 4.840 ;
        RECT 4.050 1.900 4.280 4.050 ;
        RECT 4.050 1.110 4.310 1.900 ;
        RECT 4.050 0.000 4.280 1.110 ;
    END
  END GATE1
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 2.516100 ;
    PORT
      LAYER nwell ;
        RECT 0.010 5.300 1.740 6.050 ;
        RECT 0.010 1.730 1.750 5.300 ;
        RECT 0.010 0.010 1.740 1.730 ;
      LAYER met1 ;
        RECT 0.350 0.010 0.770 6.050 ;
    END
  END VTUN
  PIN DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.105400 ;
    PORT
      LAYER met2 ;
        RECT 9.050 0.680 9.360 0.820 ;
        RECT 9.050 0.670 11.530 0.680 ;
        RECT 0.000 0.520 11.530 0.670 ;
        RECT 9.050 0.500 11.530 0.520 ;
        RECT 9.050 0.490 9.360 0.500 ;
    END
  END DRAIN2
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 1.240 2.220 1.320 ;
        RECT 0.000 1.030 2.220 1.240 ;
        RECT 1.910 0.990 2.220 1.030 ;
    END
  END VIN12
  PIN COMMONSOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 1.030400 ;
    PORT
      LAYER met2 ;
        RECT 0.000 3.330 10.460 3.550 ;
        RECT 10.140 3.190 10.460 3.330 ;
        RECT 10.180 2.850 10.440 3.190 ;
        RECT 10.140 2.590 10.460 2.850 ;
    END
  END COMMONSOURCE
  OBS
      LAYER li1 ;
        RECT 1.870 5.040 6.930 5.870 ;
        RECT 9.120 5.470 9.650 5.640 ;
        RECT 10.930 5.370 11.130 5.720 ;
        RECT 10.930 5.340 11.140 5.370 ;
        RECT 1.940 4.960 2.420 5.040 ;
        RECT 1.950 4.710 2.420 4.960 ;
        RECT 7.250 4.890 7.600 5.060 ;
        RECT 8.620 4.890 8.950 5.060 ;
        RECT 0.440 3.910 0.990 4.340 ;
        RECT 4.070 4.100 4.300 4.790 ;
        RECT 9.370 4.560 9.540 5.080 ;
        RECT 9.210 4.300 9.540 4.560 ;
        RECT 7.250 4.100 7.600 4.270 ;
        RECT 8.620 4.100 8.950 4.270 ;
        RECT 3.040 3.080 3.230 3.480 ;
        RECT 7.260 3.310 7.600 3.480 ;
        RECT 8.620 3.310 8.950 3.480 ;
        RECT 9.370 3.390 9.540 4.300 ;
        RECT 10.200 3.480 10.370 5.090 ;
        RECT 10.920 4.760 11.140 5.340 ;
        RECT 10.930 4.750 11.140 4.760 ;
        RECT 10.570 4.580 10.760 4.590 ;
        RECT 10.570 4.290 10.770 4.580 ;
        RECT 10.560 3.960 10.800 4.290 ;
        RECT 2.850 3.070 3.230 3.080 ;
        RECT 2.850 2.890 6.590 3.070 ;
        RECT 2.850 2.850 3.230 2.890 ;
        RECT 0.440 2.180 0.990 2.610 ;
        RECT 3.040 2.470 3.230 2.850 ;
        RECT 8.700 2.740 8.870 3.310 ;
        RECT 10.200 3.290 10.380 3.480 ;
        RECT 7.260 2.570 7.600 2.740 ;
        RECT 8.620 2.570 8.950 2.740 ;
        RECT 1.920 1.030 2.260 1.280 ;
        RECT 4.070 1.160 4.300 1.890 ;
        RECT 7.250 1.780 7.600 1.950 ;
        RECT 8.620 1.780 8.950 1.950 ;
        RECT 9.370 1.800 9.540 2.660 ;
        RECT 9.210 1.540 9.540 1.800 ;
        RECT 1.910 0.950 2.260 1.030 ;
        RECT 7.250 0.990 7.600 1.160 ;
        RECT 8.620 0.990 8.950 1.160 ;
        RECT 9.370 0.970 9.540 1.540 ;
        RECT 10.200 2.570 10.380 2.760 ;
        RECT 10.200 0.960 10.370 2.570 ;
        RECT 10.560 1.760 10.800 2.090 ;
        RECT 10.570 1.470 10.770 1.760 ;
        RECT 10.570 1.460 10.760 1.470 ;
        RECT 10.930 1.290 11.140 1.300 ;
        RECT 1.910 0.100 6.960 0.950 ;
        RECT 10.920 0.710 11.140 1.290 ;
        RECT 10.930 0.680 11.140 0.710 ;
        RECT 9.120 0.410 9.650 0.580 ;
        RECT 10.930 0.330 11.130 0.680 ;
      LAYER mcon ;
        RECT 10.940 5.170 11.110 5.340 ;
        RECT 2.010 4.750 2.180 4.920 ;
        RECT 4.100 4.590 4.270 4.760 ;
        RECT 0.440 3.990 0.710 4.260 ;
        RECT 4.100 4.140 4.270 4.310 ;
        RECT 9.270 4.340 9.440 4.510 ;
        RECT 10.580 4.330 10.760 4.520 ;
        RECT 2.860 2.880 3.030 3.050 ;
        RECT 0.440 2.260 0.710 2.530 ;
        RECT 4.100 1.640 4.270 1.810 ;
        RECT 9.270 1.580 9.440 1.750 ;
        RECT 1.980 1.060 2.150 1.230 ;
        RECT 4.100 1.190 4.270 1.360 ;
        RECT 10.580 1.530 10.760 1.720 ;
        RECT 10.940 0.710 11.110 0.880 ;
      LAYER met1 ;
        RECT 9.050 5.230 9.360 5.670 ;
        RECT 1.940 4.680 2.260 5.000 ;
        RECT 9.200 4.270 9.520 4.590 ;
        RECT 10.170 3.480 10.410 3.610 ;
        RECT 10.170 3.160 10.430 3.480 ;
        RECT 10.170 2.560 10.430 2.880 ;
        RECT 10.170 2.440 10.410 2.560 ;
        RECT 9.200 1.510 9.520 1.830 ;
        RECT 1.910 0.990 2.230 1.310 ;
        RECT 9.050 0.380 9.360 0.820 ;
      LAYER via ;
        RECT 9.080 5.260 9.340 5.520 ;
        RECT 1.970 4.710 2.230 4.970 ;
        RECT 9.230 4.300 9.490 4.560 ;
        RECT 10.170 3.190 10.430 3.450 ;
        RECT 10.170 2.590 10.430 2.850 ;
        RECT 9.230 1.540 9.490 1.800 ;
        RECT 1.940 1.020 2.200 1.280 ;
        RECT 9.080 0.530 9.340 0.790 ;
  END
END sky130_hilas_FGBiasWeakGate2x1cell

MACRO sky130_hilas_swc4x2cell
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x2cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.400 BY 9.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 17.090 5.950 17.470 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.090 0.000 17.470 0.150 ;
    END
  END GATE2
  PIN VTUN
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 11.960 0.000 12.360 0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.040 0.000 13.440 0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.040 5.950 13.440 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.960 5.920 12.360 6.050 ;
    END
  END VTUN
  PIN GATE1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 7.930 5.950 8.310 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 7.930 0.000 8.310 0.090 ;
    END
  END GATE1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 22.240 0.010 22.400 0.070 ;
    END
  END VINJ
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 2.160 5.930 2.470 5.950 ;
        RECT 2.840 5.930 5.690 6.010 ;
        RECT 19.730 5.930 22.560 6.010 ;
        RECT 22.930 5.930 23.240 5.950 ;
        RECT 0.000 5.910 10.060 5.930 ;
        RECT 15.340 5.910 25.400 5.930 ;
        RECT 0.000 5.760 25.400 5.910 ;
        RECT 0.000 5.750 2.560 5.760 ;
        RECT 2.160 5.620 2.470 5.750 ;
        RECT 2.840 5.710 3.260 5.760 ;
        RECT 5.250 5.730 19.930 5.760 ;
        RECT 22.240 5.710 22.560 5.760 ;
        RECT 22.840 5.750 25.400 5.760 ;
        RECT 22.930 5.620 23.240 5.750 ;
        RECT 3.070 5.380 3.390 5.460 ;
        RECT 7.000 5.380 7.320 5.390 ;
        RECT 3.070 5.200 7.320 5.380 ;
        RECT 3.070 5.140 3.390 5.200 ;
        RECT 7.000 5.130 7.320 5.200 ;
        RECT 18.080 5.380 18.400 5.390 ;
        RECT 22.010 5.380 22.330 5.460 ;
        RECT 18.080 5.200 22.330 5.380 ;
        RECT 18.080 5.130 18.400 5.200 ;
        RECT 22.010 5.140 22.330 5.200 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.110 8.710 3.350 9.870 ;
        RECT 3.100 8.050 3.370 8.710 ;
        RECT 3.110 6.050 3.350 8.050 ;
        RECT 3.000 6.010 3.350 6.050 ;
        RECT 2.840 5.710 3.350 6.010 ;
        RECT 3.110 5.460 3.350 5.710 ;
        RECT 3.100 5.140 3.360 5.460 ;
        RECT 3.110 3.820 3.350 5.140 ;
      LAYER via ;
        RECT 2.870 5.730 3.130 5.990 ;
        RECT 3.100 5.170 3.360 5.430 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.000 0.000 3.160 0.060 ;
    END
  END VINJ
  PIN GATESELECT1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 3.410 6.000 3.600 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.410 0.010 3.600 0.070 ;
    END
  END GATESELECT1
  PIN GATESELECT2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 21.800 0.010 21.990 0.070 ;
    END
  END GATESELECT2
  PIN COL1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 3.810 6.000 3.970 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.810 0.010 3.970 0.070 ;
    END
  END COL1
  PIN COL2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 21.430 0.010 21.590 0.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.430 6.000 21.590 6.050 ;
    END
  END COL2
  PIN ROW1
    USE ANALOG ;
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 2.160 4.950 2.470 5.070 ;
        RECT 2.640 4.950 2.780 5.130 ;
        RECT 2.160 4.940 10.060 4.950 ;
        RECT 0.000 4.780 10.060 4.940 ;
        RECT 0.000 4.760 2.560 4.780 ;
        RECT 2.160 4.740 2.470 4.760 ;
        RECT 7.740 4.690 9.280 4.780 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.670 4.950 22.760 5.120 ;
        RECT 22.930 4.950 23.240 5.070 ;
        RECT 15.340 4.940 23.240 4.950 ;
        RECT 15.340 4.780 25.400 4.940 ;
        RECT 16.120 4.690 17.660 4.780 ;
        RECT 22.840 4.760 25.400 4.780 ;
        RECT 22.930 4.740 23.240 4.760 ;
    END
  END ROW1
  PIN ROW2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 2.640 3.940 2.790 4.130 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.640 3.940 22.770 4.120 ;
    END
  END ROW2
  PIN DRAIN1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 2.640 5.370 2.780 5.560 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.670 5.370 22.760 5.550 ;
    END
  END DRAIN1
  PIN DRAIN2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 2.640 3.510 2.770 3.690 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.630 3.510 22.770 3.690 ;
    END
  END DRAIN2
  PIN DRAIN3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 2.640 2.360 2.710 2.540 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.680 2.360 22.770 2.540 ;
    END
  END DRAIN3
  PIN ROW3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 2.640 1.930 2.710 2.110 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.680 1.930 22.770 2.110 ;
    END
  END ROW3
  PIN ROW4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 2.640 0.940 2.710 1.120 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.680 0.940 22.770 1.120 ;
    END
  END ROW4
  PIN DRAIN4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 2.640 0.510 2.710 0.690 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.680 0.510 22.770 0.690 ;
    END
  END DRAIN4
  PIN VGND
    PORT
      LAYER met1 ;
        RECT 5.750 5.960 5.990 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.750 0.000 5.990 0.080 ;
    END
    PORT
      LAYER met1 ;
        RECT 9.680 0.000 9.920 0.070 ;
    END
    PORT
      LAYER nwell ;
        RECT 8.340 8.010 10.070 9.870 ;
        RECT 8.340 6.170 10.080 8.010 ;
        RECT 8.340 3.820 10.070 6.170 ;
      LAYER met1 ;
        RECT 9.320 6.050 9.720 9.870 ;
        RECT 9.320 5.990 9.920 6.050 ;
        RECT 9.320 3.820 9.720 5.990 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.480 0.000 15.720 0.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.410 0.000 19.650 0.060 ;
    END
    PORT
      LAYER nwell ;
        RECT 15.330 8.010 17.060 9.870 ;
        RECT 15.320 6.170 17.060 8.010 ;
        RECT 15.330 3.820 17.060 6.170 ;
      LAYER met1 ;
        RECT 15.680 6.050 16.080 9.870 ;
        RECT 15.480 6.000 16.080 6.050 ;
        RECT 15.680 3.820 16.080 6.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.410 5.980 19.650 6.050 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 0.010 9.860 2.560 9.870 ;
        RECT 0.000 3.840 2.560 9.860 ;
        RECT 0.010 3.830 2.560 3.840 ;
        RECT 4.090 3.820 6.320 9.870 ;
        RECT 19.080 3.820 21.310 9.870 ;
        RECT 22.840 9.860 25.390 9.870 ;
        RECT 22.840 3.840 25.400 9.860 ;
        RECT 22.840 3.830 25.390 3.840 ;
      LAYER li1 ;
        RECT 0.400 9.190 0.600 9.540 ;
        RECT 2.140 9.460 2.460 9.470 ;
        RECT 1.880 9.290 2.460 9.460 ;
        RECT 2.130 9.240 2.460 9.290 ;
        RECT 2.140 9.210 2.460 9.240 ;
        RECT 22.940 9.460 23.260 9.470 ;
        RECT 22.940 9.290 23.520 9.460 ;
        RECT 22.940 9.240 23.270 9.290 ;
        RECT 22.940 9.210 23.260 9.240 ;
        RECT 0.390 9.160 0.600 9.190 ;
        RECT 24.800 9.190 25.000 9.540 ;
        RECT 0.390 8.570 0.610 9.160 ;
        RECT 1.130 8.600 1.330 9.170 ;
        RECT 2.140 8.880 2.460 8.920 ;
        RECT 2.130 8.840 2.460 8.880 ;
        RECT 1.880 8.670 2.460 8.840 ;
        RECT 2.140 8.660 2.460 8.670 ;
        RECT 22.940 8.880 23.260 8.920 ;
        RECT 22.940 8.840 23.270 8.880 ;
        RECT 22.940 8.670 23.520 8.840 ;
        RECT 22.940 8.660 23.260 8.670 ;
        RECT 0.390 7.540 0.610 8.130 ;
        RECT 3.140 8.110 3.310 8.620 ;
        RECT 7.080 8.120 7.250 8.630 ;
        RECT 18.150 8.120 18.320 8.630 ;
        RECT 22.090 8.110 22.260 8.620 ;
        RECT 24.070 8.600 24.270 9.170 ;
        RECT 24.800 9.160 25.010 9.190 ;
        RECT 24.790 8.570 25.010 9.160 ;
        RECT 0.390 7.510 0.600 7.540 ;
        RECT 1.130 7.530 1.330 8.100 ;
        RECT 2.140 8.030 2.460 8.040 ;
        RECT 1.880 7.860 2.460 8.030 ;
        RECT 2.130 7.820 2.460 7.860 ;
        RECT 2.140 7.780 2.460 7.820 ;
        RECT 22.940 8.030 23.260 8.040 ;
        RECT 22.940 7.860 23.520 8.030 ;
        RECT 22.940 7.820 23.270 7.860 ;
        RECT 22.940 7.780 23.260 7.820 ;
        RECT 24.070 7.530 24.270 8.100 ;
        RECT 24.790 7.540 25.010 8.130 ;
        RECT 0.400 7.160 0.600 7.510 ;
        RECT 24.800 7.510 25.010 7.540 ;
        RECT 2.140 7.460 2.460 7.490 ;
        RECT 2.130 7.410 2.460 7.460 ;
        RECT 22.940 7.460 23.260 7.490 ;
        RECT 1.880 7.240 2.460 7.410 ;
        RECT 2.140 7.230 2.460 7.240 ;
        RECT 0.770 6.760 1.210 6.930 ;
        RECT 0.400 6.180 0.600 6.530 ;
        RECT 2.140 6.450 2.460 6.460 ;
        RECT 1.880 6.280 2.460 6.450 ;
        RECT 2.130 6.230 2.460 6.280 ;
        RECT 3.140 6.270 3.310 7.280 ;
        RECT 5.070 6.550 5.620 6.980 ;
        RECT 7.070 6.410 7.240 7.420 ;
        RECT 9.100 6.620 9.650 7.050 ;
        RECT 15.750 6.620 16.300 7.050 ;
        RECT 18.160 6.410 18.330 7.420 ;
        RECT 22.940 7.410 23.270 7.460 ;
        RECT 19.780 6.550 20.330 6.980 ;
        RECT 22.090 6.270 22.260 7.280 ;
        RECT 22.940 7.240 23.520 7.410 ;
        RECT 22.940 7.230 23.260 7.240 ;
        RECT 24.800 7.160 25.000 7.510 ;
        RECT 24.190 6.760 24.630 6.930 ;
        RECT 22.940 6.450 23.260 6.460 ;
        RECT 22.940 6.280 23.520 6.450 ;
        RECT 2.140 6.200 2.460 6.230 ;
        RECT 22.940 6.230 23.270 6.280 ;
        RECT 22.940 6.200 23.260 6.230 ;
        RECT 0.390 6.150 0.600 6.180 ;
        RECT 24.800 6.180 25.000 6.530 ;
        RECT 0.390 5.560 0.610 6.150 ;
        RECT 1.130 5.590 1.330 6.160 ;
        RECT 2.140 5.870 2.460 5.910 ;
        RECT 2.130 5.830 2.460 5.870 ;
        RECT 1.880 5.660 2.460 5.830 ;
        RECT 2.140 5.650 2.460 5.660 ;
        RECT 22.940 5.870 23.260 5.910 ;
        RECT 22.940 5.830 23.270 5.870 ;
        RECT 22.940 5.660 23.520 5.830 ;
        RECT 22.940 5.650 23.260 5.660 ;
        RECT 24.070 5.590 24.270 6.160 ;
        RECT 24.800 6.150 25.010 6.180 ;
        RECT 24.790 5.560 25.010 6.150 ;
        RECT 0.390 4.540 0.610 5.130 ;
        RECT 0.390 4.510 0.600 4.540 ;
        RECT 1.130 4.530 1.330 5.100 ;
        RECT 2.140 5.030 2.460 5.040 ;
        RECT 1.880 4.860 2.460 5.030 ;
        RECT 2.130 4.820 2.460 4.860 ;
        RECT 2.140 4.780 2.460 4.820 ;
        RECT 22.940 5.030 23.260 5.040 ;
        RECT 22.940 4.860 23.520 5.030 ;
        RECT 22.940 4.820 23.270 4.860 ;
        RECT 22.940 4.780 23.260 4.820 ;
        RECT 24.070 4.530 24.270 5.100 ;
        RECT 24.790 4.540 25.010 5.130 ;
        RECT 0.400 4.160 0.600 4.510 ;
        RECT 24.800 4.510 25.010 4.540 ;
        RECT 2.140 4.460 2.460 4.490 ;
        RECT 2.130 4.410 2.460 4.460 ;
        RECT 1.880 4.240 2.460 4.410 ;
        RECT 2.140 4.230 2.460 4.240 ;
        RECT 22.940 4.460 23.260 4.490 ;
        RECT 22.940 4.410 23.270 4.460 ;
        RECT 22.940 4.240 23.520 4.410 ;
        RECT 22.940 4.230 23.260 4.240 ;
        RECT 24.800 4.160 25.000 4.510 ;
      LAYER mcon ;
        RECT 2.230 9.250 2.400 9.420 ;
        RECT 23.000 9.250 23.170 9.420 ;
        RECT 0.420 8.990 0.590 9.160 ;
        RECT 1.150 8.960 1.320 9.130 ;
        RECT 24.080 8.960 24.250 9.130 ;
        RECT 2.230 8.700 2.400 8.870 ;
        RECT 23.000 8.700 23.170 8.870 ;
        RECT 3.140 8.450 3.310 8.620 ;
        RECT 7.080 8.460 7.250 8.630 ;
        RECT 18.150 8.460 18.320 8.630 ;
        RECT 22.090 8.450 22.260 8.620 ;
        RECT 24.810 8.990 24.980 9.160 ;
        RECT 0.420 7.540 0.590 7.710 ;
        RECT 2.230 7.830 2.400 8.000 ;
        RECT 23.000 7.830 23.170 8.000 ;
        RECT 1.150 7.570 1.320 7.740 ;
        RECT 24.080 7.570 24.250 7.740 ;
        RECT 24.810 7.540 24.980 7.710 ;
        RECT 2.230 7.280 2.400 7.450 ;
        RECT 3.140 6.860 3.310 7.030 ;
        RECT 7.070 7.000 7.240 7.170 ;
        RECT 23.000 7.280 23.170 7.450 ;
        RECT 3.140 6.520 3.310 6.690 ;
        RECT 5.350 6.630 5.620 6.900 ;
        RECT 7.070 6.660 7.240 6.830 ;
        RECT 2.230 6.240 2.400 6.410 ;
        RECT 9.380 6.700 9.650 6.970 ;
        RECT 15.750 6.700 16.020 6.970 ;
        RECT 18.160 7.000 18.330 7.170 ;
        RECT 18.160 6.660 18.330 6.830 ;
        RECT 19.780 6.630 20.050 6.900 ;
        RECT 22.090 6.860 22.260 7.030 ;
        RECT 24.450 6.760 24.630 6.930 ;
        RECT 22.090 6.520 22.260 6.690 ;
        RECT 23.000 6.240 23.170 6.410 ;
        RECT 0.420 5.980 0.590 6.150 ;
        RECT 1.150 5.950 1.320 6.120 ;
        RECT 24.080 5.950 24.250 6.120 ;
        RECT 2.230 5.690 2.400 5.860 ;
        RECT 23.000 5.690 23.170 5.860 ;
        RECT 24.810 5.980 24.980 6.150 ;
        RECT 0.420 4.540 0.590 4.710 ;
        RECT 2.230 4.830 2.400 5.000 ;
        RECT 23.000 4.830 23.170 5.000 ;
        RECT 1.150 4.570 1.320 4.740 ;
        RECT 24.080 4.570 24.250 4.740 ;
        RECT 24.810 4.540 24.980 4.710 ;
        RECT 2.230 4.280 2.400 4.450 ;
        RECT 23.000 4.280 23.170 4.450 ;
      LAYER met1 ;
        RECT 0.360 9.220 0.520 9.870 ;
        RECT 0.360 8.670 0.630 9.220 ;
        RECT 0.350 8.620 0.630 8.670 ;
        RECT 0.770 8.880 0.960 9.870 ;
        RECT 1.170 9.190 1.330 9.870 ;
        RECT 1.130 9.170 1.330 9.190 ;
        RECT 2.150 9.180 2.470 9.500 ;
        RECT 1.120 8.930 1.350 9.170 ;
        RECT 0.770 8.760 0.940 8.880 ;
        RECT 0.350 8.530 0.520 8.620 ;
        RECT 0.360 8.170 0.520 8.530 ;
        RECT 0.350 8.080 0.520 8.170 ;
        RECT 0.350 8.030 0.630 8.080 ;
        RECT 0.360 7.480 0.630 8.030 ;
        RECT 0.770 7.940 0.930 8.760 ;
        RECT 1.130 8.710 1.330 8.930 ;
        RECT 1.170 7.990 1.330 8.710 ;
        RECT 2.150 8.630 2.470 8.950 ;
        RECT 0.770 7.820 0.940 7.940 ;
        RECT 0.360 6.210 0.520 7.480 ;
        RECT 0.770 6.960 0.960 7.820 ;
        RECT 1.130 7.770 1.330 7.990 ;
        RECT 1.120 7.530 1.350 7.770 ;
        RECT 2.150 7.750 2.470 8.070 ;
        RECT 5.290 7.950 5.670 9.870 ;
        RECT 7.040 8.690 7.280 9.870 ;
        RECT 18.120 8.690 18.360 9.870 ;
        RECT 7.030 8.030 7.290 8.690 ;
        RECT 18.110 8.030 18.370 8.690 ;
        RECT 1.130 7.510 1.330 7.530 ;
        RECT 0.740 6.730 0.980 6.960 ;
        RECT 0.360 5.660 0.630 6.210 ;
        RECT 0.350 5.610 0.630 5.660 ;
        RECT 0.770 5.870 0.960 6.730 ;
        RECT 1.170 6.180 1.330 7.510 ;
        RECT 2.150 7.200 2.470 7.520 ;
        RECT 1.130 6.160 1.330 6.180 ;
        RECT 2.150 6.170 2.470 6.490 ;
        RECT 1.120 5.920 1.350 6.160 ;
        RECT 5.290 6.090 5.680 7.950 ;
        RECT 0.770 5.750 0.940 5.870 ;
        RECT 0.350 5.520 0.520 5.610 ;
        RECT 0.360 5.170 0.520 5.520 ;
        RECT 0.350 5.080 0.520 5.170 ;
        RECT 0.350 5.030 0.630 5.080 ;
        RECT 0.360 4.480 0.630 5.030 ;
        RECT 0.770 4.940 0.930 5.750 ;
        RECT 1.130 5.700 1.330 5.920 ;
        RECT 1.170 4.990 1.330 5.700 ;
        RECT 2.150 5.620 2.470 5.940 ;
        RECT 0.770 4.820 0.940 4.940 ;
        RECT 0.360 3.830 0.520 4.480 ;
        RECT 0.770 3.830 0.960 4.820 ;
        RECT 1.130 4.770 1.330 4.990 ;
        RECT 1.120 4.530 1.350 4.770 ;
        RECT 2.150 4.750 2.470 5.070 ;
        RECT 1.130 4.510 1.330 4.530 ;
        RECT 1.170 3.830 1.330 4.510 ;
        RECT 2.150 4.200 2.470 4.520 ;
        RECT 5.290 3.820 5.670 6.090 ;
        RECT 7.040 5.420 7.280 8.030 ;
        RECT 12.360 5.690 13.040 5.910 ;
        RECT 18.120 5.420 18.360 8.030 ;
        RECT 19.730 7.950 20.110 9.870 ;
        RECT 22.050 8.710 22.290 9.870 ;
        RECT 22.930 9.180 23.250 9.500 ;
        RECT 24.070 9.190 24.230 9.870 ;
        RECT 24.070 9.170 24.270 9.190 ;
        RECT 22.030 8.050 22.300 8.710 ;
        RECT 22.930 8.630 23.250 8.950 ;
        RECT 24.050 8.930 24.280 9.170 ;
        RECT 24.070 8.710 24.270 8.930 ;
        RECT 24.440 8.880 24.630 9.870 ;
        RECT 24.880 9.220 25.040 9.870 ;
        RECT 24.460 8.760 24.630 8.880 ;
        RECT 19.720 6.090 20.110 7.950 ;
        RECT 7.030 5.100 7.290 5.420 ;
        RECT 18.110 5.100 18.370 5.420 ;
        RECT 7.040 3.820 7.280 5.100 ;
        RECT 18.120 3.820 18.360 5.100 ;
        RECT 19.730 3.820 20.110 6.090 ;
        RECT 22.050 6.050 22.290 8.050 ;
        RECT 22.930 7.750 23.250 8.070 ;
        RECT 24.070 7.990 24.230 8.710 ;
        RECT 24.070 7.770 24.270 7.990 ;
        RECT 24.470 7.940 24.630 8.760 ;
        RECT 24.770 8.670 25.040 9.220 ;
        RECT 24.770 8.620 25.050 8.670 ;
        RECT 24.880 8.530 25.050 8.620 ;
        RECT 24.880 8.170 25.040 8.530 ;
        RECT 24.880 8.080 25.050 8.170 ;
        RECT 24.460 7.820 24.630 7.940 ;
        RECT 24.050 7.530 24.280 7.770 ;
        RECT 22.930 7.200 23.250 7.520 ;
        RECT 24.070 7.510 24.270 7.530 ;
        RECT 22.930 6.170 23.250 6.490 ;
        RECT 24.070 6.180 24.230 7.510 ;
        RECT 24.440 6.960 24.630 7.820 ;
        RECT 24.770 8.030 25.050 8.080 ;
        RECT 24.770 7.480 25.040 8.030 ;
        RECT 24.420 6.730 24.660 6.960 ;
        RECT 24.070 6.160 24.270 6.180 ;
        RECT 21.800 6.000 21.990 6.050 ;
        RECT 22.050 6.010 22.400 6.050 ;
        RECT 22.050 5.710 22.560 6.010 ;
        RECT 22.050 5.460 22.290 5.710 ;
        RECT 22.930 5.620 23.250 5.940 ;
        RECT 24.050 5.920 24.280 6.160 ;
        RECT 24.070 5.700 24.270 5.920 ;
        RECT 24.440 5.870 24.630 6.730 ;
        RECT 24.880 6.210 25.040 7.480 ;
        RECT 24.460 5.750 24.630 5.870 ;
        RECT 22.040 5.140 22.300 5.460 ;
        RECT 22.050 3.820 22.290 5.140 ;
        RECT 22.930 4.750 23.250 5.070 ;
        RECT 24.070 4.990 24.230 5.700 ;
        RECT 24.070 4.770 24.270 4.990 ;
        RECT 24.470 4.940 24.630 5.750 ;
        RECT 24.770 5.660 25.040 6.210 ;
        RECT 24.770 5.610 25.050 5.660 ;
        RECT 24.880 5.520 25.050 5.610 ;
        RECT 24.880 5.170 25.040 5.520 ;
        RECT 24.880 5.080 25.050 5.170 ;
        RECT 24.460 4.820 24.630 4.940 ;
        RECT 24.050 4.530 24.280 4.770 ;
        RECT 22.930 4.200 23.250 4.520 ;
        RECT 24.070 4.510 24.270 4.530 ;
        RECT 24.070 3.830 24.230 4.510 ;
        RECT 24.440 3.830 24.630 4.820 ;
        RECT 24.770 5.030 25.050 5.080 ;
        RECT 24.770 4.480 25.040 5.030 ;
        RECT 24.880 3.830 25.040 4.480 ;
      LAYER via ;
        RECT 2.180 9.210 2.440 9.470 ;
        RECT 2.180 8.660 2.440 8.920 ;
        RECT 2.180 7.780 2.440 8.040 ;
        RECT 2.180 7.230 2.440 7.490 ;
        RECT 2.180 6.200 2.440 6.460 ;
        RECT 2.180 5.650 2.440 5.910 ;
        RECT 2.180 4.780 2.440 5.040 ;
        RECT 2.180 4.230 2.440 4.490 ;
        RECT 22.960 9.210 23.220 9.470 ;
        RECT 22.960 8.660 23.220 8.920 ;
        RECT 7.030 5.130 7.290 5.390 ;
        RECT 18.110 5.130 18.370 5.390 ;
        RECT 22.960 7.780 23.220 8.040 ;
        RECT 22.960 7.230 23.220 7.490 ;
        RECT 22.960 6.200 23.220 6.460 ;
        RECT 22.270 5.730 22.530 5.990 ;
        RECT 22.960 5.650 23.220 5.910 ;
        RECT 22.040 5.170 22.300 5.430 ;
        RECT 22.960 4.780 23.220 5.040 ;
        RECT 22.960 4.230 23.220 4.490 ;
      LAYER met2 ;
        RECT 2.160 9.370 2.470 9.510 ;
        RECT 22.930 9.370 23.240 9.510 ;
        RECT 0.000 9.190 10.070 9.370 ;
        RECT 15.330 9.190 25.400 9.370 ;
        RECT 2.160 9.180 2.470 9.190 ;
        RECT 22.930 9.180 23.240 9.190 ;
        RECT 2.160 8.940 2.470 8.960 ;
        RECT 22.930 8.940 23.240 8.960 ;
        RECT 0.000 8.760 10.070 8.940 ;
        RECT 15.330 8.760 25.400 8.940 ;
        RECT 2.160 8.630 2.470 8.760 ;
        RECT 22.930 8.630 23.240 8.760 ;
        RECT 2.160 7.940 2.470 8.070 ;
        RECT 22.930 7.940 23.240 8.070 ;
        RECT 0.000 7.760 10.080 7.940 ;
        RECT 15.320 7.760 25.400 7.940 ;
        RECT 2.160 7.740 2.470 7.760 ;
        RECT 22.930 7.740 23.240 7.760 ;
        RECT 2.160 7.510 2.470 7.520 ;
        RECT 22.930 7.510 23.240 7.520 ;
        RECT 0.000 7.330 10.080 7.510 ;
        RECT 15.320 7.330 25.400 7.510 ;
        RECT 2.160 7.190 2.470 7.330 ;
        RECT 22.930 7.190 23.240 7.330 ;
        RECT 2.160 6.360 2.470 6.500 ;
        RECT 0.000 6.350 2.470 6.360 ;
        RECT 22.930 6.360 23.240 6.500 ;
        RECT 22.930 6.350 25.400 6.360 ;
        RECT 0.000 6.180 10.060 6.350 ;
        RECT 15.340 6.180 25.400 6.350 ;
        RECT 2.160 6.170 2.470 6.180 ;
        RECT 22.930 6.170 23.240 6.180 ;
        RECT 2.160 4.510 2.470 4.520 ;
        RECT 22.930 4.510 23.240 4.520 ;
        RECT 0.000 4.340 10.060 4.510 ;
        RECT 15.340 4.340 25.400 4.510 ;
        RECT 0.000 4.330 2.470 4.340 ;
        RECT 2.160 4.190 2.470 4.330 ;
        RECT 22.930 4.330 25.400 4.340 ;
        RECT 22.930 4.190 23.240 4.330 ;
        RECT 9.340 1.380 16.100 1.560 ;
  END
END sky130_hilas_swc4x2cell

MACRO sky130_hilas_polyresistorGND
  CLASS CORE ;
  FOREIGN sky130_hilas_polyresistorGND ;
  ORIGIN 0.000 0.000 ;
  SIZE 55.470 BY 10.890 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN INPUT
    PORT
      LAYER met1 ;
        RECT 21.060 10.250 23.470 10.890 ;
        RECT 21.080 8.900 21.490 10.250 ;
    END
  END INPUT
  PIN OUTPUT
    ANTENNADIFFAREA 16.454399 ;
    PORT
      LAYER met2 ;
        RECT 0.000 7.380 55.470 8.770 ;
    END
  END OUTPUT
  PIN VGND
    ANTENNADIFFAREA 16.454399 ;
    PORT
      LAYER met1 ;
        RECT 27.810 9.320 28.220 10.360 ;
        RECT 0.330 8.710 24.700 8.730 ;
        RECT 0.270 8.320 24.700 8.710 ;
        RECT 0.270 0.070 0.680 8.320 ;
        RECT 26.870 0.820 29.230 9.320 ;
        RECT 33.500 8.720 53.790 8.730 ;
        RECT 33.440 8.710 53.790 8.720 ;
        RECT 33.440 8.330 54.730 8.710 ;
        RECT 33.440 8.320 54.700 8.330 ;
        RECT 26.750 0.000 29.230 0.820 ;
      LAYER via ;
        RECT 0.820 8.410 24.620 8.670 ;
        RECT 33.500 8.410 54.360 8.670 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 21.140 9.120 21.360 10.240 ;
        RECT 21.090 8.930 21.420 9.120 ;
        RECT 27.880 8.930 28.120 10.280 ;
        RECT 0.380 8.460 55.120 8.730 ;
        RECT 0.380 8.330 24.720 8.460 ;
        RECT 33.410 8.330 55.120 8.460 ;
        RECT 0.380 0.730 0.550 8.330 ;
        RECT 54.950 1.250 55.120 8.330 ;
        RECT 26.820 0.390 29.030 0.560 ;
      LAYER mcon ;
        RECT 21.170 9.820 21.340 9.990 ;
        RECT 21.170 9.480 21.340 9.650 ;
        RECT 21.170 9.140 21.340 9.310 ;
        RECT 27.920 9.860 28.090 10.030 ;
        RECT 27.920 9.520 28.090 9.690 ;
        RECT 27.920 9.180 28.090 9.350 ;
        RECT 0.720 8.350 24.620 8.520 ;
        RECT 33.500 8.350 54.670 8.520 ;
        RECT 27.160 0.390 27.330 0.560 ;
        RECT 27.500 0.390 27.670 0.560 ;
        RECT 27.840 0.390 28.010 0.560 ;
        RECT 28.180 0.390 28.350 0.560 ;
        RECT 28.520 0.390 28.690 0.560 ;
        RECT 28.860 0.390 29.030 0.560 ;
      LAYER met2 ;
        RECT 0.000 1.080 55.470 2.480 ;
  END
END sky130_hilas_polyresistorGND

MACRO sky130_hilas_swc4x2cellOverlap
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x2cellOverlap ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.790 BY 9.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VERT1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 3.080 5.990 3.240 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.080 0.010 3.240 0.080 ;
    END
  END VERT1
  PIN HORIZ1
    USE ANALOG ;
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met2 ;
        RECT 1.910 4.940 1.990 5.120 ;
        RECT 2.160 4.950 2.470 5.070 ;
        RECT 2.160 4.940 9.350 4.950 ;
        RECT 0.000 4.780 9.350 4.940 ;
        RECT 0.000 4.760 2.560 4.780 ;
        RECT 2.160 4.740 2.470 4.760 ;
    END
    PORT
      LAYER met2 ;
        RECT 19.320 4.950 19.630 5.070 ;
        RECT 12.440 4.940 19.630 4.950 ;
        RECT 19.780 4.940 19.890 5.120 ;
        RECT 12.440 4.780 21.790 4.940 ;
        RECT 19.230 4.760 21.790 4.780 ;
        RECT 19.320 4.740 19.630 4.760 ;
    END
  END HORIZ1
  PIN DRAIN1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 5.370 1.990 5.550 ;
    END
    PORT
      LAYER met2 ;
        RECT 19.770 5.370 19.880 5.550 ;
    END
  END DRAIN1
  PIN HORIZ2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 3.940 1.990 4.120 ;
    END
    PORT
      LAYER met2 ;
        RECT 19.780 3.940 19.890 4.120 ;
    END
  END HORIZ2
  PIN DRAIN2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 3.510 1.990 3.690 ;
    END
    PORT
      LAYER met2 ;
        RECT 19.780 3.510 19.890 3.690 ;
    END
  END DRAIN2
  PIN DRAIN3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 2.360 1.980 2.540 ;
    END
    PORT
      LAYER met2 ;
        RECT 19.770 2.360 19.880 2.540 ;
    END
  END DRAIN3
  PIN HORIZ3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 1.930 1.980 2.110 ;
    END
    PORT
      LAYER met2 ;
        RECT 19.770 1.930 19.880 2.110 ;
    END
  END HORIZ3
  PIN HORIZ4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 0.940 1.980 1.120 ;
    END
    PORT
      LAYER met2 ;
        RECT 19.770 0.940 19.880 1.120 ;
    END
  END HORIZ4
  PIN DRAIN4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 1.910 0.510 1.980 0.690 ;
    END
  END DRAIN4
  PIN VINJ
    PORT
      LAYER met1 ;
        RECT 2.270 5.990 2.430 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.270 0.010 2.430 0.080 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.360 0.010 19.520 0.080 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.360 5.980 19.520 6.050 ;
    END
  END VINJ
  PIN GATESELECT1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 2.680 5.990 2.870 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.680 0.010 2.870 0.080 ;
    END
  END GATESELECT1
  PIN VERT2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 18.550 5.980 18.710 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 18.550 0.010 18.710 0.080 ;
    END
  END VERT2
  PIN GATESELECT2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 18.920 5.980 19.110 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 18.920 0.010 19.110 0.080 ;
    END
  END GATESELECT2
  PIN DRAIN
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 19.770 0.510 19.880 0.690 ;
    END
  END DRAIN
  PIN GATE2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 15.200 0.000 15.440 6.050 ;
    END
  END GATE2
  PIN GATE1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 6.350 0.000 6.600 6.050 ;
    END
  END GATE1
  PIN VTUN
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 9.960 0.000 10.260 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.540 0.000 11.840 6.050 ;
    END
  END VTUN
  OBS
      LAYER nwell ;
        RECT 0.010 9.860 6.560 9.870 ;
        RECT 0.000 3.840 6.560 9.860 ;
        RECT 0.010 3.830 6.560 3.840 ;
        RECT 2.560 3.820 6.560 3.830 ;
        RECT 15.230 9.860 21.780 9.870 ;
        RECT 15.230 3.840 21.790 9.860 ;
        RECT 15.230 3.830 21.780 3.840 ;
        RECT 15.230 3.820 19.230 3.830 ;
      LAYER li1 ;
        RECT 0.400 9.190 0.600 9.540 ;
        RECT 2.140 9.460 2.460 9.470 ;
        RECT 1.880 9.290 2.460 9.460 ;
        RECT 2.130 9.240 2.460 9.290 ;
        RECT 2.140 9.210 2.460 9.240 ;
        RECT 0.390 9.160 0.600 9.190 ;
        RECT 0.390 8.570 0.610 9.160 ;
        RECT 1.130 8.600 1.330 9.170 ;
        RECT 2.140 8.880 2.460 8.920 ;
        RECT 2.130 8.840 2.460 8.880 ;
        RECT 1.880 8.670 2.460 8.840 ;
        RECT 2.140 8.660 2.460 8.670 ;
        RECT 2.900 8.560 6.210 9.540 ;
        RECT 8.120 8.660 8.290 9.550 ;
        RECT 13.500 8.660 13.670 9.550 ;
        RECT 15.580 8.560 18.890 9.540 ;
        RECT 19.330 9.460 19.650 9.470 ;
        RECT 19.330 9.290 19.910 9.460 ;
        RECT 19.330 9.240 19.660 9.290 ;
        RECT 19.330 9.210 19.650 9.240 ;
        RECT 21.190 9.190 21.390 9.540 ;
        RECT 19.330 8.880 19.650 8.920 ;
        RECT 19.330 8.840 19.660 8.880 ;
        RECT 19.330 8.670 19.910 8.840 ;
        RECT 19.330 8.660 19.650 8.670 ;
        RECT 20.460 8.600 20.660 9.170 ;
        RECT 21.190 9.160 21.400 9.190 ;
        RECT 21.180 8.570 21.400 9.160 ;
        RECT 0.390 7.540 0.610 8.130 ;
        RECT 0.390 7.510 0.600 7.540 ;
        RECT 1.130 7.530 1.330 8.100 ;
        RECT 2.140 8.030 2.460 8.040 ;
        RECT 1.880 7.860 2.460 8.030 ;
        RECT 2.130 7.820 2.460 7.860 ;
        RECT 2.140 7.780 2.460 7.820 ;
        RECT 0.400 7.160 0.600 7.510 ;
        RECT 2.140 7.460 2.460 7.490 ;
        RECT 2.130 7.410 2.460 7.460 ;
        RECT 1.880 7.240 2.460 7.410 ;
        RECT 2.140 7.230 2.460 7.240 ;
        RECT 2.900 7.090 6.210 8.070 ;
        RECT 8.120 7.140 8.290 8.030 ;
        RECT 13.500 7.140 13.670 8.030 ;
        RECT 15.580 7.090 18.890 8.070 ;
        RECT 19.330 8.030 19.650 8.040 ;
        RECT 19.330 7.860 19.910 8.030 ;
        RECT 19.330 7.820 19.660 7.860 ;
        RECT 19.330 7.780 19.650 7.820 ;
        RECT 20.460 7.530 20.660 8.100 ;
        RECT 21.180 7.540 21.400 8.130 ;
        RECT 21.190 7.510 21.400 7.540 ;
        RECT 19.330 7.460 19.650 7.490 ;
        RECT 19.330 7.410 19.660 7.460 ;
        RECT 19.330 7.240 19.910 7.410 ;
        RECT 19.330 7.230 19.650 7.240 ;
        RECT 21.190 7.160 21.390 7.510 ;
        RECT 0.770 6.760 1.210 6.930 ;
        RECT 20.580 6.760 21.020 6.930 ;
        RECT 0.400 6.180 0.600 6.530 ;
        RECT 2.140 6.450 2.460 6.460 ;
        RECT 1.880 6.280 2.460 6.450 ;
        RECT 2.130 6.230 2.460 6.280 ;
        RECT 2.140 6.200 2.460 6.230 ;
        RECT 0.390 6.150 0.600 6.180 ;
        RECT 0.390 5.560 0.610 6.150 ;
        RECT 1.130 5.590 1.330 6.160 ;
        RECT 2.140 5.870 2.460 5.910 ;
        RECT 2.130 5.830 2.460 5.870 ;
        RECT 1.880 5.660 2.460 5.830 ;
        RECT 2.140 5.650 2.460 5.660 ;
        RECT 2.900 5.620 6.210 6.600 ;
        RECT 8.120 5.690 8.290 6.580 ;
        RECT 13.500 5.690 13.670 6.580 ;
        RECT 15.580 5.620 18.890 6.600 ;
        RECT 19.330 6.450 19.650 6.460 ;
        RECT 19.330 6.280 19.910 6.450 ;
        RECT 19.330 6.230 19.660 6.280 ;
        RECT 19.330 6.200 19.650 6.230 ;
        RECT 21.190 6.180 21.390 6.530 ;
        RECT 19.330 5.870 19.650 5.910 ;
        RECT 19.330 5.830 19.660 5.870 ;
        RECT 19.330 5.660 19.910 5.830 ;
        RECT 19.330 5.650 19.650 5.660 ;
        RECT 20.460 5.590 20.660 6.160 ;
        RECT 21.190 6.150 21.400 6.180 ;
        RECT 21.180 5.560 21.400 6.150 ;
        RECT 0.390 4.540 0.610 5.130 ;
        RECT 0.390 4.510 0.600 4.540 ;
        RECT 1.130 4.530 1.330 5.100 ;
        RECT 2.140 5.030 2.460 5.040 ;
        RECT 1.880 4.860 2.460 5.030 ;
        RECT 2.130 4.820 2.460 4.860 ;
        RECT 2.140 4.780 2.460 4.820 ;
        RECT 0.400 4.160 0.600 4.510 ;
        RECT 2.140 4.460 2.460 4.490 ;
        RECT 2.130 4.410 2.460 4.460 ;
        RECT 1.880 4.240 2.460 4.410 ;
        RECT 2.140 4.230 2.460 4.240 ;
        RECT 2.900 4.150 6.210 5.130 ;
        RECT 8.120 4.150 8.290 5.040 ;
        RECT 13.500 4.150 13.670 5.040 ;
        RECT 15.580 4.150 18.890 5.130 ;
        RECT 19.330 5.030 19.650 5.040 ;
        RECT 19.330 4.860 19.910 5.030 ;
        RECT 19.330 4.820 19.660 4.860 ;
        RECT 19.330 4.780 19.650 4.820 ;
        RECT 20.460 4.530 20.660 5.100 ;
        RECT 21.180 4.540 21.400 5.130 ;
        RECT 21.190 4.510 21.400 4.540 ;
        RECT 19.330 4.460 19.650 4.490 ;
        RECT 19.330 4.410 19.660 4.460 ;
        RECT 19.330 4.240 19.910 4.410 ;
        RECT 19.330 4.230 19.650 4.240 ;
        RECT 21.190 4.160 21.390 4.510 ;
      LAYER mcon ;
        RECT 2.230 9.250 2.400 9.420 ;
        RECT 4.470 9.310 4.640 9.480 ;
        RECT 0.420 8.990 0.590 9.160 ;
        RECT 1.150 8.960 1.320 9.130 ;
        RECT 4.470 8.960 4.640 9.130 ;
        RECT 2.230 8.700 2.400 8.870 ;
        RECT 4.470 8.620 4.640 8.790 ;
        RECT 8.120 9.350 8.290 9.520 ;
        RECT 13.500 9.350 13.670 9.520 ;
        RECT 17.150 9.310 17.320 9.480 ;
        RECT 19.390 9.250 19.560 9.420 ;
        RECT 17.150 8.960 17.320 9.130 ;
        RECT 20.470 8.960 20.640 9.130 ;
        RECT 17.150 8.620 17.320 8.790 ;
        RECT 19.390 8.700 19.560 8.870 ;
        RECT 21.200 8.990 21.370 9.160 ;
        RECT 0.420 7.540 0.590 7.710 ;
        RECT 2.230 7.830 2.400 8.000 ;
        RECT 4.470 7.840 4.640 8.010 ;
        RECT 1.150 7.570 1.320 7.740 ;
        RECT 4.470 7.490 4.640 7.660 ;
        RECT 2.230 7.280 2.400 7.450 ;
        RECT 4.470 7.150 4.640 7.320 ;
        RECT 8.120 7.830 8.290 8.000 ;
        RECT 13.500 7.830 13.670 8.000 ;
        RECT 17.150 7.840 17.320 8.010 ;
        RECT 19.390 7.830 19.560 8.000 ;
        RECT 17.150 7.490 17.320 7.660 ;
        RECT 20.470 7.570 20.640 7.740 ;
        RECT 21.200 7.540 21.370 7.710 ;
        RECT 17.150 7.150 17.320 7.320 ;
        RECT 19.390 7.280 19.560 7.450 ;
        RECT 20.840 6.760 21.020 6.930 ;
        RECT 2.230 6.240 2.400 6.410 ;
        RECT 4.470 6.370 4.640 6.540 ;
        RECT 0.420 5.980 0.590 6.150 ;
        RECT 1.150 5.950 1.320 6.120 ;
        RECT 4.470 6.020 4.640 6.190 ;
        RECT 2.230 5.690 2.400 5.860 ;
        RECT 4.470 5.680 4.640 5.850 ;
        RECT 8.120 6.380 8.290 6.550 ;
        RECT 13.500 6.380 13.670 6.550 ;
        RECT 17.150 6.370 17.320 6.540 ;
        RECT 19.390 6.240 19.560 6.410 ;
        RECT 17.150 6.020 17.320 6.190 ;
        RECT 20.470 5.950 20.640 6.120 ;
        RECT 17.150 5.680 17.320 5.850 ;
        RECT 19.390 5.690 19.560 5.860 ;
        RECT 21.200 5.980 21.370 6.150 ;
        RECT 0.420 4.540 0.590 4.710 ;
        RECT 2.230 4.830 2.400 5.000 ;
        RECT 4.470 4.900 4.640 5.070 ;
        RECT 1.150 4.570 1.320 4.740 ;
        RECT 4.470 4.550 4.640 4.720 ;
        RECT 2.230 4.280 2.400 4.450 ;
        RECT 4.470 4.210 4.640 4.380 ;
        RECT 8.120 4.840 8.290 5.010 ;
        RECT 13.500 4.840 13.670 5.010 ;
        RECT 17.150 4.900 17.320 5.070 ;
        RECT 19.390 4.830 19.560 5.000 ;
        RECT 17.150 4.550 17.320 4.720 ;
        RECT 20.470 4.570 20.640 4.740 ;
        RECT 21.200 4.540 21.370 4.710 ;
        RECT 17.150 4.210 17.320 4.380 ;
        RECT 19.390 4.280 19.560 4.450 ;
      LAYER met1 ;
        RECT 0.360 9.220 0.520 9.870 ;
        RECT 0.360 8.670 0.630 9.220 ;
        RECT 0.350 8.620 0.630 8.670 ;
        RECT 0.770 8.880 0.960 9.870 ;
        RECT 1.170 9.190 1.330 9.870 ;
        RECT 1.130 9.170 1.330 9.190 ;
        RECT 2.150 9.180 2.470 9.500 ;
        RECT 1.120 8.930 1.350 9.170 ;
        RECT 0.770 8.760 0.940 8.880 ;
        RECT 0.350 8.530 0.520 8.620 ;
        RECT 0.360 8.170 0.520 8.530 ;
        RECT 0.350 8.080 0.520 8.170 ;
        RECT 0.350 8.030 0.630 8.080 ;
        RECT 0.360 7.480 0.630 8.030 ;
        RECT 0.770 7.940 0.930 8.760 ;
        RECT 1.130 8.710 1.330 8.930 ;
        RECT 1.170 7.990 1.330 8.710 ;
        RECT 2.150 8.630 2.470 8.950 ;
        RECT 4.440 8.900 4.680 9.540 ;
        RECT 4.440 8.640 4.670 8.900 ;
        RECT 4.430 8.420 4.670 8.640 ;
        RECT 0.770 7.820 0.940 7.940 ;
        RECT 0.360 6.210 0.520 7.480 ;
        RECT 0.770 6.960 0.960 7.820 ;
        RECT 1.130 7.770 1.330 7.990 ;
        RECT 1.120 7.530 1.350 7.770 ;
        RECT 2.150 7.750 2.470 8.070 ;
        RECT 1.130 7.510 1.330 7.530 ;
        RECT 0.740 6.730 0.980 6.960 ;
        RECT 0.360 5.660 0.630 6.210 ;
        RECT 0.350 5.610 0.630 5.660 ;
        RECT 0.770 5.870 0.960 6.730 ;
        RECT 1.170 6.180 1.330 7.510 ;
        RECT 2.150 7.200 2.470 7.520 ;
        RECT 4.440 7.430 4.680 8.070 ;
        RECT 4.440 7.170 4.670 7.430 ;
        RECT 4.430 6.950 4.670 7.170 ;
        RECT 1.130 6.160 1.330 6.180 ;
        RECT 2.150 6.170 2.470 6.490 ;
        RECT 1.120 5.920 1.350 6.160 ;
        RECT 4.440 5.960 4.680 6.600 ;
        RECT 0.770 5.750 0.940 5.870 ;
        RECT 0.350 5.520 0.520 5.610 ;
        RECT 0.360 5.170 0.520 5.520 ;
        RECT 0.350 5.080 0.520 5.170 ;
        RECT 0.350 5.030 0.630 5.080 ;
        RECT 0.360 4.480 0.630 5.030 ;
        RECT 0.770 4.940 0.930 5.750 ;
        RECT 1.130 5.700 1.330 5.920 ;
        RECT 1.170 4.990 1.330 5.700 ;
        RECT 2.150 5.620 2.470 5.940 ;
        RECT 4.440 5.700 4.670 5.960 ;
        RECT 4.430 5.480 4.670 5.700 ;
        RECT 0.770 4.820 0.940 4.940 ;
        RECT 0.360 3.830 0.520 4.480 ;
        RECT 0.770 3.830 0.960 4.820 ;
        RECT 1.130 4.770 1.330 4.990 ;
        RECT 1.120 4.530 1.350 4.770 ;
        RECT 2.150 4.750 2.470 5.070 ;
        RECT 1.130 4.510 1.330 4.530 ;
        RECT 1.170 3.830 1.330 4.510 ;
        RECT 2.150 4.200 2.470 4.520 ;
        RECT 4.440 4.490 4.680 5.130 ;
        RECT 4.440 4.230 4.670 4.490 ;
        RECT 4.430 4.010 4.670 4.230 ;
        RECT 8.070 3.820 8.340 9.870 ;
        RECT 13.450 3.820 13.720 9.870 ;
        RECT 17.110 8.900 17.350 9.540 ;
        RECT 19.320 9.180 19.640 9.500 ;
        RECT 20.460 9.190 20.620 9.870 ;
        RECT 20.460 9.170 20.660 9.190 ;
        RECT 17.120 8.640 17.350 8.900 ;
        RECT 17.120 8.420 17.360 8.640 ;
        RECT 19.320 8.630 19.640 8.950 ;
        RECT 20.440 8.930 20.670 9.170 ;
        RECT 20.460 8.710 20.660 8.930 ;
        RECT 20.830 8.880 21.020 9.870 ;
        RECT 21.270 9.220 21.430 9.870 ;
        RECT 20.850 8.760 21.020 8.880 ;
        RECT 17.110 7.430 17.350 8.070 ;
        RECT 19.320 7.750 19.640 8.070 ;
        RECT 20.460 7.990 20.620 8.710 ;
        RECT 20.460 7.770 20.660 7.990 ;
        RECT 20.860 7.940 21.020 8.760 ;
        RECT 21.160 8.670 21.430 9.220 ;
        RECT 21.160 8.620 21.440 8.670 ;
        RECT 21.270 8.530 21.440 8.620 ;
        RECT 21.270 8.170 21.430 8.530 ;
        RECT 21.270 8.080 21.440 8.170 ;
        RECT 20.850 7.820 21.020 7.940 ;
        RECT 20.440 7.530 20.670 7.770 ;
        RECT 17.120 7.170 17.350 7.430 ;
        RECT 19.320 7.200 19.640 7.520 ;
        RECT 20.460 7.510 20.660 7.530 ;
        RECT 17.120 6.950 17.360 7.170 ;
        RECT 17.110 5.960 17.350 6.600 ;
        RECT 19.320 6.170 19.640 6.490 ;
        RECT 20.460 6.180 20.620 7.510 ;
        RECT 20.830 6.960 21.020 7.820 ;
        RECT 21.160 8.030 21.440 8.080 ;
        RECT 21.160 7.480 21.430 8.030 ;
        RECT 20.810 6.730 21.050 6.960 ;
        RECT 20.460 6.160 20.660 6.180 ;
        RECT 17.120 5.700 17.350 5.960 ;
        RECT 17.120 5.480 17.360 5.700 ;
        RECT 19.320 5.620 19.640 5.940 ;
        RECT 20.440 5.920 20.670 6.160 ;
        RECT 20.460 5.700 20.660 5.920 ;
        RECT 20.830 5.870 21.020 6.730 ;
        RECT 21.270 6.210 21.430 7.480 ;
        RECT 20.850 5.750 21.020 5.870 ;
        RECT 17.110 4.490 17.350 5.130 ;
        RECT 19.320 4.750 19.640 5.070 ;
        RECT 20.460 4.990 20.620 5.700 ;
        RECT 20.460 4.770 20.660 4.990 ;
        RECT 20.860 4.940 21.020 5.750 ;
        RECT 21.160 5.660 21.430 6.210 ;
        RECT 21.160 5.610 21.440 5.660 ;
        RECT 21.270 5.520 21.440 5.610 ;
        RECT 21.270 5.170 21.430 5.520 ;
        RECT 21.270 5.080 21.440 5.170 ;
        RECT 20.850 4.820 21.020 4.940 ;
        RECT 20.440 4.530 20.670 4.770 ;
        RECT 17.120 4.230 17.350 4.490 ;
        RECT 17.120 4.010 17.360 4.230 ;
        RECT 19.320 4.200 19.640 4.520 ;
        RECT 20.460 4.510 20.660 4.530 ;
        RECT 20.460 3.830 20.620 4.510 ;
        RECT 20.830 3.830 21.020 4.820 ;
        RECT 21.160 5.030 21.440 5.080 ;
        RECT 21.160 4.480 21.430 5.030 ;
        RECT 21.270 3.830 21.430 4.480 ;
      LAYER via ;
        RECT 2.180 9.210 2.440 9.470 ;
        RECT 2.180 8.660 2.440 8.920 ;
        RECT 2.180 7.780 2.440 8.040 ;
        RECT 2.180 7.230 2.440 7.490 ;
        RECT 2.180 6.200 2.440 6.460 ;
        RECT 2.180 5.650 2.440 5.910 ;
        RECT 2.180 4.780 2.440 5.040 ;
        RECT 2.180 4.230 2.440 4.490 ;
        RECT 19.350 9.210 19.610 9.470 ;
        RECT 19.350 8.660 19.610 8.920 ;
        RECT 19.350 7.780 19.610 8.040 ;
        RECT 19.350 7.230 19.610 7.490 ;
        RECT 19.350 6.200 19.610 6.460 ;
        RECT 19.350 5.650 19.610 5.910 ;
        RECT 19.350 4.780 19.610 5.040 ;
        RECT 19.350 4.230 19.610 4.490 ;
      LAYER met2 ;
        RECT 2.160 9.370 2.470 9.510 ;
        RECT 19.320 9.370 19.630 9.510 ;
        RECT 0.000 9.190 9.350 9.370 ;
        RECT 12.440 9.190 21.790 9.370 ;
        RECT 2.160 9.180 2.470 9.190 ;
        RECT 19.320 9.180 19.630 9.190 ;
        RECT 2.160 8.940 2.470 8.960 ;
        RECT 19.320 8.940 19.630 8.960 ;
        RECT 0.000 8.760 9.350 8.940 ;
        RECT 12.440 8.760 21.790 8.940 ;
        RECT 2.160 8.630 2.470 8.760 ;
        RECT 19.320 8.630 19.630 8.760 ;
        RECT 2.160 7.940 2.470 8.070 ;
        RECT 19.320 7.940 19.630 8.070 ;
        RECT 0.000 7.760 9.350 7.940 ;
        RECT 12.440 7.760 21.790 7.940 ;
        RECT 2.160 7.740 2.470 7.760 ;
        RECT 19.320 7.740 19.630 7.760 ;
        RECT 2.160 7.510 2.470 7.520 ;
        RECT 19.320 7.510 19.630 7.520 ;
        RECT 0.000 7.440 2.470 7.510 ;
        RECT 2.480 7.440 9.350 7.510 ;
        RECT 0.000 7.330 9.350 7.440 ;
        RECT 12.440 7.440 19.310 7.510 ;
        RECT 19.320 7.440 21.790 7.510 ;
        RECT 12.440 7.330 21.790 7.440 ;
        RECT 2.160 7.190 2.470 7.330 ;
        RECT 19.320 7.190 19.630 7.330 ;
        RECT 2.160 6.360 2.470 6.500 ;
        RECT 0.000 6.350 2.470 6.360 ;
        RECT 19.320 6.360 19.630 6.500 ;
        RECT 19.320 6.350 21.790 6.360 ;
        RECT 0.000 6.180 9.350 6.350 ;
        RECT 12.440 6.180 21.790 6.350 ;
        RECT 2.160 6.170 2.470 6.180 ;
        RECT 19.320 6.170 19.630 6.180 ;
        RECT 2.160 5.930 2.470 5.950 ;
        RECT 19.320 5.930 19.630 5.950 ;
        RECT 0.000 5.760 9.350 5.930 ;
        RECT 12.440 5.760 21.790 5.930 ;
        RECT 0.000 5.750 2.560 5.760 ;
        RECT 19.230 5.750 21.790 5.760 ;
        RECT 2.160 5.620 2.470 5.750 ;
        RECT 19.320 5.620 19.630 5.750 ;
        RECT 2.160 4.510 2.470 4.520 ;
        RECT 19.320 4.510 19.630 4.520 ;
        RECT 0.000 4.340 9.350 4.510 ;
        RECT 12.440 4.340 21.790 4.510 ;
        RECT 0.000 4.330 2.470 4.340 ;
        RECT 2.160 4.190 2.470 4.330 ;
        RECT 19.320 4.330 21.790 4.340 ;
        RECT 19.320 4.190 19.630 4.330 ;
        RECT 4.310 3.610 4.430 3.690 ;
        RECT 17.400 3.550 17.520 3.690 ;
  END
END sky130_hilas_swc4x2cellOverlap

MACRO sky130_hilas_FGBias2x1cell
  CLASS CORE ;
  FOREIGN sky130_hilas_FGBias2x1cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.530 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 2.516100 ;
    PORT
      LAYER nwell ;
        RECT 0.010 5.300 1.740 6.050 ;
        RECT 0.010 1.730 1.750 5.300 ;
        RECT 0.010 0.010 1.740 1.730 ;
      LAYER met1 ;
        RECT 0.350 0.000 0.770 6.050 ;
    END
  END VTUN
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2.830 0.000 3.060 6.050 ;
    END
  END VGND
  PIN GATE_CONTROL
    USE ANALOG ;
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT 3.770 3.660 6.490 5.310 ;
        RECT 3.770 3.620 6.480 3.660 ;
        RECT 3.770 2.290 6.480 2.330 ;
        RECT 3.770 0.640 6.490 2.290 ;
      LAYER met1 ;
        RECT 4.050 4.840 4.280 6.050 ;
        RECT 4.050 4.050 4.310 4.840 ;
        RECT 4.050 1.900 4.280 4.050 ;
        RECT 4.050 1.110 4.310 1.900 ;
        RECT 4.050 0.000 4.280 1.110 ;
    END
  END GATE_CONTROL
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.105400 ;
    PORT
      LAYER met2 ;
        RECT 9.050 5.550 9.360 5.560 ;
        RECT 0.000 5.370 11.530 5.550 ;
        RECT 9.050 5.230 9.360 5.370 ;
    END
  END DRAIN1
  PIN DRAIN4
    USE ANALOG ;
    ANTENNADIFFAREA 0.105400 ;
    PORT
      LAYER met2 ;
        RECT 9.050 0.680 9.360 0.820 ;
        RECT 9.050 0.670 11.530 0.680 ;
        RECT 0.000 0.520 11.530 0.670 ;
        RECT 9.050 0.500 11.530 0.520 ;
        RECT 9.050 0.490 9.360 0.500 ;
    END
  END DRAIN4
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 8.220 0.010 11.530 6.050 ;
      LAYER met2 ;
        RECT 10.140 3.190 10.460 3.450 ;
        RECT 10.180 3.170 11.360 3.190 ;
        RECT 10.180 2.910 11.400 3.170 ;
        RECT 10.180 2.850 11.360 2.910 ;
        RECT 10.140 2.840 11.360 2.850 ;
        RECT 10.140 2.590 10.460 2.840 ;
    END
  END VINJ
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 9.200 4.530 9.510 4.600 ;
        RECT 9.200 4.310 11.530 4.530 ;
        RECT 9.200 4.270 9.510 4.310 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 9.200 1.770 9.510 1.840 ;
        RECT 9.200 1.560 11.530 1.770 ;
        RECT 9.200 1.510 9.510 1.560 ;
    END
  END OUTPUT2
  PIN GATECOL
    ANTENNAGATEAREA 0.310000 ;
    PORT
      LAYER met1 ;
        RECT 10.570 4.590 10.760 6.050 ;
        RECT 10.570 4.560 10.790 4.590 ;
        RECT 10.550 4.290 10.800 4.560 ;
        RECT 10.560 4.280 10.800 4.290 ;
        RECT 10.560 4.040 10.790 4.280 ;
        RECT 10.600 2.010 10.760 4.040 ;
        RECT 10.560 1.770 10.790 2.010 ;
        RECT 10.560 1.760 10.800 1.770 ;
        RECT 10.550 1.490 10.800 1.760 ;
        RECT 10.570 1.460 10.790 1.490 ;
        RECT 10.570 0.000 10.760 1.460 ;
    END
  END GATECOL
  PIN VINJ
    ANTENNADIFFAREA 0.510000 ;
    PORT
      LAYER met1 ;
        RECT 11.010 5.400 11.290 6.050 ;
        RECT 10.900 4.800 11.290 5.400 ;
        RECT 11.010 3.200 11.290 4.800 ;
        RECT 11.010 2.880 11.370 3.200 ;
        RECT 11.010 1.250 11.290 2.880 ;
        RECT 10.900 0.650 11.290 1.250 ;
        RECT 11.010 0.000 11.290 0.650 ;
      LAYER via ;
        RECT 11.110 2.910 11.370 3.170 ;
    END
  END VINJ
  OBS
      LAYER li1 ;
        RECT 9.120 5.470 9.650 5.640 ;
        RECT 10.930 5.370 11.130 5.720 ;
        RECT 10.930 5.340 11.140 5.370 ;
        RECT 7.250 4.890 7.600 5.060 ;
        RECT 8.620 4.890 8.950 5.060 ;
        RECT 0.440 3.910 0.990 4.340 ;
        RECT 4.070 4.100 4.300 4.790 ;
        RECT 9.370 4.560 9.540 5.080 ;
        RECT 9.210 4.300 9.540 4.560 ;
        RECT 7.250 4.100 7.600 4.270 ;
        RECT 8.620 4.100 8.950 4.270 ;
        RECT 3.040 3.080 3.230 3.480 ;
        RECT 7.260 3.310 7.600 3.480 ;
        RECT 8.620 3.310 8.950 3.480 ;
        RECT 9.370 3.390 9.540 4.300 ;
        RECT 10.200 3.480 10.370 5.090 ;
        RECT 10.920 4.760 11.140 5.340 ;
        RECT 10.930 4.750 11.140 4.760 ;
        RECT 10.570 4.580 10.760 4.590 ;
        RECT 10.570 4.290 10.770 4.580 ;
        RECT 10.560 3.960 10.800 4.290 ;
        RECT 2.850 3.070 3.230 3.080 ;
        RECT 2.850 2.890 6.590 3.070 ;
        RECT 2.850 2.850 3.230 2.890 ;
        RECT 0.440 2.180 0.990 2.610 ;
        RECT 3.040 2.470 3.230 2.850 ;
        RECT 8.700 2.740 8.870 3.310 ;
        RECT 10.200 3.290 10.380 3.480 ;
        RECT 7.260 2.570 7.600 2.740 ;
        RECT 8.620 2.570 8.950 2.740 ;
        RECT 4.070 1.160 4.300 1.890 ;
        RECT 7.250 1.780 7.600 1.950 ;
        RECT 8.620 1.780 8.950 1.950 ;
        RECT 9.370 1.800 9.540 2.660 ;
        RECT 9.210 1.540 9.540 1.800 ;
        RECT 7.250 0.990 7.600 1.160 ;
        RECT 8.620 0.990 8.950 1.160 ;
        RECT 9.370 0.970 9.540 1.540 ;
        RECT 10.200 2.570 10.380 2.760 ;
        RECT 10.200 0.960 10.370 2.570 ;
        RECT 10.560 1.760 10.800 2.090 ;
        RECT 10.570 1.470 10.770 1.760 ;
        RECT 10.570 1.460 10.760 1.470 ;
        RECT 10.930 1.290 11.140 1.300 ;
        RECT 10.920 0.710 11.140 1.290 ;
        RECT 10.930 0.680 11.140 0.710 ;
        RECT 9.120 0.410 9.650 0.580 ;
        RECT 10.930 0.330 11.130 0.680 ;
      LAYER mcon ;
        RECT 10.940 5.170 11.110 5.340 ;
        RECT 4.100 4.590 4.270 4.760 ;
        RECT 0.440 3.990 0.710 4.260 ;
        RECT 4.100 4.140 4.270 4.310 ;
        RECT 9.270 4.340 9.440 4.510 ;
        RECT 10.580 4.330 10.760 4.520 ;
        RECT 2.860 2.880 3.030 3.050 ;
        RECT 0.440 2.260 0.710 2.530 ;
        RECT 4.100 1.640 4.270 1.810 ;
        RECT 9.270 1.580 9.440 1.750 ;
        RECT 4.100 1.190 4.270 1.360 ;
        RECT 10.580 1.530 10.760 1.720 ;
        RECT 10.940 0.710 11.110 0.880 ;
      LAYER met1 ;
        RECT 9.050 5.230 9.360 5.670 ;
        RECT 9.200 4.270 9.520 4.590 ;
        RECT 10.170 3.480 10.410 3.610 ;
        RECT 10.170 3.160 10.430 3.480 ;
        RECT 10.170 2.560 10.430 2.880 ;
        RECT 10.170 2.440 10.410 2.560 ;
        RECT 9.200 1.510 9.520 1.830 ;
        RECT 9.050 0.380 9.360 0.820 ;
      LAYER via ;
        RECT 9.080 5.260 9.340 5.520 ;
        RECT 9.230 4.300 9.490 4.560 ;
        RECT 10.170 3.190 10.430 3.450 ;
        RECT 10.170 2.590 10.430 2.850 ;
        RECT 9.230 1.540 9.490 1.800 ;
        RECT 9.080 0.530 9.340 0.790 ;
  END
END sky130_hilas_FGBias2x1cell

MACRO sky130_hilas_drainSelect01
  CLASS CORE ;
  FOREIGN sky130_hilas_drainSelect01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.720 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DRAIN4
    ANTENNADIFFAREA 0.275800 ;
    PORT
      LAYER met2 ;
        RECT 0.050 0.690 0.570 0.700 ;
        RECT 0.050 0.620 2.030 0.690 ;
        RECT 0.050 0.570 2.070 0.620 ;
        RECT 4.160 0.570 4.480 0.650 ;
        RECT 0.050 0.520 4.480 0.570 ;
        RECT 1.750 0.380 4.480 0.520 ;
        RECT 1.750 0.360 2.070 0.380 ;
        RECT 4.160 0.330 4.480 0.380 ;
    END
  END DRAIN4
  PIN DRAIN3
    ANTENNADIFFAREA 0.275800 ;
    PORT
      LAYER met2 ;
        RECT 1.750 2.740 2.070 2.760 ;
        RECT 4.160 2.740 4.480 2.790 ;
        RECT 1.750 2.550 4.480 2.740 ;
        RECT 0.050 2.530 0.570 2.540 ;
        RECT 0.050 2.520 1.270 2.530 ;
        RECT 1.750 2.520 2.070 2.550 ;
        RECT 0.050 2.500 2.070 2.520 ;
        RECT 0.050 2.360 2.000 2.500 ;
        RECT 4.160 2.470 4.480 2.550 ;
    END
  END DRAIN3
  PIN DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.275800 ;
    PORT
      LAYER met2 ;
        RECT 0.050 3.670 1.240 3.690 ;
        RECT 0.050 3.550 1.960 3.670 ;
        RECT 0.050 3.510 2.070 3.550 ;
        RECT 1.750 3.500 2.070 3.510 ;
        RECT 4.160 3.500 4.480 3.580 ;
        RECT 1.750 3.310 4.480 3.500 ;
        RECT 1.750 3.290 2.070 3.310 ;
        RECT 4.160 3.260 4.480 3.310 ;
    END
  END DRAIN2
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.275800 ;
    PORT
      LAYER met2 ;
        RECT 1.750 5.670 2.070 5.690 ;
        RECT 4.160 5.670 4.480 5.720 ;
        RECT 0.050 5.540 1.300 5.550 ;
        RECT 1.750 5.540 4.480 5.670 ;
        RECT 0.050 5.480 4.480 5.540 ;
        RECT 0.050 5.430 2.070 5.480 ;
        RECT 0.050 5.380 1.990 5.430 ;
        RECT 4.160 5.400 4.480 5.480 ;
        RECT 0.050 5.370 1.300 5.380 ;
    END
  END DRAIN1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.000 0.000 3.420 6.050 ;
      LAYER met1 ;
        RECT 0.580 5.830 0.830 6.050 ;
        RECT 0.190 4.760 0.830 5.830 ;
        RECT 0.580 4.220 0.830 4.760 ;
        RECT 0.190 3.150 0.830 4.220 ;
        RECT 0.580 2.900 0.830 3.150 ;
        RECT 0.190 1.830 0.830 2.900 ;
        RECT 0.580 1.290 0.830 1.830 ;
        RECT 0.190 0.220 0.830 1.290 ;
        RECT 0.580 0.000 0.830 0.220 ;
    END
  END VINJ
  PIN DRAIN_MUX
    USE ANALOG ;
    ANTENNADIFFAREA 0.719200 ;
    PORT
      LAYER met1 ;
        RECT 3.570 0.000 3.800 6.050 ;
    END
  END DRAIN_MUX
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 4.920 5.830 5.110 6.050 ;
        RECT 4.920 5.340 5.390 5.830 ;
        RECT 4.920 5.080 5.110 5.340 ;
        RECT 4.880 4.790 5.110 5.080 ;
        RECT 4.920 4.190 5.110 4.790 ;
        RECT 4.880 3.900 5.110 4.190 ;
        RECT 4.920 3.640 5.110 3.900 ;
        RECT 4.920 3.150 5.390 3.640 ;
        RECT 4.920 2.900 5.110 3.150 ;
        RECT 4.920 2.410 5.390 2.900 ;
        RECT 4.920 2.150 5.110 2.410 ;
        RECT 4.880 1.860 5.110 2.150 ;
        RECT 4.920 1.260 5.110 1.860 ;
        RECT 4.880 0.970 5.110 1.260 ;
        RECT 4.920 0.710 5.110 0.970 ;
        RECT 4.920 0.220 5.390 0.710 ;
        RECT 4.920 0.000 5.110 0.220 ;
    END
  END VGND
  PIN SELECT4
    ANTENNAGATEAREA 0.625000 ;
    PORT
      LAYER met2 ;
        RECT 5.240 1.090 5.580 1.160 ;
        RECT 5.240 0.860 5.720 1.090 ;
    END
  END SELECT4
  PIN SELECT3
    ANTENNAGATEAREA 0.625000 ;
    PORT
      LAYER met2 ;
        RECT 5.240 2.030 5.720 2.260 ;
        RECT 5.240 1.960 5.580 2.030 ;
    END
  END SELECT3
  PIN SELECT2
    ANTENNAGATEAREA 0.625000 ;
    PORT
      LAYER met2 ;
        RECT 5.240 4.020 5.580 4.090 ;
        RECT 5.240 3.790 5.720 4.020 ;
    END
  END SELECT2
  PIN SELECT1
    ANTENNAGATEAREA 0.625000 ;
    PORT
      LAYER met2 ;
        RECT 5.240 4.960 5.720 5.190 ;
        RECT 5.240 4.890 5.580 4.960 ;
    END
  END SELECT1
  OBS
      LAYER li1 ;
        RECT 0.220 4.920 0.390 5.770 ;
        RECT 0.620 4.790 0.790 5.720 ;
        RECT 4.310 5.650 4.550 5.680 ;
        RECT 1.320 5.480 2.280 5.650 ;
        RECT 2.730 5.480 4.070 5.650 ;
        RECT 4.310 5.480 4.880 5.650 ;
        RECT 1.600 5.470 1.770 5.480 ;
        RECT 4.310 5.440 4.550 5.480 ;
        RECT 5.190 5.350 5.360 5.770 ;
        RECT 1.760 5.030 2.090 5.210 ;
        RECT 5.260 5.130 5.430 5.170 ;
        RECT 4.900 5.030 5.090 5.050 ;
        RECT 1.320 4.860 4.070 5.030 ;
        RECT 4.530 4.860 5.090 5.030 ;
        RECT 4.900 4.820 5.090 4.860 ;
        RECT 5.260 4.960 5.490 5.130 ;
        RECT 5.260 4.610 5.430 4.960 ;
        RECT 0.220 3.210 0.390 4.060 ;
        RECT 0.620 3.260 0.790 4.190 ;
        RECT 4.900 4.120 5.090 4.160 ;
        RECT 1.320 3.950 4.070 4.120 ;
        RECT 4.530 3.950 5.090 4.120 ;
        RECT 1.760 3.770 2.090 3.950 ;
        RECT 4.900 3.930 5.090 3.950 ;
        RECT 5.260 4.020 5.430 4.370 ;
        RECT 5.260 3.850 5.490 4.020 ;
        RECT 5.260 3.810 5.430 3.850 ;
        RECT 1.600 3.500 1.770 3.510 ;
        RECT 4.310 3.500 4.550 3.540 ;
        RECT 1.320 3.330 2.280 3.500 ;
        RECT 2.730 3.330 4.070 3.500 ;
        RECT 4.310 3.330 4.880 3.500 ;
        RECT 4.310 3.300 4.550 3.330 ;
        RECT 5.190 3.210 5.360 3.630 ;
        RECT 0.220 1.990 0.390 2.840 ;
        RECT 0.620 1.860 0.790 2.790 ;
        RECT 4.310 2.720 4.550 2.750 ;
        RECT 1.320 2.550 2.280 2.720 ;
        RECT 2.730 2.550 4.070 2.720 ;
        RECT 4.310 2.550 4.880 2.720 ;
        RECT 1.600 2.540 1.770 2.550 ;
        RECT 4.310 2.510 4.550 2.550 ;
        RECT 5.190 2.420 5.360 2.840 ;
        RECT 1.760 2.100 2.090 2.280 ;
        RECT 5.260 2.200 5.430 2.240 ;
        RECT 4.900 2.100 5.090 2.120 ;
        RECT 1.320 1.930 4.070 2.100 ;
        RECT 4.530 1.930 5.090 2.100 ;
        RECT 4.900 1.890 5.090 1.930 ;
        RECT 5.260 2.030 5.490 2.200 ;
        RECT 5.260 1.680 5.430 2.030 ;
        RECT 0.220 0.280 0.390 1.130 ;
        RECT 0.620 0.330 0.790 1.260 ;
        RECT 4.900 1.190 5.090 1.230 ;
        RECT 1.320 1.020 4.070 1.190 ;
        RECT 4.530 1.020 5.090 1.190 ;
        RECT 1.760 0.840 2.090 1.020 ;
        RECT 4.900 1.000 5.090 1.020 ;
        RECT 5.260 1.090 5.430 1.440 ;
        RECT 5.260 0.920 5.490 1.090 ;
        RECT 5.260 0.880 5.430 0.920 ;
        RECT 1.600 0.570 1.770 0.580 ;
        RECT 4.310 0.570 4.550 0.610 ;
        RECT 1.320 0.400 2.280 0.570 ;
        RECT 2.730 0.400 4.070 0.570 ;
        RECT 4.310 0.400 4.880 0.570 ;
        RECT 4.310 0.370 4.550 0.400 ;
        RECT 5.190 0.280 5.360 0.700 ;
      LAYER mcon ;
        RECT 0.220 5.600 0.390 5.770 ;
        RECT 0.220 5.260 0.390 5.430 ;
        RECT 3.600 5.480 3.770 5.650 ;
        RECT 4.350 5.480 4.520 5.650 ;
        RECT 5.190 5.600 5.360 5.770 ;
        RECT 0.620 5.150 0.790 5.320 ;
        RECT 4.910 4.850 5.080 5.020 ;
        RECT 5.320 4.960 5.490 5.130 ;
        RECT 0.220 3.890 0.390 4.060 ;
        RECT 0.220 3.550 0.390 3.720 ;
        RECT 4.910 3.960 5.080 4.130 ;
        RECT 0.620 3.660 0.790 3.830 ;
        RECT 5.320 3.850 5.490 4.020 ;
        RECT 1.600 3.340 1.770 3.510 ;
        RECT 3.600 3.330 3.770 3.500 ;
        RECT 4.350 3.330 4.520 3.500 ;
        RECT 0.220 2.670 0.390 2.840 ;
        RECT 0.220 2.330 0.390 2.500 ;
        RECT 3.600 2.550 3.770 2.720 ;
        RECT 4.350 2.550 4.520 2.720 ;
        RECT 5.190 2.670 5.360 2.840 ;
        RECT 0.620 2.220 0.790 2.390 ;
        RECT 4.910 1.920 5.080 2.090 ;
        RECT 5.320 2.030 5.490 2.200 ;
        RECT 0.220 0.960 0.390 1.130 ;
        RECT 0.220 0.620 0.390 0.790 ;
        RECT 4.910 1.030 5.080 1.200 ;
        RECT 0.620 0.730 0.790 0.900 ;
        RECT 5.320 0.920 5.490 1.090 ;
        RECT 1.600 0.410 1.770 0.580 ;
        RECT 3.600 0.400 3.770 0.570 ;
        RECT 4.350 0.400 4.520 0.570 ;
      LAYER met1 ;
        RECT 1.730 5.670 2.070 5.720 ;
        RECT 1.510 5.650 2.070 5.670 ;
        RECT 4.160 5.690 4.530 5.710 ;
        RECT 1.510 5.480 2.190 5.650 ;
        RECT 1.510 5.440 2.070 5.480 ;
        RECT 1.730 5.400 2.070 5.440 ;
        RECT 4.160 5.430 4.580 5.690 ;
        RECT 4.160 5.420 4.530 5.430 ;
        RECT 5.250 4.900 5.570 5.180 ;
        RECT 5.250 3.800 5.570 4.080 ;
        RECT 1.730 3.540 2.070 3.580 ;
        RECT 1.510 3.500 2.070 3.540 ;
        RECT 4.160 3.550 4.530 3.560 ;
        RECT 1.510 3.330 2.190 3.500 ;
        RECT 1.510 3.310 2.070 3.330 ;
        RECT 1.730 3.260 2.070 3.310 ;
        RECT 4.160 3.290 4.580 3.550 ;
        RECT 4.160 3.270 4.530 3.290 ;
        RECT 1.730 2.740 2.070 2.790 ;
        RECT 1.510 2.720 2.070 2.740 ;
        RECT 4.160 2.760 4.530 2.780 ;
        RECT 1.510 2.550 2.190 2.720 ;
        RECT 1.510 2.510 2.070 2.550 ;
        RECT 1.730 2.470 2.070 2.510 ;
        RECT 4.160 2.500 4.580 2.760 ;
        RECT 4.160 2.490 4.530 2.500 ;
        RECT 5.250 1.970 5.570 2.250 ;
        RECT 5.250 0.870 5.570 1.150 ;
        RECT 1.730 0.610 2.070 0.650 ;
        RECT 1.510 0.570 2.070 0.610 ;
        RECT 4.160 0.620 4.530 0.630 ;
        RECT 1.510 0.400 2.190 0.570 ;
        RECT 1.510 0.380 2.070 0.400 ;
        RECT 1.730 0.330 2.070 0.380 ;
        RECT 4.160 0.360 4.580 0.620 ;
        RECT 4.160 0.340 4.530 0.360 ;
      LAYER via ;
        RECT 1.780 5.430 2.040 5.690 ;
        RECT 4.190 5.430 4.450 5.690 ;
        RECT 5.280 4.910 5.540 5.170 ;
        RECT 5.280 3.810 5.540 4.070 ;
        RECT 1.780 3.290 2.040 3.550 ;
        RECT 4.190 3.290 4.450 3.550 ;
        RECT 1.780 2.500 2.040 2.760 ;
        RECT 4.190 2.500 4.450 2.760 ;
        RECT 5.280 1.980 5.540 2.240 ;
        RECT 5.280 0.880 5.540 1.140 ;
        RECT 1.780 0.360 2.040 0.620 ;
        RECT 4.190 0.360 4.450 0.620 ;
  END
END sky130_hilas_drainSelect01

MACRO sky130_hilas_DAC5bit01
  CLASS CORE ;
  FOREIGN sky130_hilas_DAC5bit01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.580 BY 5.970 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    USE ANALOG ;
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER met2 ;
        RECT 8.260 0.990 8.580 1.020 ;
        RECT 0.000 0.790 8.580 0.990 ;
        RECT 8.260 0.760 8.580 0.790 ;
    END
  END A0
  PIN A1
    USE ANALOG ;
    ANTENNAGATEAREA 0.456300 ;
    PORT
      LAYER met2 ;
        RECT 11.590 5.630 11.910 5.950 ;
        RECT 11.710 2.110 11.860 5.630 ;
        RECT 0.000 1.910 11.870 2.110 ;
        RECT 0.000 1.900 0.140 1.910 ;
    END
  END A1
  PIN A2
    USE ANALOG ;
    ANTENNAGATEAREA 0.608400 ;
    PORT
      LAYER met2 ;
        RECT 9.980 5.650 10.300 5.950 ;
        RECT 9.980 5.630 10.310 5.650 ;
        RECT 10.110 3.090 10.310 5.630 ;
        RECT 0.000 2.880 10.310 3.090 ;
    END
  END A2
  PIN A3
    USE ANALOG ;
    ANTENNAGATEAREA 2.281500 ;
    PORT
      LAYER met2 ;
        RECT 8.370 5.620 8.690 5.940 ;
        RECT 3.540 5.420 3.860 5.570 ;
        RECT 3.480 5.250 3.860 5.420 ;
        RECT 0.000 4.960 2.060 5.020 ;
        RECT 3.480 4.960 3.700 5.250 ;
        RECT 8.400 4.970 8.650 5.620 ;
        RECT 8.400 4.960 8.680 4.970 ;
        RECT 0.000 4.810 8.680 4.960 ;
        RECT 0.260 4.630 0.460 4.810 ;
        RECT 1.900 4.660 8.680 4.810 ;
        RECT 0.210 4.310 0.530 4.630 ;
    END
  END A3
  PIN A4
    USE ANALOG ;
    ANTENNAGATEAREA 3.650400 ;
    PORT
      LAYER met2 ;
        RECT 0.000 5.940 7.050 5.970 ;
        RECT 0.000 5.780 7.070 5.940 ;
        RECT 0.000 5.760 0.150 5.780 ;
        RECT 0.350 5.620 0.670 5.780 ;
        RECT 1.940 5.630 2.260 5.780 ;
        RECT 5.140 5.620 5.460 5.780 ;
        RECT 6.750 5.620 7.070 5.780 ;
    END
  END A4
  PIN VPWR
    USE ANALOG ;
    ANTENNADIFFAREA 3.264300 ;
    PORT
      LAYER met2 ;
        RECT 12.710 5.690 13.870 5.970 ;
        RECT 12.830 5.510 13.140 5.690 ;
        RECT 13.460 5.680 13.870 5.690 ;
        RECT 13.500 5.510 13.810 5.680 ;
    END
  END VPWR
  PIN OUT
    USE ANALOG ;
    ANTENNADIFFAREA 3.264300 ;
    PORT
      LAYER met1 ;
        RECT 3.010 0.240 3.240 0.290 ;
        RECT 4.630 0.240 4.860 0.290 ;
        RECT 6.230 0.240 6.460 0.290 ;
        RECT 7.850 0.240 8.080 0.290 ;
        RECT 9.450 0.240 9.680 0.290 ;
        RECT 11.070 0.240 11.300 0.290 ;
        RECT 12.670 0.240 12.900 0.290 ;
        RECT 14.280 0.240 14.510 0.290 ;
        RECT 3.010 0.010 16.580 0.240 ;
        RECT 3.010 0.000 3.240 0.010 ;
        RECT 4.630 0.000 4.860 0.010 ;
        RECT 6.230 0.000 6.460 0.010 ;
        RECT 7.850 0.000 8.080 0.010 ;
        RECT 9.450 0.000 9.680 0.010 ;
        RECT 11.070 0.000 11.300 0.010 ;
        RECT 12.670 0.000 12.900 0.010 ;
        RECT 14.280 0.000 14.510 0.010 ;
    END
  END OUT
  OBS
      LAYER nwell ;
        RECT 0.370 0.030 16.470 5.680 ;
      LAYER li1 ;
        RECT 0.400 5.470 0.610 5.900 ;
        RECT 1.990 5.480 2.200 5.910 ;
        RECT 3.390 5.500 3.820 5.520 ;
        RECT 0.420 5.450 0.590 5.470 ;
        RECT 2.010 5.460 2.180 5.480 ;
        RECT 3.370 5.330 3.820 5.500 ;
        RECT 5.190 5.470 5.400 5.900 ;
        RECT 6.800 5.470 7.010 5.900 ;
        RECT 8.420 5.470 8.630 5.900 ;
        RECT 10.030 5.480 10.240 5.910 ;
        RECT 11.640 5.480 11.850 5.910 ;
        RECT 12.950 5.800 13.160 5.810 ;
        RECT 12.840 5.760 13.160 5.800 ;
        RECT 13.510 5.760 13.830 5.800 ;
        RECT 12.840 5.570 13.170 5.760 ;
        RECT 13.510 5.570 13.840 5.760 ;
        RECT 12.840 5.540 13.160 5.570 ;
        RECT 13.510 5.540 13.830 5.570 ;
        RECT 5.210 5.450 5.380 5.470 ;
        RECT 6.820 5.450 6.990 5.470 ;
        RECT 8.440 5.450 8.610 5.470 ;
        RECT 10.050 5.460 10.220 5.480 ;
        RECT 11.660 5.460 11.830 5.480 ;
        RECT 3.390 5.310 3.820 5.330 ;
        RECT 3.980 5.030 4.150 5.040 ;
        RECT 12.950 5.030 13.160 5.540 ;
        RECT 13.620 5.030 13.790 5.540 ;
        RECT 2.370 4.800 13.800 5.030 ;
        RECT 0.260 4.160 0.470 4.590 ;
        RECT 2.370 4.460 2.540 4.800 ;
        RECT 0.280 4.140 0.450 4.160 ;
        RECT 2.360 4.130 2.540 4.460 ;
        RECT 0.320 3.210 0.530 3.640 ;
        RECT 2.370 3.500 2.540 4.130 ;
        RECT 0.340 3.190 0.510 3.210 ;
        RECT 2.360 3.170 2.540 3.500 ;
        RECT 0.320 2.270 0.530 2.700 ;
        RECT 2.370 2.540 2.540 3.170 ;
        RECT 0.340 2.250 0.510 2.270 ;
        RECT 2.360 2.210 2.540 2.540 ;
        RECT 2.370 1.580 2.540 2.210 ;
        RECT 2.360 1.250 2.540 1.580 ;
        RECT 2.370 1.240 2.540 1.250 ;
        RECT 3.030 4.460 3.200 4.470 ;
        RECT 3.980 4.460 4.150 4.800 ;
        RECT 5.570 4.460 5.740 4.800 ;
        RECT 3.030 4.130 3.210 4.460 ;
        RECT 3.970 4.130 4.150 4.460 ;
        RECT 4.650 4.430 4.820 4.460 ;
        RECT 4.650 4.130 4.830 4.430 ;
        RECT 3.030 3.500 3.200 4.130 ;
        RECT 3.980 3.500 4.150 4.130 ;
        RECT 4.660 3.500 4.830 4.130 ;
        RECT 3.030 3.170 3.210 3.500 ;
        RECT 3.970 3.170 4.150 3.500 ;
        RECT 4.650 3.170 4.830 3.500 ;
        RECT 3.030 2.540 3.200 3.170 ;
        RECT 3.980 2.540 4.150 3.170 ;
        RECT 4.660 2.540 4.830 3.170 ;
        RECT 3.030 2.210 3.210 2.540 ;
        RECT 3.970 2.210 4.150 2.540 ;
        RECT 4.650 2.210 4.830 2.540 ;
        RECT 3.030 1.580 3.200 2.210 ;
        RECT 3.980 1.580 4.150 2.210 ;
        RECT 4.660 1.580 4.830 2.210 ;
        RECT 3.030 1.250 3.210 1.580 ;
        RECT 3.970 1.250 4.150 1.580 ;
        RECT 4.650 1.250 4.830 1.580 ;
        RECT 3.030 0.260 3.200 1.250 ;
        RECT 3.980 1.240 4.150 1.250 ;
        RECT 4.660 0.260 4.830 1.250 ;
        RECT 5.570 4.130 5.750 4.460 ;
        RECT 5.570 3.500 5.740 4.130 ;
        RECT 5.570 3.170 5.750 3.500 ;
        RECT 5.570 2.540 5.740 3.170 ;
        RECT 5.570 2.210 5.750 2.540 ;
        RECT 5.570 1.580 5.740 2.210 ;
        RECT 5.570 1.250 5.750 1.580 ;
        RECT 5.570 1.240 5.740 1.250 ;
        RECT 6.260 0.260 6.430 4.510 ;
        RECT 6.740 3.220 6.950 3.650 ;
        RECT 6.760 3.200 6.930 3.220 ;
        RECT 7.190 1.240 7.360 4.800 ;
        RECT 8.810 4.460 8.980 4.800 ;
        RECT 7.870 4.130 8.050 4.460 ;
        RECT 8.800 4.130 8.980 4.460 ;
        RECT 7.880 3.500 8.050 4.130 ;
        RECT 8.810 3.500 8.980 4.130 ;
        RECT 7.870 3.170 8.050 3.500 ;
        RECT 8.800 3.170 8.980 3.500 ;
        RECT 7.880 2.540 8.050 3.170 ;
        RECT 8.270 2.740 8.440 2.760 ;
        RECT 7.870 2.210 8.050 2.540 ;
        RECT 8.250 2.310 8.460 2.740 ;
        RECT 7.880 1.580 8.050 2.210 ;
        RECT 8.810 1.580 8.980 3.170 ;
        RECT 7.870 1.250 8.050 1.580 ;
        RECT 8.800 1.260 8.980 1.580 ;
        RECT 8.800 1.250 8.970 1.260 ;
        RECT 7.880 0.260 8.050 1.250 ;
        RECT 9.480 0.260 9.650 4.510 ;
        RECT 9.990 1.310 10.200 1.740 ;
        RECT 10.010 1.290 10.180 1.310 ;
        RECT 10.410 1.250 10.580 4.800 ;
        RECT 11.100 4.460 11.270 4.510 ;
        RECT 11.090 4.130 11.270 4.460 ;
        RECT 11.100 3.500 11.270 4.130 ;
        RECT 11.090 3.170 11.270 3.500 ;
        RECT 11.100 2.540 11.270 3.170 ;
        RECT 11.090 2.210 11.270 2.540 ;
        RECT 11.100 1.580 11.270 2.210 ;
        RECT 11.090 1.250 11.270 1.580 ;
        RECT 12.020 1.250 12.190 4.800 ;
        RECT 11.100 0.260 11.270 1.250 ;
        RECT 12.700 0.260 12.870 4.490 ;
        RECT 13.630 1.230 13.800 4.800 ;
        RECT 14.310 0.260 14.480 4.670 ;
        RECT 3.030 0.030 3.220 0.260 ;
        RECT 4.650 0.030 4.840 0.260 ;
        RECT 6.250 0.030 6.440 0.260 ;
        RECT 7.870 0.030 8.060 0.260 ;
        RECT 9.470 0.030 9.660 0.260 ;
        RECT 11.090 0.030 11.280 0.260 ;
        RECT 12.690 0.030 12.880 0.260 ;
        RECT 14.300 0.030 14.490 0.260 ;
        RECT 3.030 0.010 3.200 0.030 ;
        RECT 4.660 0.010 4.830 0.030 ;
        RECT 6.260 0.010 6.430 0.030 ;
        RECT 7.880 0.010 8.050 0.030 ;
        RECT 9.480 0.010 9.650 0.030 ;
        RECT 11.100 0.010 11.270 0.030 ;
        RECT 12.700 0.010 12.870 0.030 ;
        RECT 14.310 0.010 14.480 0.030 ;
      LAYER mcon ;
        RECT 12.900 5.580 13.070 5.750 ;
        RECT 13.570 5.580 13.740 5.750 ;
        RECT 8.270 2.590 8.440 2.760 ;
        RECT 3.040 0.060 3.210 0.230 ;
        RECT 4.660 0.060 4.830 0.230 ;
        RECT 6.260 0.060 6.430 0.230 ;
        RECT 7.880 0.060 8.050 0.230 ;
        RECT 9.480 0.060 9.650 0.230 ;
        RECT 11.100 0.060 11.270 0.230 ;
        RECT 12.700 0.060 12.870 0.230 ;
        RECT 14.310 0.060 14.480 0.230 ;
      LAYER met1 ;
        RECT 0.350 5.620 0.670 5.940 ;
        RECT 1.940 5.630 2.260 5.950 ;
        RECT 0.390 5.390 0.620 5.620 ;
        RECT 1.980 5.400 2.210 5.630 ;
        RECT 5.140 5.620 5.460 5.940 ;
        RECT 6.750 5.620 7.070 5.940 ;
        RECT 8.370 5.620 8.690 5.940 ;
        RECT 9.980 5.630 10.300 5.950 ;
        RECT 11.590 5.630 11.910 5.950 ;
        RECT 3.540 5.530 3.860 5.570 ;
        RECT 3.310 5.300 3.860 5.530 ;
        RECT 5.180 5.390 5.410 5.620 ;
        RECT 6.790 5.390 7.020 5.620 ;
        RECT 8.410 5.390 8.640 5.620 ;
        RECT 10.020 5.400 10.250 5.630 ;
        RECT 11.630 5.400 11.860 5.630 ;
        RECT 12.830 5.510 13.150 5.830 ;
        RECT 13.500 5.510 13.820 5.830 ;
        RECT 3.540 5.250 3.860 5.300 ;
        RECT 0.210 4.310 0.530 4.630 ;
        RECT 0.250 4.080 0.480 4.310 ;
        RECT 0.270 3.360 0.590 3.680 ;
        RECT 6.740 3.560 10.190 3.730 ;
        RECT 6.740 3.430 6.960 3.560 ;
        RECT 0.310 3.130 0.540 3.360 ;
        RECT 6.730 3.140 6.960 3.430 ;
        RECT 0.270 2.420 0.590 2.740 ;
        RECT 8.240 2.530 8.470 2.820 ;
        RECT 0.310 2.190 0.540 2.420 ;
        RECT 8.250 2.310 8.470 2.530 ;
        RECT 8.290 1.050 8.470 2.310 ;
        RECT 9.990 1.740 10.190 3.560 ;
        RECT 9.990 1.520 10.210 1.740 ;
        RECT 9.980 1.230 10.210 1.520 ;
        RECT 8.290 0.730 8.550 1.050 ;
      LAYER via ;
        RECT 0.380 5.650 0.640 5.910 ;
        RECT 1.970 5.660 2.230 5.920 ;
        RECT 5.170 5.650 5.430 5.910 ;
        RECT 6.780 5.650 7.040 5.910 ;
        RECT 8.400 5.650 8.660 5.910 ;
        RECT 10.010 5.660 10.270 5.920 ;
        RECT 11.620 5.660 11.880 5.920 ;
        RECT 3.570 5.280 3.830 5.540 ;
        RECT 12.860 5.540 13.120 5.800 ;
        RECT 13.530 5.540 13.790 5.800 ;
        RECT 0.240 4.340 0.500 4.600 ;
        RECT 0.300 3.390 0.560 3.650 ;
        RECT 0.300 2.450 0.560 2.710 ;
        RECT 8.290 0.760 8.550 1.020 ;
      LAYER met2 ;
        RECT 0.270 3.360 0.590 3.680 ;
        RECT 0.270 2.420 0.590 2.740 ;
  END
END sky130_hilas_DAC5bit01

MACRO sky130_hilas_capacitorSize04
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize04 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.780 BY 5.290 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAP1TERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 4.960 3.830 5.620 4.490 ;
    END
  END CAP1TERM02
  PIN CAP2TERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 4.960 0.830 5.620 1.490 ;
    END
  END CAP2TERM02
  PIN CAP2TERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 0.120 1.230 0.780 1.490 ;
        RECT 2.560 1.230 3.010 1.240 ;
        RECT 0.120 0.830 3.060 1.230 ;
        RECT 0.570 0.820 3.060 0.830 ;
        RECT 2.540 0.740 3.060 0.820 ;
    END
  END CAP2TERM01
  PIN CAP1TERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 0.090 4.240 0.750 4.490 ;
        RECT 2.560 4.240 3.010 4.250 ;
        RECT 0.090 3.830 3.060 4.240 ;
        RECT 2.540 3.750 3.060 3.830 ;
    END
  END CAP1TERM01
  OBS
      LAYER met2 ;
        RECT 0.020 4.980 5.770 5.160 ;
        RECT 0.020 4.550 5.770 4.730 ;
        RECT 0.220 4.310 0.590 4.370 ;
        RECT 0.020 4.030 0.590 4.310 ;
        RECT 0.220 3.970 0.590 4.030 ;
        RECT 5.090 4.310 5.460 4.370 ;
        RECT 5.090 4.030 5.770 4.310 ;
        RECT 5.090 3.970 5.460 4.030 ;
        RECT 0.020 3.550 5.770 3.730 ;
        RECT 0.020 3.120 5.770 3.300 ;
        RECT 0.020 1.970 5.770 2.140 ;
        RECT 0.020 1.550 5.770 1.720 ;
        RECT 0.250 1.310 0.620 1.370 ;
        RECT 0.020 1.030 0.620 1.310 ;
        RECT 0.250 0.970 0.620 1.030 ;
        RECT 5.090 1.310 5.460 1.370 ;
        RECT 5.090 1.030 5.780 1.310 ;
        RECT 5.090 0.970 5.460 1.030 ;
        RECT 0.020 0.570 5.770 0.740 ;
        RECT 0.020 0.130 5.770 0.300 ;
      LAYER via2 ;
        RECT 0.270 4.030 0.550 4.310 ;
        RECT 5.140 4.030 5.420 4.310 ;
        RECT 0.300 1.030 0.580 1.310 ;
        RECT 5.140 1.030 5.420 1.310 ;
      LAYER met3 ;
        RECT 1.710 4.520 4.010 5.290 ;
        RECT 0.000 3.770 0.790 4.520 ;
        RECT 1.710 3.770 5.660 4.520 ;
        RECT 1.710 3.010 4.010 3.770 ;
        RECT 0.030 0.770 0.820 1.520 ;
        RECT 1.710 1.510 4.010 2.280 ;
        RECT 4.870 1.510 5.660 1.520 ;
        RECT 1.710 0.780 5.660 1.510 ;
        RECT 1.710 0.000 4.010 0.780 ;
        RECT 4.870 0.770 5.660 0.780 ;
      LAYER via3 ;
        RECT 0.190 3.920 0.620 4.400 ;
        RECT 5.060 3.920 5.490 4.400 ;
        RECT 0.220 0.920 0.650 1.400 ;
        RECT 5.060 0.920 5.490 1.400 ;
  END
END sky130_hilas_capacitorSize04

MACRO sky130_hilas_capacitorArray01
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorArray01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.700 BY 9.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM2
    USE ANALOG ;
    PORT
      LAYER met3 ;
        RECT 35.230 2.200 36.380 3.840 ;
        RECT 35.680 2.190 36.380 2.200 ;
    END
  END CAPTERM2
  PIN CAPTERM1
    USE ANALOG ;
    ANTENNADIFFAREA 0.087000 ;
    PORT
      LAYER met3 ;
        RECT 11.250 5.740 11.630 6.030 ;
        RECT 11.170 4.490 11.710 5.740 ;
    END
  END CAPTERM1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 5.400 5.380 5.720 5.390 ;
        RECT 8.980 5.380 36.700 5.550 ;
        RECT 5.400 5.370 36.700 5.380 ;
        RECT 5.400 5.200 9.650 5.370 ;
        RECT 5.400 5.130 5.720 5.200 ;
        RECT 9.330 5.140 9.650 5.200 ;
    END
  END VINJ
  PIN GATESELECT
    PORT
      LAYER met1 ;
        RECT 9.120 6.000 9.310 6.050 ;
    END
  END GATESELECT
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 0.360 5.910 0.760 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.360 0.000 0.750 0.120 ;
    END
  END VTUN
  PIN GATE
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 4.420 5.970 4.790 6.050 ;
        RECT 4.410 5.920 4.790 5.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.400 0.130 4.410 0.150 ;
        RECT 4.400 0.010 4.790 0.130 ;
        RECT 4.400 0.000 4.410 0.010 ;
    END
  END GATE
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 0.000 3.510 0.120 3.690 ;
    END
    PORT
      LAYER met2 ;
        RECT 35.690 3.690 36.700 3.700 ;
        RECT 8.940 3.510 36.700 3.690 ;
    END
  END DRAIN2
  PIN DRAIN1
    PORT
      LAYER met2 ;
        RECT 0.010 5.370 0.120 5.550 ;
    END
  END DRAIN1
  PIN DRAIN4
    PORT
      LAYER met2 ;
        RECT 8.810 0.520 36.700 0.690 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.020 0.520 0.120 0.690 ;
    END
  END DRAIN4
  PIN DRAIN3
    PORT
      LAYER met2 ;
        RECT 8.770 2.360 36.700 2.530 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.020 2.360 0.120 2.530 ;
    END
  END DRAIN3
  PIN VGND
    ANTENNADIFFAREA 1.978000 ;
    PORT
      LAYER nwell ;
        RECT 2.650 8.010 4.380 9.870 ;
        RECT 2.640 6.170 4.380 8.010 ;
        RECT 2.650 3.820 4.380 6.170 ;
      LAYER met1 ;
        RECT 3.000 6.050 3.400 9.870 ;
        RECT 2.800 5.990 3.400 6.050 ;
        RECT 3.000 3.820 3.400 5.990 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.730 5.980 6.970 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.800 0.000 3.040 0.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.730 0.000 6.970 0.070 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 0.010 5.370 0.120 5.550 ;
        RECT 6.400 3.820 8.630 9.870 ;
        RECT 10.160 9.860 12.710 9.870 ;
        RECT 10.160 6.050 12.720 9.860 ;
        RECT 10.070 6.040 35.420 6.050 ;
        RECT 10.080 5.970 35.420 6.040 ;
        RECT 0.000 3.510 0.120 3.690 ;
        RECT 0.020 0.520 0.120 0.690 ;
        RECT 10.060 0.060 35.420 5.970 ;
        RECT 10.070 0.010 35.420 0.060 ;
        RECT 12.000 0.000 35.420 0.010 ;
      LAYER li1 ;
        RECT 10.260 9.460 10.580 9.470 ;
        RECT 10.260 9.290 10.840 9.460 ;
        RECT 10.260 9.240 10.590 9.290 ;
        RECT 10.260 9.210 10.580 9.240 ;
        RECT 12.120 9.190 12.320 9.540 ;
        RECT 10.260 8.880 10.580 8.920 ;
        RECT 10.260 8.840 10.590 8.880 ;
        RECT 10.260 8.670 10.840 8.840 ;
        RECT 10.260 8.660 10.580 8.670 ;
        RECT 5.470 8.120 5.640 8.630 ;
        RECT 9.410 8.110 9.580 8.620 ;
        RECT 11.390 8.600 11.590 9.170 ;
        RECT 12.120 9.160 12.330 9.190 ;
        RECT 12.110 8.570 12.330 9.160 ;
        RECT 10.260 8.030 10.580 8.040 ;
        RECT 10.260 7.860 10.840 8.030 ;
        RECT 10.260 7.820 10.590 7.860 ;
        RECT 10.260 7.780 10.580 7.820 ;
        RECT 11.390 7.530 11.590 8.100 ;
        RECT 12.110 7.540 12.330 8.130 ;
        RECT 12.120 7.510 12.330 7.540 ;
        RECT 10.260 7.460 10.580 7.490 ;
        RECT 3.070 6.620 3.620 7.050 ;
        RECT 5.480 6.410 5.650 7.420 ;
        RECT 10.260 7.410 10.590 7.460 ;
        RECT 7.100 6.550 7.650 6.980 ;
        RECT 9.410 6.270 9.580 7.280 ;
        RECT 10.260 7.240 10.840 7.410 ;
        RECT 10.260 7.230 10.580 7.240 ;
        RECT 12.120 7.160 12.320 7.510 ;
        RECT 11.510 6.760 11.950 6.930 ;
        RECT 10.260 6.450 10.580 6.460 ;
        RECT 10.260 6.280 10.840 6.450 ;
        RECT 10.260 6.230 10.590 6.280 ;
        RECT 10.260 6.200 10.580 6.230 ;
        RECT 12.120 6.180 12.320 6.530 ;
        RECT 10.260 5.870 10.580 5.910 ;
        RECT 10.260 5.830 10.590 5.870 ;
        RECT 10.260 5.660 10.840 5.830 ;
        RECT 10.260 5.650 10.580 5.660 ;
        RECT 11.390 5.590 11.590 6.160 ;
        RECT 12.120 6.150 12.330 6.180 ;
        RECT 12.110 5.560 12.330 6.150 ;
        RECT 10.260 5.030 10.580 5.040 ;
        RECT 10.260 4.860 10.840 5.030 ;
        RECT 10.260 4.820 10.590 4.860 ;
        RECT 10.260 4.780 10.580 4.820 ;
        RECT 11.390 4.530 11.590 5.100 ;
        RECT 12.110 4.540 12.330 5.130 ;
        RECT 12.120 4.510 12.330 4.540 ;
        RECT 10.260 4.460 10.580 4.490 ;
        RECT 10.260 4.410 10.590 4.460 ;
        RECT 10.260 4.240 10.840 4.410 ;
        RECT 10.260 4.230 10.580 4.240 ;
        RECT 12.120 4.160 12.320 4.510 ;
      LAYER mcon ;
        RECT 10.320 9.250 10.490 9.420 ;
        RECT 11.400 8.960 11.570 9.130 ;
        RECT 10.320 8.700 10.490 8.870 ;
        RECT 5.470 8.460 5.640 8.630 ;
        RECT 9.410 8.450 9.580 8.620 ;
        RECT 12.130 8.990 12.300 9.160 ;
        RECT 10.320 7.830 10.490 8.000 ;
        RECT 11.400 7.570 11.570 7.740 ;
        RECT 12.130 7.540 12.300 7.710 ;
        RECT 10.320 7.280 10.490 7.450 ;
        RECT 3.070 6.700 3.340 6.970 ;
        RECT 5.480 7.000 5.650 7.170 ;
        RECT 5.480 6.660 5.650 6.830 ;
        RECT 7.100 6.630 7.370 6.900 ;
        RECT 9.410 6.860 9.580 7.030 ;
        RECT 11.770 6.760 11.950 6.930 ;
        RECT 9.410 6.520 9.580 6.690 ;
        RECT 10.320 6.240 10.490 6.410 ;
        RECT 11.400 5.950 11.570 6.120 ;
        RECT 10.320 5.690 10.490 5.860 ;
        RECT 12.130 5.980 12.300 6.150 ;
        RECT 10.320 4.830 10.490 5.000 ;
        RECT 11.400 4.570 11.570 4.740 ;
        RECT 12.130 4.540 12.300 4.710 ;
        RECT 10.320 4.280 10.490 4.450 ;
      LAYER met1 ;
        RECT 5.440 8.690 5.680 9.870 ;
        RECT 5.430 8.030 5.690 8.690 ;
        RECT 5.440 5.420 5.680 8.030 ;
        RECT 7.050 7.950 7.430 9.870 ;
        RECT 9.370 8.710 9.610 9.870 ;
        RECT 10.250 9.180 10.570 9.500 ;
        RECT 11.390 9.190 11.550 9.870 ;
        RECT 11.390 9.170 11.590 9.190 ;
        RECT 9.350 8.050 9.620 8.710 ;
        RECT 10.250 8.630 10.570 8.950 ;
        RECT 11.370 8.930 11.600 9.170 ;
        RECT 11.390 8.710 11.590 8.930 ;
        RECT 11.760 8.880 11.950 9.870 ;
        RECT 12.200 9.220 12.360 9.870 ;
        RECT 11.780 8.760 11.950 8.880 ;
        RECT 7.040 6.090 7.430 7.950 ;
        RECT 5.430 5.100 5.690 5.420 ;
        RECT 5.440 3.820 5.680 5.100 ;
        RECT 7.050 3.820 7.430 6.090 ;
        RECT 9.370 6.050 9.610 8.050 ;
        RECT 10.250 7.750 10.570 8.070 ;
        RECT 11.390 7.990 11.550 8.710 ;
        RECT 11.390 7.770 11.590 7.990 ;
        RECT 11.790 7.940 11.950 8.760 ;
        RECT 12.090 8.670 12.360 9.220 ;
        RECT 12.090 8.620 12.370 8.670 ;
        RECT 12.200 8.530 12.370 8.620 ;
        RECT 12.200 8.170 12.360 8.530 ;
        RECT 12.200 8.080 12.370 8.170 ;
        RECT 11.780 7.820 11.950 7.940 ;
        RECT 11.370 7.530 11.600 7.770 ;
        RECT 10.250 7.200 10.570 7.520 ;
        RECT 11.390 7.510 11.590 7.530 ;
        RECT 10.250 6.170 10.570 6.490 ;
        RECT 11.390 6.180 11.550 7.510 ;
        RECT 11.760 6.960 11.950 7.820 ;
        RECT 12.090 8.030 12.370 8.080 ;
        RECT 12.090 7.480 12.360 8.030 ;
        RECT 11.740 6.730 11.980 6.960 ;
        RECT 11.390 6.160 11.590 6.180 ;
        RECT 8.700 5.710 8.960 6.030 ;
        RECT 9.370 6.000 9.720 6.050 ;
        RECT 9.370 5.460 9.610 6.000 ;
        RECT 10.250 5.620 10.570 5.940 ;
        RECT 11.370 5.920 11.600 6.160 ;
        RECT 11.390 5.700 11.590 5.920 ;
        RECT 11.760 5.870 11.950 6.730 ;
        RECT 12.200 6.210 12.360 7.480 ;
        RECT 11.780 5.750 11.950 5.870 ;
        RECT 9.360 5.140 9.620 5.460 ;
        RECT 9.370 3.820 9.610 5.140 ;
        RECT 10.250 4.750 10.570 5.070 ;
        RECT 11.390 4.990 11.550 5.700 ;
        RECT 11.390 4.770 11.590 4.990 ;
        RECT 11.790 4.940 11.950 5.750 ;
        RECT 12.090 5.660 12.360 6.210 ;
        RECT 12.090 5.610 12.370 5.660 ;
        RECT 12.200 5.520 12.370 5.610 ;
        RECT 12.200 5.170 12.360 5.520 ;
        RECT 12.200 5.080 12.370 5.170 ;
        RECT 11.780 4.820 11.950 4.940 ;
        RECT 11.370 4.530 11.600 4.770 ;
        RECT 10.250 4.200 10.570 4.520 ;
        RECT 11.390 4.510 11.590 4.530 ;
        RECT 11.390 3.830 11.550 4.510 ;
        RECT 11.760 3.830 11.950 4.820 ;
        RECT 12.090 5.030 12.370 5.080 ;
        RECT 12.090 4.480 12.360 5.030 ;
        RECT 12.200 3.830 12.360 4.480 ;
        RECT 8.750 0.010 8.910 0.070 ;
        RECT 9.120 0.010 9.310 0.070 ;
        RECT 9.560 0.010 9.720 0.070 ;
      LAYER via ;
        RECT 10.280 9.210 10.540 9.470 ;
        RECT 10.280 8.660 10.540 8.920 ;
        RECT 5.430 5.130 5.690 5.390 ;
        RECT 10.280 7.780 10.540 8.040 ;
        RECT 10.280 7.230 10.540 7.490 ;
        RECT 10.280 6.200 10.540 6.460 ;
        RECT 8.700 5.740 8.960 6.000 ;
        RECT 10.280 5.650 10.540 5.910 ;
        RECT 9.360 5.170 9.620 5.430 ;
        RECT 10.280 4.780 10.540 5.040 ;
        RECT 10.280 4.230 10.540 4.490 ;
      LAYER met2 ;
        RECT 10.250 9.370 10.560 9.510 ;
        RECT 2.650 9.190 12.720 9.370 ;
        RECT 10.250 9.180 10.560 9.190 ;
        RECT 10.250 8.940 10.560 8.960 ;
        RECT 2.650 8.760 12.720 8.940 ;
        RECT 10.250 8.630 10.560 8.760 ;
        RECT 10.250 7.940 10.560 8.070 ;
        RECT 2.640 7.760 12.720 7.940 ;
        RECT 10.250 7.740 10.560 7.760 ;
        RECT 10.250 7.510 10.560 7.520 ;
        RECT 2.640 7.330 12.720 7.510 ;
        RECT 10.250 7.190 10.560 7.330 ;
        RECT 10.250 6.360 10.560 6.500 ;
        RECT 10.250 6.350 12.720 6.360 ;
        RECT 2.660 6.180 12.720 6.350 ;
        RECT 10.250 6.170 10.560 6.180 ;
        RECT 10.740 6.020 11.250 6.050 ;
        RECT 8.670 5.930 8.990 6.000 ;
        RECT 10.250 5.930 10.560 5.950 ;
        RECT 10.740 5.930 11.670 6.020 ;
        RECT 2.660 5.760 12.720 5.930 ;
        RECT 8.670 5.750 12.720 5.760 ;
        RECT 8.670 5.740 11.670 5.750 ;
        RECT 10.250 5.620 10.560 5.740 ;
        RECT 11.170 5.720 11.670 5.740 ;
        RECT 8.920 4.950 36.700 5.120 ;
        RECT 2.660 4.940 36.700 4.950 ;
        RECT 2.660 4.780 12.720 4.940 ;
        RECT 3.440 4.690 4.980 4.780 ;
        RECT 10.160 4.760 12.720 4.780 ;
        RECT 10.250 4.740 10.560 4.760 ;
        RECT 10.250 4.510 10.560 4.520 ;
        RECT 2.660 4.340 12.720 4.510 ;
        RECT 10.250 4.330 12.720 4.340 ;
        RECT 10.250 4.290 10.560 4.330 ;
        RECT 9.880 4.190 10.560 4.290 ;
        RECT 9.880 4.120 10.250 4.190 ;
        RECT 8.980 3.940 36.700 4.120 ;
        RECT 9.880 3.890 10.250 3.940 ;
        RECT 36.010 2.790 36.700 3.200 ;
        RECT 9.840 2.110 10.210 2.200 ;
        RECT 8.870 1.940 36.700 2.110 ;
        RECT 9.840 1.800 10.210 1.940 ;
        RECT 10.930 1.130 11.300 1.330 ;
        RECT 8.850 0.960 36.700 1.130 ;
        RECT 10.930 0.930 11.300 0.960 ;
      LAYER via2 ;
        RECT 11.300 5.720 11.580 6.000 ;
        RECT 9.930 3.950 10.210 4.230 ;
        RECT 36.080 2.850 36.370 3.130 ;
        RECT 9.890 1.860 10.170 2.140 ;
        RECT 10.980 0.990 11.260 1.270 ;
      LAYER met3 ;
        RECT 9.660 3.690 10.450 4.440 ;
        RECT 9.620 2.300 10.410 2.350 ;
        RECT 9.620 2.000 10.550 2.300 ;
        RECT 9.620 1.600 10.410 2.000 ;
        RECT 10.710 1.090 11.500 1.480 ;
        RECT 10.710 0.790 11.640 1.090 ;
        RECT 10.710 0.730 11.500 0.790 ;
      LAYER via3 ;
        RECT 9.850 3.840 10.280 4.320 ;
        RECT 9.810 1.750 10.240 2.230 ;
        RECT 10.900 0.880 11.330 1.360 ;
      LAYER met4 ;
        RECT 12.790 5.380 16.890 5.680 ;
        RECT 11.100 4.770 13.800 4.880 ;
        RECT 11.100 4.470 14.010 4.770 ;
        RECT 9.750 4.050 10.410 4.410 ;
        RECT 13.500 4.130 14.010 4.470 ;
        RECT 16.510 4.180 16.890 5.380 ;
        RECT 19.350 4.210 22.630 4.510 ;
        RECT 9.750 3.750 11.770 4.050 ;
        RECT 11.470 3.190 11.770 3.750 ;
        RECT 19.350 3.190 19.650 4.210 ;
        RECT 22.330 3.190 22.630 4.210 ;
        RECT 11.470 2.890 22.630 3.190 ;
        RECT 25.030 4.190 33.920 4.490 ;
        RECT 9.710 2.300 10.370 2.320 ;
        RECT 13.710 2.300 16.900 2.330 ;
        RECT 19.350 2.300 19.650 2.330 ;
        RECT 9.710 2.000 22.570 2.300 ;
        RECT 9.710 1.660 10.370 2.000 ;
        RECT 13.710 1.630 14.010 2.000 ;
        RECT 16.600 1.660 16.900 2.000 ;
        RECT 19.350 1.660 19.650 2.000 ;
        RECT 16.600 1.630 19.650 1.660 ;
        RECT 22.270 1.630 22.570 2.000 ;
        RECT 10.800 1.090 11.460 1.450 ;
        RECT 13.710 1.330 22.570 1.630 ;
        RECT 25.030 1.670 25.330 4.190 ;
        RECT 27.860 4.160 30.970 4.190 ;
        RECT 27.860 1.670 28.160 4.160 ;
        RECT 30.670 1.670 30.970 4.160 ;
        RECT 33.620 1.670 33.920 4.190 ;
        RECT 25.030 1.370 33.980 1.670 ;
        RECT 30.670 1.360 33.980 1.370 ;
        RECT 10.800 0.790 11.850 1.090 ;
        RECT 11.550 0.550 11.850 0.790 ;
        RECT 33.680 0.550 33.980 1.360 ;
        RECT 11.550 0.250 33.980 0.550 ;
  END
END sky130_hilas_capacitorArray01

MACRO sky130_hilas_pFETmed
  CLASS CORE ;
  FOREIGN sky130_hilas_pFETmed ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.190 BY 2.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 0.000 0.000 1.190 2.870 ;
      LAYER li1 ;
        RECT 0.240 0.150 0.410 2.640 ;
        RECT 0.790 0.140 0.960 2.640 ;
  END
END sky130_hilas_pFETmed

MACRO sky130_hilas_swc4x1cellOverlap2
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x1cellOverlap2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.350 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 2.790 6.040 9.340 6.050 ;
        RECT 2.790 0.020 9.350 6.040 ;
        RECT 2.790 0.010 9.340 0.020 ;
        RECT 2.790 0.000 6.790 0.010 ;
      LAYER li1 ;
        RECT 1.060 4.840 1.230 5.730 ;
        RECT 3.140 4.740 6.450 5.720 ;
        RECT 6.890 5.640 7.210 5.650 ;
        RECT 6.890 5.470 7.470 5.640 ;
        RECT 6.890 5.420 7.220 5.470 ;
        RECT 6.890 5.390 7.210 5.420 ;
        RECT 8.750 5.370 8.950 5.720 ;
        RECT 6.890 5.060 7.210 5.100 ;
        RECT 6.890 5.020 7.220 5.060 ;
        RECT 6.890 4.850 7.470 5.020 ;
        RECT 6.890 4.840 7.210 4.850 ;
        RECT 8.020 4.780 8.220 5.350 ;
        RECT 8.750 5.340 8.960 5.370 ;
        RECT 8.740 4.750 8.960 5.340 ;
        RECT 1.060 3.320 1.230 4.210 ;
        RECT 3.140 3.270 6.450 4.250 ;
        RECT 6.890 4.210 7.210 4.220 ;
        RECT 6.890 4.040 7.470 4.210 ;
        RECT 6.890 4.000 7.220 4.040 ;
        RECT 6.890 3.960 7.210 4.000 ;
        RECT 8.020 3.710 8.220 4.280 ;
        RECT 8.740 3.720 8.960 4.310 ;
        RECT 8.750 3.690 8.960 3.720 ;
        RECT 6.890 3.640 7.210 3.670 ;
        RECT 6.890 3.590 7.220 3.640 ;
        RECT 6.890 3.420 7.470 3.590 ;
        RECT 6.890 3.410 7.210 3.420 ;
        RECT 8.750 3.340 8.950 3.690 ;
        RECT 8.140 2.940 8.580 3.110 ;
        RECT 1.060 1.870 1.230 2.760 ;
        RECT 3.140 1.800 6.450 2.780 ;
        RECT 6.890 2.630 7.210 2.640 ;
        RECT 6.890 2.460 7.470 2.630 ;
        RECT 6.890 2.410 7.220 2.460 ;
        RECT 6.890 2.380 7.210 2.410 ;
        RECT 8.750 2.360 8.950 2.710 ;
        RECT 6.890 2.050 7.210 2.090 ;
        RECT 6.890 2.010 7.220 2.050 ;
        RECT 6.890 1.840 7.470 2.010 ;
        RECT 6.890 1.830 7.210 1.840 ;
        RECT 8.020 1.770 8.220 2.340 ;
        RECT 8.750 2.330 8.960 2.360 ;
        RECT 8.740 1.740 8.960 2.330 ;
        RECT 1.060 0.330 1.230 1.220 ;
        RECT 3.140 0.330 6.450 1.310 ;
        RECT 6.890 1.210 7.210 1.220 ;
        RECT 6.890 1.040 7.470 1.210 ;
        RECT 6.890 1.000 7.220 1.040 ;
        RECT 6.890 0.960 7.210 1.000 ;
        RECT 8.020 0.710 8.220 1.280 ;
        RECT 8.740 0.720 8.960 1.310 ;
        RECT 8.750 0.690 8.960 0.720 ;
        RECT 6.890 0.640 7.210 0.670 ;
        RECT 6.890 0.590 7.220 0.640 ;
        RECT 6.890 0.420 7.470 0.590 ;
        RECT 6.890 0.410 7.210 0.420 ;
        RECT 8.750 0.340 8.950 0.690 ;
      LAYER mcon ;
        RECT 1.060 5.530 1.230 5.700 ;
        RECT 4.710 5.490 4.880 5.660 ;
        RECT 6.950 5.430 7.120 5.600 ;
        RECT 4.710 5.140 4.880 5.310 ;
        RECT 8.030 5.140 8.200 5.310 ;
        RECT 4.710 4.800 4.880 4.970 ;
        RECT 6.950 4.880 7.120 5.050 ;
        RECT 8.760 5.170 8.930 5.340 ;
        RECT 1.060 4.010 1.230 4.180 ;
        RECT 4.710 4.020 4.880 4.190 ;
        RECT 6.950 4.010 7.120 4.180 ;
        RECT 4.710 3.670 4.880 3.840 ;
        RECT 8.030 3.750 8.200 3.920 ;
        RECT 8.760 3.720 8.930 3.890 ;
        RECT 4.710 3.330 4.880 3.500 ;
        RECT 6.950 3.460 7.120 3.630 ;
        RECT 8.400 2.940 8.580 3.110 ;
        RECT 1.060 2.560 1.230 2.730 ;
        RECT 4.710 2.550 4.880 2.720 ;
        RECT 6.950 2.420 7.120 2.590 ;
        RECT 4.710 2.200 4.880 2.370 ;
        RECT 8.030 2.130 8.200 2.300 ;
        RECT 4.710 1.860 4.880 2.030 ;
        RECT 6.950 1.870 7.120 2.040 ;
        RECT 8.760 2.160 8.930 2.330 ;
        RECT 1.060 1.020 1.230 1.190 ;
        RECT 4.710 1.080 4.880 1.250 ;
        RECT 6.950 1.010 7.120 1.180 ;
        RECT 4.710 0.730 4.880 0.900 ;
        RECT 8.030 0.750 8.200 0.920 ;
        RECT 8.760 0.720 8.930 0.890 ;
        RECT 4.710 0.390 4.880 0.560 ;
        RECT 6.950 0.460 7.120 0.630 ;
      LAYER met1 ;
        RECT 1.010 0.000 1.280 6.050 ;
        RECT 4.670 5.080 4.910 5.720 ;
        RECT 6.880 5.360 7.200 5.680 ;
        RECT 8.020 5.370 8.180 6.050 ;
        RECT 8.020 5.350 8.220 5.370 ;
        RECT 4.680 4.820 4.910 5.080 ;
        RECT 4.680 4.600 4.920 4.820 ;
        RECT 6.880 4.810 7.200 5.130 ;
        RECT 8.000 5.110 8.230 5.350 ;
        RECT 8.020 4.890 8.220 5.110 ;
        RECT 8.390 5.060 8.580 6.050 ;
        RECT 8.830 5.400 8.990 6.050 ;
        RECT 8.410 4.940 8.580 5.060 ;
        RECT 4.670 3.610 4.910 4.250 ;
        RECT 6.880 3.930 7.200 4.250 ;
        RECT 8.020 4.170 8.180 4.890 ;
        RECT 8.020 3.950 8.220 4.170 ;
        RECT 8.420 4.120 8.580 4.940 ;
        RECT 8.720 4.850 8.990 5.400 ;
        RECT 8.720 4.800 9.000 4.850 ;
        RECT 8.830 4.710 9.000 4.800 ;
        RECT 8.830 4.350 8.990 4.710 ;
        RECT 8.830 4.260 9.000 4.350 ;
        RECT 8.410 4.000 8.580 4.120 ;
        RECT 8.000 3.710 8.230 3.950 ;
        RECT 4.680 3.350 4.910 3.610 ;
        RECT 6.880 3.380 7.200 3.700 ;
        RECT 8.020 3.690 8.220 3.710 ;
        RECT 4.680 3.130 4.920 3.350 ;
        RECT 4.670 2.140 4.910 2.780 ;
        RECT 6.880 2.350 7.200 2.670 ;
        RECT 8.020 2.360 8.180 3.690 ;
        RECT 8.390 3.140 8.580 4.000 ;
        RECT 8.720 4.210 9.000 4.260 ;
        RECT 8.720 3.660 8.990 4.210 ;
        RECT 8.370 2.910 8.610 3.140 ;
        RECT 8.020 2.340 8.220 2.360 ;
        RECT 4.680 1.880 4.910 2.140 ;
        RECT 4.680 1.660 4.920 1.880 ;
        RECT 6.880 1.800 7.200 2.120 ;
        RECT 8.000 2.100 8.230 2.340 ;
        RECT 8.020 1.880 8.220 2.100 ;
        RECT 8.390 2.050 8.580 2.910 ;
        RECT 8.830 2.390 8.990 3.660 ;
        RECT 8.410 1.930 8.580 2.050 ;
        RECT 4.670 0.670 4.910 1.310 ;
        RECT 6.880 0.930 7.200 1.250 ;
        RECT 8.020 1.170 8.180 1.880 ;
        RECT 8.020 0.950 8.220 1.170 ;
        RECT 8.420 1.120 8.580 1.930 ;
        RECT 8.720 1.840 8.990 2.390 ;
        RECT 8.720 1.790 9.000 1.840 ;
        RECT 8.830 1.700 9.000 1.790 ;
        RECT 8.830 1.350 8.990 1.700 ;
        RECT 8.830 1.260 9.000 1.350 ;
        RECT 8.410 1.000 8.580 1.120 ;
        RECT 8.000 0.710 8.230 0.950 ;
        RECT 4.680 0.410 4.910 0.670 ;
        RECT 4.680 0.190 4.920 0.410 ;
        RECT 6.880 0.380 7.200 0.700 ;
        RECT 8.020 0.690 8.220 0.710 ;
        RECT 8.020 0.010 8.180 0.690 ;
        RECT 8.390 0.010 8.580 1.000 ;
        RECT 8.720 1.210 9.000 1.260 ;
        RECT 8.720 0.660 8.990 1.210 ;
        RECT 8.830 0.010 8.990 0.660 ;
      LAYER via ;
        RECT 6.910 5.390 7.170 5.650 ;
        RECT 6.910 4.840 7.170 5.100 ;
        RECT 6.910 3.960 7.170 4.220 ;
        RECT 6.910 3.410 7.170 3.670 ;
        RECT 6.910 2.380 7.170 2.640 ;
        RECT 6.910 1.830 7.170 2.090 ;
        RECT 6.910 0.960 7.170 1.220 ;
        RECT 6.910 0.410 7.170 0.670 ;
      LAYER met2 ;
        RECT 6.880 5.550 7.190 5.690 ;
        RECT 0.000 5.370 9.350 5.550 ;
        RECT 6.880 5.360 7.190 5.370 ;
        RECT 6.880 5.120 7.190 5.140 ;
        RECT 0.000 4.940 9.350 5.120 ;
        RECT 6.880 4.810 7.190 4.940 ;
        RECT 6.880 4.120 7.190 4.250 ;
        RECT 0.000 3.940 9.350 4.120 ;
        RECT 6.880 3.920 7.190 3.940 ;
        RECT 6.880 3.690 7.190 3.700 ;
        RECT 0.000 3.620 6.870 3.690 ;
        RECT 6.880 3.620 9.350 3.690 ;
        RECT 0.000 3.510 9.350 3.620 ;
        RECT 6.880 3.370 7.190 3.510 ;
        RECT 6.880 2.540 7.190 2.680 ;
        RECT 6.880 2.530 9.350 2.540 ;
        RECT 0.000 2.360 9.350 2.530 ;
        RECT 6.880 2.350 7.190 2.360 ;
        RECT 6.880 2.110 7.190 2.130 ;
        RECT 0.000 1.940 9.350 2.110 ;
        RECT 6.790 1.930 9.350 1.940 ;
        RECT 6.880 1.800 7.190 1.930 ;
        RECT 6.880 1.130 7.190 1.250 ;
        RECT 0.000 1.120 7.190 1.130 ;
        RECT 0.000 0.960 9.350 1.120 ;
        RECT 6.790 0.940 9.350 0.960 ;
        RECT 6.880 0.920 7.190 0.940 ;
        RECT 6.880 0.690 7.190 0.700 ;
        RECT 0.000 0.520 9.350 0.690 ;
        RECT 6.880 0.510 9.350 0.520 ;
        RECT 6.880 0.370 7.190 0.510 ;
  END
END sky130_hilas_swc4x1cellOverlap2

MACRO sky130_hilas_TA2SignalBiasCell
  CLASS CORE ;
  FOREIGN sky130_hilas_TA2SignalBiasCell ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.880 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VOUT_AMP2
    USE ANALOG ;
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER met2 ;
        RECT 5.960 3.570 6.270 3.620 ;
        RECT 8.260 3.570 8.570 3.590 ;
        RECT 5.960 3.340 8.880 3.570 ;
        RECT 5.960 3.290 6.270 3.340 ;
        RECT 8.260 3.260 8.570 3.340 ;
    END
  END VOUT_AMP2
  PIN VOUT_AMP1
    USE ANALOG ;
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER met2 ;
        RECT 5.960 2.740 6.270 2.800 ;
        RECT 8.250 2.740 8.560 2.870 ;
        RECT 5.960 2.520 8.880 2.740 ;
        RECT 5.960 2.470 6.270 2.520 ;
    END
  END VOUT_AMP1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 6.920 0.000 7.260 6.050 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.000 6.040 4.040 6.050 ;
        RECT 0.000 0.010 5.600 6.040 ;
        RECT 3.740 0.000 5.600 0.010 ;
        RECT 7.600 0.000 8.880 6.050 ;
      LAYER met2 ;
        RECT 0.790 5.870 1.030 6.050 ;
        RECT 0.750 5.580 1.060 5.870 ;
        RECT 0.270 5.540 1.060 5.580 ;
        RECT 0.270 5.230 1.030 5.540 ;
        RECT 0.270 5.000 4.810 5.230 ;
        RECT 0.270 4.760 1.030 5.000 ;
        RECT 0.270 4.750 0.720 4.760 ;
        RECT 4.580 4.640 4.810 5.000 ;
        RECT 7.600 4.640 7.930 4.790 ;
        RECT 4.580 4.440 7.930 4.640 ;
        RECT 4.840 4.430 7.930 4.440 ;
        RECT 7.600 3.860 7.930 4.430 ;
        RECT 0.710 1.380 1.020 1.710 ;
    END
    PORT
      LAYER met1 ;
        RECT 7.590 4.790 7.860 6.050 ;
        RECT 7.590 3.860 7.940 4.790 ;
        RECT 7.590 1.880 7.860 3.860 ;
        RECT 7.590 1.590 7.870 1.880 ;
        RECT 7.590 0.000 7.860 1.590 ;
      LAYER via ;
        RECT 7.630 3.890 7.890 4.750 ;
    END
  END VPWR
  PIN VIN22
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT 4.390 6.030 4.640 6.040 ;
        RECT 4.990 6.030 5.300 6.040 ;
        RECT 4.390 5.780 5.300 6.030 ;
        RECT 4.990 5.710 5.300 5.780 ;
    END
  END VIN22
  PIN VIN21
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT 4.750 3.350 5.060 3.390 ;
        RECT 4.660 3.340 5.090 3.350 ;
        RECT 4.430 3.110 5.530 3.340 ;
        RECT 4.750 3.060 5.060 3.110 ;
    END
  END VIN21
  PIN VIN11
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT 3.190 2.940 3.500 2.990 ;
        RECT 2.870 2.710 3.970 2.940 ;
        RECT 2.870 2.700 3.530 2.710 ;
        RECT 3.190 2.660 3.500 2.700 ;
    END
  END VIN11
  PIN VIN12
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT 3.430 0.270 3.740 0.340 ;
        RECT 2.830 0.020 3.740 0.270 ;
        RECT 3.430 0.010 3.740 0.020 ;
    END
  END VIN12
  PIN VBIAS2
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT 1.680 0.270 1.990 0.340 ;
        RECT 1.110 0.260 1.990 0.270 ;
        RECT 0.050 0.030 1.990 0.260 ;
        RECT 1.110 0.020 1.990 0.030 ;
        RECT 1.680 0.010 1.990 0.020 ;
    END
  END VBIAS2
  PIN VBIAS1
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT 1.440 2.940 1.750 2.990 ;
        RECT 0.010 2.710 2.220 2.940 ;
        RECT 0.010 2.700 1.780 2.710 ;
        RECT 0.010 2.690 0.650 2.700 ;
        RECT 1.440 2.660 1.750 2.700 ;
    END
  END VBIAS1
  OBS
      LAYER li1 ;
        RECT 4.730 6.000 4.900 6.050 ;
        RECT 0.760 5.790 1.080 5.830 ;
        RECT 0.760 5.600 1.090 5.790 ;
        RECT 4.730 5.740 5.290 6.000 ;
        RECT 4.730 5.720 4.900 5.740 ;
        RECT 6.200 5.720 6.400 5.760 ;
        RECT 0.760 5.580 1.080 5.600 ;
        RECT 0.670 5.570 1.080 5.580 ;
        RECT 0.420 5.380 1.020 5.570 ;
        RECT 0.250 4.840 1.020 5.380 ;
        RECT 0.250 3.510 0.420 4.840 ;
        RECT 0.260 0.570 0.430 2.350 ;
        RECT 0.840 1.670 1.020 4.840 ;
        RECT 1.650 4.550 1.820 5.570 ;
        RECT 1.600 4.510 1.920 4.550 ;
        RECT 1.600 4.320 1.930 4.510 ;
        RECT 1.600 4.290 1.920 4.320 ;
        RECT 1.650 3.790 1.820 4.290 ;
        RECT 1.570 3.730 2.110 3.790 ;
        RECT 1.570 3.620 2.120 3.730 ;
        RECT 1.930 3.500 2.120 3.620 ;
        RECT 1.400 3.200 1.570 3.360 ;
        RECT 1.400 3.030 1.620 3.200 ;
        RECT 1.450 2.950 1.620 3.030 ;
        RECT 1.450 2.910 1.770 2.950 ;
        RECT 1.450 2.720 1.780 2.910 ;
        RECT 1.450 2.690 1.770 2.720 ;
        RECT 0.720 1.630 1.040 1.670 ;
        RECT 0.720 1.440 1.050 1.630 ;
        RECT 0.720 1.410 1.040 1.440 ;
        RECT 0.840 0.480 1.020 1.410 ;
        RECT 1.650 1.140 1.820 2.520 ;
        RECT 2.590 1.670 2.770 5.580 ;
        RECT 3.400 3.790 3.570 5.570 ;
        RECT 4.150 4.640 4.330 5.570 ;
        RECT 4.880 5.310 5.210 5.480 ;
        RECT 5.970 5.460 6.400 5.720 ;
        RECT 6.200 5.430 6.400 5.460 ;
        RECT 4.960 5.170 5.210 5.310 ;
        RECT 4.960 4.910 5.440 5.170 ;
        RECT 5.790 5.070 5.960 5.110 ;
        RECT 6.200 5.070 6.400 5.100 ;
        RECT 4.030 4.610 4.350 4.640 ;
        RECT 4.030 4.420 4.360 4.610 ;
        RECT 4.030 4.380 4.350 4.420 ;
        RECT 3.320 3.730 3.860 3.790 ;
        RECT 3.320 3.620 3.870 3.730 ;
        RECT 3.680 3.500 3.870 3.620 ;
        RECT 3.150 3.200 3.320 3.360 ;
        RECT 3.150 3.030 3.370 3.200 ;
        RECT 3.200 2.950 3.370 3.030 ;
        RECT 3.200 2.910 3.520 2.950 ;
        RECT 3.200 2.720 3.530 2.910 ;
        RECT 3.200 2.690 3.520 2.720 ;
        RECT 2.470 1.630 2.790 1.670 ;
        RECT 2.470 1.440 2.800 1.630 ;
        RECT 2.470 1.410 2.790 1.440 ;
        RECT 1.650 0.880 2.130 1.140 ;
        RECT 1.650 0.740 1.900 0.880 ;
        RECT 1.570 0.570 1.900 0.740 ;
        RECT 2.590 0.480 2.770 1.410 ;
        RECT 3.400 1.140 3.570 2.520 ;
        RECT 3.400 0.880 3.880 1.140 ;
        RECT 3.400 0.740 3.650 0.880 ;
        RECT 3.320 0.570 3.650 0.740 ;
        RECT 4.150 0.470 4.330 4.380 ;
        RECT 4.960 3.530 5.130 4.910 ;
        RECT 5.790 4.810 6.400 5.070 ;
        RECT 5.790 4.780 5.960 4.810 ;
        RECT 6.200 4.770 6.400 4.810 ;
        RECT 6.790 4.770 7.340 5.760 ;
        RECT 8.160 5.640 8.740 5.810 ;
        RECT 8.160 5.540 8.550 5.640 ;
        RECT 8.160 5.510 8.540 5.540 ;
        RECT 8.160 5.360 8.520 5.510 ;
        RECT 7.810 5.190 8.520 5.360 ;
        RECT 5.790 4.240 5.960 4.270 ;
        RECT 6.200 4.240 6.400 4.280 ;
        RECT 5.790 3.980 6.400 4.240 ;
        RECT 5.790 3.940 5.960 3.980 ;
        RECT 6.200 3.950 6.400 3.980 ;
        RECT 6.200 3.590 6.400 3.620 ;
        RECT 4.760 3.330 5.080 3.360 ;
        RECT 5.970 3.330 6.400 3.590 ;
        RECT 4.760 3.140 5.090 3.330 ;
        RECT 6.200 3.290 6.400 3.330 ;
        RECT 6.790 3.290 7.340 4.280 ;
        RECT 7.650 3.870 8.510 4.750 ;
        RECT 7.650 3.860 7.860 3.870 ;
        RECT 8.270 3.510 8.590 3.550 ;
        RECT 8.270 3.450 8.600 3.510 ;
        RECT 7.800 3.320 8.600 3.450 ;
        RECT 7.800 3.290 8.590 3.320 ;
        RECT 7.800 3.270 8.500 3.290 ;
        RECT 4.760 3.100 5.080 3.140 ;
        RECT 4.760 3.020 4.930 3.100 ;
        RECT 4.710 2.850 4.930 3.020 ;
        RECT 4.710 2.690 4.880 2.850 ;
        RECT 6.200 2.760 6.400 2.800 ;
        RECT 5.240 2.430 5.430 2.550 ;
        RECT 5.970 2.500 6.400 2.760 ;
        RECT 6.200 2.470 6.400 2.500 ;
        RECT 4.880 2.320 5.430 2.430 ;
        RECT 4.880 2.260 5.420 2.320 ;
        RECT 4.960 0.480 5.130 2.260 ;
        RECT 5.790 2.110 5.960 2.150 ;
        RECT 6.200 2.110 6.400 2.140 ;
        RECT 5.790 1.850 6.400 2.110 ;
        RECT 5.790 1.820 5.960 1.850 ;
        RECT 6.200 1.810 6.400 1.850 ;
        RECT 6.790 1.810 7.340 2.800 ;
        RECT 8.260 2.790 8.580 2.830 ;
        RECT 7.800 2.610 8.590 2.790 ;
        RECT 8.260 2.600 8.590 2.610 ;
        RECT 8.260 2.570 8.580 2.600 ;
        RECT 7.810 1.850 8.510 2.190 ;
        RECT 7.660 1.620 8.510 1.850 ;
        RECT 5.790 1.280 5.960 1.310 ;
        RECT 6.200 1.280 6.400 1.320 ;
        RECT 5.790 1.020 6.400 1.280 ;
        RECT 5.790 0.980 5.960 1.020 ;
        RECT 6.200 0.990 6.400 1.020 ;
        RECT 6.200 0.630 6.400 0.660 ;
        RECT 5.970 0.370 6.400 0.630 ;
        RECT 6.200 0.330 6.400 0.370 ;
        RECT 6.790 0.330 7.340 1.320 ;
        RECT 7.810 1.310 8.510 1.620 ;
        RECT 7.810 0.700 8.520 0.870 ;
        RECT 8.160 0.420 8.520 0.700 ;
        RECT 1.420 0.310 1.590 0.330 ;
        RECT 3.170 0.310 3.340 0.330 ;
        RECT 1.420 0.050 1.980 0.310 ;
        RECT 3.170 0.050 3.730 0.310 ;
        RECT 8.160 0.250 8.740 0.420 ;
        RECT 1.420 0.000 1.590 0.050 ;
        RECT 3.170 0.000 3.340 0.050 ;
      LAYER mcon ;
        RECT 0.820 5.610 0.990 5.780 ;
        RECT 5.060 5.780 5.230 5.950 ;
        RECT 0.250 5.210 0.420 5.380 ;
        RECT 0.840 5.160 1.010 5.330 ;
        RECT 0.250 4.870 0.420 5.040 ;
        RECT 0.250 4.530 0.420 4.700 ;
        RECT 0.250 4.190 0.420 4.360 ;
        RECT 0.250 3.850 0.420 4.020 ;
        RECT 0.840 4.820 1.010 4.990 ;
        RECT 0.260 2.180 0.430 2.350 ;
        RECT 0.260 1.840 0.430 2.010 ;
        RECT 1.660 4.330 1.830 4.500 ;
        RECT 1.940 3.530 2.110 3.700 ;
        RECT 1.510 2.730 1.680 2.900 ;
        RECT 0.260 1.500 0.430 1.670 ;
        RECT 0.780 1.450 0.950 1.620 ;
        RECT 0.260 1.160 0.430 1.330 ;
        RECT 0.260 0.820 0.430 0.990 ;
        RECT 6.030 5.500 6.200 5.670 ;
        RECT 8.280 5.550 8.450 5.720 ;
        RECT 7.010 5.180 7.180 5.350 ;
        RECT 5.210 4.950 5.380 5.120 ;
        RECT 4.090 4.430 4.260 4.600 ;
        RECT 3.690 3.530 3.860 3.700 ;
        RECT 3.260 2.730 3.430 2.900 ;
        RECT 2.530 1.450 2.700 1.620 ;
        RECT 1.900 0.930 2.070 1.100 ;
        RECT 3.650 0.930 3.820 1.100 ;
        RECT 5.980 4.850 6.150 5.020 ;
        RECT 7.670 4.580 7.840 4.750 ;
        RECT 5.980 4.030 6.150 4.200 ;
        RECT 7.010 3.700 7.180 3.870 ;
        RECT 7.670 4.240 7.840 4.410 ;
        RECT 7.670 3.880 7.840 4.050 ;
        RECT 6.030 3.380 6.200 3.550 ;
        RECT 4.820 3.150 4.990 3.320 ;
        RECT 8.330 3.330 8.500 3.500 ;
        RECT 5.250 2.350 5.420 2.520 ;
        RECT 6.030 2.540 6.200 2.710 ;
        RECT 8.320 2.610 8.490 2.780 ;
        RECT 7.010 2.220 7.180 2.390 ;
        RECT 5.980 1.890 6.150 2.060 ;
        RECT 7.670 1.650 7.840 1.820 ;
        RECT 5.980 1.070 6.150 1.240 ;
        RECT 7.010 0.740 7.180 0.910 ;
        RECT 6.030 0.420 6.200 0.590 ;
        RECT 8.240 0.360 8.410 0.530 ;
        RECT 1.750 0.100 1.920 0.270 ;
        RECT 3.500 0.100 3.670 0.270 ;
      LAYER met1 ;
        RECT 0.750 5.590 1.070 5.860 ;
        RECT 4.980 5.710 5.300 6.030 ;
        RECT 0.220 5.540 1.070 5.590 ;
        RECT 0.220 5.270 1.040 5.540 ;
        RECT 5.960 5.430 6.280 5.750 ;
        RECT 8.210 5.480 8.530 5.800 ;
        RECT 0.220 4.980 1.070 5.270 ;
        RECT 0.220 4.730 1.040 4.980 ;
        RECT 5.130 4.880 5.450 5.200 ;
        RECT 5.910 4.780 6.230 5.100 ;
        RECT 0.220 1.700 0.860 4.730 ;
        RECT 1.590 4.260 1.910 4.580 ;
        RECT 4.020 4.350 4.340 4.670 ;
        RECT 5.240 4.190 5.450 4.300 ;
        RECT 5.220 3.870 5.480 4.190 ;
        RECT 5.910 3.950 6.230 4.270 ;
        RECT 1.910 3.470 2.140 3.760 ;
        RECT 3.660 3.470 3.890 3.760 ;
        RECT 1.440 2.660 1.760 2.980 ;
        RECT 1.930 2.180 2.140 3.470 ;
        RECT 3.190 2.660 3.510 2.980 ;
        RECT 3.680 2.180 3.890 3.470 ;
        RECT 4.750 3.070 5.070 3.390 ;
        RECT 5.240 2.580 5.450 3.870 ;
        RECT 5.960 3.300 6.280 3.620 ;
        RECT 8.260 3.260 8.580 3.580 ;
        RECT 5.220 2.290 5.450 2.580 ;
        RECT 5.960 2.470 6.280 2.790 ;
        RECT 8.250 2.540 8.570 2.860 ;
        RECT 1.910 1.860 2.170 2.180 ;
        RECT 3.660 1.860 3.920 2.180 ;
        RECT 1.930 1.750 2.140 1.860 ;
        RECT 3.680 1.750 3.890 1.860 ;
        RECT 5.910 1.820 6.230 2.140 ;
        RECT 0.220 1.380 1.030 1.700 ;
        RECT 2.460 1.380 2.780 1.700 ;
        RECT 0.220 0.550 0.860 1.380 ;
        RECT 1.820 0.850 2.140 1.170 ;
        RECT 3.570 0.850 3.890 1.170 ;
        RECT 5.910 0.990 6.230 1.310 ;
        RECT 0.440 0.540 0.860 0.550 ;
        RECT 5.960 0.340 6.280 0.660 ;
        RECT 1.670 0.020 1.990 0.340 ;
        RECT 3.420 0.020 3.740 0.340 ;
        RECT 8.170 0.290 8.490 0.610 ;
      LAYER via ;
        RECT 0.780 5.570 1.040 5.830 ;
        RECT 5.010 5.740 5.270 6.000 ;
        RECT 0.340 4.790 0.930 5.510 ;
        RECT 5.990 5.460 6.250 5.720 ;
        RECT 8.240 5.510 8.500 5.770 ;
        RECT 5.160 4.910 5.420 5.170 ;
        RECT 5.940 4.810 6.200 5.070 ;
        RECT 1.620 4.290 1.880 4.550 ;
        RECT 4.050 4.380 4.310 4.640 ;
        RECT 5.220 3.900 5.480 4.160 ;
        RECT 5.940 3.980 6.200 4.240 ;
        RECT 1.470 2.690 1.730 2.950 ;
        RECT 3.220 2.690 3.480 2.950 ;
        RECT 4.780 3.100 5.040 3.360 ;
        RECT 5.990 3.330 6.250 3.590 ;
        RECT 8.290 3.290 8.550 3.550 ;
        RECT 5.990 2.500 6.250 2.760 ;
        RECT 8.280 2.570 8.540 2.830 ;
        RECT 1.910 1.890 2.170 2.150 ;
        RECT 3.660 1.890 3.920 2.150 ;
        RECT 5.940 1.850 6.200 2.110 ;
        RECT 0.740 1.410 1.000 1.670 ;
        RECT 2.490 1.410 2.750 1.670 ;
        RECT 1.850 0.880 2.110 1.140 ;
        RECT 3.600 0.880 3.860 1.140 ;
        RECT 5.940 1.020 6.200 1.280 ;
        RECT 5.990 0.370 6.250 0.630 ;
        RECT 1.700 0.050 1.960 0.310 ;
        RECT 3.450 0.050 3.710 0.310 ;
        RECT 8.200 0.320 8.460 0.580 ;
      LAYER met2 ;
        RECT 5.960 5.710 6.270 5.760 ;
        RECT 8.210 5.710 8.520 5.810 ;
        RECT 5.960 5.480 8.520 5.710 ;
        RECT 5.960 5.430 6.270 5.480 ;
        RECT 5.140 5.170 5.450 5.210 ;
        RECT 4.960 5.030 5.700 5.170 ;
        RECT 5.910 5.030 6.220 5.110 ;
        RECT 4.960 4.920 6.220 5.030 ;
        RECT 5.140 4.880 6.220 4.920 ;
        RECT 5.450 4.820 6.220 4.880 ;
        RECT 5.450 4.800 5.700 4.820 ;
        RECT 5.910 4.780 6.220 4.820 ;
        RECT 1.590 4.530 1.900 4.590 ;
        RECT 4.020 4.530 4.330 4.670 ;
        RECT 1.590 4.340 4.330 4.530 ;
        RECT 1.590 4.310 4.070 4.340 ;
        RECT 1.590 4.260 1.900 4.310 ;
        RECT 5.480 4.230 5.690 4.240 ;
        RECT 5.910 4.230 6.220 4.270 ;
        RECT 5.480 4.160 6.220 4.230 ;
        RECT 5.190 4.140 6.220 4.160 ;
        RECT 5.140 4.020 6.220 4.140 ;
        RECT 5.140 3.950 5.690 4.020 ;
        RECT 5.140 3.890 5.610 3.950 ;
        RECT 5.910 3.940 6.220 4.020 ;
        RECT 1.830 1.910 2.300 2.160 ;
        RECT 3.580 2.070 4.050 2.160 ;
        RECT 5.910 2.070 6.220 2.150 ;
        RECT 3.580 1.910 6.220 2.070 ;
        RECT 1.880 1.890 2.200 1.910 ;
        RECT 3.630 1.890 6.220 1.910 ;
        RECT 3.920 1.870 6.220 1.890 ;
        RECT 5.610 1.860 6.220 1.870 ;
        RECT 5.910 1.820 6.220 1.860 ;
        RECT 2.460 1.700 2.770 1.710 ;
        RECT 2.350 1.520 2.770 1.700 ;
        RECT 2.330 1.510 2.770 1.520 ;
        RECT 2.110 1.380 2.770 1.510 ;
        RECT 2.110 1.170 2.470 1.380 ;
        RECT 5.910 1.270 6.220 1.310 ;
        RECT 3.630 1.170 6.220 1.270 ;
        RECT 1.830 1.130 2.470 1.170 ;
        RECT 3.580 1.130 6.220 1.170 ;
        RECT 1.650 0.890 2.470 1.130 ;
        RECT 3.400 1.060 6.220 1.130 ;
        RECT 1.650 0.880 2.200 0.890 ;
        RECT 3.400 0.880 3.950 1.060 ;
        RECT 5.910 0.980 6.220 1.060 ;
        RECT 1.830 0.840 2.140 0.880 ;
        RECT 3.580 0.840 3.890 0.880 ;
        RECT 5.960 0.580 6.270 0.660 ;
        RECT 8.170 0.580 8.480 0.620 ;
        RECT 5.960 0.350 8.670 0.580 ;
        RECT 5.960 0.330 6.270 0.350 ;
        RECT 8.170 0.290 8.480 0.350 ;
  END
END sky130_hilas_TA2SignalBiasCell

MACRO sky130_hilas_Tgate4Single01
  CLASS CORE ;
  FOREIGN sky130_hilas_Tgate4Single01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.760 BY 6.050 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN INPUT1_4
    USE ANALOG ;
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 1.640 0.320 1.950 0.440 ;
        RECT 0.870 0.310 1.990 0.320 ;
        RECT 3.210 0.310 3.520 0.440 ;
        RECT 0.000 0.110 3.520 0.310 ;
        RECT 0.870 0.100 1.990 0.110 ;
    END
  END INPUT1_4
  PIN VPWR
    USE ANALOG ;
    ANTENNADIFFAREA 0.908800 ;
    PORT
      LAYER nwell ;
        RECT 0.120 0.000 2.880 6.050 ;
      LAYER met1 ;
        RECT 0.740 5.180 0.940 6.050 ;
        RECT 0.730 4.890 0.960 5.180 ;
        RECT 0.740 4.180 0.940 4.890 ;
        RECT 0.730 3.890 0.960 4.180 ;
        RECT 0.740 2.160 0.940 3.890 ;
        RECT 0.730 1.870 0.960 2.160 ;
        RECT 0.740 1.160 0.940 1.870 ;
        RECT 0.730 0.870 0.960 1.160 ;
        RECT 0.740 0.000 0.940 0.870 ;
    END
  END VPWR
  PIN SELECT4
    USE ANALOG ;
    ANTENNAGATEAREA 0.372000 ;
    PORT
      LAYER met2 ;
        RECT 0.290 1.290 0.610 1.380 ;
        RECT 0.000 1.090 0.610 1.290 ;
    END
  END SELECT4
  PIN SELECT3
    USE ANALOG ;
    ANTENNAGATEAREA 0.372000 ;
    PORT
      LAYER met2 ;
        RECT 0.000 1.740 0.610 1.940 ;
        RECT 0.290 1.650 0.610 1.740 ;
    END
  END SELECT3
  PIN INPUT1_3
    USE ANALOG ;
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 0.870 2.920 1.990 2.930 ;
        RECT 0.000 2.720 3.520 2.920 ;
        RECT 0.870 2.710 1.990 2.720 ;
        RECT 1.640 2.590 1.950 2.710 ;
        RECT 3.210 2.590 3.520 2.720 ;
    END
  END INPUT1_3
  PIN INPUT1_2
    USE ANALOG ;
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 1.640 3.340 1.950 3.460 ;
        RECT 0.870 3.330 1.990 3.340 ;
        RECT 3.210 3.330 3.520 3.460 ;
        RECT 0.000 3.130 3.520 3.330 ;
        RECT 0.870 3.120 1.990 3.130 ;
    END
  END INPUT1_2
  PIN SELECT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.372000 ;
    PORT
      LAYER met2 ;
        RECT 0.290 4.310 0.610 4.400 ;
        RECT 0.000 4.110 0.610 4.310 ;
    END
  END SELECT2
  PIN SELECT1
    USE ANALOG ;
    ANTENNAGATEAREA 0.372000 ;
    PORT
      LAYER met2 ;
        RECT 0.000 4.760 0.610 4.960 ;
        RECT 0.290 4.670 0.610 4.760 ;
    END
  END SELECT1
  PIN INPUT1_1
    USE ANALOG ;
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 0.870 5.940 1.990 5.950 ;
        RECT 0.000 5.740 3.520 5.940 ;
        RECT 0.870 5.730 1.990 5.740 ;
        RECT 1.640 5.610 1.950 5.730 ;
        RECT 3.210 5.610 3.520 5.740 ;
    END
  END INPUT1_1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 4.250 5.180 4.440 6.050 ;
        RECT 4.230 4.890 4.460 5.180 ;
        RECT 4.250 4.180 4.440 4.890 ;
        RECT 4.230 3.890 4.460 4.180 ;
        RECT 4.250 2.160 4.440 3.890 ;
        RECT 4.230 1.870 4.460 2.160 ;
        RECT 4.250 1.160 4.440 1.870 ;
        RECT 4.230 0.870 4.460 1.160 ;
        RECT 4.250 0.000 4.440 0.870 ;
    END
  END VGND
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.182900 ;
    PORT
      LAYER met2 ;
        RECT 2.560 4.960 2.880 5.000 ;
        RECT 3.570 4.960 3.890 4.990 ;
        RECT 2.510 4.760 4.760 4.960 ;
        RECT 2.560 4.740 2.880 4.760 ;
        RECT 3.570 4.730 3.890 4.760 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.182900 ;
    PORT
      LAYER met2 ;
        RECT 2.560 4.310 2.880 4.330 ;
        RECT 3.570 4.310 3.890 4.340 ;
        RECT 2.510 4.110 4.760 4.310 ;
        RECT 2.560 4.070 2.880 4.110 ;
        RECT 3.570 4.080 3.890 4.110 ;
    END
  END OUTPUT2
  PIN OUTPUT3
    USE ANALOG ;
    ANTENNADIFFAREA 0.182900 ;
    PORT
      LAYER met2 ;
        RECT 2.560 1.940 2.880 1.980 ;
        RECT 3.570 1.940 3.890 1.970 ;
        RECT 2.510 1.740 4.760 1.940 ;
        RECT 2.560 1.720 2.880 1.740 ;
        RECT 3.570 1.710 3.890 1.740 ;
    END
  END OUTPUT3
  PIN OUTPUT4
    USE ANALOG ;
    ANTENNADIFFAREA 0.182900 ;
    PORT
      LAYER met2 ;
        RECT 2.560 1.290 2.880 1.310 ;
        RECT 3.570 1.290 3.890 1.320 ;
        RECT 2.510 1.090 4.760 1.290 ;
        RECT 2.560 1.050 2.880 1.090 ;
        RECT 3.570 1.060 3.890 1.090 ;
    END
  END OUTPUT4
  OBS
      LAYER li1 ;
        RECT 1.650 5.880 1.970 5.910 ;
        RECT 3.220 5.880 3.540 5.910 ;
        RECT 0.430 5.540 0.600 5.820 ;
        RECT 1.650 5.690 1.980 5.880 ;
        RECT 2.660 5.740 2.850 5.760 ;
        RECT 1.650 5.650 1.970 5.690 ;
        RECT 0.430 5.500 0.640 5.540 ;
        RECT 0.430 5.480 0.660 5.500 ;
        RECT 1.780 5.490 1.950 5.650 ;
        RECT 2.390 5.570 2.850 5.740 ;
        RECT 3.220 5.690 3.550 5.880 ;
        RECT 3.790 5.740 3.980 5.770 ;
        RECT 3.220 5.650 3.540 5.690 ;
        RECT 2.640 5.560 2.850 5.570 ;
        RECT 2.660 5.530 2.850 5.560 ;
        RECT 3.280 5.490 3.450 5.650 ;
        RECT 3.790 5.570 4.230 5.740 ;
        RECT 3.790 5.540 3.980 5.570 ;
        RECT 0.430 5.460 0.690 5.480 ;
        RECT 0.430 5.410 0.770 5.460 ;
        RECT 0.430 5.350 0.920 5.410 ;
        RECT 0.430 5.320 0.940 5.350 ;
        RECT 0.470 5.290 0.940 5.320 ;
        RECT 0.600 5.240 0.940 5.290 ;
        RECT 0.720 5.230 0.940 5.240 ;
        RECT 0.730 5.200 0.940 5.230 ;
        RECT 0.750 5.120 0.940 5.200 ;
        RECT 2.110 5.120 2.440 5.240 ;
        RECT 4.510 5.150 4.680 5.830 ;
        RECT 0.260 5.070 0.430 5.090 ;
        RECT 0.240 4.640 0.450 5.070 ;
        RECT 0.750 4.950 1.270 5.120 ;
        RECT 0.750 4.920 0.940 4.950 ;
        RECT 1.620 4.940 3.520 5.120 ;
        RECT 4.250 5.110 4.680 5.150 ;
        RECT 3.900 4.950 4.680 5.110 ;
        RECT 3.900 4.940 4.440 4.950 ;
        RECT 4.250 4.920 4.440 4.940 ;
        RECT 0.240 4.000 0.450 4.430 ;
        RECT 0.750 4.120 0.940 4.150 ;
        RECT 4.250 4.130 4.440 4.150 ;
        RECT 0.260 3.980 0.430 4.000 ;
        RECT 0.750 3.950 1.270 4.120 ;
        RECT 1.620 3.950 3.520 4.130 ;
        RECT 3.900 4.120 4.440 4.130 ;
        RECT 3.900 3.960 4.680 4.120 ;
        RECT 0.750 3.870 0.940 3.950 ;
        RECT 0.730 3.840 0.940 3.870 ;
        RECT 0.720 3.830 0.940 3.840 ;
        RECT 2.110 3.830 2.440 3.950 ;
        RECT 4.250 3.920 4.680 3.960 ;
        RECT 0.600 3.780 0.940 3.830 ;
        RECT 0.470 3.750 0.940 3.780 ;
        RECT 0.430 3.720 0.940 3.750 ;
        RECT 0.430 3.660 0.920 3.720 ;
        RECT 0.430 3.610 0.770 3.660 ;
        RECT 0.430 3.590 0.690 3.610 ;
        RECT 0.430 3.570 0.660 3.590 ;
        RECT 0.430 3.530 0.640 3.570 ;
        RECT 0.430 3.250 0.600 3.530 ;
        RECT 1.780 3.420 1.950 3.580 ;
        RECT 2.660 3.510 2.850 3.540 ;
        RECT 2.640 3.500 2.850 3.510 ;
        RECT 1.650 3.380 1.970 3.420 ;
        RECT 1.650 3.190 1.980 3.380 ;
        RECT 2.390 3.330 2.850 3.500 ;
        RECT 3.280 3.420 3.450 3.580 ;
        RECT 3.790 3.500 3.980 3.530 ;
        RECT 2.660 3.310 2.850 3.330 ;
        RECT 3.220 3.380 3.540 3.420 ;
        RECT 3.220 3.190 3.550 3.380 ;
        RECT 3.790 3.330 4.230 3.500 ;
        RECT 3.790 3.300 3.980 3.330 ;
        RECT 4.510 3.240 4.680 3.920 ;
        RECT 1.650 3.160 1.970 3.190 ;
        RECT 3.220 3.160 3.540 3.190 ;
        RECT 1.650 2.860 1.970 2.890 ;
        RECT 3.220 2.860 3.540 2.890 ;
        RECT 0.430 2.520 0.600 2.800 ;
        RECT 1.650 2.670 1.980 2.860 ;
        RECT 2.660 2.720 2.850 2.740 ;
        RECT 1.650 2.630 1.970 2.670 ;
        RECT 0.430 2.480 0.640 2.520 ;
        RECT 0.430 2.460 0.660 2.480 ;
        RECT 1.780 2.470 1.950 2.630 ;
        RECT 2.390 2.550 2.850 2.720 ;
        RECT 3.220 2.670 3.550 2.860 ;
        RECT 3.790 2.720 3.980 2.750 ;
        RECT 3.220 2.630 3.540 2.670 ;
        RECT 2.640 2.540 2.850 2.550 ;
        RECT 2.660 2.510 2.850 2.540 ;
        RECT 3.280 2.470 3.450 2.630 ;
        RECT 3.790 2.550 4.230 2.720 ;
        RECT 3.790 2.520 3.980 2.550 ;
        RECT 0.430 2.440 0.690 2.460 ;
        RECT 0.430 2.390 0.770 2.440 ;
        RECT 0.430 2.330 0.920 2.390 ;
        RECT 0.430 2.300 0.940 2.330 ;
        RECT 0.470 2.270 0.940 2.300 ;
        RECT 0.600 2.220 0.940 2.270 ;
        RECT 0.720 2.210 0.940 2.220 ;
        RECT 0.730 2.180 0.940 2.210 ;
        RECT 0.750 2.100 0.940 2.180 ;
        RECT 2.110 2.100 2.440 2.220 ;
        RECT 4.510 2.130 4.680 2.810 ;
        RECT 0.260 2.050 0.430 2.070 ;
        RECT 0.240 1.620 0.450 2.050 ;
        RECT 0.750 1.930 1.270 2.100 ;
        RECT 0.750 1.900 0.940 1.930 ;
        RECT 1.620 1.920 3.520 2.100 ;
        RECT 4.250 2.090 4.680 2.130 ;
        RECT 3.900 1.930 4.680 2.090 ;
        RECT 3.900 1.920 4.440 1.930 ;
        RECT 4.250 1.900 4.440 1.920 ;
        RECT 0.240 0.980 0.450 1.410 ;
        RECT 0.750 1.100 0.940 1.130 ;
        RECT 4.250 1.110 4.440 1.130 ;
        RECT 0.260 0.960 0.430 0.980 ;
        RECT 0.750 0.930 1.270 1.100 ;
        RECT 1.620 0.930 3.520 1.110 ;
        RECT 3.900 1.100 4.440 1.110 ;
        RECT 3.900 0.940 4.680 1.100 ;
        RECT 0.750 0.850 0.940 0.930 ;
        RECT 0.730 0.820 0.940 0.850 ;
        RECT 0.720 0.810 0.940 0.820 ;
        RECT 2.110 0.810 2.440 0.930 ;
        RECT 4.250 0.900 4.680 0.940 ;
        RECT 0.600 0.760 0.940 0.810 ;
        RECT 0.470 0.730 0.940 0.760 ;
        RECT 0.430 0.700 0.940 0.730 ;
        RECT 0.430 0.640 0.920 0.700 ;
        RECT 0.430 0.590 0.770 0.640 ;
        RECT 0.430 0.570 0.690 0.590 ;
        RECT 0.430 0.550 0.660 0.570 ;
        RECT 0.430 0.510 0.640 0.550 ;
        RECT 0.430 0.230 0.600 0.510 ;
        RECT 1.780 0.400 1.950 0.560 ;
        RECT 2.660 0.490 2.850 0.520 ;
        RECT 2.640 0.480 2.850 0.490 ;
        RECT 1.650 0.360 1.970 0.400 ;
        RECT 1.650 0.170 1.980 0.360 ;
        RECT 2.390 0.310 2.850 0.480 ;
        RECT 3.280 0.400 3.450 0.560 ;
        RECT 3.790 0.480 3.980 0.510 ;
        RECT 2.660 0.290 2.850 0.310 ;
        RECT 3.220 0.360 3.540 0.400 ;
        RECT 3.220 0.170 3.550 0.360 ;
        RECT 3.790 0.310 4.230 0.480 ;
        RECT 3.790 0.280 3.980 0.310 ;
        RECT 4.510 0.220 4.680 0.900 ;
        RECT 1.650 0.140 1.970 0.170 ;
        RECT 3.220 0.140 3.540 0.170 ;
      LAYER mcon ;
        RECT 1.710 5.700 1.880 5.870 ;
        RECT 2.670 5.560 2.840 5.730 ;
        RECT 3.280 5.700 3.450 5.870 ;
        RECT 3.800 5.570 3.970 5.740 ;
        RECT 0.260 4.920 0.430 5.090 ;
        RECT 0.760 4.950 0.930 5.120 ;
        RECT 4.260 4.950 4.430 5.120 ;
        RECT 0.760 3.950 0.930 4.120 ;
        RECT 4.260 3.950 4.430 4.120 ;
        RECT 1.710 3.200 1.880 3.370 ;
        RECT 2.670 3.340 2.840 3.510 ;
        RECT 3.280 3.200 3.450 3.370 ;
        RECT 3.800 3.330 3.970 3.500 ;
        RECT 1.710 2.680 1.880 2.850 ;
        RECT 2.670 2.540 2.840 2.710 ;
        RECT 3.280 2.680 3.450 2.850 ;
        RECT 3.800 2.550 3.970 2.720 ;
        RECT 0.260 1.900 0.430 2.070 ;
        RECT 0.760 1.930 0.930 2.100 ;
        RECT 4.260 1.930 4.430 2.100 ;
        RECT 0.760 0.930 0.930 1.100 ;
        RECT 4.260 0.930 4.430 1.100 ;
        RECT 1.710 0.180 1.880 0.350 ;
        RECT 2.670 0.320 2.840 0.490 ;
        RECT 3.280 0.180 3.450 0.350 ;
        RECT 3.800 0.310 3.970 0.480 ;
      LAYER met1 ;
        RECT 1.640 5.620 1.960 5.940 ;
        RECT 2.640 5.500 2.870 5.790 ;
        RECT 3.210 5.620 3.530 5.940 ;
        RECT 3.770 5.510 4.000 5.800 ;
        RECT 0.230 4.960 0.460 5.150 ;
        RECT 2.660 5.030 2.850 5.500 ;
        RECT 0.230 4.860 0.580 4.960 ;
        RECT 0.240 4.640 0.580 4.860 ;
        RECT 2.590 4.710 2.850 5.030 ;
        RECT 3.770 5.020 3.960 5.510 ;
        RECT 3.600 4.770 3.960 5.020 ;
        RECT 3.600 4.700 3.860 4.770 ;
        RECT 0.240 4.210 0.580 4.430 ;
        RECT 0.230 4.110 0.580 4.210 ;
        RECT 0.230 3.920 0.460 4.110 ;
        RECT 2.590 4.040 2.850 4.360 ;
        RECT 3.600 4.300 3.860 4.370 ;
        RECT 3.600 4.050 3.960 4.300 ;
        RECT 2.660 3.570 2.850 4.040 ;
        RECT 1.640 3.130 1.960 3.450 ;
        RECT 2.640 3.280 2.870 3.570 ;
        RECT 3.770 3.560 3.960 4.050 ;
        RECT 3.210 3.130 3.530 3.450 ;
        RECT 3.770 3.270 4.000 3.560 ;
        RECT 1.640 2.600 1.960 2.920 ;
        RECT 2.640 2.480 2.870 2.770 ;
        RECT 3.210 2.600 3.530 2.920 ;
        RECT 3.770 2.490 4.000 2.780 ;
        RECT 0.230 1.940 0.460 2.130 ;
        RECT 2.660 2.010 2.850 2.480 ;
        RECT 0.230 1.840 0.580 1.940 ;
        RECT 0.240 1.620 0.580 1.840 ;
        RECT 2.590 1.690 2.850 2.010 ;
        RECT 3.770 2.000 3.960 2.490 ;
        RECT 3.600 1.750 3.960 2.000 ;
        RECT 3.600 1.680 3.860 1.750 ;
        RECT 0.240 1.190 0.580 1.410 ;
        RECT 0.230 1.090 0.580 1.190 ;
        RECT 0.230 0.900 0.460 1.090 ;
        RECT 2.590 1.020 2.850 1.340 ;
        RECT 3.600 1.280 3.860 1.350 ;
        RECT 3.600 1.030 3.960 1.280 ;
        RECT 2.660 0.550 2.850 1.020 ;
        RECT 1.640 0.110 1.960 0.430 ;
        RECT 2.640 0.260 2.870 0.550 ;
        RECT 3.770 0.540 3.960 1.030 ;
        RECT 3.210 0.110 3.530 0.430 ;
        RECT 3.770 0.250 4.000 0.540 ;
      LAYER via ;
        RECT 1.670 5.650 1.930 5.910 ;
        RECT 3.240 5.650 3.500 5.910 ;
        RECT 0.320 4.670 0.580 4.930 ;
        RECT 2.590 4.740 2.850 5.000 ;
        RECT 3.600 4.730 3.860 4.990 ;
        RECT 0.320 4.140 0.580 4.400 ;
        RECT 2.590 4.070 2.850 4.330 ;
        RECT 3.600 4.080 3.860 4.340 ;
        RECT 1.670 3.160 1.930 3.420 ;
        RECT 3.240 3.160 3.500 3.420 ;
        RECT 1.670 2.630 1.930 2.890 ;
        RECT 3.240 2.630 3.500 2.890 ;
        RECT 0.320 1.650 0.580 1.910 ;
        RECT 2.590 1.720 2.850 1.980 ;
        RECT 3.600 1.710 3.860 1.970 ;
        RECT 0.320 1.120 0.580 1.380 ;
        RECT 2.590 1.050 2.850 1.310 ;
        RECT 3.600 1.060 3.860 1.320 ;
        RECT 1.670 0.140 1.930 0.400 ;
        RECT 3.240 0.140 3.500 0.400 ;
  END
END sky130_hilas_Tgate4Single01

MACRO sky130_hilas_VinjDecode2to4
  CLASS CORE ;
  FOREIGN sky130_hilas_VinjDecode2to4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.320 BY 8.330 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN OUTPUT00
    PORT
      LAYER met2 ;
        RECT 12.820 6.270 12.950 6.440 ;
    END
  END OUTPUT00
  PIN OUTPUT01
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 12.940 5.010 13.310 5.090 ;
        RECT 12.940 5.000 13.970 5.010 ;
        RECT 15.850 5.000 16.160 5.160 ;
        RECT 12.940 4.930 16.320 5.000 ;
        RECT 12.820 4.830 16.320 4.930 ;
        RECT 12.820 4.760 12.950 4.830 ;
    END
  END OUTPUT01
  PIN OUTPUT10
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 12.940 3.500 13.310 3.580 ;
        RECT 12.940 3.490 13.970 3.500 ;
        RECT 15.850 3.490 16.160 3.650 ;
        RECT 12.940 3.420 16.320 3.490 ;
        RECT 12.820 3.320 16.320 3.420 ;
        RECT 12.820 3.250 12.950 3.320 ;
    END
  END OUTPUT10
  PIN OUTPUT11
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 12.940 1.990 13.310 2.070 ;
        RECT 12.940 1.980 13.970 1.990 ;
        RECT 15.850 1.980 16.160 2.140 ;
        RECT 12.940 1.920 16.320 1.980 ;
        RECT 12.820 1.810 16.320 1.920 ;
        RECT 12.820 1.750 12.950 1.810 ;
    END
  END OUTPUT11
  PIN VGND
    PORT
      LAYER met1 ;
        RECT 11.660 7.510 11.930 7.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.660 1.540 11.930 1.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.180 7.470 3.410 7.560 ;
    END
  END VGND
  PIN VINJ
    ANTENNADIFFAREA 0.691200 ;
    PORT
      LAYER met1 ;
        RECT 6.540 1.590 6.770 6.120 ;
        RECT 6.690 1.540 6.910 1.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.690 7.490 6.910 7.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.610 7.480 0.830 7.560 ;
    END
  END VINJ
  PIN IN2
    PORT
      LAYER met2 ;
        RECT 0.000 5.480 0.110 5.660 ;
    END
  END IN2
  PIN IN1
    PORT
      LAYER met2 ;
        RECT 0.000 6.990 0.110 7.170 ;
    END
  END IN1
  PIN ENABLE
    PORT
      LAYER met2 ;
        RECT 0.000 3.970 0.110 4.150 ;
    END
  END ENABLE
  OBS
      LAYER nwell ;
        RECT 6.690 7.490 6.910 7.550 ;
        RECT 3.360 1.500 5.340 6.160 ;
        RECT 6.690 1.540 6.910 1.590 ;
        RECT 9.450 0.000 12.890 6.160 ;
      LAYER li1 ;
        RECT 3.980 5.730 4.150 5.870 ;
        RECT 10.070 5.730 10.240 5.870 ;
        RECT 10.800 5.750 10.970 5.830 ;
        RECT 11.610 5.750 11.780 5.830 ;
        RECT 13.150 5.790 13.320 5.910 ;
        RECT 3.980 5.560 4.170 5.730 ;
        RECT 3.980 5.460 4.150 5.560 ;
        RECT 3.550 5.080 3.720 5.180 ;
        RECT 3.530 4.910 3.720 5.080 ;
        RECT 3.550 4.850 3.720 4.910 ;
        RECT 3.970 5.120 4.140 5.180 ;
        RECT 3.970 4.850 4.220 5.120 ;
        RECT 4.710 5.100 4.960 5.180 ;
        RECT 4.710 4.930 6.010 5.100 ;
        RECT 6.570 5.090 6.740 5.720 ;
        RECT 10.070 5.560 10.260 5.730 ;
        RECT 10.070 5.460 10.240 5.560 ;
        RECT 10.800 5.180 11.010 5.750 ;
        RECT 11.570 5.500 11.780 5.750 ;
        RECT 12.170 5.570 12.340 5.670 ;
        RECT 13.110 5.620 13.320 5.790 ;
        RECT 15.040 5.720 15.300 5.790 ;
        RECT 15.840 5.720 16.020 5.850 ;
        RECT 13.150 5.580 13.320 5.620 ;
        RECT 11.570 5.180 11.740 5.500 ;
        RECT 12.140 5.400 12.340 5.570 ;
        RECT 12.170 5.300 12.340 5.400 ;
        RECT 13.710 5.540 14.580 5.710 ;
        RECT 15.040 5.540 16.020 5.720 ;
        RECT 3.980 4.830 4.220 4.850 ;
        RECT 4.790 4.840 4.960 4.930 ;
        RECT 6.490 4.920 6.820 5.090 ;
        RECT 9.640 5.080 9.810 5.180 ;
        RECT 9.620 4.910 9.810 5.080 ;
        RECT 9.640 4.850 9.810 4.910 ;
        RECT 10.060 5.120 10.230 5.180 ;
        RECT 10.060 4.850 10.310 5.120 ;
        RECT 10.800 4.930 11.050 5.180 ;
        RECT 10.070 4.830 10.310 4.850 ;
        RECT 10.880 4.840 11.050 4.930 ;
        RECT 11.530 4.930 11.740 5.180 ;
        RECT 13.710 5.100 13.880 5.540 ;
        RECT 15.040 5.100 15.300 5.540 ;
        RECT 15.840 5.430 16.020 5.540 ;
        RECT 12.250 4.930 13.880 5.100 ;
        RECT 14.330 4.930 15.300 5.100 ;
        RECT 15.750 4.930 16.090 5.100 ;
        RECT 11.530 4.850 11.700 4.930 ;
        RECT 13.020 4.890 13.190 4.930 ;
        RECT 3.980 4.220 4.150 4.360 ;
        RECT 10.070 4.220 10.240 4.360 ;
        RECT 10.800 4.240 10.970 4.320 ;
        RECT 11.610 4.240 11.780 4.320 ;
        RECT 13.150 4.280 13.320 4.400 ;
        RECT 3.980 4.050 4.170 4.220 ;
        RECT 3.980 3.950 4.150 4.050 ;
        RECT 3.550 3.570 3.720 3.670 ;
        RECT 3.530 3.400 3.720 3.570 ;
        RECT 3.550 3.340 3.720 3.400 ;
        RECT 3.970 3.610 4.140 3.670 ;
        RECT 3.970 3.340 4.220 3.610 ;
        RECT 4.710 3.590 4.960 3.670 ;
        RECT 4.710 3.420 6.010 3.590 ;
        RECT 6.570 3.580 6.740 4.210 ;
        RECT 10.070 4.050 10.260 4.220 ;
        RECT 10.070 3.950 10.240 4.050 ;
        RECT 10.800 3.670 11.010 4.240 ;
        RECT 11.570 3.990 11.780 4.240 ;
        RECT 12.170 4.060 12.340 4.160 ;
        RECT 13.110 4.110 13.320 4.280 ;
        RECT 15.040 4.210 15.300 4.280 ;
        RECT 15.840 4.210 16.020 4.340 ;
        RECT 13.150 4.070 13.320 4.110 ;
        RECT 11.570 3.670 11.740 3.990 ;
        RECT 12.140 3.890 12.340 4.060 ;
        RECT 12.170 3.790 12.340 3.890 ;
        RECT 13.710 4.030 14.580 4.200 ;
        RECT 15.040 4.030 16.020 4.210 ;
        RECT 3.980 3.320 4.220 3.340 ;
        RECT 4.790 3.330 4.960 3.420 ;
        RECT 6.490 3.410 6.820 3.580 ;
        RECT 9.640 3.570 9.810 3.670 ;
        RECT 9.620 3.400 9.810 3.570 ;
        RECT 9.640 3.340 9.810 3.400 ;
        RECT 10.060 3.610 10.230 3.670 ;
        RECT 10.060 3.340 10.310 3.610 ;
        RECT 10.800 3.420 11.050 3.670 ;
        RECT 10.070 3.320 10.310 3.340 ;
        RECT 10.880 3.330 11.050 3.420 ;
        RECT 11.530 3.420 11.740 3.670 ;
        RECT 13.710 3.590 13.880 4.030 ;
        RECT 15.040 3.590 15.300 4.030 ;
        RECT 15.840 3.920 16.020 4.030 ;
        RECT 12.250 3.420 13.880 3.590 ;
        RECT 14.330 3.420 15.300 3.590 ;
        RECT 15.750 3.420 16.090 3.590 ;
        RECT 11.530 3.340 11.700 3.420 ;
        RECT 13.020 3.380 13.190 3.420 ;
        RECT 3.980 2.710 4.150 2.850 ;
        RECT 10.070 2.710 10.240 2.850 ;
        RECT 10.800 2.730 10.970 2.810 ;
        RECT 11.610 2.730 11.780 2.810 ;
        RECT 13.150 2.770 13.320 2.890 ;
        RECT 3.980 2.540 4.170 2.710 ;
        RECT 3.980 2.440 4.150 2.540 ;
        RECT 3.550 2.060 3.720 2.160 ;
        RECT 3.530 1.890 3.720 2.060 ;
        RECT 3.550 1.830 3.720 1.890 ;
        RECT 3.970 2.100 4.140 2.160 ;
        RECT 3.970 1.830 4.220 2.100 ;
        RECT 4.710 2.080 4.960 2.160 ;
        RECT 4.710 1.910 6.010 2.080 ;
        RECT 6.570 2.070 6.740 2.700 ;
        RECT 10.070 2.540 10.260 2.710 ;
        RECT 10.070 2.440 10.240 2.540 ;
        RECT 10.800 2.160 11.010 2.730 ;
        RECT 11.570 2.480 11.780 2.730 ;
        RECT 12.170 2.550 12.340 2.650 ;
        RECT 13.110 2.600 13.320 2.770 ;
        RECT 15.040 2.700 15.300 2.770 ;
        RECT 15.840 2.700 16.020 2.830 ;
        RECT 13.150 2.560 13.320 2.600 ;
        RECT 11.570 2.160 11.740 2.480 ;
        RECT 12.140 2.380 12.340 2.550 ;
        RECT 12.170 2.280 12.340 2.380 ;
        RECT 13.710 2.520 14.580 2.690 ;
        RECT 15.040 2.520 16.020 2.700 ;
        RECT 3.980 1.810 4.220 1.830 ;
        RECT 4.790 1.820 4.960 1.910 ;
        RECT 6.490 1.900 6.820 2.070 ;
        RECT 9.640 2.060 9.810 2.160 ;
        RECT 9.620 1.890 9.810 2.060 ;
        RECT 9.640 1.830 9.810 1.890 ;
        RECT 10.060 2.100 10.230 2.160 ;
        RECT 10.060 1.830 10.310 2.100 ;
        RECT 10.800 1.910 11.050 2.160 ;
        RECT 10.070 1.810 10.310 1.830 ;
        RECT 10.880 1.820 11.050 1.910 ;
        RECT 11.530 1.910 11.740 2.160 ;
        RECT 13.710 2.080 13.880 2.520 ;
        RECT 15.040 2.080 15.300 2.520 ;
        RECT 15.840 2.410 16.020 2.520 ;
        RECT 12.250 1.910 13.880 2.080 ;
        RECT 14.330 1.910 15.300 2.080 ;
        RECT 15.750 1.910 16.090 2.080 ;
        RECT 11.530 1.830 11.700 1.910 ;
        RECT 13.020 1.870 13.190 1.910 ;
        RECT 10.070 1.210 10.240 1.350 ;
        RECT 10.800 1.230 10.970 1.310 ;
        RECT 11.610 1.230 11.780 1.310 ;
        RECT 13.150 1.270 13.320 1.390 ;
        RECT 10.070 1.040 10.260 1.210 ;
        RECT 10.070 0.940 10.240 1.040 ;
        RECT 10.800 0.660 11.010 1.230 ;
        RECT 11.570 0.980 11.780 1.230 ;
        RECT 12.170 1.050 12.340 1.150 ;
        RECT 13.110 1.100 13.320 1.270 ;
        RECT 15.040 1.200 15.300 1.270 ;
        RECT 15.840 1.200 16.020 1.330 ;
        RECT 13.150 1.060 13.320 1.100 ;
        RECT 11.570 0.660 11.740 0.980 ;
        RECT 12.140 0.880 12.340 1.050 ;
        RECT 12.170 0.780 12.340 0.880 ;
        RECT 13.710 1.020 14.580 1.190 ;
        RECT 15.040 1.020 16.020 1.200 ;
        RECT 9.640 0.560 9.810 0.660 ;
        RECT 9.620 0.390 9.810 0.560 ;
        RECT 9.640 0.330 9.810 0.390 ;
        RECT 10.060 0.600 10.230 0.660 ;
        RECT 10.060 0.330 10.310 0.600 ;
        RECT 10.800 0.410 11.050 0.660 ;
        RECT 10.070 0.310 10.310 0.330 ;
        RECT 10.880 0.320 11.050 0.410 ;
        RECT 11.530 0.410 11.740 0.660 ;
        RECT 13.710 0.580 13.880 1.020 ;
        RECT 15.040 0.580 15.300 1.020 ;
        RECT 15.840 0.910 16.020 1.020 ;
        RECT 12.250 0.410 13.880 0.580 ;
        RECT 14.330 0.410 15.300 0.580 ;
        RECT 15.750 0.410 16.090 0.580 ;
        RECT 11.530 0.330 11.700 0.410 ;
        RECT 13.020 0.370 13.190 0.410 ;
      LAYER mcon ;
        RECT 4.000 5.560 4.170 5.730 ;
        RECT 10.090 5.560 10.260 5.730 ;
        RECT 6.570 5.200 6.740 5.370 ;
        RECT 4.010 4.880 4.180 5.050 ;
        RECT 5.350 4.930 5.520 5.100 ;
        RECT 10.100 4.880 10.270 5.050 ;
        RECT 15.070 5.220 15.250 5.400 ;
        RECT 4.000 4.050 4.170 4.220 ;
        RECT 10.090 4.050 10.260 4.220 ;
        RECT 6.570 3.690 6.740 3.860 ;
        RECT 4.010 3.370 4.180 3.540 ;
        RECT 5.350 3.420 5.520 3.590 ;
        RECT 10.100 3.370 10.270 3.540 ;
        RECT 15.070 3.710 15.250 3.890 ;
        RECT 4.000 2.540 4.170 2.710 ;
        RECT 10.090 2.540 10.260 2.710 ;
        RECT 6.570 2.180 6.740 2.350 ;
        RECT 4.010 1.860 4.180 2.030 ;
        RECT 5.350 1.910 5.520 2.080 ;
        RECT 10.100 1.860 10.270 2.030 ;
        RECT 15.070 2.200 15.250 2.380 ;
        RECT 10.090 1.040 10.260 1.210 ;
        RECT 10.100 0.360 10.270 0.530 ;
        RECT 15.070 0.700 15.250 0.880 ;
      LAYER met1 ;
        RECT 3.670 7.210 3.940 7.500 ;
        RECT 3.630 6.940 3.960 7.210 ;
        RECT 3.670 6.160 3.940 6.940 ;
        RECT 3.660 5.830 3.940 6.160 ;
        RECT 4.130 6.120 4.400 6.600 ;
        RECT 3.670 5.800 3.940 5.830 ;
        RECT 3.440 4.840 3.750 5.190 ;
        RECT 3.440 3.330 3.750 3.680 ;
        RECT 3.970 2.980 4.400 6.120 ;
        RECT 4.590 5.610 4.860 7.070 ;
        RECT 5.540 6.570 5.830 6.620 ;
        RECT 5.520 6.220 5.830 6.570 ;
        RECT 4.540 5.340 4.870 5.610 ;
        RECT 4.590 4.030 4.860 5.340 ;
        RECT 5.540 5.140 5.830 6.220 ;
        RECT 10.060 5.780 10.280 6.120 ;
        RECT 10.060 5.520 10.290 5.780 ;
        RECT 5.270 5.130 5.830 5.140 ;
        RECT 4.570 3.700 4.860 4.030 ;
        RECT 4.590 3.680 4.860 3.700 ;
        RECT 5.060 4.880 5.830 5.130 ;
        RECT 5.060 4.740 5.340 4.880 ;
        RECT 5.060 3.630 5.330 4.740 ;
        RECT 5.540 3.630 5.830 4.880 ;
        RECT 9.530 4.840 9.840 5.190 ;
        RECT 10.060 5.120 10.280 5.520 ;
        RECT 12.080 5.360 12.410 5.620 ;
        RECT 13.050 5.580 13.480 5.870 ;
        RECT 10.060 4.810 10.310 5.120 ;
        RECT 12.920 4.830 13.310 5.100 ;
        RECT 10.060 4.270 10.280 4.810 ;
        RECT 10.060 4.010 10.290 4.270 ;
        RECT 5.060 3.570 5.830 3.630 ;
        RECT 5.060 3.370 5.840 3.570 ;
        RECT 3.970 2.650 4.430 2.980 ;
        RECT 3.970 2.600 4.400 2.650 ;
        RECT 3.970 2.500 4.200 2.600 ;
        RECT 5.060 2.530 5.330 3.370 ;
        RECT 3.440 1.820 3.750 2.170 ;
        RECT 3.970 2.100 4.190 2.500 ;
        RECT 5.040 2.200 5.330 2.530 ;
        RECT 5.060 2.170 5.330 2.200 ;
        RECT 5.540 3.220 5.840 3.370 ;
        RECT 9.530 3.330 9.840 3.680 ;
        RECT 10.060 3.610 10.280 4.010 ;
        RECT 12.080 3.850 12.410 4.110 ;
        RECT 13.050 4.070 13.480 4.360 ;
        RECT 10.060 3.300 10.310 3.610 ;
        RECT 12.920 3.320 13.310 3.590 ;
        RECT 5.540 2.120 5.830 3.220 ;
        RECT 10.060 2.760 10.280 3.300 ;
        RECT 10.060 2.500 10.290 2.760 ;
        RECT 3.970 1.790 4.220 2.100 ;
        RECT 5.270 1.860 5.830 2.120 ;
        RECT 3.970 1.590 4.190 1.790 ;
        RECT 5.540 1.680 5.830 1.860 ;
        RECT 9.530 1.820 9.840 2.170 ;
        RECT 10.060 2.100 10.280 2.500 ;
        RECT 12.080 2.340 12.410 2.600 ;
        RECT 13.050 2.560 13.480 2.850 ;
        RECT 10.060 1.790 10.310 2.100 ;
        RECT 12.920 1.810 13.310 2.080 ;
        RECT 10.060 1.260 10.280 1.790 ;
        RECT 10.060 1.000 10.290 1.260 ;
        RECT 9.530 0.320 9.840 0.670 ;
        RECT 10.060 0.600 10.280 1.000 ;
        RECT 12.080 0.840 12.410 1.100 ;
        RECT 13.050 1.060 13.480 1.350 ;
        RECT 10.060 0.290 10.310 0.600 ;
        RECT 12.920 0.310 13.310 0.580 ;
        RECT 10.060 0.090 10.280 0.290 ;
        RECT 15.030 0.090 15.300 6.130 ;
        RECT 15.850 4.840 16.160 5.160 ;
        RECT 15.850 3.330 16.160 3.650 ;
        RECT 15.850 1.820 16.160 2.140 ;
        RECT 15.850 0.320 16.160 0.640 ;
      LAYER via ;
        RECT 3.660 6.940 3.930 7.210 ;
        RECT 4.590 6.750 4.860 7.020 ;
        RECT 3.660 5.860 3.930 6.130 ;
        RECT 4.130 6.260 4.400 6.530 ;
        RECT 3.470 4.870 3.730 5.130 ;
        RECT 5.520 6.250 5.810 6.540 ;
        RECT 4.570 5.340 4.840 5.610 ;
        RECT 4.120 4.180 4.390 4.450 ;
        RECT 3.470 3.360 3.730 3.620 ;
        RECT 4.570 3.730 4.840 4.000 ;
        RECT 5.300 5.040 5.560 5.140 ;
        RECT 5.070 5.000 5.560 5.040 ;
        RECT 5.070 4.880 5.820 5.000 ;
        RECT 5.070 4.770 5.340 4.880 ;
        RECT 5.560 4.740 5.820 4.880 ;
        RECT 9.560 4.870 9.820 5.130 ;
        RECT 12.120 5.360 12.380 5.620 ;
        RECT 13.110 5.610 13.370 5.870 ;
        RECT 12.980 4.830 13.240 5.090 ;
        RECT 5.300 3.540 5.560 3.630 ;
        RECT 5.300 3.370 5.840 3.540 ;
        RECT 4.160 2.680 4.430 2.950 ;
        RECT 3.470 1.850 3.730 2.110 ;
        RECT 5.040 2.230 5.310 2.500 ;
        RECT 5.550 3.250 5.840 3.370 ;
        RECT 9.560 3.360 9.820 3.620 ;
        RECT 12.120 3.850 12.380 4.110 ;
        RECT 13.110 4.100 13.370 4.360 ;
        RECT 12.980 3.320 13.240 3.580 ;
        RECT 5.300 2.000 5.560 2.120 ;
        RECT 5.300 1.860 5.830 2.000 ;
        RECT 5.540 1.710 5.830 1.860 ;
        RECT 9.560 1.850 9.820 2.110 ;
        RECT 12.120 2.340 12.380 2.600 ;
        RECT 13.110 2.590 13.370 2.850 ;
        RECT 12.980 1.810 13.240 2.070 ;
        RECT 9.560 0.350 9.820 0.610 ;
        RECT 12.120 0.840 12.380 1.100 ;
        RECT 13.110 1.090 13.370 1.350 ;
        RECT 12.980 0.310 13.240 0.570 ;
        RECT 15.880 4.870 16.140 5.130 ;
        RECT 15.880 3.360 16.140 3.620 ;
        RECT 15.880 1.850 16.140 2.110 ;
        RECT 15.880 0.350 16.140 0.610 ;
      LAYER met2 ;
        RECT 3.710 7.400 6.080 7.410 ;
        RECT 3.690 7.250 6.080 7.400 ;
        RECT 3.690 7.240 3.960 7.250 ;
        RECT 3.660 7.170 3.960 7.240 ;
        RECT 3.430 6.990 3.960 7.170 ;
        RECT 3.660 6.910 3.930 6.990 ;
        RECT 4.560 6.960 4.890 7.020 ;
        RECT 4.560 6.800 6.080 6.960 ;
        RECT 4.560 6.750 4.890 6.800 ;
        RECT 4.100 6.500 4.430 6.530 ;
        RECT 3.430 6.320 4.450 6.500 ;
        RECT 4.100 6.310 4.450 6.320 ;
        RECT 5.490 6.470 5.840 6.540 ;
        RECT 5.490 6.310 6.080 6.470 ;
        RECT 4.100 6.260 4.430 6.310 ;
        RECT 5.490 6.250 5.840 6.310 ;
        RECT 3.630 6.070 3.960 6.130 ;
        RECT 3.630 5.910 5.270 6.070 ;
        RECT 3.630 5.860 3.960 5.910 ;
        RECT 5.110 5.900 5.270 5.910 ;
        RECT 5.110 5.740 6.070 5.900 ;
        RECT 9.440 5.810 13.480 5.970 ;
        RECT 3.360 5.550 6.970 5.730 ;
        RECT 3.430 5.480 4.840 5.550 ;
        RECT 12.080 5.540 12.410 5.620 ;
        RECT 13.060 5.580 13.480 5.810 ;
        RECT 11.810 5.520 12.410 5.540 ;
        RECT 4.570 5.450 4.840 5.480 ;
        RECT 4.570 5.310 4.850 5.450 ;
        RECT 4.620 5.290 4.850 5.310 ;
        RECT 5.120 5.290 6.080 5.450 ;
        RECT 9.450 5.360 12.410 5.520 ;
        RECT 5.120 5.140 5.280 5.290 ;
        RECT 3.440 5.030 3.760 5.130 ;
        RECT 5.120 5.060 5.590 5.140 ;
        RECT 5.120 5.040 6.970 5.060 ;
        RECT 3.430 4.990 3.760 5.030 ;
        RECT 5.040 4.990 6.970 5.040 ;
        RECT 9.530 5.030 9.850 5.130 ;
        RECT 3.430 4.880 6.970 4.990 ;
        RECT 3.430 4.810 5.370 4.880 ;
        RECT 5.040 4.770 5.370 4.810 ;
        RECT 5.530 4.800 6.080 4.880 ;
        RECT 9.450 4.870 9.850 5.030 ;
        RECT 5.530 4.740 5.850 4.800 ;
        RECT 4.090 4.390 4.420 4.450 ;
        RECT 4.090 4.230 6.080 4.390 ;
        RECT 9.440 4.300 13.480 4.460 ;
        RECT 4.090 4.220 4.420 4.230 ;
        RECT 3.360 4.040 6.970 4.220 ;
        RECT 12.080 4.030 12.410 4.110 ;
        RECT 13.060 4.070 13.480 4.300 ;
        RECT 11.810 4.010 12.410 4.030 ;
        RECT 4.540 3.940 4.870 4.000 ;
        RECT 4.540 3.780 6.080 3.940 ;
        RECT 9.450 3.850 12.410 4.010 ;
        RECT 4.540 3.730 4.870 3.780 ;
        RECT 3.440 3.520 3.760 3.620 ;
        RECT 3.430 3.480 3.760 3.520 ;
        RECT 5.270 3.550 5.590 3.630 ;
        RECT 5.270 3.480 6.970 3.550 ;
        RECT 9.530 3.520 9.850 3.620 ;
        RECT 3.430 3.370 6.970 3.480 ;
        RECT 3.430 3.300 6.080 3.370 ;
        RECT 9.450 3.360 9.850 3.520 ;
        RECT 5.520 3.290 6.080 3.300 ;
        RECT 5.520 3.250 5.870 3.290 ;
        RECT 4.130 2.890 4.460 2.950 ;
        RECT 4.130 2.730 6.080 2.890 ;
        RECT 9.440 2.790 13.480 2.950 ;
        RECT 4.130 2.710 4.460 2.730 ;
        RECT 3.360 2.530 6.970 2.710 ;
        RECT 12.080 2.520 12.410 2.600 ;
        RECT 13.060 2.560 13.480 2.790 ;
        RECT 11.810 2.500 12.410 2.520 ;
        RECT 5.010 2.440 5.340 2.500 ;
        RECT 5.010 2.280 6.080 2.440 ;
        RECT 9.450 2.340 12.410 2.500 ;
        RECT 5.010 2.230 5.340 2.280 ;
        RECT 3.440 2.010 3.760 2.110 ;
        RECT 3.430 1.850 3.760 2.010 ;
        RECT 5.270 2.040 5.590 2.120 ;
        RECT 5.270 1.860 6.970 2.040 ;
        RECT 9.530 2.010 9.850 2.110 ;
        RECT 5.510 1.790 6.080 1.860 ;
        RECT 9.450 1.850 9.850 2.010 ;
        RECT 5.510 1.710 5.860 1.790 ;
        RECT 9.440 1.290 13.480 1.450 ;
        RECT 12.080 1.020 12.410 1.100 ;
        RECT 13.060 1.060 13.480 1.290 ;
        RECT 11.810 1.000 12.410 1.020 ;
        RECT 9.450 0.840 12.410 1.000 ;
        RECT 9.530 0.510 9.850 0.610 ;
        RECT 9.450 0.350 9.850 0.510 ;
        RECT 12.940 0.490 13.310 0.570 ;
        RECT 12.940 0.480 13.970 0.490 ;
        RECT 15.850 0.480 16.160 0.640 ;
        RECT 12.940 0.310 16.320 0.480 ;
  END
END sky130_hilas_VinjDecode2to4

MACRO sky130_hilas_TA2Cell_1FG
  CLASS CORE ;
  FOREIGN sky130_hilas_TA2Cell_1FG ;
  ORIGIN 0.000 0.000 ;
  SIZE 32.050 BY 9.870 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 12.810 1.250 13.290 1.260 ;
        RECT 12.810 1.010 13.700 1.250 ;
    END
  END VIN12
  PIN VIN11
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 12.860 4.770 13.700 4.970 ;
    END
  END VIN11
  PIN VIN21
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT 27.920 3.350 28.230 3.390 ;
        RECT 27.600 3.340 28.260 3.350 ;
        RECT 27.600 3.110 28.700 3.340 ;
        RECT 27.920 3.060 28.230 3.110 ;
    END
  END VIN21
  PIN VIN22
    USE ANALOG ;
    ANTENNAGATEAREA 4.342100 ;
    ANTENNADIFFAREA 8.158800 ;
    PORT
      LAYER nwell ;
        RECT 27.570 6.050 30.880 9.870 ;
        RECT 26.920 6.040 32.050 6.050 ;
        RECT 26.910 3.830 32.050 6.040 ;
        RECT 26.910 0.000 28.770 3.830 ;
        RECT 30.770 0.000 32.050 3.830 ;
      LAYER met2 ;
        RECT 29.490 7.010 29.810 7.270 ;
        RECT 29.530 6.990 30.710 7.010 ;
        RECT 29.530 6.730 30.750 6.990 ;
        RECT 29.530 6.670 30.710 6.730 ;
        RECT 29.490 6.660 30.710 6.670 ;
        RECT 29.490 6.410 29.810 6.660 ;
        RECT 28.160 6.030 28.470 6.040 ;
        RECT 27.590 6.020 28.470 6.030 ;
        RECT 27.520 5.780 28.470 6.020 ;
        RECT 28.160 5.710 28.470 5.780 ;
        RECT 29.130 5.710 29.440 5.760 ;
        RECT 31.380 5.710 31.690 5.810 ;
        RECT 28.550 5.590 28.860 5.660 ;
        RECT 29.130 5.590 31.690 5.710 ;
        RECT 28.550 5.480 31.690 5.590 ;
        RECT 28.550 5.380 30.880 5.480 ;
        RECT 28.550 5.330 28.860 5.380 ;
        RECT 28.310 5.170 28.620 5.210 ;
        RECT 28.130 5.030 28.850 5.170 ;
        RECT 29.080 5.030 29.390 5.110 ;
        RECT 28.130 4.920 29.390 5.030 ;
        RECT 28.310 4.880 29.390 4.920 ;
        RECT 28.580 4.820 29.390 4.880 ;
        RECT 28.580 4.810 28.850 4.820 ;
        RECT 29.080 4.780 29.390 4.820 ;
        RECT 27.190 4.530 27.500 4.670 ;
        RECT 13.310 4.490 23.450 4.520 ;
        RECT 26.840 4.490 27.500 4.530 ;
        RECT 28.400 4.500 28.710 4.640 ;
        RECT 28.400 4.490 30.880 4.500 ;
        RECT 13.310 4.340 30.880 4.490 ;
        RECT 13.310 4.300 23.450 4.340 ;
        RECT 26.840 4.310 27.190 4.340 ;
        RECT 28.400 4.320 30.880 4.340 ;
        RECT 28.400 4.310 28.710 4.320 ;
        RECT 23.230 3.100 23.450 4.300 ;
        RECT 28.650 4.240 28.850 4.250 ;
        RECT 28.650 4.230 28.870 4.240 ;
        RECT 29.080 4.230 29.390 4.270 ;
        RECT 28.650 4.160 29.390 4.230 ;
        RECT 28.360 4.140 29.390 4.160 ;
        RECT 28.310 4.020 29.390 4.140 ;
        RECT 28.310 3.900 28.870 4.020 ;
        RECT 29.080 3.940 29.390 4.020 ;
        RECT 28.310 3.890 28.780 3.900 ;
        RECT 23.200 3.060 23.450 3.100 ;
        RECT 23.200 2.420 23.460 3.060 ;
        RECT 23.200 2.210 27.330 2.420 ;
        RECT 27.120 2.070 27.330 2.210 ;
        RECT 29.080 2.070 29.390 2.150 ;
        RECT 27.120 1.860 29.390 2.070 ;
        RECT 29.080 1.820 29.390 1.860 ;
        RECT 18.140 0.350 18.460 0.360 ;
        RECT 28.580 0.350 28.910 0.490 ;
        RECT 18.140 0.190 28.910 0.350 ;
        RECT 18.140 0.180 18.830 0.190 ;
        RECT 18.140 0.060 18.460 0.180 ;
    END
  END VIN22
  PIN VPWR
    USE ANALOG ;
    ANTENNADIFFAREA 1.373600 ;
    PORT
      LAYER met1 ;
        RECT 30.750 5.900 31.030 6.050 ;
        RECT 30.760 4.470 31.030 5.900 ;
        RECT 30.760 4.180 31.040 4.470 ;
        RECT 30.760 1.880 31.030 4.180 ;
        RECT 30.760 1.590 31.040 1.880 ;
        RECT 30.760 0.000 31.030 1.590 ;
    END
  END VPWR
  PIN VGND
    USE ANALOG ;
    ANTENNAGATEAREA 3.745100 ;
    ANTENNADIFFAREA 3.678400 ;
    PORT
      LAYER met1 ;
        RECT 29.920 8.410 30.110 9.870 ;
        RECT 30.360 9.220 30.640 9.870 ;
        RECT 30.250 8.620 30.640 9.220 ;
        RECT 29.920 8.380 30.140 8.410 ;
        RECT 29.900 8.110 30.150 8.380 ;
        RECT 29.910 8.100 30.150 8.110 ;
        RECT 29.910 7.860 30.140 8.100 ;
        RECT 29.520 6.380 29.780 6.700 ;
        RECT 29.520 6.260 29.760 6.380 ;
        RECT 29.950 6.050 30.110 7.860 ;
        RECT 30.360 7.020 30.640 8.620 ;
        RECT 30.360 6.700 30.720 7.020 ;
        RECT 30.360 6.050 30.640 6.700 ;
        RECT 28.150 5.710 28.470 6.030 ;
        RECT 29.950 5.830 30.640 6.050 ;
        RECT 29.130 5.430 29.450 5.750 ;
        RECT 29.910 5.580 30.640 5.830 ;
        RECT 29.900 5.310 30.640 5.580 ;
        RECT 29.080 4.780 29.400 5.100 ;
        RECT 28.400 4.200 28.710 4.640 ;
        RECT 28.410 4.190 28.620 4.200 ;
        RECT 28.390 3.870 28.650 4.190 ;
        RECT 29.080 3.950 29.400 4.270 ;
        RECT 28.410 2.580 28.620 3.870 ;
        RECT 29.920 3.820 30.640 5.310 ;
        RECT 28.390 2.290 28.620 2.580 ;
        RECT 28.580 0.200 28.910 0.490 ;
        RECT 30.090 0.200 30.430 3.820 ;
        RECT 28.570 0.060 30.430 0.200 ;
        RECT 30.090 0.000 30.430 0.060 ;
      LAYER via ;
        RECT 29.520 6.410 29.780 6.670 ;
        RECT 30.460 6.730 30.720 6.990 ;
        RECT 28.180 5.740 28.440 6.000 ;
        RECT 29.160 5.460 29.420 5.720 ;
        RECT 29.110 4.810 29.370 5.070 ;
        RECT 28.430 4.350 28.690 4.610 ;
        RECT 28.390 3.900 28.650 4.160 ;
        RECT 29.110 3.980 29.370 4.240 ;
        RECT 28.610 0.210 28.880 0.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 12.430 5.960 12.660 6.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 18.220 5.960 18.450 6.050 ;
    END
  END VGND
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 4.200 5.880 4.520 6.000 ;
        RECT 26.400 5.880 26.720 6.000 ;
        RECT 4.200 5.700 26.720 5.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 26.400 0.000 26.680 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.200 6.000 4.480 6.050 ;
        RECT 4.200 5.720 4.520 6.000 ;
      LAYER via ;
        RECT 4.230 5.730 4.490 5.990 ;
    END
  END VINJ
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER met2 ;
        RECT 29.130 3.570 29.440 3.620 ;
        RECT 31.430 3.570 31.740 3.590 ;
        RECT 29.130 3.340 32.050 3.570 ;
        RECT 29.130 3.290 29.440 3.340 ;
        RECT 31.430 3.260 31.740 3.340 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.305700 ;
    PORT
      LAYER met2 ;
        RECT 29.130 2.740 29.440 2.800 ;
        RECT 31.420 2.740 31.730 2.870 ;
        RECT 29.130 2.520 32.050 2.740 ;
        RECT 29.130 2.470 29.440 2.520 ;
    END
  END OUTPUT2
  PIN DRAIN1
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 2.020 5.590 2.330 5.660 ;
        RECT 0.000 5.380 11.530 5.590 ;
        RECT 1.310 5.370 11.530 5.380 ;
        RECT 2.020 5.330 2.330 5.370 ;
    END
  END DRAIN1
  PIN DRAIN2
    PORT
      LAYER met2 ;
        RECT 3.960 0.500 4.040 0.680 ;
    END
  END DRAIN2
  PIN COLSEL2
    PORT
      LAYER met1 ;
        RECT 4.730 5.990 4.920 6.050 ;
    END
  END COLSEL2
  PIN GATE2
    PORT
      LAYER met1 ;
        RECT 11.210 5.960 11.440 6.040 ;
    END
  END GATE2
  PIN GATE1
    PORT
      LAYER met1 ;
        RECT 19.440 5.970 19.670 6.050 ;
    END
  END GATE1
  PIN COLSEL1
    PORT
      LAYER met1 ;
        RECT 25.960 5.970 26.150 6.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.960 0.000 26.150 0.050 ;
    END
  END COLSEL1
  PIN VTUN
    PORT
      LAYER met1 ;
        RECT 14.720 5.890 16.160 6.050 ;
    END
  END VTUN
  OBS
      LAYER nwell ;
        RECT 0.000 3.830 3.310 9.860 ;
        RECT 5.040 7.480 7.760 9.130 ;
        RECT 9.790 9.120 11.520 9.870 ;
        RECT 5.050 7.440 7.760 7.480 ;
        RECT 5.050 6.110 7.760 6.150 ;
        RECT 5.040 6.050 7.760 6.110 ;
        RECT 3.960 6.040 7.760 6.050 ;
        RECT 3.960 5.370 4.030 5.550 ;
        RECT 5.040 4.460 7.760 6.040 ;
        RECT 9.780 5.550 11.520 9.120 ;
        RECT 9.790 3.830 11.520 5.550 ;
        RECT 19.360 9.120 21.090 9.870 ;
        RECT 19.360 5.550 21.100 9.120 ;
        RECT 23.120 7.480 25.840 9.130 ;
        RECT 23.120 7.440 25.830 7.480 ;
        RECT 23.120 6.110 25.830 6.150 ;
        RECT 19.360 3.830 21.090 5.550 ;
        RECT 23.120 4.460 25.840 6.110 ;
        RECT 3.960 0.500 4.040 0.680 ;
      LAYER li1 ;
        RECT 0.400 9.190 0.600 9.540 ;
        RECT 1.880 9.290 2.410 9.460 ;
        RECT 0.390 9.160 0.600 9.190 ;
        RECT 0.390 8.580 0.610 9.160 ;
        RECT 0.390 8.570 0.600 8.580 ;
        RECT 0.770 8.400 0.960 8.410 ;
        RECT 0.760 8.110 0.960 8.400 ;
        RECT 0.730 7.780 0.970 8.110 ;
        RECT 1.160 7.300 1.330 8.910 ;
        RECT 1.150 7.110 1.330 7.300 ;
        RECT 1.990 8.380 2.160 8.900 ;
        RECT 2.580 8.710 2.910 8.880 ;
        RECT 3.930 8.710 4.280 8.880 ;
        RECT 4.600 8.860 9.660 9.690 ;
        RECT 28.470 9.290 29.000 9.460 ;
        RECT 30.280 9.190 30.480 9.540 ;
        RECT 30.280 9.160 30.490 9.190 ;
        RECT 9.110 8.780 9.590 8.860 ;
        RECT 1.990 8.120 2.320 8.380 ;
        RECT 1.990 7.210 2.160 8.120 ;
        RECT 2.580 7.920 2.910 8.090 ;
        RECT 3.930 7.920 4.280 8.090 ;
        RECT 7.230 7.920 7.460 8.610 ;
        RECT 9.110 8.530 9.580 8.780 ;
        RECT 26.600 8.710 26.950 8.880 ;
        RECT 27.970 8.710 28.300 8.880 ;
        RECT 10.540 7.730 11.090 8.160 ;
        RECT 19.790 7.730 20.340 8.160 ;
        RECT 23.420 7.920 23.650 8.610 ;
        RECT 28.720 8.380 28.890 8.900 ;
        RECT 28.560 8.120 28.890 8.380 ;
        RECT 26.600 7.920 26.950 8.090 ;
        RECT 27.970 7.920 28.300 8.090 ;
        RECT 2.580 7.130 2.910 7.300 ;
        RECT 3.930 7.130 4.270 7.300 ;
        RECT 1.150 6.390 1.330 6.580 ;
        RECT 2.660 6.560 2.830 7.130 ;
        RECT 8.300 6.900 8.490 7.300 ;
        RECT 22.390 6.900 22.580 7.300 ;
        RECT 26.610 7.130 26.950 7.300 ;
        RECT 27.970 7.130 28.300 7.300 ;
        RECT 28.720 7.210 28.890 8.120 ;
        RECT 29.550 7.300 29.720 8.910 ;
        RECT 30.270 8.580 30.490 9.160 ;
        RECT 30.280 8.570 30.490 8.580 ;
        RECT 29.920 8.400 30.110 8.410 ;
        RECT 29.920 8.110 30.120 8.400 ;
        RECT 29.910 7.780 30.150 8.110 ;
        RECT 8.300 6.890 8.680 6.900 ;
        RECT 4.940 6.710 8.680 6.890 ;
        RECT 8.300 6.670 8.680 6.710 ;
        RECT 22.200 6.890 22.580 6.900 ;
        RECT 22.200 6.710 25.940 6.890 ;
        RECT 22.200 6.670 22.580 6.710 ;
        RECT 0.730 5.580 0.970 5.910 ;
        RECT 0.760 5.290 0.960 5.580 ;
        RECT 0.770 5.280 0.960 5.290 ;
        RECT 0.390 5.110 0.600 5.120 ;
        RECT 0.390 4.530 0.610 5.110 ;
        RECT 1.160 4.780 1.330 6.390 ;
        RECT 1.990 5.620 2.160 6.480 ;
        RECT 2.580 6.390 2.910 6.560 ;
        RECT 3.930 6.390 4.270 6.560 ;
        RECT 8.300 6.290 8.490 6.670 ;
        RECT 10.540 6.000 11.090 6.430 ;
        RECT 19.790 6.000 20.340 6.430 ;
        RECT 22.390 6.290 22.580 6.670 ;
        RECT 28.050 6.560 28.220 7.130 ;
        RECT 29.550 7.110 29.730 7.300 ;
        RECT 26.610 6.390 26.950 6.560 ;
        RECT 27.970 6.390 28.300 6.560 ;
        RECT 27.900 6.000 28.070 6.050 ;
        RECT 1.990 5.360 2.320 5.620 ;
        RECT 2.580 5.600 2.910 5.770 ;
        RECT 3.930 5.600 4.280 5.770 ;
        RECT 1.990 4.790 2.160 5.360 ;
        RECT 7.230 4.980 7.460 5.710 ;
        RECT 2.580 4.810 2.910 4.980 ;
        RECT 3.930 4.810 4.280 4.980 ;
        RECT 9.270 4.850 9.610 5.100 ;
        RECT 23.420 4.980 23.650 5.710 ;
        RECT 26.600 5.600 26.950 5.770 ;
        RECT 27.900 5.740 28.460 6.000 ;
        RECT 27.900 5.720 28.300 5.740 ;
        RECT 27.970 5.600 28.300 5.720 ;
        RECT 28.720 5.620 28.890 6.480 ;
        RECT 29.550 6.390 29.730 6.580 ;
        RECT 29.550 5.760 29.720 6.390 ;
        RECT 29.370 5.720 29.720 5.760 ;
        RECT 9.270 4.770 9.620 4.850 ;
        RECT 26.600 4.810 26.950 4.980 ;
        RECT 0.390 4.500 0.600 4.530 ;
        RECT 0.400 4.150 0.600 4.500 ;
        RECT 1.880 4.230 2.410 4.400 ;
        RECT 4.570 3.920 9.620 4.770 ;
        RECT 27.320 4.640 27.500 5.570 ;
        RECT 28.050 5.310 28.380 5.480 ;
        RECT 28.560 5.360 28.890 5.620 ;
        RECT 29.140 5.460 29.720 5.720 ;
        RECT 29.910 5.760 30.150 5.910 ;
        RECT 29.910 5.580 30.510 5.760 ;
        RECT 29.370 5.430 29.720 5.460 ;
        RECT 28.130 5.170 28.380 5.310 ;
        RECT 28.130 4.980 28.610 5.170 ;
        RECT 27.970 4.910 28.610 4.980 ;
        RECT 27.970 4.810 28.300 4.910 ;
        RECT 27.200 4.610 27.520 4.640 ;
        RECT 27.200 4.420 27.530 4.610 ;
        RECT 27.200 4.380 27.520 4.420 ;
        RECT 12.450 2.470 12.650 3.480 ;
        RECT 18.200 2.470 18.490 3.480 ;
        RECT 27.320 0.470 27.500 4.380 ;
        RECT 28.130 3.530 28.300 4.810 ;
        RECT 28.720 4.790 28.890 5.360 ;
        RECT 28.960 5.070 29.130 5.110 ;
        RECT 29.550 5.100 29.720 5.430 ;
        RECT 29.920 5.280 30.510 5.580 ;
        RECT 31.330 5.640 31.910 5.810 ;
        RECT 31.330 5.540 31.720 5.640 ;
        RECT 31.330 5.510 31.710 5.540 ;
        RECT 31.330 5.360 31.690 5.510 ;
        RECT 29.370 5.070 29.720 5.100 ;
        RECT 28.960 4.810 29.720 5.070 ;
        RECT 28.960 4.780 29.130 4.810 ;
        RECT 29.370 4.780 29.720 4.810 ;
        RECT 29.370 4.770 29.570 4.780 ;
        RECT 29.960 4.770 30.510 5.280 ;
        RECT 30.980 5.190 31.690 5.360 ;
        RECT 30.270 4.530 30.490 4.770 ;
        RECT 30.280 4.500 30.490 4.530 ;
        RECT 28.470 4.270 29.000 4.400 ;
        RECT 30.280 4.280 30.480 4.500 ;
        RECT 30.980 4.440 31.680 4.750 ;
        RECT 28.470 4.240 29.130 4.270 ;
        RECT 29.370 4.240 29.570 4.280 ;
        RECT 28.470 4.230 29.570 4.240 ;
        RECT 28.960 3.980 29.570 4.230 ;
        RECT 28.960 3.940 29.130 3.980 ;
        RECT 29.370 3.950 29.570 3.980 ;
        RECT 29.370 3.590 29.570 3.620 ;
        RECT 27.930 3.330 28.250 3.360 ;
        RECT 29.140 3.330 29.570 3.590 ;
        RECT 27.930 3.140 28.260 3.330 ;
        RECT 29.370 3.290 29.570 3.330 ;
        RECT 29.960 3.290 30.510 4.280 ;
        RECT 30.830 4.210 31.680 4.440 ;
        RECT 30.980 3.870 31.680 4.210 ;
        RECT 31.440 3.510 31.760 3.550 ;
        RECT 31.440 3.450 31.770 3.510 ;
        RECT 30.970 3.320 31.770 3.450 ;
        RECT 30.970 3.290 31.760 3.320 ;
        RECT 30.970 3.270 31.670 3.290 ;
        RECT 27.930 3.100 28.250 3.140 ;
        RECT 27.930 3.020 28.100 3.100 ;
        RECT 27.880 2.850 28.100 3.020 ;
        RECT 27.880 2.690 28.050 2.850 ;
        RECT 29.370 2.760 29.570 2.800 ;
        RECT 28.410 2.430 28.600 2.550 ;
        RECT 29.140 2.500 29.570 2.760 ;
        RECT 29.370 2.470 29.570 2.500 ;
        RECT 28.050 2.320 28.600 2.430 ;
        RECT 28.050 2.260 28.590 2.320 ;
        RECT 28.130 0.480 28.300 2.260 ;
        RECT 28.960 2.110 29.130 2.150 ;
        RECT 29.370 2.110 29.570 2.140 ;
        RECT 28.960 1.850 29.570 2.110 ;
        RECT 28.960 1.820 29.130 1.850 ;
        RECT 29.370 1.810 29.570 1.850 ;
        RECT 29.960 1.810 30.510 2.800 ;
        RECT 31.430 2.790 31.750 2.830 ;
        RECT 30.970 2.610 31.760 2.790 ;
        RECT 31.430 2.600 31.760 2.610 ;
        RECT 31.430 2.570 31.750 2.600 ;
        RECT 30.980 1.850 31.680 2.190 ;
        RECT 30.830 1.620 31.680 1.850 ;
        RECT 28.960 1.280 29.130 1.310 ;
        RECT 29.370 1.280 29.570 1.320 ;
        RECT 28.960 1.020 29.570 1.280 ;
        RECT 28.960 0.980 29.130 1.020 ;
        RECT 29.370 0.990 29.570 1.020 ;
        RECT 29.370 0.630 29.570 0.660 ;
        RECT 29.140 0.370 29.570 0.630 ;
        RECT 29.370 0.330 29.570 0.370 ;
        RECT 29.960 0.330 30.510 1.320 ;
        RECT 30.980 1.310 31.680 1.620 ;
        RECT 30.980 0.700 31.690 0.870 ;
        RECT 31.330 0.420 31.690 0.700 ;
        RECT 31.330 0.250 31.910 0.420 ;
      LAYER mcon ;
        RECT 2.230 9.290 2.410 9.460 ;
        RECT 0.420 8.990 0.590 9.160 ;
        RECT 0.770 8.150 0.950 8.340 ;
        RECT 30.290 8.990 30.460 9.160 ;
        RECT 7.260 8.410 7.430 8.580 ;
        RECT 9.350 8.570 9.520 8.740 ;
        RECT 2.090 8.160 2.260 8.330 ;
        RECT 23.450 8.410 23.620 8.580 ;
        RECT 7.260 7.960 7.430 8.130 ;
        RECT 10.820 7.810 11.090 8.080 ;
        RECT 19.790 7.810 20.060 8.080 ;
        RECT 23.450 7.960 23.620 8.130 ;
        RECT 28.620 8.160 28.790 8.330 ;
        RECT 29.930 8.150 30.110 8.340 ;
        RECT 8.500 6.700 8.670 6.870 ;
        RECT 22.210 6.700 22.380 6.870 ;
        RECT 0.770 5.350 0.950 5.540 ;
        RECT 10.820 6.080 11.090 6.350 ;
        RECT 19.790 6.080 20.060 6.350 ;
        RECT 28.230 5.780 28.400 5.950 ;
        RECT 2.090 5.400 2.260 5.570 ;
        RECT 7.260 5.460 7.430 5.630 ;
        RECT 7.260 5.010 7.430 5.180 ;
        RECT 23.450 5.460 23.620 5.630 ;
        RECT 9.380 4.880 9.550 5.050 ;
        RECT 23.450 5.010 23.620 5.180 ;
        RECT 0.420 4.530 0.590 4.700 ;
        RECT 2.230 4.230 2.410 4.400 ;
        RECT 28.620 5.400 28.790 5.570 ;
        RECT 29.200 5.500 29.370 5.670 ;
        RECT 28.380 4.950 28.550 5.120 ;
        RECT 27.260 4.430 27.430 4.600 ;
        RECT 12.460 3.230 12.630 3.400 ;
        RECT 12.470 2.540 12.640 2.710 ;
        RECT 18.250 3.230 18.420 3.400 ;
        RECT 18.250 2.550 18.420 2.720 ;
        RECT 29.930 5.350 30.110 5.540 ;
        RECT 31.450 5.550 31.620 5.720 ;
        RECT 29.150 4.850 29.320 5.020 ;
        RECT 30.180 5.180 30.350 5.350 ;
        RECT 30.290 4.530 30.460 4.700 ;
        RECT 29.150 4.030 29.320 4.200 ;
        RECT 30.840 4.240 31.010 4.410 ;
        RECT 30.180 3.700 30.350 3.870 ;
        RECT 29.200 3.380 29.370 3.550 ;
        RECT 27.990 3.150 28.160 3.320 ;
        RECT 31.500 3.330 31.670 3.500 ;
        RECT 28.420 2.350 28.590 2.520 ;
        RECT 29.200 2.540 29.370 2.710 ;
        RECT 31.490 2.610 31.660 2.780 ;
        RECT 30.180 2.220 30.350 2.390 ;
        RECT 29.150 1.890 29.320 2.060 ;
        RECT 30.840 1.650 31.010 1.820 ;
        RECT 29.150 1.070 29.320 1.240 ;
        RECT 30.180 0.740 30.350 0.910 ;
        RECT 29.200 0.420 29.370 0.590 ;
        RECT 31.410 0.360 31.580 0.530 ;
      LAYER met1 ;
        RECT 0.240 9.220 0.520 9.870 ;
        RECT 0.240 8.620 0.630 9.220 ;
        RECT 0.240 5.070 0.520 8.620 ;
        RECT 0.770 8.410 0.960 9.870 ;
        RECT 2.170 9.050 2.480 9.490 ;
        RECT 7.250 8.660 7.480 9.870 ;
        RECT 8.470 8.900 8.700 9.870 ;
        RECT 0.740 8.380 0.960 8.410 ;
        RECT 0.730 8.110 0.980 8.380 ;
        RECT 0.730 8.100 0.970 8.110 ;
        RECT 0.740 7.860 0.970 8.100 ;
        RECT 2.010 8.090 2.330 8.410 ;
        RECT 7.220 7.870 7.480 8.660 ;
        RECT 8.460 8.650 8.700 8.900 ;
        RECT 0.770 5.830 0.930 7.860 ;
        RECT 1.120 7.300 1.360 7.430 ;
        RECT 1.100 6.980 1.360 7.300 ;
        RECT 1.100 6.380 1.360 6.700 ;
        RECT 1.120 6.260 1.360 6.380 ;
        RECT 0.740 5.590 0.970 5.830 ;
        RECT 7.250 5.720 7.480 7.870 ;
        RECT 0.730 5.580 0.970 5.590 ;
        RECT 0.730 5.310 0.980 5.580 ;
        RECT 2.010 5.330 2.330 5.650 ;
        RECT 0.740 5.280 0.960 5.310 ;
        RECT 0.240 4.470 0.630 5.070 ;
        RECT 0.240 3.820 0.520 4.470 ;
        RECT 0.770 3.820 0.960 5.280 ;
        RECT 7.220 4.930 7.480 5.720 ;
        RECT 2.170 4.200 2.480 4.640 ;
        RECT 7.250 3.820 7.480 4.930 ;
        RECT 8.470 3.820 8.700 8.650 ;
        RECT 9.270 8.500 9.590 8.820 ;
        RECT 9.300 4.810 9.620 5.130 ;
        RECT 10.760 3.830 11.180 9.870 ;
        RECT 19.700 3.820 20.120 9.870 ;
        RECT 22.180 3.820 22.410 9.870 ;
        RECT 23.400 8.660 23.630 9.870 ;
        RECT 28.400 9.050 28.710 9.490 ;
        RECT 23.400 7.870 23.660 8.660 ;
        RECT 28.550 8.090 28.870 8.410 ;
        RECT 23.400 5.720 23.630 7.870 ;
        RECT 29.520 7.300 29.760 7.430 ;
        RECT 29.520 6.980 29.780 7.300 ;
        RECT 26.400 6.000 26.680 6.050 ;
        RECT 23.400 4.930 23.660 5.720 ;
        RECT 26.400 5.700 26.720 6.000 ;
        RECT 28.550 5.330 28.870 5.650 ;
        RECT 31.380 5.480 31.700 5.800 ;
        RECT 23.400 3.820 23.630 4.930 ;
        RECT 28.300 4.880 28.620 5.200 ;
        RECT 27.190 4.350 27.510 4.670 ;
        RECT 12.460 3.230 12.630 3.400 ;
        RECT 18.250 3.230 18.420 3.400 ;
        RECT 27.920 3.070 28.240 3.390 ;
        RECT 29.130 3.300 29.450 3.620 ;
        RECT 31.430 3.260 31.750 3.580 ;
        RECT 12.440 2.640 12.760 2.940 ;
        RECT 12.470 2.540 12.640 2.640 ;
        RECT 18.140 2.570 18.460 2.890 ;
        RECT 18.250 2.550 18.420 2.570 ;
        RECT 29.130 2.470 29.450 2.790 ;
        RECT 31.420 2.540 31.740 2.860 ;
        RECT 29.080 1.820 29.400 2.140 ;
        RECT 29.080 0.990 29.400 1.310 ;
        RECT 18.140 0.060 18.460 0.360 ;
        RECT 29.130 0.340 29.450 0.660 ;
        RECT 31.340 0.290 31.660 0.610 ;
      LAYER via ;
        RECT 2.190 9.080 2.450 9.340 ;
        RECT 2.040 8.120 2.300 8.380 ;
        RECT 1.100 7.010 1.360 7.270 ;
        RECT 1.100 6.410 1.360 6.670 ;
        RECT 2.040 5.360 2.300 5.620 ;
        RECT 2.190 4.350 2.450 4.610 ;
        RECT 9.300 8.530 9.560 8.790 ;
        RECT 9.330 4.840 9.590 5.100 ;
        RECT 28.430 9.080 28.690 9.340 ;
        RECT 28.580 8.120 28.840 8.380 ;
        RECT 29.520 7.010 29.780 7.270 ;
        RECT 26.430 5.720 26.690 5.980 ;
        RECT 28.580 5.360 28.840 5.620 ;
        RECT 31.410 5.510 31.670 5.770 ;
        RECT 28.330 4.910 28.590 5.170 ;
        RECT 27.220 4.380 27.480 4.640 ;
        RECT 27.950 3.100 28.210 3.360 ;
        RECT 29.160 3.330 29.420 3.590 ;
        RECT 31.460 3.290 31.720 3.550 ;
        RECT 12.470 2.660 12.730 2.920 ;
        RECT 18.170 2.600 18.430 2.860 ;
        RECT 29.160 2.500 29.420 2.760 ;
        RECT 31.450 2.570 31.710 2.830 ;
        RECT 29.110 1.850 29.370 2.110 ;
        RECT 29.110 1.020 29.370 1.280 ;
        RECT 29.160 0.370 29.420 0.630 ;
        RECT 18.170 0.080 18.430 0.340 ;
        RECT 31.370 0.320 31.630 0.580 ;
      LAYER met2 ;
        RECT 2.170 9.370 2.480 9.380 ;
        RECT 28.400 9.370 28.710 9.380 ;
        RECT 0.000 9.190 11.530 9.370 ;
        RECT 19.350 9.190 30.880 9.370 ;
        RECT 2.170 9.050 2.480 9.190 ;
        RECT 28.400 9.050 28.710 9.190 ;
        RECT 9.280 8.780 9.590 8.830 ;
        RECT 9.280 8.770 9.740 8.780 ;
        RECT 9.280 8.590 11.530 8.770 ;
        RECT 9.280 8.500 9.590 8.590 ;
        RECT 2.020 8.350 2.330 8.420 ;
        RECT 0.000 8.340 2.330 8.350 ;
        RECT 28.550 8.350 28.860 8.420 ;
        RECT 0.000 8.130 11.530 8.340 ;
        RECT 1.310 8.120 11.530 8.130 ;
        RECT 28.550 8.130 30.880 8.350 ;
        RECT 2.020 8.090 2.330 8.120 ;
        RECT 28.550 8.090 28.860 8.130 ;
        RECT 1.070 7.150 11.530 7.370 ;
        RECT 1.070 7.010 1.390 7.150 ;
        RECT 1.090 6.670 1.350 7.010 ;
        RECT 1.070 6.410 1.390 6.670 ;
        RECT 9.310 5.060 9.620 5.140 ;
        RECT 9.310 4.850 11.530 5.060 ;
        RECT 9.310 4.810 9.620 4.850 ;
        RECT 2.170 4.500 2.480 4.640 ;
        RECT 0.000 4.490 2.480 4.500 ;
        RECT 0.000 4.340 11.530 4.490 ;
        RECT 0.000 4.320 2.480 4.340 ;
        RECT 2.170 4.310 2.480 4.320 ;
        RECT 13.260 3.330 22.270 3.550 ;
        RECT 12.440 2.890 12.760 2.940 ;
        RECT 12.440 2.640 18.460 2.890 ;
        RECT 18.140 2.570 18.460 2.640 ;
        RECT 13.310 1.550 18.970 1.770 ;
        RECT 18.750 1.220 18.970 1.550 ;
        RECT 22.050 1.720 22.270 3.330 ;
        RECT 22.050 1.500 24.900 1.720 ;
        RECT 29.080 1.270 29.390 1.310 ;
        RECT 23.120 1.220 29.390 1.270 ;
        RECT 18.750 1.060 29.390 1.220 ;
        RECT 18.750 1.000 23.510 1.060 ;
        RECT 29.080 0.980 29.390 1.060 ;
        RECT 29.130 0.580 29.440 0.660 ;
        RECT 31.340 0.580 31.650 0.620 ;
        RECT 29.130 0.350 31.840 0.580 ;
        RECT 29.130 0.330 29.440 0.350 ;
        RECT 31.340 0.290 31.650 0.350 ;
  END
END sky130_hilas_TA2Cell_1FG

MACRO sky130_hilas_swc4x1cellOverlap
  CLASS CORE ;
  FOREIGN sky130_hilas_swc4x1cellOverlap ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 6.710 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
      LAYER nwell ;
        RECT 4.870 6.360 7.590 6.650 ;
        RECT 0.010 4.500 1.740 6.360 ;
        RECT 0.000 2.660 1.740 4.500 ;
        RECT 4.870 6.350 10.070 6.360 ;
        RECT 4.870 3.560 10.080 6.350 ;
        RECT 0.010 0.310 1.740 2.660 ;
        RECT 4.860 0.330 10.080 3.560 ;
        RECT 4.860 0.320 10.070 0.330 ;
        RECT 4.860 0.060 7.580 0.320 ;
      LAYER li1 ;
        RECT 5.270 5.080 7.220 6.250 ;
        RECT 7.620 5.950 7.940 5.960 ;
        RECT 7.620 5.780 8.200 5.950 ;
        RECT 7.620 5.730 7.950 5.780 ;
        RECT 7.620 5.700 7.940 5.730 ;
        RECT 9.480 5.680 9.680 6.030 ;
        RECT 7.620 5.370 7.940 5.410 ;
        RECT 7.620 5.330 7.950 5.370 ;
        RECT 7.620 5.160 8.200 5.330 ;
        RECT 7.620 5.150 7.940 5.160 ;
        RECT 8.750 5.090 8.950 5.660 ;
        RECT 9.480 5.650 9.690 5.680 ;
        RECT 9.470 5.060 9.690 5.650 ;
        RECT 5.270 3.550 7.220 4.720 ;
        RECT 7.620 4.520 7.940 4.530 ;
        RECT 7.620 4.350 8.200 4.520 ;
        RECT 7.620 4.310 7.950 4.350 ;
        RECT 7.620 4.270 7.940 4.310 ;
        RECT 8.750 4.020 8.950 4.590 ;
        RECT 9.470 4.030 9.690 4.620 ;
        RECT 9.480 4.000 9.690 4.030 ;
        RECT 7.620 3.950 7.940 3.980 ;
        RECT 7.620 3.900 7.950 3.950 ;
        RECT 7.620 3.730 8.200 3.900 ;
        RECT 7.620 3.720 7.940 3.730 ;
        RECT 9.480 3.650 9.680 4.000 ;
        RECT 0.430 3.110 0.980 3.540 ;
        RECT 8.870 3.250 9.310 3.420 ;
        RECT 5.260 1.990 7.210 3.160 ;
        RECT 7.620 2.940 7.940 2.950 ;
        RECT 7.620 2.770 8.200 2.940 ;
        RECT 7.620 2.720 7.950 2.770 ;
        RECT 7.620 2.690 7.940 2.720 ;
        RECT 9.480 2.670 9.680 3.020 ;
        RECT 7.620 2.360 7.940 2.400 ;
        RECT 7.620 2.320 7.950 2.360 ;
        RECT 7.620 2.150 8.200 2.320 ;
        RECT 7.620 2.140 7.940 2.150 ;
        RECT 8.750 2.080 8.950 2.650 ;
        RECT 9.480 2.640 9.690 2.670 ;
        RECT 9.470 2.050 9.690 2.640 ;
        RECT 5.260 0.450 7.210 1.620 ;
        RECT 7.620 1.520 7.940 1.530 ;
        RECT 7.620 1.350 8.200 1.520 ;
        RECT 7.620 1.310 7.950 1.350 ;
        RECT 7.620 1.270 7.940 1.310 ;
        RECT 8.750 1.020 8.950 1.590 ;
        RECT 9.470 1.030 9.690 1.620 ;
        RECT 9.480 1.000 9.690 1.030 ;
        RECT 7.620 0.950 7.940 0.980 ;
        RECT 7.620 0.900 7.950 0.950 ;
        RECT 7.620 0.730 8.200 0.900 ;
        RECT 7.620 0.720 7.940 0.730 ;
        RECT 9.480 0.650 9.680 1.000 ;
      LAYER mcon ;
        RECT 5.750 5.910 5.920 6.080 ;
        RECT 5.750 5.570 5.920 5.740 ;
        RECT 7.680 5.740 7.850 5.910 ;
        RECT 8.760 5.450 8.930 5.620 ;
        RECT 5.750 5.230 5.920 5.400 ;
        RECT 7.680 5.190 7.850 5.360 ;
        RECT 9.490 5.480 9.660 5.650 ;
        RECT 5.750 4.380 5.920 4.550 ;
        RECT 7.680 4.320 7.850 4.490 ;
        RECT 5.750 4.040 5.920 4.210 ;
        RECT 8.760 4.060 8.930 4.230 ;
        RECT 9.490 4.030 9.660 4.200 ;
        RECT 5.750 3.700 5.920 3.870 ;
        RECT 7.680 3.770 7.850 3.940 ;
        RECT 0.430 3.190 0.700 3.460 ;
        RECT 9.130 3.250 9.310 3.420 ;
        RECT 5.740 2.820 5.910 2.990 ;
        RECT 7.680 2.730 7.850 2.900 ;
        RECT 5.740 2.480 5.910 2.650 ;
        RECT 8.760 2.440 8.930 2.610 ;
        RECT 5.740 2.140 5.910 2.310 ;
        RECT 7.680 2.180 7.850 2.350 ;
        RECT 9.490 2.470 9.660 2.640 ;
        RECT 5.740 1.280 5.910 1.450 ;
        RECT 7.680 1.320 7.850 1.490 ;
        RECT 5.740 0.940 5.910 1.110 ;
        RECT 8.760 1.060 8.930 1.230 ;
        RECT 9.490 1.030 9.660 1.200 ;
        RECT 5.740 0.600 5.910 0.770 ;
        RECT 7.680 0.770 7.850 0.940 ;
      LAYER met1 ;
        RECT 0.360 0.310 0.760 6.300 ;
        RECT 5.710 5.660 5.970 6.140 ;
        RECT 7.610 5.670 7.930 5.990 ;
        RECT 8.750 5.680 8.910 6.360 ;
        RECT 8.750 5.660 8.950 5.680 ;
        RECT 5.700 5.140 5.970 5.660 ;
        RECT 5.700 4.690 5.960 5.140 ;
        RECT 7.610 5.120 7.930 5.440 ;
        RECT 8.730 5.420 8.960 5.660 ;
        RECT 8.750 5.200 8.950 5.420 ;
        RECT 9.120 5.370 9.310 6.360 ;
        RECT 9.560 5.710 9.720 6.360 ;
        RECT 9.140 5.250 9.310 5.370 ;
        RECT 5.710 4.130 5.970 4.610 ;
        RECT 7.610 4.240 7.930 4.560 ;
        RECT 8.750 4.480 8.910 5.200 ;
        RECT 8.750 4.260 8.950 4.480 ;
        RECT 9.150 4.430 9.310 5.250 ;
        RECT 9.450 5.160 9.720 5.710 ;
        RECT 9.450 5.110 9.730 5.160 ;
        RECT 9.560 5.020 9.730 5.110 ;
        RECT 9.560 4.660 9.720 5.020 ;
        RECT 9.560 4.570 9.730 4.660 ;
        RECT 9.140 4.310 9.310 4.430 ;
        RECT 5.700 3.610 5.970 4.130 ;
        RECT 8.730 4.020 8.960 4.260 ;
        RECT 7.610 3.690 7.930 4.010 ;
        RECT 8.750 4.000 8.950 4.020 ;
        RECT 5.700 3.160 5.960 3.610 ;
        RECT 5.700 2.570 5.960 3.050 ;
        RECT 7.610 2.660 7.930 2.980 ;
        RECT 8.750 2.670 8.910 4.000 ;
        RECT 9.120 3.450 9.310 4.310 ;
        RECT 9.450 4.520 9.730 4.570 ;
        RECT 9.450 3.970 9.720 4.520 ;
        RECT 9.100 3.220 9.340 3.450 ;
        RECT 8.750 2.650 8.950 2.670 ;
        RECT 5.690 2.050 5.960 2.570 ;
        RECT 7.610 2.110 7.930 2.430 ;
        RECT 8.730 2.410 8.960 2.650 ;
        RECT 8.750 2.190 8.950 2.410 ;
        RECT 9.120 2.360 9.310 3.220 ;
        RECT 9.560 2.700 9.720 3.970 ;
        RECT 9.140 2.240 9.310 2.360 ;
        RECT 5.690 1.600 5.950 2.050 ;
        RECT 5.700 1.030 5.960 1.510 ;
        RECT 7.610 1.240 7.930 1.560 ;
        RECT 8.750 1.480 8.910 2.190 ;
        RECT 8.750 1.260 8.950 1.480 ;
        RECT 9.150 1.430 9.310 2.240 ;
        RECT 9.450 2.150 9.720 2.700 ;
        RECT 9.450 2.100 9.730 2.150 ;
        RECT 9.560 2.010 9.730 2.100 ;
        RECT 9.560 1.660 9.720 2.010 ;
        RECT 9.560 1.570 9.730 1.660 ;
        RECT 9.140 1.310 9.310 1.430 ;
        RECT 5.690 0.510 5.960 1.030 ;
        RECT 8.730 1.020 8.960 1.260 ;
        RECT 7.610 0.690 7.930 1.010 ;
        RECT 8.750 1.000 8.950 1.020 ;
        RECT 5.690 0.060 5.950 0.510 ;
        RECT 8.750 0.320 8.910 1.000 ;
        RECT 9.120 0.320 9.310 1.310 ;
        RECT 9.450 1.520 9.730 1.570 ;
        RECT 9.450 0.970 9.720 1.520 ;
        RECT 9.560 0.320 9.720 0.970 ;
      LAYER via ;
        RECT 7.640 5.700 7.900 5.960 ;
        RECT 7.640 5.150 7.900 5.410 ;
        RECT 7.640 4.270 7.900 4.530 ;
        RECT 7.640 3.720 7.900 3.980 ;
        RECT 7.640 2.690 7.900 2.950 ;
        RECT 7.640 2.140 7.900 2.400 ;
        RECT 7.640 1.270 7.900 1.530 ;
        RECT 7.640 0.720 7.900 0.980 ;
      LAYER met2 ;
        RECT 7.610 5.860 7.920 6.000 ;
        RECT 0.000 5.680 10.080 5.860 ;
        RECT 7.610 5.670 7.920 5.680 ;
        RECT 7.610 5.430 7.920 5.450 ;
        RECT 0.000 5.250 10.080 5.430 ;
        RECT 7.610 5.120 7.920 5.250 ;
        RECT 7.610 4.430 7.920 4.560 ;
        RECT 0.000 4.250 10.080 4.430 ;
        RECT 7.610 4.230 7.920 4.250 ;
        RECT 7.610 4.000 7.920 4.010 ;
        RECT 0.000 3.930 7.600 4.000 ;
        RECT 7.610 3.930 10.080 4.000 ;
        RECT 0.000 3.820 10.080 3.930 ;
        RECT 7.610 3.680 7.920 3.820 ;
        RECT 7.610 2.850 7.920 2.990 ;
        RECT 7.610 2.840 10.080 2.850 ;
        RECT 0.020 2.670 10.080 2.840 ;
        RECT 7.610 2.660 7.920 2.670 ;
        RECT 7.610 2.420 7.920 2.440 ;
        RECT 0.020 2.250 10.080 2.420 ;
        RECT 7.520 2.240 10.080 2.250 ;
        RECT 7.610 2.110 7.920 2.240 ;
        RECT 7.610 1.440 7.920 1.560 ;
        RECT 0.020 1.430 7.920 1.440 ;
        RECT 0.020 1.270 10.080 1.430 ;
        RECT 0.800 1.180 2.340 1.270 ;
        RECT 7.520 1.250 10.080 1.270 ;
        RECT 7.610 1.230 7.920 1.250 ;
        RECT 7.610 1.000 7.920 1.010 ;
        RECT 0.020 0.830 10.080 1.000 ;
        RECT 7.610 0.820 10.080 0.830 ;
        RECT 7.610 0.680 7.920 0.820 ;
  END
END sky130_hilas_swc4x1cellOverlap

MACRO sky130_hilas_capacitorSize02
  CLASS CORE ;
  FOREIGN sky130_hilas_capacitorSize02 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.970 BY 5.830 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 7.230 2.620 7.890 3.280 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 0.110 3.200 0.770 3.260 ;
        RECT 1.160 3.200 2.170 3.210 ;
        RECT 0.110 2.700 3.800 3.200 ;
        RECT 0.110 2.690 1.520 2.700 ;
        RECT 0.110 2.600 0.770 2.690 ;
        RECT 3.160 1.580 3.790 2.700 ;
        RECT 3.160 1.570 5.310 1.580 ;
        RECT 1.840 1.270 5.310 1.570 ;
        RECT 1.840 1.100 4.850 1.270 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 0.000 5.280 7.970 5.460 ;
        RECT 0.000 4.850 7.970 5.030 ;
        RECT 0.030 3.850 7.970 4.030 ;
        RECT 0.030 3.420 7.970 3.600 ;
        RECT 0.240 3.080 0.610 3.140 ;
        RECT 0.020 2.800 0.610 3.080 ;
        RECT 0.240 2.740 0.610 2.800 ;
        RECT 7.360 3.100 7.730 3.160 ;
        RECT 7.360 2.820 7.970 3.100 ;
        RECT 7.360 2.760 7.730 2.820 ;
        RECT 0.030 2.270 7.970 2.440 ;
        RECT 0.030 1.850 7.970 2.020 ;
        RECT 0.030 0.870 7.970 1.040 ;
        RECT 0.030 0.430 7.970 0.600 ;
      LAYER via2 ;
        RECT 0.290 2.800 0.570 3.080 ;
        RECT 7.410 2.820 7.690 3.100 ;
      LAYER met3 ;
        RECT 1.460 5.800 3.770 5.830 ;
        RECT 1.460 3.310 5.690 5.800 ;
        RECT 0.020 2.540 0.810 3.290 ;
        RECT 1.460 2.560 7.930 3.310 ;
        RECT 1.460 0.020 5.690 2.560 ;
        RECT 3.740 0.000 5.690 0.020 ;
      LAYER via3 ;
        RECT 0.210 2.690 0.640 3.170 ;
        RECT 7.330 2.710 7.760 3.190 ;
  END
END sky130_hilas_capacitorSize02

MACRO sky130_hilas_TopProtectStructure
  CLASS CORE ;
  FOREIGN sky130_hilas_TopProtectStructure ;
  ORIGIN 0.000 0.000 ;
  SIZE 373.410 BY 389.400 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN IO07
    ANTENNAGATEAREA 54.899799 ;
    ANTENNADIFFAREA 1293.556030 ;
    PORT
      LAYER nwell ;
        RECT 128.920 378.090 131.660 381.590 ;
        RECT 134.530 377.000 144.220 381.600 ;
        RECT 151.360 381.580 154.070 381.620 ;
        RECT 133.930 375.610 144.220 377.000 ;
        RECT 145.800 375.590 149.800 381.580 ;
        RECT 151.350 379.930 154.070 381.580 ;
        RECT 156.550 379.880 158.770 381.570 ;
        RECT 179.660 380.440 191.710 386.380 ;
        RECT 208.250 380.440 220.300 386.380 ;
        RECT 236.840 380.440 248.890 386.380 ;
        RECT 265.430 380.440 277.480 386.380 ;
        RECT 294.020 380.440 306.070 386.380 ;
        RECT 322.610 380.440 334.660 386.380 ;
        RECT 351.200 380.440 363.250 386.380 ;
        RECT 151.360 378.590 154.070 378.630 ;
        RECT 151.350 375.930 154.070 378.590 ;
        RECT 185.420 357.320 188.840 363.370 ;
        RECT 205.190 357.080 208.500 369.140 ;
        RECT 214.980 368.400 216.710 369.150 ;
        RECT 214.970 364.830 216.710 368.400 ;
        RECT 210.230 360.730 212.950 362.380 ;
        RECT 214.980 362.370 216.710 364.830 ;
        RECT 210.240 360.690 212.950 360.730 ;
        RECT 210.240 359.360 212.950 359.400 ;
        RECT 210.230 359.300 212.950 359.360 ;
        RECT 209.150 359.290 212.950 359.300 ;
        RECT 210.230 357.710 212.950 359.290 ;
        RECT 214.970 358.800 216.710 362.370 ;
        RECT 214.980 357.210 216.710 358.800 ;
        RECT 213.350 357.080 216.710 357.210 ;
        RECT 224.550 368.400 226.280 369.150 ;
        RECT 224.550 364.830 226.290 368.400 ;
        RECT 228.310 366.760 231.030 368.410 ;
        RECT 228.310 366.720 231.020 366.760 ;
        RECT 232.760 365.440 236.070 369.150 ;
        RECT 364.450 366.940 370.390 378.990 ;
        RECT 230.750 365.430 236.070 365.440 ;
        RECT 228.310 365.330 236.070 365.430 ;
        RECT 224.550 362.370 226.280 364.830 ;
        RECT 228.310 363.740 237.240 365.330 ;
        RECT 230.750 362.380 237.240 363.740 ;
        RECT 224.550 358.800 226.290 362.370 ;
        RECT 228.310 360.690 237.240 362.380 ;
        RECT 230.750 359.400 237.240 360.690 ;
        RECT 228.310 359.390 237.240 359.400 ;
        RECT 228.310 359.360 231.020 359.390 ;
        RECT 224.550 357.080 226.280 358.800 ;
        RECT 228.310 357.710 231.030 359.360 ;
        RECT 232.100 357.080 237.240 359.390 ;
        RECT 205.840 355.350 207.570 357.080 ;
        RECT 205.830 353.510 207.570 355.350 ;
        RECT 205.840 351.160 207.570 353.510 ;
        RECT 213.350 351.180 215.910 357.080 ;
        RECT 232.100 353.250 233.960 357.080 ;
        RECT 235.960 353.250 237.240 357.080 ;
        RECT 213.350 351.170 215.900 351.180 ;
        RECT 142.730 339.210 143.290 341.180 ;
        RECT 169.590 336.310 172.100 342.550 ;
        RECT 364.450 338.350 370.390 350.400 ;
        RECT 137.560 324.850 138.180 330.550 ;
        RECT 175.840 326.160 176.860 331.860 ;
        RECT 185.650 326.190 186.670 331.890 ;
        RECT 232.870 314.260 234.220 329.730 ;
        RECT 232.860 313.790 234.220 314.260 ;
        RECT 364.450 309.760 370.390 321.810 ;
        RECT 364.450 281.170 370.390 293.220 ;
        RECT 364.450 252.580 370.390 264.630 ;
        RECT 364.450 223.990 370.390 236.040 ;
        RECT 364.450 195.400 370.390 207.450 ;
      LAYER met3 ;
        RECT 202.240 366.860 202.690 367.610 ;
        RECT 202.240 360.700 202.610 366.860 ;
        RECT 203.280 366.850 203.730 367.600 ;
        RECT 203.360 364.210 203.730 366.850 ;
        RECT 203.360 363.610 203.800 364.210 ;
        RECT 202.240 360.370 202.730 360.700 ;
        RECT 202.290 360.210 202.730 360.370 ;
        RECT 203.360 358.500 203.730 363.610 ;
        RECT 203.350 357.630 203.820 358.500 ;
    END
  END IO07
  PIN IO08
    ANTENNAGATEAREA 54.899799 ;
    ANTENNADIFFAREA 1281.299683 ;
    PORT
      LAYER met2 ;
        RECT 164.790 385.910 364.920 387.310 ;
        RECT 165.260 385.900 166.190 385.910 ;
        RECT 193.850 385.900 194.780 385.910 ;
        RECT 222.440 385.900 223.370 385.910 ;
        RECT 251.030 385.900 251.960 385.910 ;
        RECT 279.620 385.900 280.550 385.910 ;
        RECT 308.210 385.900 309.140 385.910 ;
        RECT 336.800 385.900 337.730 385.910 ;
        RECT 165.510 385.580 165.680 385.900 ;
        RECT 129.360 384.190 184.830 385.580 ;
        RECT 194.100 384.790 194.270 385.900 ;
        RECT 222.690 384.790 222.860 385.900 ;
        RECT 251.280 384.790 251.450 385.900 ;
        RECT 279.870 384.790 280.040 385.900 ;
        RECT 308.460 384.790 308.630 385.900 ;
        RECT 337.050 384.790 337.220 385.900 ;
        RECT 368.720 385.020 369.910 385.030 ;
        RECT 356.920 384.500 369.910 385.020 ;
        RECT 125.780 382.380 126.460 383.600 ;
        RECT 127.010 382.380 127.460 382.480 ;
        RECT 125.780 382.150 127.460 382.380 ;
        RECT 125.780 381.280 126.460 382.150 ;
        RECT 127.010 382.050 127.460 382.150 ;
        RECT 132.290 381.410 132.610 381.460 ;
        RECT 129.430 381.170 132.610 381.410 ;
        RECT 129.430 381.150 129.750 381.170 ;
        RECT 191.130 381.010 191.770 384.020 ;
        RECT 209.630 381.810 210.090 381.830 ;
        RECT 219.720 381.810 220.360 384.020 ;
        RECT 240.500 381.810 241.360 383.160 ;
        RECT 209.630 381.440 241.360 381.810 ;
        RECT 209.630 381.420 210.090 381.440 ;
        RECT 219.720 381.010 220.360 381.440 ;
        RECT 240.500 381.060 241.360 381.440 ;
        RECT 248.310 381.010 248.950 384.020 ;
        RECT 276.900 381.010 277.540 384.020 ;
        RECT 305.490 381.010 306.130 384.020 ;
        RECT 334.080 381.010 334.720 384.020 ;
        RECT 356.710 383.740 369.910 384.500 ;
        RECT 362.670 381.010 363.310 383.740 ;
        RECT 367.750 382.420 369.910 383.740 ;
        RECT 164.790 380.660 364.920 381.010 ;
        RECT 125.630 380.180 128.110 380.190 ;
        RECT 129.420 380.180 129.740 380.380 ;
        RECT 130.150 380.180 130.460 380.390 ;
        RECT 130.830 380.180 131.150 380.390 ;
        RECT 131.490 380.180 146.140 380.310 ;
        RECT 125.630 380.100 146.140 380.180 ;
        RECT 125.630 379.930 131.630 380.100 ;
        RECT 145.560 380.090 146.310 380.100 ;
        RECT 125.630 379.790 131.490 379.930 ;
        RECT 127.900 379.420 131.490 379.790 ;
        RECT 131.980 379.630 132.300 379.950 ;
        RECT 145.560 379.790 147.180 380.090 ;
        RECT 164.790 379.860 365.020 380.660 ;
        RECT 145.560 379.650 145.800 379.790 ;
        RECT 146.880 379.730 147.180 379.790 ;
        RECT 129.420 379.290 129.740 379.420 ;
        RECT 130.150 379.290 130.460 379.420 ;
        RECT 130.850 379.290 131.170 379.420 ;
        RECT 132.000 379.290 132.270 379.630 ;
        RECT 145.540 379.320 145.850 379.650 ;
        RECT 146.880 379.410 147.210 379.730 ;
        RECT 147.610 379.720 365.020 379.860 ;
        RECT 146.900 379.400 147.210 379.410 ;
        RECT 147.590 379.610 365.020 379.720 ;
        RECT 147.590 379.560 170.480 379.610 ;
        RECT 147.590 379.400 147.910 379.560 ;
        RECT 170.000 379.500 170.480 379.560 ;
        RECT 170.010 379.480 170.460 379.500 ;
        RECT 190.230 379.480 192.860 379.610 ;
        RECT 218.820 379.480 221.450 379.610 ;
        RECT 247.410 379.480 250.040 379.610 ;
        RECT 276.000 379.480 278.630 379.610 ;
        RECT 304.590 379.480 307.220 379.610 ;
        RECT 333.180 379.480 335.810 379.610 ;
        RECT 147.590 379.390 147.900 379.400 ;
        RECT 129.360 379.150 184.830 379.290 ;
        RECT 190.230 379.190 192.780 379.480 ;
        RECT 189.770 379.150 192.780 379.190 ;
        RECT 125.780 378.190 126.460 379.070 ;
        RECT 127.110 378.580 127.540 379.050 ;
        RECT 129.360 378.970 192.780 379.150 ;
        RECT 218.820 378.970 221.370 379.480 ;
        RECT 247.410 378.970 249.960 379.480 ;
        RECT 276.000 378.970 278.550 379.480 ;
        RECT 304.590 378.970 307.140 379.480 ;
        RECT 333.180 378.970 335.730 379.480 ;
        RECT 361.770 379.050 365.020 379.610 ;
        RECT 367.750 379.050 369.030 382.420 ;
        RECT 361.770 378.970 369.030 379.050 ;
        RECT 129.360 378.750 191.240 378.970 ;
        RECT 218.820 378.900 219.440 378.970 ;
        RECT 247.410 378.900 248.030 378.970 ;
        RECT 276.000 378.900 276.620 378.970 ;
        RECT 304.590 378.900 305.210 378.970 ;
        RECT 333.180 378.900 333.800 378.970 ;
        RECT 361.770 378.900 362.390 378.970 ;
        RECT 129.360 378.580 184.830 378.750 ;
        RECT 189.770 378.710 191.190 378.750 ;
        RECT 127.110 378.570 184.830 378.580 ;
        RECT 127.200 378.350 184.830 378.570 ;
        RECT 129.360 378.190 184.830 378.350 ;
        RECT 125.780 377.890 184.830 378.190 ;
        RECT 362.980 378.410 369.030 378.970 ;
        RECT 362.980 378.130 365.020 378.410 ;
        RECT 125.780 377.870 129.440 377.890 ;
        RECT 125.780 376.750 126.460 377.870 ;
        RECT 131.560 377.710 131.870 377.890 ;
        RECT 128.470 377.610 131.870 377.710 ;
        RECT 128.470 377.480 131.850 377.610 ;
        RECT 171.670 377.540 172.170 377.570 ;
        RECT 177.390 377.540 177.890 377.570 ;
        RECT 128.470 377.450 128.790 377.480 ;
        RECT 171.670 377.130 201.830 377.540 ;
        RECT 362.910 377.510 365.020 378.130 ;
        RECT 171.820 377.100 201.830 377.130 ;
        RECT 130.130 376.540 130.440 376.750 ;
        RECT 131.560 376.540 131.870 376.770 ;
        RECT 127.780 376.380 132.700 376.540 ;
        RECT 125.970 376.210 132.700 376.380 ;
        RECT 167.250 376.530 167.750 376.550 ;
        RECT 172.990 376.530 173.430 376.580 ;
        RECT 187.360 376.530 187.860 376.550 ;
        RECT 125.970 376.160 132.710 376.210 ;
        RECT 125.970 376.050 132.730 376.160 ;
        RECT 167.250 376.110 193.760 376.530 ;
        RECT 167.400 376.090 193.760 376.110 ;
        RECT 172.990 376.080 173.430 376.090 ;
        RECT 193.160 376.070 193.660 376.090 ;
        RECT 125.970 375.980 128.240 376.050 ;
        RECT 125.970 375.780 126.370 375.980 ;
        RECT 129.340 375.840 129.650 376.050 ;
        RECT 130.270 375.840 130.580 376.050 ;
        RECT 130.970 375.840 131.280 376.050 ;
        RECT 131.710 375.870 132.730 376.050 ;
        RECT 144.820 375.870 145.130 375.990 ;
        RECT 154.680 375.870 154.990 376.010 ;
        RECT 131.710 375.840 154.990 375.870 ;
        RECT 125.620 375.380 126.370 375.780 ;
        RECT 131.730 375.680 154.990 375.840 ;
        RECT 131.730 375.660 154.960 375.680 ;
        RECT 237.880 375.170 238.650 375.320 ;
        RECT 128.390 374.750 238.650 375.170 ;
        RECT 237.880 374.610 238.650 374.750 ;
        RECT 125.330 373.930 126.010 374.600 ;
        RECT 134.250 373.930 134.720 373.950 ;
        RECT 85.990 373.240 90.080 373.490 ;
        RECT 125.330 373.350 134.720 373.930 ;
        RECT 125.330 373.240 126.050 373.350 ;
        RECT 134.250 373.330 134.720 373.350 ;
        RECT 164.500 373.320 164.800 373.380 ;
        RECT 205.820 373.320 206.120 373.350 ;
        RECT 85.990 371.780 127.960 373.240 ;
        RECT 164.500 373.090 206.190 373.320 ;
        RECT 164.500 373.060 164.800 373.090 ;
        RECT 205.820 373.010 206.120 373.090 ;
        RECT 157.420 372.660 157.730 372.680 ;
        RECT 147.630 372.580 147.950 372.590 ;
        RECT 157.420 372.580 157.740 372.660 ;
        RECT 181.600 372.590 181.920 372.610 ;
        RECT 181.600 372.580 181.930 372.590 ;
        RECT 188.370 372.580 188.690 372.610 ;
        RECT 203.140 372.580 203.460 372.600 ;
        RECT 217.800 372.580 218.360 372.720 ;
        RECT 147.630 372.350 218.360 372.580 ;
        RECT 147.630 372.270 147.950 372.350 ;
        RECT 157.420 372.340 157.730 372.350 ;
        RECT 181.600 372.330 181.930 372.350 ;
        RECT 188.370 372.330 188.690 372.350 ;
        RECT 203.140 372.340 203.460 372.350 ;
        RECT 217.800 372.210 218.360 372.350 ;
        RECT 153.420 372.130 153.790 372.190 ;
        RECT 216.620 372.130 217.160 372.150 ;
        RECT 153.420 371.900 217.160 372.130 ;
        RECT 153.420 371.840 153.790 371.900 ;
        RECT 85.990 371.480 128.430 371.780 ;
        RECT 185.220 371.680 185.500 371.690 ;
        RECT 156.250 371.670 156.560 371.680 ;
        RECT 185.200 371.670 185.520 371.680 ;
        RECT 187.930 371.670 188.250 371.700 ;
        RECT 202.250 371.670 202.570 371.730 ;
        RECT 215.540 371.670 216.080 371.680 ;
        RECT 85.990 370.990 127.960 371.480 ;
        RECT 156.250 371.440 216.080 371.670 ;
        RECT 216.620 371.590 217.160 371.900 ;
        RECT 156.250 371.410 156.580 371.440 ;
        RECT 185.200 371.420 185.520 371.440 ;
        RECT 187.930 371.420 188.250 371.440 ;
        RECT 185.220 371.410 185.500 371.420 ;
        RECT 156.250 371.390 156.560 371.410 ;
        RECT 150.170 371.210 150.490 371.220 ;
        RECT 214.600 371.210 215.130 371.240 ;
        RECT 85.990 370.390 90.080 370.990 ;
        RECT 125.290 370.980 125.800 370.990 ;
        RECT 144.930 370.980 145.330 370.990 ;
        RECT 125.290 370.630 145.330 370.980 ;
        RECT 150.170 370.980 215.130 371.210 ;
        RECT 215.540 371.120 216.080 371.440 ;
        RECT 150.170 370.920 150.490 370.980 ;
        RECT 125.290 370.590 125.800 370.630 ;
        RECT 144.930 370.600 145.330 370.630 ;
        RECT 182.070 370.630 182.390 370.670 ;
        RECT 197.720 370.630 199.000 370.730 ;
        RECT 214.600 370.630 215.130 370.980 ;
        RECT 165.570 369.670 165.830 370.470 ;
        RECT 182.070 370.420 199.000 370.630 ;
        RECT 182.070 370.390 182.390 370.420 ;
        RECT 194.490 370.050 194.770 370.070 ;
        RECT 194.470 370.020 194.790 370.050 ;
        RECT 226.610 370.020 227.950 370.560 ;
        RECT 194.470 369.810 227.950 370.020 ;
        RECT 194.470 369.790 194.790 369.810 ;
        RECT 194.490 369.770 194.770 369.790 ;
        RECT 167.570 369.670 167.910 369.730 ;
        RECT 165.470 369.450 167.910 369.670 ;
        RECT 226.610 369.280 227.950 369.810 ;
        RECT 207.600 368.660 207.920 368.670 ;
        RECT 207.360 368.650 207.920 368.660 ;
        RECT 233.590 368.650 233.900 368.660 ;
        RECT 205.190 368.570 216.710 368.650 ;
        RECT 224.540 368.570 236.070 368.650 ;
        RECT 240.470 368.570 241.330 370.550 ;
        RECT 205.190 368.470 241.330 368.570 ;
        RECT 207.360 368.330 207.670 368.470 ;
        RECT 212.120 368.450 241.330 368.470 ;
        RECT 140.810 368.160 141.120 368.250 ;
        RECT 140.210 367.990 141.120 368.160 ;
        RECT 140.810 367.970 141.120 367.990 ;
        RECT 141.900 368.170 142.210 368.260 ;
        RECT 212.120 368.200 241.220 368.450 ;
        RECT 212.120 368.170 212.530 368.200 ;
        RECT 141.900 368.000 143.010 368.170 ;
        RECT 141.900 367.970 142.210 368.000 ;
        RECT 145.310 367.970 145.600 367.990 ;
        RECT 132.860 367.570 145.620 367.970 ;
        RECT 102.040 365.460 102.520 365.490 ;
        RECT 125.300 365.460 126.570 365.750 ;
        RECT 27.330 364.260 29.970 365.440 ;
        RECT 102.040 365.080 127.830 365.460 ;
        RECT 102.040 365.060 102.520 365.080 ;
        RECT 125.300 364.880 126.570 365.080 ;
        RECT 132.860 364.880 133.260 367.570 ;
        RECT 140.340 367.510 140.660 367.570 ;
        RECT 145.310 367.560 145.600 367.570 ;
        RECT 202.190 367.260 202.770 367.700 ;
        RECT 202.190 367.070 202.830 367.260 ;
        RECT 136.660 366.890 137.030 366.900 ;
        RECT 134.870 366.660 137.030 366.890 ;
        RECT 140.340 366.830 140.660 366.910 ;
        RECT 140.210 366.660 140.660 366.830 ;
        RECT 145.320 366.670 145.640 366.720 ;
        RECT 134.870 366.530 142.290 366.660 ;
        RECT 134.870 365.830 135.490 366.530 ;
        RECT 136.660 366.490 142.290 366.530 ;
        RECT 144.750 366.500 145.700 366.670 ;
        RECT 145.320 366.460 145.640 366.500 ;
        RECT 202.590 366.460 202.830 367.070 ;
        RECT 203.210 367.060 203.790 367.690 ;
        RECT 233.740 367.630 234.050 367.700 ;
        RECT 206.030 367.550 206.500 367.610 ;
        RECT 230.930 367.560 231.220 367.570 ;
        RECT 230.930 367.550 231.230 367.560 ;
        RECT 233.740 367.550 236.070 367.630 ;
        RECT 241.460 367.550 241.910 367.570 ;
        RECT 206.030 367.120 241.920 367.550 ;
        RECT 206.970 367.110 207.280 367.120 ;
        RECT 230.930 367.110 231.230 367.120 ;
        RECT 206.970 366.920 216.710 367.110 ;
        RECT 230.930 367.090 231.220 367.110 ;
        RECT 206.970 366.800 207.280 366.920 ;
        RECT 140.810 366.320 141.120 366.410 ;
        RECT 140.210 366.150 141.120 366.320 ;
        RECT 141.900 366.330 142.210 366.420 ;
        RECT 140.810 366.080 141.120 366.150 ;
        RECT 141.550 366.250 141.870 366.300 ;
        RECT 141.900 366.250 143.010 366.330 ;
        RECT 234.680 366.290 235.000 366.550 ;
        RECT 240.960 366.440 241.320 366.450 ;
        RECT 227.110 366.260 227.410 366.280 ;
        RECT 234.720 366.270 235.900 366.290 ;
        RECT 234.720 366.260 235.940 366.270 ;
        RECT 240.400 366.260 241.320 366.440 ;
        RECT 141.550 366.160 143.010 366.250 ;
        RECT 206.250 366.230 206.570 366.260 ;
        RECT 141.550 366.080 142.290 366.160 ;
        RECT 141.550 366.040 141.870 366.080 ;
        RECT 206.250 366.000 216.710 366.230 ;
        RECT 227.100 366.160 241.320 366.260 ;
        RECT 140.340 365.910 140.660 365.990 ;
        RECT 136.660 365.830 137.030 365.870 ;
        RECT 125.300 364.480 133.260 364.880 ;
        RECT 134.340 365.740 137.030 365.830 ;
        RECT 140.210 365.740 140.660 365.910 ;
        RECT 227.100 365.840 241.360 366.160 ;
        RECT 227.110 365.820 227.410 365.840 ;
        RECT 145.320 365.750 145.640 365.800 ;
        RECT 134.340 365.570 142.290 365.740 ;
        RECT 144.750 365.580 145.700 365.750 ;
        RECT 234.680 365.690 235.000 365.840 ;
        RECT 134.340 365.460 137.030 365.570 ;
        RECT 145.320 365.540 145.640 365.580 ;
        RECT 240.400 365.500 241.360 365.840 ;
        RECT 134.340 365.350 135.490 365.460 ;
        RECT 134.340 364.900 135.450 365.350 ;
        RECT 140.620 365.320 140.930 365.430 ;
        RECT 140.210 365.130 140.930 365.320 ;
        RECT 140.620 365.100 140.930 365.130 ;
        RECT 141.520 365.330 141.840 365.380 ;
        RECT 141.520 365.260 142.290 365.330 ;
        RECT 141.520 365.160 143.010 365.260 ;
        RECT 141.520 365.120 141.840 365.160 ;
        RECT 141.920 365.060 143.010 365.160 ;
        RECT 206.960 365.250 207.270 365.440 ;
        RECT 231.500 365.330 232.620 365.340 ;
        RECT 209.340 365.250 209.660 365.310 ;
        RECT 206.960 365.190 216.710 365.250 ;
        RECT 230.630 365.190 234.150 365.330 ;
        RECT 206.960 365.130 234.150 365.190 ;
        RECT 206.960 365.120 232.620 365.130 ;
        RECT 206.960 365.110 231.930 365.120 ;
        RECT 206.990 365.060 231.930 365.110 ;
        RECT 141.920 365.000 142.230 365.060 ;
        RECT 209.340 365.010 231.930 365.060 ;
        RECT 232.270 365.000 232.580 365.120 ;
        RECT 232.710 365.060 233.660 365.130 ;
        RECT 233.350 364.990 233.660 365.060 ;
        RECT 233.840 365.000 234.150 365.130 ;
        RECT 234.320 364.990 234.630 365.040 ;
        RECT 236.570 364.990 236.880 365.090 ;
        RECT 136.660 364.900 137.030 364.940 ;
        RECT 140.620 364.900 140.940 364.960 ;
        RECT 134.340 364.820 137.030 364.900 ;
        RECT 140.210 364.820 140.940 364.900 ;
        RECT 145.290 364.830 145.610 364.880 ;
        RECT 233.740 364.870 234.050 364.940 ;
        RECT 234.320 364.870 236.880 364.990 ;
        RECT 134.340 364.650 142.290 364.820 ;
        RECT 144.750 364.660 145.700 364.830 ;
        RECT 233.740 364.760 236.880 364.870 ;
        RECT 233.740 364.660 236.070 364.760 ;
        RECT 134.340 364.530 137.030 364.650 ;
        RECT 140.620 364.640 140.940 364.650 ;
        RECT 145.290 364.620 145.610 364.660 ;
        RECT 233.740 364.610 234.050 364.660 ;
        RECT 134.340 364.490 135.240 364.530 ;
        RECT 125.300 364.260 126.570 364.480 ;
        RECT 27.250 362.010 127.560 364.260 ;
        RECT 15.100 359.920 17.990 361.880 ;
        RECT 27.330 361.840 29.970 362.010 ;
        RECT 102.040 360.690 102.580 360.720 ;
        RECT 125.730 360.690 127.000 360.820 ;
        RECT 102.040 360.280 127.470 360.690 ;
        RECT 102.040 360.240 102.580 360.280 ;
        RECT 125.730 359.940 127.000 360.280 ;
        RECT 134.340 359.940 134.710 364.490 ;
        RECT 140.620 364.360 140.930 364.470 ;
        RECT 140.210 364.170 140.930 364.360 ;
        RECT 141.530 364.410 141.850 364.460 ;
        RECT 233.500 364.450 233.810 364.490 ;
        RECT 141.530 364.300 142.290 364.410 ;
        RECT 233.320 364.390 234.040 364.450 ;
        RECT 233.190 364.350 234.040 364.390 ;
        RECT 234.270 364.380 234.580 364.390 ;
        RECT 234.200 364.350 234.580 364.380 ;
        RECT 141.530 364.240 143.010 364.300 ;
        RECT 141.530 364.200 141.850 364.240 ;
        RECT 140.620 364.140 140.930 364.170 ;
        RECT 141.920 364.100 143.010 364.240 ;
        RECT 141.920 364.040 142.230 364.100 ;
        RECT 212.490 364.020 221.640 364.250 ;
        RECT 230.630 364.150 231.240 364.350 ;
        RECT 233.140 364.150 235.390 364.350 ;
        RECT 230.920 364.060 231.240 364.150 ;
        RECT 233.190 364.130 233.510 364.150 ;
        RECT 233.770 364.100 234.580 364.150 ;
        RECT 233.770 364.090 234.040 364.100 ;
        RECT 234.270 364.060 234.580 364.100 ;
        RECT 240.460 364.070 241.360 365.500 ;
        RECT 140.620 363.940 140.940 364.000 ;
        RECT 140.210 363.820 140.940 363.940 ;
        RECT 221.350 363.920 221.640 364.020 ;
        RECT 135.820 363.800 142.310 363.820 ;
        RECT 125.730 359.920 134.710 359.940 ;
        RECT 15.070 359.570 134.710 359.920 ;
        RECT 135.530 363.630 142.310 363.800 ;
        RECT 221.350 363.770 230.470 363.920 ;
        RECT 232.380 363.810 232.690 363.950 ;
        RECT 230.920 363.770 231.240 363.790 ;
        RECT 232.030 363.770 232.690 363.810 ;
        RECT 233.590 363.780 233.900 363.920 ;
        RECT 233.590 363.770 236.070 363.780 ;
        RECT 221.350 363.720 236.070 363.770 ;
        RECT 221.350 363.710 221.640 363.720 ;
        RECT 135.530 363.450 137.030 363.630 ;
        RECT 224.540 363.620 236.070 363.720 ;
        RECT 135.530 362.860 136.190 363.450 ;
        RECT 136.660 363.410 137.030 363.450 ;
        RECT 140.620 363.440 140.930 363.510 ;
        RECT 230.630 363.500 231.240 363.620 ;
        RECT 232.030 363.590 232.380 363.620 ;
        RECT 233.140 363.600 236.070 363.620 ;
        RECT 233.140 363.500 235.390 363.600 ;
        RECT 233.190 363.460 233.510 363.500 ;
        RECT 233.840 363.440 234.580 363.500 ;
        RECT 140.620 363.400 141.200 363.440 ;
        RECT 233.550 363.420 234.580 363.440 ;
        RECT 141.920 363.400 142.230 363.410 ;
        RECT 140.210 363.340 142.310 363.400 ;
        RECT 140.210 363.210 143.010 363.340 ;
        RECT 140.620 363.180 141.200 363.210 ;
        RECT 141.920 363.140 143.010 363.210 ;
        RECT 212.490 363.300 220.700 363.420 ;
        RECT 233.500 363.300 234.580 363.420 ;
        RECT 212.490 363.200 228.640 363.300 ;
        RECT 141.920 363.080 142.230 363.140 ;
        RECT 220.480 363.100 228.640 363.200 ;
        RECT 233.500 363.180 234.060 363.300 ;
        RECT 234.270 363.220 234.580 363.300 ;
        RECT 233.500 363.170 233.970 363.180 ;
        RECT 140.620 362.980 140.940 363.040 ;
        RECT 140.210 362.860 140.940 362.980 ;
        RECT 135.530 362.670 142.310 362.860 ;
        RECT 135.530 362.490 137.030 362.670 ;
        RECT 135.530 362.480 136.200 362.490 ;
        RECT 135.530 362.440 136.190 362.480 ;
        RECT 136.660 362.450 137.030 362.490 ;
        RECT 140.840 362.440 141.160 362.480 ;
        RECT 15.070 358.060 127.190 359.570 ;
        RECT 125.670 355.480 126.940 356.070 ;
        RECT 23.960 355.180 127.480 355.480 ;
        RECT 135.530 355.180 135.900 362.440 ;
        RECT 140.840 362.250 142.310 362.440 ;
        RECT 220.480 362.420 220.700 363.100 ;
        RECT 223.100 362.940 223.560 363.070 ;
        RECT 228.420 362.940 228.640 363.100 ;
        RECT 223.100 362.740 230.470 362.940 ;
        RECT 234.320 362.850 234.630 362.900 ;
        RECT 234.830 362.850 236.540 362.940 ;
        RECT 236.620 362.850 236.930 362.870 ;
        RECT 223.100 362.620 223.560 362.740 ;
        RECT 228.420 362.620 228.640 362.740 ;
        RECT 232.270 362.730 232.580 362.850 ;
        RECT 231.500 362.720 232.620 362.730 ;
        RECT 233.840 362.720 234.150 362.850 ;
        RECT 230.630 362.620 234.150 362.720 ;
        RECT 234.320 362.620 237.240 362.850 ;
        RECT 224.540 362.440 236.070 362.620 ;
        RECT 227.240 362.420 227.460 362.430 ;
        RECT 220.480 362.290 227.490 362.420 ;
        RECT 228.420 362.380 228.640 362.440 ;
        RECT 232.790 362.390 233.900 362.440 ;
        RECT 228.390 362.340 228.640 362.380 ;
        RECT 233.110 362.340 233.420 362.390 ;
        RECT 228.390 362.290 228.650 362.340 ;
        RECT 231.500 362.310 232.620 362.320 ;
        RECT 233.590 362.310 233.900 362.390 ;
        RECT 140.840 362.220 141.160 362.250 ;
        RECT 220.480 362.170 230.470 362.290 ;
        RECT 214.470 362.030 214.780 362.080 ;
        RECT 214.470 362.020 214.930 362.030 ;
        RECT 214.470 361.840 216.720 362.020 ;
        RECT 214.470 361.750 214.780 361.840 ;
        RECT 140.880 361.480 141.200 361.520 ;
        RECT 140.880 361.290 142.310 361.480 ;
        RECT 220.480 361.440 220.700 362.170 ;
        RECT 224.110 362.090 230.470 362.170 ;
        RECT 230.630 362.110 234.150 362.310 ;
        RECT 236.340 362.290 236.540 362.620 ;
        RECT 236.620 362.540 236.930 362.620 ;
        RECT 231.500 362.100 232.620 362.110 ;
        RECT 224.110 361.970 224.470 362.090 ;
        RECT 220.480 361.310 224.170 361.440 ;
        RECT 227.200 361.310 227.490 362.090 ;
        RECT 228.390 361.700 228.650 362.090 ;
        RECT 232.270 361.980 232.580 362.100 ;
        RECT 233.840 361.980 234.150 362.110 ;
        RECT 234.830 362.090 236.540 362.290 ;
        RECT 234.320 362.020 234.630 362.080 ;
        RECT 236.340 362.020 236.540 362.090 ;
        RECT 236.610 362.020 236.920 362.150 ;
        RECT 234.320 361.800 237.240 362.020 ;
        RECT 234.320 361.750 234.630 361.800 ;
        RECT 228.390 361.490 232.520 361.700 ;
        RECT 232.310 361.350 232.520 361.490 ;
        RECT 233.740 361.600 234.050 361.670 ;
        RECT 233.740 361.380 236.070 361.600 ;
        RECT 233.190 361.350 233.510 361.370 ;
        RECT 233.740 361.350 234.050 361.380 ;
        RECT 234.270 361.360 234.580 361.380 ;
        RECT 234.200 361.350 234.580 361.360 ;
        RECT 232.310 361.330 234.580 361.350 ;
        RECT 140.880 361.260 141.200 361.290 ;
        RECT 220.480 361.110 230.470 361.310 ;
        RECT 230.630 361.130 231.240 361.330 ;
        RECT 232.310 361.140 235.390 361.330 ;
        RECT 233.140 361.130 235.390 361.140 ;
        RECT 220.480 361.100 222.080 361.110 ;
        RECT 185.200 361.010 185.510 361.020 ;
        RECT 185.190 360.950 185.520 361.010 ;
        RECT 184.840 360.900 185.520 360.950 ;
        RECT 181.610 360.820 185.520 360.900 ;
        RECT 186.840 360.870 188.790 361.010 ;
        RECT 223.940 360.900 224.170 361.110 ;
        RECT 227.200 361.000 227.490 361.110 ;
        RECT 230.920 361.040 231.240 361.130 ;
        RECT 233.190 361.110 233.510 361.130 ;
        RECT 234.200 361.100 234.580 361.130 ;
        RECT 236.340 361.040 236.540 361.800 ;
        RECT 240.430 361.040 241.330 361.710 ;
        RECT 227.200 360.900 230.090 361.000 ;
        RECT 186.770 360.850 188.790 360.870 ;
        RECT 186.770 360.820 187.090 360.850 ;
        RECT 187.570 360.840 188.790 360.850 ;
        RECT 188.270 360.830 188.790 360.840 ;
        RECT 181.610 360.680 187.090 360.820 ;
        RECT 212.490 360.700 230.470 360.900 ;
        RECT 184.360 360.630 187.090 360.680 ;
        RECT 184.360 360.580 184.680 360.630 ;
        RECT 186.770 360.610 187.090 360.630 ;
        RECT 223.940 360.650 224.170 360.700 ;
        RECT 230.920 360.680 231.240 360.770 ;
        RECT 233.190 360.680 233.510 360.700 ;
        RECT 234.200 360.680 234.520 360.710 ;
        RECT 223.940 360.500 224.160 360.650 ;
        RECT 230.630 360.550 231.240 360.680 ;
        RECT 233.140 360.550 235.390 360.680 ;
        RECT 228.310 360.500 235.390 360.550 ;
        RECT 223.940 360.480 235.390 360.500 ;
        RECT 236.340 360.610 241.330 361.040 ;
        RECT 223.940 360.340 234.580 360.480 ;
        RECT 223.940 360.280 228.700 360.340 ;
        RECT 234.270 360.260 234.580 360.340 ;
        RECT 234.680 360.260 235.000 360.480 ;
        RECT 234.720 360.240 235.900 360.260 ;
        RECT 225.030 360.030 225.420 360.050 ;
        RECT 225.020 359.920 225.430 360.030 ;
        RECT 234.720 359.980 235.940 360.240 ;
        RECT 225.020 359.720 230.470 359.920 ;
        RECT 234.320 359.860 234.630 359.940 ;
        RECT 234.720 359.920 235.900 359.980 ;
        RECT 236.340 359.920 236.540 360.610 ;
        RECT 234.680 359.900 236.540 359.920 ;
        RECT 234.680 359.860 236.840 359.900 ;
        RECT 225.020 359.630 225.430 359.720 ;
        RECT 232.270 359.710 232.580 359.830 ;
        RECT 233.840 359.780 234.150 359.830 ;
        RECT 231.500 359.700 232.620 359.710 ;
        RECT 233.750 359.700 234.150 359.780 ;
        RECT 230.630 359.630 234.150 359.700 ;
        RECT 217.560 359.500 234.150 359.630 ;
        RECT 234.320 359.630 237.030 359.860 ;
        RECT 234.320 359.610 234.630 359.630 ;
        RECT 236.340 359.570 236.840 359.630 ;
        RECT 240.430 359.620 241.330 360.610 ;
        RECT 217.560 359.480 234.070 359.500 ;
        RECT 217.560 359.330 217.880 359.480 ;
        RECT 223.360 359.330 223.680 359.480 ;
        RECT 225.850 359.330 226.250 359.340 ;
        RECT 225.830 359.270 226.270 359.330 ;
        RECT 233.350 359.280 233.660 359.290 ;
        RECT 232.780 359.270 233.660 359.280 ;
        RECT 236.340 359.270 236.540 359.570 ;
        RECT 209.390 359.130 209.710 359.250 ;
        RECT 225.830 359.130 230.470 359.270 ;
        RECT 231.590 359.130 231.910 359.250 ;
        RECT 209.390 358.950 231.910 359.130 ;
        RECT 232.710 359.030 233.660 359.270 ;
        RECT 234.830 359.150 236.540 359.270 ;
        RECT 234.830 359.070 236.510 359.150 ;
        RECT 233.350 358.960 233.660 359.030 ;
        RECT 234.320 358.960 234.630 359.010 ;
        RECT 236.570 358.960 236.880 359.060 ;
        RECT 233.740 358.840 234.050 358.910 ;
        RECT 234.320 358.840 236.880 358.960 ;
        RECT 233.740 358.730 236.880 358.840 ;
        RECT 233.740 358.630 236.070 358.730 ;
        RECT 233.740 358.580 234.050 358.630 ;
        RECT 233.500 358.420 233.810 358.460 ;
        RECT 214.500 358.310 214.810 358.390 ;
        RECT 214.500 358.290 216.720 358.310 ;
        RECT 212.490 358.090 230.470 358.290 ;
        RECT 233.320 358.280 234.040 358.420 ;
        RECT 234.270 358.280 234.580 358.360 ;
        RECT 233.320 358.170 234.580 358.280 ;
        RECT 233.500 358.130 234.580 358.170 ;
        RECT 214.500 358.060 214.810 358.090 ;
        RECT 218.050 358.020 218.890 358.090 ;
        RECT 233.770 358.070 234.580 358.130 ;
        RECT 233.770 358.060 234.040 358.070 ;
        RECT 234.270 358.030 234.580 358.070 ;
        RECT 232.380 357.780 232.690 357.920 ;
        RECT 218.500 357.740 228.640 357.770 ;
        RECT 232.030 357.740 232.690 357.780 ;
        RECT 233.590 357.750 233.900 357.890 ;
        RECT 233.590 357.740 236.070 357.750 ;
        RECT 218.500 357.590 236.070 357.740 ;
        RECT 218.500 357.550 228.640 357.590 ;
        RECT 232.030 357.560 232.380 357.590 ;
        RECT 233.590 357.570 236.070 357.590 ;
        RECT 233.590 357.560 233.900 357.570 ;
        RECT 228.420 356.350 228.640 357.550 ;
        RECT 233.840 357.490 234.040 357.500 ;
        RECT 233.840 357.480 234.060 357.490 ;
        RECT 234.270 357.480 234.580 357.520 ;
        RECT 233.840 357.410 234.580 357.480 ;
        RECT 233.550 357.390 234.580 357.410 ;
        RECT 233.500 357.270 234.580 357.390 ;
        RECT 233.500 357.150 234.060 357.270 ;
        RECT 234.270 357.190 234.580 357.270 ;
        RECT 233.500 357.140 233.970 357.150 ;
        RECT 228.390 356.310 228.640 356.350 ;
        RECT 217.630 356.140 217.950 356.190 ;
        RECT 217.630 355.890 223.650 356.140 ;
        RECT 223.330 355.820 223.650 355.890 ;
        RECT 228.390 355.670 228.650 356.310 ;
        RECT 228.390 355.460 232.520 355.670 ;
        RECT 23.960 354.810 135.900 355.180 ;
        RECT 232.310 355.320 232.520 355.460 ;
        RECT 237.690 355.410 238.470 355.560 ;
        RECT 240.430 355.410 241.330 356.330 ;
        RECT 234.270 355.320 234.580 355.400 ;
        RECT 232.310 355.110 234.580 355.320 ;
        RECT 234.270 355.070 234.580 355.110 ;
        RECT 237.690 354.940 241.330 355.410 ;
        RECT 23.960 353.400 127.480 354.810 ;
        RECT 237.690 354.790 238.470 354.940 ;
        RECT 181.840 354.390 182.160 354.400 ;
        RECT 209.650 354.390 210.110 354.460 ;
        RECT 181.840 354.110 210.110 354.390 ;
        RECT 240.430 354.240 241.330 354.940 ;
        RECT 181.840 354.060 182.160 354.110 ;
        RECT 209.650 354.050 210.110 354.110 ;
        RECT 223.330 353.600 223.650 353.610 ;
        RECT 233.770 353.600 234.100 353.740 ;
        RECT 223.330 353.440 234.100 353.600 ;
        RECT 223.330 353.430 224.020 353.440 ;
        RECT 23.960 333.290 26.040 353.400 ;
        RECT 192.670 353.270 192.980 353.290 ;
        RECT 193.350 353.270 196.200 353.350 ;
        RECT 210.240 353.270 213.070 353.350 ;
        RECT 223.330 353.310 223.650 353.430 ;
        RECT 213.440 353.270 213.750 353.290 ;
        RECT 190.510 353.250 200.570 353.270 ;
        RECT 205.850 353.250 215.910 353.270 ;
        RECT 190.510 353.100 215.910 353.250 ;
        RECT 190.510 353.090 193.070 353.100 ;
        RECT 192.670 352.960 192.980 353.090 ;
        RECT 193.350 353.050 193.770 353.100 ;
        RECT 195.760 353.070 210.440 353.100 ;
        RECT 212.750 353.050 213.070 353.100 ;
        RECT 213.350 353.090 215.910 353.100 ;
        RECT 213.440 352.960 213.750 353.090 ;
        RECT 193.580 352.720 193.900 352.800 ;
        RECT 197.510 352.720 197.830 352.730 ;
        RECT 193.580 352.540 197.830 352.720 ;
        RECT 193.580 352.480 193.900 352.540 ;
        RECT 197.510 352.470 197.830 352.540 ;
        RECT 208.590 352.720 208.910 352.730 ;
        RECT 212.520 352.720 212.840 352.800 ;
        RECT 208.590 352.540 212.840 352.720 ;
        RECT 208.590 352.470 208.910 352.540 ;
        RECT 212.520 352.480 212.840 352.540 ;
        RECT 363.620 351.550 365.020 377.510 ;
        RECT 367.750 373.190 369.030 378.410 ;
        RECT 368.270 372.450 369.030 373.190 ;
        RECT 369.920 353.470 371.320 380.660 ;
        RECT 369.910 352.960 371.320 353.470 ;
        RECT 368.800 352.790 371.320 352.960 ;
        RECT 369.910 352.540 371.320 352.790 ;
        RECT 363.490 351.470 365.020 351.550 ;
        RECT 217.710 350.420 218.310 350.480 ;
        RECT 240.430 350.420 241.330 351.450 ;
        RECT 217.710 349.950 241.330 350.420 ;
        RECT 217.710 349.900 218.310 349.950 ;
        RECT 240.430 349.360 241.330 349.950 ;
        RECT 362.980 350.460 365.020 351.470 ;
        RECT 362.980 349.820 368.030 350.460 ;
        RECT 362.980 349.540 365.020 349.820 ;
        RECT 362.910 348.920 365.020 349.540 ;
        RECT 193.250 347.320 193.560 347.460 ;
        RECT 191.090 347.140 193.660 347.320 ;
        RECT 193.250 347.130 193.560 347.140 ;
        RECT 193.250 346.890 193.560 346.910 ;
        RECT 191.090 346.710 201.170 346.890 ;
        RECT 193.250 346.580 193.560 346.710 ;
        RECT 201.020 346.700 201.170 346.710 ;
        RECT 140.840 346.450 141.150 346.470 ;
        RECT 141.500 346.450 141.810 346.470 ;
        RECT 140.840 345.980 148.160 346.450 ;
        RECT 140.840 345.960 141.150 345.980 ;
        RECT 141.500 345.960 141.810 345.980 ;
        RECT 147.690 345.300 148.160 345.980 ;
        RECT 174.460 346.310 174.770 346.330 ;
        RECT 212.100 346.310 212.550 346.340 ;
        RECT 174.460 345.900 212.550 346.310 ;
        RECT 174.460 345.880 174.770 345.900 ;
        RECT 193.250 345.890 193.560 345.900 ;
        RECT 201.050 345.890 201.190 345.900 ;
        RECT 191.080 345.710 201.190 345.890 ;
        RECT 212.100 345.880 212.550 345.900 ;
        RECT 193.250 345.690 193.560 345.710 ;
        RECT 193.250 345.460 193.560 345.470 ;
        RECT 191.090 345.420 193.560 345.460 ;
        RECT 191.090 345.300 193.650 345.420 ;
        RECT 240.460 345.300 241.360 346.270 ;
        RECT 139.510 345.170 139.770 345.240 ;
        RECT 141.560 345.170 141.880 345.190 ;
        RECT 143.320 345.170 143.650 345.210 ;
        RECT 139.510 344.980 143.650 345.170 ;
        RECT 139.510 344.920 139.770 344.980 ;
        RECT 141.560 344.930 141.880 344.980 ;
        RECT 143.320 344.940 143.650 344.980 ;
        RECT 147.690 344.830 241.360 345.300 ;
        RECT 138.960 344.770 139.280 344.810 ;
        RECT 140.900 344.770 141.220 344.830 ;
        RECT 143.820 344.770 144.140 344.810 ;
        RECT 138.960 344.580 144.140 344.770 ;
        RECT 216.620 344.710 217.190 344.830 ;
        RECT 138.960 344.550 139.280 344.580 ;
        RECT 140.900 344.570 141.220 344.580 ;
        RECT 143.820 344.550 144.140 344.580 ;
        RECT 142.300 344.190 142.610 344.260 ;
        RECT 145.300 344.210 145.600 344.230 ;
        RECT 145.290 344.190 145.610 344.210 ;
        RECT 142.300 343.980 145.610 344.190 ;
        RECT 240.460 344.180 241.360 344.830 ;
        RECT 142.300 343.930 142.610 343.980 ;
        RECT 143.070 343.970 145.610 343.980 ;
        RECT 141.130 343.750 141.440 343.820 ;
        RECT 143.070 343.750 143.290 343.970 ;
        RECT 145.290 343.950 145.610 343.970 ;
        RECT 145.300 343.930 145.600 343.950 ;
        RECT 141.130 343.530 143.290 343.750 ;
        RECT 141.130 343.490 141.440 343.530 ;
        RECT 142.810 343.030 143.130 343.090 ;
        RECT 144.680 343.060 144.970 343.080 ;
        RECT 142.810 343.020 143.290 343.030 ;
        RECT 144.670 343.020 144.990 343.060 ;
        RECT 142.810 342.830 144.990 343.020 ;
        RECT 142.810 342.820 143.290 342.830 ;
        RECT 142.810 342.770 143.130 342.820 ;
        RECT 144.670 342.800 144.990 342.830 ;
        RECT 144.680 342.780 144.970 342.800 ;
        RECT 139.980 342.420 140.300 342.440 ;
        RECT 139.760 342.200 140.300 342.420 ;
        RECT 139.980 342.180 140.300 342.200 ;
        RECT 142.730 341.840 143.050 341.960 ;
        RECT 139.760 341.640 143.050 341.840 ;
        RECT 139.760 341.630 142.740 341.640 ;
        RECT 139.760 341.420 142.740 341.440 ;
        RECT 139.760 341.230 143.060 341.420 ;
        RECT 142.740 341.100 143.060 341.230 ;
        RECT 138.990 340.900 139.280 340.910 ;
        RECT 138.980 340.880 139.300 340.900 ;
        RECT 139.980 340.880 140.300 340.890 ;
        RECT 138.980 340.660 140.300 340.880 ;
        RECT 138.980 340.640 139.300 340.660 ;
        RECT 138.990 340.620 139.280 340.640 ;
        RECT 139.980 340.630 140.300 340.660 ;
        RECT 142.790 340.420 143.110 340.470 ;
        RECT 144.250 340.420 144.570 340.470 ;
        RECT 142.790 340.210 144.570 340.420 ;
        RECT 142.790 340.150 143.110 340.210 ;
        RECT 144.250 340.170 144.570 340.210 ;
        RECT 215.500 340.060 216.050 340.070 ;
        RECT 215.500 340.040 216.060 340.060 ;
        RECT 240.430 340.040 241.330 341.190 ;
        RECT 215.500 339.570 241.330 340.040 ;
        RECT 215.500 339.560 216.060 339.570 ;
        RECT 215.500 339.540 216.050 339.560 ;
        RECT 240.430 339.100 241.330 339.570 ;
        RECT 140.090 337.840 140.400 337.850 ;
        RECT 141.180 337.840 141.490 337.850 ;
        RECT 138.770 337.830 141.490 337.840 ;
        RECT 138.540 337.520 141.490 337.830 ;
        RECT 138.540 337.510 141.480 337.520 ;
        RECT 41.350 335.890 127.960 336.820 ;
        RECT 138.540 335.890 138.890 337.510 ;
        RECT 165.470 337.450 167.910 337.670 ;
        RECT 139.540 337.160 139.850 337.170 ;
        RECT 140.640 337.160 140.950 337.170 ;
        RECT 141.740 337.160 142.050 337.170 ;
        RECT 139.510 336.840 142.670 337.160 ;
        RECT 142.350 335.890 142.670 336.840 ;
        RECT 165.570 336.650 165.830 337.450 ;
        RECT 167.570 337.390 167.910 337.450 ;
        RECT 220.690 337.230 221.250 337.300 ;
        RECT 233.410 337.230 234.090 337.290 ;
        RECT 240.940 337.230 241.600 337.870 ;
        RECT 171.750 336.970 172.080 336.990 ;
        RECT 171.740 336.890 172.090 336.970 ;
        RECT 177.490 336.890 177.810 336.950 ;
        RECT 170.400 336.830 170.720 336.840 ;
        RECT 171.740 336.830 177.810 336.890 ;
        RECT 170.400 336.730 177.810 336.830 ;
        RECT 220.690 336.820 241.600 337.230 ;
        RECT 220.690 336.770 221.250 336.820 ;
        RECT 233.410 336.760 234.090 336.820 ;
        RECT 170.400 336.660 172.090 336.730 ;
        RECT 177.490 336.680 177.810 336.730 ;
        RECT 240.940 336.720 241.600 336.820 ;
        RECT 170.400 336.630 172.030 336.660 ;
        RECT 170.400 336.580 170.720 336.630 ;
        RECT 167.320 336.270 167.650 336.510 ;
        RECT 171.800 336.270 171.910 336.430 ;
        RECT 173.180 336.400 173.480 336.410 ;
        RECT 173.170 336.270 173.490 336.400 ;
        RECT 183.710 336.270 183.990 336.570 ;
        RECT 187.740 336.270 188.040 336.550 ;
        RECT 167.320 336.250 188.040 336.270 ;
        RECT 167.320 336.220 188.030 336.250 ;
        RECT 167.320 336.110 187.970 336.220 ;
        RECT 171.130 335.890 171.570 335.900 ;
        RECT 41.350 335.880 171.570 335.890 ;
        RECT 41.350 335.470 171.590 335.880 ;
        RECT 41.350 334.920 127.960 335.470 ;
        RECT 138.540 335.070 138.890 335.470 ;
        RECT 138.540 334.920 141.490 335.070 ;
        RECT 142.350 334.920 142.670 335.470 ;
        RECT 164.280 335.460 164.760 335.470 ;
        RECT 171.110 335.460 171.590 335.470 ;
        RECT 171.130 335.450 171.570 335.460 ;
        RECT 41.350 334.740 167.770 334.920 ;
        RECT 23.890 329.920 26.230 333.290 ;
        RECT 23.960 329.050 26.040 329.920 ;
        RECT 41.350 218.980 43.430 334.740 ;
        RECT 125.790 334.500 167.770 334.740 ;
        RECT 214.450 334.740 215.050 334.790 ;
        RECT 240.860 334.740 242.960 335.680 ;
        RECT 138.540 333.870 138.890 334.500 ;
        RECT 138.540 333.740 138.920 333.870 ;
        RECT 138.540 333.700 139.290 333.740 ;
        RECT 140.090 333.700 140.400 333.720 ;
        RECT 138.540 333.400 141.490 333.700 ;
        RECT 140.090 333.390 140.400 333.400 ;
        RECT 141.180 333.370 141.490 333.400 ;
        RECT 139.540 333.020 139.850 333.030 ;
        RECT 142.350 333.020 142.670 334.500 ;
        RECT 148.840 334.000 149.670 334.500 ;
        RECT 214.450 334.270 242.960 334.740 ;
        RECT 214.450 334.230 215.050 334.270 ;
        RECT 240.860 333.600 242.960 334.270 ;
        RECT 240.880 333.590 241.650 333.600 ;
        RECT 139.520 332.690 142.670 333.020 ;
        RECT 139.520 332.680 142.580 332.690 ;
        RECT 142.430 332.480 142.720 332.500 ;
        RECT 144.660 332.480 144.970 332.500 ;
        RECT 142.420 332.120 144.970 332.480 ;
        RECT 142.430 332.100 142.720 332.120 ;
        RECT 144.660 332.100 144.970 332.120 ;
        RECT 181.960 331.610 185.020 331.620 ;
        RECT 172.150 331.580 175.210 331.590 ;
        RECT 172.060 331.250 175.210 331.580 ;
        RECT 177.490 331.580 180.550 331.590 ;
        RECT 177.490 331.250 180.640 331.580 ;
        RECT 139.380 330.280 139.690 330.290 ;
        RECT 140.470 330.280 140.780 330.290 ;
        RECT 138.060 330.270 140.780 330.280 ;
        RECT 137.830 329.960 140.780 330.270 ;
        RECT 137.830 329.950 140.770 329.960 ;
        RECT 136.620 329.520 136.990 329.530 ;
        RECT 137.830 329.520 138.180 329.950 ;
        RECT 138.830 329.600 139.140 329.610 ;
        RECT 139.930 329.600 140.240 329.610 ;
        RECT 141.030 329.600 141.340 329.610 ;
        RECT 125.730 328.700 127.000 329.400 ;
        RECT 135.300 329.140 138.180 329.520 ;
        RECT 138.800 329.280 141.960 329.600 ;
        RECT 135.300 328.700 135.680 329.140 ;
        RECT 136.620 329.120 136.990 329.140 ;
        RECT 125.730 328.600 135.680 328.700 ;
        RECT 49.850 328.320 135.680 328.600 ;
        RECT 49.850 326.520 127.960 328.320 ;
        RECT 137.830 327.510 138.180 329.140 ;
        RECT 141.640 328.820 141.960 329.280 ;
        RECT 172.060 329.160 172.380 331.250 ;
        RECT 174.880 331.240 175.190 331.250 ;
        RECT 177.510 331.240 177.820 331.250 ;
        RECT 173.240 330.870 173.550 330.900 ;
        RECT 174.330 330.870 174.640 330.880 ;
        RECT 178.060 330.870 178.370 330.880 ;
        RECT 179.150 330.870 179.460 330.900 ;
        RECT 173.240 330.570 176.190 330.870 ;
        RECT 174.330 330.550 174.640 330.570 ;
        RECT 175.440 330.530 176.190 330.570 ;
        RECT 175.810 330.400 176.190 330.530 ;
        RECT 175.840 329.970 176.190 330.400 ;
        RECT 176.510 330.570 179.460 330.870 ;
        RECT 176.510 330.530 177.260 330.570 ;
        RECT 178.060 330.550 178.370 330.570 ;
        RECT 176.510 330.400 176.890 330.530 ;
        RECT 176.510 329.970 176.860 330.400 ;
        RECT 180.320 329.970 180.640 331.250 ;
        RECT 181.870 331.280 185.020 331.610 ;
        RECT 187.300 331.610 190.360 331.620 ;
        RECT 187.300 331.280 190.450 331.610 ;
        RECT 181.870 329.970 182.190 331.280 ;
        RECT 184.690 331.270 185.000 331.280 ;
        RECT 187.320 331.270 187.630 331.280 ;
        RECT 183.050 330.900 183.360 330.930 ;
        RECT 184.140 330.900 184.450 330.910 ;
        RECT 187.870 330.900 188.180 330.910 ;
        RECT 188.960 330.900 189.270 330.930 ;
        RECT 183.050 330.600 186.000 330.900 ;
        RECT 184.140 330.580 184.450 330.600 ;
        RECT 185.250 330.560 186.000 330.600 ;
        RECT 185.620 330.430 186.000 330.560 ;
        RECT 185.650 329.970 186.000 330.430 ;
        RECT 186.320 330.600 189.270 330.900 ;
        RECT 186.320 330.560 187.070 330.600 ;
        RECT 187.870 330.580 188.180 330.600 ;
        RECT 186.320 330.430 186.700 330.560 ;
        RECT 186.320 329.970 186.670 330.430 ;
        RECT 175.820 329.940 186.720 329.970 ;
        RECT 175.810 329.690 186.720 329.940 ;
        RECT 175.810 329.660 176.190 329.690 ;
        RECT 175.840 329.530 176.190 329.660 ;
        RECT 173.240 329.200 176.190 329.530 ;
        RECT 171.890 329.150 172.390 329.160 ;
        RECT 175.840 329.150 176.190 329.200 ;
        RECT 176.510 329.680 176.890 329.690 ;
        RECT 176.510 329.530 176.860 329.680 ;
        RECT 176.510 329.200 179.460 329.530 ;
        RECT 176.510 329.150 176.860 329.200 ;
        RECT 180.320 329.150 180.640 329.690 ;
        RECT 181.870 329.150 182.190 329.690 ;
        RECT 185.620 329.660 186.000 329.690 ;
        RECT 185.650 329.560 186.000 329.660 ;
        RECT 183.050 329.230 186.000 329.560 ;
        RECT 185.650 329.150 186.000 329.230 ;
        RECT 186.320 329.560 186.670 329.690 ;
        RECT 186.320 329.230 189.270 329.560 ;
        RECT 186.320 329.150 186.670 329.230 ;
        RECT 190.130 329.150 190.450 331.280 ;
        RECT 193.790 331.590 196.850 331.600 ;
        RECT 193.790 331.260 196.940 331.590 ;
        RECT 193.810 331.250 194.120 331.260 ;
        RECT 194.360 330.880 194.670 330.890 ;
        RECT 195.450 330.880 195.760 330.910 ;
        RECT 192.810 330.580 195.760 330.880 ;
        RECT 192.810 330.540 193.560 330.580 ;
        RECT 194.360 330.560 194.670 330.580 ;
        RECT 192.810 330.410 193.190 330.540 ;
        RECT 192.810 329.540 193.160 330.410 ;
        RECT 192.810 329.210 195.760 329.540 ;
        RECT 192.810 329.150 193.160 329.210 ;
        RECT 196.620 329.150 196.940 331.260 ;
        RECT 217.820 329.150 218.380 329.170 ;
        RECT 145.290 328.820 145.570 328.830 ;
        RECT 141.640 328.490 145.590 328.820 ;
        RECT 171.890 328.690 218.380 329.150 ;
        RECT 171.890 328.610 175.220 328.690 ;
        RECT 141.640 328.240 141.960 328.490 ;
        RECT 145.290 328.470 145.570 328.490 ;
        RECT 172.060 328.470 175.220 328.610 ;
        RECT 138.800 327.910 141.960 328.240 ;
        RECT 137.830 327.180 140.780 327.510 ;
        RECT 137.830 327.170 138.180 327.180 ;
        RECT 137.830 327.140 138.220 327.170 ;
        RECT 141.640 327.140 141.960 327.910 ;
        RECT 172.060 327.430 172.380 328.470 ;
        RECT 144.250 327.160 144.580 327.200 ;
        RECT 144.240 327.140 144.590 327.160 ;
        RECT 137.830 326.850 147.900 327.140 ;
        RECT 172.060 327.110 175.220 327.430 ;
        RECT 172.680 327.100 172.990 327.110 ;
        RECT 173.780 327.100 174.090 327.110 ;
        RECT 174.880 327.100 175.190 327.110 ;
        RECT 41.170 215.460 43.620 218.980 ;
        RECT 41.350 215.340 43.430 215.460 ;
        RECT 49.850 161.840 51.930 326.520 ;
        RECT 137.830 326.310 138.180 326.850 ;
        RECT 141.640 326.510 141.960 326.850 ;
        RECT 144.250 326.830 144.580 326.850 ;
        RECT 137.830 326.180 138.210 326.310 ;
        RECT 137.830 326.140 138.580 326.180 ;
        RECT 141.640 326.170 144.050 326.510 ;
        RECT 139.380 326.140 139.690 326.160 ;
        RECT 137.830 325.840 140.780 326.140 ;
        RECT 139.380 325.830 139.690 325.840 ;
        RECT 140.470 325.810 140.780 325.840 ;
        RECT 141.640 325.930 144.090 326.170 ;
        RECT 141.640 325.910 144.050 325.930 ;
        RECT 138.830 325.460 139.140 325.470 ;
        RECT 141.640 325.460 141.960 325.910 ;
        RECT 143.080 325.840 143.740 325.910 ;
        RECT 143.110 325.830 143.710 325.840 ;
        RECT 138.810 325.130 141.960 325.460 ;
        RECT 138.810 325.120 141.870 325.130 ;
        RECT 147.600 324.770 147.890 326.850 ;
        RECT 175.840 326.760 176.190 328.690 ;
        RECT 173.250 326.750 176.190 326.760 ;
        RECT 173.240 326.440 176.190 326.750 ;
        RECT 176.510 326.760 176.860 328.690 ;
        RECT 177.480 328.470 180.640 328.690 ;
        RECT 180.320 328.240 180.640 328.470 ;
        RECT 181.870 328.500 185.030 328.690 ;
        RECT 181.870 328.240 182.190 328.500 ;
        RECT 185.650 328.240 186.000 328.690 ;
        RECT 186.320 328.240 186.670 328.690 ;
        RECT 187.290 328.500 190.450 328.690 ;
        RECT 190.130 328.240 190.450 328.500 ;
        RECT 192.810 328.240 193.160 328.690 ;
        RECT 193.780 328.480 196.940 328.690 ;
        RECT 217.820 328.670 218.380 328.690 ;
        RECT 196.620 328.240 196.940 328.480 ;
        RECT 180.200 327.780 217.280 328.240 ;
        RECT 180.270 327.680 180.790 327.780 ;
        RECT 180.320 327.430 180.640 327.680 ;
        RECT 177.480 327.110 180.640 327.430 ;
        RECT 181.870 327.460 182.190 327.780 ;
        RECT 181.870 327.330 185.030 327.460 ;
        RECT 185.650 327.330 186.000 327.780 ;
        RECT 186.320 327.330 186.670 327.780 ;
        RECT 190.130 327.460 190.450 327.780 ;
        RECT 187.290 327.330 190.450 327.460 ;
        RECT 192.810 327.330 193.160 327.780 ;
        RECT 196.620 327.440 196.940 327.780 ;
        RECT 216.630 327.720 217.190 327.780 ;
        RECT 193.780 327.330 196.940 327.440 ;
        RECT 181.640 327.260 216.190 327.330 ;
        RECT 177.510 327.100 177.820 327.110 ;
        RECT 178.610 327.100 178.920 327.110 ;
        RECT 179.710 327.100 180.020 327.110 ;
        RECT 181.630 326.870 216.190 327.260 ;
        RECT 176.510 326.750 179.450 326.760 ;
        RECT 176.510 326.440 179.460 326.750 ;
        RECT 173.240 326.430 175.960 326.440 ;
        RECT 176.740 326.430 179.460 326.440 ;
        RECT 173.240 326.420 173.550 326.430 ;
        RECT 174.330 326.420 174.640 326.430 ;
        RECT 178.060 326.420 178.370 326.430 ;
        RECT 179.150 326.420 179.460 326.430 ;
        RECT 181.630 326.740 182.280 326.870 ;
        RECT 185.650 326.790 186.000 326.870 ;
        RECT 183.060 326.780 186.000 326.790 ;
        RECT 181.630 326.350 182.230 326.740 ;
        RECT 183.050 326.470 186.000 326.780 ;
        RECT 186.320 326.790 186.670 326.870 ;
        RECT 186.320 326.780 189.260 326.790 ;
        RECT 186.320 326.470 189.270 326.780 ;
        RECT 183.050 326.460 185.770 326.470 ;
        RECT 186.550 326.460 189.270 326.470 ;
        RECT 183.050 326.450 183.360 326.460 ;
        RECT 184.140 326.450 184.450 326.460 ;
        RECT 187.870 326.450 188.180 326.460 ;
        RECT 188.960 326.450 189.270 326.460 ;
        RECT 190.090 326.410 190.690 326.840 ;
        RECT 192.810 326.770 193.160 326.870 ;
        RECT 215.500 326.850 216.060 326.870 ;
        RECT 192.810 326.760 195.750 326.770 ;
        RECT 192.810 326.450 195.760 326.760 ;
        RECT 193.040 326.440 195.760 326.450 ;
        RECT 194.360 326.430 194.670 326.440 ;
        RECT 195.450 326.430 195.760 326.440 ;
        RECT 190.080 326.390 190.690 326.410 ;
        RECT 196.580 326.390 197.180 326.820 ;
        RECT 214.570 326.390 215.130 326.400 ;
        RECT 181.630 326.020 182.240 326.350 ;
        RECT 190.080 325.930 215.220 326.390 ;
        RECT 190.080 325.880 190.610 325.930 ;
        RECT 190.080 325.830 190.600 325.880 ;
        RECT 164.020 324.770 164.340 324.790 ;
        RECT 220.020 324.770 221.180 324.800 ;
        RECT 102.100 324.610 102.560 324.620 ;
        RECT 102.100 324.170 127.970 324.610 ;
        RECT 102.100 324.150 102.560 324.170 ;
        RECT 125.730 323.470 127.000 324.170 ;
        RECT 147.410 323.650 221.180 324.770 ;
        RECT 164.020 323.630 164.340 323.650 ;
        RECT 175.390 323.570 177.310 323.650 ;
        RECT 185.200 323.540 187.130 323.650 ;
        RECT 220.020 323.620 221.180 323.650 ;
        RECT 125.730 323.450 135.700 323.470 ;
        RECT 54.100 323.090 135.700 323.450 ;
        RECT 54.100 321.370 127.960 323.090 ;
        RECT 135.320 322.240 135.700 323.090 ;
        RECT 363.620 322.960 365.020 348.920 ;
        RECT 369.920 324.880 371.320 352.540 ;
        RECT 369.910 324.370 371.320 324.880 ;
        RECT 368.800 324.200 371.320 324.370 ;
        RECT 369.910 323.950 371.320 324.200 ;
        RECT 363.490 322.880 365.020 322.960 ;
        RECT 136.620 322.240 136.990 322.250 ;
        RECT 135.320 321.860 138.040 322.240 ;
        RECT 362.980 321.870 365.020 322.880 ;
        RECT 136.620 321.840 136.990 321.860 ;
        RECT 223.860 321.470 224.060 321.480 ;
        RECT 227.580 321.470 227.900 321.520 ;
        RECT 49.430 158.170 52.140 161.840 ;
        RECT 49.850 157.450 51.930 158.170 ;
        RECT 54.100 133.220 56.180 321.370 ;
        RECT 223.860 321.320 227.900 321.470 ;
        RECT 126.940 320.320 127.440 320.430 ;
        RECT 195.910 320.350 196.300 320.360 ;
        RECT 195.900 320.320 196.300 320.350 ;
        RECT 126.940 320.040 196.300 320.320 ;
        RECT 126.940 319.960 127.440 320.040 ;
        RECT 195.900 320.020 196.300 320.040 ;
        RECT 195.910 320.010 196.300 320.020 ;
        RECT 223.180 319.230 223.610 319.250 ;
        RECT 204.680 319.200 206.640 319.230 ;
        RECT 223.160 319.200 223.620 319.230 ;
        RECT 204.680 318.850 223.620 319.200 ;
        RECT 204.680 312.750 206.640 318.850 ;
        RECT 223.160 318.830 223.620 318.850 ;
        RECT 223.180 318.820 223.610 318.830 ;
        RECT 223.860 318.410 224.060 321.320 ;
        RECT 227.580 321.200 227.900 321.320 ;
        RECT 362.980 321.230 368.030 321.870 ;
        RECT 362.980 320.950 365.020 321.230 ;
        RECT 362.910 320.330 365.020 320.950 ;
        RECT 224.830 319.910 227.600 319.920 ;
        RECT 224.830 319.720 227.900 319.910 ;
        RECT 224.080 318.420 224.510 318.440 ;
        RECT 224.070 318.410 224.520 318.420 ;
        RECT 208.610 318.030 224.520 318.410 ;
        RECT 204.650 312.100 206.680 312.750 ;
        RECT 208.610 312.730 210.570 318.030 ;
        RECT 222.710 317.870 222.970 318.030 ;
        RECT 222.740 317.590 222.940 317.870 ;
        RECT 223.860 317.590 224.060 318.030 ;
        RECT 224.080 318.010 224.510 318.030 ;
        RECT 224.830 317.600 225.040 319.720 ;
        RECT 227.580 319.590 227.900 319.720 ;
        RECT 226.610 318.260 226.920 318.290 ;
        RECT 227.570 318.260 227.890 318.300 ;
        RECT 226.610 318.010 227.890 318.260 ;
        RECT 224.830 317.590 225.450 317.600 ;
        RECT 212.760 317.210 225.450 317.590 ;
        RECT 212.760 312.750 214.740 317.210 ;
        RECT 222.740 316.800 222.940 317.210 ;
        RECT 223.860 316.800 224.060 317.210 ;
        RECT 224.830 316.800 225.040 317.210 ;
        RECT 225.840 316.800 226.260 316.830 ;
        RECT 216.870 316.420 226.260 316.800 ;
        RECT 208.600 312.080 210.630 312.730 ;
        RECT 212.720 312.100 214.750 312.750 ;
        RECT 216.870 312.720 218.850 316.420 ;
        RECT 222.740 313.630 222.940 316.420 ;
        RECT 223.860 313.630 224.060 316.420 ;
        RECT 224.830 313.630 225.040 316.420 ;
        RECT 225.840 316.390 226.260 316.420 ;
        RECT 226.610 313.630 226.910 318.010 ;
        RECT 227.570 317.980 227.890 318.010 ;
        RECT 227.570 316.660 227.890 316.680 ;
        RECT 227.570 316.360 227.920 316.660 ;
        RECT 227.730 315.070 227.920 316.360 ;
        RECT 227.570 314.750 227.920 315.070 ;
        RECT 227.730 313.630 227.920 314.750 ;
        RECT 221.940 313.430 228.180 313.630 ;
        RECT 221.940 312.750 222.140 313.430 ;
        RECT 222.740 312.750 222.940 313.430 ;
        RECT 216.860 312.070 218.890 312.720 ;
        RECT 220.850 312.100 222.940 312.750 ;
        RECT 222.740 309.610 222.940 312.100 ;
        RECT 223.860 309.750 224.060 313.430 ;
        RECT 223.850 309.610 224.060 309.750 ;
        RECT 224.830 312.750 225.040 313.430 ;
        RECT 226.610 313.310 226.910 313.430 ;
        RECT 227.200 313.310 227.520 313.430 ;
        RECT 226.610 313.220 227.520 313.310 ;
        RECT 227.730 313.220 227.920 313.430 ;
        RECT 229.100 313.220 229.300 313.630 ;
        RECT 226.610 313.020 229.300 313.220 ;
        RECT 226.610 312.750 227.070 313.020 ;
        RECT 224.830 312.450 227.070 312.750 ;
        RECT 224.830 312.100 226.910 312.450 ;
        RECT 224.830 309.610 225.040 312.100 ;
        RECT 226.610 311.670 226.910 312.100 ;
        RECT 227.730 311.870 227.920 313.020 ;
        RECT 226.610 311.510 226.970 311.670 ;
        RECT 227.580 311.550 227.920 311.870 ;
        RECT 226.260 310.070 226.580 310.140 ;
        RECT 226.760 310.070 226.970 311.510 ;
        RECT 227.730 310.280 227.920 311.550 ;
        RECT 226.260 309.870 226.970 310.070 ;
        RECT 227.570 309.960 227.920 310.280 ;
        RECT 226.260 309.820 226.580 309.870 ;
        RECT 226.760 309.610 226.970 309.870 ;
        RECT 227.730 309.760 227.920 309.960 ;
        RECT 227.710 309.610 227.920 309.760 ;
        RECT 363.620 294.370 365.020 320.330 ;
        RECT 369.920 296.290 371.320 323.950 ;
        RECT 369.910 295.780 371.320 296.290 ;
        RECT 368.800 295.610 371.320 295.780 ;
        RECT 369.910 295.360 371.320 295.610 ;
        RECT 363.490 294.290 365.020 294.370 ;
        RECT 362.980 293.280 365.020 294.290 ;
        RECT 362.980 292.640 368.030 293.280 ;
        RECT 362.980 292.360 365.020 292.640 ;
        RECT 362.910 291.740 365.020 292.360 ;
        RECT 363.620 265.780 365.020 291.740 ;
        RECT 369.920 267.700 371.320 295.360 ;
        RECT 369.910 267.190 371.320 267.700 ;
        RECT 368.800 267.020 371.320 267.190 ;
        RECT 369.910 266.770 371.320 267.020 ;
        RECT 363.490 265.700 365.020 265.780 ;
        RECT 362.980 264.690 365.020 265.700 ;
        RECT 362.980 264.050 368.030 264.690 ;
        RECT 362.980 263.770 365.020 264.050 ;
        RECT 362.910 263.150 365.020 263.770 ;
        RECT 363.620 237.190 365.020 263.150 ;
        RECT 369.920 239.110 371.320 266.770 ;
        RECT 369.910 238.600 371.320 239.110 ;
        RECT 368.800 238.430 371.320 238.600 ;
        RECT 369.910 238.180 371.320 238.430 ;
        RECT 363.490 237.110 365.020 237.190 ;
        RECT 362.980 236.100 365.020 237.110 ;
        RECT 362.980 235.460 368.030 236.100 ;
        RECT 362.980 235.180 365.020 235.460 ;
        RECT 362.910 234.560 365.020 235.180 ;
        RECT 363.620 208.600 365.020 234.560 ;
        RECT 369.920 210.520 371.320 238.180 ;
        RECT 369.910 210.010 371.320 210.520 ;
        RECT 368.800 209.840 371.320 210.010 ;
        RECT 369.910 209.590 371.320 209.840 ;
        RECT 363.490 208.520 365.020 208.600 ;
        RECT 362.980 207.510 365.020 208.520 ;
        RECT 362.980 206.870 368.030 207.510 ;
        RECT 362.980 206.590 365.020 206.870 ;
        RECT 362.910 205.970 365.020 206.590 ;
        RECT 363.620 180.530 365.020 205.970 ;
        RECT 369.920 181.930 371.320 209.590 ;
        RECT 369.910 181.420 371.320 181.930 ;
        RECT 368.800 181.250 371.320 181.420 ;
        RECT 369.910 181.000 371.320 181.250 ;
        RECT 369.920 180.530 371.320 181.000 ;
        RECT 53.770 129.740 56.510 133.220 ;
        RECT 54.100 128.930 56.180 129.740 ;
      LAYER via2 ;
        RECT 202.310 367.230 202.630 367.550 ;
        RECT 203.340 367.220 203.660 367.540 ;
    END
  END IO08
  PIN IO09
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 369.830 265.620 370.820 265.630 ;
        RECT 369.830 265.100 371.220 265.620 ;
        RECT 370.730 261.490 371.220 265.100 ;
        RECT 371.100 240.520 373.060 241.870 ;
        RECT 370.670 240.460 373.060 240.520 ;
        RECT 370.650 239.880 373.060 240.460 ;
        RECT 370.670 239.130 373.060 239.880 ;
        RECT 363.040 238.410 373.060 239.130 ;
        RECT 368.710 238.180 373.060 238.410 ;
        RECT 370.670 238.150 373.060 238.180 ;
        RECT 371.100 237.980 373.060 238.150 ;
      LAYER via ;
        RECT 370.020 265.190 370.780 265.540 ;
        RECT 370.820 261.760 371.170 264.750 ;
        RECT 369.960 238.310 370.580 239.010 ;
        RECT 370.820 238.370 371.150 240.400 ;
    END
  END IO09
  PIN IO10
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 369.830 294.210 370.820 294.220 ;
        RECT 369.830 293.690 371.220 294.210 ;
        RECT 370.730 290.080 371.220 293.690 ;
        RECT 371.830 270.470 373.080 270.480 ;
        RECT 371.110 269.110 373.080 270.470 ;
        RECT 370.670 269.050 373.080 269.110 ;
        RECT 370.650 268.470 373.080 269.050 ;
        RECT 370.670 267.720 373.080 268.470 ;
        RECT 363.040 267.000 373.080 267.720 ;
        RECT 368.710 266.770 373.080 267.000 ;
        RECT 370.670 266.740 373.080 266.770 ;
        RECT 371.110 266.590 373.080 266.740 ;
        RECT 371.110 266.580 371.830 266.590 ;
      LAYER via ;
        RECT 370.020 293.780 370.780 294.130 ;
        RECT 370.820 290.350 371.170 293.340 ;
        RECT 369.960 266.900 370.580 267.600 ;
        RECT 370.820 266.960 371.150 268.990 ;
    END
  END IO10
  PIN IO11
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 369.830 322.800 370.820 322.810 ;
        RECT 369.830 322.280 371.220 322.800 ;
        RECT 370.730 318.670 371.220 322.280 ;
        RECT 371.110 297.700 373.070 299.040 ;
        RECT 370.670 297.640 373.070 297.700 ;
        RECT 370.650 297.060 373.070 297.640 ;
        RECT 370.670 296.310 373.070 297.060 ;
        RECT 363.040 295.590 373.070 296.310 ;
        RECT 368.710 295.360 373.070 295.590 ;
        RECT 370.670 295.330 373.070 295.360 ;
        RECT 371.110 295.150 373.070 295.330 ;
      LAYER via ;
        RECT 370.020 322.370 370.780 322.720 ;
        RECT 370.820 318.940 371.170 321.930 ;
        RECT 369.960 295.490 370.580 296.190 ;
        RECT 370.820 295.550 371.150 297.580 ;
    END
  END IO11
  PIN IO12
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 369.830 351.390 370.820 351.400 ;
        RECT 369.830 350.870 371.220 351.390 ;
        RECT 370.730 347.260 371.220 350.870 ;
        RECT 371.110 326.290 373.070 327.640 ;
        RECT 370.670 326.230 373.070 326.290 ;
        RECT 370.650 325.650 373.070 326.230 ;
        RECT 370.670 324.900 373.070 325.650 ;
        RECT 363.040 324.180 373.070 324.900 ;
        RECT 368.710 323.950 373.070 324.180 ;
        RECT 370.670 323.920 373.070 323.950 ;
        RECT 371.110 323.750 373.070 323.920 ;
      LAYER via ;
        RECT 370.020 350.960 370.780 351.310 ;
        RECT 370.820 347.530 371.170 350.520 ;
        RECT 369.960 324.080 370.580 324.780 ;
        RECT 370.820 324.140 371.150 326.170 ;
    END
  END IO12
  PIN IO13
    ANTENNADIFFAREA 97.647797 ;
    PORT
      LAYER met1 ;
        RECT 336.600 387.110 340.490 389.070 ;
        RECT 336.770 386.660 339.140 387.110 ;
        RECT 360.110 386.810 364.240 387.210 ;
        RECT 360.110 386.720 364.250 386.810 ;
        RECT 336.800 384.700 337.750 386.660 ;
        RECT 338.500 386.640 339.080 386.660 ;
        RECT 363.720 385.820 364.250 386.720 ;
        RECT 337.030 379.030 337.750 384.700 ;
        RECT 369.830 379.980 370.820 379.990 ;
        RECT 369.830 379.460 371.220 379.980 ;
        RECT 370.730 375.850 371.220 379.460 ;
        RECT 371.830 356.230 373.080 356.240 ;
        RECT 371.110 354.880 373.080 356.230 ;
        RECT 370.670 354.820 373.080 354.880 ;
        RECT 370.650 354.240 373.080 354.820 ;
        RECT 370.670 353.490 373.080 354.240 ;
        RECT 363.040 352.770 373.080 353.490 ;
        RECT 368.710 352.540 373.080 352.770 ;
        RECT 370.670 352.510 373.080 352.540 ;
        RECT 371.110 352.350 373.080 352.510 ;
        RECT 371.110 352.340 371.830 352.350 ;
      LAYER via ;
        RECT 336.990 386.810 339.020 387.140 ;
        RECT 360.380 386.810 363.370 387.160 ;
        RECT 336.930 385.950 337.630 386.570 ;
        RECT 363.810 386.010 364.160 386.770 ;
        RECT 370.020 379.550 370.780 379.900 ;
        RECT 370.820 376.120 371.170 379.110 ;
        RECT 369.960 352.670 370.580 353.370 ;
        RECT 370.820 352.730 371.150 354.760 ;
    END
  END IO13
  PIN IO25
    ANTENNADIFFAREA 636.910278 ;
    PORT
      LAYER met2 ;
        RECT 2.090 354.190 3.490 381.380 ;
        RECT 2.090 353.680 3.500 354.190 ;
        RECT 2.090 353.510 4.610 353.680 ;
        RECT 2.090 353.260 3.500 353.510 ;
        RECT 2.090 325.600 3.490 353.260 ;
        RECT 2.090 325.090 3.500 325.600 ;
        RECT 2.090 324.920 4.610 325.090 ;
        RECT 2.090 324.670 3.500 324.920 ;
        RECT 2.090 297.010 3.490 324.670 ;
        RECT 2.090 296.500 3.500 297.010 ;
        RECT 2.090 296.330 4.610 296.500 ;
        RECT 2.090 296.080 3.500 296.330 ;
        RECT 2.090 268.420 3.490 296.080 ;
        RECT 2.090 267.910 3.500 268.420 ;
        RECT 2.090 267.740 4.610 267.910 ;
        RECT 2.090 267.490 3.500 267.740 ;
        RECT 2.090 239.830 3.490 267.490 ;
        RECT 2.090 239.320 3.500 239.830 ;
        RECT 2.090 239.150 4.610 239.320 ;
        RECT 2.090 238.900 3.500 239.150 ;
        RECT 2.090 211.240 3.490 238.900 ;
        RECT 2.090 210.730 3.500 211.240 ;
        RECT 2.090 210.560 4.610 210.730 ;
        RECT 2.090 210.310 3.500 210.560 ;
        RECT 2.090 182.650 3.490 210.310 ;
        RECT 2.090 182.140 3.500 182.650 ;
        RECT 2.090 181.970 4.610 182.140 ;
        RECT 2.090 181.720 3.500 181.970 ;
        RECT 2.090 154.060 3.490 181.720 ;
        RECT 2.090 153.550 3.500 154.060 ;
        RECT 2.090 153.380 4.610 153.550 ;
        RECT 2.090 153.130 3.500 153.380 ;
        RECT 2.090 125.470 3.490 153.130 ;
        RECT 2.090 124.960 3.500 125.470 ;
        RECT 2.090 124.790 4.610 124.960 ;
        RECT 2.090 124.540 3.500 124.790 ;
        RECT 2.090 96.880 3.490 124.540 ;
        RECT 2.090 96.370 3.500 96.880 ;
        RECT 2.090 96.200 4.610 96.370 ;
        RECT 2.090 95.950 3.500 96.200 ;
        RECT 2.090 68.290 3.490 95.950 ;
        RECT 2.090 67.780 3.500 68.290 ;
        RECT 2.090 67.610 4.610 67.780 ;
        RECT 2.090 67.360 3.500 67.610 ;
        RECT 2.090 39.700 3.490 67.360 ;
        RECT 2.090 39.190 3.500 39.700 ;
        RECT 2.090 39.020 4.610 39.190 ;
        RECT 2.090 38.770 3.500 39.020 ;
        RECT 2.090 11.110 3.490 38.770 ;
        RECT 2.090 10.600 3.500 11.110 ;
        RECT 2.090 10.430 4.610 10.600 ;
        RECT 2.090 10.180 3.500 10.430 ;
        RECT 2.090 9.710 3.490 10.180 ;
    END
  END IO25
  PIN IO26
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 2.590 352.110 3.580 352.120 ;
        RECT 2.190 351.590 3.580 352.110 ;
        RECT 2.190 347.980 2.680 351.590 ;
        RECT 0.240 327.010 2.290 328.360 ;
        RECT 0.240 326.950 2.740 327.010 ;
        RECT 0.240 326.370 2.760 326.950 ;
        RECT 0.240 325.620 2.740 326.370 ;
        RECT 0.240 324.900 10.370 325.620 ;
        RECT 0.240 324.670 4.700 324.900 ;
        RECT 0.240 324.640 2.740 324.670 ;
        RECT 0.240 324.470 2.290 324.640 ;
        RECT 1.480 324.460 2.290 324.470 ;
      LAYER via ;
        RECT 2.630 351.680 3.390 352.030 ;
        RECT 2.240 348.250 2.590 351.240 ;
        RECT 2.260 324.860 2.590 326.890 ;
        RECT 2.830 324.800 3.450 325.500 ;
    END
  END IO26
  PIN IO27
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 2.590 323.520 3.580 323.530 ;
        RECT 2.190 323.000 3.580 323.520 ;
        RECT 2.190 319.390 2.680 323.000 ;
        RECT 1.480 299.760 2.290 299.770 ;
        RECT 0.230 298.420 2.290 299.760 ;
        RECT 0.230 298.360 2.740 298.420 ;
        RECT 0.230 297.780 2.760 298.360 ;
        RECT 0.230 297.030 2.740 297.780 ;
        RECT 0.230 296.310 10.370 297.030 ;
        RECT 0.230 296.080 4.700 296.310 ;
        RECT 0.230 296.050 2.740 296.080 ;
        RECT 0.230 295.870 2.290 296.050 ;
      LAYER via ;
        RECT 2.630 323.090 3.390 323.440 ;
        RECT 2.240 319.660 2.590 322.650 ;
        RECT 2.260 296.270 2.590 298.300 ;
        RECT 2.830 296.210 3.450 296.910 ;
    END
  END IO27
  PIN IO28
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 2.590 294.930 3.580 294.940 ;
        RECT 2.190 294.410 3.580 294.930 ;
        RECT 2.190 290.800 2.680 294.410 ;
        RECT 1.490 271.170 2.300 271.180 ;
        RECT 0.250 269.830 2.300 271.170 ;
        RECT 0.250 269.770 2.740 269.830 ;
        RECT 0.250 269.190 2.760 269.770 ;
        RECT 0.250 268.440 2.740 269.190 ;
        RECT 0.250 267.720 10.370 268.440 ;
        RECT 0.250 267.490 4.700 267.720 ;
        RECT 0.250 267.460 2.740 267.490 ;
        RECT 0.250 267.280 2.300 267.460 ;
      LAYER via ;
        RECT 2.630 294.500 3.390 294.850 ;
        RECT 2.240 291.070 2.590 294.060 ;
        RECT 2.260 267.680 2.590 269.710 ;
        RECT 2.830 267.620 3.450 268.320 ;
    END
  END IO28
  PIN IO29
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 2.590 266.340 3.580 266.350 ;
        RECT 2.190 265.820 3.580 266.340 ;
        RECT 2.190 262.210 2.680 265.820 ;
        RECT 0.240 241.240 2.290 242.590 ;
        RECT 0.240 241.180 2.740 241.240 ;
        RECT 0.240 240.600 2.760 241.180 ;
        RECT 0.240 239.850 2.740 240.600 ;
        RECT 0.240 239.130 10.370 239.850 ;
        RECT 0.240 238.900 4.700 239.130 ;
        RECT 0.240 238.870 2.740 238.900 ;
        RECT 0.240 238.700 2.290 238.870 ;
        RECT 1.480 238.690 2.290 238.700 ;
      LAYER via ;
        RECT 2.630 265.910 3.390 266.260 ;
        RECT 2.240 262.480 2.590 265.470 ;
        RECT 2.260 239.090 2.590 241.120 ;
        RECT 2.830 239.030 3.450 239.730 ;
    END
  END IO29
  PIN IO30
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 2.590 237.750 3.580 237.760 ;
        RECT 2.190 237.230 3.580 237.750 ;
        RECT 2.190 233.620 2.680 237.230 ;
        RECT 1.480 213.990 2.290 214.000 ;
        RECT 0.230 212.650 2.290 213.990 ;
        RECT 0.230 212.590 2.740 212.650 ;
        RECT 0.230 212.010 2.760 212.590 ;
        RECT 0.230 211.260 2.740 212.010 ;
        RECT 0.230 210.540 10.370 211.260 ;
        RECT 0.230 210.310 4.700 210.540 ;
        RECT 0.230 210.280 2.740 210.310 ;
        RECT 0.230 210.100 2.290 210.280 ;
      LAYER via ;
        RECT 2.630 237.320 3.390 237.670 ;
        RECT 2.240 233.890 2.590 236.880 ;
        RECT 2.260 210.500 2.590 212.530 ;
        RECT 2.830 210.440 3.450 211.140 ;
    END
  END IO30
  PIN IO31
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 2.590 209.160 3.580 209.170 ;
        RECT 2.190 208.640 3.580 209.160 ;
        RECT 2.190 205.030 2.680 208.640 ;
        RECT 1.480 185.410 2.290 185.420 ;
        RECT 0.240 184.060 2.290 185.410 ;
        RECT 0.240 184.000 2.740 184.060 ;
        RECT 0.240 183.420 2.760 184.000 ;
        RECT 0.240 182.670 2.740 183.420 ;
        RECT 0.240 181.950 10.370 182.670 ;
        RECT 0.240 181.720 4.700 181.950 ;
        RECT 0.240 181.690 2.740 181.720 ;
        RECT 0.240 181.520 2.290 181.690 ;
      LAYER via ;
        RECT 2.630 208.730 3.390 209.080 ;
        RECT 2.240 205.300 2.590 208.290 ;
        RECT 2.260 181.910 2.590 183.940 ;
        RECT 2.830 181.850 3.450 182.550 ;
    END
  END IO31
  PIN IO32
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 2.590 180.570 3.580 180.580 ;
        RECT 2.190 180.050 3.580 180.570 ;
        RECT 2.190 176.440 2.680 180.050 ;
        RECT 0.270 155.470 2.310 156.830 ;
        RECT 0.270 155.410 2.740 155.470 ;
        RECT 0.270 154.830 2.760 155.410 ;
        RECT 0.270 154.080 2.740 154.830 ;
        RECT 0.270 153.360 10.370 154.080 ;
        RECT 0.270 153.130 4.700 153.360 ;
        RECT 0.270 153.100 2.740 153.130 ;
        RECT 0.270 152.940 2.310 153.100 ;
        RECT 1.500 152.930 2.310 152.940 ;
      LAYER via ;
        RECT 2.630 180.140 3.390 180.490 ;
        RECT 2.240 176.710 2.590 179.700 ;
        RECT 2.260 153.320 2.590 155.350 ;
        RECT 2.830 153.260 3.450 153.960 ;
    END
  END IO32
  PIN IO33
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 2.590 151.980 3.580 151.990 ;
        RECT 2.190 151.460 3.580 151.980 ;
        RECT 2.190 147.850 2.680 151.460 ;
        RECT 1.490 128.220 2.300 128.230 ;
        RECT 0.250 126.880 2.300 128.220 ;
        RECT 0.250 126.820 2.740 126.880 ;
        RECT 0.250 126.240 2.760 126.820 ;
        RECT 0.250 125.490 2.740 126.240 ;
        RECT 0.250 124.770 10.370 125.490 ;
        RECT 0.250 124.540 4.700 124.770 ;
        RECT 0.250 124.510 2.740 124.540 ;
        RECT 0.250 124.330 2.300 124.510 ;
      LAYER via ;
        RECT 2.630 151.550 3.390 151.900 ;
        RECT 2.240 148.120 2.590 151.110 ;
        RECT 2.260 124.730 2.590 126.760 ;
        RECT 2.830 124.670 3.450 125.370 ;
    END
  END IO33
  PIN IO34
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 2.590 123.390 3.580 123.400 ;
        RECT 2.190 122.870 3.580 123.390 ;
        RECT 2.190 119.260 2.680 122.870 ;
        RECT 1.490 99.630 2.300 99.640 ;
        RECT 0.240 98.290 2.300 99.630 ;
        RECT 0.240 98.230 2.740 98.290 ;
        RECT 0.240 97.650 2.760 98.230 ;
        RECT 0.240 96.900 2.740 97.650 ;
        RECT 0.240 96.180 10.370 96.900 ;
        RECT 0.240 95.950 4.700 96.180 ;
        RECT 0.240 95.920 2.740 95.950 ;
        RECT 0.240 95.740 2.300 95.920 ;
      LAYER via ;
        RECT 2.630 122.960 3.390 123.310 ;
        RECT 2.240 119.530 2.590 122.520 ;
        RECT 2.260 96.140 2.590 98.170 ;
        RECT 2.830 96.080 3.450 96.780 ;
    END
  END IO34
  PIN IO35
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 2.590 94.800 3.580 94.810 ;
        RECT 2.190 94.280 3.580 94.800 ;
        RECT 2.190 90.670 2.680 94.280 ;
        RECT 1.490 71.040 2.300 71.050 ;
        RECT 0.240 69.700 2.300 71.040 ;
        RECT 0.240 69.640 2.740 69.700 ;
        RECT 0.240 69.060 2.760 69.640 ;
        RECT 0.240 68.310 2.740 69.060 ;
        RECT 0.240 67.590 10.370 68.310 ;
        RECT 0.240 67.360 4.700 67.590 ;
        RECT 0.240 67.330 2.740 67.360 ;
        RECT 0.240 67.150 2.300 67.330 ;
      LAYER via ;
        RECT 2.630 94.370 3.390 94.720 ;
        RECT 2.240 90.940 2.590 93.930 ;
        RECT 2.260 67.550 2.590 69.580 ;
        RECT 2.830 67.490 3.450 68.190 ;
    END
  END IO35
  PIN IO36
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 2.590 66.210 3.580 66.220 ;
        RECT 2.190 65.690 3.580 66.210 ;
        RECT 2.190 62.080 2.680 65.690 ;
        RECT 1.500 42.450 2.310 42.460 ;
        RECT 0.250 41.110 2.310 42.450 ;
        RECT 0.250 41.050 2.740 41.110 ;
        RECT 0.250 40.470 2.760 41.050 ;
        RECT 0.250 39.720 2.740 40.470 ;
        RECT 0.250 39.000 10.370 39.720 ;
        RECT 0.250 38.770 4.700 39.000 ;
        RECT 0.250 38.740 2.740 38.770 ;
        RECT 0.250 38.560 2.310 38.740 ;
      LAYER via ;
        RECT 2.630 65.780 3.390 66.130 ;
        RECT 2.240 62.350 2.590 65.340 ;
        RECT 2.260 38.960 2.590 40.990 ;
        RECT 2.830 38.900 3.450 39.600 ;
    END
  END IO36
  PIN IO37
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 2.590 37.620 3.580 37.630 ;
        RECT 2.190 37.100 3.580 37.620 ;
        RECT 2.190 33.490 2.680 37.100 ;
        RECT 0.250 12.520 2.290 13.870 ;
        RECT 0.250 12.460 2.740 12.520 ;
        RECT 0.250 11.880 2.760 12.460 ;
        RECT 0.250 11.130 2.740 11.880 ;
        RECT 0.250 10.410 10.370 11.130 ;
        RECT 0.250 10.180 4.700 10.410 ;
        RECT 0.250 10.150 2.740 10.180 ;
        RECT 0.250 9.980 2.290 10.150 ;
        RECT 1.480 9.970 2.290 9.980 ;
      LAYER via ;
        RECT 2.630 37.190 3.390 37.540 ;
        RECT 2.240 33.760 2.590 36.750 ;
        RECT 2.260 10.370 2.590 12.400 ;
        RECT 2.830 10.310 3.450 11.010 ;
    END
  END IO37
  PIN VSSA1
    ANTENNADIFFAREA 118.154396 ;
    PORT
      LAYER nwell ;
        RECT 3.020 367.660 8.960 379.710 ;
        RECT 3.020 339.070 8.960 351.120 ;
        RECT 3.020 310.480 8.960 322.530 ;
        RECT 3.020 281.890 8.960 293.940 ;
        RECT 3.020 253.300 8.960 265.350 ;
        RECT 3.020 224.710 8.960 236.760 ;
        RECT 3.020 196.120 8.960 208.170 ;
        RECT 3.020 167.530 8.960 179.580 ;
        RECT 3.020 138.940 8.960 150.990 ;
        RECT 3.020 110.350 8.960 122.400 ;
        RECT 3.020 81.760 8.960 93.810 ;
        RECT 3.020 53.170 8.960 65.220 ;
        RECT 3.020 24.580 8.960 36.630 ;
      LAYER met2 ;
        RECT 3.650 385.010 16.580 385.020 ;
        RECT 3.520 383.620 16.580 385.010 ;
        RECT 3.520 382.100 5.810 383.620 ;
        RECT 3.970 382.060 5.810 382.100 ;
        RECT 4.410 379.770 5.810 382.060 ;
        RECT 8.390 380.860 9.790 381.380 ;
        RECT 8.390 380.780 9.920 380.860 ;
        RECT 8.390 379.770 10.430 380.780 ;
        RECT 4.410 379.130 10.430 379.770 ;
        RECT 4.410 373.540 5.810 379.130 ;
        RECT 8.390 378.850 10.430 379.130 ;
        RECT 8.390 378.230 10.500 378.850 ;
        RECT 8.390 352.270 9.790 378.230 ;
        RECT 8.390 352.190 9.920 352.270 ;
        RECT 8.390 351.180 10.430 352.190 ;
        RECT 5.380 350.540 10.430 351.180 ;
        RECT 8.390 350.260 10.430 350.540 ;
        RECT 8.390 349.640 10.500 350.260 ;
        RECT 8.390 323.680 9.790 349.640 ;
        RECT 8.390 323.600 9.920 323.680 ;
        RECT 8.390 322.590 10.430 323.600 ;
        RECT 5.380 321.950 10.430 322.590 ;
        RECT 8.390 321.670 10.430 321.950 ;
        RECT 8.390 321.050 10.500 321.670 ;
        RECT 8.390 295.090 9.790 321.050 ;
        RECT 8.390 295.010 9.920 295.090 ;
        RECT 8.390 294.000 10.430 295.010 ;
        RECT 5.380 293.360 10.430 294.000 ;
        RECT 8.390 293.080 10.430 293.360 ;
        RECT 8.390 292.460 10.500 293.080 ;
        RECT 8.390 266.500 9.790 292.460 ;
        RECT 8.390 266.420 9.920 266.500 ;
        RECT 8.390 265.410 10.430 266.420 ;
        RECT 5.380 264.770 10.430 265.410 ;
        RECT 8.390 264.490 10.430 264.770 ;
        RECT 8.390 263.870 10.500 264.490 ;
        RECT 8.390 237.910 9.790 263.870 ;
        RECT 8.390 237.830 9.920 237.910 ;
        RECT 8.390 236.820 10.430 237.830 ;
        RECT 5.380 236.180 10.430 236.820 ;
        RECT 8.390 235.900 10.430 236.180 ;
        RECT 8.390 235.280 10.500 235.900 ;
        RECT 8.390 209.320 9.790 235.280 ;
        RECT 8.390 209.240 9.920 209.320 ;
        RECT 8.390 208.230 10.430 209.240 ;
        RECT 5.380 207.590 10.430 208.230 ;
        RECT 8.390 207.310 10.430 207.590 ;
        RECT 8.390 206.690 10.500 207.310 ;
        RECT 8.390 180.730 9.790 206.690 ;
        RECT 8.390 180.650 9.920 180.730 ;
        RECT 8.390 179.640 10.430 180.650 ;
        RECT 5.380 179.000 10.430 179.640 ;
        RECT 8.390 178.720 10.430 179.000 ;
        RECT 8.390 178.100 10.500 178.720 ;
        RECT 8.390 152.140 9.790 178.100 ;
        RECT 8.390 152.060 9.920 152.140 ;
        RECT 8.390 151.050 10.430 152.060 ;
        RECT 5.380 150.410 10.430 151.050 ;
        RECT 8.390 150.130 10.430 150.410 ;
        RECT 8.390 149.510 10.500 150.130 ;
        RECT 8.390 123.550 9.790 149.510 ;
        RECT 8.390 123.470 9.920 123.550 ;
        RECT 8.390 122.460 10.430 123.470 ;
        RECT 5.380 121.820 10.430 122.460 ;
        RECT 8.390 121.540 10.430 121.820 ;
        RECT 8.390 120.920 10.500 121.540 ;
        RECT 8.390 94.960 9.790 120.920 ;
        RECT 8.390 94.880 9.920 94.960 ;
        RECT 8.390 93.870 10.430 94.880 ;
        RECT 5.380 93.230 10.430 93.870 ;
        RECT 8.390 92.950 10.430 93.230 ;
        RECT 8.390 92.330 10.500 92.950 ;
        RECT 8.390 66.370 9.790 92.330 ;
        RECT 8.390 66.290 9.920 66.370 ;
        RECT 8.390 65.280 10.430 66.290 ;
        RECT 5.380 64.640 10.430 65.280 ;
        RECT 8.390 64.360 10.430 64.640 ;
        RECT 8.390 63.740 10.500 64.360 ;
        RECT 8.390 37.780 9.790 63.740 ;
        RECT 8.390 37.700 9.920 37.780 ;
        RECT 8.390 36.690 10.430 37.700 ;
        RECT 5.380 36.050 10.430 36.690 ;
        RECT 8.390 35.770 10.430 36.050 ;
        RECT 8.390 35.150 10.500 35.770 ;
        RECT 8.390 9.710 9.790 35.150 ;
    END
  END VSSA1
  PIN ANALOG10
    ANTENNADIFFAREA 146.979294 ;
    PORT
      LAYER met2 ;
        RECT 23.590 385.910 109.360 387.310 ;
        RECT 24.060 385.900 24.990 385.910 ;
        RECT 52.650 385.900 53.580 385.910 ;
        RECT 81.240 385.900 82.170 385.910 ;
        RECT 24.310 384.790 24.480 385.900 ;
        RECT 52.900 384.790 53.070 385.900 ;
        RECT 81.490 384.790 81.660 385.900 ;
    END
  END ANALOG10
  PIN ANALOG09
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 52.440 387.110 56.330 389.070 ;
        RECT 52.620 386.660 54.990 387.110 ;
        RECT 75.960 386.810 80.090 387.210 ;
        RECT 75.960 386.720 80.100 386.810 ;
        RECT 52.650 384.700 53.600 386.660 ;
        RECT 54.350 386.640 54.930 386.660 ;
        RECT 79.570 385.820 80.100 386.720 ;
        RECT 52.880 379.030 53.600 384.700 ;
      LAYER via ;
        RECT 52.840 386.810 54.870 387.140 ;
        RECT 76.230 386.810 79.220 387.160 ;
        RECT 52.780 385.950 53.480 386.570 ;
        RECT 79.660 386.010 80.010 386.770 ;
    END
  END ANALOG09
  PIN ANALOG08
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 81.030 387.110 84.920 389.070 ;
        RECT 81.210 386.660 83.580 387.110 ;
        RECT 104.550 386.810 108.680 387.210 ;
        RECT 104.550 386.720 108.690 386.810 ;
        RECT 81.240 384.700 82.190 386.660 ;
        RECT 82.940 386.640 83.520 386.660 ;
        RECT 108.160 385.820 108.690 386.720 ;
        RECT 81.470 379.030 82.190 384.700 ;
      LAYER via ;
        RECT 81.430 386.810 83.460 387.140 ;
        RECT 104.820 386.810 107.810 387.160 ;
        RECT 81.370 385.950 82.070 386.570 ;
        RECT 108.250 386.010 108.600 386.770 ;
    END
  END ANALOG08
  PIN ANALOG07
    PORT
      LAYER met1 ;
        RECT 122.930 387.130 126.820 389.100 ;
    END
  END ANALOG07
  PIN ANALOG06
    ANTENNAGATEAREA 12.719800 ;
    ANTENNADIFFAREA 129.537796 ;
    PORT
      LAYER met1 ;
        RECT 157.170 386.130 157.580 387.170 ;
        RECT 165.050 387.110 168.940 389.080 ;
        RECT 179.140 388.780 179.490 388.930 ;
        RECT 179.130 387.830 179.500 388.780 ;
        RECT 177.350 387.460 181.250 387.830 ;
        RECT 165.230 386.660 167.600 387.110 ;
        RECT 129.690 385.520 154.060 385.540 ;
        RECT 129.630 385.130 154.060 385.520 ;
        RECT 129.630 381.440 130.040 385.130 ;
        RECT 153.090 382.860 154.430 383.310 ;
        RECT 156.230 382.860 158.590 386.130 ;
        RECT 165.260 385.540 166.210 386.660 ;
        RECT 166.960 386.640 167.540 386.660 ;
        RECT 177.340 386.000 181.250 387.460 ;
        RECT 188.570 386.810 192.700 387.210 ;
        RECT 188.570 386.720 192.710 386.810 ;
        RECT 167.630 385.990 181.250 386.000 ;
        RECT 166.960 385.540 181.250 385.990 ;
        RECT 192.180 385.820 192.710 386.720 ;
        RECT 162.860 385.530 183.150 385.540 ;
        RECT 162.800 385.520 183.150 385.530 ;
        RECT 162.800 385.430 184.090 385.520 ;
        RECT 162.800 385.130 190.310 385.430 ;
        RECT 165.260 384.700 166.210 385.130 ;
        RECT 165.490 382.860 166.210 384.700 ;
        RECT 153.090 382.440 166.610 382.860 ;
        RECT 153.090 382.300 154.430 382.440 ;
        RECT 129.460 381.240 130.040 381.440 ;
        RECT 147.680 381.700 150.450 381.940 ;
        RECT 129.400 380.930 130.040 381.240 ;
        RECT 130.810 380.930 131.840 381.240 ;
        RECT 129.630 380.410 130.040 380.930 ;
        RECT 129.450 380.140 130.040 380.410 ;
        RECT 130.140 380.140 130.460 380.380 ;
        RECT 130.860 380.140 131.120 380.420 ;
        RECT 129.410 379.480 131.160 380.140 ;
        RECT 129.450 379.220 130.040 379.480 ;
        RECT 130.140 379.220 130.460 379.480 ;
        RECT 130.880 379.240 131.140 379.480 ;
        RECT 129.630 378.710 130.040 379.220 ;
        RECT 129.470 378.190 130.040 378.710 ;
        RECT 129.450 377.870 130.040 378.190 ;
        RECT 131.600 378.160 131.840 380.930 ;
        RECT 147.680 380.610 147.920 381.700 ;
        RECT 147.680 380.350 147.910 380.610 ;
        RECT 147.670 380.130 147.910 380.350 ;
        RECT 131.980 379.630 132.300 379.950 ;
        RECT 132.030 379.400 132.260 379.630 ;
        RECT 128.500 377.420 128.760 377.740 ;
        RECT 128.510 376.240 128.750 377.420 ;
        RECT 129.470 377.300 130.040 377.870 ;
        RECT 131.560 377.620 131.880 377.940 ;
        RECT 147.680 377.810 147.920 378.450 ;
        RECT 147.680 377.550 147.910 377.810 ;
        RECT 129.630 376.880 130.040 377.300 ;
        RECT 147.670 376.900 147.910 377.550 ;
        RECT 130.120 376.630 130.440 376.740 ;
        RECT 129.250 376.420 130.440 376.630 ;
        RECT 131.550 376.440 131.870 376.760 ;
        RECT 129.250 376.240 130.410 376.420 ;
        RECT 128.510 376.160 131.100 376.240 ;
        RECT 128.510 375.840 131.280 376.160 ;
        RECT 131.700 375.840 132.020 376.160 ;
        RECT 128.510 375.470 131.100 375.840 ;
        RECT 132.410 375.830 132.730 376.150 ;
        RECT 128.510 375.200 128.750 375.470 ;
        RECT 128.420 374.720 128.840 375.200 ;
        RECT 129.250 374.720 130.410 375.470 ;
        RECT 134.310 374.720 134.600 376.650 ;
        RECT 147.670 376.260 147.920 376.900 ;
        RECT 147.670 374.720 147.910 376.260 ;
        RECT 150.210 374.720 150.450 381.700 ;
        RECT 156.230 381.640 158.590 382.440 ;
        RECT 153.520 381.370 158.590 381.640 ;
        RECT 153.520 380.390 153.790 381.370 ;
        RECT 153.530 378.180 153.790 378.200 ;
        RECT 153.490 374.720 153.800 378.180 ;
        RECT 156.230 377.630 158.590 381.370 ;
        RECT 165.490 379.190 166.610 382.440 ;
        RECT 166.960 381.130 190.310 385.130 ;
        RECT 191.080 384.010 191.650 384.020 ;
        RECT 166.960 380.850 181.250 381.130 ;
        RECT 170.000 379.950 170.420 380.850 ;
        RECT 170.000 379.470 170.470 379.950 ;
        RECT 177.340 379.300 181.250 380.850 ;
        RECT 165.490 379.030 166.630 379.190 ;
        RECT 166.150 378.710 166.630 379.030 ;
        RECT 177.320 378.530 181.270 379.300 ;
        RECT 156.110 376.810 158.590 377.630 ;
        RECT 179.210 377.060 179.940 378.530 ;
        RECT 156.280 374.720 156.550 376.810 ;
        RECT 157.450 375.770 157.700 376.810 ;
        RECT 157.450 375.590 157.710 375.770 ;
        RECT 129.250 373.590 156.610 374.720 ;
        RECT 129.250 373.390 156.800 373.590 ;
        RECT 134.290 373.290 134.700 373.390 ;
        RECT 147.670 372.600 147.910 373.390 ;
        RECT 147.620 372.260 147.960 372.600 ;
        RECT 150.210 371.230 150.450 373.390 ;
        RECT 153.490 372.200 153.800 373.390 ;
        RECT 153.410 371.830 153.800 372.200 ;
        RECT 155.280 371.990 156.610 373.390 ;
        RECT 157.450 372.690 157.700 375.590 ;
        RECT 157.410 372.330 157.740 372.690 ;
        RECT 156.280 371.690 156.550 371.990 ;
        RECT 156.240 371.380 156.580 371.690 ;
        RECT 150.160 370.910 150.500 371.230 ;
        RECT 179.370 366.670 179.540 377.060 ;
        RECT 184.370 376.530 185.340 381.130 ;
        RECT 191.080 380.590 191.700 384.010 ;
        RECT 191.080 380.580 191.650 380.590 ;
        RECT 184.350 376.060 185.360 376.530 ;
      LAYER via ;
        RECT 165.450 386.810 167.480 387.140 ;
        RECT 130.180 385.220 153.980 385.480 ;
        RECT 165.390 385.950 166.090 386.570 ;
        RECT 188.840 386.810 191.830 387.160 ;
        RECT 192.270 386.010 192.620 386.770 ;
        RECT 162.860 385.220 183.720 385.480 ;
        RECT 129.460 381.150 129.720 381.410 ;
        RECT 129.450 380.120 129.710 380.380 ;
        RECT 130.170 380.090 130.430 380.350 ;
        RECT 130.860 380.130 131.120 380.390 ;
        RECT 129.450 379.670 129.710 379.930 ;
        RECT 130.860 379.690 131.120 379.950 ;
        RECT 129.450 379.250 129.710 379.510 ;
        RECT 130.170 379.250 130.430 379.510 ;
        RECT 130.880 379.270 131.140 379.530 ;
        RECT 132.010 379.660 132.270 379.920 ;
        RECT 129.450 377.900 129.710 378.160 ;
        RECT 128.500 377.450 128.760 377.710 ;
        RECT 131.590 377.650 131.850 377.910 ;
        RECT 130.150 376.450 130.410 376.710 ;
        RECT 131.580 376.470 131.840 376.730 ;
        RECT 129.360 375.870 129.620 376.130 ;
        RECT 130.290 375.870 130.550 376.130 ;
        RECT 130.990 375.870 131.250 376.130 ;
        RECT 131.730 375.870 131.990 376.130 ;
        RECT 132.440 375.860 132.700 376.120 ;
        RECT 128.420 374.750 128.840 375.170 ;
        RECT 170.030 379.500 170.450 379.920 ;
        RECT 166.180 378.740 166.600 379.160 ;
        RECT 179.240 377.100 179.680 377.540 ;
        RECT 134.370 373.350 134.660 373.930 ;
        RECT 147.660 372.290 147.920 372.550 ;
        RECT 153.450 371.860 153.760 372.170 ;
        RECT 157.450 372.400 157.710 372.660 ;
        RECT 156.280 371.410 156.550 371.670 ;
        RECT 150.200 370.940 150.460 371.200 ;
        RECT 191.240 380.720 191.660 383.890 ;
        RECT 184.380 376.100 185.330 376.510 ;
    END
  END ANALOG06
  PIN ANALOG05
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 193.640 387.110 197.530 389.080 ;
        RECT 193.820 386.660 196.190 387.110 ;
        RECT 217.160 386.810 221.290 387.210 ;
        RECT 217.160 386.720 221.300 386.810 ;
        RECT 193.850 384.700 194.800 386.660 ;
        RECT 195.550 386.640 196.130 386.660 ;
        RECT 220.770 385.820 221.300 386.720 ;
        RECT 194.080 379.030 194.800 384.700 ;
      LAYER via ;
        RECT 194.040 386.810 196.070 387.140 ;
        RECT 217.430 386.810 220.420 387.160 ;
        RECT 193.980 385.950 194.680 386.570 ;
        RECT 220.860 386.010 221.210 386.770 ;
    END
  END ANALOG05
  PIN ANALOG04
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 222.240 387.110 226.130 389.080 ;
        RECT 222.410 386.660 224.780 387.110 ;
        RECT 245.750 386.810 249.880 387.210 ;
        RECT 245.750 386.720 249.890 386.810 ;
        RECT 222.440 384.700 223.390 386.660 ;
        RECT 224.140 386.640 224.720 386.660 ;
        RECT 249.360 385.820 249.890 386.720 ;
        RECT 222.670 379.030 223.390 384.700 ;
      LAYER via ;
        RECT 222.630 386.810 224.660 387.140 ;
        RECT 246.020 386.810 249.010 387.160 ;
        RECT 222.570 385.950 223.270 386.570 ;
        RECT 249.450 386.010 249.800 386.770 ;
    END
  END ANALOG04
  PIN ANALOG03
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 250.830 387.110 254.720 389.080 ;
        RECT 251.000 386.660 253.370 387.110 ;
        RECT 274.340 386.810 278.470 387.210 ;
        RECT 274.340 386.720 278.480 386.810 ;
        RECT 251.030 384.700 251.980 386.660 ;
        RECT 252.730 386.640 253.310 386.660 ;
        RECT 277.950 385.820 278.480 386.720 ;
        RECT 251.260 379.030 251.980 384.700 ;
      LAYER via ;
        RECT 251.220 386.810 253.250 387.140 ;
        RECT 274.610 386.810 277.600 387.160 ;
        RECT 251.160 385.950 251.860 386.570 ;
        RECT 278.040 386.010 278.390 386.770 ;
    END
  END ANALOG03
  PIN ANALOG02
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 279.420 387.910 283.310 389.080 ;
        RECT 279.410 387.110 283.300 387.910 ;
        RECT 279.590 386.660 281.960 387.110 ;
        RECT 302.930 386.810 307.060 387.210 ;
        RECT 302.930 386.720 307.070 386.810 ;
        RECT 279.620 384.700 280.570 386.660 ;
        RECT 281.320 386.640 281.900 386.660 ;
        RECT 306.540 385.820 307.070 386.720 ;
        RECT 279.850 379.030 280.570 384.700 ;
      LAYER via ;
        RECT 279.810 386.810 281.840 387.140 ;
        RECT 303.200 386.810 306.190 387.160 ;
        RECT 279.750 385.950 280.450 386.570 ;
        RECT 306.630 386.010 306.980 386.770 ;
    END
  END ANALOG02
  PIN ANALOG01
    ANTENNADIFFAREA 48.993099 ;
    PORT
      LAYER met1 ;
        RECT 308.010 387.910 311.900 389.070 ;
        RECT 308.000 387.900 311.900 387.910 ;
        RECT 308.000 387.110 311.890 387.900 ;
        RECT 308.180 386.660 310.550 387.110 ;
        RECT 331.520 386.810 335.650 387.210 ;
        RECT 331.520 386.720 335.660 386.810 ;
        RECT 308.210 384.700 309.160 386.660 ;
        RECT 309.910 386.640 310.490 386.660 ;
        RECT 335.130 385.820 335.660 386.720 ;
        RECT 308.440 379.030 309.160 384.700 ;
      LAYER via ;
        RECT 308.400 386.810 310.430 387.140 ;
        RECT 331.790 386.810 334.780 387.160 ;
        RECT 308.340 385.950 309.040 386.570 ;
        RECT 335.220 386.010 335.570 386.770 ;
    END
  END ANALOG01
  PIN VSSA1
    PORT
      LAYER met2 ;
        RECT 4.380 0.330 5.780 2.300 ;
    END
    PORT
      LAYER met2 ;
        RECT 368.290 173.390 369.030 173.730 ;
        RECT 367.630 172.990 369.040 173.390 ;
        RECT 367.650 172.300 369.030 172.990 ;
        RECT 367.640 171.130 369.040 172.300 ;
    END
  END VSSA1
  PIN VDDA1
    PORT
      LAYER met2 ;
        RECT 10.680 0.000 12.080 3.660 ;
    END
    PORT
      LAYER met2 ;
        RECT 361.310 172.360 362.710 173.140 ;
        RECT 361.300 172.240 362.710 172.360 ;
        RECT 361.290 172.090 362.710 172.240 ;
        RECT 361.290 171.190 362.700 172.090 ;
    END
  END VDDA1
  PIN LADATAOUT01
    PORT
      LAYER met2 ;
        RECT 146.280 6.780 148.300 301.800 ;
        RECT 146.280 5.220 148.310 6.780 ;
        RECT 146.280 5.210 148.300 5.220 ;
    END
  END LADATAOUT01
  PIN LADATAOUT00
    PORT
      LAYER met2 ;
        RECT 142.220 5.210 144.240 301.800 ;
    END
  END LADATAOUT00
  PIN LADATAOUT02
    PORT
      LAYER met2 ;
        RECT 150.250 6.770 152.270 301.800 ;
        RECT 150.240 5.210 152.270 6.770 ;
    END
  END LADATAOUT02
  PIN LADATAOUT03
    PORT
      LAYER met2 ;
        RECT 154.250 6.770 156.270 301.800 ;
        RECT 154.240 5.210 156.270 6.770 ;
    END
  END LADATAOUT03
  PIN LADATAOUT04
    PORT
      LAYER met2 ;
        RECT 158.300 5.210 160.320 301.800 ;
    END
  END LADATAOUT04
  PIN LADATAOUT05
    PORT
      LAYER met2 ;
        RECT 162.310 6.780 164.330 301.800 ;
        RECT 162.300 5.220 164.330 6.780 ;
        RECT 162.310 5.210 164.330 5.220 ;
    END
  END LADATAOUT05
  PIN LADATAOUT06
    PORT
      LAYER met2 ;
        RECT 166.310 5.210 168.330 301.800 ;
    END
  END LADATAOUT06
  PIN LADATAOUT07
    PORT
      LAYER met2 ;
        RECT 170.400 5.210 172.420 301.800 ;
    END
  END LADATAOUT07
  PIN LADATAOUT08
    PORT
      LAYER met2 ;
        RECT 174.530 6.770 176.550 301.800 ;
        RECT 174.520 5.210 176.550 6.770 ;
    END
  END LADATAOUT08
  PIN LADATAOUT09
    PORT
      LAYER met2 ;
        RECT 178.530 6.770 180.550 301.800 ;
        RECT 178.520 5.210 180.550 6.770 ;
    END
  END LADATAOUT09
  PIN LADATAOUT10
    PORT
      LAYER met2 ;
        RECT 182.490 6.770 184.510 301.800 ;
        RECT 182.480 5.210 184.510 6.770 ;
    END
  END LADATAOUT10
  PIN LADATAOUT11
    PORT
      LAYER met2 ;
        RECT 186.540 6.780 188.560 301.800 ;
        RECT 186.540 5.220 188.570 6.780 ;
        RECT 186.540 5.210 188.560 5.220 ;
    END
  END LADATAOUT11
  PIN LADATAOUT12
    PORT
      LAYER met2 ;
        RECT 190.630 5.210 192.650 301.800 ;
    END
  END LADATAOUT12
  PIN LADATAOUT13
    PORT
      LAYER met2 ;
        RECT 194.640 6.760 196.660 301.800 ;
        RECT 194.640 5.210 196.670 6.760 ;
        RECT 194.650 5.200 196.670 5.210 ;
    END
  END LADATAOUT13
  PIN LADATAOUT14
    PORT
      LAYER met2 ;
        RECT 198.680 6.770 200.700 301.800 ;
        RECT 198.680 5.210 200.710 6.770 ;
    END
  END LADATAOUT14
  PIN LADATAOUT15
    PORT
      LAYER met2 ;
        RECT 202.770 6.750 204.790 301.800 ;
        RECT 202.770 5.210 204.800 6.750 ;
        RECT 202.780 5.190 204.800 5.210 ;
    END
  END LADATAOUT15
  PIN LADATA16
    PORT
      LAYER met2 ;
        RECT 206.820 5.210 208.840 301.800 ;
    END
  END LADATA16
  PIN LADATAOUT17
    PORT
      LAYER met2 ;
        RECT 210.790 5.210 212.810 301.800 ;
    END
  END LADATAOUT17
  PIN LADATAOUT18
    PORT
      LAYER met2 ;
        RECT 214.910 5.210 216.930 301.800 ;
    END
  END LADATAOUT18
  PIN LADATAOUT19
    PORT
      LAYER met2 ;
        RECT 219.040 5.200 221.060 301.800 ;
    END
  END LADATAOUT19
  PIN LADATAOUT20
    PORT
      LAYER met2 ;
        RECT 223.050 5.210 225.070 301.800 ;
    END
  END LADATAOUT20
  PIN LADATAOUT21
    PORT
      LAYER met2 ;
        RECT 227.060 6.890 229.080 301.800 ;
        RECT 227.060 5.230 229.100 6.890 ;
    END
  END LADATAOUT21
  PIN LADATAOUT22
    PORT
      LAYER met2 ;
        RECT 231.150 6.870 233.170 301.800 ;
        RECT 231.150 5.210 233.180 6.870 ;
    END
  END LADATAOUT22
  PIN LADATAOUT23
    PORT
      LAYER met2 ;
        RECT 235.320 5.210 237.340 301.800 ;
    END
  END LADATAOUT23
  PIN LADATAOUT24
    PORT
      LAYER met2 ;
        RECT 239.320 6.870 241.340 301.800 ;
        RECT 239.320 5.210 241.350 6.870 ;
    END
  END LADATAOUT24
  PIN LADATAIN00
    PORT
      LAYER met2 ;
        RECT 243.330 6.870 245.350 301.800 ;
        RECT 243.300 5.210 245.350 6.870 ;
    END
  END LADATAIN00
  PIN LADATAIN01
    PORT
      LAYER met2 ;
        RECT 247.290 6.870 249.310 301.800 ;
        RECT 247.280 5.210 249.310 6.870 ;
    END
  END LADATAIN01
  PIN LADATAIN02
    PORT
      LAYER met2 ;
        RECT 251.340 6.870 253.360 301.800 ;
        RECT 251.340 5.210 253.380 6.870 ;
    END
  END LADATAIN02
  PIN LADATAIN03
    PORT
      LAYER met2 ;
        RECT 255.400 6.870 257.420 301.800 ;
        RECT 255.400 5.210 257.440 6.870 ;
    END
  END LADATAIN03
  PIN VCCA
    ANTENNAGATEAREA 0.354000 ;
    ANTENNADIFFAREA 4.549800 ;
    PORT
      LAYER nwell ;
        RECT 191.100 347.810 193.650 347.820 ;
        RECT 191.090 344.000 193.650 347.810 ;
        RECT 195.180 344.000 197.410 347.820 ;
        RECT 191.090 343.990 197.410 344.000 ;
        RECT 191.090 343.840 193.760 343.990 ;
        RECT 191.090 343.830 193.940 343.840 ;
        RECT 191.090 341.790 193.760 343.830 ;
        RECT 191.100 341.780 193.760 341.790 ;
        RECT 193.240 340.920 193.760 341.780 ;
        RECT 195.180 341.770 197.410 343.990 ;
        RECT 193.350 337.960 193.760 340.920 ;
      LAYER met2 ;
        RECT 243.670 356.810 267.000 357.240 ;
        RECT 193.250 343.880 193.560 343.900 ;
        RECT 191.090 343.720 201.160 343.880 ;
        RECT 191.090 343.710 201.150 343.720 ;
        RECT 191.090 343.700 193.650 343.710 ;
        RECT 193.250 343.570 193.560 343.700 ;
        RECT 196.510 343.690 196.830 343.710 ;
        RECT 196.510 343.500 204.430 343.690 ;
        RECT 204.590 343.500 204.900 343.540 ;
        RECT 196.510 343.480 204.900 343.500 ;
        RECT 196.510 343.450 196.830 343.480 ;
        RECT 204.220 343.290 204.900 343.480 ;
        RECT 204.590 343.210 204.900 343.290 ;
        RECT 193.240 343.020 193.390 343.070 ;
        RECT 193.240 342.900 193.560 343.020 ;
        RECT 193.240 342.890 201.160 342.900 ;
        RECT 191.090 342.730 201.160 342.890 ;
        RECT 191.090 342.710 193.650 342.730 ;
        RECT 193.240 342.690 193.560 342.710 ;
        RECT 193.240 342.560 193.390 342.690 ;
        RECT 196.490 342.560 196.810 342.660 ;
        RECT 198.830 342.640 200.370 342.730 ;
        RECT 193.240 342.460 196.810 342.560 ;
        RECT 191.090 342.400 196.810 342.460 ;
        RECT 191.090 342.370 193.660 342.400 ;
        RECT 198.740 342.370 199.060 342.420 ;
        RECT 191.090 342.280 199.060 342.370 ;
        RECT 192.670 342.210 199.060 342.280 ;
        RECT 193.250 342.160 193.560 342.210 ;
        RECT 198.740 342.160 199.060 342.210 ;
        RECT 193.220 342.140 193.560 342.160 ;
        RECT 193.220 341.900 193.540 342.140 ;
        RECT 193.290 341.890 193.460 341.900 ;
        RECT 198.220 341.440 198.540 341.490 ;
        RECT 192.680 341.420 198.540 341.440 ;
        RECT 192.680 341.390 204.020 341.420 ;
        RECT 192.680 341.280 204.080 341.390 ;
        RECT 196.450 341.220 204.080 341.280 ;
        RECT 204.590 341.220 204.900 341.300 ;
        RECT 193.200 341.120 193.520 341.150 ;
        RECT 196.450 341.120 196.690 341.220 ;
        RECT 193.200 340.940 196.690 341.120 ;
        RECT 203.890 341.020 204.900 341.220 ;
        RECT 204.490 341.010 204.900 341.020 ;
        RECT 204.590 340.970 204.900 341.010 ;
        RECT 193.200 340.920 196.610 340.940 ;
        RECT 193.200 340.890 193.520 340.920 ;
        RECT 196.490 340.740 196.810 340.780 ;
        RECT 196.490 340.720 204.040 340.740 ;
        RECT 204.590 340.730 204.900 340.770 ;
        RECT 204.490 340.720 204.900 340.730 ;
        RECT 196.490 340.520 204.900 340.720 ;
        RECT 196.590 340.510 196.910 340.520 ;
        RECT 204.590 340.440 204.900 340.520 ;
        RECT 193.180 339.600 193.380 340.060 ;
        RECT 197.750 339.600 198.070 339.650 ;
        RECT 192.670 339.440 198.070 339.600 ;
        RECT 193.180 339.360 196.730 339.440 ;
        RECT 197.750 339.390 198.070 339.440 ;
        RECT 196.330 339.340 196.650 339.360 ;
        RECT 198.720 333.210 254.550 333.250 ;
        RECT 198.720 332.750 255.260 333.210 ;
        RECT 249.160 332.350 251.170 332.370 ;
        RECT 198.180 331.850 251.170 332.350 ;
        RECT 197.710 331.430 246.980 331.450 ;
        RECT 197.710 330.950 247.090 331.430 ;
        RECT 245.080 330.890 247.090 330.950 ;
        RECT 249.160 330.890 251.170 331.850 ;
        RECT 253.250 330.890 255.260 332.750 ;
        RECT 243.490 328.800 333.540 330.890 ;
        RECT 245.080 327.580 247.090 328.800 ;
        RECT 249.160 327.580 251.170 328.800 ;
        RECT 253.250 327.580 255.260 328.800 ;
        RECT 264.460 327.580 268.990 327.660 ;
        RECT 243.770 326.430 269.060 327.580 ;
        RECT 245.080 325.380 247.090 326.430 ;
        RECT 249.160 325.380 251.170 326.430 ;
        RECT 253.250 325.380 255.260 326.430 ;
        RECT 264.460 326.410 268.990 326.430 ;
        RECT 243.810 323.290 329.300 325.380 ;
        RECT 245.080 312.750 247.090 323.290 ;
        RECT 245.080 312.100 247.150 312.750 ;
        RECT 249.160 312.730 251.170 323.290 ;
        RECT 253.250 312.750 255.260 323.290 ;
        RECT 245.080 312.060 247.090 312.100 ;
        RECT 249.160 312.080 251.200 312.730 ;
        RECT 253.220 312.170 255.260 312.750 ;
        RECT 253.220 312.100 255.250 312.170 ;
        RECT 249.160 312.000 251.170 312.080 ;
        RECT 327.210 191.860 329.300 323.290 ;
        RECT 331.450 218.330 333.540 328.800 ;
        RECT 331.280 214.620 333.710 218.330 ;
        RECT 327.220 189.960 329.300 191.860 ;
        RECT 327.220 189.840 329.310 189.960 ;
        RECT 327.110 189.780 329.310 189.840 ;
        RECT 326.850 186.100 329.380 189.780 ;
        RECT 327.110 186.080 329.200 186.100 ;
        RECT 263.620 164.230 268.220 165.010 ;
        RECT 263.620 162.550 362.770 164.230 ;
        RECT 263.620 161.260 362.900 162.550 ;
        RECT 263.620 160.440 268.220 161.260 ;
    END
  END VCCA
  OBS
      LAYER nwell ;
        RECT 38.460 380.440 50.510 386.380 ;
        RECT 67.050 380.440 79.100 386.380 ;
        RECT 95.640 380.440 107.690 386.380 ;
        RECT 140.280 362.510 142.850 365.600 ;
        RECT 163.860 364.570 165.630 370.810 ;
        RECT 169.590 364.570 172.100 370.810 ;
        RECT 210.230 366.760 212.950 368.410 ;
        RECT 210.230 366.720 212.940 366.760 ;
        RECT 210.230 365.390 212.940 365.430 ;
        RECT 210.230 365.330 212.950 365.390 ;
        RECT 209.140 365.320 212.950 365.330 ;
        RECT 209.340 365.010 209.660 365.310 ;
        RECT 210.230 363.740 212.950 365.320 ;
        RECT 164.700 363.560 164.940 363.610 ;
        RECT 164.460 363.550 165.930 363.560 ;
        RECT 164.160 363.470 165.930 363.550 ;
        RECT 170.190 363.470 172.400 363.560 ;
        RECT 178.340 363.310 179.020 363.320 ;
        RECT 163.860 356.210 165.630 362.450 ;
        RECT 169.590 356.210 172.100 362.450 ;
        RECT 178.330 357.260 179.030 363.310 ;
        RECT 202.230 360.160 202.790 360.700 ;
        RECT 209.150 358.620 209.220 358.800 ;
        RECT 190.520 357.200 193.070 357.210 ;
        RECT 163.860 346.080 165.630 352.320 ;
        RECT 169.590 346.080 172.100 352.320 ;
        RECT 185.420 347.250 188.840 353.300 ;
        RECT 190.510 351.180 193.070 357.200 ;
        RECT 190.520 351.170 193.070 351.180 ;
        RECT 194.600 351.160 196.830 357.210 ;
        RECT 198.850 355.350 200.580 357.210 ;
        RECT 198.850 353.510 200.590 355.350 ;
        RECT 209.150 353.750 209.230 353.930 ;
        RECT 198.850 351.160 200.580 353.510 ;
        RECT 209.590 351.160 211.820 357.210 ;
        RECT 199.430 347.190 201.160 347.820 ;
        RECT 199.430 344.120 201.170 347.190 ;
        RECT 199.040 343.900 199.420 344.000 ;
        RECT 138.890 338.290 141.260 341.160 ;
        RECT 163.860 336.310 165.630 342.550 ;
        RECT 178.330 337.510 180.080 343.510 ;
        RECT 185.420 337.490 188.840 343.540 ;
        RECT 199.430 341.770 201.160 344.120 ;
        RECT 203.070 343.860 203.470 344.000 ;
        RECT 180.230 332.110 182.250 336.070 ;
        RECT 180.230 332.080 184.270 332.110 ;
        RECT 138.550 327.630 138.560 327.670 ;
        RECT 139.560 324.630 142.950 330.330 ;
        RECT 171.070 326.380 174.460 332.080 ;
        RECT 175.460 329.040 175.470 329.080 ;
        RECT 177.230 329.040 177.240 329.080 ;
        RECT 178.240 326.410 184.270 332.080 ;
        RECT 185.270 329.070 185.280 329.110 ;
        RECT 187.040 329.070 187.050 329.110 ;
        RECT 188.050 326.410 191.440 332.110 ;
        RECT 178.240 326.380 181.630 326.410 ;
        RECT 221.980 309.980 227.630 326.080 ;
      LAYER li1 ;
        RECT 31.320 387.460 31.570 388.920 ;
        RECT 31.360 387.450 31.530 387.460 ;
        RECT 38.000 387.430 38.250 388.900 ;
        RECT 59.910 387.460 60.160 388.920 ;
        RECT 59.950 387.450 60.120 387.460 ;
        RECT 66.590 387.430 66.840 388.900 ;
        RECT 88.500 387.460 88.750 388.920 ;
        RECT 88.540 387.450 88.710 387.460 ;
        RECT 95.180 387.430 95.430 388.900 ;
        RECT 172.520 387.460 172.770 388.920 ;
        RECT 172.560 387.450 172.730 387.460 ;
        RECT 179.200 387.430 179.450 388.900 ;
        RECT 201.110 387.460 201.360 388.920 ;
        RECT 201.150 387.450 201.320 387.460 ;
        RECT 207.790 387.430 208.040 388.900 ;
        RECT 229.700 387.460 229.950 388.920 ;
        RECT 229.740 387.450 229.910 387.460 ;
        RECT 236.380 387.430 236.630 388.900 ;
        RECT 258.290 387.460 258.540 388.920 ;
        RECT 258.330 387.450 258.500 387.460 ;
        RECT 264.970 387.430 265.220 388.900 ;
        RECT 286.880 387.460 287.130 388.920 ;
        RECT 286.920 387.450 287.090 387.460 ;
        RECT 293.560 387.430 293.810 388.900 ;
        RECT 315.470 387.460 315.720 388.920 ;
        RECT 315.510 387.450 315.680 387.460 ;
        RECT 322.150 387.430 322.400 388.900 ;
        RECT 344.060 387.460 344.310 388.920 ;
        RECT 344.100 387.450 344.270 387.460 ;
        RECT 350.740 387.430 350.990 388.900 ;
        RECT 24.140 386.710 51.520 387.220 ;
        RECT 24.140 384.780 24.940 386.710 ;
        RECT 25.520 386.260 25.690 386.340 ;
        RECT 36.760 386.260 36.990 386.350 ;
        RECT 25.520 386.250 36.990 386.260 ;
        RECT 2.180 380.170 9.710 380.720 ;
        RECT 0.500 367.200 1.970 367.450 ;
        RECT 2.180 367.260 2.690 380.170 ;
        RECT 9.040 380.160 9.710 380.170 ;
        RECT 5.340 379.270 8.800 379.710 ;
        RECT 3.410 379.170 8.800 379.270 ;
        RECT 3.410 379.100 8.690 379.170 ;
        RECT 3.410 368.190 3.580 379.100 ;
        RECT 3.910 378.690 8.140 378.710 ;
        RECT 3.890 368.580 8.220 378.690 ;
        RECT 3.950 368.530 4.120 368.580 ;
        RECT 8.520 368.190 8.690 379.100 ;
        RECT 3.410 368.020 8.690 368.190 ;
        RECT 8.450 368.010 8.690 368.020 ;
        RECT 9.200 367.260 9.710 380.160 ;
        RECT 24.140 380.200 24.650 384.780 ;
        RECT 25.510 380.780 36.990 386.250 ;
        RECT 25.440 380.610 36.990 380.780 ;
        RECT 25.510 380.550 25.700 380.610 ;
        RECT 36.760 380.370 36.990 380.610 ;
        RECT 25.390 380.200 27.190 380.210 ;
        RECT 37.550 380.200 38.060 386.710 ;
        RECT 38.820 385.820 50.070 385.990 ;
        RECT 38.820 380.950 38.990 385.820 ;
        RECT 39.380 385.490 49.490 385.510 ;
        RECT 39.380 385.450 49.510 385.490 ;
        RECT 39.330 385.280 49.510 385.450 ;
        RECT 39.380 381.260 49.510 385.280 ;
        RECT 49.900 384.060 50.070 385.820 ;
        RECT 39.380 381.180 49.490 381.260 ;
        RECT 38.810 380.880 38.990 380.950 ;
        RECT 49.900 380.880 50.510 384.060 ;
        RECT 38.810 380.710 50.510 380.880 ;
        RECT 49.970 380.600 50.510 380.710 ;
        RECT 50.970 380.360 51.520 386.710 ;
        RECT 50.960 380.200 51.520 380.360 ;
        RECT 24.140 379.860 51.520 380.200 ;
        RECT 52.730 386.710 80.110 387.220 ;
        RECT 52.730 384.780 53.530 386.710 ;
        RECT 54.110 386.260 54.280 386.340 ;
        RECT 65.350 386.260 65.580 386.350 ;
        RECT 54.110 386.250 65.580 386.260 ;
        RECT 52.730 380.200 53.240 384.780 ;
        RECT 54.100 380.780 65.580 386.250 ;
        RECT 54.030 380.610 65.580 380.780 ;
        RECT 54.100 380.550 54.290 380.610 ;
        RECT 65.350 380.370 65.580 380.610 ;
        RECT 53.980 380.200 55.780 380.210 ;
        RECT 66.140 380.200 66.650 386.710 ;
        RECT 67.410 385.820 78.660 385.990 ;
        RECT 67.410 380.950 67.580 385.820 ;
        RECT 67.970 385.490 78.080 385.510 ;
        RECT 67.970 385.450 78.100 385.490 ;
        RECT 67.920 385.280 78.100 385.450 ;
        RECT 67.970 381.260 78.100 385.280 ;
        RECT 78.490 384.060 78.660 385.820 ;
        RECT 67.970 381.180 78.080 381.260 ;
        RECT 67.400 380.880 67.580 380.950 ;
        RECT 78.490 380.880 79.100 384.060 ;
        RECT 67.400 380.710 79.100 380.880 ;
        RECT 78.560 380.600 79.100 380.710 ;
        RECT 79.560 380.360 80.110 386.710 ;
        RECT 79.550 380.200 80.110 380.360 ;
        RECT 52.730 379.860 80.110 380.200 ;
        RECT 81.320 386.710 108.700 387.220 ;
        RECT 81.320 384.780 82.120 386.710 ;
        RECT 82.700 386.260 82.870 386.340 ;
        RECT 93.940 386.260 94.170 386.350 ;
        RECT 82.700 386.250 94.170 386.260 ;
        RECT 81.320 380.200 81.830 384.780 ;
        RECT 82.690 380.780 94.170 386.250 ;
        RECT 82.620 380.610 94.170 380.780 ;
        RECT 82.690 380.550 82.880 380.610 ;
        RECT 93.940 380.370 94.170 380.610 ;
        RECT 82.570 380.200 84.370 380.210 ;
        RECT 94.730 380.200 95.240 386.710 ;
        RECT 96.000 385.820 107.250 385.990 ;
        RECT 96.000 380.950 96.170 385.820 ;
        RECT 96.560 385.490 106.670 385.510 ;
        RECT 96.560 385.450 106.690 385.490 ;
        RECT 96.510 385.280 106.690 385.450 ;
        RECT 96.560 381.260 106.690 385.280 ;
        RECT 107.080 384.060 107.250 385.820 ;
        RECT 96.560 381.180 106.670 381.260 ;
        RECT 95.990 380.880 96.170 380.950 ;
        RECT 107.080 380.880 107.690 384.060 ;
        RECT 95.990 380.710 107.690 380.880 ;
        RECT 107.150 380.600 107.690 380.710 ;
        RECT 108.150 380.360 108.700 386.710 ;
        RECT 150.500 385.930 150.720 387.050 ;
        RECT 150.450 385.740 150.780 385.930 ;
        RECT 157.240 385.740 157.480 387.090 ;
        RECT 165.340 386.710 192.720 387.220 ;
        RECT 165.340 385.540 166.140 386.710 ;
        RECT 166.720 386.260 166.890 386.340 ;
        RECT 177.960 386.260 178.190 386.350 ;
        RECT 166.720 386.250 178.190 386.260 ;
        RECT 166.710 385.540 178.190 386.250 ;
        RECT 178.750 385.540 179.260 386.710 ;
        RECT 180.020 385.820 191.270 385.990 ;
        RECT 180.020 385.540 180.190 385.820 ;
        RECT 129.740 385.510 184.480 385.540 ;
        RECT 129.740 385.490 190.690 385.510 ;
        RECT 129.740 385.270 190.710 385.490 ;
        RECT 129.740 385.140 154.080 385.270 ;
        RECT 162.770 385.140 190.710 385.270 ;
        RECT 128.920 381.170 129.090 381.470 ;
        RECT 129.740 381.170 129.910 385.140 ;
        RECT 165.340 384.780 166.140 385.140 ;
        RECT 128.920 380.990 129.920 381.170 ;
        RECT 130.320 381.160 130.490 381.470 ;
        RECT 132.120 381.200 132.790 381.370 ;
        RECT 130.320 380.990 131.330 381.160 ;
        RECT 108.140 380.200 108.700 380.360 ;
        RECT 129.740 380.310 129.910 380.990 ;
        RECT 132.120 380.410 132.790 380.580 ;
        RECT 130.130 380.310 130.450 380.350 ;
        RECT 81.320 379.860 108.700 380.200 ;
        RECT 129.250 380.140 131.330 380.310 ;
        RECT 146.140 380.270 149.450 381.250 ;
        RECT 153.540 380.450 153.770 381.140 ;
        RECT 158.240 380.400 158.470 381.090 ;
        RECT 165.340 380.200 165.850 384.780 ;
        RECT 166.710 380.780 178.190 385.140 ;
        RECT 166.640 380.610 178.190 380.780 ;
        RECT 166.710 380.550 166.900 380.610 ;
        RECT 177.960 380.370 178.190 380.610 ;
        RECT 166.590 380.200 168.390 380.210 ;
        RECT 178.750 380.200 179.260 385.140 ;
        RECT 180.020 380.950 180.190 385.140 ;
        RECT 180.580 381.260 190.710 385.140 ;
        RECT 191.100 384.060 191.270 385.820 ;
        RECT 180.580 381.180 190.690 381.260 ;
        RECT 180.010 380.880 180.190 380.950 ;
        RECT 184.310 380.880 184.480 381.180 ;
        RECT 191.100 380.880 191.710 384.060 ;
        RECT 180.010 380.710 191.710 380.880 ;
        RECT 184.310 380.200 184.480 380.710 ;
        RECT 191.170 380.600 191.710 380.710 ;
        RECT 192.170 380.360 192.720 386.710 ;
        RECT 192.160 380.200 192.720 380.360 ;
        RECT 129.740 379.900 129.910 380.140 ;
        RECT 130.120 380.120 130.450 380.140 ;
        RECT 130.130 380.090 130.450 380.120 ;
        RECT 24.170 379.690 51.520 379.860 ;
        RECT 52.760 379.690 80.110 379.860 ;
        RECT 81.350 379.690 108.700 379.860 ;
        RECT 129.430 379.730 131.250 379.900 ;
        RECT 24.170 379.670 24.860 379.690 ;
        RECT 25.370 379.680 27.170 379.690 ;
        RECT 52.760 379.670 53.450 379.690 ;
        RECT 53.960 379.680 55.760 379.690 ;
        RECT 81.350 379.670 82.040 379.690 ;
        RECT 82.550 379.680 84.350 379.690 ;
        RECT 129.740 379.490 129.910 379.730 ;
        RECT 130.130 379.490 130.450 379.510 ;
        RECT 129.250 379.320 131.330 379.490 ;
        RECT 132.040 379.480 132.250 379.910 ;
        RECT 146.250 379.610 146.420 379.960 ;
        RECT 165.340 379.860 192.720 380.200 ;
        RECT 193.930 386.710 221.310 387.220 ;
        RECT 193.930 384.780 194.730 386.710 ;
        RECT 195.310 386.260 195.480 386.340 ;
        RECT 206.550 386.260 206.780 386.350 ;
        RECT 195.310 386.250 206.780 386.260 ;
        RECT 193.930 380.200 194.440 384.780 ;
        RECT 195.300 380.780 206.780 386.250 ;
        RECT 195.230 380.610 206.780 380.780 ;
        RECT 195.300 380.550 195.490 380.610 ;
        RECT 206.550 380.370 206.780 380.610 ;
        RECT 195.180 380.200 196.980 380.210 ;
        RECT 207.340 380.200 207.850 386.710 ;
        RECT 208.610 385.820 219.860 385.990 ;
        RECT 208.610 380.950 208.780 385.820 ;
        RECT 209.170 385.490 219.280 385.510 ;
        RECT 209.170 385.450 219.300 385.490 ;
        RECT 209.120 385.280 219.300 385.450 ;
        RECT 209.170 381.260 219.300 385.280 ;
        RECT 219.690 384.060 219.860 385.820 ;
        RECT 209.170 381.180 219.280 381.260 ;
        RECT 208.600 380.880 208.780 380.950 ;
        RECT 219.690 380.880 220.300 384.060 ;
        RECT 208.600 380.710 220.300 380.880 ;
        RECT 219.760 380.600 220.300 380.710 ;
        RECT 220.760 380.360 221.310 386.710 ;
        RECT 220.750 380.200 221.310 380.360 ;
        RECT 193.930 379.860 221.310 380.200 ;
        RECT 222.520 386.710 249.900 387.220 ;
        RECT 222.520 384.780 223.320 386.710 ;
        RECT 223.900 386.260 224.070 386.340 ;
        RECT 235.140 386.260 235.370 386.350 ;
        RECT 223.900 386.250 235.370 386.260 ;
        RECT 222.520 380.200 223.030 384.780 ;
        RECT 223.890 380.780 235.370 386.250 ;
        RECT 223.820 380.610 235.370 380.780 ;
        RECT 223.890 380.550 224.080 380.610 ;
        RECT 235.140 380.370 235.370 380.610 ;
        RECT 223.770 380.200 225.570 380.210 ;
        RECT 235.930 380.200 236.440 386.710 ;
        RECT 237.200 385.820 248.450 385.990 ;
        RECT 237.200 380.950 237.370 385.820 ;
        RECT 237.760 385.490 247.870 385.510 ;
        RECT 237.760 385.450 247.890 385.490 ;
        RECT 237.710 385.280 247.890 385.450 ;
        RECT 237.760 381.260 247.890 385.280 ;
        RECT 248.280 384.060 248.450 385.820 ;
        RECT 237.760 381.180 247.870 381.260 ;
        RECT 237.190 380.880 237.370 380.950 ;
        RECT 248.280 380.880 248.890 384.060 ;
        RECT 237.190 380.710 248.890 380.880 ;
        RECT 248.350 380.600 248.890 380.710 ;
        RECT 249.350 380.360 249.900 386.710 ;
        RECT 249.340 380.200 249.900 380.360 ;
        RECT 222.520 379.860 249.900 380.200 ;
        RECT 251.110 386.710 278.490 387.220 ;
        RECT 251.110 384.780 251.910 386.710 ;
        RECT 252.490 386.260 252.660 386.340 ;
        RECT 263.730 386.260 263.960 386.350 ;
        RECT 252.490 386.250 263.960 386.260 ;
        RECT 251.110 380.200 251.620 384.780 ;
        RECT 252.480 380.780 263.960 386.250 ;
        RECT 252.410 380.610 263.960 380.780 ;
        RECT 252.480 380.550 252.670 380.610 ;
        RECT 263.730 380.370 263.960 380.610 ;
        RECT 252.360 380.200 254.160 380.210 ;
        RECT 264.520 380.200 265.030 386.710 ;
        RECT 265.790 385.820 277.040 385.990 ;
        RECT 265.790 380.950 265.960 385.820 ;
        RECT 266.350 385.490 276.460 385.510 ;
        RECT 266.350 385.450 276.480 385.490 ;
        RECT 266.300 385.280 276.480 385.450 ;
        RECT 266.350 381.260 276.480 385.280 ;
        RECT 276.870 384.060 277.040 385.820 ;
        RECT 266.350 381.180 276.460 381.260 ;
        RECT 265.780 380.880 265.960 380.950 ;
        RECT 276.870 380.880 277.480 384.060 ;
        RECT 265.780 380.710 277.480 380.880 ;
        RECT 276.940 380.600 277.480 380.710 ;
        RECT 277.940 380.360 278.490 386.710 ;
        RECT 277.930 380.200 278.490 380.360 ;
        RECT 251.110 379.860 278.490 380.200 ;
        RECT 279.700 386.710 307.080 387.220 ;
        RECT 279.700 384.780 280.500 386.710 ;
        RECT 281.080 386.260 281.250 386.340 ;
        RECT 292.320 386.260 292.550 386.350 ;
        RECT 281.080 386.250 292.550 386.260 ;
        RECT 279.700 380.200 280.210 384.780 ;
        RECT 281.070 380.780 292.550 386.250 ;
        RECT 281.000 380.610 292.550 380.780 ;
        RECT 281.070 380.550 281.260 380.610 ;
        RECT 292.320 380.370 292.550 380.610 ;
        RECT 280.950 380.200 282.750 380.210 ;
        RECT 293.110 380.200 293.620 386.710 ;
        RECT 294.380 385.820 305.630 385.990 ;
        RECT 294.380 380.950 294.550 385.820 ;
        RECT 294.940 385.490 305.050 385.510 ;
        RECT 294.940 385.450 305.070 385.490 ;
        RECT 294.890 385.280 305.070 385.450 ;
        RECT 294.940 381.260 305.070 385.280 ;
        RECT 305.460 384.060 305.630 385.820 ;
        RECT 294.940 381.180 305.050 381.260 ;
        RECT 294.370 380.880 294.550 380.950 ;
        RECT 305.460 380.880 306.070 384.060 ;
        RECT 294.370 380.710 306.070 380.880 ;
        RECT 305.530 380.600 306.070 380.710 ;
        RECT 306.530 380.360 307.080 386.710 ;
        RECT 306.520 380.200 307.080 380.360 ;
        RECT 279.700 379.860 307.080 380.200 ;
        RECT 308.290 386.710 335.670 387.220 ;
        RECT 308.290 384.780 309.090 386.710 ;
        RECT 309.670 386.260 309.840 386.340 ;
        RECT 320.910 386.260 321.140 386.350 ;
        RECT 309.670 386.250 321.140 386.260 ;
        RECT 308.290 380.200 308.800 384.780 ;
        RECT 309.660 380.780 321.140 386.250 ;
        RECT 309.590 380.610 321.140 380.780 ;
        RECT 309.660 380.550 309.850 380.610 ;
        RECT 320.910 380.370 321.140 380.610 ;
        RECT 309.540 380.200 311.340 380.210 ;
        RECT 321.700 380.200 322.210 386.710 ;
        RECT 322.970 385.820 334.220 385.990 ;
        RECT 322.970 380.950 323.140 385.820 ;
        RECT 323.530 385.490 333.640 385.510 ;
        RECT 323.530 385.450 333.660 385.490 ;
        RECT 323.480 385.280 333.660 385.450 ;
        RECT 323.530 381.260 333.660 385.280 ;
        RECT 334.050 384.060 334.220 385.820 ;
        RECT 323.530 381.180 333.640 381.260 ;
        RECT 322.960 380.880 323.140 380.950 ;
        RECT 334.050 380.880 334.660 384.060 ;
        RECT 322.960 380.710 334.660 380.880 ;
        RECT 334.120 380.600 334.660 380.710 ;
        RECT 335.120 380.360 335.670 386.710 ;
        RECT 335.110 380.200 335.670 380.360 ;
        RECT 308.290 379.860 335.670 380.200 ;
        RECT 336.880 386.710 364.260 387.220 ;
        RECT 336.880 384.780 337.680 386.710 ;
        RECT 338.260 386.260 338.430 386.340 ;
        RECT 349.500 386.260 349.730 386.350 ;
        RECT 338.260 386.250 349.730 386.260 ;
        RECT 336.880 380.200 337.390 384.780 ;
        RECT 338.250 380.780 349.730 386.250 ;
        RECT 338.180 380.610 349.730 380.780 ;
        RECT 338.250 380.550 338.440 380.610 ;
        RECT 349.500 380.370 349.730 380.610 ;
        RECT 338.130 380.200 339.930 380.210 ;
        RECT 350.290 380.200 350.800 386.710 ;
        RECT 351.560 385.820 362.810 385.990 ;
        RECT 351.560 380.950 351.730 385.820 ;
        RECT 352.120 385.490 362.230 385.510 ;
        RECT 352.120 385.450 362.250 385.490 ;
        RECT 352.070 385.280 362.250 385.450 ;
        RECT 352.120 381.260 362.250 385.280 ;
        RECT 362.640 384.060 362.810 385.820 ;
        RECT 352.120 381.180 362.230 381.260 ;
        RECT 351.550 380.880 351.730 380.950 ;
        RECT 362.640 380.880 363.250 384.060 ;
        RECT 351.550 380.710 363.250 380.880 ;
        RECT 362.710 380.600 363.250 380.710 ;
        RECT 363.710 380.360 364.260 386.710 ;
        RECT 363.700 380.200 364.260 380.360 ;
        RECT 336.880 380.000 364.260 380.200 ;
        RECT 336.880 379.860 371.230 380.000 ;
        RECT 146.970 379.690 147.140 379.720 ;
        RECT 146.880 379.650 147.200 379.690 ;
        RECT 147.650 379.680 147.820 379.720 ;
        RECT 165.370 379.690 192.720 379.860 ;
        RECT 193.960 379.690 221.310 379.860 ;
        RECT 222.550 379.690 249.900 379.860 ;
        RECT 251.140 379.690 278.490 379.860 ;
        RECT 279.730 379.690 307.080 379.860 ;
        RECT 308.320 379.690 335.670 379.860 ;
        RECT 336.910 379.690 371.230 379.860 ;
        RECT 145.520 379.570 146.420 379.610 ;
        RECT 132.060 379.460 132.230 379.480 ;
        RECT 145.510 379.380 146.420 379.570 ;
        RECT 146.870 379.460 147.200 379.650 ;
        RECT 147.570 379.640 147.890 379.680 ;
        RECT 165.370 379.670 166.060 379.690 ;
        RECT 166.570 379.680 168.370 379.690 ;
        RECT 146.880 379.430 147.200 379.460 ;
        RECT 147.560 379.450 147.890 379.640 ;
        RECT 146.970 379.390 147.140 379.430 ;
        RECT 147.570 379.420 147.890 379.450 ;
        RECT 147.650 379.390 147.820 379.420 ;
        RECT 145.520 379.350 146.420 379.380 ;
        RECT 154.750 379.370 154.920 379.390 ;
        RECT 129.740 378.650 129.910 379.320 ;
        RECT 130.120 379.280 130.450 379.320 ;
        RECT 130.130 379.250 130.450 379.280 ;
        RECT 132.120 378.980 132.790 379.150 ;
        RECT 129.250 378.480 129.920 378.650 ;
        RECT 130.650 378.480 131.330 378.650 ;
        RECT 129.740 377.540 129.910 378.480 ;
        RECT 131.630 378.360 131.820 378.420 ;
        RECT 131.630 378.190 132.800 378.360 ;
        RECT 131.560 377.910 131.730 377.940 ;
        RECT 131.560 377.880 131.890 377.910 ;
        RECT 131.560 377.690 131.900 377.880 ;
        RECT 131.560 377.650 131.890 377.690 ;
        RECT 131.560 377.610 131.730 377.650 ;
        RECT 130.310 377.530 130.480 377.590 ;
        RECT 132.130 377.580 132.800 377.750 ;
        RECT 129.250 377.360 129.920 377.530 ;
        RECT 130.310 377.360 131.330 377.530 ;
        RECT 130.310 377.260 130.480 377.360 ;
        RECT 130.110 376.690 130.430 376.710 ;
        RECT 131.540 376.690 131.860 376.730 ;
        RECT 129.240 376.520 132.820 376.690 ;
        RECT 130.100 376.480 130.430 376.520 ;
        RECT 131.530 376.500 131.860 376.520 ;
        RECT 130.110 376.450 130.430 376.480 ;
        RECT 131.540 376.470 131.860 376.500 ;
        RECT 129.320 376.090 129.640 376.130 ;
        RECT 130.250 376.090 130.570 376.130 ;
        RECT 130.950 376.090 131.270 376.130 ;
        RECT 131.690 376.090 132.010 376.130 ;
        RECT 129.310 376.020 129.640 376.090 ;
        RECT 130.240 376.020 130.570 376.090 ;
        RECT 130.940 376.020 131.270 376.090 ;
        RECT 131.680 376.070 132.010 376.090 ;
        RECT 132.400 376.080 132.720 376.120 ;
        RECT 132.390 376.070 132.720 376.080 ;
        RECT 131.680 376.020 132.720 376.070 ;
        RECT 129.290 375.850 132.720 376.020 ;
        RECT 134.390 375.910 134.560 376.580 ;
        RECT 144.880 376.490 145.050 379.140 ;
        RECT 146.250 378.950 146.420 379.350 ;
        RECT 151.860 379.200 154.920 379.370 ;
        RECT 154.750 378.550 154.920 379.200 ;
        RECT 146.140 377.470 149.450 378.450 ;
        RECT 154.750 378.380 156.020 378.550 ;
        RECT 153.540 377.460 153.770 378.150 ;
        RECT 144.880 375.950 145.060 376.490 ;
        RECT 144.800 375.910 145.120 375.950 ;
        RECT 146.140 375.920 149.450 376.900 ;
        RECT 153.540 376.450 153.770 377.140 ;
        RECT 154.750 375.970 154.920 378.380 ;
        RECT 184.310 378.060 184.480 379.690 ;
        RECT 193.960 379.670 194.650 379.690 ;
        RECT 195.160 379.680 196.960 379.690 ;
        RECT 222.550 379.670 223.240 379.690 ;
        RECT 223.750 379.680 225.550 379.690 ;
        RECT 251.140 379.670 251.830 379.690 ;
        RECT 252.340 379.680 254.140 379.690 ;
        RECT 279.730 379.670 280.420 379.690 ;
        RECT 280.930 379.680 282.730 379.690 ;
        RECT 308.320 379.670 309.010 379.690 ;
        RECT 309.520 379.680 311.320 379.690 ;
        RECT 336.910 379.670 337.600 379.690 ;
        RECT 338.110 379.680 339.910 379.690 ;
        RECT 363.700 379.450 371.230 379.690 ;
        RECT 363.700 379.440 364.370 379.450 ;
        RECT 157.490 377.370 157.660 377.620 ;
        RECT 156.180 377.200 158.390 377.370 ;
        RECT 157.490 376.730 157.660 377.200 ;
        RECT 154.660 375.930 154.980 375.970 ;
        RECT 131.870 375.840 132.720 375.850 ;
        RECT 144.790 375.720 145.120 375.910 ;
        RECT 154.650 375.740 154.980 375.930 ;
        RECT 144.800 375.690 145.120 375.720 ;
        RECT 154.660 375.710 154.980 375.740 ;
        RECT 144.830 372.130 146.350 372.140 ;
        RECT 144.830 371.340 146.380 372.130 ;
        RECT 165.520 370.340 165.870 370.440 ;
        RECT 168.590 370.420 170.820 370.570 ;
        RECT 168.590 370.400 170.970 370.420 ;
        RECT 168.590 370.390 168.770 370.400 ;
        RECT 168.130 370.370 168.770 370.390 ;
        RECT 167.180 370.340 167.640 370.370 ;
        RECT 164.110 370.170 164.870 370.340 ;
        RECT 165.120 370.170 166.290 370.340 ;
        RECT 166.530 370.200 167.640 370.340 ;
        RECT 168.090 370.200 168.770 370.370 ;
        RECT 170.370 370.250 170.970 370.400 ;
        RECT 171.430 370.240 171.760 370.410 ;
        RECT 166.530 370.170 167.350 370.200 ;
        RECT 164.110 370.160 164.340 370.170 ;
        RECT 164.070 369.720 164.340 370.160 ;
        RECT 167.090 370.030 167.350 370.170 ;
        RECT 168.590 370.140 168.770 370.200 ;
        RECT 169.710 370.050 170.040 370.220 ;
        RECT 165.550 369.720 165.880 369.980 ;
        RECT 167.090 369.860 168.270 370.030 ;
        RECT 167.090 369.720 167.350 369.860 ;
        RECT 163.520 369.580 163.690 369.640 ;
        RECT 163.490 369.360 163.710 369.580 ;
        RECT 164.040 369.540 164.370 369.720 ;
        RECT 164.620 369.550 166.780 369.720 ;
        RECT 167.020 369.550 167.350 369.720 ;
        RECT 167.180 369.500 167.350 369.550 ;
        RECT 167.640 369.360 167.850 369.690 ;
        RECT 168.090 369.420 168.270 369.860 ;
        RECT 169.790 369.800 170.040 370.050 ;
        RECT 169.790 369.700 170.260 369.800 ;
        RECT 171.510 369.780 171.690 370.240 ;
        RECT 169.620 369.690 170.260 369.700 ;
        RECT 168.820 369.630 170.260 369.690 ;
        RECT 168.820 369.520 170.180 369.630 ;
        RECT 170.730 369.610 171.690 369.780 ;
        RECT 163.520 369.310 163.690 369.360 ;
        RECT 165.520 368.790 165.870 368.890 ;
        RECT 168.590 368.870 170.820 369.020 ;
        RECT 168.590 368.850 170.970 368.870 ;
        RECT 168.590 368.840 168.770 368.850 ;
        RECT 168.130 368.820 168.770 368.840 ;
        RECT 167.180 368.790 167.640 368.820 ;
        RECT 164.110 368.620 164.870 368.790 ;
        RECT 165.120 368.620 166.290 368.790 ;
        RECT 166.530 368.650 167.640 368.790 ;
        RECT 168.090 368.650 168.770 368.820 ;
        RECT 170.370 368.700 170.970 368.850 ;
        RECT 171.430 368.690 171.760 368.860 ;
        RECT 166.530 368.620 167.350 368.650 ;
        RECT 164.110 368.610 164.340 368.620 ;
        RECT 141.130 368.210 141.330 368.250 ;
        RECT 140.820 367.950 141.330 368.210 ;
        RECT 141.130 367.920 141.330 367.950 ;
        RECT 141.720 368.220 141.920 368.250 ;
        RECT 141.720 368.180 142.230 368.220 ;
        RECT 141.720 367.990 142.240 368.180 ;
        RECT 164.070 368.170 164.340 368.610 ;
        RECT 167.090 368.480 167.350 368.620 ;
        RECT 168.590 368.590 168.770 368.650 ;
        RECT 169.710 368.500 170.040 368.670 ;
        RECT 165.550 368.170 165.880 368.430 ;
        RECT 167.090 368.310 168.270 368.480 ;
        RECT 167.090 368.170 167.350 368.310 ;
        RECT 163.520 368.030 163.690 368.090 ;
        RECT 141.720 367.960 142.230 367.990 ;
        RECT 141.720 367.920 141.920 367.960 ;
        RECT 142.410 367.770 142.580 367.820 ;
        RECT 163.490 367.810 163.710 368.030 ;
        RECT 164.040 367.990 164.370 368.170 ;
        RECT 164.620 368.000 166.780 368.170 ;
        RECT 167.020 368.000 167.350 368.170 ;
        RECT 167.180 367.950 167.350 368.000 ;
        RECT 167.640 367.810 167.850 368.140 ;
        RECT 168.090 367.870 168.270 368.310 ;
        RECT 169.790 368.250 170.040 368.500 ;
        RECT 169.790 368.150 170.260 368.250 ;
        RECT 171.510 368.230 171.690 368.690 ;
        RECT 169.620 368.140 170.260 368.150 ;
        RECT 168.820 368.080 170.260 368.140 ;
        RECT 168.820 367.970 170.180 368.080 ;
        RECT 170.730 368.060 171.690 368.230 ;
        RECT 192.800 368.180 193.470 369.050 ;
        RECT 205.080 368.740 207.180 369.050 ;
        RECT 205.080 368.570 207.600 368.740 ;
        RECT 207.840 368.720 208.030 368.750 ;
        RECT 205.080 368.200 207.180 368.570 ;
        RECT 207.840 368.550 208.900 368.720 ;
        RECT 233.660 368.570 234.190 368.740 ;
        RECT 207.840 368.520 208.030 368.550 ;
        RECT 205.580 367.860 205.800 368.200 ;
        RECT 205.580 367.850 205.790 367.860 ;
        RECT 140.380 367.750 140.810 367.770 ;
        RECT 140.380 367.580 140.830 367.750 ;
        RECT 142.400 367.740 142.580 367.770 ;
        RECT 163.520 367.760 163.690 367.810 ;
        RECT 142.400 367.730 142.830 367.740 ;
        RECT 140.380 367.560 140.810 367.580 ;
        RECT 142.400 367.500 142.990 367.730 ;
        RECT 205.960 367.680 206.150 367.690 ;
        RECT 142.400 367.490 142.830 367.500 ;
        RECT 142.400 367.430 142.570 367.490 ;
        RECT 141.130 367.290 141.330 367.330 ;
        RECT 2.180 366.750 9.710 367.260 ;
        RECT 140.820 367.030 141.330 367.290 ;
        RECT 141.130 367.000 141.330 367.030 ;
        RECT 141.720 367.300 141.920 367.330 ;
        RECT 141.720 367.260 142.230 367.300 ;
        RECT 141.720 367.070 142.240 367.260 ;
        RECT 165.520 367.240 165.870 367.340 ;
        RECT 168.590 367.320 170.820 367.470 ;
        RECT 205.950 367.390 206.150 367.680 ;
        RECT 168.590 367.300 170.970 367.320 ;
        RECT 168.590 367.290 168.770 367.300 ;
        RECT 168.130 367.270 168.770 367.290 ;
        RECT 167.180 367.240 167.640 367.270 ;
        RECT 164.110 367.070 164.870 367.240 ;
        RECT 165.120 367.070 166.290 367.240 ;
        RECT 166.530 367.100 167.640 367.240 ;
        RECT 168.090 367.100 168.770 367.270 ;
        RECT 170.370 367.150 170.970 367.300 ;
        RECT 171.430 367.140 171.760 367.310 ;
        RECT 166.530 367.070 167.350 367.100 ;
        RECT 141.720 367.040 142.230 367.070 ;
        RECT 164.110 367.060 164.340 367.070 ;
        RECT 141.720 367.000 141.920 367.040 ;
        RECT 0.480 360.730 1.940 360.770 ;
        RECT 0.480 360.560 1.950 360.730 ;
        RECT 0.480 360.520 1.940 360.560 ;
        RECT 2.180 354.140 2.690 366.750 ;
        RECT 3.050 365.960 9.030 366.190 ;
        RECT 3.140 354.900 8.790 365.960 ;
        RECT 9.200 356.390 9.710 366.750 ;
        RECT 140.380 366.830 140.810 366.850 ;
        RECT 140.380 366.660 140.830 366.830 ;
        RECT 140.380 366.640 140.810 366.660 ;
        RECT 164.070 366.620 164.340 367.060 ;
        RECT 167.090 366.930 167.350 367.070 ;
        RECT 168.590 367.040 168.770 367.100 ;
        RECT 169.710 366.950 170.040 367.120 ;
        RECT 165.550 366.620 165.880 366.880 ;
        RECT 167.090 366.760 168.270 366.930 ;
        RECT 167.090 366.620 167.350 366.760 ;
        RECT 163.520 366.480 163.690 366.540 ;
        RECT 141.130 366.370 141.330 366.410 ;
        RECT 140.820 366.110 141.330 366.370 ;
        RECT 141.130 366.080 141.330 366.110 ;
        RECT 141.720 366.380 141.920 366.410 ;
        RECT 141.720 366.340 142.230 366.380 ;
        RECT 141.720 366.150 142.240 366.340 ;
        RECT 163.490 366.260 163.710 366.480 ;
        RECT 164.040 366.440 164.370 366.620 ;
        RECT 164.620 366.450 166.780 366.620 ;
        RECT 167.020 366.450 167.350 366.620 ;
        RECT 167.180 366.400 167.350 366.450 ;
        RECT 167.640 366.260 167.850 366.590 ;
        RECT 168.090 366.320 168.270 366.760 ;
        RECT 169.790 366.700 170.040 366.950 ;
        RECT 169.790 366.600 170.260 366.700 ;
        RECT 171.510 366.680 171.690 367.140 ;
        RECT 205.920 367.060 206.160 367.390 ;
        RECT 169.620 366.590 170.260 366.600 ;
        RECT 168.820 366.530 170.260 366.590 ;
        RECT 168.820 366.420 170.180 366.530 ;
        RECT 170.730 366.510 171.690 366.680 ;
        RECT 206.350 366.580 206.520 368.190 ;
        RECT 207.180 367.090 207.350 368.180 ;
        RECT 208.310 368.160 208.500 368.190 ;
        RECT 207.770 367.990 208.500 368.160 ;
        RECT 208.730 368.160 208.900 368.550 ;
        RECT 235.470 368.470 235.670 368.820 ;
        RECT 235.470 368.440 235.680 368.470 ;
        RECT 208.730 367.990 209.470 368.160 ;
        RECT 231.790 367.990 232.140 368.160 ;
        RECT 233.160 367.990 233.490 368.160 ;
        RECT 208.310 367.960 208.500 367.990 ;
        RECT 210.530 367.370 210.760 367.890 ;
        RECT 207.770 367.200 210.760 367.370 ;
        RECT 206.950 367.050 207.350 367.090 ;
        RECT 206.940 366.860 207.350 367.050 ;
        RECT 215.730 367.010 216.280 367.440 ;
        RECT 224.980 367.010 225.530 367.440 ;
        RECT 228.610 367.200 228.840 367.890 ;
        RECT 233.910 367.660 234.080 368.180 ;
        RECT 233.750 367.400 234.080 367.660 ;
        RECT 231.790 367.200 232.140 367.370 ;
        RECT 233.160 367.200 233.490 367.370 ;
        RECT 206.950 366.830 207.350 366.860 ;
        RECT 206.340 366.390 206.520 366.580 ;
        RECT 207.180 366.490 207.350 366.830 ;
        RECT 207.840 366.580 208.030 366.760 ;
        RECT 207.770 366.410 208.120 366.580 ;
        RECT 163.520 366.210 163.690 366.260 ;
        RECT 141.720 366.120 142.230 366.150 ;
        RECT 141.720 366.080 141.920 366.120 ;
        RECT 208.690 366.000 208.900 366.430 ;
        RECT 209.120 366.410 209.460 366.580 ;
        RECT 208.710 365.980 208.880 366.000 ;
        RECT 140.380 365.910 140.810 365.930 ;
        RECT 140.380 365.740 140.830 365.910 ;
        RECT 140.380 365.720 140.810 365.740 ;
        RECT 165.520 365.690 165.870 365.790 ;
        RECT 168.590 365.770 170.820 365.920 ;
        RECT 168.590 365.750 170.970 365.770 ;
        RECT 168.590 365.740 168.770 365.750 ;
        RECT 168.130 365.720 168.770 365.740 ;
        RECT 167.180 365.690 167.640 365.720 ;
        RECT 164.110 365.520 164.870 365.690 ;
        RECT 165.120 365.520 166.290 365.690 ;
        RECT 166.530 365.550 167.640 365.690 ;
        RECT 168.090 365.550 168.770 365.720 ;
        RECT 170.370 365.600 170.970 365.750 ;
        RECT 171.430 365.590 171.760 365.760 ;
        RECT 206.340 365.670 206.520 365.860 ;
        RECT 166.530 365.520 167.350 365.550 ;
        RECT 164.110 365.510 164.340 365.520 ;
        RECT 140.630 365.350 140.950 365.390 ;
        RECT 140.630 365.330 140.960 365.350 ;
        RECT 140.630 365.130 141.250 365.330 ;
        RECT 141.080 365.000 141.250 365.130 ;
        RECT 141.760 365.290 141.930 365.330 ;
        RECT 141.760 365.250 142.250 365.290 ;
        RECT 141.760 365.060 142.260 365.250 ;
        RECT 164.070 365.070 164.340 365.510 ;
        RECT 167.090 365.380 167.350 365.520 ;
        RECT 168.590 365.490 168.770 365.550 ;
        RECT 169.710 365.400 170.040 365.570 ;
        RECT 165.550 365.070 165.880 365.330 ;
        RECT 167.090 365.210 168.270 365.380 ;
        RECT 167.090 365.070 167.350 365.210 ;
        RECT 141.760 365.030 142.250 365.060 ;
        RECT 141.760 365.000 141.930 365.030 ;
        RECT 163.520 364.930 163.690 364.990 ;
        RECT 140.470 364.890 140.900 364.910 ;
        RECT 140.450 364.720 140.900 364.890 ;
        RECT 140.470 364.700 140.900 364.720 ;
        RECT 163.490 364.710 163.710 364.930 ;
        RECT 164.040 364.890 164.370 365.070 ;
        RECT 164.620 364.900 166.780 365.070 ;
        RECT 167.020 364.900 167.350 365.070 ;
        RECT 167.180 364.850 167.350 364.900 ;
        RECT 167.640 364.710 167.850 365.040 ;
        RECT 168.090 364.770 168.270 365.210 ;
        RECT 169.790 365.150 170.040 365.400 ;
        RECT 169.790 365.050 170.260 365.150 ;
        RECT 171.510 365.130 171.690 365.590 ;
        RECT 169.620 365.040 170.260 365.050 ;
        RECT 168.820 364.980 170.260 365.040 ;
        RECT 168.820 364.870 170.180 364.980 ;
        RECT 170.730 364.960 171.690 365.130 ;
        RECT 205.920 364.860 206.160 365.190 ;
        RECT 163.520 364.660 163.690 364.710 ;
        RECT 205.950 364.570 206.150 364.860 ;
        RECT 205.960 364.560 206.150 364.570 ;
        RECT 140.630 364.390 140.950 364.430 ;
        RECT 205.580 364.390 205.790 364.400 ;
        RECT 140.630 364.370 140.960 364.390 ;
        RECT 140.630 364.170 141.250 364.370 ;
        RECT 141.080 364.040 141.250 364.170 ;
        RECT 141.760 364.330 141.930 364.370 ;
        RECT 141.760 364.290 142.250 364.330 ;
        RECT 141.760 364.100 142.260 364.290 ;
        RECT 141.760 364.070 142.250 364.100 ;
        RECT 141.760 364.040 141.930 364.070 ;
        RECT 140.470 363.930 140.900 363.950 ;
        RECT 140.450 363.760 140.900 363.930 ;
        RECT 205.580 363.810 205.800 364.390 ;
        RECT 206.350 364.060 206.520 365.670 ;
        RECT 207.180 365.400 207.350 365.760 ;
        RECT 207.770 365.670 208.120 365.840 ;
        RECT 208.310 365.820 208.500 365.870 ;
        RECT 209.210 365.840 209.380 366.410 ;
        RECT 213.490 366.180 213.680 366.580 ;
        RECT 227.580 366.180 227.770 366.580 ;
        RECT 231.800 366.410 232.140 366.580 ;
        RECT 233.160 366.410 233.490 366.580 ;
        RECT 233.910 366.490 234.080 367.400 ;
        RECT 234.740 366.580 234.910 368.190 ;
        RECT 235.460 367.860 235.680 368.440 ;
        RECT 235.470 367.850 235.680 367.860 ;
        RECT 235.110 367.680 235.300 367.690 ;
        RECT 235.110 367.390 235.310 367.680 ;
        RECT 235.100 367.060 235.340 367.390 ;
        RECT 213.490 366.170 213.870 366.180 ;
        RECT 210.130 365.990 213.870 366.170 ;
        RECT 213.490 365.950 213.870 365.990 ;
        RECT 227.390 366.170 227.770 366.180 ;
        RECT 227.390 365.990 231.130 366.170 ;
        RECT 227.390 365.950 227.770 365.990 ;
        RECT 208.310 365.810 208.540 365.820 ;
        RECT 209.120 365.810 209.460 365.840 ;
        RECT 208.310 365.670 209.460 365.810 ;
        RECT 207.850 365.460 208.040 365.670 ;
        RECT 208.310 365.640 209.290 365.670 ;
        RECT 208.450 365.610 209.290 365.640 ;
        RECT 213.490 365.570 213.680 365.950 ;
        RECT 206.940 365.360 207.350 365.400 ;
        RECT 206.930 365.170 207.350 365.360 ;
        RECT 215.730 365.280 216.280 365.710 ;
        RECT 224.980 365.280 225.530 365.710 ;
        RECT 227.580 365.570 227.770 365.950 ;
        RECT 233.240 365.840 233.410 366.410 ;
        RECT 234.740 366.390 234.920 366.580 ;
        RECT 363.700 366.540 364.210 379.440 ;
        RECT 364.610 378.550 368.070 378.990 ;
        RECT 364.610 378.450 370.000 378.550 ;
        RECT 364.720 378.380 370.000 378.450 ;
        RECT 364.720 367.470 364.890 378.380 ;
        RECT 365.270 377.970 369.500 377.990 ;
        RECT 365.190 367.860 369.520 377.970 ;
        RECT 369.290 367.810 369.460 367.860 ;
        RECT 369.830 367.470 370.000 378.380 ;
        RECT 364.720 367.300 370.000 367.470 ;
        RECT 364.720 367.290 364.960 367.300 ;
        RECT 370.720 366.540 371.230 379.450 ;
        RECT 363.700 366.030 371.230 366.540 ;
        RECT 371.440 366.480 372.910 366.730 ;
        RECT 231.800 365.670 232.140 365.840 ;
        RECT 233.160 365.670 233.490 365.840 ;
        RECT 232.280 365.270 232.600 365.300 ;
        RECT 233.090 365.280 233.260 365.330 ;
        RECT 233.910 365.300 234.080 365.760 ;
        RECT 234.740 365.670 234.920 365.860 ;
        RECT 206.940 365.140 207.350 365.170 ;
        RECT 207.180 364.070 207.350 365.140 ;
        RECT 207.770 364.950 210.700 365.050 ;
        RECT 207.770 364.880 210.760 364.950 ;
        RECT 209.790 364.560 209.960 364.620 ;
        RECT 209.770 364.350 209.980 364.560 ;
        RECT 208.300 364.260 208.490 364.290 ;
        RECT 209.790 364.280 209.960 364.350 ;
        RECT 210.530 364.260 210.760 364.880 ;
        RECT 228.610 364.260 228.840 364.990 ;
        RECT 231.060 364.930 231.230 365.210 ;
        RECT 232.280 365.080 232.610 365.270 ;
        RECT 233.090 365.130 233.650 365.280 ;
        RECT 231.060 364.890 231.270 364.930 ;
        RECT 231.060 364.870 231.290 364.890 ;
        RECT 231.790 364.880 232.140 365.050 ;
        RECT 232.280 365.040 232.600 365.080 ;
        RECT 232.410 364.880 232.580 365.040 ;
        RECT 233.020 365.020 233.650 365.130 ;
        RECT 233.850 365.270 234.170 365.300 ;
        RECT 233.850 365.080 234.180 365.270 ;
        RECT 234.420 365.130 234.610 365.160 ;
        RECT 234.740 365.130 234.910 365.670 ;
        RECT 235.140 365.190 235.310 365.220 ;
        RECT 233.850 365.040 234.170 365.080 ;
        RECT 233.020 364.960 233.490 365.020 ;
        RECT 233.160 364.880 233.490 364.960 ;
        RECT 233.910 364.900 234.080 365.040 ;
        RECT 234.420 365.000 234.910 365.130 ;
        RECT 231.060 364.850 231.320 364.870 ;
        RECT 231.060 364.800 231.400 364.850 ;
        RECT 231.060 364.740 231.550 364.800 ;
        RECT 231.060 364.710 231.570 364.740 ;
        RECT 231.100 364.680 231.570 364.710 ;
        RECT 231.230 364.630 231.570 364.680 ;
        RECT 231.350 364.620 231.570 364.630 ;
        RECT 231.360 364.590 231.570 364.620 ;
        RECT 231.380 364.510 231.570 364.590 ;
        RECT 232.510 364.510 232.690 364.850 ;
        RECT 232.740 364.510 233.070 364.630 ;
        RECT 233.240 364.590 233.570 364.760 ;
        RECT 233.750 364.640 234.080 364.900 ;
        RECT 234.330 364.740 234.910 365.000 ;
        RECT 235.100 365.040 235.340 365.190 ;
        RECT 235.100 364.860 235.700 365.040 ;
        RECT 234.560 364.710 234.910 364.740 ;
        RECT 233.320 364.510 233.570 364.590 ;
        RECT 233.910 364.510 234.080 364.640 ;
        RECT 234.740 364.540 234.910 364.710 ;
        RECT 235.110 364.560 235.700 364.860 ;
        RECT 236.520 364.920 237.100 365.090 ;
        RECT 236.520 364.820 236.910 364.920 ;
        RECT 236.520 364.790 236.900 364.820 ;
        RECT 236.520 364.640 236.880 364.790 ;
        RECT 235.140 364.540 235.700 364.560 ;
        RECT 230.890 364.460 231.060 364.480 ;
        RECT 207.770 364.090 208.490 364.260 ;
        RECT 208.300 364.060 208.490 364.090 ;
        RECT 208.660 364.090 209.470 364.260 ;
        RECT 205.580 363.780 205.790 363.810 ;
        RECT 140.470 363.740 140.900 363.760 ;
        RECT 140.630 363.430 140.950 363.470 ;
        RECT 205.590 363.430 205.790 363.780 ;
        RECT 207.870 363.750 208.060 363.780 ;
        RECT 208.660 363.750 208.850 364.090 ;
        RECT 230.870 364.030 231.080 364.460 ;
        RECT 231.380 364.340 231.900 364.510 ;
        RECT 232.250 364.390 234.150 364.510 ;
        RECT 234.740 364.500 235.700 364.540 ;
        RECT 232.250 364.350 234.320 364.390 ;
        RECT 234.530 364.350 235.700 364.500 ;
        RECT 236.170 364.470 236.880 364.640 ;
        RECT 232.250 364.340 235.700 364.350 ;
        RECT 231.380 364.310 231.570 364.340 ;
        RECT 232.250 364.330 235.070 364.340 ;
        RECT 231.790 364.090 232.140 364.260 ;
        RECT 232.510 363.920 232.690 364.330 ;
        RECT 233.320 364.260 233.800 364.330 ;
        RECT 233.160 364.190 233.800 364.260 ;
        RECT 233.160 364.090 233.490 364.190 ;
        RECT 232.390 363.890 232.710 363.920 ;
        RECT 207.070 363.510 207.600 363.680 ;
        RECT 207.870 363.570 208.850 363.750 ;
        RECT 207.870 363.550 208.060 363.570 ;
        RECT 140.630 363.410 140.960 363.430 ;
        RECT 140.630 363.210 141.250 363.410 ;
        RECT 141.080 363.080 141.250 363.210 ;
        RECT 141.760 363.370 141.930 363.410 ;
        RECT 230.870 363.390 231.080 363.820 ;
        RECT 232.390 363.700 232.720 363.890 ;
        RECT 232.390 363.660 232.710 363.700 ;
        RECT 231.380 363.510 231.570 363.540 ;
        RECT 232.510 363.520 232.690 363.660 ;
        RECT 233.320 363.520 233.490 364.090 ;
        RECT 233.910 364.070 234.080 364.330 ;
        RECT 234.150 364.310 235.070 364.330 ;
        RECT 234.150 364.090 234.910 364.310 ;
        RECT 234.150 364.060 234.320 364.090 ;
        RECT 234.560 364.060 234.910 364.090 ;
        RECT 234.560 364.050 234.760 364.060 ;
        RECT 235.150 364.050 235.700 364.340 ;
        RECT 235.460 363.810 235.680 364.050 ;
        RECT 235.470 363.780 235.680 363.810 ;
        RECT 233.660 363.550 234.190 363.680 ;
        RECT 235.470 363.560 235.670 363.780 ;
        RECT 236.170 363.720 236.870 364.030 ;
        RECT 233.660 363.520 234.320 363.550 ;
        RECT 234.560 363.520 234.760 363.560 ;
        RECT 234.880 363.520 235.070 363.540 ;
        RECT 232.250 363.510 235.070 363.520 ;
        RECT 235.150 363.510 235.700 363.560 ;
        RECT 230.890 363.370 231.060 363.390 ;
        RECT 141.760 363.330 142.250 363.370 ;
        RECT 231.380 363.340 231.900 363.510 ;
        RECT 232.250 363.350 235.700 363.510 ;
        RECT 236.020 363.490 236.870 363.720 ;
        RECT 232.250 363.340 234.760 363.350 ;
        RECT 141.760 363.140 142.260 363.330 ;
        RECT 231.380 363.260 231.570 363.340 ;
        RECT 231.360 363.230 231.570 363.260 ;
        RECT 231.350 363.220 231.570 363.230 ;
        RECT 231.230 363.170 231.570 363.220 ;
        RECT 231.100 363.140 231.570 363.170 ;
        RECT 141.760 363.110 142.250 363.140 ;
        RECT 231.060 363.110 231.570 363.140 ;
        RECT 141.760 363.080 141.930 363.110 ;
        RECT 140.470 362.970 140.900 362.990 ;
        RECT 140.450 362.800 140.900 362.970 ;
        RECT 140.470 362.780 140.900 362.800 ;
        RECT 142.260 362.740 142.680 362.910 ;
        RECT 142.360 362.700 142.590 362.740 ;
        RECT 183.480 362.670 183.650 363.090 ;
        RECT 184.290 362.970 184.530 363.000 ;
        RECT 183.960 362.800 184.530 362.970 ;
        RECT 184.770 362.800 186.110 362.970 ;
        RECT 186.560 362.800 187.520 362.970 ;
        RECT 184.290 362.760 184.530 362.800 ;
        RECT 187.070 362.790 187.240 362.800 ;
        RECT 183.410 362.450 183.580 362.490 ;
        RECT 163.520 362.310 163.690 362.360 ;
        RECT 163.490 362.090 163.710 362.310 ;
        RECT 163.520 362.030 163.690 362.090 ;
        RECT 164.040 361.950 164.370 362.130 ;
        RECT 167.180 362.120 167.350 362.170 ;
        RECT 164.620 361.950 166.780 362.120 ;
        RECT 167.020 361.950 167.350 362.120 ;
        RECT 167.640 361.980 167.850 362.310 ;
        RECT 183.350 362.280 183.580 362.450 ;
        RECT 164.070 361.510 164.340 361.950 ;
        RECT 165.550 361.690 165.880 361.950 ;
        RECT 167.090 361.810 167.350 361.950 ;
        RECT 168.090 361.810 168.270 362.250 ;
        RECT 168.820 362.040 170.180 362.150 ;
        RECT 168.820 361.980 170.260 362.040 ;
        RECT 169.620 361.970 170.260 361.980 ;
        RECT 164.110 361.500 164.340 361.510 ;
        RECT 167.090 361.640 168.270 361.810 ;
        RECT 169.790 361.870 170.260 361.970 ;
        RECT 170.730 361.890 171.690 362.060 ;
        RECT 183.410 361.930 183.580 362.280 ;
        RECT 183.750 362.350 183.940 362.370 ;
        RECT 186.750 362.350 187.080 362.530 ;
        RECT 183.750 362.180 184.310 362.350 ;
        RECT 184.770 362.180 187.520 362.350 ;
        RECT 183.750 362.140 183.940 362.180 ;
        RECT 188.050 362.110 188.220 363.040 ;
        RECT 188.450 362.240 188.620 363.090 ;
        RECT 231.060 363.050 231.550 363.110 ;
        RECT 231.060 363.000 231.400 363.050 ;
        RECT 231.060 362.980 231.320 363.000 ;
        RECT 231.060 362.960 231.290 362.980 ;
        RECT 232.510 362.970 232.690 363.340 ;
        RECT 232.740 363.220 233.070 363.340 ;
        RECT 205.590 362.440 205.790 362.790 ;
        RECT 207.070 362.540 207.600 362.710 ;
        RECT 205.580 362.410 205.790 362.440 ;
        RECT 167.090 361.500 167.350 361.640 ;
        RECT 169.790 361.620 170.040 361.870 ;
        RECT 164.110 361.330 164.870 361.500 ;
        RECT 165.120 361.330 166.290 361.500 ;
        RECT 166.530 361.470 167.350 361.500 ;
        RECT 168.590 361.470 168.770 361.530 ;
        RECT 166.530 361.330 167.640 361.470 ;
        RECT 165.520 361.230 165.870 361.330 ;
        RECT 167.180 361.300 167.640 361.330 ;
        RECT 168.090 361.300 168.770 361.470 ;
        RECT 169.710 361.450 170.040 361.620 ;
        RECT 171.510 361.430 171.690 361.890 ;
        RECT 205.580 361.830 205.800 362.410 ;
        RECT 205.580 361.820 205.790 361.830 ;
        RECT 168.130 361.280 168.770 361.300 ;
        RECT 168.590 361.270 168.770 361.280 ;
        RECT 170.370 361.270 170.970 361.420 ;
        RECT 168.590 361.250 170.970 361.270 ;
        RECT 171.430 361.260 171.760 361.430 ;
        RECT 183.410 361.340 183.580 361.690 ;
        RECT 205.960 361.650 206.150 361.660 ;
        RECT 168.590 361.100 170.820 361.250 ;
        RECT 183.350 361.170 183.580 361.340 ;
        RECT 183.750 361.440 183.940 361.480 ;
        RECT 183.750 361.270 184.310 361.440 ;
        RECT 184.770 361.270 187.520 361.440 ;
        RECT 183.750 361.250 183.940 361.270 ;
        RECT 183.410 361.130 183.580 361.170 ;
        RECT 186.750 361.090 187.080 361.270 ;
        RECT 163.520 360.760 163.690 360.810 ;
        RECT 163.490 360.540 163.710 360.760 ;
        RECT 163.520 360.480 163.690 360.540 ;
        RECT 164.040 360.400 164.370 360.580 ;
        RECT 167.180 360.570 167.350 360.620 ;
        RECT 164.620 360.400 166.780 360.570 ;
        RECT 167.020 360.400 167.350 360.570 ;
        RECT 167.640 360.430 167.850 360.760 ;
        RECT 164.070 359.960 164.340 360.400 ;
        RECT 165.550 360.140 165.880 360.400 ;
        RECT 167.090 360.260 167.350 360.400 ;
        RECT 168.090 360.260 168.270 360.700 ;
        RECT 168.820 360.490 170.180 360.600 ;
        RECT 183.480 360.530 183.650 360.950 ;
        RECT 184.290 360.820 184.530 360.860 ;
        RECT 187.070 360.820 187.240 360.830 ;
        RECT 183.960 360.650 184.530 360.820 ;
        RECT 184.770 360.650 186.110 360.820 ;
        RECT 186.560 360.650 187.520 360.820 ;
        RECT 184.290 360.620 184.530 360.650 ;
        RECT 188.050 360.580 188.220 361.510 ;
        RECT 188.450 360.530 188.620 361.380 ;
        RECT 205.950 361.360 206.150 361.650 ;
        RECT 205.920 361.030 206.160 361.360 ;
        RECT 206.350 360.550 206.520 362.160 ;
        RECT 168.820 360.430 170.260 360.490 ;
        RECT 169.620 360.420 170.260 360.430 ;
        RECT 164.110 359.950 164.340 359.960 ;
        RECT 167.090 360.090 168.270 360.260 ;
        RECT 169.790 360.320 170.260 360.420 ;
        RECT 170.730 360.340 171.690 360.510 ;
        RECT 206.340 360.360 206.520 360.550 ;
        RECT 207.180 361.630 207.350 362.150 ;
        RECT 207.770 361.960 208.100 362.130 ;
        RECT 209.120 361.960 209.470 362.130 ;
        RECT 209.790 362.110 214.850 362.940 ;
        RECT 231.060 362.920 231.270 362.960 ;
        RECT 231.060 362.640 231.230 362.920 ;
        RECT 232.410 362.810 232.690 362.970 ;
        RECT 233.320 362.930 233.490 363.340 ;
        RECT 234.150 363.260 234.760 363.340 ;
        RECT 234.880 363.310 235.700 363.350 ;
        RECT 234.150 363.220 234.320 363.260 ;
        RECT 234.560 363.230 234.760 363.260 ;
        RECT 233.290 362.900 233.490 362.930 ;
        RECT 233.270 362.890 233.490 362.900 ;
        RECT 232.280 362.550 232.690 362.810 ;
        RECT 233.020 362.810 233.490 362.890 ;
        RECT 233.910 362.810 234.080 362.970 ;
        RECT 234.420 362.900 234.610 362.920 ;
        RECT 234.420 362.890 234.760 362.900 ;
        RECT 234.420 362.870 234.860 362.890 ;
        RECT 233.020 362.720 233.480 362.810 ;
        RECT 233.290 362.700 233.480 362.720 ;
        RECT 233.850 362.770 234.170 362.810 ;
        RECT 233.850 362.710 234.180 362.770 ;
        RECT 234.330 362.720 234.860 362.870 ;
        RECT 232.510 362.280 232.690 362.550 ;
        RECT 233.120 362.610 233.440 362.640 ;
        RECT 233.120 362.420 233.450 362.610 ;
        RECT 233.660 362.540 234.190 362.710 ;
        RECT 234.330 362.610 234.760 362.720 ;
        RECT 235.140 362.630 235.700 363.310 ;
        RECT 236.170 363.150 236.870 363.490 ;
        RECT 236.630 362.790 236.950 362.830 ;
        RECT 236.630 362.730 236.960 362.790 ;
        RECT 234.560 362.570 234.760 362.610 ;
        RECT 235.150 362.570 235.700 362.630 ;
        RECT 236.160 362.600 236.960 362.730 ;
        RECT 236.160 362.570 236.950 362.600 ;
        RECT 235.470 362.440 235.670 362.570 ;
        RECT 236.160 362.550 236.860 362.570 ;
        RECT 233.120 362.380 233.440 362.420 ;
        RECT 235.470 362.410 235.680 362.440 ;
        RECT 233.120 362.300 233.290 362.380 ;
        RECT 214.300 362.030 214.780 362.110 ;
        RECT 207.180 361.370 207.510 361.630 ;
        RECT 207.180 360.460 207.350 361.370 ;
        RECT 207.770 361.170 208.100 361.340 ;
        RECT 209.120 361.170 209.470 361.340 ;
        RECT 212.420 361.170 212.650 361.860 ;
        RECT 214.300 361.780 214.770 362.030 ;
        RECT 231.060 361.910 231.230 362.190 ;
        RECT 231.790 361.960 232.140 362.130 ;
        RECT 232.280 362.020 232.690 362.280 ;
        RECT 233.070 362.130 233.290 362.300 ;
        RECT 233.850 362.250 234.170 362.280 ;
        RECT 233.070 362.110 233.490 362.130 ;
        RECT 231.060 361.870 231.270 361.910 ;
        RECT 215.730 360.980 216.280 361.410 ;
        RECT 224.980 360.980 225.530 361.410 ;
        RECT 228.610 361.170 228.840 361.860 ;
        RECT 231.060 361.850 231.290 361.870 ;
        RECT 232.410 361.860 232.690 362.020 ;
        RECT 233.020 361.960 233.490 362.110 ;
        RECT 233.850 362.060 234.180 362.250 ;
        RECT 234.420 362.110 234.610 362.140 ;
        RECT 234.740 362.110 234.910 362.160 ;
        RECT 233.850 362.020 234.170 362.060 ;
        RECT 234.420 362.040 234.910 362.110 ;
        RECT 233.020 361.940 233.480 361.960 ;
        RECT 233.270 361.930 233.480 361.940 ;
        RECT 233.290 361.900 233.480 361.930 ;
        RECT 231.060 361.830 231.320 361.850 ;
        RECT 231.060 361.780 231.400 361.830 ;
        RECT 231.060 361.720 231.550 361.780 ;
        RECT 231.060 361.690 231.570 361.720 ;
        RECT 231.100 361.660 231.570 361.690 ;
        RECT 231.230 361.610 231.570 361.660 ;
        RECT 231.350 361.600 231.570 361.610 ;
        RECT 231.360 361.570 231.570 361.600 ;
        RECT 231.380 361.490 231.570 361.570 ;
        RECT 232.510 361.490 232.690 361.860 ;
        RECT 233.600 361.710 233.790 361.830 ;
        RECT 233.240 361.630 233.790 361.710 ;
        RECT 233.910 361.630 234.080 362.020 ;
        RECT 234.330 361.780 234.910 362.040 ;
        RECT 234.560 361.750 234.910 361.780 ;
        RECT 232.740 361.490 233.070 361.610 ;
        RECT 233.240 361.540 234.080 361.630 ;
        RECT 233.320 361.490 233.490 361.540 ;
        RECT 233.750 361.490 234.080 361.540 ;
        RECT 234.740 361.520 234.910 361.750 ;
        RECT 235.140 362.080 235.310 362.200 ;
        RECT 235.460 362.080 235.680 362.410 ;
        RECT 235.140 361.660 235.700 362.080 ;
        RECT 236.620 362.070 236.940 362.110 ;
        RECT 236.160 361.890 236.950 362.070 ;
        RECT 236.620 361.880 236.950 361.890 ;
        RECT 236.620 361.850 236.940 361.880 ;
        RECT 235.110 361.520 235.700 361.660 ;
        RECT 230.890 361.440 231.060 361.460 ;
        RECT 230.870 361.010 231.080 361.440 ;
        RECT 231.380 361.340 231.900 361.490 ;
        RECT 232.250 361.430 234.150 361.490 ;
        RECT 234.740 361.480 235.700 361.520 ;
        RECT 232.250 361.390 234.320 361.430 ;
        RECT 234.530 361.390 235.700 361.480 ;
        RECT 231.380 361.320 232.140 361.340 ;
        RECT 231.380 361.290 231.570 361.320 ;
        RECT 231.790 361.170 232.140 361.320 ;
        RECT 232.250 361.320 235.700 361.390 ;
        RECT 232.250 361.310 235.070 361.320 ;
        RECT 207.770 360.380 208.100 360.550 ;
        RECT 209.120 360.380 209.460 360.550 ;
        RECT 167.090 359.950 167.350 360.090 ;
        RECT 169.790 360.070 170.040 360.320 ;
        RECT 164.110 359.780 164.870 359.950 ;
        RECT 165.120 359.780 166.290 359.950 ;
        RECT 166.530 359.920 167.350 359.950 ;
        RECT 168.590 359.920 168.770 359.980 ;
        RECT 166.530 359.780 167.640 359.920 ;
        RECT 165.520 359.680 165.870 359.780 ;
        RECT 167.180 359.750 167.640 359.780 ;
        RECT 168.090 359.750 168.770 359.920 ;
        RECT 169.710 359.900 170.040 360.070 ;
        RECT 171.510 359.880 171.690 360.340 ;
        RECT 168.130 359.730 168.770 359.750 ;
        RECT 168.590 359.720 168.770 359.730 ;
        RECT 170.370 359.720 170.970 359.870 ;
        RECT 168.590 359.700 170.970 359.720 ;
        RECT 171.430 359.710 171.760 359.880 ;
        RECT 183.480 359.740 183.650 360.160 ;
        RECT 184.290 360.040 184.530 360.070 ;
        RECT 183.960 359.870 184.530 360.040 ;
        RECT 184.770 359.870 186.110 360.040 ;
        RECT 186.560 359.870 187.520 360.040 ;
        RECT 184.290 359.830 184.530 359.870 ;
        RECT 187.070 359.860 187.240 359.870 ;
        RECT 168.590 359.550 170.820 359.700 ;
        RECT 183.410 359.520 183.580 359.560 ;
        RECT 183.350 359.350 183.580 359.520 ;
        RECT 163.520 359.210 163.690 359.260 ;
        RECT 163.490 358.990 163.710 359.210 ;
        RECT 163.520 358.930 163.690 358.990 ;
        RECT 164.040 358.850 164.370 359.030 ;
        RECT 167.180 359.020 167.350 359.070 ;
        RECT 164.620 358.850 166.780 359.020 ;
        RECT 167.020 358.850 167.350 359.020 ;
        RECT 167.640 358.880 167.850 359.210 ;
        RECT 164.070 358.410 164.340 358.850 ;
        RECT 165.550 358.590 165.880 358.850 ;
        RECT 167.090 358.710 167.350 358.850 ;
        RECT 168.090 358.710 168.270 359.150 ;
        RECT 168.820 358.940 170.180 359.050 ;
        RECT 183.410 359.000 183.580 359.350 ;
        RECT 183.750 359.420 183.940 359.440 ;
        RECT 186.750 359.420 187.080 359.600 ;
        RECT 183.750 359.250 184.310 359.420 ;
        RECT 184.770 359.250 187.520 359.420 ;
        RECT 183.750 359.210 183.940 359.250 ;
        RECT 188.050 359.180 188.220 360.110 ;
        RECT 188.450 359.310 188.620 360.160 ;
        RECT 206.340 359.640 206.520 359.830 ;
        RECT 207.850 359.810 208.020 360.380 ;
        RECT 213.490 360.150 213.680 360.550 ;
        RECT 227.580 360.150 227.770 360.550 ;
        RECT 230.870 360.370 231.080 360.800 ;
        RECT 231.380 360.490 231.570 360.520 ;
        RECT 231.800 360.490 232.140 360.550 ;
        RECT 232.510 360.500 232.690 361.310 ;
        RECT 233.160 361.170 233.490 361.310 ;
        RECT 233.320 360.550 233.490 361.170 ;
        RECT 233.160 360.500 233.490 360.550 ;
        RECT 233.910 360.500 234.080 361.310 ;
        RECT 234.150 361.290 235.070 361.310 ;
        RECT 234.150 361.130 234.910 361.290 ;
        RECT 234.150 361.100 234.320 361.130 ;
        RECT 234.560 361.090 234.910 361.130 ;
        RECT 234.740 360.600 234.910 361.090 ;
        RECT 235.100 361.090 235.700 361.320 ;
        RECT 236.170 361.130 236.870 361.470 ;
        RECT 235.100 361.030 235.340 361.090 ;
        RECT 236.020 360.900 236.870 361.130 ;
        RECT 234.150 360.560 234.320 360.590 ;
        RECT 234.560 360.560 234.910 360.600 ;
        RECT 234.150 360.550 234.910 360.560 ;
        RECT 234.150 360.520 234.920 360.550 ;
        RECT 234.150 360.500 235.070 360.520 ;
        RECT 231.380 360.380 232.140 360.490 ;
        RECT 232.250 360.490 235.070 360.500 ;
        RECT 235.150 360.490 235.700 360.600 ;
        RECT 236.170 360.590 236.870 360.900 ;
        RECT 230.890 360.350 231.060 360.370 ;
        RECT 231.380 360.320 231.900 360.380 ;
        RECT 232.250 360.330 235.700 360.490 ;
        RECT 232.250 360.320 234.760 360.330 ;
        RECT 231.380 360.240 231.570 360.320 ;
        RECT 231.360 360.210 231.570 360.240 ;
        RECT 231.350 360.200 231.570 360.210 ;
        RECT 231.230 360.150 231.570 360.200 ;
        RECT 213.490 360.140 213.870 360.150 ;
        RECT 210.130 359.960 213.870 360.140 ;
        RECT 213.490 359.920 213.870 359.960 ;
        RECT 227.390 360.140 227.770 360.150 ;
        RECT 231.100 360.140 231.570 360.150 ;
        RECT 227.390 360.090 231.570 360.140 ;
        RECT 227.390 360.030 231.550 360.090 ;
        RECT 227.390 359.980 231.400 360.030 ;
        RECT 227.390 359.960 231.320 359.980 ;
        RECT 227.390 359.920 227.770 359.960 ;
        RECT 168.820 358.880 170.260 358.940 ;
        RECT 169.620 358.870 170.260 358.880 ;
        RECT 164.110 358.400 164.340 358.410 ;
        RECT 167.090 358.540 168.270 358.710 ;
        RECT 169.790 358.770 170.260 358.870 ;
        RECT 170.730 358.790 171.690 358.960 ;
        RECT 205.920 358.830 206.160 359.160 ;
        RECT 167.090 358.400 167.350 358.540 ;
        RECT 169.790 358.520 170.040 358.770 ;
        RECT 164.110 358.230 164.870 358.400 ;
        RECT 165.120 358.230 166.290 358.400 ;
        RECT 166.530 358.370 167.350 358.400 ;
        RECT 168.590 358.370 168.770 358.430 ;
        RECT 166.530 358.230 167.640 358.370 ;
        RECT 165.520 358.130 165.870 358.230 ;
        RECT 167.180 358.200 167.640 358.230 ;
        RECT 168.090 358.200 168.770 358.370 ;
        RECT 169.710 358.350 170.040 358.520 ;
        RECT 171.510 358.330 171.690 358.790 ;
        RECT 183.410 358.410 183.580 358.760 ;
        RECT 168.130 358.180 168.770 358.200 ;
        RECT 168.590 358.170 168.770 358.180 ;
        RECT 170.370 358.170 170.970 358.320 ;
        RECT 168.590 358.150 170.970 358.170 ;
        RECT 171.430 358.160 171.760 358.330 ;
        RECT 183.350 358.240 183.580 358.410 ;
        RECT 183.750 358.510 183.940 358.550 ;
        RECT 183.750 358.340 184.310 358.510 ;
        RECT 184.770 358.340 187.520 358.510 ;
        RECT 183.750 358.320 183.940 358.340 ;
        RECT 183.410 358.200 183.580 358.240 ;
        RECT 186.750 358.160 187.080 358.340 ;
        RECT 168.590 358.000 170.820 358.150 ;
        RECT 163.520 357.660 163.690 357.710 ;
        RECT 163.490 357.440 163.710 357.660 ;
        RECT 163.520 357.380 163.690 357.440 ;
        RECT 164.040 357.300 164.370 357.480 ;
        RECT 167.180 357.470 167.350 357.520 ;
        RECT 164.620 357.300 166.780 357.470 ;
        RECT 167.020 357.300 167.350 357.470 ;
        RECT 167.640 357.330 167.850 357.660 ;
        RECT 183.480 357.600 183.650 358.020 ;
        RECT 184.290 357.890 184.530 357.930 ;
        RECT 187.070 357.890 187.240 357.900 ;
        RECT 183.960 357.720 184.530 357.890 ;
        RECT 184.770 357.720 186.110 357.890 ;
        RECT 186.560 357.720 187.520 357.890 ;
        RECT 184.290 357.690 184.530 357.720 ;
        RECT 188.050 357.650 188.220 358.580 ;
        RECT 205.950 358.540 206.150 358.830 ;
        RECT 205.960 358.530 206.150 358.540 ;
        RECT 188.450 357.600 188.620 358.450 ;
        RECT 205.580 358.360 205.790 358.370 ;
        RECT 205.580 357.780 205.800 358.360 ;
        RECT 206.350 358.030 206.520 359.640 ;
        RECT 207.180 358.870 207.350 359.730 ;
        RECT 207.770 359.640 208.100 359.810 ;
        RECT 209.120 359.640 209.460 359.810 ;
        RECT 213.490 359.540 213.680 359.920 ;
        RECT 215.730 359.250 216.280 359.680 ;
        RECT 224.980 359.250 225.530 359.680 ;
        RECT 227.580 359.540 227.770 359.920 ;
        RECT 231.060 359.940 231.290 359.960 ;
        RECT 232.510 359.950 232.690 360.320 ;
        RECT 232.740 360.200 233.070 360.320 ;
        RECT 231.060 359.900 231.270 359.940 ;
        RECT 231.060 359.620 231.230 359.900 ;
        RECT 231.800 359.640 232.140 359.810 ;
        RECT 232.410 359.790 232.690 359.950 ;
        RECT 233.240 359.870 233.490 360.320 ;
        RECT 234.150 360.300 234.760 360.320 ;
        RECT 234.150 360.260 234.320 360.300 ;
        RECT 234.560 360.270 234.760 360.300 ;
        RECT 234.880 360.290 235.700 360.330 ;
        RECT 232.280 359.750 232.690 359.790 ;
        RECT 232.280 359.560 232.610 359.750 ;
        RECT 233.020 359.700 233.490 359.870 ;
        RECT 233.910 359.790 234.080 359.950 ;
        RECT 234.560 359.910 234.760 359.940 ;
        RECT 234.330 359.870 234.760 359.910 ;
        RECT 234.330 359.830 234.860 359.870 ;
        RECT 233.160 359.640 233.490 359.700 ;
        RECT 233.850 359.750 234.170 359.790 ;
        RECT 233.850 359.560 234.180 359.750 ;
        RECT 234.330 359.650 234.920 359.830 ;
        RECT 234.560 359.640 234.920 359.650 ;
        RECT 234.560 359.610 234.910 359.640 ;
        RECT 235.140 359.610 235.700 360.290 ;
        RECT 236.170 359.980 236.880 360.150 ;
        RECT 236.520 359.700 236.880 359.980 ;
        RECT 232.280 359.530 232.600 359.560 ;
        RECT 233.850 359.530 234.170 359.560 ;
        RECT 233.090 359.250 233.260 359.300 ;
        RECT 207.180 358.610 207.510 358.870 ;
        RECT 207.770 358.850 208.100 359.020 ;
        RECT 209.120 358.850 209.470 359.020 ;
        RECT 207.180 358.040 207.350 358.610 ;
        RECT 212.420 358.230 212.650 358.960 ;
        RECT 207.770 358.060 208.100 358.230 ;
        RECT 209.120 358.060 209.470 358.230 ;
        RECT 214.460 358.100 214.800 358.350 ;
        RECT 228.610 358.230 228.840 358.960 ;
        RECT 231.790 358.850 232.140 359.020 ;
        RECT 233.090 358.990 233.650 359.250 ;
        RECT 233.090 358.970 233.490 358.990 ;
        RECT 233.160 358.850 233.490 358.970 ;
        RECT 233.910 358.870 234.080 359.530 ;
        RECT 234.740 359.010 234.910 359.610 ;
        RECT 236.520 359.530 237.100 359.700 ;
        RECT 234.560 358.970 234.910 359.010 ;
        RECT 214.460 358.020 214.810 358.100 ;
        RECT 231.790 358.060 232.140 358.230 ;
        RECT 205.580 357.750 205.790 357.780 ;
        RECT 164.070 356.860 164.340 357.300 ;
        RECT 165.550 357.040 165.880 357.300 ;
        RECT 167.090 357.160 167.350 357.300 ;
        RECT 168.090 357.160 168.270 357.600 ;
        RECT 168.820 357.390 170.180 357.500 ;
        RECT 168.820 357.330 170.260 357.390 ;
        RECT 169.620 357.320 170.260 357.330 ;
        RECT 164.110 356.850 164.340 356.860 ;
        RECT 167.090 356.990 168.270 357.160 ;
        RECT 169.790 357.220 170.260 357.320 ;
        RECT 170.730 357.240 171.690 357.410 ;
        RECT 205.590 357.400 205.790 357.750 ;
        RECT 207.070 357.480 207.600 357.650 ;
        RECT 167.090 356.850 167.350 356.990 ;
        RECT 169.790 356.970 170.040 357.220 ;
        RECT 164.110 356.680 164.870 356.850 ;
        RECT 165.120 356.680 166.290 356.850 ;
        RECT 166.530 356.820 167.350 356.850 ;
        RECT 168.590 356.820 168.770 356.880 ;
        RECT 166.530 356.680 167.640 356.820 ;
        RECT 165.520 356.580 165.870 356.680 ;
        RECT 167.180 356.650 167.640 356.680 ;
        RECT 168.090 356.650 168.770 356.820 ;
        RECT 169.710 356.800 170.040 356.970 ;
        RECT 171.510 356.780 171.690 357.240 ;
        RECT 209.760 357.170 214.810 358.020 ;
        RECT 232.510 357.890 232.690 358.820 ;
        RECT 233.240 358.560 233.570 358.730 ;
        RECT 233.750 358.610 234.080 358.870 ;
        RECT 234.330 358.710 234.910 358.970 ;
        RECT 235.100 359.010 235.340 359.160 ;
        RECT 235.100 358.830 235.700 359.010 ;
        RECT 234.560 358.680 234.910 358.710 ;
        RECT 233.320 358.420 233.570 358.560 ;
        RECT 233.320 358.230 233.800 358.420 ;
        RECT 233.160 358.160 233.800 358.230 ;
        RECT 233.160 358.060 233.490 358.160 ;
        RECT 232.390 357.860 232.710 357.890 ;
        RECT 232.390 357.670 232.720 357.860 ;
        RECT 232.390 357.630 232.710 357.670 ;
        RECT 168.130 356.630 168.770 356.650 ;
        RECT 168.590 356.620 168.770 356.630 ;
        RECT 170.370 356.620 170.970 356.770 ;
        RECT 168.590 356.600 170.970 356.620 ;
        RECT 171.430 356.610 171.760 356.780 ;
        RECT 168.590 356.450 170.820 356.600 ;
        RECT 190.910 356.530 191.110 356.880 ;
        RECT 192.650 356.800 192.970 356.810 ;
        RECT 192.390 356.630 192.970 356.800 ;
        RECT 192.640 356.580 192.970 356.630 ;
        RECT 192.650 356.550 192.970 356.580 ;
        RECT 213.450 356.800 213.770 356.810 ;
        RECT 213.450 356.630 214.030 356.800 ;
        RECT 213.450 356.580 213.780 356.630 ;
        RECT 213.450 356.550 213.770 356.580 ;
        RECT 190.900 356.500 191.110 356.530 ;
        RECT 215.310 356.530 215.510 356.880 ;
        RECT 9.190 356.370 9.710 356.390 ;
        RECT 3.140 354.890 8.850 354.900 ;
        RECT 3.060 354.720 8.850 354.890 ;
        RECT 3.150 354.710 8.850 354.720 ;
        RECT 8.620 354.640 8.790 354.710 ;
        RECT 9.190 354.590 9.720 356.370 ;
        RECT 190.900 355.910 191.120 356.500 ;
        RECT 191.640 355.940 191.840 356.510 ;
        RECT 192.650 356.220 192.970 356.260 ;
        RECT 192.640 356.180 192.970 356.220 ;
        RECT 192.390 356.010 192.970 356.180 ;
        RECT 192.650 356.000 192.970 356.010 ;
        RECT 213.450 356.220 213.770 356.260 ;
        RECT 213.450 356.180 213.780 356.220 ;
        RECT 213.450 356.010 214.030 356.180 ;
        RECT 213.450 356.000 213.770 356.010 ;
        RECT 190.900 354.880 191.120 355.470 ;
        RECT 193.650 355.450 193.820 355.960 ;
        RECT 197.590 355.460 197.760 355.970 ;
        RECT 208.660 355.460 208.830 355.970 ;
        RECT 212.600 355.450 212.770 355.960 ;
        RECT 214.580 355.940 214.780 356.510 ;
        RECT 215.310 356.500 215.520 356.530 ;
        RECT 215.300 355.910 215.520 356.500 ;
        RECT 217.640 355.720 217.840 356.730 ;
        RECT 223.390 355.720 223.680 356.730 ;
        RECT 190.900 354.850 191.110 354.880 ;
        RECT 191.640 354.870 191.840 355.440 ;
        RECT 192.650 355.370 192.970 355.380 ;
        RECT 192.390 355.200 192.970 355.370 ;
        RECT 192.640 355.160 192.970 355.200 ;
        RECT 192.650 355.120 192.970 355.160 ;
        RECT 213.450 355.370 213.770 355.380 ;
        RECT 213.450 355.200 214.030 355.370 ;
        RECT 213.450 355.160 213.780 355.200 ;
        RECT 213.450 355.120 213.770 355.160 ;
        RECT 214.580 354.870 214.780 355.440 ;
        RECT 215.300 354.880 215.520 355.470 ;
        RECT 9.200 354.570 9.720 354.590 ;
        RECT 2.180 353.850 4.620 354.140 ;
        RECT 9.200 354.060 9.710 354.570 ;
        RECT 190.910 354.500 191.110 354.850 ;
        RECT 215.310 354.850 215.520 354.880 ;
        RECT 192.650 354.800 192.970 354.830 ;
        RECT 192.640 354.750 192.970 354.800 ;
        RECT 213.450 354.800 213.770 354.830 ;
        RECT 192.390 354.580 192.970 354.750 ;
        RECT 192.650 354.570 192.970 354.580 ;
        RECT 191.280 354.100 191.720 354.270 ;
        RECT 9.200 353.850 9.730 354.060 ;
        RECT 2.180 353.370 9.730 353.850 ;
        RECT 190.910 353.520 191.110 353.870 ;
        RECT 192.650 353.790 192.970 353.800 ;
        RECT 192.390 353.620 192.970 353.790 ;
        RECT 192.640 353.570 192.970 353.620 ;
        RECT 193.650 353.610 193.820 354.620 ;
        RECT 195.580 353.890 196.130 354.320 ;
        RECT 197.580 353.750 197.750 354.760 ;
        RECT 199.610 353.960 200.160 354.390 ;
        RECT 206.260 353.960 206.810 354.390 ;
        RECT 208.670 353.750 208.840 354.760 ;
        RECT 213.450 354.750 213.780 354.800 ;
        RECT 210.290 353.890 210.840 354.320 ;
        RECT 212.600 353.610 212.770 354.620 ;
        RECT 213.450 354.580 214.030 354.750 ;
        RECT 213.450 354.570 213.770 354.580 ;
        RECT 215.310 354.500 215.510 354.850 ;
        RECT 214.700 354.100 215.140 354.270 ;
        RECT 213.450 353.790 213.770 353.800 ;
        RECT 213.450 353.620 214.030 353.790 ;
        RECT 192.650 353.540 192.970 353.570 ;
        RECT 213.450 353.570 213.780 353.620 ;
        RECT 213.450 353.540 213.770 353.570 ;
        RECT 190.900 353.490 191.110 353.520 ;
        RECT 215.310 353.520 215.510 353.870 ;
        RECT 232.510 353.720 232.690 357.630 ;
        RECT 233.320 356.780 233.490 358.060 ;
        RECT 233.910 358.040 234.080 358.610 ;
        RECT 234.150 358.320 234.320 358.360 ;
        RECT 234.740 358.350 234.910 358.680 ;
        RECT 235.110 358.530 235.700 358.830 ;
        RECT 236.520 358.890 237.100 359.060 ;
        RECT 236.520 358.790 236.910 358.890 ;
        RECT 236.520 358.760 236.900 358.790 ;
        RECT 236.520 358.610 236.880 358.760 ;
        RECT 234.560 358.320 234.910 358.350 ;
        RECT 234.150 358.060 234.910 358.320 ;
        RECT 234.150 358.030 234.320 358.060 ;
        RECT 234.560 358.030 234.910 358.060 ;
        RECT 234.560 358.020 234.760 358.030 ;
        RECT 235.150 358.020 235.700 358.530 ;
        RECT 236.170 358.440 236.880 358.610 ;
        RECT 235.460 357.780 235.680 358.020 ;
        RECT 235.470 357.750 235.680 357.780 ;
        RECT 233.660 357.520 234.190 357.650 ;
        RECT 235.470 357.530 235.670 357.750 ;
        RECT 236.170 357.690 236.870 358.000 ;
        RECT 233.660 357.490 234.320 357.520 ;
        RECT 234.560 357.490 234.760 357.530 ;
        RECT 233.660 357.480 234.760 357.490 ;
        RECT 234.150 357.230 234.760 357.480 ;
        RECT 234.150 357.190 234.320 357.230 ;
        RECT 234.560 357.200 234.760 357.230 ;
        RECT 234.560 356.840 234.760 356.870 ;
        RECT 233.120 356.580 233.440 356.610 ;
        RECT 234.330 356.580 234.760 356.840 ;
        RECT 233.120 356.390 233.450 356.580 ;
        RECT 234.560 356.540 234.760 356.580 ;
        RECT 235.150 356.540 235.700 357.530 ;
        RECT 236.020 357.460 236.870 357.690 ;
        RECT 236.170 357.120 236.870 357.460 ;
        RECT 236.630 356.760 236.950 356.800 ;
        RECT 236.630 356.700 236.960 356.760 ;
        RECT 236.160 356.570 236.960 356.700 ;
        RECT 236.160 356.540 236.950 356.570 ;
        RECT 236.160 356.520 236.860 356.540 ;
        RECT 233.120 356.350 233.440 356.390 ;
        RECT 233.120 356.270 233.290 356.350 ;
        RECT 233.070 356.100 233.290 356.270 ;
        RECT 233.070 355.940 233.240 356.100 ;
        RECT 234.560 356.010 234.760 356.050 ;
        RECT 233.600 355.680 233.790 355.800 ;
        RECT 234.330 355.750 234.760 356.010 ;
        RECT 234.560 355.720 234.760 355.750 ;
        RECT 233.240 355.570 233.790 355.680 ;
        RECT 233.240 355.510 233.780 355.570 ;
        RECT 233.320 353.730 233.490 355.510 ;
        RECT 234.150 355.360 234.320 355.400 ;
        RECT 234.560 355.360 234.760 355.390 ;
        RECT 234.150 355.100 234.760 355.360 ;
        RECT 234.150 355.070 234.320 355.100 ;
        RECT 234.560 355.060 234.760 355.100 ;
        RECT 235.150 355.060 235.700 356.050 ;
        RECT 236.620 356.040 236.940 356.080 ;
        RECT 236.160 355.860 236.950 356.040 ;
        RECT 236.620 355.850 236.950 355.860 ;
        RECT 236.620 355.820 236.940 355.850 ;
        RECT 363.700 355.670 364.210 366.030 ;
        RECT 364.380 365.240 370.360 365.470 ;
        RECT 363.700 355.650 364.220 355.670 ;
        RECT 236.170 355.100 236.870 355.440 ;
        RECT 236.020 354.870 236.870 355.100 ;
        RECT 234.150 354.530 234.320 354.560 ;
        RECT 234.560 354.530 234.760 354.570 ;
        RECT 234.150 354.270 234.760 354.530 ;
        RECT 234.150 354.230 234.320 354.270 ;
        RECT 234.560 354.240 234.760 354.270 ;
        RECT 234.560 353.880 234.760 353.910 ;
        RECT 234.330 353.620 234.760 353.880 ;
        RECT 234.560 353.580 234.760 353.620 ;
        RECT 235.150 353.580 235.700 354.570 ;
        RECT 236.170 354.560 236.870 354.870 ;
        RECT 236.170 353.950 236.880 354.120 ;
        RECT 236.520 353.670 236.880 353.950 ;
        RECT 363.690 353.870 364.220 355.650 ;
        RECT 364.620 354.180 370.270 365.240 ;
        RECT 364.560 354.170 370.270 354.180 ;
        RECT 364.560 354.000 370.350 354.170 ;
        RECT 364.560 353.990 370.260 354.000 ;
        RECT 364.620 353.920 364.790 353.990 ;
        RECT 363.690 353.850 364.210 353.870 ;
        RECT 2.180 353.340 9.540 353.370 ;
        RECT 183.480 352.600 183.650 353.020 ;
        RECT 184.290 352.900 184.530 352.930 ;
        RECT 183.960 352.730 184.530 352.900 ;
        RECT 184.770 352.730 186.110 352.900 ;
        RECT 186.560 352.730 187.520 352.900 ;
        RECT 184.290 352.690 184.530 352.730 ;
        RECT 187.070 352.720 187.240 352.730 ;
        RECT 183.410 352.380 183.580 352.420 ;
        RECT 163.520 352.180 163.690 352.230 ;
        RECT 183.350 352.210 183.580 352.380 ;
        RECT 2.180 351.580 9.710 352.130 ;
        RECT 163.490 351.960 163.710 352.180 ;
        RECT 163.520 351.900 163.690 351.960 ;
        RECT 164.040 351.820 164.370 352.000 ;
        RECT 167.180 351.990 167.350 352.040 ;
        RECT 164.620 351.820 166.780 351.990 ;
        RECT 167.020 351.820 167.350 351.990 ;
        RECT 167.640 351.850 167.850 352.180 ;
        RECT 0.500 338.610 1.970 338.860 ;
        RECT 2.180 338.670 2.690 351.580 ;
        RECT 9.040 351.570 9.710 351.580 ;
        RECT 5.340 350.680 8.800 351.120 ;
        RECT 3.410 350.580 8.800 350.680 ;
        RECT 3.410 350.510 8.690 350.580 ;
        RECT 3.410 339.600 3.580 350.510 ;
        RECT 3.910 350.100 8.140 350.120 ;
        RECT 3.890 339.990 8.220 350.100 ;
        RECT 3.950 339.940 4.120 339.990 ;
        RECT 8.520 339.600 8.690 350.510 ;
        RECT 3.410 339.430 8.690 339.600 ;
        RECT 8.450 339.420 8.690 339.430 ;
        RECT 9.200 338.670 9.710 351.570 ;
        RECT 164.070 351.380 164.340 351.820 ;
        RECT 165.550 351.560 165.880 351.820 ;
        RECT 167.090 351.680 167.350 351.820 ;
        RECT 168.090 351.680 168.270 352.120 ;
        RECT 168.820 351.910 170.180 352.020 ;
        RECT 168.820 351.850 170.260 351.910 ;
        RECT 169.620 351.840 170.260 351.850 ;
        RECT 164.110 351.370 164.340 351.380 ;
        RECT 167.090 351.510 168.270 351.680 ;
        RECT 169.790 351.740 170.260 351.840 ;
        RECT 170.730 351.760 171.690 351.930 ;
        RECT 183.410 351.860 183.580 352.210 ;
        RECT 183.750 352.280 183.940 352.300 ;
        RECT 186.750 352.280 187.080 352.460 ;
        RECT 183.750 352.110 184.310 352.280 ;
        RECT 184.770 352.110 187.520 352.280 ;
        RECT 183.750 352.070 183.940 352.110 ;
        RECT 188.050 352.040 188.220 352.970 ;
        RECT 188.450 352.170 188.620 353.020 ;
        RECT 190.900 352.900 191.120 353.490 ;
        RECT 191.640 352.930 191.840 353.500 ;
        RECT 192.650 353.210 192.970 353.250 ;
        RECT 192.640 353.170 192.970 353.210 ;
        RECT 192.390 353.000 192.970 353.170 ;
        RECT 192.650 352.990 192.970 353.000 ;
        RECT 213.450 353.210 213.770 353.250 ;
        RECT 213.450 353.170 213.780 353.210 ;
        RECT 213.450 353.000 214.030 353.170 ;
        RECT 213.450 352.990 213.770 353.000 ;
        RECT 214.580 352.930 214.780 353.500 ;
        RECT 215.310 353.490 215.520 353.520 ;
        RECT 236.520 353.500 237.100 353.670 ;
        RECT 215.300 352.900 215.520 353.490 ;
        RECT 363.700 353.340 364.210 353.850 ;
        RECT 370.720 353.420 371.230 366.030 ;
        RECT 371.470 360.010 372.930 360.050 ;
        RECT 371.460 359.840 372.930 360.010 ;
        RECT 371.470 359.800 372.930 359.840 ;
        RECT 363.680 353.130 364.210 353.340 ;
        RECT 368.790 353.130 371.230 353.420 ;
        RECT 363.680 352.650 371.230 353.130 ;
        RECT 363.870 352.620 371.230 352.650 ;
        RECT 190.900 351.880 191.120 352.470 ;
        RECT 190.900 351.850 191.110 351.880 ;
        RECT 191.640 351.870 191.840 352.440 ;
        RECT 192.650 352.370 192.970 352.380 ;
        RECT 192.390 352.200 192.970 352.370 ;
        RECT 192.640 352.160 192.970 352.200 ;
        RECT 192.650 352.120 192.970 352.160 ;
        RECT 213.450 352.370 213.770 352.380 ;
        RECT 213.450 352.200 214.030 352.370 ;
        RECT 213.450 352.160 213.780 352.200 ;
        RECT 213.450 352.120 213.770 352.160 ;
        RECT 214.580 351.870 214.780 352.440 ;
        RECT 215.300 351.880 215.520 352.470 ;
        RECT 167.090 351.370 167.350 351.510 ;
        RECT 169.790 351.490 170.040 351.740 ;
        RECT 164.110 351.200 164.870 351.370 ;
        RECT 165.120 351.200 166.290 351.370 ;
        RECT 166.530 351.340 167.350 351.370 ;
        RECT 168.590 351.340 168.770 351.400 ;
        RECT 166.530 351.200 167.640 351.340 ;
        RECT 165.520 351.100 165.870 351.200 ;
        RECT 167.180 351.170 167.640 351.200 ;
        RECT 168.090 351.170 168.770 351.340 ;
        RECT 169.710 351.320 170.040 351.490 ;
        RECT 171.510 351.300 171.690 351.760 ;
        RECT 168.130 351.150 168.770 351.170 ;
        RECT 168.590 351.140 168.770 351.150 ;
        RECT 170.370 351.140 170.970 351.290 ;
        RECT 168.590 351.120 170.970 351.140 ;
        RECT 171.430 351.130 171.760 351.300 ;
        RECT 183.410 351.270 183.580 351.620 ;
        RECT 190.910 351.500 191.110 351.850 ;
        RECT 215.310 351.850 215.520 351.880 ;
        RECT 192.650 351.800 192.970 351.830 ;
        RECT 192.640 351.750 192.970 351.800 ;
        RECT 192.390 351.580 192.970 351.750 ;
        RECT 192.650 351.570 192.970 351.580 ;
        RECT 213.450 351.800 213.770 351.830 ;
        RECT 213.450 351.750 213.780 351.800 ;
        RECT 213.450 351.580 214.030 351.750 ;
        RECT 213.450 351.570 213.770 351.580 ;
        RECT 215.310 351.500 215.510 351.850 ;
        RECT 168.590 350.970 170.820 351.120 ;
        RECT 183.350 351.100 183.580 351.270 ;
        RECT 183.750 351.370 183.940 351.410 ;
        RECT 183.750 351.200 184.310 351.370 ;
        RECT 184.770 351.200 187.520 351.370 ;
        RECT 183.750 351.180 183.940 351.200 ;
        RECT 183.410 351.060 183.580 351.100 ;
        RECT 186.750 351.020 187.080 351.200 ;
        RECT 163.520 350.630 163.690 350.680 ;
        RECT 163.490 350.410 163.710 350.630 ;
        RECT 163.520 350.350 163.690 350.410 ;
        RECT 164.040 350.270 164.370 350.450 ;
        RECT 167.180 350.440 167.350 350.490 ;
        RECT 164.620 350.270 166.780 350.440 ;
        RECT 167.020 350.270 167.350 350.440 ;
        RECT 167.640 350.300 167.850 350.630 ;
        RECT 164.070 349.830 164.340 350.270 ;
        RECT 165.550 350.010 165.880 350.270 ;
        RECT 167.090 350.130 167.350 350.270 ;
        RECT 168.090 350.130 168.270 350.570 ;
        RECT 168.820 350.360 170.180 350.470 ;
        RECT 183.480 350.460 183.650 350.880 ;
        RECT 184.290 350.750 184.530 350.790 ;
        RECT 187.070 350.750 187.240 350.760 ;
        RECT 183.960 350.580 184.530 350.750 ;
        RECT 184.770 350.580 186.110 350.750 ;
        RECT 186.560 350.580 187.520 350.750 ;
        RECT 184.290 350.550 184.530 350.580 ;
        RECT 188.050 350.510 188.220 351.440 ;
        RECT 188.450 350.460 188.620 351.310 ;
        RECT 363.700 350.860 371.230 351.410 ;
        RECT 363.700 350.850 364.370 350.860 ;
        RECT 168.820 350.300 170.260 350.360 ;
        RECT 169.620 350.290 170.260 350.300 ;
        RECT 164.110 349.820 164.340 349.830 ;
        RECT 167.090 349.960 168.270 350.130 ;
        RECT 169.790 350.190 170.260 350.290 ;
        RECT 170.730 350.210 171.690 350.380 ;
        RECT 167.090 349.820 167.350 349.960 ;
        RECT 169.790 349.940 170.040 350.190 ;
        RECT 164.110 349.650 164.870 349.820 ;
        RECT 165.120 349.650 166.290 349.820 ;
        RECT 166.530 349.790 167.350 349.820 ;
        RECT 168.590 349.790 168.770 349.850 ;
        RECT 166.530 349.650 167.640 349.790 ;
        RECT 165.520 349.550 165.870 349.650 ;
        RECT 167.180 349.620 167.640 349.650 ;
        RECT 168.090 349.620 168.770 349.790 ;
        RECT 169.710 349.770 170.040 349.940 ;
        RECT 171.510 349.750 171.690 350.210 ;
        RECT 168.130 349.600 168.770 349.620 ;
        RECT 168.590 349.590 168.770 349.600 ;
        RECT 170.370 349.590 170.970 349.740 ;
        RECT 168.590 349.570 170.970 349.590 ;
        RECT 171.430 349.580 171.760 349.750 ;
        RECT 183.480 349.670 183.650 350.090 ;
        RECT 184.290 349.970 184.530 350.000 ;
        RECT 183.960 349.800 184.530 349.970 ;
        RECT 184.770 349.800 186.110 349.970 ;
        RECT 186.560 349.800 187.520 349.970 ;
        RECT 184.290 349.760 184.530 349.800 ;
        RECT 187.070 349.790 187.240 349.800 ;
        RECT 168.590 349.420 170.820 349.570 ;
        RECT 183.410 349.450 183.580 349.490 ;
        RECT 183.350 349.280 183.580 349.450 ;
        RECT 163.520 349.080 163.690 349.130 ;
        RECT 163.490 348.860 163.710 349.080 ;
        RECT 163.520 348.800 163.690 348.860 ;
        RECT 164.040 348.720 164.370 348.900 ;
        RECT 167.180 348.890 167.350 348.940 ;
        RECT 164.620 348.720 166.780 348.890 ;
        RECT 167.020 348.720 167.350 348.890 ;
        RECT 167.640 348.750 167.850 349.080 ;
        RECT 164.070 348.280 164.340 348.720 ;
        RECT 165.550 348.460 165.880 348.720 ;
        RECT 167.090 348.580 167.350 348.720 ;
        RECT 168.090 348.580 168.270 349.020 ;
        RECT 183.410 348.930 183.580 349.280 ;
        RECT 183.750 349.350 183.940 349.370 ;
        RECT 186.750 349.350 187.080 349.530 ;
        RECT 183.750 349.180 184.310 349.350 ;
        RECT 184.770 349.180 187.520 349.350 ;
        RECT 183.750 349.140 183.940 349.180 ;
        RECT 188.050 349.110 188.220 350.040 ;
        RECT 188.450 349.240 188.620 350.090 ;
        RECT 168.820 348.810 170.180 348.920 ;
        RECT 168.820 348.750 170.260 348.810 ;
        RECT 169.620 348.740 170.260 348.750 ;
        RECT 164.110 348.270 164.340 348.280 ;
        RECT 167.090 348.410 168.270 348.580 ;
        RECT 169.790 348.640 170.260 348.740 ;
        RECT 170.730 348.660 171.690 348.830 ;
        RECT 167.090 348.270 167.350 348.410 ;
        RECT 169.790 348.390 170.040 348.640 ;
        RECT 164.110 348.100 164.870 348.270 ;
        RECT 165.120 348.100 166.290 348.270 ;
        RECT 166.530 348.240 167.350 348.270 ;
        RECT 168.590 348.240 168.770 348.300 ;
        RECT 166.530 348.100 167.640 348.240 ;
        RECT 165.520 348.000 165.870 348.100 ;
        RECT 167.180 348.070 167.640 348.100 ;
        RECT 168.090 348.070 168.770 348.240 ;
        RECT 169.710 348.220 170.040 348.390 ;
        RECT 171.510 348.200 171.690 348.660 ;
        RECT 183.410 348.340 183.580 348.690 ;
        RECT 168.130 348.050 168.770 348.070 ;
        RECT 168.590 348.040 168.770 348.050 ;
        RECT 170.370 348.040 170.970 348.190 ;
        RECT 168.590 348.020 170.970 348.040 ;
        RECT 171.430 348.030 171.760 348.200 ;
        RECT 183.350 348.170 183.580 348.340 ;
        RECT 183.750 348.440 183.940 348.480 ;
        RECT 183.750 348.270 184.310 348.440 ;
        RECT 184.770 348.270 187.520 348.440 ;
        RECT 183.750 348.250 183.940 348.270 ;
        RECT 183.410 348.130 183.580 348.170 ;
        RECT 186.750 348.090 187.080 348.270 ;
        RECT 168.590 347.870 170.820 348.020 ;
        RECT 163.520 347.530 163.690 347.580 ;
        RECT 183.480 347.530 183.650 347.950 ;
        RECT 184.290 347.820 184.530 347.860 ;
        RECT 187.070 347.820 187.240 347.830 ;
        RECT 183.960 347.650 184.530 347.820 ;
        RECT 184.770 347.650 186.110 347.820 ;
        RECT 186.560 347.650 187.520 347.820 ;
        RECT 184.290 347.620 184.530 347.650 ;
        RECT 188.050 347.580 188.220 348.510 ;
        RECT 188.450 347.530 188.620 348.380 ;
        RECT 163.490 347.310 163.710 347.530 ;
        RECT 163.520 347.250 163.690 347.310 ;
        RECT 164.040 347.170 164.370 347.350 ;
        RECT 167.180 347.340 167.350 347.390 ;
        RECT 164.620 347.170 166.780 347.340 ;
        RECT 167.020 347.170 167.350 347.340 ;
        RECT 167.640 347.200 167.850 347.530 ;
        RECT 164.070 346.730 164.340 347.170 ;
        RECT 165.550 346.910 165.880 347.170 ;
        RECT 167.090 347.030 167.350 347.170 ;
        RECT 168.090 347.030 168.270 347.470 ;
        RECT 168.820 347.260 170.180 347.370 ;
        RECT 168.820 347.200 170.260 347.260 ;
        RECT 169.620 347.190 170.260 347.200 ;
        RECT 164.110 346.720 164.340 346.730 ;
        RECT 167.090 346.860 168.270 347.030 ;
        RECT 169.790 347.090 170.260 347.190 ;
        RECT 170.730 347.110 171.690 347.280 ;
        RECT 191.490 347.140 191.690 347.490 ;
        RECT 193.230 347.410 193.550 347.420 ;
        RECT 192.970 347.240 193.550 347.410 ;
        RECT 193.220 347.190 193.550 347.240 ;
        RECT 193.230 347.160 193.550 347.190 ;
        RECT 167.090 346.720 167.350 346.860 ;
        RECT 169.790 346.840 170.040 347.090 ;
        RECT 164.110 346.550 164.870 346.720 ;
        RECT 165.120 346.550 166.290 346.720 ;
        RECT 166.530 346.690 167.350 346.720 ;
        RECT 168.590 346.690 168.770 346.750 ;
        RECT 166.530 346.550 167.640 346.690 ;
        RECT 165.520 346.450 165.870 346.550 ;
        RECT 167.180 346.520 167.640 346.550 ;
        RECT 168.090 346.520 168.770 346.690 ;
        RECT 169.710 346.670 170.040 346.840 ;
        RECT 171.510 346.650 171.690 347.110 ;
        RECT 191.480 347.110 191.690 347.140 ;
        RECT 168.130 346.500 168.770 346.520 ;
        RECT 168.590 346.490 168.770 346.500 ;
        RECT 170.370 346.490 170.970 346.640 ;
        RECT 168.590 346.470 170.970 346.490 ;
        RECT 171.430 346.480 171.760 346.650 ;
        RECT 191.480 346.520 191.700 347.110 ;
        RECT 192.220 346.550 192.420 347.120 ;
        RECT 193.230 346.830 193.550 346.870 ;
        RECT 193.220 346.790 193.550 346.830 ;
        RECT 192.970 346.620 193.550 346.790 ;
        RECT 193.230 346.610 193.550 346.620 ;
        RECT 168.590 346.320 170.820 346.470 ;
        RECT 191.480 345.490 191.700 346.080 ;
        RECT 191.480 345.460 191.690 345.490 ;
        RECT 192.220 345.480 192.420 346.050 ;
        RECT 194.360 346.040 194.530 346.550 ;
        RECT 198.380 346.070 198.550 346.580 ;
        RECT 193.230 345.980 193.550 345.990 ;
        RECT 192.970 345.810 193.550 345.980 ;
        RECT 193.220 345.770 193.550 345.810 ;
        RECT 193.230 345.730 193.550 345.770 ;
        RECT 191.490 345.110 191.690 345.460 ;
        RECT 193.230 345.410 193.550 345.440 ;
        RECT 193.220 345.360 193.550 345.410 ;
        RECT 192.970 345.190 193.550 345.360 ;
        RECT 193.230 345.180 193.550 345.190 ;
        RECT 191.860 344.710 192.300 344.880 ;
        RECT 140.590 343.790 140.760 344.280 ;
        RECT 140.440 343.760 140.760 343.790 ;
        RECT 141.140 343.790 141.310 344.280 ;
        RECT 141.780 344.230 141.950 344.280 ;
        RECT 142.330 344.230 142.500 344.280 ;
        RECT 141.660 344.200 141.980 344.230 ;
        RECT 142.310 344.200 142.630 344.230 ;
        RECT 141.660 344.010 141.990 344.200 ;
        RECT 142.310 344.010 142.640 344.200 ;
        RECT 191.490 344.130 191.690 344.480 ;
        RECT 193.230 344.400 193.550 344.410 ;
        RECT 192.970 344.230 193.550 344.400 ;
        RECT 193.220 344.180 193.550 344.230 ;
        RECT 194.350 344.180 194.520 345.370 ;
        RECT 196.160 344.500 196.710 344.930 ;
        RECT 193.230 344.150 193.550 344.180 ;
        RECT 191.480 344.100 191.690 344.130 ;
        RECT 198.370 344.120 198.540 345.310 ;
        RECT 200.190 344.570 200.740 345.000 ;
        RECT 141.660 343.970 141.980 344.010 ;
        RECT 142.310 343.970 142.630 344.010 ;
        RECT 141.140 343.760 141.460 343.790 ;
        RECT 140.440 343.570 140.770 343.760 ;
        RECT 141.140 343.570 141.470 343.760 ;
        RECT 140.440 343.530 140.760 343.570 ;
        RECT 140.050 342.070 140.220 342.090 ;
        RECT 140.030 341.640 140.240 342.070 ;
        RECT 140.590 341.880 140.760 343.530 ;
        RECT 141.140 343.530 141.460 343.570 ;
        RECT 141.140 341.880 141.310 343.530 ;
        RECT 141.780 341.880 141.950 343.970 ;
        RECT 142.330 341.880 142.500 343.970 ;
        RECT 191.480 343.510 191.700 344.100 ;
        RECT 192.220 343.540 192.420 344.110 ;
        RECT 193.230 343.820 193.550 343.860 ;
        RECT 193.220 343.780 193.550 343.820 ;
        RECT 192.970 343.610 193.550 343.780 ;
        RECT 193.230 343.600 193.550 343.610 ;
        RECT 204.600 343.480 204.920 343.510 ;
        RECT 142.880 342.520 143.050 343.370 ;
        RECT 204.600 343.310 206.390 343.480 ;
        RECT 204.600 343.290 204.930 343.310 ;
        RECT 183.480 342.840 183.650 343.260 ;
        RECT 184.290 343.140 184.530 343.170 ;
        RECT 183.960 342.970 184.530 343.140 ;
        RECT 184.770 342.970 186.110 343.140 ;
        RECT 186.560 342.970 187.520 343.140 ;
        RECT 184.290 342.930 184.530 342.970 ;
        RECT 187.070 342.960 187.240 342.970 ;
        RECT 183.410 342.620 183.580 342.660 ;
        RECT 163.520 342.410 163.690 342.460 ;
        RECT 183.350 342.450 183.580 342.620 ;
        RECT 163.490 342.190 163.710 342.410 ;
        RECT 163.520 342.130 163.690 342.190 ;
        RECT 164.040 342.050 164.370 342.230 ;
        RECT 167.180 342.220 167.350 342.270 ;
        RECT 164.620 342.050 166.780 342.220 ;
        RECT 167.020 342.050 167.350 342.220 ;
        RECT 167.640 342.080 167.850 342.410 ;
        RECT 142.770 341.890 143.200 341.910 ;
        RECT 142.770 341.720 143.220 341.890 ;
        RECT 142.770 341.700 143.200 341.720 ;
        RECT 164.070 341.610 164.340 342.050 ;
        RECT 165.550 341.790 165.880 342.050 ;
        RECT 167.090 341.910 167.350 342.050 ;
        RECT 168.090 341.910 168.270 342.350 ;
        RECT 168.820 342.140 170.180 342.250 ;
        RECT 168.820 342.080 170.260 342.140 ;
        RECT 169.620 342.070 170.260 342.080 ;
        RECT 164.110 341.600 164.340 341.610 ;
        RECT 167.090 341.740 168.270 341.910 ;
        RECT 169.790 341.970 170.260 342.070 ;
        RECT 170.730 341.990 171.690 342.160 ;
        RECT 183.410 342.100 183.580 342.450 ;
        RECT 183.750 342.520 183.940 342.540 ;
        RECT 186.750 342.520 187.080 342.700 ;
        RECT 183.750 342.350 184.310 342.520 ;
        RECT 184.770 342.350 187.520 342.520 ;
        RECT 183.750 342.310 183.940 342.350 ;
        RECT 188.050 342.280 188.220 343.210 ;
        RECT 188.450 342.410 188.620 343.260 ;
        RECT 204.600 343.250 204.920 343.290 ;
        RECT 206.220 343.080 206.390 343.310 ;
        RECT 191.480 342.490 191.700 343.080 ;
        RECT 191.480 342.460 191.690 342.490 ;
        RECT 192.220 342.480 192.420 343.050 ;
        RECT 193.230 342.980 193.550 342.990 ;
        RECT 192.970 342.810 193.550 342.980 ;
        RECT 205.070 342.830 205.410 343.080 ;
        RECT 205.580 342.910 205.910 343.080 ;
        RECT 206.130 342.910 206.470 343.080 ;
        RECT 193.220 342.770 193.550 342.810 ;
        RECT 193.230 342.730 193.550 342.770 ;
        RECT 204.750 342.570 205.410 342.830 ;
        RECT 205.660 342.740 205.830 342.910 ;
        RECT 206.220 342.740 206.390 342.910 ;
        RECT 205.580 342.570 205.910 342.740 ;
        RECT 206.130 342.570 206.470 342.740 ;
        RECT 191.490 342.110 191.690 342.460 ;
        RECT 193.230 342.410 193.550 342.440 ;
        RECT 193.220 342.360 193.550 342.410 ;
        RECT 192.970 342.190 193.550 342.360 ;
        RECT 193.230 342.180 193.550 342.190 ;
        RECT 205.660 342.340 205.910 342.570 ;
        RECT 206.790 342.490 207.300 343.160 ;
        RECT 205.660 342.170 206.330 342.340 ;
        RECT 167.090 341.600 167.350 341.740 ;
        RECT 169.790 341.720 170.040 341.970 ;
        RECT 164.110 341.430 164.870 341.600 ;
        RECT 165.120 341.430 166.290 341.600 ;
        RECT 166.530 341.570 167.350 341.600 ;
        RECT 168.590 341.570 168.770 341.630 ;
        RECT 166.530 341.430 167.640 341.570 ;
        RECT 2.180 338.160 9.710 338.670 ;
        RECT 139.130 338.520 139.300 341.010 ;
        RECT 139.680 338.520 139.850 341.020 ;
        RECT 140.040 341.000 140.250 341.430 ;
        RECT 142.780 341.350 143.210 341.370 ;
        RECT 142.780 341.180 143.230 341.350 ;
        RECT 165.520 341.330 165.870 341.430 ;
        RECT 167.180 341.400 167.640 341.430 ;
        RECT 168.090 341.400 168.770 341.570 ;
        RECT 169.710 341.550 170.040 341.720 ;
        RECT 171.510 341.530 171.690 341.990 ;
        RECT 205.660 341.940 205.910 342.170 ;
        RECT 168.130 341.380 168.770 341.400 ;
        RECT 168.590 341.370 168.770 341.380 ;
        RECT 170.370 341.370 170.970 341.520 ;
        RECT 168.590 341.350 170.970 341.370 ;
        RECT 171.430 341.360 171.760 341.530 ;
        RECT 183.410 341.510 183.580 341.860 ;
        RECT 204.750 341.680 205.410 341.940 ;
        RECT 205.580 341.770 205.910 341.940 ;
        RECT 206.130 341.770 206.470 341.940 ;
        RECT 168.590 341.200 170.820 341.350 ;
        RECT 183.350 341.340 183.580 341.510 ;
        RECT 183.750 341.610 183.940 341.650 ;
        RECT 183.750 341.440 184.310 341.610 ;
        RECT 184.770 341.440 187.520 341.610 ;
        RECT 183.750 341.420 183.940 341.440 ;
        RECT 183.410 341.300 183.580 341.340 ;
        RECT 186.750 341.260 187.080 341.440 ;
        RECT 142.780 341.160 143.210 341.180 ;
        RECT 140.060 340.980 140.230 341.000 ;
        RECT 140.310 339.910 140.480 341.010 ;
        RECT 140.310 339.880 140.790 339.910 ;
        RECT 140.310 339.690 140.800 339.880 ;
        RECT 140.310 339.650 140.790 339.690 ;
        RECT 140.310 338.520 140.480 339.650 ;
        RECT 140.860 338.520 141.030 341.020 ;
        RECT 163.520 340.860 163.690 340.910 ;
        RECT 163.490 340.640 163.710 340.860 ;
        RECT 142.870 339.970 143.040 340.640 ;
        RECT 163.520 340.580 163.690 340.640 ;
        RECT 164.040 340.500 164.370 340.680 ;
        RECT 167.180 340.670 167.350 340.720 ;
        RECT 164.620 340.500 166.780 340.670 ;
        RECT 167.020 340.500 167.350 340.670 ;
        RECT 167.640 340.530 167.850 340.860 ;
        RECT 164.070 340.060 164.340 340.500 ;
        RECT 165.550 340.240 165.880 340.500 ;
        RECT 167.090 340.360 167.350 340.500 ;
        RECT 168.090 340.360 168.270 340.800 ;
        RECT 183.480 340.700 183.650 341.120 ;
        RECT 184.290 340.990 184.530 341.030 ;
        RECT 187.070 340.990 187.240 341.000 ;
        RECT 183.960 340.820 184.530 340.990 ;
        RECT 184.770 340.820 186.110 340.990 ;
        RECT 186.560 340.820 187.520 340.990 ;
        RECT 184.290 340.790 184.530 340.820 ;
        RECT 188.050 340.750 188.220 341.680 ;
        RECT 188.450 340.700 188.620 341.550 ;
        RECT 205.070 341.430 205.410 341.680 ;
        RECT 205.660 341.600 205.830 341.770 ;
        RECT 206.220 341.600 206.390 341.770 ;
        RECT 205.580 341.430 205.910 341.600 ;
        RECT 206.130 341.430 206.470 341.600 ;
        RECT 204.600 341.220 204.920 341.260 ;
        RECT 204.600 341.200 204.930 341.220 ;
        RECT 206.220 341.200 206.390 341.430 ;
        RECT 206.790 341.350 207.300 342.020 ;
        RECT 204.600 341.030 206.390 341.200 ;
        RECT 204.600 341.000 204.920 341.030 ;
        RECT 204.600 340.710 204.920 340.740 ;
        RECT 168.820 340.590 170.180 340.700 ;
        RECT 168.820 340.530 170.260 340.590 ;
        RECT 169.620 340.520 170.260 340.530 ;
        RECT 164.110 340.050 164.340 340.060 ;
        RECT 167.090 340.190 168.270 340.360 ;
        RECT 169.790 340.420 170.260 340.520 ;
        RECT 170.730 340.440 171.690 340.610 ;
        RECT 204.600 340.540 206.390 340.710 ;
        RECT 204.600 340.520 204.930 340.540 ;
        RECT 204.600 340.480 204.920 340.520 ;
        RECT 167.090 340.050 167.350 340.190 ;
        RECT 169.790 340.170 170.040 340.420 ;
        RECT 141.160 339.870 141.480 339.900 ;
        RECT 164.110 339.880 164.870 340.050 ;
        RECT 165.120 339.880 166.290 340.050 ;
        RECT 166.530 340.020 167.350 340.050 ;
        RECT 168.590 340.020 168.770 340.080 ;
        RECT 166.530 339.880 167.640 340.020 ;
        RECT 141.160 339.680 141.490 339.870 ;
        RECT 165.520 339.780 165.870 339.880 ;
        RECT 167.180 339.850 167.640 339.880 ;
        RECT 168.090 339.850 168.770 340.020 ;
        RECT 169.710 340.000 170.040 340.170 ;
        RECT 171.510 339.980 171.690 340.440 ;
        RECT 168.130 339.830 168.770 339.850 ;
        RECT 168.590 339.820 168.770 339.830 ;
        RECT 170.370 339.820 170.970 339.970 ;
        RECT 168.590 339.800 170.970 339.820 ;
        RECT 171.430 339.810 171.760 339.980 ;
        RECT 183.480 339.910 183.650 340.330 ;
        RECT 184.290 340.210 184.530 340.240 ;
        RECT 183.960 340.040 184.530 340.210 ;
        RECT 184.770 340.040 186.110 340.210 ;
        RECT 186.560 340.040 187.520 340.210 ;
        RECT 184.290 340.000 184.530 340.040 ;
        RECT 187.070 340.030 187.240 340.040 ;
        RECT 141.160 339.640 141.480 339.680 ;
        RECT 168.590 339.650 170.820 339.800 ;
        RECT 183.410 339.690 183.580 339.730 ;
        RECT 183.350 339.520 183.580 339.690 ;
        RECT 163.520 339.310 163.690 339.360 ;
        RECT 141.640 339.100 141.960 339.130 ;
        RECT 141.640 338.910 141.970 339.100 ;
        RECT 163.490 339.090 163.710 339.310 ;
        RECT 142.350 339.040 142.670 339.070 ;
        RECT 141.640 338.870 141.960 338.910 ;
        RECT 142.350 338.850 142.680 339.040 ;
        RECT 163.520 339.030 163.690 339.090 ;
        RECT 164.040 338.950 164.370 339.130 ;
        RECT 167.180 339.120 167.350 339.170 ;
        RECT 164.620 338.950 166.780 339.120 ;
        RECT 167.020 338.950 167.350 339.120 ;
        RECT 167.640 338.980 167.850 339.310 ;
        RECT 142.350 338.810 142.670 338.850 ;
        RECT 164.070 338.510 164.340 338.950 ;
        RECT 165.550 338.690 165.880 338.950 ;
        RECT 167.090 338.810 167.350 338.950 ;
        RECT 168.090 338.810 168.270 339.250 ;
        RECT 183.410 339.170 183.580 339.520 ;
        RECT 183.750 339.590 183.940 339.610 ;
        RECT 186.750 339.590 187.080 339.770 ;
        RECT 183.750 339.420 184.310 339.590 ;
        RECT 184.770 339.420 187.520 339.590 ;
        RECT 183.750 339.380 183.940 339.420 ;
        RECT 188.050 339.350 188.220 340.280 ;
        RECT 188.450 339.480 188.620 340.330 ;
        RECT 206.220 340.310 206.390 340.540 ;
        RECT 205.070 340.060 205.410 340.310 ;
        RECT 205.580 340.140 205.910 340.310 ;
        RECT 206.130 340.140 206.470 340.310 ;
        RECT 204.750 339.800 205.410 340.060 ;
        RECT 205.660 339.970 205.830 340.140 ;
        RECT 206.220 339.970 206.390 340.140 ;
        RECT 205.580 339.800 205.910 339.970 ;
        RECT 206.130 339.800 206.470 339.970 ;
        RECT 205.660 339.570 205.910 339.800 ;
        RECT 206.790 339.720 207.300 340.390 ;
        RECT 205.660 339.400 206.330 339.570 ;
        RECT 205.660 339.170 205.910 339.400 ;
        RECT 168.820 339.040 170.180 339.150 ;
        RECT 193.160 339.070 193.480 339.110 ;
        RECT 168.820 338.980 170.260 339.040 ;
        RECT 169.620 338.970 170.260 338.980 ;
        RECT 164.110 338.500 164.340 338.510 ;
        RECT 167.090 338.640 168.270 338.810 ;
        RECT 169.790 338.870 170.260 338.970 ;
        RECT 170.730 338.890 171.690 339.060 ;
        RECT 167.090 338.500 167.350 338.640 ;
        RECT 169.790 338.620 170.040 338.870 ;
        RECT 164.110 338.330 164.870 338.500 ;
        RECT 165.120 338.330 166.290 338.500 ;
        RECT 166.530 338.470 167.350 338.500 ;
        RECT 168.590 338.470 168.770 338.530 ;
        RECT 166.530 338.330 167.640 338.470 ;
        RECT 0.480 332.140 1.940 332.180 ;
        RECT 0.480 331.970 1.950 332.140 ;
        RECT 0.480 331.930 1.940 331.970 ;
        RECT 2.180 325.550 2.690 338.160 ;
        RECT 3.050 337.370 9.030 337.600 ;
        RECT 3.140 326.310 8.790 337.370 ;
        RECT 9.200 327.800 9.710 338.160 ;
        RECT 139.040 337.810 139.210 337.880 ;
        RECT 138.970 337.780 139.290 337.810 ;
        RECT 138.960 337.590 139.290 337.780 ;
        RECT 138.970 337.550 139.290 337.590 ;
        RECT 139.040 335.040 139.210 337.550 ;
        RECT 139.590 337.140 139.760 337.880 ;
        RECT 140.140 337.820 140.310 337.880 ;
        RECT 140.070 337.790 140.390 337.820 ;
        RECT 140.060 337.600 140.390 337.790 ;
        RECT 140.070 337.560 140.390 337.600 ;
        RECT 139.520 337.110 139.840 337.140 ;
        RECT 139.510 336.920 139.840 337.110 ;
        RECT 139.520 336.880 139.840 336.920 ;
        RECT 139.590 335.770 139.760 336.880 ;
        RECT 139.520 335.740 139.840 335.770 ;
        RECT 139.510 335.550 139.840 335.740 ;
        RECT 139.520 335.510 139.840 335.550 ;
        RECT 138.970 335.010 139.290 335.040 ;
        RECT 138.960 334.820 139.290 335.010 ;
        RECT 138.970 334.780 139.290 334.820 ;
        RECT 139.040 333.700 139.210 334.780 ;
        RECT 138.960 333.670 139.280 333.700 ;
        RECT 138.950 333.480 139.280 333.670 ;
        RECT 138.960 333.440 139.280 333.480 ;
        RECT 139.040 332.700 139.210 333.440 ;
        RECT 139.590 333.000 139.760 335.510 ;
        RECT 140.140 335.040 140.310 337.560 ;
        RECT 140.690 337.140 140.860 337.880 ;
        RECT 141.240 337.820 141.410 337.880 ;
        RECT 141.160 337.790 141.480 337.820 ;
        RECT 141.150 337.600 141.480 337.790 ;
        RECT 141.160 337.560 141.480 337.600 ;
        RECT 140.620 337.110 140.940 337.140 ;
        RECT 140.610 336.920 140.940 337.110 ;
        RECT 140.620 336.880 140.940 336.920 ;
        RECT 140.690 335.770 140.860 336.880 ;
        RECT 140.620 335.740 140.940 335.770 ;
        RECT 140.610 335.550 140.940 335.740 ;
        RECT 140.620 335.510 140.940 335.550 ;
        RECT 140.070 335.010 140.390 335.040 ;
        RECT 140.060 334.820 140.390 335.010 ;
        RECT 140.070 334.780 140.390 334.820 ;
        RECT 140.140 333.690 140.310 334.780 ;
        RECT 140.070 333.660 140.390 333.690 ;
        RECT 140.060 333.470 140.390 333.660 ;
        RECT 140.070 333.430 140.390 333.470 ;
        RECT 139.520 332.970 139.840 333.000 ;
        RECT 139.510 332.780 139.840 332.970 ;
        RECT 139.520 332.740 139.840 332.780 ;
        RECT 139.590 332.700 139.760 332.740 ;
        RECT 140.140 332.700 140.310 333.430 ;
        RECT 140.690 332.990 140.860 335.510 ;
        RECT 141.240 335.040 141.410 337.560 ;
        RECT 141.790 337.140 141.960 337.880 ;
        RECT 142.200 337.600 142.710 338.280 ;
        RECT 165.520 338.230 165.870 338.330 ;
        RECT 167.180 338.300 167.640 338.330 ;
        RECT 168.090 338.300 168.770 338.470 ;
        RECT 169.710 338.450 170.040 338.620 ;
        RECT 171.510 338.430 171.690 338.890 ;
        RECT 183.410 338.580 183.580 338.930 ;
        RECT 193.160 338.880 193.490 339.070 ;
        RECT 204.750 338.910 205.410 339.170 ;
        RECT 205.580 339.000 205.910 339.170 ;
        RECT 206.130 339.000 206.470 339.170 ;
        RECT 193.160 338.850 193.480 338.880 ;
        RECT 168.130 338.280 168.770 338.300 ;
        RECT 168.590 338.270 168.770 338.280 ;
        RECT 170.370 338.270 170.970 338.420 ;
        RECT 168.590 338.250 170.970 338.270 ;
        RECT 171.430 338.260 171.760 338.430 ;
        RECT 183.350 338.410 183.580 338.580 ;
        RECT 183.750 338.680 183.940 338.720 ;
        RECT 183.750 338.510 184.310 338.680 ;
        RECT 184.770 338.510 187.520 338.680 ;
        RECT 183.750 338.490 183.940 338.510 ;
        RECT 183.410 338.370 183.580 338.410 ;
        RECT 186.750 338.330 187.080 338.510 ;
        RECT 168.590 338.100 170.820 338.250 ;
        RECT 163.520 337.760 163.690 337.810 ;
        RECT 183.480 337.770 183.650 338.190 ;
        RECT 184.290 338.060 184.530 338.100 ;
        RECT 187.070 338.060 187.240 338.070 ;
        RECT 183.960 337.890 184.530 338.060 ;
        RECT 184.770 337.890 186.110 338.060 ;
        RECT 186.560 337.890 187.520 338.060 ;
        RECT 184.290 337.860 184.530 337.890 ;
        RECT 188.050 337.820 188.220 338.750 ;
        RECT 188.450 337.770 188.620 338.620 ;
        RECT 193.210 338.260 193.390 338.850 ;
        RECT 205.070 338.660 205.410 338.910 ;
        RECT 205.660 338.830 205.830 339.000 ;
        RECT 206.220 338.830 206.390 339.000 ;
        RECT 205.580 338.660 205.910 338.830 ;
        RECT 206.130 338.660 206.470 338.830 ;
        RECT 204.600 338.450 204.920 338.490 ;
        RECT 204.600 338.430 204.930 338.450 ;
        RECT 206.220 338.430 206.390 338.660 ;
        RECT 206.790 338.580 207.300 339.250 ;
        RECT 204.600 338.260 206.390 338.430 ;
        RECT 193.210 338.220 193.530 338.260 ;
        RECT 204.600 338.230 204.920 338.260 ;
        RECT 193.210 338.030 193.540 338.220 ;
        RECT 193.210 338.000 193.530 338.030 ;
        RECT 363.700 337.950 364.210 350.850 ;
        RECT 364.610 349.960 368.070 350.400 ;
        RECT 364.610 349.860 370.000 349.960 ;
        RECT 364.720 349.790 370.000 349.860 ;
        RECT 364.720 338.880 364.890 349.790 ;
        RECT 365.270 349.380 369.500 349.400 ;
        RECT 365.190 339.270 369.520 349.380 ;
        RECT 369.290 339.220 369.460 339.270 ;
        RECT 369.830 338.880 370.000 349.790 ;
        RECT 364.720 338.710 370.000 338.880 ;
        RECT 364.720 338.700 364.960 338.710 ;
        RECT 370.720 337.950 371.230 350.860 ;
        RECT 142.200 337.530 142.720 337.600 ;
        RECT 163.490 337.540 163.710 337.760 ;
        RECT 142.210 337.270 142.720 337.530 ;
        RECT 163.520 337.480 163.690 337.540 ;
        RECT 164.040 337.400 164.370 337.580 ;
        RECT 167.180 337.570 167.350 337.620 ;
        RECT 164.620 337.400 166.780 337.570 ;
        RECT 167.020 337.400 167.350 337.570 ;
        RECT 167.640 337.430 167.850 337.760 ;
        RECT 141.720 337.110 142.040 337.140 ;
        RECT 141.710 336.920 142.040 337.110 ;
        RECT 141.720 336.880 142.040 336.920 ;
        RECT 141.790 335.770 141.960 336.880 ;
        RECT 142.500 335.890 142.670 337.080 ;
        RECT 164.070 336.960 164.340 337.400 ;
        RECT 165.550 337.140 165.880 337.400 ;
        RECT 167.090 337.260 167.350 337.400 ;
        RECT 168.090 337.260 168.270 337.700 ;
        RECT 168.820 337.490 170.180 337.600 ;
        RECT 168.820 337.430 170.260 337.490 ;
        RECT 169.620 337.420 170.260 337.430 ;
        RECT 164.110 336.950 164.340 336.960 ;
        RECT 167.090 337.090 168.270 337.260 ;
        RECT 169.790 337.320 170.260 337.420 ;
        RECT 170.730 337.340 171.690 337.510 ;
        RECT 167.090 336.950 167.350 337.090 ;
        RECT 169.790 337.070 170.040 337.320 ;
        RECT 164.110 336.780 164.870 336.950 ;
        RECT 165.120 336.780 166.290 336.950 ;
        RECT 166.530 336.920 167.350 336.950 ;
        RECT 168.590 336.920 168.770 336.980 ;
        RECT 166.530 336.780 167.640 336.920 ;
        RECT 165.520 336.680 165.870 336.780 ;
        RECT 167.180 336.750 167.640 336.780 ;
        RECT 168.090 336.750 168.770 336.920 ;
        RECT 169.710 336.900 170.040 337.070 ;
        RECT 171.510 336.880 171.690 337.340 ;
        RECT 363.700 337.440 371.230 337.950 ;
        RECT 371.440 337.890 372.910 338.140 ;
        RECT 168.130 336.730 168.770 336.750 ;
        RECT 168.590 336.720 168.770 336.730 ;
        RECT 170.370 336.720 170.970 336.870 ;
        RECT 168.590 336.700 170.970 336.720 ;
        RECT 171.430 336.710 171.760 336.880 ;
        RECT 168.590 336.550 170.820 336.700 ;
        RECT 141.720 335.740 142.040 335.770 ;
        RECT 141.710 335.550 142.040 335.740 ;
        RECT 141.720 335.510 142.040 335.550 ;
        RECT 141.160 335.010 141.480 335.040 ;
        RECT 141.150 334.820 141.480 335.010 ;
        RECT 141.160 334.780 141.480 334.820 ;
        RECT 141.240 333.670 141.410 334.780 ;
        RECT 141.160 333.640 141.480 333.670 ;
        RECT 141.150 333.450 141.480 333.640 ;
        RECT 141.160 333.410 141.480 333.450 ;
        RECT 140.620 332.960 140.940 332.990 ;
        RECT 140.610 332.770 140.940 332.960 ;
        RECT 140.620 332.730 140.940 332.770 ;
        RECT 140.690 332.700 140.860 332.730 ;
        RECT 141.240 332.700 141.410 333.410 ;
        RECT 141.790 332.990 141.960 335.510 ;
        RECT 148.830 333.580 149.590 334.000 ;
        RECT 141.710 332.960 142.030 332.990 ;
        RECT 141.700 332.770 142.030 332.960 ;
        RECT 148.850 332.790 149.590 333.580 ;
        RECT 141.710 332.730 142.030 332.770 ;
        RECT 141.790 332.700 141.960 332.730 ;
        RECT 181.120 331.850 181.290 331.880 ;
        RECT 138.260 330.220 138.580 330.250 ;
        RECT 139.360 330.230 139.680 330.260 ;
        RECT 140.450 330.230 140.770 330.260 ;
        RECT 138.250 330.030 138.580 330.220 ;
        RECT 139.350 330.040 139.680 330.230 ;
        RECT 140.440 330.190 140.770 330.230 ;
        RECT 141.490 330.190 142.000 330.720 ;
        RECT 138.260 329.990 138.580 330.030 ;
        RECT 139.360 330.000 139.680 330.040 ;
        RECT 139.790 329.580 139.960 330.190 ;
        RECT 140.340 330.000 140.770 330.190 ;
        RECT 138.810 329.550 139.130 329.580 ;
        RECT 138.800 329.360 139.130 329.550 ;
        RECT 138.810 329.320 139.130 329.360 ;
        RECT 139.790 329.320 140.230 329.580 ;
        RECT 139.790 328.210 139.960 329.320 ;
        RECT 138.810 328.180 139.130 328.210 ;
        RECT 138.800 327.990 139.130 328.180 ;
        RECT 138.810 327.950 139.130 327.990 ;
        RECT 139.790 327.950 140.230 328.210 ;
        RECT 138.330 327.910 138.490 327.920 ;
        RECT 138.880 327.910 139.040 327.920 ;
        RECT 139.430 327.910 139.590 327.920 ;
        RECT 9.190 327.780 9.710 327.800 ;
        RECT 3.140 326.300 8.850 326.310 ;
        RECT 3.060 326.130 8.850 326.300 ;
        RECT 3.150 326.120 8.850 326.130 ;
        RECT 8.620 326.050 8.790 326.120 ;
        RECT 9.190 326.000 9.720 327.780 ;
        RECT 138.320 327.560 138.490 327.910 ;
        RECT 138.870 327.580 139.040 327.910 ;
        RECT 139.420 327.580 139.590 327.910 ;
        RECT 139.790 327.690 139.960 327.950 ;
        RECT 139.980 327.910 140.140 327.920 ;
        RECT 138.330 327.540 138.490 327.560 ;
        RECT 138.880 327.540 139.040 327.580 ;
        RECT 139.430 327.540 139.590 327.580 ;
        RECT 139.970 327.510 140.140 327.910 ;
        RECT 140.340 327.690 140.510 330.000 ;
        RECT 140.890 329.580 141.060 330.190 ;
        RECT 141.440 329.710 142.160 330.190 ;
        RECT 140.890 329.320 141.330 329.580 ;
        RECT 140.890 328.210 141.060 329.320 ;
        RECT 140.890 327.950 141.330 328.210 ;
        RECT 140.530 327.910 140.690 327.920 ;
        RECT 140.520 327.580 140.690 327.910 ;
        RECT 140.890 327.690 141.060 327.950 ;
        RECT 141.080 327.910 141.240 327.920 ;
        RECT 140.530 327.540 140.690 327.580 ;
        RECT 141.070 327.570 141.240 327.910 ;
        RECT 141.440 327.690 141.610 329.710 ;
        RECT 141.990 327.690 142.160 329.710 ;
        RECT 142.540 327.690 142.710 330.180 ;
        RECT 171.310 329.360 171.480 331.850 ;
        RECT 171.860 329.350 172.030 331.850 ;
        RECT 172.410 329.350 172.580 331.850 ;
        RECT 172.960 331.540 173.130 331.850 ;
        RECT 172.700 331.280 173.130 331.540 ;
        RECT 172.960 329.350 173.130 331.280 ;
        RECT 173.510 330.860 173.680 331.850 ;
        RECT 174.060 331.540 174.230 331.850 ;
        RECT 173.790 331.280 174.230 331.540 ;
        RECT 173.250 330.600 173.680 330.860 ;
        RECT 173.510 329.490 173.680 330.600 ;
        RECT 173.250 329.350 173.680 329.490 ;
        RECT 174.060 329.350 174.230 331.280 ;
        RECT 174.890 331.490 175.210 331.530 ;
        RECT 174.890 331.300 175.220 331.490 ;
        RECT 174.890 331.270 175.210 331.300 ;
        RECT 176.070 330.900 176.240 331.660 ;
        RECT 176.460 330.900 176.630 331.660 ;
        RECT 178.470 331.540 178.640 331.850 ;
        RECT 177.490 331.490 177.810 331.530 ;
        RECT 177.480 331.300 177.810 331.490 ;
        RECT 177.490 331.270 177.810 331.300 ;
        RECT 178.470 331.280 178.910 331.540 ;
        RECT 174.340 330.800 174.660 330.840 ;
        RECT 174.340 330.610 174.670 330.800 ;
        RECT 175.450 330.790 175.770 330.830 ;
        RECT 176.930 330.790 177.250 330.830 ;
        RECT 178.040 330.800 178.360 330.840 ;
        RECT 174.340 330.580 174.660 330.610 ;
        RECT 175.450 330.600 175.780 330.790 ;
        RECT 176.920 330.600 177.250 330.790 ;
        RECT 178.030 330.610 178.360 330.800 ;
        RECT 175.450 330.570 175.770 330.600 ;
        RECT 176.930 330.570 177.250 330.600 ;
        RECT 178.040 330.580 178.360 330.610 ;
        RECT 174.340 329.450 174.660 329.490 ;
        RECT 175.440 329.450 175.760 329.490 ;
        RECT 176.940 329.450 177.260 329.490 ;
        RECT 178.040 329.450 178.360 329.490 ;
        RECT 173.250 329.260 173.580 329.350 ;
        RECT 174.340 329.260 174.670 329.450 ;
        RECT 175.440 329.260 175.770 329.450 ;
        RECT 176.930 329.260 177.260 329.450 ;
        RECT 178.030 329.260 178.360 329.450 ;
        RECT 178.470 329.350 178.640 331.280 ;
        RECT 179.020 330.860 179.190 331.850 ;
        RECT 179.570 331.540 179.740 331.850 ;
        RECT 179.570 331.280 180.000 331.540 ;
        RECT 179.020 330.600 179.450 330.860 ;
        RECT 179.020 329.490 179.190 330.600 ;
        RECT 179.020 329.350 179.450 329.490 ;
        RECT 179.570 329.350 179.740 331.280 ;
        RECT 180.120 329.350 180.290 331.850 ;
        RECT 180.670 329.350 180.840 331.850 ;
        RECT 181.120 329.390 181.390 331.850 ;
        RECT 181.220 329.360 181.390 329.390 ;
        RECT 181.670 329.380 181.840 331.880 ;
        RECT 182.220 329.380 182.390 331.880 ;
        RECT 182.770 331.570 182.940 331.880 ;
        RECT 182.510 331.310 182.940 331.570 ;
        RECT 182.770 329.380 182.940 331.310 ;
        RECT 183.320 330.890 183.490 331.880 ;
        RECT 183.870 331.570 184.040 331.880 ;
        RECT 183.600 331.310 184.040 331.570 ;
        RECT 183.060 330.630 183.490 330.890 ;
        RECT 183.320 329.520 183.490 330.630 ;
        RECT 183.060 329.380 183.490 329.520 ;
        RECT 183.870 329.380 184.040 331.310 ;
        RECT 184.700 331.520 185.020 331.560 ;
        RECT 184.700 331.330 185.030 331.520 ;
        RECT 184.700 331.300 185.020 331.330 ;
        RECT 185.880 330.930 186.050 331.690 ;
        RECT 186.270 330.930 186.440 331.690 ;
        RECT 188.280 331.570 188.450 331.880 ;
        RECT 187.300 331.520 187.620 331.560 ;
        RECT 187.290 331.330 187.620 331.520 ;
        RECT 187.300 331.300 187.620 331.330 ;
        RECT 188.280 331.310 188.720 331.570 ;
        RECT 184.150 330.830 184.470 330.870 ;
        RECT 184.150 330.640 184.480 330.830 ;
        RECT 185.260 330.820 185.580 330.860 ;
        RECT 186.740 330.820 187.060 330.860 ;
        RECT 187.850 330.830 188.170 330.870 ;
        RECT 184.150 330.610 184.470 330.640 ;
        RECT 185.260 330.630 185.590 330.820 ;
        RECT 186.730 330.630 187.060 330.820 ;
        RECT 187.840 330.640 188.170 330.830 ;
        RECT 185.260 330.600 185.580 330.630 ;
        RECT 186.740 330.600 187.060 330.630 ;
        RECT 187.850 330.610 188.170 330.640 ;
        RECT 184.150 329.480 184.470 329.520 ;
        RECT 185.250 329.480 185.570 329.520 ;
        RECT 186.750 329.480 187.070 329.520 ;
        RECT 187.850 329.480 188.170 329.520 ;
        RECT 179.120 329.260 179.450 329.350 ;
        RECT 183.060 329.290 183.390 329.380 ;
        RECT 184.150 329.290 184.480 329.480 ;
        RECT 185.250 329.290 185.580 329.480 ;
        RECT 186.740 329.290 187.070 329.480 ;
        RECT 187.840 329.290 188.170 329.480 ;
        RECT 188.280 329.380 188.450 331.310 ;
        RECT 188.830 330.890 189.000 331.880 ;
        RECT 189.380 331.570 189.550 331.880 ;
        RECT 189.380 331.310 189.810 331.570 ;
        RECT 188.830 330.630 189.260 330.890 ;
        RECT 188.830 329.520 189.000 330.630 ;
        RECT 188.830 329.380 189.260 329.520 ;
        RECT 189.380 329.380 189.550 331.310 ;
        RECT 189.930 329.380 190.100 331.880 ;
        RECT 190.480 329.380 190.650 331.880 ;
        RECT 191.030 329.390 191.200 331.880 ;
        RECT 193.310 330.840 193.480 331.580 ;
        RECT 193.860 331.540 194.030 331.580 ;
        RECT 193.790 331.500 194.110 331.540 ;
        RECT 193.780 331.310 194.110 331.500 ;
        RECT 193.790 331.280 194.110 331.310 ;
        RECT 193.230 330.800 193.550 330.840 ;
        RECT 193.220 330.610 193.550 330.800 ;
        RECT 193.230 330.580 193.550 330.610 ;
        RECT 193.310 329.500 193.480 330.580 ;
        RECT 193.240 329.460 193.560 329.500 ;
        RECT 188.930 329.290 189.260 329.380 ;
        RECT 183.060 329.260 183.380 329.290 ;
        RECT 184.150 329.260 184.470 329.290 ;
        RECT 185.250 329.260 185.570 329.290 ;
        RECT 186.750 329.260 187.070 329.290 ;
        RECT 187.850 329.260 188.170 329.290 ;
        RECT 188.940 329.260 189.260 329.290 ;
        RECT 193.230 329.270 193.560 329.460 ;
        RECT 173.250 329.230 173.570 329.260 ;
        RECT 174.340 329.230 174.660 329.260 ;
        RECT 175.440 329.230 175.760 329.260 ;
        RECT 176.940 329.230 177.260 329.260 ;
        RECT 178.040 329.230 178.360 329.260 ;
        RECT 179.130 329.230 179.450 329.260 ;
        RECT 193.240 329.240 193.560 329.270 ;
        RECT 172.780 329.140 172.940 329.170 ;
        RECT 141.080 327.540 141.240 327.570 ;
        RECT 138.260 327.450 138.580 327.480 ;
        RECT 139.360 327.450 139.680 327.480 ;
        RECT 140.450 327.450 140.770 327.480 ;
        RECT 138.250 327.260 138.580 327.450 ;
        RECT 139.350 327.260 139.680 327.450 ;
        RECT 140.440 327.360 140.770 327.450 ;
        RECT 138.260 327.220 138.580 327.260 ;
        RECT 139.360 327.220 139.680 327.260 ;
        RECT 138.250 326.110 138.570 326.140 ;
        RECT 9.200 325.980 9.720 326.000 ;
        RECT 2.180 325.260 4.620 325.550 ;
        RECT 9.200 325.470 9.710 325.980 ;
        RECT 138.240 325.920 138.570 326.110 ;
        RECT 139.360 326.100 139.680 326.130 ;
        RECT 138.250 325.880 138.570 325.920 ;
        RECT 139.350 325.910 139.680 326.100 ;
        RECT 139.360 325.870 139.680 325.910 ;
        RECT 9.200 325.260 9.730 325.470 ;
        RECT 2.180 324.780 9.730 325.260 ;
        RECT 137.780 325.050 137.950 325.810 ;
        RECT 138.810 325.410 139.130 325.440 ;
        RECT 138.800 325.220 139.130 325.410 ;
        RECT 138.810 325.180 139.130 325.220 ;
        RECT 139.790 325.430 139.960 327.360 ;
        RECT 140.340 327.220 140.770 327.360 ;
        RECT 140.340 326.110 140.510 327.220 ;
        RECT 140.340 325.850 140.770 326.110 ;
        RECT 139.790 325.170 140.230 325.430 ;
        RECT 139.790 324.860 139.960 325.170 ;
        RECT 140.340 324.860 140.510 325.850 ;
        RECT 140.890 325.430 141.060 327.360 ;
        RECT 140.890 325.170 141.320 325.430 ;
        RECT 140.890 324.860 141.060 325.170 ;
        RECT 141.440 324.860 141.610 327.360 ;
        RECT 141.990 324.860 142.160 327.360 ;
        RECT 142.540 324.860 142.710 327.350 ;
        RECT 171.310 326.530 171.480 329.020 ;
        RECT 171.860 327.000 172.030 329.020 ;
        RECT 172.410 327.000 172.580 329.020 ;
        RECT 172.780 328.800 172.950 329.140 ;
        RECT 173.330 329.130 173.490 329.170 ;
        RECT 172.780 328.790 172.940 328.800 ;
        RECT 172.960 328.760 173.130 329.020 ;
        RECT 173.330 328.800 173.500 329.130 ;
        RECT 173.330 328.790 173.490 328.800 ;
        RECT 172.690 328.500 173.130 328.760 ;
        RECT 172.960 327.390 173.130 328.500 ;
        RECT 172.690 327.130 173.130 327.390 ;
        RECT 171.860 326.520 172.580 327.000 ;
        RECT 172.960 326.520 173.130 327.130 ;
        RECT 173.510 326.710 173.680 329.020 ;
        RECT 173.880 328.800 174.050 329.200 ;
        RECT 174.430 329.130 174.590 329.170 ;
        RECT 174.980 329.130 175.140 329.170 ;
        RECT 175.530 329.150 175.690 329.170 ;
        RECT 177.010 329.150 177.170 329.170 ;
        RECT 173.880 328.790 174.040 328.800 ;
        RECT 174.060 328.760 174.230 329.020 ;
        RECT 174.430 328.800 174.600 329.130 ;
        RECT 174.980 328.800 175.150 329.130 ;
        RECT 175.530 328.800 175.700 329.150 ;
        RECT 177.000 328.800 177.170 329.150 ;
        RECT 177.560 329.130 177.720 329.170 ;
        RECT 178.110 329.130 178.270 329.170 ;
        RECT 177.550 328.800 177.720 329.130 ;
        RECT 178.100 328.800 178.270 329.130 ;
        RECT 174.430 328.790 174.590 328.800 ;
        RECT 174.980 328.790 175.140 328.800 ;
        RECT 175.530 328.790 175.690 328.800 ;
        RECT 177.010 328.790 177.170 328.800 ;
        RECT 177.560 328.790 177.720 328.800 ;
        RECT 178.110 328.790 178.270 328.800 ;
        RECT 178.470 328.760 178.640 329.020 ;
        RECT 178.650 328.800 178.820 329.200 ;
        RECT 182.590 329.170 182.750 329.200 ;
        RECT 179.210 329.130 179.370 329.170 ;
        RECT 179.760 329.140 179.920 329.170 ;
        RECT 178.660 328.790 178.820 328.800 ;
        RECT 173.790 328.500 174.230 328.760 ;
        RECT 174.890 328.720 175.210 328.760 ;
        RECT 177.490 328.720 177.810 328.760 ;
        RECT 174.890 328.530 175.220 328.720 ;
        RECT 177.480 328.530 177.810 328.720 ;
        RECT 174.890 328.500 175.210 328.530 ;
        RECT 177.490 328.500 177.810 328.530 ;
        RECT 178.470 328.500 178.910 328.760 ;
        RECT 174.060 327.390 174.230 328.500 ;
        RECT 178.470 327.390 178.640 328.500 ;
        RECT 173.790 327.130 174.230 327.390 ;
        RECT 174.890 327.350 175.210 327.390 ;
        RECT 177.490 327.350 177.810 327.390 ;
        RECT 174.890 327.160 175.220 327.350 ;
        RECT 177.480 327.160 177.810 327.350 ;
        RECT 174.890 327.130 175.210 327.160 ;
        RECT 177.490 327.130 177.810 327.160 ;
        RECT 178.470 327.130 178.910 327.390 ;
        RECT 173.250 326.520 173.680 326.710 ;
        RECT 174.060 326.520 174.230 327.130 ;
        RECT 174.340 326.670 174.660 326.710 ;
        RECT 175.440 326.680 175.760 326.720 ;
        RECT 176.940 326.680 177.260 326.720 ;
        RECT 172.020 325.990 172.530 326.520 ;
        RECT 173.250 326.480 173.580 326.520 ;
        RECT 174.340 326.480 174.670 326.670 ;
        RECT 175.440 326.490 175.770 326.680 ;
        RECT 176.930 326.490 177.260 326.680 ;
        RECT 178.040 326.670 178.360 326.710 ;
        RECT 173.250 326.450 173.570 326.480 ;
        RECT 174.340 326.450 174.660 326.480 ;
        RECT 175.440 326.460 175.760 326.490 ;
        RECT 176.940 326.460 177.260 326.490 ;
        RECT 178.030 326.480 178.360 326.670 ;
        RECT 178.470 326.520 178.640 327.130 ;
        RECT 179.020 326.710 179.190 329.020 ;
        RECT 179.200 328.800 179.370 329.130 ;
        RECT 179.210 328.790 179.370 328.800 ;
        RECT 179.570 328.760 179.740 329.020 ;
        RECT 179.750 328.800 179.920 329.140 ;
        RECT 181.120 329.020 181.290 329.050 ;
        RECT 179.760 328.790 179.920 328.800 ;
        RECT 179.570 328.500 180.010 328.760 ;
        RECT 179.570 327.390 179.740 328.500 ;
        RECT 179.570 327.130 180.010 327.390 ;
        RECT 179.020 326.520 179.450 326.710 ;
        RECT 179.570 326.520 179.740 327.130 ;
        RECT 180.120 327.000 180.290 329.020 ;
        RECT 180.670 327.000 180.840 329.020 ;
        RECT 180.120 326.520 180.840 327.000 ;
        RECT 181.120 326.560 181.390 329.020 ;
        RECT 181.220 326.530 181.390 326.560 ;
        RECT 181.670 327.030 181.840 329.050 ;
        RECT 182.220 327.030 182.390 329.050 ;
        RECT 182.590 328.830 182.760 329.170 ;
        RECT 183.140 329.160 183.300 329.200 ;
        RECT 182.590 328.820 182.750 328.830 ;
        RECT 182.770 328.790 182.940 329.050 ;
        RECT 183.140 328.830 183.310 329.160 ;
        RECT 183.140 328.820 183.300 328.830 ;
        RECT 182.500 328.530 182.940 328.790 ;
        RECT 182.770 327.420 182.940 328.530 ;
        RECT 182.500 327.160 182.940 327.420 ;
        RECT 181.670 326.550 182.390 327.030 ;
        RECT 182.770 326.550 182.940 327.160 ;
        RECT 183.320 326.740 183.490 329.050 ;
        RECT 183.690 328.830 183.860 329.230 ;
        RECT 184.240 329.160 184.400 329.200 ;
        RECT 184.790 329.160 184.950 329.200 ;
        RECT 185.340 329.180 185.500 329.200 ;
        RECT 186.820 329.180 186.980 329.200 ;
        RECT 183.690 328.820 183.850 328.830 ;
        RECT 183.870 328.790 184.040 329.050 ;
        RECT 184.240 328.830 184.410 329.160 ;
        RECT 184.790 328.830 184.960 329.160 ;
        RECT 185.340 328.830 185.510 329.180 ;
        RECT 186.810 328.830 186.980 329.180 ;
        RECT 187.370 329.160 187.530 329.200 ;
        RECT 187.920 329.160 188.080 329.200 ;
        RECT 187.360 328.830 187.530 329.160 ;
        RECT 187.910 328.830 188.080 329.160 ;
        RECT 184.240 328.820 184.400 328.830 ;
        RECT 184.790 328.820 184.950 328.830 ;
        RECT 185.340 328.820 185.500 328.830 ;
        RECT 186.820 328.820 186.980 328.830 ;
        RECT 187.370 328.820 187.530 328.830 ;
        RECT 187.920 328.820 188.080 328.830 ;
        RECT 188.280 328.790 188.450 329.050 ;
        RECT 188.460 328.830 188.630 329.230 ;
        RECT 189.020 329.160 189.180 329.200 ;
        RECT 189.570 329.170 189.730 329.200 ;
        RECT 188.470 328.820 188.630 328.830 ;
        RECT 183.600 328.530 184.040 328.790 ;
        RECT 184.700 328.750 185.020 328.790 ;
        RECT 187.300 328.750 187.620 328.790 ;
        RECT 184.700 328.560 185.030 328.750 ;
        RECT 187.290 328.560 187.620 328.750 ;
        RECT 184.700 328.530 185.020 328.560 ;
        RECT 187.300 328.530 187.620 328.560 ;
        RECT 188.280 328.530 188.720 328.790 ;
        RECT 183.870 327.420 184.040 328.530 ;
        RECT 188.280 327.420 188.450 328.530 ;
        RECT 183.600 327.160 184.040 327.420 ;
        RECT 184.700 327.380 185.020 327.420 ;
        RECT 187.300 327.380 187.620 327.420 ;
        RECT 184.700 327.190 185.030 327.380 ;
        RECT 187.290 327.190 187.620 327.380 ;
        RECT 184.700 327.160 185.020 327.190 ;
        RECT 187.300 327.160 187.620 327.190 ;
        RECT 188.280 327.160 188.720 327.420 ;
        RECT 183.060 326.550 183.490 326.740 ;
        RECT 183.870 326.550 184.040 327.160 ;
        RECT 184.150 326.700 184.470 326.740 ;
        RECT 185.250 326.710 185.570 326.750 ;
        RECT 186.750 326.710 187.070 326.750 ;
        RECT 179.120 326.480 179.450 326.520 ;
        RECT 178.040 326.450 178.360 326.480 ;
        RECT 179.130 326.450 179.450 326.480 ;
        RECT 180.170 325.990 180.680 326.520 ;
        RECT 181.830 326.020 182.340 326.550 ;
        RECT 183.060 326.510 183.390 326.550 ;
        RECT 184.150 326.510 184.480 326.700 ;
        RECT 185.250 326.520 185.580 326.710 ;
        RECT 186.740 326.520 187.070 326.710 ;
        RECT 187.850 326.700 188.170 326.740 ;
        RECT 183.060 326.480 183.380 326.510 ;
        RECT 184.150 326.480 184.470 326.510 ;
        RECT 185.250 326.490 185.570 326.520 ;
        RECT 186.750 326.490 187.070 326.520 ;
        RECT 187.840 326.510 188.170 326.700 ;
        RECT 188.280 326.550 188.450 327.160 ;
        RECT 188.830 326.740 189.000 329.050 ;
        RECT 189.010 328.830 189.180 329.160 ;
        RECT 189.020 328.820 189.180 328.830 ;
        RECT 189.380 328.790 189.550 329.050 ;
        RECT 189.560 328.830 189.730 329.170 ;
        RECT 189.570 328.820 189.730 328.830 ;
        RECT 189.380 328.530 189.820 328.790 ;
        RECT 189.380 327.420 189.550 328.530 ;
        RECT 189.380 327.160 189.820 327.420 ;
        RECT 188.830 326.550 189.260 326.740 ;
        RECT 189.380 326.550 189.550 327.160 ;
        RECT 189.930 327.030 190.100 329.050 ;
        RECT 190.480 327.030 190.650 329.050 ;
        RECT 189.930 326.550 190.650 327.030 ;
        RECT 191.030 326.560 191.200 329.050 ;
        RECT 193.310 326.730 193.480 329.240 ;
        RECT 193.860 328.770 194.030 331.280 ;
        RECT 194.410 330.850 194.580 331.580 ;
        RECT 194.960 331.550 195.130 331.580 ;
        RECT 194.890 331.510 195.210 331.550 ;
        RECT 194.880 331.320 195.210 331.510 ;
        RECT 194.890 331.290 195.210 331.320 ;
        RECT 194.340 330.810 194.660 330.850 ;
        RECT 194.330 330.620 194.660 330.810 ;
        RECT 194.340 330.590 194.660 330.620 ;
        RECT 194.410 329.500 194.580 330.590 ;
        RECT 194.340 329.460 194.660 329.500 ;
        RECT 194.330 329.270 194.660 329.460 ;
        RECT 194.340 329.240 194.660 329.270 ;
        RECT 193.790 328.730 194.110 328.770 ;
        RECT 193.780 328.540 194.110 328.730 ;
        RECT 193.790 328.510 194.110 328.540 ;
        RECT 193.860 327.400 194.030 328.510 ;
        RECT 193.790 327.360 194.110 327.400 ;
        RECT 193.780 327.170 194.110 327.360 ;
        RECT 193.790 327.140 194.110 327.170 ;
        RECT 193.240 326.690 193.560 326.730 ;
        RECT 188.930 326.510 189.260 326.550 ;
        RECT 187.850 326.480 188.170 326.510 ;
        RECT 188.940 326.480 189.260 326.510 ;
        RECT 189.980 326.020 190.490 326.550 ;
        RECT 193.230 326.500 193.560 326.690 ;
        RECT 193.240 326.470 193.560 326.500 ;
        RECT 193.310 326.400 193.480 326.470 ;
        RECT 193.860 326.400 194.030 327.140 ;
        RECT 194.410 326.720 194.580 329.240 ;
        RECT 194.960 328.770 195.130 331.290 ;
        RECT 195.510 330.870 195.680 331.580 ;
        RECT 196.060 331.550 196.230 331.580 ;
        RECT 195.980 331.510 196.300 331.550 ;
        RECT 195.970 331.320 196.300 331.510 ;
        RECT 195.980 331.290 196.300 331.320 ;
        RECT 195.430 330.830 195.750 330.870 ;
        RECT 195.420 330.640 195.750 330.830 ;
        RECT 195.430 330.610 195.750 330.640 ;
        RECT 195.510 329.500 195.680 330.610 ;
        RECT 195.430 329.460 195.750 329.500 ;
        RECT 195.420 329.270 195.750 329.460 ;
        RECT 195.430 329.240 195.750 329.270 ;
        RECT 194.890 328.730 195.210 328.770 ;
        RECT 194.880 328.540 195.210 328.730 ;
        RECT 194.890 328.510 195.210 328.540 ;
        RECT 194.960 327.400 195.130 328.510 ;
        RECT 194.890 327.360 195.210 327.400 ;
        RECT 194.880 327.170 195.210 327.360 ;
        RECT 194.890 327.140 195.210 327.170 ;
        RECT 194.340 326.680 194.660 326.720 ;
        RECT 194.330 326.490 194.660 326.680 ;
        RECT 194.340 326.460 194.660 326.490 ;
        RECT 194.410 326.400 194.580 326.460 ;
        RECT 194.960 326.400 195.130 327.140 ;
        RECT 195.510 326.720 195.680 329.240 ;
        RECT 196.060 328.770 196.230 331.290 ;
        RECT 195.990 328.730 196.310 328.770 ;
        RECT 195.980 328.540 196.310 328.730 ;
        RECT 195.990 328.510 196.310 328.540 ;
        RECT 196.060 327.400 196.230 328.510 ;
        RECT 195.990 327.360 196.310 327.400 ;
        RECT 195.980 327.170 196.310 327.360 ;
        RECT 196.770 327.200 196.940 328.390 ;
        RECT 195.990 327.140 196.310 327.170 ;
        RECT 195.430 326.680 195.750 326.720 ;
        RECT 195.420 326.490 195.750 326.680 ;
        RECT 195.430 326.460 195.750 326.490 ;
        RECT 195.510 326.400 195.680 326.460 ;
        RECT 196.060 326.400 196.230 327.140 ;
        RECT 196.480 326.750 196.990 327.010 ;
        RECT 196.470 326.680 196.990 326.750 ;
        RECT 196.470 326.000 196.980 326.680 ;
        RECT 143.180 324.890 145.570 325.260 ;
        RECT 2.180 324.750 9.540 324.780 ;
        RECT 2.180 322.990 9.710 323.540 ;
        RECT 0.500 310.020 1.970 310.270 ;
        RECT 2.180 310.080 2.690 322.990 ;
        RECT 9.040 322.980 9.710 322.990 ;
        RECT 5.340 322.090 8.800 322.530 ;
        RECT 3.410 321.990 8.800 322.090 ;
        RECT 3.410 321.920 8.690 321.990 ;
        RECT 3.410 311.010 3.580 321.920 ;
        RECT 3.910 321.510 8.140 321.530 ;
        RECT 3.890 311.400 8.220 321.510 ;
        RECT 3.950 311.350 4.120 311.400 ;
        RECT 8.520 311.010 8.690 321.920 ;
        RECT 3.410 310.840 8.690 311.010 ;
        RECT 8.450 310.830 8.690 310.840 ;
        RECT 9.200 310.080 9.710 322.980 ;
        RECT 143.230 321.630 145.570 324.890 ;
        RECT 221.980 324.090 222.210 324.100 ;
        RECT 221.960 323.920 226.620 324.090 ;
        RECT 221.980 323.910 222.210 323.920 ;
        RECT 227.520 323.440 227.710 323.450 ;
        RECT 223.180 323.400 226.980 323.410 ;
        RECT 227.490 323.400 227.750 323.440 ;
        RECT 223.180 323.240 227.750 323.400 ;
        RECT 226.750 323.230 227.750 323.240 ;
        RECT 226.750 322.770 226.980 323.230 ;
        RECT 227.490 323.120 227.750 323.230 ;
        RECT 227.520 322.770 227.710 322.780 ;
        RECT 226.750 322.560 227.760 322.770 ;
        RECT 221.980 322.480 222.210 322.490 ;
        RECT 221.960 322.310 226.440 322.480 ;
        RECT 221.980 322.300 222.210 322.310 ;
        RECT 226.750 321.800 226.980 322.560 ;
        RECT 227.490 322.450 227.750 322.560 ;
        RECT 223.200 321.630 226.980 321.800 ;
        RECT 143.230 321.620 145.560 321.630 ;
        RECT 221.980 320.880 222.210 320.890 ;
        RECT 221.960 320.710 226.460 320.880 ;
        RECT 221.980 320.700 222.210 320.710 ;
        RECT 223.200 320.700 223.530 320.710 ;
        RECT 224.160 320.700 224.490 320.710 ;
        RECT 225.120 320.700 225.450 320.710 ;
        RECT 226.080 320.700 226.410 320.710 ;
        RECT 226.750 320.190 226.980 321.630 ;
        RECT 227.430 321.440 227.860 321.460 ;
        RECT 227.410 321.270 227.860 321.440 ;
        RECT 227.430 321.250 227.860 321.270 ;
        RECT 223.200 320.020 226.980 320.190 ;
        RECT 223.260 319.790 223.690 319.810 ;
        RECT 223.240 319.620 223.690 319.790 ;
        RECT 223.260 319.600 223.690 319.620 ;
        RECT 221.980 319.260 222.210 319.270 ;
        RECT 221.960 319.090 226.460 319.260 ;
        RECT 221.980 319.080 222.210 319.090 ;
        RECT 226.750 318.590 226.980 320.020 ;
        RECT 227.430 319.830 227.860 319.850 ;
        RECT 227.410 319.660 227.860 319.830 ;
        RECT 227.430 319.640 227.860 319.660 ;
        RECT 223.210 318.580 226.980 318.590 ;
        RECT 223.200 318.420 226.980 318.580 ;
        RECT 223.200 318.410 223.530 318.420 ;
        RECT 225.120 318.410 225.450 318.420 ;
        RECT 226.080 318.410 226.410 318.420 ;
        RECT 224.260 318.050 224.690 318.070 ;
        RECT 224.260 317.880 224.710 318.050 ;
        RECT 224.260 317.860 224.690 317.880 ;
        RECT 221.980 317.660 222.210 317.670 ;
        RECT 221.960 317.490 226.410 317.660 ;
        RECT 221.980 317.480 222.210 317.490 ;
        RECT 223.200 317.480 223.530 317.490 ;
        RECT 224.160 317.480 224.490 317.490 ;
        RECT 225.120 317.480 225.450 317.490 ;
        RECT 226.080 317.480 226.410 317.490 ;
        RECT 226.750 316.970 226.980 318.420 ;
        RECT 227.420 318.220 227.850 318.240 ;
        RECT 227.400 318.050 227.850 318.220 ;
        RECT 227.420 318.030 227.850 318.050 ;
        RECT 223.190 316.800 226.980 316.970 ;
        RECT 225.170 316.540 225.600 316.560 ;
        RECT 225.150 316.370 225.600 316.540 ;
        RECT 225.170 316.350 225.600 316.370 ;
        RECT 221.980 316.040 222.210 316.050 ;
        RECT 221.960 315.870 226.460 316.040 ;
        RECT 221.980 315.860 222.210 315.870 ;
        RECT 223.200 315.350 223.530 315.360 ;
        RECT 224.160 315.350 224.490 315.360 ;
        RECT 225.120 315.350 225.450 315.360 ;
        RECT 226.080 315.350 226.410 315.360 ;
        RECT 226.750 315.350 226.980 316.800 ;
        RECT 227.420 316.600 227.850 316.620 ;
        RECT 227.400 316.430 227.850 316.600 ;
        RECT 227.420 316.410 227.850 316.430 ;
        RECT 223.190 315.180 226.980 315.350 ;
        RECT 221.980 314.440 222.210 314.450 ;
        RECT 221.960 314.430 226.380 314.440 ;
        RECT 221.960 314.270 226.410 314.430 ;
        RECT 221.980 314.260 222.210 314.270 ;
        RECT 223.200 314.260 223.530 314.270 ;
        RECT 224.160 314.260 224.490 314.270 ;
        RECT 225.120 314.260 225.450 314.270 ;
        RECT 226.080 314.260 226.410 314.270 ;
        RECT 226.750 313.760 226.980 315.180 ;
        RECT 227.420 314.990 227.850 315.010 ;
        RECT 227.400 314.820 227.850 314.990 ;
        RECT 227.420 314.800 227.850 314.820 ;
        RECT 233.410 314.630 233.780 329.500 ;
        RECT 363.700 327.080 364.210 337.440 ;
        RECT 364.380 336.650 370.360 336.880 ;
        RECT 363.700 327.060 364.220 327.080 ;
        RECT 363.690 325.280 364.220 327.060 ;
        RECT 364.620 325.590 370.270 336.650 ;
        RECT 364.560 325.580 370.270 325.590 ;
        RECT 364.560 325.410 370.350 325.580 ;
        RECT 364.560 325.400 370.260 325.410 ;
        RECT 364.620 325.330 364.790 325.400 ;
        RECT 363.690 325.260 364.210 325.280 ;
        RECT 363.700 324.750 364.210 325.260 ;
        RECT 370.720 324.830 371.230 337.440 ;
        RECT 371.470 331.420 372.930 331.460 ;
        RECT 371.460 331.250 372.930 331.420 ;
        RECT 371.470 331.210 372.930 331.250 ;
        RECT 363.680 324.540 364.210 324.750 ;
        RECT 368.790 324.540 371.230 324.830 ;
        RECT 363.680 324.060 371.230 324.540 ;
        RECT 363.870 324.030 371.230 324.060 ;
        RECT 363.700 322.270 371.230 322.820 ;
        RECT 363.700 322.260 364.370 322.270 ;
        RECT 233.410 314.380 233.790 314.630 ;
        RECT 223.190 313.590 226.990 313.760 ;
        RECT 223.200 313.580 223.530 313.590 ;
        RECT 224.160 313.580 224.490 313.590 ;
        RECT 225.120 313.580 225.450 313.590 ;
        RECT 226.080 313.580 226.410 313.590 ;
        RECT 221.980 312.810 222.210 312.830 ;
        RECT 223.200 312.810 223.530 312.820 ;
        RECT 224.160 312.810 224.490 312.820 ;
        RECT 225.120 312.810 225.450 312.820 ;
        RECT 226.080 312.810 226.410 312.820 ;
        RECT 221.960 312.640 226.420 312.810 ;
        RECT 226.750 312.150 226.980 313.590 ;
        RECT 227.260 313.000 227.470 313.430 ;
        RECT 227.280 312.980 227.450 313.000 ;
        RECT 223.190 311.980 226.980 312.150 ;
        RECT 223.200 311.970 223.530 311.980 ;
        RECT 224.160 311.970 224.490 311.980 ;
        RECT 225.120 311.970 225.450 311.980 ;
        RECT 226.080 311.970 226.410 311.980 ;
        RECT 227.430 311.790 227.860 311.810 ;
        RECT 227.410 311.620 227.860 311.790 ;
        RECT 227.430 311.600 227.860 311.620 ;
        RECT 227.420 310.200 227.850 310.220 ;
        RECT 224.220 310.120 224.650 310.140 ;
        RECT 225.160 310.120 225.590 310.140 ;
        RECT 2.180 309.570 9.710 310.080 ;
        RECT 224.200 309.950 224.650 310.120 ;
        RECT 225.140 309.950 225.590 310.120 ;
        RECT 226.110 310.060 226.540 310.080 ;
        RECT 224.220 309.930 224.650 309.950 ;
        RECT 225.160 309.930 225.590 309.950 ;
        RECT 226.090 309.890 226.540 310.060 ;
        RECT 227.400 310.030 227.850 310.200 ;
        RECT 227.420 310.010 227.850 310.030 ;
        RECT 226.110 309.870 226.540 309.890 ;
        RECT 0.480 303.550 1.940 303.590 ;
        RECT 0.480 303.380 1.950 303.550 ;
        RECT 0.480 303.340 1.940 303.380 ;
        RECT 2.180 296.960 2.690 309.570 ;
        RECT 3.050 308.780 9.030 309.010 ;
        RECT 3.140 297.720 8.790 308.780 ;
        RECT 9.200 299.210 9.710 309.570 ;
        RECT 9.190 299.190 9.710 299.210 ;
        RECT 363.700 309.360 364.210 322.260 ;
        RECT 364.610 321.370 368.070 321.810 ;
        RECT 364.610 321.270 370.000 321.370 ;
        RECT 364.720 321.200 370.000 321.270 ;
        RECT 364.720 310.290 364.890 321.200 ;
        RECT 365.270 320.790 369.500 320.810 ;
        RECT 365.190 310.680 369.520 320.790 ;
        RECT 369.290 310.630 369.460 310.680 ;
        RECT 369.830 310.290 370.000 321.200 ;
        RECT 364.720 310.120 370.000 310.290 ;
        RECT 364.720 310.110 364.960 310.120 ;
        RECT 370.720 309.360 371.230 322.270 ;
        RECT 363.700 308.850 371.230 309.360 ;
        RECT 371.440 309.300 372.910 309.550 ;
        RECT 3.140 297.710 8.850 297.720 ;
        RECT 3.060 297.540 8.850 297.710 ;
        RECT 3.150 297.530 8.850 297.540 ;
        RECT 8.620 297.460 8.790 297.530 ;
        RECT 9.190 297.410 9.720 299.190 ;
        RECT 363.700 298.490 364.210 308.850 ;
        RECT 364.380 308.060 370.360 308.290 ;
        RECT 363.700 298.470 364.220 298.490 ;
        RECT 9.200 297.390 9.720 297.410 ;
        RECT 2.180 296.670 4.620 296.960 ;
        RECT 9.200 296.880 9.710 297.390 ;
        RECT 9.200 296.670 9.730 296.880 ;
        RECT 363.690 296.690 364.220 298.470 ;
        RECT 364.620 297.000 370.270 308.060 ;
        RECT 364.560 296.990 370.270 297.000 ;
        RECT 364.560 296.820 370.350 296.990 ;
        RECT 364.560 296.810 370.260 296.820 ;
        RECT 364.620 296.740 364.790 296.810 ;
        RECT 363.690 296.670 364.210 296.690 ;
        RECT 2.180 296.190 9.730 296.670 ;
        RECT 2.180 296.160 9.540 296.190 ;
        RECT 363.700 296.160 364.210 296.670 ;
        RECT 370.720 296.240 371.230 308.850 ;
        RECT 371.470 302.830 372.930 302.870 ;
        RECT 371.460 302.660 372.930 302.830 ;
        RECT 371.470 302.620 372.930 302.660 ;
        RECT 363.680 295.950 364.210 296.160 ;
        RECT 368.790 295.950 371.230 296.240 ;
        RECT 363.680 295.470 371.230 295.950 ;
        RECT 363.870 295.440 371.230 295.470 ;
        RECT 2.180 294.400 9.710 294.950 ;
        RECT 0.500 281.430 1.970 281.680 ;
        RECT 2.180 281.490 2.690 294.400 ;
        RECT 9.040 294.390 9.710 294.400 ;
        RECT 5.340 293.500 8.800 293.940 ;
        RECT 3.410 293.400 8.800 293.500 ;
        RECT 3.410 293.330 8.690 293.400 ;
        RECT 3.410 282.420 3.580 293.330 ;
        RECT 3.910 292.920 8.140 292.940 ;
        RECT 3.890 282.810 8.220 292.920 ;
        RECT 3.950 282.760 4.120 282.810 ;
        RECT 8.520 282.420 8.690 293.330 ;
        RECT 3.410 282.250 8.690 282.420 ;
        RECT 8.450 282.240 8.690 282.250 ;
        RECT 9.200 281.490 9.710 294.390 ;
        RECT 2.180 280.980 9.710 281.490 ;
        RECT 0.480 274.960 1.940 275.000 ;
        RECT 0.480 274.790 1.950 274.960 ;
        RECT 0.480 274.750 1.940 274.790 ;
        RECT 2.180 268.370 2.690 280.980 ;
        RECT 3.050 280.190 9.030 280.420 ;
        RECT 3.140 269.130 8.790 280.190 ;
        RECT 9.200 270.620 9.710 280.980 ;
        RECT 9.190 270.600 9.710 270.620 ;
        RECT 363.700 293.680 371.230 294.230 ;
        RECT 363.700 293.670 364.370 293.680 ;
        RECT 363.700 280.770 364.210 293.670 ;
        RECT 364.610 292.780 368.070 293.220 ;
        RECT 364.610 292.680 370.000 292.780 ;
        RECT 364.720 292.610 370.000 292.680 ;
        RECT 364.720 281.700 364.890 292.610 ;
        RECT 365.270 292.200 369.500 292.220 ;
        RECT 365.190 282.090 369.520 292.200 ;
        RECT 369.290 282.040 369.460 282.090 ;
        RECT 369.830 281.700 370.000 292.610 ;
        RECT 364.720 281.530 370.000 281.700 ;
        RECT 364.720 281.520 364.960 281.530 ;
        RECT 370.720 280.770 371.230 293.680 ;
        RECT 363.700 280.260 371.230 280.770 ;
        RECT 371.440 280.710 372.910 280.960 ;
        RECT 3.140 269.120 8.850 269.130 ;
        RECT 3.060 268.950 8.850 269.120 ;
        RECT 3.150 268.940 8.850 268.950 ;
        RECT 8.620 268.870 8.790 268.940 ;
        RECT 9.190 268.820 9.720 270.600 ;
        RECT 363.700 269.900 364.210 280.260 ;
        RECT 364.380 279.470 370.360 279.700 ;
        RECT 363.700 269.880 364.220 269.900 ;
        RECT 9.200 268.800 9.720 268.820 ;
        RECT 2.180 268.080 4.620 268.370 ;
        RECT 9.200 268.290 9.710 268.800 ;
        RECT 9.200 268.080 9.730 268.290 ;
        RECT 363.690 268.100 364.220 269.880 ;
        RECT 364.620 268.410 370.270 279.470 ;
        RECT 364.560 268.400 370.270 268.410 ;
        RECT 364.560 268.230 370.350 268.400 ;
        RECT 364.560 268.220 370.260 268.230 ;
        RECT 364.620 268.150 364.790 268.220 ;
        RECT 363.690 268.080 364.210 268.100 ;
        RECT 2.180 267.600 9.730 268.080 ;
        RECT 2.180 267.570 9.540 267.600 ;
        RECT 363.700 267.570 364.210 268.080 ;
        RECT 370.720 267.650 371.230 280.260 ;
        RECT 371.470 274.240 372.930 274.280 ;
        RECT 371.460 274.070 372.930 274.240 ;
        RECT 371.470 274.030 372.930 274.070 ;
        RECT 363.680 267.360 364.210 267.570 ;
        RECT 368.790 267.360 371.230 267.650 ;
        RECT 363.680 266.880 371.230 267.360 ;
        RECT 363.870 266.850 371.230 266.880 ;
        RECT 2.180 265.810 9.710 266.360 ;
        RECT 0.500 252.840 1.970 253.090 ;
        RECT 2.180 252.900 2.690 265.810 ;
        RECT 9.040 265.800 9.710 265.810 ;
        RECT 5.340 264.910 8.800 265.350 ;
        RECT 3.410 264.810 8.800 264.910 ;
        RECT 3.410 264.740 8.690 264.810 ;
        RECT 3.410 253.830 3.580 264.740 ;
        RECT 3.910 264.330 8.140 264.350 ;
        RECT 3.890 254.220 8.220 264.330 ;
        RECT 3.950 254.170 4.120 254.220 ;
        RECT 8.520 253.830 8.690 264.740 ;
        RECT 3.410 253.660 8.690 253.830 ;
        RECT 8.450 253.650 8.690 253.660 ;
        RECT 9.200 252.900 9.710 265.800 ;
        RECT 2.180 252.390 9.710 252.900 ;
        RECT 0.480 246.370 1.940 246.410 ;
        RECT 0.480 246.200 1.950 246.370 ;
        RECT 0.480 246.160 1.940 246.200 ;
        RECT 2.180 239.780 2.690 252.390 ;
        RECT 3.050 251.600 9.030 251.830 ;
        RECT 3.140 240.540 8.790 251.600 ;
        RECT 9.200 242.030 9.710 252.390 ;
        RECT 9.190 242.010 9.710 242.030 ;
        RECT 363.700 265.090 371.230 265.640 ;
        RECT 363.700 265.080 364.370 265.090 ;
        RECT 363.700 252.180 364.210 265.080 ;
        RECT 364.610 264.190 368.070 264.630 ;
        RECT 364.610 264.090 370.000 264.190 ;
        RECT 364.720 264.020 370.000 264.090 ;
        RECT 364.720 253.110 364.890 264.020 ;
        RECT 365.270 263.610 369.500 263.630 ;
        RECT 365.190 253.500 369.520 263.610 ;
        RECT 369.290 253.450 369.460 253.500 ;
        RECT 369.830 253.110 370.000 264.020 ;
        RECT 364.720 252.940 370.000 253.110 ;
        RECT 364.720 252.930 364.960 252.940 ;
        RECT 370.720 252.180 371.230 265.090 ;
        RECT 363.700 251.670 371.230 252.180 ;
        RECT 371.440 252.120 372.910 252.370 ;
        RECT 3.140 240.530 8.850 240.540 ;
        RECT 3.060 240.360 8.850 240.530 ;
        RECT 3.150 240.350 8.850 240.360 ;
        RECT 8.620 240.280 8.790 240.350 ;
        RECT 9.190 240.230 9.720 242.010 ;
        RECT 363.700 241.310 364.210 251.670 ;
        RECT 364.380 250.880 370.360 251.110 ;
        RECT 363.700 241.290 364.220 241.310 ;
        RECT 9.200 240.210 9.720 240.230 ;
        RECT 2.180 239.490 4.620 239.780 ;
        RECT 9.200 239.700 9.710 240.210 ;
        RECT 9.200 239.490 9.730 239.700 ;
        RECT 363.690 239.510 364.220 241.290 ;
        RECT 364.620 239.820 370.270 250.880 ;
        RECT 364.560 239.810 370.270 239.820 ;
        RECT 364.560 239.640 370.350 239.810 ;
        RECT 364.560 239.630 370.260 239.640 ;
        RECT 364.620 239.560 364.790 239.630 ;
        RECT 363.690 239.490 364.210 239.510 ;
        RECT 2.180 239.010 9.730 239.490 ;
        RECT 2.180 238.980 9.540 239.010 ;
        RECT 363.700 238.980 364.210 239.490 ;
        RECT 370.720 239.060 371.230 251.670 ;
        RECT 371.470 245.650 372.930 245.690 ;
        RECT 371.460 245.480 372.930 245.650 ;
        RECT 371.470 245.440 372.930 245.480 ;
        RECT 363.680 238.770 364.210 238.980 ;
        RECT 368.790 238.770 371.230 239.060 ;
        RECT 363.680 238.290 371.230 238.770 ;
        RECT 363.870 238.260 371.230 238.290 ;
        RECT 2.180 237.220 9.710 237.770 ;
        RECT 0.500 224.250 1.970 224.500 ;
        RECT 2.180 224.310 2.690 237.220 ;
        RECT 9.040 237.210 9.710 237.220 ;
        RECT 5.340 236.320 8.800 236.760 ;
        RECT 3.410 236.220 8.800 236.320 ;
        RECT 3.410 236.150 8.690 236.220 ;
        RECT 3.410 225.240 3.580 236.150 ;
        RECT 3.910 235.740 8.140 235.760 ;
        RECT 3.890 225.630 8.220 235.740 ;
        RECT 3.950 225.580 4.120 225.630 ;
        RECT 8.520 225.240 8.690 236.150 ;
        RECT 3.410 225.070 8.690 225.240 ;
        RECT 8.450 225.060 8.690 225.070 ;
        RECT 9.200 224.310 9.710 237.210 ;
        RECT 2.180 223.800 9.710 224.310 ;
        RECT 0.480 217.780 1.940 217.820 ;
        RECT 0.480 217.610 1.950 217.780 ;
        RECT 0.480 217.570 1.940 217.610 ;
        RECT 2.180 211.190 2.690 223.800 ;
        RECT 3.050 223.010 9.030 223.240 ;
        RECT 3.140 211.950 8.790 223.010 ;
        RECT 9.200 213.440 9.710 223.800 ;
        RECT 9.190 213.420 9.710 213.440 ;
        RECT 363.700 236.500 371.230 237.050 ;
        RECT 363.700 236.490 364.370 236.500 ;
        RECT 363.700 223.590 364.210 236.490 ;
        RECT 364.610 235.600 368.070 236.040 ;
        RECT 364.610 235.500 370.000 235.600 ;
        RECT 364.720 235.430 370.000 235.500 ;
        RECT 364.720 224.520 364.890 235.430 ;
        RECT 365.270 235.020 369.500 235.040 ;
        RECT 365.190 224.910 369.520 235.020 ;
        RECT 369.290 224.860 369.460 224.910 ;
        RECT 369.830 224.520 370.000 235.430 ;
        RECT 364.720 224.350 370.000 224.520 ;
        RECT 364.720 224.340 364.960 224.350 ;
        RECT 370.720 223.590 371.230 236.500 ;
        RECT 363.700 223.080 371.230 223.590 ;
        RECT 371.440 223.530 372.910 223.780 ;
        RECT 3.140 211.940 8.850 211.950 ;
        RECT 3.060 211.770 8.850 211.940 ;
        RECT 3.150 211.760 8.850 211.770 ;
        RECT 8.620 211.690 8.790 211.760 ;
        RECT 9.190 211.640 9.720 213.420 ;
        RECT 363.700 212.720 364.210 223.080 ;
        RECT 364.380 222.290 370.360 222.520 ;
        RECT 363.700 212.700 364.220 212.720 ;
        RECT 9.200 211.620 9.720 211.640 ;
        RECT 2.180 210.900 4.620 211.190 ;
        RECT 9.200 211.110 9.710 211.620 ;
        RECT 9.200 210.900 9.730 211.110 ;
        RECT 363.690 210.920 364.220 212.700 ;
        RECT 364.620 211.230 370.270 222.290 ;
        RECT 364.560 211.220 370.270 211.230 ;
        RECT 364.560 211.050 370.350 211.220 ;
        RECT 364.560 211.040 370.260 211.050 ;
        RECT 364.620 210.970 364.790 211.040 ;
        RECT 363.690 210.900 364.210 210.920 ;
        RECT 2.180 210.420 9.730 210.900 ;
        RECT 2.180 210.390 9.540 210.420 ;
        RECT 363.700 210.390 364.210 210.900 ;
        RECT 370.720 210.470 371.230 223.080 ;
        RECT 371.470 217.060 372.930 217.100 ;
        RECT 371.460 216.890 372.930 217.060 ;
        RECT 371.470 216.850 372.930 216.890 ;
        RECT 363.680 210.180 364.210 210.390 ;
        RECT 368.790 210.180 371.230 210.470 ;
        RECT 363.680 209.700 371.230 210.180 ;
        RECT 363.870 209.670 371.230 209.700 ;
        RECT 2.180 208.630 9.710 209.180 ;
        RECT 0.500 195.660 1.970 195.910 ;
        RECT 2.180 195.720 2.690 208.630 ;
        RECT 9.040 208.620 9.710 208.630 ;
        RECT 5.340 207.730 8.800 208.170 ;
        RECT 3.410 207.630 8.800 207.730 ;
        RECT 3.410 207.560 8.690 207.630 ;
        RECT 3.410 196.650 3.580 207.560 ;
        RECT 3.910 207.150 8.140 207.170 ;
        RECT 3.890 197.040 8.220 207.150 ;
        RECT 3.950 196.990 4.120 197.040 ;
        RECT 8.520 196.650 8.690 207.560 ;
        RECT 3.410 196.480 8.690 196.650 ;
        RECT 8.450 196.470 8.690 196.480 ;
        RECT 9.200 195.720 9.710 208.620 ;
        RECT 2.180 195.210 9.710 195.720 ;
        RECT 0.480 189.190 1.940 189.230 ;
        RECT 0.480 189.020 1.950 189.190 ;
        RECT 0.480 188.980 1.940 189.020 ;
        RECT 2.180 182.600 2.690 195.210 ;
        RECT 3.050 194.420 9.030 194.650 ;
        RECT 3.140 183.360 8.790 194.420 ;
        RECT 9.200 184.850 9.710 195.210 ;
        RECT 9.190 184.830 9.710 184.850 ;
        RECT 363.700 207.910 371.230 208.460 ;
        RECT 363.700 207.900 364.370 207.910 ;
        RECT 363.700 195.000 364.210 207.900 ;
        RECT 364.610 207.010 368.070 207.450 ;
        RECT 364.610 206.910 370.000 207.010 ;
        RECT 364.720 206.840 370.000 206.910 ;
        RECT 364.720 195.930 364.890 206.840 ;
        RECT 365.270 206.430 369.500 206.450 ;
        RECT 365.190 196.320 369.520 206.430 ;
        RECT 369.290 196.270 369.460 196.320 ;
        RECT 369.830 195.930 370.000 206.840 ;
        RECT 364.720 195.760 370.000 195.930 ;
        RECT 364.720 195.750 364.960 195.760 ;
        RECT 370.720 195.000 371.230 207.910 ;
        RECT 363.700 194.490 371.230 195.000 ;
        RECT 371.440 194.940 372.910 195.190 ;
        RECT 3.140 183.350 8.850 183.360 ;
        RECT 3.060 183.180 8.850 183.350 ;
        RECT 3.150 183.170 8.850 183.180 ;
        RECT 8.620 183.100 8.790 183.170 ;
        RECT 9.190 183.050 9.720 184.830 ;
        RECT 363.700 184.130 364.210 194.490 ;
        RECT 364.380 193.700 370.360 193.930 ;
        RECT 363.700 184.110 364.220 184.130 ;
        RECT 9.200 183.030 9.720 183.050 ;
        RECT 2.180 182.310 4.620 182.600 ;
        RECT 9.200 182.520 9.710 183.030 ;
        RECT 9.200 182.310 9.730 182.520 ;
        RECT 363.690 182.330 364.220 184.110 ;
        RECT 364.620 182.640 370.270 193.700 ;
        RECT 364.560 182.630 370.270 182.640 ;
        RECT 364.560 182.460 370.350 182.630 ;
        RECT 364.560 182.450 370.260 182.460 ;
        RECT 364.620 182.380 364.790 182.450 ;
        RECT 363.690 182.310 364.210 182.330 ;
        RECT 2.180 181.830 9.730 182.310 ;
        RECT 2.180 181.800 9.540 181.830 ;
        RECT 363.700 181.800 364.210 182.310 ;
        RECT 370.720 181.880 371.230 194.490 ;
        RECT 371.470 188.470 372.930 188.510 ;
        RECT 371.460 188.300 372.930 188.470 ;
        RECT 371.470 188.260 372.930 188.300 ;
        RECT 363.680 181.590 364.210 181.800 ;
        RECT 368.790 181.590 371.230 181.880 ;
        RECT 363.680 181.110 371.230 181.590 ;
        RECT 363.870 181.080 371.230 181.110 ;
        RECT 2.180 180.040 9.710 180.590 ;
        RECT 0.500 167.070 1.970 167.320 ;
        RECT 2.180 167.130 2.690 180.040 ;
        RECT 9.040 180.030 9.710 180.040 ;
        RECT 5.340 179.140 8.800 179.580 ;
        RECT 3.410 179.040 8.800 179.140 ;
        RECT 3.410 178.970 8.690 179.040 ;
        RECT 3.410 168.060 3.580 178.970 ;
        RECT 3.910 178.560 8.140 178.580 ;
        RECT 3.890 168.450 8.220 178.560 ;
        RECT 3.950 168.400 4.120 168.450 ;
        RECT 8.520 168.060 8.690 178.970 ;
        RECT 3.410 167.890 8.690 168.060 ;
        RECT 8.450 167.880 8.690 167.890 ;
        RECT 9.200 167.130 9.710 180.030 ;
        RECT 2.180 166.620 9.710 167.130 ;
        RECT 0.480 160.600 1.940 160.640 ;
        RECT 0.480 160.430 1.950 160.600 ;
        RECT 0.480 160.390 1.940 160.430 ;
        RECT 2.180 154.010 2.690 166.620 ;
        RECT 3.050 165.830 9.030 166.060 ;
        RECT 3.140 154.770 8.790 165.830 ;
        RECT 9.200 156.260 9.710 166.620 ;
        RECT 9.190 156.240 9.710 156.260 ;
        RECT 3.140 154.760 8.850 154.770 ;
        RECT 3.060 154.590 8.850 154.760 ;
        RECT 3.150 154.580 8.850 154.590 ;
        RECT 8.620 154.510 8.790 154.580 ;
        RECT 9.190 154.460 9.720 156.240 ;
        RECT 9.200 154.440 9.720 154.460 ;
        RECT 2.180 153.720 4.620 154.010 ;
        RECT 9.200 153.930 9.710 154.440 ;
        RECT 9.200 153.720 9.730 153.930 ;
        RECT 2.180 153.240 9.730 153.720 ;
        RECT 2.180 153.210 9.540 153.240 ;
        RECT 2.180 151.450 9.710 152.000 ;
        RECT 0.500 138.480 1.970 138.730 ;
        RECT 2.180 138.540 2.690 151.450 ;
        RECT 9.040 151.440 9.710 151.450 ;
        RECT 5.340 150.550 8.800 150.990 ;
        RECT 3.410 150.450 8.800 150.550 ;
        RECT 3.410 150.380 8.690 150.450 ;
        RECT 3.410 139.470 3.580 150.380 ;
        RECT 3.910 149.970 8.140 149.990 ;
        RECT 3.890 139.860 8.220 149.970 ;
        RECT 3.950 139.810 4.120 139.860 ;
        RECT 8.520 139.470 8.690 150.380 ;
        RECT 3.410 139.300 8.690 139.470 ;
        RECT 8.450 139.290 8.690 139.300 ;
        RECT 9.200 138.540 9.710 151.440 ;
        RECT 2.180 138.030 9.710 138.540 ;
        RECT 0.480 132.010 1.940 132.050 ;
        RECT 0.480 131.840 1.950 132.010 ;
        RECT 0.480 131.800 1.940 131.840 ;
        RECT 2.180 125.420 2.690 138.030 ;
        RECT 3.050 137.240 9.030 137.470 ;
        RECT 3.140 126.180 8.790 137.240 ;
        RECT 9.200 127.670 9.710 138.030 ;
        RECT 9.190 127.650 9.710 127.670 ;
        RECT 3.140 126.170 8.850 126.180 ;
        RECT 3.060 126.000 8.850 126.170 ;
        RECT 3.150 125.990 8.850 126.000 ;
        RECT 8.620 125.920 8.790 125.990 ;
        RECT 9.190 125.870 9.720 127.650 ;
        RECT 9.200 125.850 9.720 125.870 ;
        RECT 2.180 125.130 4.620 125.420 ;
        RECT 9.200 125.340 9.710 125.850 ;
        RECT 9.200 125.130 9.730 125.340 ;
        RECT 2.180 124.650 9.730 125.130 ;
        RECT 2.180 124.620 9.540 124.650 ;
        RECT 2.180 122.860 9.710 123.410 ;
        RECT 0.500 109.890 1.970 110.140 ;
        RECT 2.180 109.950 2.690 122.860 ;
        RECT 9.040 122.850 9.710 122.860 ;
        RECT 5.340 121.960 8.800 122.400 ;
        RECT 3.410 121.860 8.800 121.960 ;
        RECT 3.410 121.790 8.690 121.860 ;
        RECT 3.410 110.880 3.580 121.790 ;
        RECT 3.910 121.380 8.140 121.400 ;
        RECT 3.890 111.270 8.220 121.380 ;
        RECT 3.950 111.220 4.120 111.270 ;
        RECT 8.520 110.880 8.690 121.790 ;
        RECT 3.410 110.710 8.690 110.880 ;
        RECT 8.450 110.700 8.690 110.710 ;
        RECT 9.200 109.950 9.710 122.850 ;
        RECT 2.180 109.440 9.710 109.950 ;
        RECT 0.480 103.420 1.940 103.460 ;
        RECT 0.480 103.250 1.950 103.420 ;
        RECT 0.480 103.210 1.940 103.250 ;
        RECT 2.180 96.830 2.690 109.440 ;
        RECT 3.050 108.650 9.030 108.880 ;
        RECT 3.140 97.590 8.790 108.650 ;
        RECT 9.200 99.080 9.710 109.440 ;
        RECT 9.190 99.060 9.710 99.080 ;
        RECT 3.140 97.580 8.850 97.590 ;
        RECT 3.060 97.410 8.850 97.580 ;
        RECT 3.150 97.400 8.850 97.410 ;
        RECT 8.620 97.330 8.790 97.400 ;
        RECT 9.190 97.280 9.720 99.060 ;
        RECT 9.200 97.260 9.720 97.280 ;
        RECT 2.180 96.540 4.620 96.830 ;
        RECT 9.200 96.750 9.710 97.260 ;
        RECT 9.200 96.540 9.730 96.750 ;
        RECT 2.180 96.060 9.730 96.540 ;
        RECT 2.180 96.030 9.540 96.060 ;
        RECT 2.180 94.270 9.710 94.820 ;
        RECT 0.500 81.300 1.970 81.550 ;
        RECT 2.180 81.360 2.690 94.270 ;
        RECT 9.040 94.260 9.710 94.270 ;
        RECT 5.340 93.370 8.800 93.810 ;
        RECT 3.410 93.270 8.800 93.370 ;
        RECT 3.410 93.200 8.690 93.270 ;
        RECT 3.410 82.290 3.580 93.200 ;
        RECT 3.910 92.790 8.140 92.810 ;
        RECT 3.890 82.680 8.220 92.790 ;
        RECT 3.950 82.630 4.120 82.680 ;
        RECT 8.520 82.290 8.690 93.200 ;
        RECT 3.410 82.120 8.690 82.290 ;
        RECT 8.450 82.110 8.690 82.120 ;
        RECT 9.200 81.360 9.710 94.260 ;
        RECT 2.180 80.850 9.710 81.360 ;
        RECT 0.480 74.830 1.940 74.870 ;
        RECT 0.480 74.660 1.950 74.830 ;
        RECT 0.480 74.620 1.940 74.660 ;
        RECT 2.180 68.240 2.690 80.850 ;
        RECT 3.050 80.060 9.030 80.290 ;
        RECT 3.140 69.000 8.790 80.060 ;
        RECT 9.200 70.490 9.710 80.850 ;
        RECT 9.190 70.470 9.710 70.490 ;
        RECT 3.140 68.990 8.850 69.000 ;
        RECT 3.060 68.820 8.850 68.990 ;
        RECT 3.150 68.810 8.850 68.820 ;
        RECT 8.620 68.740 8.790 68.810 ;
        RECT 9.190 68.690 9.720 70.470 ;
        RECT 9.200 68.670 9.720 68.690 ;
        RECT 2.180 67.950 4.620 68.240 ;
        RECT 9.200 68.160 9.710 68.670 ;
        RECT 9.200 67.950 9.730 68.160 ;
        RECT 2.180 67.470 9.730 67.950 ;
        RECT 2.180 67.440 9.540 67.470 ;
        RECT 2.180 65.680 9.710 66.230 ;
        RECT 0.500 52.710 1.970 52.960 ;
        RECT 2.180 52.770 2.690 65.680 ;
        RECT 9.040 65.670 9.710 65.680 ;
        RECT 5.340 64.780 8.800 65.220 ;
        RECT 3.410 64.680 8.800 64.780 ;
        RECT 3.410 64.610 8.690 64.680 ;
        RECT 3.410 53.700 3.580 64.610 ;
        RECT 3.910 64.200 8.140 64.220 ;
        RECT 3.890 54.090 8.220 64.200 ;
        RECT 3.950 54.040 4.120 54.090 ;
        RECT 8.520 53.700 8.690 64.610 ;
        RECT 3.410 53.530 8.690 53.700 ;
        RECT 8.450 53.520 8.690 53.530 ;
        RECT 9.200 52.770 9.710 65.670 ;
        RECT 2.180 52.260 9.710 52.770 ;
        RECT 0.480 46.240 1.940 46.280 ;
        RECT 0.480 46.070 1.950 46.240 ;
        RECT 0.480 46.030 1.940 46.070 ;
        RECT 2.180 39.650 2.690 52.260 ;
        RECT 3.050 51.470 9.030 51.700 ;
        RECT 3.140 40.410 8.790 51.470 ;
        RECT 9.200 41.900 9.710 52.260 ;
        RECT 9.190 41.880 9.710 41.900 ;
        RECT 3.140 40.400 8.850 40.410 ;
        RECT 3.060 40.230 8.850 40.400 ;
        RECT 3.150 40.220 8.850 40.230 ;
        RECT 8.620 40.150 8.790 40.220 ;
        RECT 9.190 40.100 9.720 41.880 ;
        RECT 9.200 40.080 9.720 40.100 ;
        RECT 2.180 39.360 4.620 39.650 ;
        RECT 9.200 39.570 9.710 40.080 ;
        RECT 9.200 39.360 9.730 39.570 ;
        RECT 2.180 38.880 9.730 39.360 ;
        RECT 2.180 38.850 9.540 38.880 ;
        RECT 2.180 37.090 9.710 37.640 ;
        RECT 0.500 24.120 1.970 24.370 ;
        RECT 2.180 24.180 2.690 37.090 ;
        RECT 9.040 37.080 9.710 37.090 ;
        RECT 5.340 36.190 8.800 36.630 ;
        RECT 3.410 36.090 8.800 36.190 ;
        RECT 3.410 36.020 8.690 36.090 ;
        RECT 3.410 25.110 3.580 36.020 ;
        RECT 3.910 35.610 8.140 35.630 ;
        RECT 3.890 25.500 8.220 35.610 ;
        RECT 3.950 25.450 4.120 25.500 ;
        RECT 8.520 25.110 8.690 36.020 ;
        RECT 3.410 24.940 8.690 25.110 ;
        RECT 8.450 24.930 8.690 24.940 ;
        RECT 9.200 24.180 9.710 37.080 ;
        RECT 2.180 23.670 9.710 24.180 ;
        RECT 0.480 17.650 1.940 17.690 ;
        RECT 0.480 17.480 1.950 17.650 ;
        RECT 0.480 17.440 1.940 17.480 ;
        RECT 2.180 11.060 2.690 23.670 ;
        RECT 3.050 22.880 9.030 23.110 ;
        RECT 3.140 11.820 8.790 22.880 ;
        RECT 9.200 13.310 9.710 23.670 ;
        RECT 9.190 13.290 9.710 13.310 ;
        RECT 3.140 11.810 8.850 11.820 ;
        RECT 3.060 11.640 8.850 11.810 ;
        RECT 3.150 11.630 8.850 11.640 ;
        RECT 8.620 11.560 8.790 11.630 ;
        RECT 9.190 11.510 9.720 13.290 ;
        RECT 9.200 11.490 9.720 11.510 ;
        RECT 2.180 10.770 4.620 11.060 ;
        RECT 9.200 10.980 9.710 11.490 ;
        RECT 9.200 10.770 9.730 10.980 ;
        RECT 2.180 10.290 9.730 10.770 ;
        RECT 2.180 10.260 9.540 10.290 ;
      LAYER mcon ;
        RECT 31.360 388.720 31.530 388.890 ;
        RECT 31.360 388.380 31.530 388.550 ;
        RECT 31.360 388.040 31.530 388.210 ;
        RECT 31.360 387.700 31.530 387.870 ;
        RECT 38.040 388.700 38.210 388.870 ;
        RECT 38.040 388.360 38.210 388.530 ;
        RECT 38.040 388.020 38.210 388.190 ;
        RECT 38.040 387.680 38.210 387.850 ;
        RECT 59.950 388.720 60.120 388.890 ;
        RECT 59.950 388.380 60.120 388.550 ;
        RECT 59.950 388.040 60.120 388.210 ;
        RECT 59.950 387.700 60.120 387.870 ;
        RECT 66.630 388.700 66.800 388.870 ;
        RECT 66.630 388.360 66.800 388.530 ;
        RECT 66.630 388.020 66.800 388.190 ;
        RECT 66.630 387.680 66.800 387.850 ;
        RECT 88.540 388.720 88.710 388.890 ;
        RECT 88.540 388.380 88.710 388.550 ;
        RECT 88.540 388.040 88.710 388.210 ;
        RECT 88.540 387.700 88.710 387.870 ;
        RECT 95.220 388.700 95.390 388.870 ;
        RECT 95.220 388.360 95.390 388.530 ;
        RECT 95.220 388.020 95.390 388.190 ;
        RECT 95.220 387.680 95.390 387.850 ;
        RECT 172.560 388.720 172.730 388.890 ;
        RECT 172.560 388.380 172.730 388.550 ;
        RECT 172.560 388.040 172.730 388.210 ;
        RECT 172.560 387.700 172.730 387.870 ;
        RECT 179.240 388.700 179.410 388.870 ;
        RECT 179.240 388.360 179.410 388.530 ;
        RECT 179.240 388.020 179.410 388.190 ;
        RECT 179.240 387.680 179.410 387.850 ;
        RECT 201.150 388.720 201.320 388.890 ;
        RECT 201.150 388.380 201.320 388.550 ;
        RECT 201.150 388.040 201.320 388.210 ;
        RECT 201.150 387.700 201.320 387.870 ;
        RECT 207.830 388.700 208.000 388.870 ;
        RECT 207.830 388.360 208.000 388.530 ;
        RECT 207.830 388.020 208.000 388.190 ;
        RECT 207.830 387.680 208.000 387.850 ;
        RECT 229.740 388.720 229.910 388.890 ;
        RECT 229.740 388.380 229.910 388.550 ;
        RECT 229.740 388.040 229.910 388.210 ;
        RECT 229.740 387.700 229.910 387.870 ;
        RECT 236.420 388.700 236.590 388.870 ;
        RECT 236.420 388.360 236.590 388.530 ;
        RECT 236.420 388.020 236.590 388.190 ;
        RECT 236.420 387.680 236.590 387.850 ;
        RECT 258.330 388.720 258.500 388.890 ;
        RECT 258.330 388.380 258.500 388.550 ;
        RECT 258.330 388.040 258.500 388.210 ;
        RECT 258.330 387.700 258.500 387.870 ;
        RECT 265.010 388.700 265.180 388.870 ;
        RECT 265.010 388.360 265.180 388.530 ;
        RECT 265.010 388.020 265.180 388.190 ;
        RECT 265.010 387.680 265.180 387.850 ;
        RECT 286.920 388.720 287.090 388.890 ;
        RECT 286.920 388.380 287.090 388.550 ;
        RECT 286.920 388.040 287.090 388.210 ;
        RECT 286.920 387.700 287.090 387.870 ;
        RECT 293.600 388.700 293.770 388.870 ;
        RECT 293.600 388.360 293.770 388.530 ;
        RECT 293.600 388.020 293.770 388.190 ;
        RECT 293.600 387.680 293.770 387.850 ;
        RECT 315.510 388.720 315.680 388.890 ;
        RECT 315.510 388.380 315.680 388.550 ;
        RECT 315.510 388.040 315.680 388.210 ;
        RECT 315.510 387.700 315.680 387.870 ;
        RECT 322.190 388.700 322.360 388.870 ;
        RECT 322.190 388.360 322.360 388.530 ;
        RECT 322.190 388.020 322.360 388.190 ;
        RECT 322.190 387.680 322.360 387.850 ;
        RECT 344.100 388.720 344.270 388.890 ;
        RECT 344.100 388.380 344.270 388.550 ;
        RECT 344.100 388.040 344.270 388.210 ;
        RECT 344.100 387.700 344.270 387.870 ;
        RECT 350.780 388.700 350.950 388.870 ;
        RECT 350.780 388.360 350.950 388.530 ;
        RECT 350.780 388.020 350.950 388.190 ;
        RECT 350.780 387.680 350.950 387.850 ;
        RECT 24.220 387.050 26.080 387.060 ;
        RECT 24.220 386.880 26.090 387.050 ;
        RECT 47.580 386.870 50.740 387.050 ;
        RECT 24.300 385.920 24.480 386.710 ;
        RECT 24.310 384.790 24.480 385.920 ;
        RECT 24.660 384.780 24.840 386.700 ;
        RECT 25.850 385.750 36.830 385.920 ;
        RECT 25.850 385.130 36.830 385.300 ;
        RECT 2.580 380.350 3.510 380.550 ;
        RECT 2.350 376.780 2.530 379.940 ;
        RECT 5.450 379.280 8.750 379.630 ;
        RECT 0.530 367.240 0.700 367.410 ;
        RECT 0.870 367.240 1.040 367.410 ;
        RECT 1.210 367.240 1.380 367.410 ;
        RECT 1.550 367.240 1.720 367.410 ;
        RECT 4.240 368.780 4.410 378.230 ;
        RECT 4.990 368.770 5.160 378.160 ;
        RECT 5.710 368.800 5.880 378.200 ;
        RECT 6.370 368.810 6.540 378.180 ;
        RECT 7.020 368.800 7.190 378.250 ;
        RECT 7.660 368.810 7.830 378.200 ;
        RECT 25.860 384.510 36.840 384.680 ;
        RECT 25.880 383.930 36.860 384.100 ;
        RECT 25.890 383.340 36.870 383.510 ;
        RECT 25.890 382.740 36.870 382.910 ;
        RECT 25.840 382.140 36.820 382.310 ;
        RECT 25.850 381.530 36.830 381.700 ;
        RECT 25.840 380.930 36.820 381.100 ;
        RECT 39.580 384.990 49.030 385.160 ;
        RECT 39.570 384.240 48.960 384.410 ;
        RECT 39.600 383.520 49.000 383.690 ;
        RECT 39.610 382.860 48.980 383.030 ;
        RECT 39.600 382.210 49.050 382.380 ;
        RECT 39.610 381.570 49.000 381.740 ;
        RECT 51.150 385.890 51.350 386.820 ;
        RECT 50.080 380.650 50.430 383.950 ;
        RECT 52.810 387.050 54.670 387.060 ;
        RECT 52.810 386.880 54.680 387.050 ;
        RECT 76.170 386.870 79.330 387.050 ;
        RECT 52.890 385.920 53.070 386.710 ;
        RECT 52.900 384.790 53.070 385.920 ;
        RECT 53.250 384.780 53.430 386.700 ;
        RECT 54.440 385.750 65.420 385.920 ;
        RECT 54.440 385.130 65.420 385.300 ;
        RECT 54.450 384.510 65.430 384.680 ;
        RECT 54.470 383.930 65.450 384.100 ;
        RECT 54.480 383.340 65.460 383.510 ;
        RECT 54.480 382.740 65.460 382.910 ;
        RECT 54.430 382.140 65.410 382.310 ;
        RECT 54.440 381.530 65.420 381.700 ;
        RECT 54.430 380.930 65.410 381.100 ;
        RECT 68.170 384.990 77.620 385.160 ;
        RECT 68.160 384.240 77.550 384.410 ;
        RECT 68.190 383.520 77.590 383.690 ;
        RECT 68.200 382.860 77.570 383.030 ;
        RECT 68.190 382.210 77.640 382.380 ;
        RECT 68.200 381.570 77.590 381.740 ;
        RECT 79.740 385.890 79.940 386.820 ;
        RECT 78.670 380.650 79.020 383.950 ;
        RECT 81.400 387.050 83.260 387.060 ;
        RECT 81.400 386.880 83.270 387.050 ;
        RECT 104.760 386.870 107.920 387.050 ;
        RECT 81.480 385.920 81.660 386.710 ;
        RECT 81.490 384.790 81.660 385.920 ;
        RECT 81.840 384.780 82.020 386.700 ;
        RECT 83.030 385.750 94.010 385.920 ;
        RECT 83.030 385.130 94.010 385.300 ;
        RECT 83.040 384.510 94.020 384.680 ;
        RECT 83.060 383.930 94.040 384.100 ;
        RECT 83.070 383.340 94.050 383.510 ;
        RECT 83.070 382.740 94.050 382.910 ;
        RECT 83.020 382.140 94.000 382.310 ;
        RECT 83.030 381.530 94.010 381.700 ;
        RECT 83.020 380.930 94.000 381.100 ;
        RECT 96.760 384.990 106.210 385.160 ;
        RECT 96.750 384.240 106.140 384.410 ;
        RECT 96.780 383.520 106.180 383.690 ;
        RECT 96.790 382.860 106.160 383.030 ;
        RECT 96.780 382.210 106.230 382.380 ;
        RECT 96.790 381.570 106.180 381.740 ;
        RECT 108.330 385.890 108.530 386.820 ;
        RECT 150.530 386.630 150.700 386.800 ;
        RECT 150.530 386.290 150.700 386.460 ;
        RECT 150.530 385.950 150.700 386.120 ;
        RECT 157.280 386.670 157.450 386.840 ;
        RECT 157.280 386.330 157.450 386.500 ;
        RECT 157.280 385.990 157.450 386.160 ;
        RECT 107.260 380.650 107.610 383.950 ;
        RECT 165.420 387.050 167.280 387.060 ;
        RECT 165.420 386.880 167.290 387.050 ;
        RECT 188.780 386.870 191.940 387.050 ;
        RECT 165.500 385.920 165.680 386.710 ;
        RECT 165.510 385.330 165.680 385.920 ;
        RECT 165.860 385.330 166.040 386.700 ;
        RECT 167.050 385.750 178.030 385.920 ;
        RECT 130.080 385.160 153.980 385.330 ;
        RECT 162.860 385.160 184.030 385.330 ;
        RECT 165.510 384.790 165.680 385.160 ;
        RECT 165.860 384.780 166.040 385.160 ;
        RECT 167.050 385.130 178.030 385.160 ;
        RECT 129.500 380.990 129.670 381.160 ;
        RECT 132.370 381.200 132.540 381.370 ;
        RECT 130.910 380.990 131.080 381.160 ;
        RECT 147.710 381.020 147.880 381.190 ;
        RECT 147.710 380.670 147.880 380.840 ;
        RECT 132.370 380.410 132.540 380.580 ;
        RECT 147.710 380.330 147.880 380.500 ;
        RECT 153.570 380.930 153.740 381.100 ;
        RECT 153.570 380.480 153.740 380.650 ;
        RECT 158.270 380.880 158.440 381.050 ;
        RECT 158.270 380.430 158.440 380.600 ;
        RECT 129.500 380.140 129.670 380.310 ;
        RECT 130.220 380.130 130.390 380.300 ;
        RECT 130.910 380.140 131.080 380.310 ;
        RECT 167.060 384.510 178.040 384.680 ;
        RECT 167.080 383.930 178.060 384.100 ;
        RECT 167.090 383.340 178.070 383.510 ;
        RECT 167.090 382.740 178.070 382.910 ;
        RECT 167.040 382.140 178.020 382.310 ;
        RECT 167.050 381.530 178.030 381.700 ;
        RECT 167.040 380.930 178.020 381.100 ;
        RECT 180.780 384.990 190.230 385.160 ;
        RECT 180.770 384.240 190.160 384.410 ;
        RECT 180.800 383.520 190.200 383.690 ;
        RECT 180.810 382.860 190.180 383.030 ;
        RECT 180.800 382.210 190.250 382.380 ;
        RECT 180.810 381.570 190.200 381.740 ;
        RECT 192.350 385.890 192.550 386.820 ;
        RECT 191.280 380.650 191.630 383.950 ;
        RECT 129.680 379.730 129.850 379.900 ;
        RECT 130.740 379.730 130.910 379.900 ;
        RECT 129.500 379.320 129.670 379.490 ;
        RECT 130.220 379.290 130.390 379.460 ;
        RECT 130.910 379.320 131.080 379.490 ;
        RECT 194.010 387.050 195.870 387.060 ;
        RECT 194.010 386.880 195.880 387.050 ;
        RECT 217.370 386.870 220.530 387.050 ;
        RECT 194.090 385.920 194.270 386.710 ;
        RECT 194.100 384.790 194.270 385.920 ;
        RECT 194.450 384.780 194.630 386.700 ;
        RECT 195.640 385.750 206.620 385.920 ;
        RECT 195.640 385.130 206.620 385.300 ;
        RECT 195.650 384.510 206.630 384.680 ;
        RECT 195.670 383.930 206.650 384.100 ;
        RECT 195.680 383.340 206.660 383.510 ;
        RECT 195.680 382.740 206.660 382.910 ;
        RECT 195.630 382.140 206.610 382.310 ;
        RECT 195.640 381.530 206.620 381.700 ;
        RECT 195.630 380.930 206.610 381.100 ;
        RECT 209.370 384.990 218.820 385.160 ;
        RECT 209.360 384.240 218.750 384.410 ;
        RECT 209.390 383.520 218.790 383.690 ;
        RECT 209.400 382.860 218.770 383.030 ;
        RECT 209.390 382.210 218.840 382.380 ;
        RECT 209.400 381.570 218.790 381.740 ;
        RECT 220.940 385.890 221.140 386.820 ;
        RECT 219.870 380.650 220.220 383.950 ;
        RECT 222.600 387.050 224.460 387.060 ;
        RECT 222.600 386.880 224.470 387.050 ;
        RECT 245.960 386.870 249.120 387.050 ;
        RECT 222.680 385.920 222.860 386.710 ;
        RECT 222.690 384.790 222.860 385.920 ;
        RECT 223.040 384.780 223.220 386.700 ;
        RECT 224.230 385.750 235.210 385.920 ;
        RECT 224.230 385.130 235.210 385.300 ;
        RECT 224.240 384.510 235.220 384.680 ;
        RECT 224.260 383.930 235.240 384.100 ;
        RECT 224.270 383.340 235.250 383.510 ;
        RECT 224.270 382.740 235.250 382.910 ;
        RECT 224.220 382.140 235.200 382.310 ;
        RECT 224.230 381.530 235.210 381.700 ;
        RECT 224.220 380.930 235.200 381.100 ;
        RECT 237.960 384.990 247.410 385.160 ;
        RECT 237.950 384.240 247.340 384.410 ;
        RECT 237.980 383.520 247.380 383.690 ;
        RECT 237.990 382.860 247.360 383.030 ;
        RECT 237.980 382.210 247.430 382.380 ;
        RECT 237.990 381.570 247.380 381.740 ;
        RECT 249.530 385.890 249.730 386.820 ;
        RECT 248.460 380.650 248.810 383.950 ;
        RECT 251.190 387.050 253.050 387.060 ;
        RECT 251.190 386.880 253.060 387.050 ;
        RECT 274.550 386.870 277.710 387.050 ;
        RECT 251.270 385.920 251.450 386.710 ;
        RECT 251.280 384.790 251.450 385.920 ;
        RECT 251.630 384.780 251.810 386.700 ;
        RECT 252.820 385.750 263.800 385.920 ;
        RECT 252.820 385.130 263.800 385.300 ;
        RECT 252.830 384.510 263.810 384.680 ;
        RECT 252.850 383.930 263.830 384.100 ;
        RECT 252.860 383.340 263.840 383.510 ;
        RECT 252.860 382.740 263.840 382.910 ;
        RECT 252.810 382.140 263.790 382.310 ;
        RECT 252.820 381.530 263.800 381.700 ;
        RECT 252.810 380.930 263.790 381.100 ;
        RECT 266.550 384.990 276.000 385.160 ;
        RECT 266.540 384.240 275.930 384.410 ;
        RECT 266.570 383.520 275.970 383.690 ;
        RECT 266.580 382.860 275.950 383.030 ;
        RECT 266.570 382.210 276.020 382.380 ;
        RECT 266.580 381.570 275.970 381.740 ;
        RECT 278.120 385.890 278.320 386.820 ;
        RECT 277.050 380.650 277.400 383.950 ;
        RECT 279.780 387.050 281.640 387.060 ;
        RECT 279.780 386.880 281.650 387.050 ;
        RECT 303.140 386.870 306.300 387.050 ;
        RECT 279.860 385.920 280.040 386.710 ;
        RECT 279.870 384.790 280.040 385.920 ;
        RECT 280.220 384.780 280.400 386.700 ;
        RECT 281.410 385.750 292.390 385.920 ;
        RECT 281.410 385.130 292.390 385.300 ;
        RECT 281.420 384.510 292.400 384.680 ;
        RECT 281.440 383.930 292.420 384.100 ;
        RECT 281.450 383.340 292.430 383.510 ;
        RECT 281.450 382.740 292.430 382.910 ;
        RECT 281.400 382.140 292.380 382.310 ;
        RECT 281.410 381.530 292.390 381.700 ;
        RECT 281.400 380.930 292.380 381.100 ;
        RECT 295.140 384.990 304.590 385.160 ;
        RECT 295.130 384.240 304.520 384.410 ;
        RECT 295.160 383.520 304.560 383.690 ;
        RECT 295.170 382.860 304.540 383.030 ;
        RECT 295.160 382.210 304.610 382.380 ;
        RECT 295.170 381.570 304.560 381.740 ;
        RECT 306.710 385.890 306.910 386.820 ;
        RECT 305.640 380.650 305.990 383.950 ;
        RECT 308.370 387.050 310.230 387.060 ;
        RECT 308.370 386.880 310.240 387.050 ;
        RECT 331.730 386.870 334.890 387.050 ;
        RECT 308.450 385.920 308.630 386.710 ;
        RECT 308.460 384.790 308.630 385.920 ;
        RECT 308.810 384.780 308.990 386.700 ;
        RECT 310.000 385.750 320.980 385.920 ;
        RECT 310.000 385.130 320.980 385.300 ;
        RECT 310.010 384.510 320.990 384.680 ;
        RECT 310.030 383.930 321.010 384.100 ;
        RECT 310.040 383.340 321.020 383.510 ;
        RECT 310.040 382.740 321.020 382.910 ;
        RECT 309.990 382.140 320.970 382.310 ;
        RECT 310.000 381.530 320.980 381.700 ;
        RECT 309.990 380.930 320.970 381.100 ;
        RECT 323.730 384.990 333.180 385.160 ;
        RECT 323.720 384.240 333.110 384.410 ;
        RECT 323.750 383.520 333.150 383.690 ;
        RECT 323.760 382.860 333.130 383.030 ;
        RECT 323.750 382.210 333.200 382.380 ;
        RECT 323.760 381.570 333.150 381.740 ;
        RECT 335.300 385.890 335.500 386.820 ;
        RECT 334.230 380.650 334.580 383.950 ;
        RECT 336.960 387.050 338.820 387.060 ;
        RECT 336.960 386.880 338.830 387.050 ;
        RECT 360.320 386.870 363.480 387.050 ;
        RECT 337.040 385.920 337.220 386.710 ;
        RECT 337.050 384.790 337.220 385.920 ;
        RECT 337.400 384.780 337.580 386.700 ;
        RECT 338.590 385.750 349.570 385.920 ;
        RECT 338.590 385.130 349.570 385.300 ;
        RECT 338.600 384.510 349.580 384.680 ;
        RECT 338.620 383.930 349.600 384.100 ;
        RECT 338.630 383.340 349.610 383.510 ;
        RECT 338.630 382.740 349.610 382.910 ;
        RECT 338.580 382.140 349.560 382.310 ;
        RECT 338.590 381.530 349.570 381.700 ;
        RECT 338.580 380.930 349.560 381.100 ;
        RECT 352.320 384.990 361.770 385.160 ;
        RECT 352.310 384.240 361.700 384.410 ;
        RECT 352.340 383.520 361.740 383.690 ;
        RECT 352.350 382.860 361.720 383.030 ;
        RECT 352.340 382.210 361.790 382.380 ;
        RECT 352.350 381.570 361.740 381.740 ;
        RECT 363.890 385.890 364.090 386.820 ;
        RECT 362.820 380.650 363.170 383.950 ;
        RECT 145.610 379.390 145.780 379.560 ;
        RECT 146.970 379.470 147.140 379.640 ;
        RECT 147.660 379.460 147.830 379.630 ;
        RECT 132.370 378.980 132.540 379.150 ;
        RECT 129.500 378.480 129.670 378.650 ;
        RECT 130.910 378.480 131.080 378.650 ;
        RECT 131.640 378.220 131.810 378.390 ;
        RECT 131.630 377.700 131.800 377.870 ;
        RECT 132.380 377.580 132.550 377.750 ;
        RECT 129.500 377.360 129.670 377.530 ;
        RECT 130.910 377.360 131.080 377.530 ;
        RECT 130.200 376.490 130.370 376.660 ;
        RECT 131.630 376.510 131.800 376.680 ;
        RECT 134.390 376.160 134.560 376.330 ;
        RECT 129.410 375.910 129.580 376.080 ;
        RECT 130.340 375.910 130.510 376.080 ;
        RECT 131.040 375.910 131.210 376.080 ;
        RECT 131.780 375.910 131.950 376.080 ;
        RECT 132.490 375.900 132.660 376.070 ;
        RECT 147.710 378.220 147.880 378.390 ;
        RECT 147.710 377.870 147.880 378.040 ;
        RECT 147.710 377.530 147.880 377.700 ;
        RECT 153.570 377.940 153.740 378.110 ;
        RECT 153.570 377.490 153.740 377.660 ;
        RECT 153.570 376.930 153.740 377.100 ;
        RECT 147.710 376.670 147.880 376.840 ;
        RECT 147.710 376.320 147.880 376.490 ;
        RECT 153.570 376.480 153.740 376.650 ;
        RECT 147.710 375.980 147.880 376.150 ;
        RECT 369.900 379.630 370.830 379.830 ;
        RECT 157.490 377.420 157.660 377.590 ;
        RECT 156.520 377.200 156.690 377.370 ;
        RECT 156.860 377.200 157.030 377.370 ;
        RECT 157.200 377.200 157.370 377.370 ;
        RECT 157.540 377.200 157.710 377.370 ;
        RECT 157.880 377.200 158.050 377.370 ;
        RECT 158.220 377.200 158.390 377.370 ;
        RECT 144.890 375.730 145.060 375.900 ;
        RECT 154.750 375.750 154.920 375.920 ;
        RECT 144.900 371.370 145.330 372.110 ;
        RECT 165.600 370.210 165.810 370.420 ;
        RECT 170.480 370.320 170.650 370.490 ;
        RECT 164.130 369.840 164.300 370.010 ;
        RECT 171.520 369.970 171.690 370.140 ;
        RECT 171.520 369.620 171.690 369.790 ;
        RECT 165.600 368.660 165.810 368.870 ;
        RECT 170.480 368.770 170.650 368.940 ;
        RECT 164.130 368.290 164.300 368.460 ;
        RECT 140.880 367.990 141.050 368.160 ;
        RECT 141.970 368.000 142.140 368.170 ;
        RECT 171.520 368.420 171.690 368.590 ;
        RECT 171.520 368.070 171.690 368.240 ;
        RECT 193.190 368.210 193.450 369.030 ;
        RECT 205.140 368.240 205.460 369.030 ;
        RECT 207.420 368.570 207.600 368.740 ;
        RECT 207.850 368.550 208.020 368.720 ;
        RECT 205.610 368.270 205.780 368.440 ;
        RECT 140.660 367.580 140.830 367.750 ;
        RECT 142.810 367.530 142.980 367.700 ;
        RECT 205.960 367.430 206.140 367.620 ;
        RECT 140.880 367.070 141.050 367.240 ;
        RECT 141.970 367.080 142.140 367.250 ;
        RECT 165.600 367.110 165.810 367.320 ;
        RECT 170.480 367.220 170.650 367.390 ;
        RECT 0.510 360.560 0.680 360.730 ;
        RECT 0.850 360.560 1.020 360.730 ;
        RECT 1.190 360.560 1.360 360.730 ;
        RECT 1.530 360.560 1.700 360.730 ;
        RECT 2.350 355.280 2.520 355.290 ;
        RECT 2.340 353.420 2.520 355.280 ;
        RECT 3.480 355.050 3.650 366.030 ;
        RECT 4.100 355.050 4.270 366.030 ;
        RECT 4.720 355.060 4.890 366.040 ;
        RECT 5.300 355.080 5.470 366.060 ;
        RECT 5.890 355.090 6.060 366.070 ;
        RECT 6.490 355.090 6.660 366.070 ;
        RECT 7.090 355.040 7.260 366.020 ;
        RECT 7.700 355.050 7.870 366.030 ;
        RECT 8.300 355.040 8.470 366.020 ;
        RECT 140.660 366.660 140.830 366.830 ;
        RECT 164.130 366.740 164.300 366.910 ;
        RECT 140.880 366.150 141.050 366.320 ;
        RECT 141.970 366.160 142.140 366.330 ;
        RECT 171.520 366.870 171.690 367.040 ;
        RECT 171.520 366.520 171.690 366.690 ;
        RECT 208.320 367.990 208.490 368.160 ;
        RECT 235.480 368.270 235.650 368.440 ;
        RECT 210.560 367.690 210.730 367.860 ;
        RECT 228.640 367.690 228.810 367.860 ;
        RECT 210.560 367.240 210.730 367.410 ;
        RECT 207.040 366.870 207.210 367.040 ;
        RECT 216.010 367.090 216.280 367.360 ;
        RECT 224.980 367.090 225.250 367.360 ;
        RECT 228.640 367.240 228.810 367.410 ;
        RECT 233.810 367.440 233.980 367.610 ;
        RECT 207.850 366.560 208.020 366.730 ;
        RECT 140.660 365.740 140.830 365.910 ;
        RECT 165.600 365.560 165.810 365.770 ;
        RECT 170.480 365.670 170.650 365.840 ;
        RECT 235.120 367.430 235.300 367.620 ;
        RECT 213.690 365.980 213.860 366.150 ;
        RECT 227.400 365.980 227.570 366.150 ;
        RECT 140.690 365.170 140.860 365.340 ;
        RECT 141.990 365.070 142.160 365.240 ;
        RECT 164.130 365.190 164.300 365.360 ;
        RECT 171.520 365.320 171.690 365.490 ;
        RECT 171.520 364.970 171.690 365.140 ;
        RECT 205.960 364.630 206.140 364.820 ;
        RECT 140.690 364.210 140.860 364.380 ;
        RECT 141.990 364.110 142.160 364.280 ;
        RECT 208.320 365.670 208.490 365.840 ;
        RECT 207.860 365.490 208.030 365.660 ;
        RECT 207.030 365.180 207.200 365.350 ;
        RECT 216.010 365.360 216.280 365.630 ;
        RECT 224.980 365.360 225.250 365.630 ;
        RECT 364.660 378.560 367.960 378.910 ;
        RECT 365.580 368.090 365.750 377.480 ;
        RECT 366.220 368.080 366.390 377.530 ;
        RECT 366.870 368.090 367.040 377.460 ;
        RECT 367.530 368.080 367.700 377.480 ;
        RECT 368.250 368.050 368.420 377.440 ;
        RECT 369.000 368.060 369.170 377.510 ;
        RECT 370.880 376.060 371.060 379.220 ;
        RECT 371.690 366.520 371.860 366.690 ;
        RECT 372.030 366.520 372.200 366.690 ;
        RECT 372.370 366.520 372.540 366.690 ;
        RECT 372.710 366.520 372.880 366.690 ;
        RECT 210.560 364.740 210.730 364.910 ;
        RECT 210.560 364.290 210.730 364.460 ;
        RECT 228.640 364.740 228.810 364.910 ;
        RECT 232.340 365.090 232.510 365.260 ;
        RECT 233.420 365.120 233.590 365.230 ;
        RECT 233.300 365.060 233.590 365.120 ;
        RECT 233.300 364.950 233.470 365.060 ;
        RECT 233.910 365.090 234.080 365.260 ;
        RECT 233.810 364.680 233.980 364.850 ;
        RECT 234.430 364.960 234.600 365.130 ;
        RECT 234.390 364.780 234.560 364.950 ;
        RECT 235.120 364.630 235.300 364.820 ;
        RECT 236.640 364.830 236.810 365.000 ;
        RECT 228.640 364.290 228.810 364.460 ;
        RECT 230.890 364.310 231.060 364.480 ;
        RECT 231.390 364.340 231.560 364.510 ;
        RECT 208.310 364.090 208.480 364.260 ;
        RECT 205.610 363.810 205.780 363.980 ;
        RECT 233.570 364.230 233.740 364.400 ;
        RECT 234.890 364.340 235.060 364.510 ;
        RECT 235.370 364.460 235.540 364.630 ;
        RECT 207.420 363.510 207.600 363.680 ;
        RECT 207.880 363.580 208.050 363.750 ;
        RECT 232.450 363.710 232.620 363.880 ;
        RECT 140.690 363.250 140.860 363.420 ;
        RECT 234.340 364.130 234.510 364.300 ;
        RECT 235.480 363.810 235.650 363.980 ;
        RECT 233.660 363.510 233.840 363.680 ;
        RECT 231.390 363.340 231.560 363.510 ;
        RECT 141.990 363.150 142.160 363.320 ;
        RECT 183.480 362.920 183.650 363.090 ;
        RECT 142.390 362.710 142.560 362.880 ;
        RECT 184.320 362.800 184.490 362.970 ;
        RECT 185.070 362.800 185.240 362.970 ;
        RECT 164.130 361.660 164.300 361.830 ;
        RECT 171.520 361.880 171.690 362.050 ;
        RECT 188.050 362.470 188.220 362.640 ;
        RECT 183.760 362.170 183.930 362.340 ;
        RECT 188.450 362.920 188.620 363.090 ;
        RECT 188.450 362.580 188.620 362.750 ;
        RECT 207.420 362.540 207.600 362.710 ;
        RECT 205.610 362.240 205.780 362.410 ;
        RECT 165.600 361.250 165.810 361.460 ;
        RECT 171.520 361.530 171.690 361.700 ;
        RECT 170.480 361.180 170.650 361.350 ;
        RECT 183.760 361.280 183.930 361.450 ;
        RECT 205.960 361.400 206.140 361.590 ;
        RECT 188.050 360.980 188.220 361.150 ;
        RECT 164.130 360.110 164.300 360.280 ;
        RECT 184.320 360.650 184.490 360.820 ;
        RECT 185.070 360.650 185.240 360.820 ;
        RECT 187.070 360.660 187.240 360.830 ;
        RECT 188.450 361.210 188.620 361.380 ;
        RECT 188.450 360.870 188.620 361.040 ;
        RECT 171.520 360.330 171.690 360.500 ;
        RECT 234.340 363.310 234.510 363.480 ;
        RECT 234.890 363.340 235.060 363.510 ;
        RECT 236.030 363.520 236.200 363.690 ;
        RECT 235.370 362.980 235.540 363.150 ;
        RECT 232.340 362.590 232.510 362.760 ;
        RECT 233.300 362.730 233.470 362.900 ;
        RECT 234.430 362.830 234.600 362.890 ;
        RECT 233.180 362.430 233.350 362.600 ;
        RECT 233.910 362.590 234.080 362.760 ;
        RECT 234.390 362.720 234.600 362.830 ;
        RECT 234.390 362.660 234.560 362.720 ;
        RECT 236.690 362.610 236.860 362.780 ;
        RECT 212.450 361.660 212.620 361.830 ;
        RECT 214.540 361.820 214.710 361.990 ;
        RECT 232.340 362.070 232.510 362.240 ;
        RECT 207.280 361.410 207.450 361.580 ;
        RECT 228.640 361.660 228.810 361.830 ;
        RECT 233.300 361.930 233.470 362.100 ;
        RECT 233.910 362.070 234.080 362.240 ;
        RECT 235.480 362.240 235.650 362.410 ;
        RECT 212.450 361.210 212.620 361.380 ;
        RECT 216.010 361.060 216.280 361.330 ;
        RECT 224.980 361.060 225.250 361.330 ;
        RECT 233.610 361.630 233.780 361.800 ;
        RECT 234.430 361.990 234.600 362.110 ;
        RECT 234.390 361.940 234.600 361.990 ;
        RECT 234.390 361.820 234.560 361.940 ;
        RECT 228.640 361.210 228.810 361.380 ;
        RECT 230.890 361.290 231.060 361.460 ;
        RECT 231.390 361.320 231.560 361.490 ;
        RECT 233.810 361.410 233.980 361.580 ;
        RECT 236.680 361.890 236.850 362.060 ;
        RECT 165.600 359.700 165.810 359.910 ;
        RECT 171.520 359.980 171.690 360.150 ;
        RECT 183.480 359.990 183.650 360.160 ;
        RECT 170.480 359.630 170.650 359.800 ;
        RECT 184.320 359.870 184.490 360.040 ;
        RECT 185.070 359.870 185.240 360.040 ;
        RECT 164.130 358.560 164.300 358.730 ;
        RECT 188.050 359.540 188.220 359.710 ;
        RECT 183.760 359.240 183.930 359.410 ;
        RECT 188.450 359.990 188.620 360.160 ;
        RECT 188.450 359.650 188.620 359.820 ;
        RECT 234.340 361.170 234.510 361.340 ;
        RECT 234.890 361.320 235.060 361.490 ;
        RECT 235.120 361.400 235.300 361.590 ;
        RECT 235.370 361.500 235.540 361.670 ;
        RECT 236.030 360.930 236.200 361.100 ;
        RECT 231.390 360.320 231.560 360.490 ;
        RECT 234.340 360.350 234.510 360.520 ;
        RECT 234.740 360.490 234.920 360.550 ;
        RECT 234.740 360.360 235.060 360.490 ;
        RECT 213.690 359.950 213.860 360.120 ;
        RECT 227.400 359.950 227.570 360.120 ;
        RECT 171.520 358.780 171.690 358.950 ;
        RECT 165.600 358.150 165.810 358.360 ;
        RECT 171.520 358.430 171.690 358.600 ;
        RECT 205.960 358.600 206.140 358.790 ;
        RECT 170.480 358.080 170.650 358.250 ;
        RECT 183.760 358.350 183.930 358.520 ;
        RECT 188.050 358.050 188.220 358.220 ;
        RECT 184.320 357.720 184.490 357.890 ;
        RECT 185.070 357.720 185.240 357.890 ;
        RECT 187.070 357.730 187.240 357.900 ;
        RECT 188.450 358.280 188.620 358.450 ;
        RECT 188.450 357.940 188.620 358.110 ;
        RECT 216.010 359.330 216.280 359.600 ;
        RECT 224.980 359.330 225.250 359.600 ;
        RECT 234.890 360.320 235.060 360.360 ;
        RECT 235.370 360.020 235.540 360.190 ;
        RECT 232.340 359.570 232.510 359.740 ;
        RECT 233.300 359.710 233.470 359.880 ;
        RECT 233.910 359.570 234.080 359.740 ;
        RECT 234.390 359.700 234.600 359.870 ;
        RECT 234.740 359.640 234.920 359.830 ;
        RECT 236.600 359.640 236.770 359.810 ;
        RECT 233.420 359.030 233.590 359.200 ;
        RECT 207.280 358.650 207.450 358.820 ;
        RECT 212.450 358.710 212.620 358.880 ;
        RECT 212.450 358.260 212.620 358.430 ;
        RECT 228.640 358.710 228.810 358.880 ;
        RECT 214.570 358.130 214.740 358.300 ;
        RECT 228.640 358.260 228.810 358.430 ;
        RECT 205.610 357.780 205.780 357.950 ;
        RECT 164.130 357.010 164.300 357.180 ;
        RECT 207.420 357.480 207.600 357.650 ;
        RECT 171.520 357.230 171.690 357.400 ;
        RECT 165.600 356.600 165.810 356.810 ;
        RECT 233.810 358.650 233.980 358.820 ;
        RECT 234.390 358.750 234.560 358.920 ;
        RECT 233.570 358.200 233.740 358.370 ;
        RECT 232.450 357.680 232.620 357.850 ;
        RECT 171.520 356.880 171.690 357.050 ;
        RECT 170.480 356.530 170.650 356.700 ;
        RECT 192.740 356.590 192.910 356.760 ;
        RECT 213.510 356.590 213.680 356.760 ;
        RECT 190.930 356.330 191.100 356.500 ;
        RECT 191.660 356.300 191.830 356.470 ;
        RECT 214.590 356.300 214.760 356.470 ;
        RECT 192.740 356.040 192.910 356.210 ;
        RECT 213.510 356.040 213.680 356.210 ;
        RECT 193.650 355.790 193.820 355.960 ;
        RECT 197.590 355.800 197.760 355.970 ;
        RECT 208.660 355.800 208.830 355.970 ;
        RECT 212.600 355.790 212.770 355.960 ;
        RECT 215.320 356.330 215.490 356.500 ;
        RECT 217.650 356.480 217.820 356.650 ;
        RECT 217.660 355.790 217.830 355.960 ;
        RECT 223.440 356.480 223.610 356.650 ;
        RECT 223.440 355.800 223.610 355.970 ;
        RECT 190.930 354.880 191.100 355.050 ;
        RECT 192.740 355.170 192.910 355.340 ;
        RECT 213.510 355.170 213.680 355.340 ;
        RECT 191.660 354.910 191.830 355.080 ;
        RECT 214.590 354.910 214.760 355.080 ;
        RECT 215.320 354.880 215.490 355.050 ;
        RECT 2.700 353.860 4.620 354.040 ;
        RECT 192.740 354.620 192.910 354.790 ;
        RECT 193.650 354.200 193.820 354.370 ;
        RECT 197.580 354.340 197.750 354.510 ;
        RECT 213.510 354.620 213.680 354.790 ;
        RECT 2.690 353.510 4.610 353.680 ;
        RECT 193.650 353.860 193.820 354.030 ;
        RECT 195.860 353.970 196.130 354.240 ;
        RECT 197.580 354.000 197.750 354.170 ;
        RECT 192.740 353.580 192.910 353.750 ;
        RECT 199.890 354.040 200.160 354.310 ;
        RECT 206.260 354.040 206.530 354.310 ;
        RECT 208.670 354.340 208.840 354.510 ;
        RECT 208.670 354.000 208.840 354.170 ;
        RECT 210.290 353.970 210.560 354.240 ;
        RECT 212.600 354.200 212.770 354.370 ;
        RECT 214.960 354.100 215.140 354.270 ;
        RECT 212.600 353.860 212.770 354.030 ;
        RECT 213.510 353.580 213.680 353.750 ;
        RECT 2.690 353.500 3.480 353.510 ;
        RECT 235.120 358.600 235.300 358.790 ;
        RECT 236.640 358.800 236.810 358.970 ;
        RECT 234.340 358.100 234.510 358.270 ;
        RECT 235.370 358.430 235.540 358.600 ;
        RECT 235.480 357.780 235.650 357.950 ;
        RECT 234.340 357.280 234.510 357.450 ;
        RECT 236.030 357.490 236.200 357.660 ;
        RECT 235.370 356.950 235.540 357.120 ;
        RECT 234.390 356.630 234.560 356.800 ;
        RECT 233.180 356.400 233.350 356.570 ;
        RECT 236.690 356.580 236.860 356.750 ;
        RECT 233.610 355.600 233.780 355.770 ;
        RECT 234.390 355.790 234.560 355.960 ;
        RECT 236.680 355.860 236.850 356.030 ;
        RECT 235.370 355.470 235.540 355.640 ;
        RECT 234.340 355.140 234.510 355.310 ;
        RECT 236.030 354.900 236.200 355.070 ;
        RECT 234.340 354.320 234.510 354.490 ;
        RECT 235.370 353.990 235.540 354.160 ;
        RECT 234.390 353.670 234.560 353.840 ;
        RECT 364.940 354.320 365.110 365.300 ;
        RECT 365.540 354.330 365.710 365.310 ;
        RECT 366.150 354.320 366.320 365.300 ;
        RECT 366.750 354.370 366.920 365.350 ;
        RECT 367.350 354.370 367.520 365.350 ;
        RECT 367.940 354.360 368.110 365.340 ;
        RECT 368.520 354.340 368.690 365.320 ;
        RECT 369.140 354.330 369.310 365.310 ;
        RECT 369.760 354.330 369.930 365.310 ;
        RECT 371.710 359.840 371.880 360.010 ;
        RECT 372.050 359.840 372.220 360.010 ;
        RECT 372.390 359.840 372.560 360.010 ;
        RECT 372.730 359.840 372.900 360.010 ;
        RECT 236.600 353.610 236.770 353.780 ;
        RECT 190.930 353.320 191.100 353.490 ;
        RECT 183.480 352.850 183.650 353.020 ;
        RECT 184.320 352.730 184.490 352.900 ;
        RECT 185.070 352.730 185.240 352.900 ;
        RECT 2.580 351.760 3.510 351.960 ;
        RECT 2.350 348.190 2.530 351.350 ;
        RECT 5.450 350.690 8.750 351.040 ;
        RECT 0.530 338.650 0.700 338.820 ;
        RECT 0.870 338.650 1.040 338.820 ;
        RECT 1.210 338.650 1.380 338.820 ;
        RECT 1.550 338.650 1.720 338.820 ;
        RECT 4.240 340.190 4.410 349.640 ;
        RECT 4.990 340.180 5.160 349.570 ;
        RECT 5.710 340.210 5.880 349.610 ;
        RECT 6.370 340.220 6.540 349.590 ;
        RECT 7.020 340.210 7.190 349.660 ;
        RECT 7.660 340.220 7.830 349.610 ;
        RECT 164.130 351.530 164.300 351.700 ;
        RECT 171.520 351.750 171.690 351.920 ;
        RECT 188.050 352.400 188.220 352.570 ;
        RECT 183.760 352.100 183.930 352.270 ;
        RECT 188.450 352.850 188.620 353.020 ;
        RECT 191.660 353.290 191.830 353.460 ;
        RECT 214.590 353.290 214.760 353.460 ;
        RECT 192.740 353.030 192.910 353.200 ;
        RECT 213.510 353.030 213.680 353.200 ;
        RECT 215.320 353.320 215.490 353.490 ;
        RECT 370.890 354.560 371.060 354.570 ;
        RECT 368.790 353.140 370.710 353.320 ;
        RECT 188.450 352.510 188.620 352.680 ;
        RECT 368.800 352.790 370.720 352.960 ;
        RECT 369.930 352.780 370.720 352.790 ;
        RECT 370.890 352.700 371.070 354.560 ;
        RECT 190.930 351.880 191.100 352.050 ;
        RECT 192.740 352.170 192.910 352.340 ;
        RECT 213.510 352.170 213.680 352.340 ;
        RECT 191.660 351.910 191.830 352.080 ;
        RECT 214.590 351.910 214.760 352.080 ;
        RECT 215.320 351.880 215.490 352.050 ;
        RECT 165.600 351.120 165.810 351.330 ;
        RECT 171.520 351.400 171.690 351.570 ;
        RECT 170.480 351.050 170.650 351.220 ;
        RECT 192.740 351.620 192.910 351.790 ;
        RECT 213.510 351.620 213.680 351.790 ;
        RECT 183.760 351.210 183.930 351.380 ;
        RECT 188.050 350.910 188.220 351.080 ;
        RECT 164.130 349.980 164.300 350.150 ;
        RECT 184.320 350.580 184.490 350.750 ;
        RECT 185.070 350.580 185.240 350.750 ;
        RECT 187.070 350.590 187.240 350.760 ;
        RECT 188.450 351.140 188.620 351.310 ;
        RECT 188.450 350.800 188.620 350.970 ;
        RECT 369.900 351.040 370.830 351.240 ;
        RECT 171.520 350.200 171.690 350.370 ;
        RECT 165.600 349.570 165.810 349.780 ;
        RECT 171.520 349.850 171.690 350.020 ;
        RECT 183.480 349.920 183.650 350.090 ;
        RECT 170.480 349.500 170.650 349.670 ;
        RECT 184.320 349.800 184.490 349.970 ;
        RECT 185.070 349.800 185.240 349.970 ;
        RECT 164.130 348.430 164.300 348.600 ;
        RECT 188.050 349.470 188.220 349.640 ;
        RECT 183.760 349.170 183.930 349.340 ;
        RECT 188.450 349.920 188.620 350.090 ;
        RECT 188.450 349.580 188.620 349.750 ;
        RECT 171.520 348.650 171.690 348.820 ;
        RECT 165.600 348.020 165.810 348.230 ;
        RECT 171.520 348.300 171.690 348.470 ;
        RECT 170.480 347.950 170.650 348.120 ;
        RECT 183.760 348.280 183.930 348.450 ;
        RECT 188.050 347.980 188.220 348.150 ;
        RECT 184.320 347.650 184.490 347.820 ;
        RECT 185.070 347.650 185.240 347.820 ;
        RECT 187.070 347.660 187.240 347.830 ;
        RECT 188.450 348.210 188.620 348.380 ;
        RECT 188.450 347.870 188.620 348.040 ;
        RECT 164.130 346.880 164.300 347.050 ;
        RECT 171.520 347.100 171.690 347.270 ;
        RECT 193.320 347.200 193.490 347.370 ;
        RECT 165.600 346.470 165.810 346.680 ;
        RECT 171.520 346.750 171.690 346.920 ;
        RECT 191.510 346.940 191.680 347.110 ;
        RECT 170.480 346.400 170.650 346.570 ;
        RECT 192.240 346.910 192.410 347.080 ;
        RECT 193.320 346.650 193.490 346.820 ;
        RECT 194.360 346.380 194.530 346.550 ;
        RECT 191.510 345.490 191.680 345.660 ;
        RECT 198.380 346.410 198.550 346.580 ;
        RECT 193.320 345.780 193.490 345.950 ;
        RECT 192.240 345.520 192.410 345.690 ;
        RECT 193.320 345.230 193.490 345.400 ;
        RECT 194.350 345.200 194.520 345.370 ;
        RECT 194.350 344.860 194.520 345.030 ;
        RECT 198.370 345.140 198.540 345.310 ;
        RECT 194.350 344.520 194.520 344.690 ;
        RECT 141.720 344.020 141.890 344.190 ;
        RECT 142.370 344.020 142.540 344.190 ;
        RECT 193.320 344.190 193.490 344.360 ;
        RECT 196.440 344.580 196.710 344.850 ;
        RECT 198.370 344.800 198.540 344.970 ;
        RECT 198.370 344.460 198.540 344.630 ;
        RECT 200.470 344.650 200.740 344.920 ;
        RECT 140.500 343.580 140.670 343.750 ;
        RECT 141.200 343.580 141.370 343.750 ;
        RECT 140.050 341.920 140.220 342.090 ;
        RECT 191.510 343.930 191.680 344.100 ;
        RECT 192.240 343.900 192.410 344.070 ;
        RECT 193.320 343.640 193.490 343.810 ;
        RECT 142.880 343.200 143.050 343.370 ;
        RECT 204.660 343.300 204.830 343.470 ;
        RECT 142.880 342.860 143.050 343.030 ;
        RECT 183.480 343.090 183.650 343.260 ;
        RECT 184.320 342.970 184.490 343.140 ;
        RECT 185.070 342.970 185.240 343.140 ;
        RECT 143.050 341.720 143.220 341.890 ;
        RECT 164.130 341.760 164.300 341.930 ;
        RECT 171.520 341.980 171.690 342.150 ;
        RECT 188.050 342.640 188.220 342.810 ;
        RECT 183.760 342.340 183.930 342.510 ;
        RECT 188.450 343.090 188.620 343.260 ;
        RECT 188.450 342.750 188.620 342.920 ;
        RECT 191.510 342.490 191.680 342.660 ;
        RECT 193.320 342.780 193.490 342.950 ;
        RECT 192.240 342.520 192.410 342.690 ;
        RECT 204.810 342.620 204.980 342.790 ;
        RECT 206.960 342.740 207.130 342.910 ;
        RECT 193.320 342.230 193.490 342.400 ;
        RECT 205.700 342.170 205.870 342.340 ;
        RECT 165.600 341.350 165.810 341.560 ;
        RECT 171.520 341.630 171.690 341.800 ;
        RECT 143.060 341.180 143.230 341.350 ;
        RECT 170.480 341.280 170.650 341.450 ;
        RECT 204.810 341.720 204.980 341.890 ;
        RECT 183.760 341.450 183.930 341.620 ;
        RECT 188.050 341.150 188.220 341.320 ;
        RECT 140.530 339.700 140.700 339.870 ;
        RECT 142.870 340.220 143.040 340.390 ;
        RECT 164.130 340.210 164.300 340.380 ;
        RECT 184.320 340.820 184.490 340.990 ;
        RECT 185.070 340.820 185.240 340.990 ;
        RECT 187.070 340.830 187.240 341.000 ;
        RECT 188.450 341.380 188.620 341.550 ;
        RECT 206.960 341.600 207.130 341.770 ;
        RECT 188.450 341.040 188.620 341.210 ;
        RECT 204.660 341.040 204.830 341.210 ;
        RECT 171.520 340.430 171.690 340.600 ;
        RECT 204.660 340.530 204.830 340.700 ;
        RECT 141.220 339.690 141.390 339.860 ;
        RECT 165.600 339.800 165.810 340.010 ;
        RECT 171.520 340.080 171.690 340.250 ;
        RECT 183.480 340.160 183.650 340.330 ;
        RECT 170.480 339.730 170.650 339.900 ;
        RECT 184.320 340.040 184.490 340.210 ;
        RECT 185.070 340.040 185.240 340.210 ;
        RECT 141.700 338.920 141.870 339.090 ;
        RECT 142.410 338.860 142.580 339.030 ;
        RECT 164.130 338.660 164.300 338.830 ;
        RECT 188.050 339.710 188.220 339.880 ;
        RECT 183.760 339.410 183.930 339.580 ;
        RECT 188.450 340.160 188.620 340.330 ;
        RECT 188.450 339.820 188.620 339.990 ;
        RECT 204.810 339.850 204.980 340.020 ;
        RECT 206.960 339.970 207.130 340.140 ;
        RECT 205.700 339.400 205.870 339.570 ;
        RECT 171.520 338.880 171.690 339.050 ;
        RECT 0.510 331.970 0.680 332.140 ;
        RECT 0.850 331.970 1.020 332.140 ;
        RECT 1.190 331.970 1.360 332.140 ;
        RECT 1.530 331.970 1.700 332.140 ;
        RECT 2.350 326.690 2.520 326.700 ;
        RECT 2.340 324.830 2.520 326.690 ;
        RECT 3.480 326.460 3.650 337.440 ;
        RECT 4.100 326.460 4.270 337.440 ;
        RECT 4.720 326.470 4.890 337.450 ;
        RECT 5.300 326.490 5.470 337.470 ;
        RECT 5.890 326.500 6.060 337.480 ;
        RECT 6.490 326.500 6.660 337.480 ;
        RECT 7.090 326.450 7.260 337.430 ;
        RECT 7.700 326.460 7.870 337.440 ;
        RECT 8.300 326.450 8.470 337.430 ;
        RECT 165.600 338.250 165.810 338.460 ;
        RECT 171.520 338.530 171.690 338.700 ;
        RECT 193.220 338.890 193.390 339.060 ;
        RECT 204.810 338.950 204.980 339.120 ;
        RECT 142.370 338.040 142.540 338.210 ;
        RECT 170.480 338.180 170.650 338.350 ;
        RECT 183.760 338.520 183.930 338.690 ;
        RECT 188.050 338.220 188.220 338.390 ;
        RECT 139.060 337.600 139.230 337.770 ;
        RECT 140.160 337.610 140.330 337.780 ;
        RECT 139.610 336.930 139.780 337.100 ;
        RECT 139.610 335.560 139.780 335.730 ;
        RECT 139.060 334.830 139.230 335.000 ;
        RECT 139.050 333.490 139.220 333.660 ;
        RECT 141.250 337.610 141.420 337.780 ;
        RECT 140.710 336.930 140.880 337.100 ;
        RECT 140.710 335.560 140.880 335.730 ;
        RECT 140.160 334.830 140.330 335.000 ;
        RECT 140.160 333.480 140.330 333.650 ;
        RECT 139.610 332.790 139.780 332.960 ;
        RECT 184.320 337.890 184.490 338.060 ;
        RECT 185.070 337.890 185.240 338.060 ;
        RECT 187.070 337.900 187.240 338.070 ;
        RECT 188.450 338.450 188.620 338.620 ;
        RECT 188.450 338.110 188.620 338.280 ;
        RECT 206.960 338.830 207.130 339.000 ;
        RECT 204.660 338.270 204.830 338.440 ;
        RECT 193.270 338.040 193.440 338.210 ;
        RECT 364.660 349.970 367.960 350.320 ;
        RECT 365.580 339.500 365.750 348.890 ;
        RECT 366.220 339.490 366.390 348.940 ;
        RECT 366.870 339.500 367.040 348.870 ;
        RECT 367.530 339.490 367.700 348.890 ;
        RECT 368.250 339.460 368.420 348.850 ;
        RECT 369.000 339.470 369.170 348.920 ;
        RECT 370.880 347.470 371.060 350.630 ;
        RECT 142.380 337.570 142.550 337.740 ;
        RECT 141.810 336.930 141.980 337.100 ;
        RECT 164.130 337.110 164.300 337.280 ;
        RECT 142.500 336.910 142.670 337.080 ;
        RECT 171.520 337.330 171.690 337.500 ;
        RECT 142.500 336.570 142.670 336.740 ;
        RECT 165.600 336.700 165.810 336.910 ;
        RECT 171.520 336.980 171.690 337.150 ;
        RECT 371.690 337.930 371.860 338.100 ;
        RECT 372.030 337.930 372.200 338.100 ;
        RECT 372.370 337.930 372.540 338.100 ;
        RECT 372.710 337.930 372.880 338.100 ;
        RECT 170.480 336.630 170.650 336.800 ;
        RECT 142.500 336.230 142.670 336.400 ;
        RECT 141.810 335.560 141.980 335.730 ;
        RECT 141.250 334.830 141.420 335.000 ;
        RECT 141.250 333.460 141.420 333.630 ;
        RECT 140.710 332.780 140.880 332.950 ;
        RECT 149.080 333.660 149.250 334.000 ;
        RECT 149.420 333.660 149.590 334.000 ;
        RECT 141.800 332.780 141.970 332.950 ;
        RECT 141.660 330.480 141.830 330.650 ;
        RECT 138.350 330.040 138.520 330.210 ;
        RECT 139.450 330.050 139.620 330.220 ;
        RECT 140.540 330.050 140.710 330.220 ;
        RECT 138.900 329.370 139.070 329.540 ;
        RECT 140.000 329.370 140.170 329.540 ;
        RECT 138.900 328.000 139.070 328.170 ;
        RECT 140.000 328.000 140.170 328.170 ;
        RECT 141.670 330.010 141.840 330.180 ;
        RECT 141.100 329.370 141.270 329.540 ;
        RECT 141.100 328.000 141.270 328.170 ;
        RECT 172.760 331.320 172.930 331.490 ;
        RECT 173.850 331.320 174.020 331.490 ;
        RECT 173.310 330.640 173.480 330.810 ;
        RECT 173.310 329.270 173.480 329.440 ;
        RECT 176.070 331.490 176.240 331.660 ;
        RECT 174.950 331.310 175.120 331.480 ;
        RECT 176.070 331.150 176.240 331.320 ;
        RECT 176.460 331.490 176.630 331.660 ;
        RECT 176.460 331.150 176.630 331.320 ;
        RECT 177.580 331.310 177.750 331.480 ;
        RECT 178.680 331.320 178.850 331.490 ;
        RECT 174.400 330.620 174.570 330.790 ;
        RECT 175.510 330.610 175.680 330.780 ;
        RECT 177.020 330.610 177.190 330.780 ;
        RECT 178.130 330.620 178.300 330.790 ;
        RECT 174.400 329.270 174.570 329.440 ;
        RECT 175.500 329.270 175.670 329.440 ;
        RECT 177.030 329.270 177.200 329.440 ;
        RECT 178.130 329.270 178.300 329.440 ;
        RECT 179.770 331.320 179.940 331.490 ;
        RECT 179.220 330.640 179.390 330.810 ;
        RECT 179.220 329.270 179.390 329.440 ;
        RECT 182.570 331.350 182.740 331.520 ;
        RECT 183.660 331.350 183.830 331.520 ;
        RECT 183.120 330.670 183.290 330.840 ;
        RECT 183.120 329.300 183.290 329.470 ;
        RECT 185.880 331.520 186.050 331.690 ;
        RECT 184.760 331.340 184.930 331.510 ;
        RECT 185.880 331.180 186.050 331.350 ;
        RECT 186.270 331.520 186.440 331.690 ;
        RECT 186.270 331.180 186.440 331.350 ;
        RECT 187.390 331.340 187.560 331.510 ;
        RECT 188.490 331.350 188.660 331.520 ;
        RECT 184.210 330.650 184.380 330.820 ;
        RECT 185.320 330.640 185.490 330.810 ;
        RECT 186.830 330.640 187.000 330.810 ;
        RECT 187.940 330.650 188.110 330.820 ;
        RECT 184.210 329.300 184.380 329.470 ;
        RECT 185.310 329.300 185.480 329.470 ;
        RECT 186.840 329.300 187.010 329.470 ;
        RECT 187.940 329.300 188.110 329.470 ;
        RECT 189.580 331.350 189.750 331.520 ;
        RECT 189.030 330.670 189.200 330.840 ;
        RECT 189.030 329.300 189.200 329.470 ;
        RECT 193.880 331.320 194.050 331.490 ;
        RECT 193.320 330.620 193.490 330.790 ;
        RECT 193.330 329.280 193.500 329.450 ;
        RECT 138.350 327.270 138.520 327.440 ;
        RECT 139.450 327.270 139.620 327.440 ;
        RECT 2.700 325.270 4.620 325.450 ;
        RECT 138.340 325.930 138.510 326.100 ;
        RECT 139.450 325.920 139.620 326.090 ;
        RECT 2.690 324.920 4.610 325.090 ;
        RECT 137.780 325.390 137.950 325.560 ;
        RECT 138.900 325.230 139.070 325.400 ;
        RECT 140.540 327.270 140.710 327.440 ;
        RECT 140.540 325.900 140.710 326.070 ;
        RECT 140.000 325.220 140.170 325.390 ;
        RECT 2.690 324.910 3.480 324.920 ;
        RECT 141.090 325.220 141.260 325.390 ;
        RECT 172.750 328.540 172.920 328.710 ;
        RECT 172.750 327.170 172.920 327.340 ;
        RECT 172.180 326.530 172.350 326.700 ;
        RECT 173.850 328.540 174.020 328.710 ;
        RECT 174.950 328.540 175.120 328.710 ;
        RECT 177.580 328.540 177.750 328.710 ;
        RECT 178.680 328.540 178.850 328.710 ;
        RECT 173.850 327.170 174.020 327.340 ;
        RECT 174.950 327.170 175.120 327.340 ;
        RECT 177.580 327.170 177.750 327.340 ;
        RECT 178.680 327.170 178.850 327.340 ;
        RECT 173.310 326.490 173.480 326.660 ;
        RECT 174.400 326.490 174.570 326.660 ;
        RECT 175.500 326.500 175.670 326.670 ;
        RECT 177.030 326.500 177.200 326.670 ;
        RECT 178.130 326.490 178.300 326.660 ;
        RECT 179.780 328.540 179.950 328.710 ;
        RECT 179.780 327.170 179.950 327.340 ;
        RECT 179.220 326.490 179.390 326.660 ;
        RECT 180.350 326.530 180.520 326.700 ;
        RECT 182.560 328.570 182.730 328.740 ;
        RECT 182.560 327.200 182.730 327.370 ;
        RECT 181.990 326.560 182.160 326.730 ;
        RECT 183.660 328.570 183.830 328.740 ;
        RECT 184.760 328.570 184.930 328.740 ;
        RECT 187.390 328.570 187.560 328.740 ;
        RECT 188.490 328.570 188.660 328.740 ;
        RECT 183.660 327.200 183.830 327.370 ;
        RECT 184.760 327.200 184.930 327.370 ;
        RECT 187.390 327.200 187.560 327.370 ;
        RECT 188.490 327.200 188.660 327.370 ;
        RECT 172.190 326.060 172.360 326.230 ;
        RECT 180.340 326.060 180.510 326.230 ;
        RECT 183.120 326.520 183.290 326.690 ;
        RECT 184.210 326.520 184.380 326.690 ;
        RECT 185.310 326.530 185.480 326.700 ;
        RECT 186.840 326.530 187.010 326.700 ;
        RECT 187.940 326.520 188.110 326.690 ;
        RECT 189.590 328.570 189.760 328.740 ;
        RECT 189.590 327.200 189.760 327.370 ;
        RECT 189.030 326.520 189.200 326.690 ;
        RECT 190.160 326.560 190.330 326.730 ;
        RECT 194.980 331.330 195.150 331.500 ;
        RECT 194.430 330.630 194.600 330.800 ;
        RECT 194.430 329.280 194.600 329.450 ;
        RECT 193.880 328.550 194.050 328.720 ;
        RECT 193.880 327.180 194.050 327.350 ;
        RECT 182.000 326.090 182.170 326.260 ;
        RECT 193.330 326.510 193.500 326.680 ;
        RECT 196.070 331.330 196.240 331.500 ;
        RECT 195.520 330.650 195.690 330.820 ;
        RECT 195.520 329.280 195.690 329.450 ;
        RECT 194.980 328.550 195.150 328.720 ;
        RECT 194.980 327.180 195.150 327.350 ;
        RECT 194.430 326.500 194.600 326.670 ;
        RECT 196.080 328.550 196.250 328.720 ;
        RECT 196.770 328.220 196.940 328.390 ;
        RECT 196.770 327.880 196.940 328.050 ;
        RECT 196.770 327.540 196.940 327.710 ;
        RECT 196.080 327.180 196.250 327.350 ;
        RECT 195.520 326.500 195.690 326.670 ;
        RECT 196.650 326.540 196.820 326.710 ;
        RECT 190.150 326.090 190.320 326.260 ;
        RECT 196.640 326.070 196.810 326.240 ;
        RECT 2.580 323.170 3.510 323.370 ;
        RECT 2.350 319.600 2.530 322.760 ;
        RECT 5.450 322.100 8.750 322.450 ;
        RECT 0.530 310.060 0.700 310.230 ;
        RECT 0.870 310.060 1.040 310.230 ;
        RECT 1.210 310.060 1.380 310.230 ;
        RECT 1.550 310.060 1.720 310.230 ;
        RECT 4.240 311.600 4.410 321.050 ;
        RECT 4.990 311.590 5.160 320.980 ;
        RECT 5.710 311.620 5.880 321.020 ;
        RECT 6.370 311.630 6.540 321.000 ;
        RECT 7.020 311.620 7.190 321.070 ;
        RECT 7.660 311.630 7.830 321.020 ;
        RECT 143.240 321.690 143.410 325.210 ;
        RECT 143.610 321.690 143.780 325.210 ;
        RECT 143.960 321.690 144.130 325.210 ;
        RECT 144.300 321.690 144.470 325.210 ;
        RECT 144.650 321.690 144.820 325.210 ;
        RECT 145.010 321.690 145.180 325.210 ;
        RECT 145.370 321.690 145.540 325.210 ;
        RECT 222.010 323.920 222.180 324.090 ;
        RECT 227.530 323.180 227.700 323.350 ;
        RECT 222.010 322.310 222.180 322.480 ;
        RECT 227.530 322.510 227.700 322.680 ;
        RECT 222.010 320.710 222.180 320.880 ;
        RECT 222.010 319.090 222.180 319.260 ;
        RECT 224.540 317.880 224.710 318.050 ;
        RECT 222.010 317.490 222.180 317.660 ;
        RECT 222.010 315.870 222.180 316.040 ;
        RECT 222.010 314.270 222.180 314.440 ;
        RECT 233.610 314.480 233.780 329.430 ;
        RECT 364.940 325.730 365.110 336.710 ;
        RECT 365.540 325.740 365.710 336.720 ;
        RECT 366.150 325.730 366.320 336.710 ;
        RECT 366.750 325.780 366.920 336.760 ;
        RECT 367.350 325.780 367.520 336.760 ;
        RECT 367.940 325.770 368.110 336.750 ;
        RECT 368.520 325.750 368.690 336.730 ;
        RECT 369.140 325.740 369.310 336.720 ;
        RECT 369.760 325.740 369.930 336.720 ;
        RECT 371.710 331.250 371.880 331.420 ;
        RECT 372.050 331.250 372.220 331.420 ;
        RECT 372.390 331.250 372.560 331.420 ;
        RECT 372.730 331.250 372.900 331.420 ;
        RECT 370.890 325.970 371.060 325.980 ;
        RECT 368.790 324.550 370.710 324.730 ;
        RECT 368.800 324.200 370.720 324.370 ;
        RECT 369.930 324.190 370.720 324.200 ;
        RECT 370.890 324.110 371.070 325.970 ;
        RECT 369.900 322.450 370.830 322.650 ;
        RECT 222.010 312.650 222.180 312.820 ;
        RECT 0.510 303.380 0.680 303.550 ;
        RECT 0.850 303.380 1.020 303.550 ;
        RECT 1.190 303.380 1.360 303.550 ;
        RECT 1.530 303.380 1.700 303.550 ;
        RECT 2.350 298.100 2.520 298.110 ;
        RECT 2.340 296.240 2.520 298.100 ;
        RECT 3.480 297.870 3.650 308.850 ;
        RECT 4.100 297.870 4.270 308.850 ;
        RECT 4.720 297.880 4.890 308.860 ;
        RECT 5.300 297.900 5.470 308.880 ;
        RECT 5.890 297.910 6.060 308.890 ;
        RECT 6.490 297.910 6.660 308.890 ;
        RECT 7.090 297.860 7.260 308.840 ;
        RECT 7.700 297.870 7.870 308.850 ;
        RECT 8.300 297.860 8.470 308.840 ;
        RECT 364.660 321.380 367.960 321.730 ;
        RECT 365.580 310.910 365.750 320.300 ;
        RECT 366.220 310.900 366.390 320.350 ;
        RECT 366.870 310.910 367.040 320.280 ;
        RECT 367.530 310.900 367.700 320.300 ;
        RECT 368.250 310.870 368.420 320.260 ;
        RECT 369.000 310.880 369.170 320.330 ;
        RECT 370.880 318.880 371.060 322.040 ;
        RECT 371.690 309.340 371.860 309.510 ;
        RECT 372.030 309.340 372.200 309.510 ;
        RECT 372.370 309.340 372.540 309.510 ;
        RECT 372.710 309.340 372.880 309.510 ;
        RECT 2.700 296.680 4.620 296.860 ;
        RECT 364.940 297.140 365.110 308.120 ;
        RECT 365.540 297.150 365.710 308.130 ;
        RECT 366.150 297.140 366.320 308.120 ;
        RECT 366.750 297.190 366.920 308.170 ;
        RECT 367.350 297.190 367.520 308.170 ;
        RECT 367.940 297.180 368.110 308.160 ;
        RECT 368.520 297.160 368.690 308.140 ;
        RECT 369.140 297.150 369.310 308.130 ;
        RECT 369.760 297.150 369.930 308.130 ;
        RECT 371.710 302.660 371.880 302.830 ;
        RECT 372.050 302.660 372.220 302.830 ;
        RECT 372.390 302.660 372.560 302.830 ;
        RECT 372.730 302.660 372.900 302.830 ;
        RECT 2.690 296.330 4.610 296.500 ;
        RECT 2.690 296.320 3.480 296.330 ;
        RECT 370.890 297.380 371.060 297.390 ;
        RECT 368.790 295.960 370.710 296.140 ;
        RECT 368.800 295.610 370.720 295.780 ;
        RECT 369.930 295.600 370.720 295.610 ;
        RECT 370.890 295.520 371.070 297.380 ;
        RECT 2.580 294.580 3.510 294.780 ;
        RECT 2.350 291.010 2.530 294.170 ;
        RECT 5.450 293.510 8.750 293.860 ;
        RECT 0.530 281.470 0.700 281.640 ;
        RECT 0.870 281.470 1.040 281.640 ;
        RECT 1.210 281.470 1.380 281.640 ;
        RECT 1.550 281.470 1.720 281.640 ;
        RECT 4.240 283.010 4.410 292.460 ;
        RECT 4.990 283.000 5.160 292.390 ;
        RECT 5.710 283.030 5.880 292.430 ;
        RECT 6.370 283.040 6.540 292.410 ;
        RECT 7.020 283.030 7.190 292.480 ;
        RECT 7.660 283.040 7.830 292.430 ;
        RECT 0.510 274.790 0.680 274.960 ;
        RECT 0.850 274.790 1.020 274.960 ;
        RECT 1.190 274.790 1.360 274.960 ;
        RECT 1.530 274.790 1.700 274.960 ;
        RECT 2.350 269.510 2.520 269.520 ;
        RECT 2.340 267.650 2.520 269.510 ;
        RECT 3.480 269.280 3.650 280.260 ;
        RECT 4.100 269.280 4.270 280.260 ;
        RECT 4.720 269.290 4.890 280.270 ;
        RECT 5.300 269.310 5.470 280.290 ;
        RECT 5.890 269.320 6.060 280.300 ;
        RECT 6.490 269.320 6.660 280.300 ;
        RECT 7.090 269.270 7.260 280.250 ;
        RECT 7.700 269.280 7.870 280.260 ;
        RECT 8.300 269.270 8.470 280.250 ;
        RECT 369.900 293.860 370.830 294.060 ;
        RECT 364.660 292.790 367.960 293.140 ;
        RECT 365.580 282.320 365.750 291.710 ;
        RECT 366.220 282.310 366.390 291.760 ;
        RECT 366.870 282.320 367.040 291.690 ;
        RECT 367.530 282.310 367.700 291.710 ;
        RECT 368.250 282.280 368.420 291.670 ;
        RECT 369.000 282.290 369.170 291.740 ;
        RECT 370.880 290.290 371.060 293.450 ;
        RECT 371.690 280.750 371.860 280.920 ;
        RECT 372.030 280.750 372.200 280.920 ;
        RECT 372.370 280.750 372.540 280.920 ;
        RECT 372.710 280.750 372.880 280.920 ;
        RECT 2.700 268.090 4.620 268.270 ;
        RECT 364.940 268.550 365.110 279.530 ;
        RECT 365.540 268.560 365.710 279.540 ;
        RECT 366.150 268.550 366.320 279.530 ;
        RECT 366.750 268.600 366.920 279.580 ;
        RECT 367.350 268.600 367.520 279.580 ;
        RECT 367.940 268.590 368.110 279.570 ;
        RECT 368.520 268.570 368.690 279.550 ;
        RECT 369.140 268.560 369.310 279.540 ;
        RECT 369.760 268.560 369.930 279.540 ;
        RECT 371.710 274.070 371.880 274.240 ;
        RECT 372.050 274.070 372.220 274.240 ;
        RECT 372.390 274.070 372.560 274.240 ;
        RECT 372.730 274.070 372.900 274.240 ;
        RECT 2.690 267.740 4.610 267.910 ;
        RECT 2.690 267.730 3.480 267.740 ;
        RECT 370.890 268.790 371.060 268.800 ;
        RECT 368.790 267.370 370.710 267.550 ;
        RECT 368.800 267.020 370.720 267.190 ;
        RECT 369.930 267.010 370.720 267.020 ;
        RECT 370.890 266.930 371.070 268.790 ;
        RECT 2.580 265.990 3.510 266.190 ;
        RECT 2.350 262.420 2.530 265.580 ;
        RECT 5.450 264.920 8.750 265.270 ;
        RECT 0.530 252.880 0.700 253.050 ;
        RECT 0.870 252.880 1.040 253.050 ;
        RECT 1.210 252.880 1.380 253.050 ;
        RECT 1.550 252.880 1.720 253.050 ;
        RECT 4.240 254.420 4.410 263.870 ;
        RECT 4.990 254.410 5.160 263.800 ;
        RECT 5.710 254.440 5.880 263.840 ;
        RECT 6.370 254.450 6.540 263.820 ;
        RECT 7.020 254.440 7.190 263.890 ;
        RECT 7.660 254.450 7.830 263.840 ;
        RECT 0.510 246.200 0.680 246.370 ;
        RECT 0.850 246.200 1.020 246.370 ;
        RECT 1.190 246.200 1.360 246.370 ;
        RECT 1.530 246.200 1.700 246.370 ;
        RECT 2.350 240.920 2.520 240.930 ;
        RECT 2.340 239.060 2.520 240.920 ;
        RECT 3.480 240.690 3.650 251.670 ;
        RECT 4.100 240.690 4.270 251.670 ;
        RECT 4.720 240.700 4.890 251.680 ;
        RECT 5.300 240.720 5.470 251.700 ;
        RECT 5.890 240.730 6.060 251.710 ;
        RECT 6.490 240.730 6.660 251.710 ;
        RECT 7.090 240.680 7.260 251.660 ;
        RECT 7.700 240.690 7.870 251.670 ;
        RECT 8.300 240.680 8.470 251.660 ;
        RECT 369.900 265.270 370.830 265.470 ;
        RECT 364.660 264.200 367.960 264.550 ;
        RECT 365.580 253.730 365.750 263.120 ;
        RECT 366.220 253.720 366.390 263.170 ;
        RECT 366.870 253.730 367.040 263.100 ;
        RECT 367.530 253.720 367.700 263.120 ;
        RECT 368.250 253.690 368.420 263.080 ;
        RECT 369.000 253.700 369.170 263.150 ;
        RECT 370.880 261.700 371.060 264.860 ;
        RECT 371.690 252.160 371.860 252.330 ;
        RECT 372.030 252.160 372.200 252.330 ;
        RECT 372.370 252.160 372.540 252.330 ;
        RECT 372.710 252.160 372.880 252.330 ;
        RECT 2.700 239.500 4.620 239.680 ;
        RECT 364.940 239.960 365.110 250.940 ;
        RECT 365.540 239.970 365.710 250.950 ;
        RECT 366.150 239.960 366.320 250.940 ;
        RECT 366.750 240.010 366.920 250.990 ;
        RECT 367.350 240.010 367.520 250.990 ;
        RECT 367.940 240.000 368.110 250.980 ;
        RECT 368.520 239.980 368.690 250.960 ;
        RECT 369.140 239.970 369.310 250.950 ;
        RECT 369.760 239.970 369.930 250.950 ;
        RECT 371.710 245.480 371.880 245.650 ;
        RECT 372.050 245.480 372.220 245.650 ;
        RECT 372.390 245.480 372.560 245.650 ;
        RECT 372.730 245.480 372.900 245.650 ;
        RECT 2.690 239.150 4.610 239.320 ;
        RECT 2.690 239.140 3.480 239.150 ;
        RECT 370.890 240.200 371.060 240.210 ;
        RECT 368.790 238.780 370.710 238.960 ;
        RECT 368.800 238.430 370.720 238.600 ;
        RECT 369.930 238.420 370.720 238.430 ;
        RECT 370.890 238.340 371.070 240.200 ;
        RECT 2.580 237.400 3.510 237.600 ;
        RECT 2.350 233.830 2.530 236.990 ;
        RECT 5.450 236.330 8.750 236.680 ;
        RECT 0.530 224.290 0.700 224.460 ;
        RECT 0.870 224.290 1.040 224.460 ;
        RECT 1.210 224.290 1.380 224.460 ;
        RECT 1.550 224.290 1.720 224.460 ;
        RECT 4.240 225.830 4.410 235.280 ;
        RECT 4.990 225.820 5.160 235.210 ;
        RECT 5.710 225.850 5.880 235.250 ;
        RECT 6.370 225.860 6.540 235.230 ;
        RECT 7.020 225.850 7.190 235.300 ;
        RECT 7.660 225.860 7.830 235.250 ;
        RECT 0.510 217.610 0.680 217.780 ;
        RECT 0.850 217.610 1.020 217.780 ;
        RECT 1.190 217.610 1.360 217.780 ;
        RECT 1.530 217.610 1.700 217.780 ;
        RECT 2.350 212.330 2.520 212.340 ;
        RECT 2.340 210.470 2.520 212.330 ;
        RECT 3.480 212.100 3.650 223.080 ;
        RECT 4.100 212.100 4.270 223.080 ;
        RECT 4.720 212.110 4.890 223.090 ;
        RECT 5.300 212.130 5.470 223.110 ;
        RECT 5.890 212.140 6.060 223.120 ;
        RECT 6.490 212.140 6.660 223.120 ;
        RECT 7.090 212.090 7.260 223.070 ;
        RECT 7.700 212.100 7.870 223.080 ;
        RECT 8.300 212.090 8.470 223.070 ;
        RECT 369.900 236.680 370.830 236.880 ;
        RECT 364.660 235.610 367.960 235.960 ;
        RECT 365.580 225.140 365.750 234.530 ;
        RECT 366.220 225.130 366.390 234.580 ;
        RECT 366.870 225.140 367.040 234.510 ;
        RECT 367.530 225.130 367.700 234.530 ;
        RECT 368.250 225.100 368.420 234.490 ;
        RECT 369.000 225.110 369.170 234.560 ;
        RECT 370.880 233.110 371.060 236.270 ;
        RECT 371.690 223.570 371.860 223.740 ;
        RECT 372.030 223.570 372.200 223.740 ;
        RECT 372.370 223.570 372.540 223.740 ;
        RECT 372.710 223.570 372.880 223.740 ;
        RECT 2.700 210.910 4.620 211.090 ;
        RECT 364.940 211.370 365.110 222.350 ;
        RECT 365.540 211.380 365.710 222.360 ;
        RECT 366.150 211.370 366.320 222.350 ;
        RECT 366.750 211.420 366.920 222.400 ;
        RECT 367.350 211.420 367.520 222.400 ;
        RECT 367.940 211.410 368.110 222.390 ;
        RECT 368.520 211.390 368.690 222.370 ;
        RECT 369.140 211.380 369.310 222.360 ;
        RECT 369.760 211.380 369.930 222.360 ;
        RECT 371.710 216.890 371.880 217.060 ;
        RECT 372.050 216.890 372.220 217.060 ;
        RECT 372.390 216.890 372.560 217.060 ;
        RECT 372.730 216.890 372.900 217.060 ;
        RECT 2.690 210.560 4.610 210.730 ;
        RECT 2.690 210.550 3.480 210.560 ;
        RECT 370.890 211.610 371.060 211.620 ;
        RECT 368.790 210.190 370.710 210.370 ;
        RECT 368.800 209.840 370.720 210.010 ;
        RECT 369.930 209.830 370.720 209.840 ;
        RECT 370.890 209.750 371.070 211.610 ;
        RECT 2.580 208.810 3.510 209.010 ;
        RECT 2.350 205.240 2.530 208.400 ;
        RECT 5.450 207.740 8.750 208.090 ;
        RECT 0.530 195.700 0.700 195.870 ;
        RECT 0.870 195.700 1.040 195.870 ;
        RECT 1.210 195.700 1.380 195.870 ;
        RECT 1.550 195.700 1.720 195.870 ;
        RECT 4.240 197.240 4.410 206.690 ;
        RECT 4.990 197.230 5.160 206.620 ;
        RECT 5.710 197.260 5.880 206.660 ;
        RECT 6.370 197.270 6.540 206.640 ;
        RECT 7.020 197.260 7.190 206.710 ;
        RECT 7.660 197.270 7.830 206.660 ;
        RECT 0.510 189.020 0.680 189.190 ;
        RECT 0.850 189.020 1.020 189.190 ;
        RECT 1.190 189.020 1.360 189.190 ;
        RECT 1.530 189.020 1.700 189.190 ;
        RECT 2.350 183.740 2.520 183.750 ;
        RECT 2.340 181.880 2.520 183.740 ;
        RECT 3.480 183.510 3.650 194.490 ;
        RECT 4.100 183.510 4.270 194.490 ;
        RECT 4.720 183.520 4.890 194.500 ;
        RECT 5.300 183.540 5.470 194.520 ;
        RECT 5.890 183.550 6.060 194.530 ;
        RECT 6.490 183.550 6.660 194.530 ;
        RECT 7.090 183.500 7.260 194.480 ;
        RECT 7.700 183.510 7.870 194.490 ;
        RECT 8.300 183.500 8.470 194.480 ;
        RECT 369.900 208.090 370.830 208.290 ;
        RECT 364.660 207.020 367.960 207.370 ;
        RECT 365.580 196.550 365.750 205.940 ;
        RECT 366.220 196.540 366.390 205.990 ;
        RECT 366.870 196.550 367.040 205.920 ;
        RECT 367.530 196.540 367.700 205.940 ;
        RECT 368.250 196.510 368.420 205.900 ;
        RECT 369.000 196.520 369.170 205.970 ;
        RECT 370.880 204.520 371.060 207.680 ;
        RECT 371.690 194.980 371.860 195.150 ;
        RECT 372.030 194.980 372.200 195.150 ;
        RECT 372.370 194.980 372.540 195.150 ;
        RECT 372.710 194.980 372.880 195.150 ;
        RECT 2.700 182.320 4.620 182.500 ;
        RECT 364.940 182.780 365.110 193.760 ;
        RECT 365.540 182.790 365.710 193.770 ;
        RECT 366.150 182.780 366.320 193.760 ;
        RECT 366.750 182.830 366.920 193.810 ;
        RECT 367.350 182.830 367.520 193.810 ;
        RECT 367.940 182.820 368.110 193.800 ;
        RECT 368.520 182.800 368.690 193.780 ;
        RECT 369.140 182.790 369.310 193.770 ;
        RECT 369.760 182.790 369.930 193.770 ;
        RECT 371.710 188.300 371.880 188.470 ;
        RECT 372.050 188.300 372.220 188.470 ;
        RECT 372.390 188.300 372.560 188.470 ;
        RECT 372.730 188.300 372.900 188.470 ;
        RECT 2.690 181.970 4.610 182.140 ;
        RECT 2.690 181.960 3.480 181.970 ;
        RECT 370.890 183.020 371.060 183.030 ;
        RECT 368.790 181.600 370.710 181.780 ;
        RECT 368.800 181.250 370.720 181.420 ;
        RECT 369.930 181.240 370.720 181.250 ;
        RECT 370.890 181.160 371.070 183.020 ;
        RECT 2.580 180.220 3.510 180.420 ;
        RECT 2.350 176.650 2.530 179.810 ;
        RECT 5.450 179.150 8.750 179.500 ;
        RECT 0.530 167.110 0.700 167.280 ;
        RECT 0.870 167.110 1.040 167.280 ;
        RECT 1.210 167.110 1.380 167.280 ;
        RECT 1.550 167.110 1.720 167.280 ;
        RECT 4.240 168.650 4.410 178.100 ;
        RECT 4.990 168.640 5.160 178.030 ;
        RECT 5.710 168.670 5.880 178.070 ;
        RECT 6.370 168.680 6.540 178.050 ;
        RECT 7.020 168.670 7.190 178.120 ;
        RECT 7.660 168.680 7.830 178.070 ;
        RECT 0.510 160.430 0.680 160.600 ;
        RECT 0.850 160.430 1.020 160.600 ;
        RECT 1.190 160.430 1.360 160.600 ;
        RECT 1.530 160.430 1.700 160.600 ;
        RECT 2.350 155.150 2.520 155.160 ;
        RECT 2.340 153.290 2.520 155.150 ;
        RECT 3.480 154.920 3.650 165.900 ;
        RECT 4.100 154.920 4.270 165.900 ;
        RECT 4.720 154.930 4.890 165.910 ;
        RECT 5.300 154.950 5.470 165.930 ;
        RECT 5.890 154.960 6.060 165.940 ;
        RECT 6.490 154.960 6.660 165.940 ;
        RECT 7.090 154.910 7.260 165.890 ;
        RECT 7.700 154.920 7.870 165.900 ;
        RECT 8.300 154.910 8.470 165.890 ;
        RECT 2.700 153.730 4.620 153.910 ;
        RECT 2.690 153.380 4.610 153.550 ;
        RECT 2.690 153.370 3.480 153.380 ;
        RECT 2.580 151.630 3.510 151.830 ;
        RECT 2.350 148.060 2.530 151.220 ;
        RECT 5.450 150.560 8.750 150.910 ;
        RECT 0.530 138.520 0.700 138.690 ;
        RECT 0.870 138.520 1.040 138.690 ;
        RECT 1.210 138.520 1.380 138.690 ;
        RECT 1.550 138.520 1.720 138.690 ;
        RECT 4.240 140.060 4.410 149.510 ;
        RECT 4.990 140.050 5.160 149.440 ;
        RECT 5.710 140.080 5.880 149.480 ;
        RECT 6.370 140.090 6.540 149.460 ;
        RECT 7.020 140.080 7.190 149.530 ;
        RECT 7.660 140.090 7.830 149.480 ;
        RECT 0.510 131.840 0.680 132.010 ;
        RECT 0.850 131.840 1.020 132.010 ;
        RECT 1.190 131.840 1.360 132.010 ;
        RECT 1.530 131.840 1.700 132.010 ;
        RECT 2.350 126.560 2.520 126.570 ;
        RECT 2.340 124.700 2.520 126.560 ;
        RECT 3.480 126.330 3.650 137.310 ;
        RECT 4.100 126.330 4.270 137.310 ;
        RECT 4.720 126.340 4.890 137.320 ;
        RECT 5.300 126.360 5.470 137.340 ;
        RECT 5.890 126.370 6.060 137.350 ;
        RECT 6.490 126.370 6.660 137.350 ;
        RECT 7.090 126.320 7.260 137.300 ;
        RECT 7.700 126.330 7.870 137.310 ;
        RECT 8.300 126.320 8.470 137.300 ;
        RECT 2.700 125.140 4.620 125.320 ;
        RECT 2.690 124.790 4.610 124.960 ;
        RECT 2.690 124.780 3.480 124.790 ;
        RECT 2.580 123.040 3.510 123.240 ;
        RECT 2.350 119.470 2.530 122.630 ;
        RECT 5.450 121.970 8.750 122.320 ;
        RECT 0.530 109.930 0.700 110.100 ;
        RECT 0.870 109.930 1.040 110.100 ;
        RECT 1.210 109.930 1.380 110.100 ;
        RECT 1.550 109.930 1.720 110.100 ;
        RECT 4.240 111.470 4.410 120.920 ;
        RECT 4.990 111.460 5.160 120.850 ;
        RECT 5.710 111.490 5.880 120.890 ;
        RECT 6.370 111.500 6.540 120.870 ;
        RECT 7.020 111.490 7.190 120.940 ;
        RECT 7.660 111.500 7.830 120.890 ;
        RECT 0.510 103.250 0.680 103.420 ;
        RECT 0.850 103.250 1.020 103.420 ;
        RECT 1.190 103.250 1.360 103.420 ;
        RECT 1.530 103.250 1.700 103.420 ;
        RECT 2.350 97.970 2.520 97.980 ;
        RECT 2.340 96.110 2.520 97.970 ;
        RECT 3.480 97.740 3.650 108.720 ;
        RECT 4.100 97.740 4.270 108.720 ;
        RECT 4.720 97.750 4.890 108.730 ;
        RECT 5.300 97.770 5.470 108.750 ;
        RECT 5.890 97.780 6.060 108.760 ;
        RECT 6.490 97.780 6.660 108.760 ;
        RECT 7.090 97.730 7.260 108.710 ;
        RECT 7.700 97.740 7.870 108.720 ;
        RECT 8.300 97.730 8.470 108.710 ;
        RECT 2.700 96.550 4.620 96.730 ;
        RECT 2.690 96.200 4.610 96.370 ;
        RECT 2.690 96.190 3.480 96.200 ;
        RECT 2.580 94.450 3.510 94.650 ;
        RECT 2.350 90.880 2.530 94.040 ;
        RECT 5.450 93.380 8.750 93.730 ;
        RECT 0.530 81.340 0.700 81.510 ;
        RECT 0.870 81.340 1.040 81.510 ;
        RECT 1.210 81.340 1.380 81.510 ;
        RECT 1.550 81.340 1.720 81.510 ;
        RECT 4.240 82.880 4.410 92.330 ;
        RECT 4.990 82.870 5.160 92.260 ;
        RECT 5.710 82.900 5.880 92.300 ;
        RECT 6.370 82.910 6.540 92.280 ;
        RECT 7.020 82.900 7.190 92.350 ;
        RECT 7.660 82.910 7.830 92.300 ;
        RECT 0.510 74.660 0.680 74.830 ;
        RECT 0.850 74.660 1.020 74.830 ;
        RECT 1.190 74.660 1.360 74.830 ;
        RECT 1.530 74.660 1.700 74.830 ;
        RECT 2.350 69.380 2.520 69.390 ;
        RECT 2.340 67.520 2.520 69.380 ;
        RECT 3.480 69.150 3.650 80.130 ;
        RECT 4.100 69.150 4.270 80.130 ;
        RECT 4.720 69.160 4.890 80.140 ;
        RECT 5.300 69.180 5.470 80.160 ;
        RECT 5.890 69.190 6.060 80.170 ;
        RECT 6.490 69.190 6.660 80.170 ;
        RECT 7.090 69.140 7.260 80.120 ;
        RECT 7.700 69.150 7.870 80.130 ;
        RECT 8.300 69.140 8.470 80.120 ;
        RECT 2.700 67.960 4.620 68.140 ;
        RECT 2.690 67.610 4.610 67.780 ;
        RECT 2.690 67.600 3.480 67.610 ;
        RECT 2.580 65.860 3.510 66.060 ;
        RECT 2.350 62.290 2.530 65.450 ;
        RECT 5.450 64.790 8.750 65.140 ;
        RECT 0.530 52.750 0.700 52.920 ;
        RECT 0.870 52.750 1.040 52.920 ;
        RECT 1.210 52.750 1.380 52.920 ;
        RECT 1.550 52.750 1.720 52.920 ;
        RECT 4.240 54.290 4.410 63.740 ;
        RECT 4.990 54.280 5.160 63.670 ;
        RECT 5.710 54.310 5.880 63.710 ;
        RECT 6.370 54.320 6.540 63.690 ;
        RECT 7.020 54.310 7.190 63.760 ;
        RECT 7.660 54.320 7.830 63.710 ;
        RECT 0.510 46.070 0.680 46.240 ;
        RECT 0.850 46.070 1.020 46.240 ;
        RECT 1.190 46.070 1.360 46.240 ;
        RECT 1.530 46.070 1.700 46.240 ;
        RECT 2.350 40.790 2.520 40.800 ;
        RECT 2.340 38.930 2.520 40.790 ;
        RECT 3.480 40.560 3.650 51.540 ;
        RECT 4.100 40.560 4.270 51.540 ;
        RECT 4.720 40.570 4.890 51.550 ;
        RECT 5.300 40.590 5.470 51.570 ;
        RECT 5.890 40.600 6.060 51.580 ;
        RECT 6.490 40.600 6.660 51.580 ;
        RECT 7.090 40.550 7.260 51.530 ;
        RECT 7.700 40.560 7.870 51.540 ;
        RECT 8.300 40.550 8.470 51.530 ;
        RECT 2.700 39.370 4.620 39.550 ;
        RECT 2.690 39.020 4.610 39.190 ;
        RECT 2.690 39.010 3.480 39.020 ;
        RECT 2.580 37.270 3.510 37.470 ;
        RECT 2.350 33.700 2.530 36.860 ;
        RECT 5.450 36.200 8.750 36.550 ;
        RECT 0.530 24.160 0.700 24.330 ;
        RECT 0.870 24.160 1.040 24.330 ;
        RECT 1.210 24.160 1.380 24.330 ;
        RECT 1.550 24.160 1.720 24.330 ;
        RECT 4.240 25.700 4.410 35.150 ;
        RECT 4.990 25.690 5.160 35.080 ;
        RECT 5.710 25.720 5.880 35.120 ;
        RECT 6.370 25.730 6.540 35.100 ;
        RECT 7.020 25.720 7.190 35.170 ;
        RECT 7.660 25.730 7.830 35.120 ;
        RECT 0.510 17.480 0.680 17.650 ;
        RECT 0.850 17.480 1.020 17.650 ;
        RECT 1.190 17.480 1.360 17.650 ;
        RECT 1.530 17.480 1.700 17.650 ;
        RECT 2.350 12.200 2.520 12.210 ;
        RECT 2.340 10.340 2.520 12.200 ;
        RECT 3.480 11.970 3.650 22.950 ;
        RECT 4.100 11.970 4.270 22.950 ;
        RECT 4.720 11.980 4.890 22.960 ;
        RECT 5.300 12.000 5.470 22.980 ;
        RECT 5.890 12.010 6.060 22.990 ;
        RECT 6.490 12.010 6.660 22.990 ;
        RECT 7.090 11.960 7.260 22.940 ;
        RECT 7.700 11.970 7.870 22.950 ;
        RECT 8.300 11.960 8.470 22.940 ;
        RECT 2.700 10.780 4.620 10.960 ;
        RECT 2.690 10.430 4.610 10.600 ;
        RECT 2.690 10.420 3.480 10.430 ;
      LAYER met1 ;
        RECT 23.850 387.110 27.740 389.080 ;
        RECT 31.300 388.810 35.200 389.400 ;
        RECT 31.300 387.460 31.590 388.810 ;
        RECT 37.940 388.780 38.290 388.930 ;
        RECT 59.890 388.810 63.790 389.400 ;
        RECT 37.930 387.830 38.300 388.780 ;
        RECT 36.150 387.460 40.050 387.830 ;
        RECT 59.890 387.460 60.180 388.810 ;
        RECT 66.530 388.780 66.880 388.930 ;
        RECT 88.480 388.810 92.380 389.400 ;
        RECT 66.520 387.830 66.890 388.780 ;
        RECT 64.740 387.460 68.640 387.830 ;
        RECT 88.480 387.460 88.770 388.810 ;
        RECT 95.120 388.780 95.470 388.930 ;
        RECT 172.500 388.810 176.400 389.400 ;
        RECT 201.090 388.810 204.990 389.400 ;
        RECT 95.110 387.830 95.480 388.780 ;
        RECT 93.330 387.460 97.230 387.830 ;
        RECT 24.030 386.660 26.400 387.110 ;
        RECT 24.060 384.700 25.010 386.660 ;
        RECT 25.760 386.640 26.340 386.660 ;
        RECT 36.140 386.000 40.050 387.460 ;
        RECT 47.370 386.810 51.500 387.210 ;
        RECT 47.370 386.720 51.510 386.810 ;
        RECT 26.430 385.990 40.050 386.000 ;
        RECT 2.590 380.700 3.580 380.710 ;
        RECT 2.190 380.180 3.580 380.700 ;
        RECT 2.190 376.570 2.680 380.180 ;
        RECT 5.390 379.650 8.810 379.700 ;
        RECT 5.380 379.080 8.820 379.650 ;
        RECT 24.290 379.030 25.010 384.700 ;
        RECT 25.760 385.430 40.050 385.990 ;
        RECT 50.980 385.820 51.510 386.720 ;
        RECT 64.730 386.000 68.640 387.460 ;
        RECT 93.320 386.000 97.230 387.460 ;
        RECT 150.420 387.060 152.830 387.700 ;
        RECT 172.500 387.460 172.790 388.810 ;
        RECT 201.090 387.460 201.380 388.810 ;
        RECT 207.730 388.780 208.080 388.930 ;
        RECT 229.680 388.810 233.580 389.400 ;
        RECT 207.720 387.830 208.090 388.780 ;
        RECT 205.940 387.460 209.840 387.830 ;
        RECT 55.020 385.990 68.640 386.000 ;
        RECT 83.610 385.990 97.230 386.000 ;
        RECT 54.350 385.430 68.640 385.990 ;
        RECT 82.940 385.430 97.230 385.990 ;
        RECT 150.440 385.710 150.850 387.060 ;
        RECT 205.160 386.030 205.500 386.170 ;
        RECT 205.930 386.030 209.840 387.460 ;
        RECT 213.040 386.030 213.760 387.770 ;
        RECT 229.680 387.460 229.970 388.810 ;
        RECT 236.320 388.780 236.670 388.930 ;
        RECT 258.270 388.810 262.170 389.400 ;
        RECT 236.310 387.830 236.680 388.780 ;
        RECT 234.530 387.460 238.430 387.830 ;
        RECT 258.270 387.460 258.560 388.810 ;
        RECT 264.910 388.780 265.260 388.930 ;
        RECT 286.860 388.810 290.760 389.400 ;
        RECT 264.900 387.830 265.270 388.780 ;
        RECT 263.120 387.460 267.020 387.830 ;
        RECT 286.860 387.460 287.150 388.810 ;
        RECT 293.500 388.780 293.850 388.930 ;
        RECT 315.450 388.810 319.350 389.400 ;
        RECT 293.490 387.830 293.860 388.780 ;
        RECT 291.710 387.460 295.610 387.830 ;
        RECT 315.450 387.460 315.740 388.810 ;
        RECT 322.090 388.780 322.440 388.930 ;
        RECT 344.040 388.810 347.940 389.400 ;
        RECT 322.080 387.830 322.450 388.780 ;
        RECT 320.300 387.460 324.200 387.830 ;
        RECT 344.040 387.460 344.330 388.810 ;
        RECT 350.680 388.780 351.030 388.930 ;
        RECT 350.670 387.830 351.040 388.780 ;
        RECT 348.890 387.460 352.790 387.830 ;
        RECT 205.160 386.000 213.760 386.030 ;
        RECT 234.520 386.000 238.430 387.460 ;
        RECT 263.110 386.000 267.020 387.460 ;
        RECT 291.700 386.000 295.610 387.460 ;
        RECT 320.290 386.000 324.200 387.460 ;
        RECT 348.880 386.000 352.790 387.460 ;
        RECT 196.220 385.990 213.760 386.000 ;
        RECT 224.810 385.990 238.430 386.000 ;
        RECT 253.400 385.990 267.020 386.000 ;
        RECT 281.990 385.990 295.610 386.000 ;
        RECT 310.580 385.990 324.200 386.000 ;
        RECT 339.170 385.990 352.790 386.000 ;
        RECT 195.550 385.430 213.760 385.990 ;
        RECT 224.140 385.430 238.430 385.990 ;
        RECT 252.730 385.430 267.020 385.990 ;
        RECT 281.320 385.430 295.610 385.990 ;
        RECT 309.910 385.430 324.200 385.990 ;
        RECT 338.500 385.430 352.790 385.990 ;
        RECT 25.760 381.130 49.110 385.430 ;
        RECT 49.880 384.010 50.450 384.020 ;
        RECT 25.760 380.850 40.050 381.130 ;
        RECT 36.140 379.300 40.050 380.850 ;
        RECT 49.880 380.590 50.500 384.010 ;
        RECT 54.350 381.130 77.700 385.430 ;
        RECT 78.470 384.010 79.040 384.020 ;
        RECT 54.350 380.850 68.640 381.130 ;
        RECT 49.880 380.580 50.450 380.590 ;
        RECT 3.970 369.250 8.270 378.310 ;
        RECT 9.950 378.260 10.670 378.810 ;
        RECT 9.950 378.250 10.450 378.260 ;
        RECT 29.370 376.240 32.600 378.700 ;
        RECT 36.120 378.530 40.070 379.300 ;
        RECT 49.050 378.950 49.610 379.450 ;
        RECT 64.730 379.300 68.640 380.850 ;
        RECT 78.470 380.590 79.090 384.010 ;
        RECT 82.940 381.130 106.290 385.430 ;
        RECT 107.060 384.010 107.630 384.020 ;
        RECT 82.940 380.850 97.230 381.130 ;
        RECT 78.470 380.580 79.040 380.590 ;
        RECT 49.060 378.730 49.610 378.950 ;
        RECT 57.960 376.240 61.190 378.700 ;
        RECT 64.710 378.530 68.660 379.300 ;
        RECT 77.640 378.950 78.200 379.450 ;
        RECT 93.320 379.300 97.230 380.850 ;
        RECT 107.060 380.590 107.680 384.010 ;
        RECT 126.990 382.020 127.490 382.500 ;
        RECT 107.060 380.580 107.630 380.590 ;
        RECT 77.650 378.730 78.200 378.950 ;
        RECT 86.550 376.240 89.780 378.700 ;
        RECT 93.300 378.530 97.250 379.300 ;
        RECT 106.230 378.950 106.790 379.450 ;
        RECT 106.240 378.730 106.790 378.950 ;
        RECT 127.090 379.060 127.480 382.020 ;
        RECT 132.320 381.400 132.580 381.490 ;
        RECT 132.310 381.170 132.600 381.400 ;
        RECT 195.550 381.130 218.900 385.430 ;
        RECT 219.670 384.010 220.240 384.020 ;
        RECT 195.550 380.850 210.030 381.130 ;
        RECT 132.260 380.480 132.650 380.610 ;
        RECT 132.260 380.190 132.680 380.480 ;
        RECT 132.450 379.250 132.680 380.190 ;
        RECT 145.530 379.320 145.850 379.640 ;
        RECT 146.890 379.400 147.210 379.720 ;
        RECT 147.580 379.390 147.900 379.710 ;
        RECT 132.320 379.180 132.680 379.250 ;
        RECT 190.250 379.220 190.810 379.450 ;
        RECT 132.260 379.070 132.680 379.180 ;
        RECT 127.090 378.570 127.560 379.060 ;
        RECT 132.260 378.950 132.650 379.070 ;
        RECT 127.090 378.560 127.540 378.570 ;
        RECT 99.090 376.490 99.260 376.610 ;
        RECT 28.670 375.470 32.620 376.240 ;
        RECT 57.270 375.470 61.220 376.240 ;
        RECT 85.850 375.470 89.800 376.240 ;
        RECT 10.100 369.250 10.870 369.270 ;
        RECT 1.570 367.500 10.870 369.250 ;
        RECT 0.620 367.490 10.870 367.500 ;
        RECT 0.470 367.140 10.870 367.490 ;
        RECT 0.620 367.130 10.870 367.140 ;
        RECT 1.570 365.350 10.870 367.130 ;
        RECT 29.370 365.590 32.600 375.470 ;
        RECT 57.960 369.000 61.190 375.470 ;
        RECT 86.550 373.290 89.780 375.470 ;
        RECT 86.120 370.550 89.950 373.290 ;
        RECT 98.740 369.930 99.260 376.490 ;
        RECT 98.680 369.420 99.330 369.930 ;
        RECT 57.800 366.110 61.300 369.000 ;
        RECT 1.940 365.340 10.870 365.350 ;
        RECT 0.000 360.790 0.590 364.400 ;
        RECT 0.000 360.500 1.940 360.790 ;
        RECT 1.480 356.940 2.290 356.950 ;
        RECT 0.230 355.600 2.290 356.940 ;
        RECT 3.400 355.630 8.550 365.340 ;
        RECT 10.100 365.320 10.870 365.340 ;
        RECT 27.200 361.970 32.600 365.590 ;
        RECT 14.760 361.890 18.150 361.960 ;
        RECT 13.790 361.810 18.150 361.890 ;
        RECT 13.150 361.800 18.150 361.810 ;
        RECT 10.560 358.570 18.150 361.800 ;
        RECT 27.200 361.790 30.140 361.970 ;
        RECT 98.740 361.740 99.260 369.420 ;
        RECT 102.140 365.510 102.550 376.720 ;
        RECT 102.020 365.040 102.550 365.510 ;
        RECT 98.540 361.010 99.260 361.740 ;
        RECT 13.150 357.890 18.150 358.570 ;
        RECT 13.150 357.870 13.790 357.890 ;
        RECT 0.230 355.540 2.740 355.600 ;
        RECT 0.230 354.960 2.760 355.540 ;
        RECT 3.410 354.960 8.550 355.630 ;
        RECT 0.230 354.210 2.740 354.960 ;
        RECT 0.230 353.490 10.370 354.210 ;
        RECT 0.230 353.260 4.700 353.490 ;
        RECT 0.230 353.230 2.740 353.260 ;
        RECT 0.230 353.050 2.290 353.230 ;
        RECT 5.390 351.060 8.810 351.110 ;
        RECT 5.380 350.490 8.820 351.060 ;
        RECT 3.970 340.660 8.270 349.720 ;
        RECT 9.950 349.670 10.670 350.220 ;
        RECT 9.950 349.660 10.450 349.670 ;
        RECT 10.100 340.660 10.870 340.680 ;
        RECT 1.570 338.910 10.870 340.660 ;
        RECT 0.620 338.900 10.870 338.910 ;
        RECT 0.470 338.550 10.870 338.900 ;
        RECT 0.620 338.540 10.870 338.550 ;
        RECT 1.570 336.760 10.870 338.540 ;
        RECT 1.940 336.750 10.870 336.760 ;
        RECT 0.000 332.200 0.590 335.810 ;
        RECT 0.000 331.910 1.940 332.200 ;
        RECT 3.400 327.040 8.550 336.750 ;
        RECT 10.100 336.730 10.870 336.750 ;
        RECT 13.150 333.210 13.790 333.230 ;
        RECT 23.930 333.210 26.190 333.250 ;
        RECT 10.560 329.980 26.190 333.210 ;
        RECT 13.150 329.290 13.790 329.980 ;
        RECT 23.930 329.940 26.190 329.980 ;
        RECT 3.410 326.370 8.550 327.040 ;
        RECT 98.740 325.660 99.260 361.010 ;
        RECT 102.140 360.790 102.550 365.040 ;
        RECT 102.000 360.200 102.620 360.790 ;
        RECT 98.660 325.060 99.290 325.660 ;
        RECT 102.140 324.640 102.550 360.200 ;
        RECT 102.090 324.140 102.570 324.640 ;
        RECT 5.390 322.470 8.810 322.520 ;
        RECT 5.380 321.900 8.820 322.470 ;
        RECT 3.970 312.070 8.270 321.130 ;
        RECT 9.950 321.080 10.670 321.630 ;
        RECT 9.950 321.070 10.450 321.080 ;
        RECT 127.090 320.450 127.480 378.560 ;
        RECT 130.880 377.300 131.110 378.710 ;
        RECT 132.320 377.780 132.590 378.950 ;
        RECT 132.320 377.550 132.650 377.780 ;
        RECT 167.280 376.080 167.720 376.580 ;
        RECT 170.570 376.250 173.800 378.710 ;
        RECT 189.760 378.690 191.230 379.220 ;
        RECT 177.420 377.100 177.860 377.600 ;
        RECT 144.810 375.660 145.130 375.980 ;
        RECT 154.670 375.680 154.990 376.000 ;
        RECT 164.490 373.340 164.810 373.390 ;
        RECT 164.400 373.050 164.810 373.340 ;
        RECT 144.870 372.160 145.360 372.170 ;
        RECT 140.810 367.920 141.130 368.240 ;
        RECT 141.900 367.930 142.220 368.250 ;
        RECT 140.340 367.780 140.660 367.830 ;
        RECT 140.340 367.550 140.890 367.780 ;
        RECT 140.340 367.510 140.660 367.550 ;
        RECT 140.810 367.000 141.130 367.320 ;
        RECT 141.900 367.010 142.220 367.330 ;
        RECT 140.340 366.860 140.660 366.910 ;
        RECT 140.340 366.630 140.890 366.860 ;
        RECT 140.340 366.590 140.660 366.630 ;
        RECT 140.940 366.400 141.170 366.950 ;
        RECT 140.810 366.080 141.170 366.400 ;
        RECT 141.610 366.330 141.830 366.950 ;
        RECT 140.340 365.940 140.660 365.990 ;
        RECT 140.340 365.710 140.890 365.940 ;
        RECT 140.340 365.670 140.660 365.710 ;
        RECT 140.940 365.420 141.170 366.080 ;
        RECT 141.580 366.010 141.840 366.330 ;
        RECT 141.900 366.090 142.220 366.410 ;
        RECT 140.620 365.100 141.170 365.420 ;
        RECT 141.610 365.410 141.830 366.010 ;
        RECT 140.940 364.960 141.170 365.100 ;
        RECT 141.550 365.090 141.830 365.410 ;
        RECT 140.620 364.920 141.170 364.960 ;
        RECT 140.390 364.690 141.170 364.920 ;
        RECT 140.620 364.640 141.170 364.690 ;
        RECT 140.940 364.460 141.170 364.640 ;
        RECT 141.610 364.490 141.830 365.090 ;
        RECT 141.920 365.000 142.240 365.320 ;
        RECT 140.620 364.140 141.170 364.460 ;
        RECT 141.560 364.170 141.830 364.490 ;
        RECT 140.940 364.000 141.170 364.140 ;
        RECT 140.620 363.960 141.170 364.000 ;
        RECT 140.390 363.730 141.170 363.960 ;
        RECT 140.620 363.680 141.170 363.730 ;
        RECT 140.940 363.500 141.170 363.680 ;
        RECT 140.620 363.180 141.170 363.500 ;
        RECT 140.910 363.150 141.170 363.180 ;
        RECT 140.940 363.040 141.170 363.150 ;
        RECT 140.620 363.000 141.170 363.040 ;
        RECT 140.390 362.770 141.170 363.000 ;
        RECT 140.620 362.720 141.170 362.770 ;
        RECT 140.940 362.510 141.170 362.720 ;
        RECT 140.870 362.190 141.170 362.510 ;
        RECT 140.940 361.550 141.170 362.190 ;
        RECT 140.910 361.230 141.170 361.550 ;
        RECT 140.940 346.480 141.170 361.230 ;
        RECT 141.610 346.480 141.830 364.170 ;
        RECT 141.920 364.040 142.240 364.360 ;
        RECT 141.920 363.080 142.240 363.400 ;
        RECT 142.390 362.910 142.610 368.390 ;
        RECT 142.790 367.760 143.010 368.390 ;
        RECT 142.780 367.470 143.010 367.760 ;
        RECT 142.330 362.680 142.620 362.910 ;
        RECT 142.390 362.510 142.610 362.680 ;
        RECT 142.790 362.510 143.010 367.470 ;
        RECT 144.300 366.670 144.520 371.220 ;
        RECT 144.860 371.010 145.370 372.160 ;
        RECT 163.910 371.160 164.150 371.210 ;
        RECT 144.810 370.910 145.370 371.010 ;
        RECT 144.700 370.510 145.370 370.910 ;
        RECT 144.700 370.480 145.360 370.510 ;
        RECT 144.700 366.670 144.920 370.480 ;
        RECT 163.360 369.310 163.770 369.640 ;
        RECT 145.920 368.360 146.270 368.820 ;
        RECT 162.350 368.380 162.720 368.690 ;
        RECT 145.320 368.000 145.570 368.120 ;
        RECT 145.290 367.540 145.610 368.000 ;
        RECT 145.320 366.750 145.570 367.540 ;
        RECT 145.320 366.430 145.610 366.750 ;
        RECT 145.320 365.830 145.570 366.430 ;
        RECT 145.320 365.510 145.610 365.830 ;
        RECT 145.320 364.910 145.570 365.510 ;
        RECT 145.320 364.590 145.580 364.910 ;
        RECT 140.830 345.950 141.170 346.480 ;
        RECT 141.490 345.950 141.830 346.480 ;
        RECT 139.520 345.210 139.750 345.280 ;
        RECT 139.480 344.950 139.800 345.210 ;
        RECT 139.030 344.840 139.260 344.880 ;
        RECT 138.990 344.520 139.260 344.840 ;
        RECT 129.680 343.280 130.400 343.980 ;
        RECT 129.690 338.130 130.350 343.280 ;
        RECT 139.030 341.000 139.260 344.520 ;
        RECT 139.520 342.480 139.750 344.950 ;
        RECT 140.940 344.860 141.170 345.950 ;
        RECT 141.610 345.220 141.830 345.950 ;
        RECT 143.370 345.240 143.640 345.280 ;
        RECT 141.590 344.900 141.850 345.220 ;
        RECT 143.350 344.910 143.640 345.240 ;
        RECT 140.930 344.540 141.190 344.860 ;
        RECT 141.650 343.940 141.970 344.260 ;
        RECT 142.300 343.940 142.620 344.260 ;
        RECT 140.430 343.500 140.750 343.820 ;
        RECT 141.130 343.500 141.450 343.820 ;
        RECT 142.820 342.490 143.110 343.400 ;
        RECT 139.520 342.470 140.250 342.480 ;
        RECT 139.520 342.150 140.270 342.470 ;
        RECT 139.520 342.110 140.250 342.150 ;
        RECT 139.030 340.930 139.290 341.000 ;
        RECT 139.010 340.920 139.290 340.930 ;
        RECT 138.980 340.610 139.300 340.920 ;
        RECT 134.880 338.750 135.310 339.180 ;
        RECT 129.690 337.410 130.430 338.130 ;
        RECT 134.930 332.940 135.300 338.750 ;
        RECT 138.980 337.520 139.300 337.840 ;
        RECT 139.520 337.170 139.750 342.110 ;
        RECT 140.020 341.860 140.250 342.110 ;
        RECT 142.730 341.920 143.050 341.960 ;
        RECT 143.370 341.940 143.640 344.910 ;
        RECT 143.250 341.920 143.640 341.940 ;
        RECT 140.020 341.640 140.240 341.860 ;
        RECT 142.730 341.690 143.640 341.920 ;
        RECT 143.850 344.840 144.090 344.880 ;
        RECT 143.850 344.520 144.110 344.840 ;
        RECT 142.730 341.640 143.050 341.690 ;
        RECT 140.040 341.210 140.260 341.430 ;
        RECT 140.030 340.920 140.260 341.210 ;
        RECT 142.740 341.380 143.060 341.420 ;
        RECT 143.850 341.380 144.090 344.520 ;
        RECT 142.740 341.150 144.090 341.380 ;
        RECT 142.740 341.100 143.060 341.150 ;
        RECT 140.010 340.600 140.270 340.920 ;
        RECT 142.810 340.470 143.080 340.650 ;
        RECT 142.790 340.150 143.110 340.470 ;
        RECT 142.810 339.980 143.080 340.150 ;
        RECT 140.460 339.620 140.780 339.940 ;
        RECT 141.150 339.610 141.470 339.930 ;
        RECT 141.630 338.840 141.950 339.160 ;
        RECT 142.340 338.780 142.660 339.100 ;
        RECT 142.290 337.960 142.610 338.280 ;
        RECT 140.080 337.530 140.400 337.850 ;
        RECT 141.170 337.530 141.490 337.850 ;
        RECT 142.300 337.490 142.620 337.810 ;
        RECT 139.520 336.850 139.850 337.170 ;
        RECT 140.630 336.850 140.950 337.170 ;
        RECT 141.730 336.850 142.050 337.170 ;
        RECT 139.520 335.800 139.750 336.850 ;
        RECT 142.440 336.680 142.730 337.110 ;
        RECT 142.440 336.660 142.910 336.680 ;
        RECT 142.450 336.360 142.910 336.660 ;
        RECT 142.450 335.830 142.730 336.360 ;
        RECT 139.520 335.480 139.850 335.800 ;
        RECT 140.630 335.480 140.950 335.800 ;
        RECT 141.730 335.480 142.050 335.800 ;
        RECT 138.980 334.750 139.300 335.070 ;
        RECT 139.520 334.610 139.750 335.480 ;
        RECT 140.080 334.750 140.400 335.070 ;
        RECT 141.170 334.750 141.490 335.070 ;
        RECT 139.520 334.380 141.970 334.610 ;
        RECT 141.650 334.050 141.970 334.380 ;
        RECT 138.970 333.410 139.290 333.730 ;
        RECT 140.080 333.400 140.400 333.720 ;
        RECT 141.170 333.380 141.490 333.700 ;
        RECT 134.890 332.510 135.320 332.940 ;
        RECT 139.530 332.710 139.850 333.030 ;
        RECT 140.630 332.700 140.950 333.020 ;
        RECT 141.720 332.700 142.040 333.020 ;
        RECT 142.410 332.480 142.740 332.510 ;
        RECT 142.270 332.400 142.740 332.480 ;
        RECT 142.030 332.160 142.740 332.400 ;
        RECT 142.410 332.090 142.740 332.160 ;
        RECT 137.800 327.200 138.060 330.730 ;
        RECT 141.580 330.400 141.900 330.720 ;
        RECT 138.270 329.960 138.590 330.280 ;
        RECT 139.370 329.970 139.690 330.290 ;
        RECT 140.460 329.970 140.780 330.290 ;
        RECT 141.590 329.930 141.910 330.250 ;
        RECT 138.820 329.290 139.140 329.610 ;
        RECT 139.920 329.290 140.240 329.610 ;
        RECT 141.020 329.290 141.340 329.610 ;
        RECT 138.820 327.920 139.140 328.240 ;
        RECT 139.920 327.920 140.240 328.240 ;
        RECT 141.020 327.920 141.340 328.240 ;
        RECT 137.800 326.850 138.190 327.200 ;
        RECT 138.270 327.190 138.590 327.510 ;
        RECT 139.370 327.190 139.690 327.510 ;
        RECT 140.460 327.190 140.780 327.510 ;
        RECT 137.800 326.280 138.170 326.850 ;
        RECT 143.850 326.490 144.090 341.150 ;
        RECT 144.300 340.480 144.520 361.230 ;
        RECT 144.700 343.090 144.920 361.230 ;
        RECT 145.320 344.240 145.570 364.590 ;
        RECT 145.940 363.820 146.200 368.360 ;
        RECT 161.710 366.660 162.100 367.030 ;
        RECT 161.130 365.170 161.520 365.560 ;
        RECT 145.940 363.500 146.220 363.820 ;
        RECT 160.490 363.580 160.880 363.960 ;
        RECT 160.520 363.570 160.860 363.580 ;
        RECT 145.940 362.860 146.200 363.500 ;
        RECT 159.880 363.380 160.220 363.390 ;
        RECT 159.870 362.990 160.230 363.380 ;
        RECT 145.940 362.540 146.230 362.860 ;
        RECT 145.940 361.900 146.200 362.540 ;
        RECT 145.940 361.580 146.220 361.900 ;
        RECT 145.320 344.220 145.580 344.240 ;
        RECT 145.310 343.940 145.590 344.220 ;
        RECT 145.320 343.920 145.580 343.940 ;
        RECT 144.660 342.770 144.980 343.090 ;
        RECT 144.260 340.160 144.540 340.480 ;
        RECT 144.300 327.190 144.520 340.160 ;
        RECT 144.700 334.950 144.920 342.770 ;
        RECT 144.700 334.470 144.990 334.950 ;
        RECT 144.700 332.510 144.920 334.470 ;
        RECT 144.680 332.090 144.940 332.510 ;
        RECT 144.700 327.470 144.920 332.090 ;
        RECT 145.320 328.850 145.570 343.920 ;
        RECT 145.940 339.910 146.200 361.580 ;
        RECT 159.260 361.430 159.620 361.820 ;
        RECT 158.610 359.890 159.020 360.290 ;
        RECT 158.080 358.330 158.440 358.720 ;
        RECT 157.500 353.270 157.830 353.290 ;
        RECT 157.440 352.850 157.830 353.270 ;
        RECT 156.870 351.660 157.200 351.680 ;
        RECT 156.820 351.270 157.210 351.660 ;
        RECT 156.250 350.110 156.580 350.120 ;
        RECT 156.220 349.720 156.580 350.110 ;
        RECT 155.600 348.240 155.990 348.640 ;
        RECT 154.930 343.070 155.360 343.470 ;
        RECT 154.270 341.500 154.680 341.900 ;
        RECT 145.930 339.590 146.240 339.910 ;
        RECT 153.660 339.860 154.050 340.260 ;
        RECT 145.280 328.450 145.580 328.850 ;
        RECT 144.700 327.330 144.940 327.470 ;
        RECT 144.260 326.840 144.570 327.190 ;
        RECT 144.710 326.700 144.940 327.330 ;
        RECT 137.800 325.750 138.060 326.280 ;
        RECT 138.260 325.850 138.580 326.170 ;
        RECT 139.370 325.840 139.690 326.160 ;
        RECT 140.460 325.820 140.780 326.140 ;
        RECT 143.060 325.930 144.090 326.490 ;
        RECT 144.700 326.670 144.940 326.700 ;
        RECT 143.060 325.820 143.850 325.930 ;
        RECT 137.750 324.940 138.060 325.750 ;
        RECT 138.820 325.150 139.140 325.470 ;
        RECT 139.920 325.140 140.240 325.460 ;
        RECT 141.010 325.140 141.330 325.460 ;
        RECT 144.700 325.280 144.920 326.670 ;
        RECT 137.800 324.740 138.060 324.940 ;
        RECT 143.170 321.600 145.590 325.280 ;
        RECT 145.940 321.310 146.200 339.590 ;
        RECT 152.970 338.420 153.380 338.810 ;
        RECT 148.760 333.270 149.690 334.920 ;
        RECT 148.850 332.790 149.590 333.270 ;
        RECT 145.850 320.900 146.200 321.310 ;
        RECT 126.920 319.930 127.480 320.450 ;
        RECT 153.030 315.080 153.360 338.420 ;
        RECT 152.980 315.070 153.410 315.080 ;
        RECT 152.950 314.610 153.440 315.070 ;
        RECT 152.980 314.590 153.410 314.610 ;
        RECT 153.680 314.290 154.010 339.860 ;
        RECT 153.590 313.800 154.080 314.290 ;
        RECT 154.330 313.580 154.660 341.500 ;
        RECT 154.300 313.120 154.700 313.580 ;
        RECT 154.090 312.630 154.670 312.740 ;
        RECT 155.000 312.630 155.330 343.070 ;
        RECT 155.640 317.210 155.970 348.240 ;
        RECT 155.640 312.750 155.960 317.210 ;
        RECT 156.250 313.360 156.580 349.720 ;
        RECT 156.870 313.610 157.200 351.270 ;
        RECT 157.500 314.640 157.830 352.850 ;
        RECT 158.100 314.940 158.430 358.330 ;
        RECT 158.680 315.510 159.010 359.890 ;
        RECT 159.290 316.540 159.620 361.430 ;
        RECT 159.880 317.150 160.210 362.990 ;
        RECT 160.520 317.820 160.850 363.570 ;
        RECT 161.140 318.470 161.470 365.170 ;
        RECT 161.740 319.100 162.070 366.660 ;
        RECT 162.370 319.710 162.700 368.380 ;
        RECT 163.360 367.760 163.770 368.090 ;
        RECT 163.360 366.210 163.770 366.540 ;
        RECT 164.100 365.020 164.340 370.810 ;
        RECT 164.400 369.550 164.640 373.050 ;
        RECT 166.850 371.140 167.160 371.210 ;
        RECT 167.340 370.810 167.650 376.080 ;
        RECT 169.870 375.480 173.820 376.250 ;
        RECT 170.570 372.480 173.800 375.480 ;
        RECT 171.280 371.160 171.570 371.210 ;
        RECT 165.520 370.170 165.870 370.460 ;
        RECT 165.520 370.150 165.720 370.170 ;
        RECT 167.040 369.750 167.650 370.810 ;
        RECT 170.400 370.270 170.720 370.570 ;
        RECT 167.040 369.480 167.880 369.750 ;
        RECT 165.520 368.620 165.870 368.910 ;
        RECT 165.520 368.600 165.720 368.620 ;
        RECT 165.520 367.070 165.870 367.360 ;
        RECT 165.520 367.050 165.720 367.070 ;
        RECT 165.520 365.520 165.870 365.810 ;
        RECT 165.520 365.500 165.720 365.520 ;
        RECT 167.040 365.030 167.350 369.480 ;
        RECT 167.600 369.420 167.880 369.480 ;
        RECT 170.400 368.720 170.720 369.020 ;
        RECT 167.600 367.870 167.880 368.200 ;
        RECT 170.400 367.170 170.720 367.470 ;
        RECT 167.600 366.320 167.880 366.650 ;
        RECT 170.400 365.620 170.720 365.920 ;
        RECT 163.360 364.660 163.770 364.990 ;
        RECT 163.910 364.970 164.340 365.020 ;
        RECT 166.850 364.970 167.350 365.030 ;
        RECT 164.100 364.570 164.340 364.970 ;
        RECT 167.040 364.570 167.350 364.970 ;
        RECT 167.600 364.770 167.880 365.100 ;
        RECT 171.470 365.020 171.760 370.810 ;
        RECT 171.770 369.500 172.060 372.480 ;
        RECT 171.280 364.970 171.760 365.020 ;
        RECT 171.470 364.570 171.760 364.970 ;
        RECT 167.640 363.550 167.650 363.560 ;
        RECT 164.400 363.470 164.640 363.550 ;
        RECT 167.340 363.470 167.650 363.550 ;
        RECT 171.770 363.470 172.060 363.550 ;
        RECT 173.230 363.110 173.420 372.480 ;
        RECT 177.510 363.070 177.760 377.100 ;
        RECT 182.210 376.630 182.820 376.770 ;
        RECT 182.190 374.670 183.370 376.630 ;
        RECT 181.390 373.760 183.370 374.670 ;
        RECT 181.390 373.580 183.200 373.760 ;
        RECT 186.630 373.600 187.350 377.460 ;
        RECT 187.390 376.080 187.830 376.580 ;
        RECT 181.390 372.890 182.120 373.580 ;
        RECT 181.590 372.330 181.930 372.620 ;
        RECT 181.640 372.300 181.900 372.330 ;
        RECT 179.760 368.770 180.020 369.090 ;
        RECT 179.790 366.540 179.980 368.770 ;
        RECT 181.660 366.520 181.870 372.300 ;
        RECT 185.230 371.700 185.490 371.710 ;
        RECT 185.210 371.400 185.510 371.700 ;
        RECT 185.230 371.390 185.490 371.400 ;
        RECT 182.060 370.370 182.400 370.690 ;
        RECT 182.130 366.540 182.320 370.370 ;
        RECT 182.500 368.280 182.790 368.600 ;
        RECT 182.540 366.520 182.750 368.280 ;
        RECT 183.540 367.800 183.880 368.120 ;
        RECT 183.620 366.550 183.800 367.800 ;
        RECT 185.260 363.370 185.460 371.390 ;
        RECT 187.490 366.500 187.720 376.080 ;
        RECT 188.390 372.310 188.670 372.630 ;
        RECT 187.950 371.400 188.230 371.720 ;
        RECT 183.730 363.150 183.920 363.370 ;
        RECT 183.450 362.660 183.920 363.150 ;
        RECT 184.310 363.010 184.680 363.030 ;
        RECT 184.260 362.750 184.680 363.010 ;
        RECT 184.310 362.740 184.680 362.750 ;
        RECT 163.360 362.030 163.770 362.360 ;
        RECT 164.100 362.050 164.340 362.450 ;
        RECT 167.040 362.050 167.350 362.450 ;
        RECT 163.910 362.000 164.340 362.050 ;
        RECT 163.360 360.480 163.770 360.810 ;
        RECT 163.360 358.930 163.770 359.260 ;
        RECT 163.360 357.380 163.770 357.710 ;
        RECT 164.100 356.210 164.340 362.000 ;
        RECT 166.850 361.990 167.350 362.050 ;
        RECT 165.520 361.500 165.720 361.520 ;
        RECT 165.520 361.210 165.870 361.500 ;
        RECT 165.520 359.950 165.720 359.970 ;
        RECT 165.520 359.660 165.870 359.950 ;
        RECT 165.520 358.400 165.720 358.420 ;
        RECT 165.520 358.110 165.870 358.400 ;
        RECT 167.040 357.540 167.350 361.990 ;
        RECT 167.600 361.920 167.880 362.250 ;
        RECT 171.470 362.050 171.760 362.450 ;
        RECT 183.270 362.220 183.590 362.500 ;
        RECT 183.730 362.400 183.920 362.660 ;
        RECT 171.280 362.000 171.760 362.050 ;
        RECT 170.400 361.100 170.720 361.400 ;
        RECT 167.600 360.370 167.880 360.700 ;
        RECT 170.400 359.550 170.720 359.850 ;
        RECT 167.600 358.820 167.880 359.150 ;
        RECT 170.400 358.000 170.720 358.300 ;
        RECT 167.600 357.540 167.880 357.600 ;
        RECT 163.910 355.810 164.150 355.860 ;
        RECT 164.400 353.100 164.640 357.470 ;
        RECT 167.040 357.270 167.880 357.540 ;
        RECT 165.520 356.850 165.720 356.870 ;
        RECT 165.520 356.560 165.870 356.850 ;
        RECT 167.040 356.210 167.650 357.270 ;
        RECT 170.400 356.450 170.720 356.750 ;
        RECT 171.470 356.210 171.760 362.000 ;
        RECT 183.730 362.110 183.960 362.400 ;
        RECT 183.730 361.510 183.920 362.110 ;
        RECT 183.270 361.120 183.590 361.400 ;
        RECT 183.730 361.220 183.960 361.510 ;
        RECT 183.730 360.960 183.920 361.220 ;
        RECT 183.450 360.470 183.920 360.960 ;
        RECT 185.040 361.030 185.460 363.370 ;
        RECT 187.980 363.370 188.200 371.400 ;
        RECT 187.980 363.150 188.260 363.370 ;
        RECT 188.410 363.150 188.640 372.310 ;
        RECT 189.780 366.310 190.200 378.690 ;
        RECT 190.810 366.310 191.230 378.690 ;
        RECT 193.190 376.040 193.630 376.540 ;
        RECT 197.710 376.240 198.990 380.850 ;
        RECT 199.160 376.240 202.390 378.700 ;
        RECT 193.290 369.060 193.520 376.040 ;
        RECT 197.710 375.470 202.410 376.240 ;
        RECT 197.710 370.790 198.990 375.470 ;
        RECT 199.160 372.480 202.390 375.470 ;
        RECT 197.710 370.710 199.010 370.790 ;
        RECT 197.700 370.410 199.010 370.710 ;
        RECT 194.480 369.760 194.780 370.080 ;
        RECT 193.160 369.050 193.520 369.060 ;
        RECT 193.130 368.200 193.520 369.050 ;
        RECT 193.160 368.190 193.520 368.200 ;
        RECT 193.290 366.500 193.520 368.190 ;
        RECT 194.510 366.500 194.740 369.760 ;
        RECT 200.790 369.210 201.220 369.550 ;
        RECT 201.030 366.540 201.220 369.210 ;
        RECT 201.470 366.450 201.750 372.480 ;
        RECT 203.170 372.310 203.430 372.630 ;
        RECT 202.280 371.440 202.540 371.760 ;
        RECT 202.310 367.720 202.500 371.440 ;
        RECT 203.190 367.720 203.410 372.310 ;
        RECT 205.160 369.090 205.500 380.850 ;
        RECT 205.930 379.300 210.030 380.850 ;
        RECT 219.670 380.590 220.290 384.010 ;
        RECT 224.140 381.130 247.490 385.430 ;
        RECT 248.260 384.010 248.830 384.020 ;
        RECT 224.140 380.850 238.430 381.130 ;
        RECT 219.670 380.580 220.240 380.590 ;
        RECT 205.910 378.530 210.030 379.300 ;
        RECT 218.840 378.950 219.400 379.450 ;
        RECT 218.850 378.730 219.400 378.950 ;
        RECT 205.810 372.990 206.130 373.360 ;
        RECT 205.830 369.150 206.100 372.990 ;
        RECT 205.110 369.010 205.500 369.090 ;
        RECT 205.100 368.240 205.500 369.010 ;
        RECT 205.110 368.170 205.500 368.240 ;
        RECT 202.140 367.030 202.820 367.720 ;
        RECT 203.180 367.030 203.860 367.720 ;
        RECT 205.160 366.390 205.500 368.170 ;
        RECT 205.550 368.500 205.710 369.150 ;
        RECT 205.550 367.950 205.820 368.500 ;
        RECT 205.540 367.900 205.820 367.950 ;
        RECT 205.540 367.810 205.710 367.900 ;
        RECT 205.550 364.440 205.710 367.810 ;
        RECT 205.830 367.660 206.150 369.150 ;
        RECT 207.830 368.780 208.040 369.150 ;
        RECT 207.360 368.330 207.670 368.770 ;
        RECT 207.820 368.490 208.050 368.780 ;
        RECT 205.830 367.610 206.170 367.660 ;
        RECT 205.830 367.110 206.510 367.610 ;
        RECT 205.830 366.460 206.120 367.110 ;
        RECT 206.960 366.800 207.280 367.120 ;
        RECT 207.830 366.790 208.040 368.490 ;
        RECT 208.300 368.220 208.490 369.150 ;
        RECT 208.290 367.930 208.520 368.220 ;
        RECT 205.960 365.110 206.120 366.460 ;
        RECT 206.310 366.290 206.550 366.710 ;
        RECT 207.820 366.500 208.050 366.790 ;
        RECT 207.830 366.360 208.040 366.500 ;
        RECT 206.280 365.970 206.550 366.290 ;
        RECT 206.310 365.540 206.550 365.970 ;
        RECT 208.300 365.900 208.490 367.930 ;
        RECT 208.710 366.430 208.920 369.150 ;
        RECT 208.680 365.920 208.920 366.430 ;
        RECT 207.850 365.720 208.040 365.850 ;
        RECT 207.830 365.430 208.060 365.720 ;
        RECT 208.290 365.610 208.520 365.900 ;
        RECT 206.950 365.110 207.270 365.430 ;
        RECT 205.930 364.870 206.160 365.110 ;
        RECT 205.920 364.860 206.160 364.870 ;
        RECT 205.920 364.590 206.170 364.860 ;
        RECT 205.930 364.560 206.150 364.590 ;
        RECT 205.540 364.350 205.710 364.440 ;
        RECT 205.540 364.300 205.820 364.350 ;
        RECT 205.550 363.750 205.820 364.300 ;
        RECT 186.770 362.990 187.110 363.040 ;
        RECT 186.770 362.970 187.330 362.990 ;
        RECT 186.650 362.800 187.330 362.970 ;
        RECT 186.770 362.760 187.330 362.800 ;
        RECT 186.770 362.720 187.110 362.760 ;
        RECT 187.980 362.080 188.650 363.150 ;
        RECT 205.550 363.120 205.710 363.750 ;
        RECT 205.430 362.470 205.710 363.120 ;
        RECT 187.980 361.540 188.260 362.080 ;
        RECT 188.410 361.540 188.640 362.080 ;
        RECT 205.430 361.870 205.820 362.470 ;
        RECT 184.310 360.870 184.680 360.880 ;
        RECT 184.260 360.610 184.680 360.870 ;
        RECT 184.310 360.590 184.680 360.610 ;
        RECT 185.040 360.700 185.520 361.030 ;
        RECT 186.770 360.860 187.110 360.900 ;
        RECT 186.770 360.820 187.330 360.860 ;
        RECT 183.730 360.220 183.920 360.470 ;
        RECT 183.450 359.730 183.920 360.220 ;
        RECT 184.310 360.080 184.680 360.100 ;
        RECT 184.260 359.820 184.680 360.080 ;
        RECT 184.310 359.810 184.680 359.820 ;
        RECT 183.270 359.290 183.590 359.570 ;
        RECT 183.730 359.470 183.920 359.730 ;
        RECT 183.730 359.180 183.960 359.470 ;
        RECT 183.730 358.580 183.920 359.180 ;
        RECT 183.270 358.190 183.590 358.470 ;
        RECT 183.730 358.290 183.960 358.580 ;
        RECT 183.730 358.030 183.920 358.290 ;
        RECT 183.450 357.540 183.920 358.030 ;
        RECT 184.310 357.940 184.680 357.950 ;
        RECT 184.260 357.680 184.680 357.940 ;
        RECT 184.310 357.660 184.680 357.680 ;
        RECT 166.850 355.810 167.160 355.880 ;
        RECT 167.340 353.030 167.650 356.210 ;
        RECT 171.280 355.810 171.570 355.860 ;
        RECT 171.770 353.050 172.060 357.520 ;
        RECT 173.230 353.060 173.420 357.460 ;
        RECT 174.540 353.250 174.770 357.500 ;
        RECT 177.510 353.250 177.760 357.520 ;
        RECT 183.730 357.320 183.920 357.540 ;
        RECT 185.040 357.320 185.270 360.700 ;
        RECT 186.650 360.650 187.330 360.820 ;
        RECT 186.770 360.630 187.330 360.650 ;
        RECT 186.770 360.580 187.110 360.630 ;
        RECT 187.980 360.470 188.650 361.540 ;
        RECT 187.980 360.220 188.260 360.470 ;
        RECT 188.410 360.220 188.640 360.470 ;
        RECT 186.770 360.060 187.110 360.110 ;
        RECT 186.770 360.040 187.330 360.060 ;
        RECT 186.650 359.870 187.330 360.040 ;
        RECT 186.770 359.830 187.330 359.870 ;
        RECT 187.980 359.860 188.650 360.220 ;
        RECT 186.770 359.790 187.110 359.830 ;
        RECT 187.970 359.790 188.650 359.860 ;
        RECT 187.960 359.190 188.650 359.790 ;
        RECT 187.970 359.160 188.650 359.190 ;
        RECT 187.980 359.150 188.650 359.160 ;
        RECT 187.980 358.610 188.260 359.150 ;
        RECT 186.770 357.930 187.110 357.970 ;
        RECT 186.770 357.890 187.330 357.930 ;
        RECT 186.650 357.720 187.330 357.890 ;
        RECT 186.770 357.700 187.330 357.720 ;
        RECT 186.770 357.650 187.110 357.700 ;
        RECT 187.980 357.540 188.650 358.610 ;
        RECT 205.430 358.320 205.710 361.870 ;
        RECT 205.960 361.660 206.150 364.560 ;
        RECT 207.360 363.480 207.670 363.920 ;
        RECT 207.850 363.810 208.040 365.430 ;
        RECT 208.300 364.320 208.490 365.610 ;
        RECT 208.280 364.030 208.510 364.320 ;
        RECT 207.850 363.600 208.080 363.810 ;
        RECT 207.840 363.520 208.080 363.600 ;
        RECT 207.840 363.100 208.070 363.520 ;
        RECT 208.300 363.100 208.490 364.030 ;
        RECT 208.710 363.100 208.920 365.920 ;
        RECT 209.660 365.330 210.030 378.530 ;
        RECT 226.650 378.700 227.930 380.850 ;
        RECT 234.520 379.300 238.430 380.850 ;
        RECT 248.260 380.590 248.880 384.010 ;
        RECT 252.730 381.130 276.080 385.430 ;
        RECT 276.850 384.010 277.420 384.020 ;
        RECT 252.730 380.850 267.020 381.130 ;
        RECT 248.260 380.580 248.830 380.590 ;
        RECT 210.450 377.950 210.910 378.380 ;
        RECT 209.500 365.310 210.100 365.330 ;
        RECT 209.340 365.270 210.100 365.310 ;
        RECT 209.340 365.010 210.030 365.270 ;
        RECT 207.360 362.300 207.670 362.740 ;
        RECT 205.930 361.630 206.150 361.660 ;
        RECT 205.920 361.360 206.170 361.630 ;
        RECT 205.920 361.350 206.160 361.360 ;
        RECT 205.930 361.110 206.160 361.350 ;
        RECT 207.200 361.340 207.520 361.660 ;
        RECT 205.960 359.080 206.120 361.110 ;
        RECT 206.310 360.550 206.550 360.680 ;
        RECT 206.290 360.230 206.550 360.550 ;
        RECT 206.290 359.630 206.550 359.950 ;
        RECT 206.310 359.510 206.550 359.630 ;
        RECT 209.660 359.300 210.030 365.010 ;
        RECT 209.390 359.240 210.110 359.300 ;
        RECT 205.930 358.840 206.160 359.080 ;
        RECT 209.390 358.970 210.030 359.240 ;
        RECT 205.920 358.830 206.160 358.840 ;
        RECT 205.920 358.560 206.170 358.830 ;
        RECT 207.200 358.580 207.520 358.900 ;
        RECT 205.930 358.530 206.150 358.560 ;
        RECT 205.430 357.720 205.820 358.320 ;
        RECT 187.980 357.320 188.260 357.540 ;
        RECT 187.980 355.960 188.200 357.320 ;
        RECT 190.870 356.560 191.030 357.210 ;
        RECT 190.870 356.010 191.140 356.560 ;
        RECT 190.860 355.960 191.140 356.010 ;
        RECT 191.280 356.220 191.470 357.210 ;
        RECT 191.680 356.530 191.840 357.210 ;
        RECT 191.640 356.510 191.840 356.530 ;
        RECT 192.660 356.520 192.980 356.840 ;
        RECT 191.630 356.270 191.860 356.510 ;
        RECT 191.280 356.100 191.450 356.220 ;
        RECT 187.980 355.870 188.330 355.960 ;
        RECT 190.860 355.870 191.030 355.960 ;
        RECT 187.980 355.650 188.490 355.870 ;
        RECT 190.870 355.510 191.030 355.870 ;
        RECT 190.860 355.420 191.030 355.510 ;
        RECT 190.860 355.370 191.140 355.420 ;
        RECT 190.870 355.070 191.140 355.370 ;
        RECT 191.280 355.280 191.440 356.100 ;
        RECT 191.640 356.050 191.840 356.270 ;
        RECT 191.680 355.330 191.840 356.050 ;
        RECT 192.660 355.970 192.980 356.290 ;
        RECT 193.620 356.050 193.860 357.210 ;
        RECT 191.280 355.160 191.450 355.280 ;
        RECT 179.270 353.820 179.550 354.930 ;
        RECT 179.800 354.240 179.990 354.840 ;
        RECT 181.800 354.400 182.190 354.420 ;
        RECT 181.790 354.310 182.190 354.400 ;
        RECT 179.800 354.050 181.430 354.240 ;
        RECT 179.270 353.540 180.990 353.820 ;
        RECT 180.710 353.310 180.990 353.540 ;
        RECT 181.240 353.270 181.430 354.050 ;
        RECT 181.640 354.060 182.190 354.310 ;
        RECT 181.640 354.040 182.180 354.060 ;
        RECT 181.640 353.190 181.800 354.040 ;
        RECT 185.760 353.970 186.140 353.990 ;
        RECT 186.280 353.970 186.510 354.880 ;
        RECT 185.760 353.740 186.510 353.970 ;
        RECT 187.500 353.880 187.730 354.880 ;
        RECT 190.810 353.890 191.230 355.070 ;
        RECT 191.280 354.300 191.470 355.160 ;
        RECT 191.640 355.110 191.840 355.330 ;
        RECT 191.630 354.870 191.860 355.110 ;
        RECT 192.660 355.090 192.980 355.410 ;
        RECT 193.610 355.390 193.880 356.050 ;
        RECT 191.640 354.850 191.840 354.870 ;
        RECT 191.250 354.070 191.490 354.300 ;
        RECT 183.730 353.080 183.920 353.300 ;
        RECT 183.450 352.590 183.920 353.080 ;
        RECT 184.310 352.940 184.680 352.960 ;
        RECT 184.260 352.680 184.680 352.940 ;
        RECT 184.310 352.670 184.680 352.680 ;
        RECT 163.360 351.900 163.770 352.230 ;
        RECT 164.100 351.920 164.340 352.320 ;
        RECT 167.040 351.920 167.350 352.320 ;
        RECT 163.910 351.870 164.340 351.920 ;
        RECT 163.360 350.350 163.770 350.680 ;
        RECT 163.360 348.800 163.770 349.130 ;
        RECT 163.360 347.250 163.770 347.580 ;
        RECT 164.100 346.080 164.340 351.870 ;
        RECT 166.850 351.860 167.350 351.920 ;
        RECT 165.520 351.370 165.720 351.390 ;
        RECT 165.520 351.080 165.870 351.370 ;
        RECT 165.520 349.820 165.720 349.840 ;
        RECT 165.520 349.530 165.870 349.820 ;
        RECT 165.520 348.270 165.720 348.290 ;
        RECT 165.520 347.980 165.870 348.270 ;
        RECT 167.040 347.410 167.350 351.860 ;
        RECT 167.600 351.790 167.880 352.120 ;
        RECT 171.470 351.920 171.760 352.320 ;
        RECT 183.270 352.150 183.590 352.430 ;
        RECT 183.730 352.330 183.920 352.590 ;
        RECT 171.280 351.870 171.760 351.920 ;
        RECT 170.400 350.970 170.720 351.270 ;
        RECT 167.600 350.240 167.880 350.570 ;
        RECT 170.400 349.420 170.720 349.720 ;
        RECT 167.600 348.690 167.880 349.020 ;
        RECT 170.400 347.870 170.720 348.170 ;
        RECT 167.600 347.410 167.880 347.470 ;
        RECT 163.910 345.680 164.150 345.730 ;
        RECT 164.400 343.570 164.640 347.340 ;
        RECT 167.040 347.140 167.880 347.410 ;
        RECT 165.520 346.720 165.720 346.740 ;
        RECT 165.520 346.430 165.870 346.720 ;
        RECT 167.040 346.080 167.650 347.140 ;
        RECT 170.400 346.320 170.720 346.620 ;
        RECT 171.470 346.080 171.760 351.870 ;
        RECT 183.730 352.040 183.960 352.330 ;
        RECT 183.730 351.440 183.920 352.040 ;
        RECT 183.270 351.050 183.590 351.330 ;
        RECT 183.730 351.150 183.960 351.440 ;
        RECT 183.730 350.890 183.920 351.150 ;
        RECT 183.450 350.400 183.920 350.890 ;
        RECT 184.310 350.800 184.680 350.810 ;
        RECT 184.260 350.540 184.680 350.800 ;
        RECT 184.310 350.520 184.680 350.540 ;
        RECT 183.730 350.150 183.920 350.400 ;
        RECT 183.450 349.660 183.920 350.150 ;
        RECT 184.310 350.010 184.680 350.030 ;
        RECT 184.260 349.750 184.680 350.010 ;
        RECT 184.310 349.740 184.680 349.750 ;
        RECT 183.270 349.220 183.590 349.500 ;
        RECT 183.730 349.400 183.920 349.660 ;
        RECT 183.730 349.110 183.960 349.400 ;
        RECT 183.730 348.510 183.920 349.110 ;
        RECT 183.270 348.120 183.590 348.400 ;
        RECT 183.730 348.220 183.960 348.510 ;
        RECT 183.730 347.960 183.920 348.220 ;
        RECT 183.450 347.470 183.920 347.960 ;
        RECT 184.310 347.870 184.680 347.880 ;
        RECT 184.260 347.610 184.680 347.870 ;
        RECT 184.310 347.590 184.680 347.610 ;
        RECT 166.850 345.680 167.160 345.750 ;
        RECT 167.340 343.570 167.650 346.080 ;
        RECT 171.280 345.680 171.570 345.730 ;
        RECT 171.770 343.570 172.060 347.390 ;
        RECT 173.230 343.300 173.420 347.390 ;
        RECT 174.540 346.350 174.770 347.430 ;
        RECT 174.450 345.870 174.780 346.350 ;
        RECT 174.540 343.260 174.770 345.870 ;
        RECT 177.510 343.470 177.760 347.450 ;
        RECT 180.830 343.410 180.990 347.460 ;
        RECT 183.580 347.250 183.920 347.470 ;
        RECT 185.040 347.250 185.270 353.300 ;
        RECT 185.760 352.970 186.140 353.740 ;
        RECT 187.500 353.580 187.750 353.880 ;
        RECT 187.510 353.110 187.750 353.580 ;
        RECT 190.810 353.500 191.270 353.890 ;
        RECT 188.010 353.080 188.260 353.300 ;
        RECT 186.770 352.920 187.110 352.970 ;
        RECT 186.770 352.900 187.330 352.920 ;
        RECT 186.650 352.730 187.330 352.900 ;
        RECT 186.770 352.690 187.330 352.730 ;
        RECT 186.770 352.650 187.110 352.690 ;
        RECT 188.010 352.010 188.650 353.080 ;
        RECT 190.870 353.000 191.270 353.500 ;
        RECT 190.860 352.950 191.270 353.000 ;
        RECT 191.280 353.210 191.470 354.070 ;
        RECT 191.680 353.520 191.840 354.850 ;
        RECT 192.660 354.540 192.980 354.860 ;
        RECT 193.290 353.900 193.520 354.880 ;
        RECT 191.640 353.500 191.840 353.520 ;
        RECT 192.660 353.510 192.980 353.830 ;
        RECT 193.290 353.550 193.550 353.900 ;
        RECT 191.630 353.260 191.860 353.500 ;
        RECT 193.310 353.390 193.550 353.550 ;
        RECT 193.620 353.390 193.860 355.390 ;
        RECT 195.800 355.290 196.180 357.210 ;
        RECT 197.550 356.030 197.790 357.210 ;
        RECT 197.540 355.370 197.800 356.030 ;
        RECT 194.510 353.990 194.740 354.880 ;
        RECT 194.490 353.610 195.300 353.990 ;
        RECT 191.280 353.090 191.450 353.210 ;
        RECT 190.860 352.860 191.030 352.950 ;
        RECT 190.870 352.510 191.030 352.860 ;
        RECT 190.860 352.420 191.030 352.510 ;
        RECT 190.860 352.370 191.140 352.420 ;
        RECT 188.010 351.470 188.260 352.010 ;
        RECT 190.870 351.820 191.140 352.370 ;
        RECT 191.280 352.280 191.440 353.090 ;
        RECT 191.640 353.040 191.840 353.260 ;
        RECT 191.680 352.330 191.840 353.040 ;
        RECT 192.660 352.960 192.980 353.280 ;
        RECT 193.310 353.110 193.860 353.390 ;
        RECT 193.920 353.340 194.110 353.390 ;
        RECT 194.320 353.340 194.480 353.390 ;
        RECT 193.350 353.050 193.860 353.110 ;
        RECT 193.620 352.800 193.860 353.050 ;
        RECT 194.920 352.970 195.300 353.610 ;
        RECT 195.800 353.430 196.190 355.290 ;
        RECT 193.610 352.480 193.870 352.800 ;
        RECT 191.280 352.160 191.450 352.280 ;
        RECT 186.770 350.790 187.110 350.830 ;
        RECT 186.770 350.750 187.330 350.790 ;
        RECT 186.650 350.580 187.330 350.750 ;
        RECT 186.770 350.560 187.330 350.580 ;
        RECT 186.770 350.510 187.110 350.560 ;
        RECT 188.010 350.400 188.650 351.470 ;
        RECT 190.870 351.170 191.030 351.820 ;
        RECT 191.280 351.170 191.470 352.160 ;
        RECT 191.640 352.110 191.840 352.330 ;
        RECT 191.630 351.870 191.860 352.110 ;
        RECT 192.660 352.090 192.980 352.410 ;
        RECT 191.640 351.850 191.840 351.870 ;
        RECT 191.680 351.170 191.840 351.850 ;
        RECT 192.660 351.540 192.980 351.860 ;
        RECT 193.620 351.160 193.860 352.480 ;
        RECT 195.800 351.160 196.180 353.430 ;
        RECT 196.260 353.300 196.500 353.390 ;
        RECT 197.550 352.760 197.790 355.370 ;
        RECT 199.830 353.860 200.230 357.210 ;
        RECT 205.430 357.070 205.710 357.720 ;
        RECT 205.960 357.070 206.150 358.530 ;
        RECT 207.360 357.450 207.670 357.890 ;
        RECT 201.030 353.860 201.220 354.840 ;
        RECT 199.200 353.490 199.480 353.810 ;
        RECT 199.630 353.670 201.220 353.860 ;
        RECT 198.440 353.290 198.820 353.390 ;
        RECT 199.260 353.190 199.420 353.490 ;
        RECT 199.630 353.320 199.820 353.670 ;
        RECT 199.830 353.480 200.230 353.670 ;
        RECT 201.470 353.480 201.750 354.930 ;
        RECT 199.830 353.200 201.750 353.480 ;
        RECT 206.190 353.390 206.590 357.210 ;
        RECT 208.630 356.030 208.870 357.210 ;
        RECT 208.620 355.370 208.880 356.030 ;
        RECT 202.470 353.260 202.870 353.390 ;
        RECT 203.550 353.290 203.950 353.390 ;
        RECT 205.990 353.340 206.590 353.390 ;
        RECT 197.540 352.440 197.800 352.760 ;
        RECT 197.550 351.160 197.790 352.440 ;
        RECT 199.830 351.160 200.230 353.200 ;
        RECT 202.870 353.030 203.550 353.250 ;
        RECT 206.190 351.160 206.590 353.340 ;
        RECT 207.600 353.290 207.980 353.390 ;
        RECT 208.630 352.760 208.870 355.370 ;
        RECT 209.660 354.490 210.030 358.970 ;
        RECT 210.470 357.210 210.840 377.950 ;
        RECT 226.650 376.240 230.980 378.700 ;
        RECT 234.500 378.530 238.450 379.300 ;
        RECT 247.430 378.950 247.990 379.450 ;
        RECT 263.110 379.300 267.020 380.850 ;
        RECT 276.850 380.590 277.470 384.010 ;
        RECT 281.320 381.130 304.670 385.430 ;
        RECT 305.440 384.010 306.010 384.020 ;
        RECT 281.320 380.850 295.610 381.130 ;
        RECT 276.850 380.580 277.420 380.590 ;
        RECT 247.440 378.730 247.990 378.950 ;
        RECT 226.650 375.470 231.000 376.240 ;
        RECT 211.220 373.240 211.670 373.670 ;
        RECT 210.240 355.290 210.840 357.210 ;
        RECT 209.630 354.030 210.080 354.490 ;
        RECT 209.660 353.990 210.030 354.030 ;
        RECT 210.230 353.900 210.840 355.290 ;
        RECT 210.230 353.440 210.880 353.900 ;
        RECT 210.230 353.430 210.840 353.440 ;
        RECT 210.240 353.390 210.840 353.430 ;
        RECT 209.920 353.320 210.160 353.390 ;
        RECT 208.620 352.440 208.880 352.760 ;
        RECT 208.630 351.160 208.870 352.440 ;
        RECT 210.240 351.160 210.620 353.390 ;
        RECT 211.240 351.550 211.610 373.240 ;
        RECT 217.790 372.190 218.370 372.750 ;
        RECT 226.650 372.480 230.980 375.470 ;
        RECT 214.580 370.620 215.140 371.270 ;
        RECT 215.530 371.110 216.090 371.690 ;
        RECT 216.610 371.570 217.170 372.160 ;
        RECT 212.110 368.160 212.540 368.600 ;
        RECT 211.780 365.220 211.990 365.330 ;
        RECT 212.120 363.120 212.490 368.160 ;
        RECT 213.660 365.330 213.890 369.150 ;
        RECT 212.660 365.270 212.870 365.330 ;
        RECT 213.660 365.260 213.920 365.330 ;
        RECT 211.790 359.290 212.020 359.410 ;
        RECT 212.120 357.210 212.670 363.120 ;
        RECT 213.660 362.150 213.890 365.260 ;
        RECT 213.650 361.900 213.890 362.150 ;
        RECT 214.600 362.070 215.100 370.620 ;
        RECT 212.120 357.070 212.800 357.210 ;
        RECT 213.660 357.070 213.890 361.900 ;
        RECT 214.460 361.750 215.100 362.070 ;
        RECT 214.600 358.380 215.100 361.750 ;
        RECT 214.490 358.060 215.100 358.380 ;
        RECT 214.600 357.210 215.100 358.060 ;
        RECT 215.530 369.150 216.030 371.110 ;
        RECT 215.530 357.210 216.370 369.150 ;
        RECT 216.400 359.210 216.630 359.290 ;
        RECT 212.120 353.390 212.490 357.070 ;
        RECT 212.560 356.050 212.800 357.070 ;
        RECT 213.440 356.520 213.760 356.840 ;
        RECT 214.580 356.510 215.140 357.210 ;
        RECT 215.390 357.080 216.370 357.210 ;
        RECT 215.390 356.560 216.030 357.080 ;
        RECT 212.540 355.390 212.810 356.050 ;
        RECT 213.440 355.970 213.760 356.290 ;
        RECT 214.560 356.270 215.140 356.510 ;
        RECT 212.560 353.390 212.800 355.390 ;
        RECT 213.440 355.090 213.760 355.410 ;
        RECT 214.580 355.110 215.140 356.270 ;
        RECT 215.280 355.960 216.030 356.560 ;
        RECT 215.390 355.420 216.030 355.960 ;
        RECT 214.560 354.870 215.140 355.110 ;
        RECT 213.440 354.540 213.760 354.860 ;
        RECT 214.580 354.300 215.140 354.870 ;
        RECT 215.280 354.820 216.030 355.420 ;
        RECT 214.580 354.070 215.170 354.300 ;
        RECT 213.440 353.510 213.760 353.830 ;
        RECT 214.580 353.500 215.140 354.070 ;
        RECT 215.390 353.550 216.030 354.820 ;
        RECT 211.940 353.340 212.100 353.390 ;
        RECT 212.120 353.340 212.500 353.390 ;
        RECT 212.560 353.350 212.910 353.390 ;
        RECT 211.210 351.540 211.610 351.550 ;
        RECT 211.200 351.120 211.620 351.540 ;
        RECT 211.240 351.110 211.610 351.120 ;
        RECT 188.010 350.150 188.260 350.400 ;
        RECT 186.770 349.990 187.110 350.040 ;
        RECT 186.770 349.970 187.330 349.990 ;
        RECT 186.650 349.800 187.330 349.970 ;
        RECT 186.770 349.760 187.330 349.800 ;
        RECT 186.770 349.720 187.110 349.760 ;
        RECT 188.010 349.080 188.650 350.150 ;
        RECT 188.010 348.540 188.260 349.080 ;
        RECT 186.770 347.860 187.110 347.900 ;
        RECT 186.770 347.820 187.330 347.860 ;
        RECT 183.580 343.820 183.820 347.250 ;
        RECT 183.560 343.570 183.950 343.820 ;
        RECT 183.700 343.320 183.950 343.570 ;
        RECT 183.450 342.830 183.920 343.320 ;
        RECT 184.310 343.180 184.680 343.200 ;
        RECT 184.260 342.920 184.680 343.180 ;
        RECT 184.310 342.910 184.680 342.920 ;
        RECT 163.360 342.130 163.770 342.460 ;
        RECT 164.100 342.150 164.340 342.550 ;
        RECT 167.040 342.150 167.350 342.550 ;
        RECT 163.910 342.100 164.340 342.150 ;
        RECT 163.360 340.580 163.770 340.910 ;
        RECT 163.360 339.030 163.770 339.360 ;
        RECT 163.360 337.480 163.770 337.810 ;
        RECT 164.100 336.310 164.340 342.100 ;
        RECT 166.850 342.090 167.350 342.150 ;
        RECT 165.520 341.600 165.720 341.620 ;
        RECT 165.520 341.310 165.870 341.600 ;
        RECT 165.520 340.050 165.720 340.070 ;
        RECT 165.520 339.760 165.870 340.050 ;
        RECT 165.520 338.500 165.720 338.520 ;
        RECT 165.520 338.210 165.870 338.500 ;
        RECT 167.040 337.640 167.350 342.090 ;
        RECT 167.600 342.020 167.880 342.350 ;
        RECT 171.470 342.150 171.760 342.550 ;
        RECT 171.280 342.100 171.760 342.150 ;
        RECT 178.860 342.140 179.180 342.480 ;
        RECT 183.270 342.390 183.590 342.670 ;
        RECT 183.730 342.570 183.920 342.830 ;
        RECT 183.730 342.280 183.960 342.570 ;
        RECT 170.400 341.200 170.720 341.500 ;
        RECT 167.600 340.470 167.880 340.800 ;
        RECT 170.400 339.650 170.720 339.950 ;
        RECT 167.600 338.920 167.880 339.250 ;
        RECT 170.400 338.100 170.720 338.400 ;
        RECT 167.600 337.640 167.880 337.700 ;
        RECT 163.910 335.910 164.150 335.960 ;
        RECT 164.400 324.940 164.640 337.570 ;
        RECT 167.040 337.370 167.880 337.640 ;
        RECT 165.520 336.950 165.720 336.970 ;
        RECT 165.520 336.660 165.870 336.950 ;
        RECT 167.040 336.490 167.650 337.370 ;
        RECT 171.470 337.000 171.760 342.100 ;
        RECT 171.770 337.000 172.060 337.620 ;
        RECT 172.270 337.020 172.610 337.340 ;
        RECT 170.400 336.550 170.720 336.850 ;
        RECT 171.470 336.650 172.090 337.000 ;
        RECT 167.040 336.310 167.670 336.490 ;
        RECT 171.470 336.310 171.760 336.650 ;
        RECT 167.300 336.160 167.670 336.310 ;
        RECT 171.770 336.190 172.060 336.650 ;
        RECT 172.270 336.410 172.520 337.020 ;
        RECT 173.230 336.430 173.420 337.630 ;
        RECT 177.510 336.960 177.760 337.690 ;
        RECT 178.940 337.380 179.150 342.140 ;
        RECT 183.730 341.680 183.920 342.280 ;
        RECT 183.270 341.290 183.590 341.570 ;
        RECT 183.730 341.390 183.960 341.680 ;
        RECT 183.730 341.130 183.920 341.390 ;
        RECT 180.200 340.450 180.590 340.700 ;
        RECT 183.450 340.640 183.920 341.130 ;
        RECT 184.310 341.040 184.680 341.050 ;
        RECT 184.260 340.780 184.680 341.040 ;
        RECT 184.310 340.760 184.680 340.780 ;
        RECT 179.480 339.350 179.820 339.690 ;
        RECT 179.520 339.330 179.740 339.350 ;
        RECT 178.910 337.060 179.190 337.380 ;
        RECT 179.520 337.050 179.720 339.330 ;
        RECT 179.980 337.370 180.170 337.870 ;
        RECT 177.480 336.670 177.820 336.960 ;
        RECT 179.480 336.730 179.760 337.050 ;
        RECT 179.940 337.040 180.220 337.370 ;
        RECT 166.850 335.910 167.160 335.980 ;
        RECT 167.340 334.950 167.650 336.160 ;
        RECT 171.200 335.910 172.060 336.190 ;
        RECT 171.120 335.900 172.060 335.910 ;
        RECT 172.220 336.300 172.520 336.410 ;
        RECT 171.120 335.430 171.580 335.900 ;
        RECT 167.290 334.470 167.710 334.950 ;
        RECT 172.220 334.790 172.410 336.300 ;
        RECT 173.170 336.110 173.490 336.430 ;
        RECT 175.850 335.900 176.600 336.090 ;
        RECT 176.100 335.060 176.600 335.900 ;
        RECT 180.410 335.820 180.590 340.450 ;
        RECT 183.730 340.390 183.920 340.640 ;
        RECT 183.450 339.900 183.920 340.390 ;
        RECT 184.310 340.250 184.680 340.270 ;
        RECT 184.260 339.990 184.680 340.250 ;
        RECT 184.310 339.980 184.680 339.990 ;
        RECT 183.270 339.460 183.590 339.740 ;
        RECT 183.730 339.640 183.920 339.900 ;
        RECT 183.730 339.350 183.960 339.640 ;
        RECT 183.730 338.750 183.920 339.350 ;
        RECT 183.270 338.360 183.590 338.640 ;
        RECT 183.730 338.460 183.960 338.750 ;
        RECT 183.730 338.200 183.920 338.460 ;
        RECT 183.450 337.770 183.920 338.200 ;
        RECT 184.310 338.110 184.680 338.120 ;
        RECT 184.260 337.850 184.680 338.110 ;
        RECT 184.310 337.830 184.680 337.850 ;
        RECT 183.450 337.710 183.950 337.770 ;
        RECT 181.730 336.980 181.990 337.010 ;
        RECT 181.710 336.680 182.010 336.980 ;
        RECT 181.730 336.670 181.990 336.680 ;
        RECT 180.410 335.520 180.890 335.820 ;
        RECT 181.740 335.750 181.960 336.670 ;
        RECT 183.700 336.540 183.950 337.710 ;
        RECT 185.040 337.490 185.270 343.540 ;
        RECT 185.760 343.190 186.140 347.680 ;
        RECT 186.650 347.650 187.330 347.820 ;
        RECT 186.770 347.630 187.330 347.650 ;
        RECT 186.770 347.580 187.110 347.630 ;
        RECT 187.510 343.800 187.750 347.540 ;
        RECT 188.010 347.470 188.650 348.540 ;
        RECT 188.010 347.250 188.260 347.470 ;
        RECT 187.510 343.530 187.980 343.800 ;
        RECT 187.710 343.300 187.980 343.530 ;
        RECT 188.010 343.320 188.260 343.540 ;
        RECT 186.770 343.160 187.110 343.210 ;
        RECT 186.770 343.140 187.330 343.160 ;
        RECT 186.650 342.970 187.330 343.140 ;
        RECT 186.770 342.930 187.330 342.970 ;
        RECT 186.770 342.890 187.110 342.930 ;
        RECT 188.010 342.250 188.650 343.320 ;
        RECT 189.790 343.170 190.190 347.700 ;
        RECT 191.450 347.170 191.610 347.820 ;
        RECT 191.450 346.620 191.720 347.170 ;
        RECT 191.440 346.570 191.720 346.620 ;
        RECT 191.860 346.830 192.050 347.820 ;
        RECT 192.260 347.140 192.420 347.820 ;
        RECT 193.310 347.450 193.550 347.540 ;
        RECT 192.220 347.120 192.420 347.140 ;
        RECT 193.240 347.400 193.560 347.450 ;
        RECT 193.240 347.340 193.670 347.400 ;
        RECT 193.920 347.350 194.110 347.410 ;
        RECT 193.240 347.130 193.560 347.340 ;
        RECT 192.210 346.880 192.440 347.120 ;
        RECT 193.310 346.900 193.550 347.130 ;
        RECT 191.860 346.710 192.030 346.830 ;
        RECT 191.440 346.480 191.610 346.570 ;
        RECT 191.450 346.120 191.610 346.480 ;
        RECT 191.440 346.030 191.610 346.120 ;
        RECT 191.440 345.980 191.720 346.030 ;
        RECT 191.450 345.430 191.720 345.980 ;
        RECT 191.860 345.890 192.020 346.710 ;
        RECT 192.220 346.660 192.420 346.880 ;
        RECT 192.260 345.940 192.420 346.660 ;
        RECT 193.240 346.580 193.560 346.900 ;
        RECT 193.310 346.020 193.550 346.580 ;
        RECT 191.860 345.770 192.030 345.890 ;
        RECT 191.450 344.160 191.610 345.430 ;
        RECT 191.860 344.910 192.050 345.770 ;
        RECT 192.220 345.720 192.420 345.940 ;
        RECT 192.210 345.480 192.440 345.720 ;
        RECT 193.240 345.700 193.560 346.020 ;
        RECT 192.220 345.460 192.420 345.480 ;
        RECT 193.310 345.470 193.550 345.700 ;
        RECT 191.830 344.680 192.070 344.910 ;
        RECT 191.450 343.610 191.720 344.160 ;
        RECT 191.440 343.560 191.720 343.610 ;
        RECT 191.860 343.820 192.050 344.680 ;
        RECT 192.260 344.130 192.420 345.460 ;
        RECT 193.240 345.150 193.560 345.470 ;
        RECT 193.310 345.030 193.550 345.150 ;
        RECT 193.310 344.790 193.890 345.030 ;
        RECT 192.220 344.110 192.420 344.130 ;
        RECT 193.240 344.120 193.560 344.440 ;
        RECT 192.210 343.870 192.440 344.110 ;
        RECT 191.860 343.700 192.030 343.820 ;
        RECT 191.440 343.470 191.610 343.560 ;
        RECT 191.450 343.120 191.610 343.470 ;
        RECT 191.440 343.030 191.610 343.120 ;
        RECT 191.440 342.980 191.720 343.030 ;
        RECT 191.450 342.430 191.720 342.980 ;
        RECT 191.860 342.890 192.020 343.700 ;
        RECT 192.220 343.650 192.420 343.870 ;
        RECT 192.260 342.940 192.420 343.650 ;
        RECT 193.240 343.570 193.560 343.890 ;
        RECT 193.650 343.450 193.890 344.790 ;
        RECT 194.320 344.000 194.570 347.820 ;
        RECT 196.380 347.420 196.760 347.820 ;
        RECT 196.260 347.340 196.760 347.420 ;
        RECT 196.380 345.900 196.760 347.340 ;
        RECT 198.330 347.430 198.600 347.820 ;
        RECT 198.330 347.340 198.820 347.430 ;
        RECT 200.410 347.410 200.810 347.820 ;
        RECT 200.190 347.340 200.810 347.410 ;
        RECT 202.470 347.340 202.870 347.460 ;
        RECT 203.550 347.340 203.950 347.460 ;
        RECT 205.990 347.340 206.230 347.410 ;
        RECT 207.600 347.340 207.980 347.490 ;
        RECT 212.120 347.410 212.490 353.340 ;
        RECT 212.560 353.050 213.070 353.350 ;
        RECT 212.560 352.800 212.800 353.050 ;
        RECT 213.440 352.960 213.760 353.280 ;
        RECT 214.560 353.260 215.140 353.500 ;
        RECT 212.550 352.480 212.810 352.800 ;
        RECT 212.560 351.160 212.800 352.480 ;
        RECT 213.440 352.090 213.760 352.410 ;
        RECT 214.580 352.110 215.140 353.260 ;
        RECT 215.280 352.950 216.030 353.550 ;
        RECT 215.390 352.420 216.030 352.950 ;
        RECT 214.560 351.870 215.140 352.110 ;
        RECT 213.440 351.540 213.760 351.860 ;
        RECT 214.580 351.170 215.140 351.870 ;
        RECT 215.280 351.820 216.030 352.420 ;
        RECT 215.390 351.170 216.030 351.820 ;
        RECT 209.920 347.340 210.160 347.400 ;
        RECT 211.940 347.350 212.100 347.410 ;
        RECT 212.120 347.350 212.500 347.410 ;
        RECT 212.750 347.350 212.910 347.410 ;
        RECT 196.380 344.040 196.770 345.900 ;
        RECT 194.110 343.930 194.270 344.000 ;
        RECT 194.320 343.930 194.710 344.000 ;
        RECT 194.920 343.930 195.080 344.000 ;
        RECT 194.320 343.380 194.570 343.930 ;
        RECT 196.380 343.740 196.760 344.040 ;
        RECT 196.380 343.420 196.800 343.740 ;
        RECT 194.300 343.350 194.580 343.380 ;
        RECT 194.290 343.070 194.590 343.350 ;
        RECT 194.300 343.050 194.580 343.070 ;
        RECT 191.860 342.770 192.030 342.890 ;
        RECT 188.010 341.710 188.260 342.250 ;
        RECT 191.450 341.780 191.610 342.430 ;
        RECT 191.860 341.780 192.050 342.770 ;
        RECT 192.220 342.720 192.420 342.940 ;
        RECT 192.210 342.480 192.440 342.720 ;
        RECT 193.240 342.700 193.560 343.020 ;
        RECT 192.220 342.460 192.420 342.480 ;
        RECT 192.260 341.780 192.420 342.460 ;
        RECT 193.240 342.150 193.560 342.470 ;
        RECT 193.250 342.070 193.510 342.150 ;
        RECT 193.240 341.870 193.510 342.070 ;
        RECT 186.770 341.030 187.110 341.070 ;
        RECT 186.770 340.990 187.330 341.030 ;
        RECT 186.650 340.820 187.330 340.990 ;
        RECT 186.770 340.800 187.330 340.820 ;
        RECT 186.770 340.750 187.110 340.800 ;
        RECT 188.010 340.640 188.650 341.710 ;
        RECT 193.240 341.180 193.450 341.870 ;
        RECT 194.320 341.770 194.570 343.050 ;
        RECT 196.380 342.690 196.760 343.420 ;
        RECT 198.330 343.350 198.600 347.340 ;
        RECT 199.040 343.900 199.420 344.000 ;
        RECT 198.310 343.040 198.620 343.350 ;
        RECT 196.380 342.370 196.780 342.690 ;
        RECT 196.380 341.770 196.760 342.370 ;
        RECT 198.330 341.770 198.600 343.040 ;
        RECT 198.770 342.390 199.030 342.450 ;
        RECT 198.760 342.130 199.030 342.390 ;
        RECT 198.250 341.200 198.510 341.520 ;
        RECT 193.230 340.860 193.490 341.180 ;
        RECT 188.010 340.390 188.260 340.640 ;
        RECT 196.520 340.490 196.780 340.810 ;
        RECT 186.770 340.230 187.110 340.280 ;
        RECT 186.770 340.210 187.330 340.230 ;
        RECT 186.650 340.040 187.330 340.210 ;
        RECT 186.770 340.000 187.330 340.040 ;
        RECT 186.770 339.960 187.110 340.000 ;
        RECT 188.010 339.320 188.650 340.390 ;
        RECT 196.520 339.630 196.680 340.490 ;
        RECT 188.010 338.780 188.260 339.320 ;
        RECT 196.360 339.310 196.680 339.630 ;
        RECT 197.780 339.360 198.040 339.680 ;
        RECT 193.150 338.820 193.470 339.140 ;
        RECT 186.770 338.100 187.110 338.140 ;
        RECT 186.770 338.060 187.330 338.100 ;
        RECT 186.650 337.890 187.330 338.060 ;
        RECT 186.770 337.870 187.330 337.890 ;
        RECT 186.770 337.820 187.110 337.870 ;
        RECT 187.710 336.560 187.980 337.790 ;
        RECT 188.010 337.710 188.650 338.780 ;
        RECT 197.280 338.430 197.540 338.750 ;
        RECT 193.200 337.970 193.520 338.290 ;
        RECT 188.010 337.490 188.260 337.710 ;
        RECT 190.530 336.990 190.960 337.390 ;
        RECT 183.690 336.280 184.010 336.540 ;
        RECT 187.710 336.250 188.060 336.560 ;
        RECT 180.490 335.410 180.890 335.520 ;
        RECT 181.680 335.350 182.020 335.750 ;
        RECT 181.740 335.270 181.960 335.350 ;
        RECT 185.690 335.080 186.630 336.010 ;
        RECT 190.570 335.200 190.920 336.990 ;
        RECT 192.390 336.430 192.610 337.750 ;
        RECT 193.650 337.030 193.880 337.750 ;
        RECT 193.650 336.800 196.860 337.030 ;
        RECT 193.650 336.790 193.880 336.800 ;
        RECT 192.100 336.190 192.610 336.430 ;
        RECT 171.780 334.470 172.410 334.790 ;
        RECT 175.610 334.740 175.850 335.060 ;
        RECT 176.850 334.740 177.090 335.060 ;
        RECT 185.420 334.760 185.660 335.080 ;
        RECT 186.660 334.760 186.900 335.080 ;
        RECT 192.100 334.940 192.330 336.190 ;
        RECT 196.630 335.830 196.860 336.800 ;
        RECT 196.580 335.430 196.890 335.830 ;
        RECT 191.990 334.500 192.450 334.940 ;
        RECT 171.780 334.370 172.220 334.470 ;
        RECT 175.610 333.400 175.850 333.720 ;
        RECT 176.850 333.390 177.090 333.710 ;
        RECT 185.420 333.420 185.660 333.740 ;
        RECT 186.660 333.410 186.900 333.730 ;
        RECT 196.630 332.260 196.860 335.430 ;
        RECT 196.500 332.040 196.860 332.260 ;
        RECT 175.960 331.770 176.220 331.970 ;
        RECT 176.480 331.770 176.740 331.970 ;
        RECT 172.690 331.250 173.010 331.570 ;
        RECT 173.780 331.250 174.100 331.570 ;
        RECT 174.880 331.240 175.200 331.560 ;
        RECT 175.960 330.960 176.270 331.770 ;
        RECT 176.430 330.960 176.740 331.770 ;
        RECT 185.770 331.800 186.030 332.000 ;
        RECT 186.290 331.800 186.550 332.000 ;
        RECT 196.300 331.810 196.860 332.040 ;
        RECT 196.300 331.800 196.840 331.810 ;
        RECT 177.500 331.240 177.820 331.560 ;
        RECT 178.600 331.250 178.920 331.570 ;
        RECT 179.690 331.250 180.010 331.570 ;
        RECT 182.500 331.280 182.820 331.600 ;
        RECT 183.590 331.280 183.910 331.600 ;
        RECT 184.690 331.270 185.010 331.590 ;
        RECT 185.770 330.990 186.080 331.800 ;
        RECT 186.240 330.990 186.550 331.800 ;
        RECT 187.310 331.270 187.630 331.590 ;
        RECT 188.410 331.280 188.730 331.600 ;
        RECT 189.500 331.280 189.820 331.600 ;
        RECT 193.800 331.250 194.120 331.570 ;
        RECT 194.900 331.260 195.220 331.580 ;
        RECT 195.990 331.260 196.310 331.580 ;
        RECT 171.990 329.190 172.310 330.940 ;
        RECT 173.240 330.570 173.560 330.890 ;
        RECT 174.330 330.550 174.650 330.870 ;
        RECT 175.610 330.860 175.850 330.950 ;
        RECT 175.440 330.630 175.850 330.860 ;
        RECT 175.440 330.540 175.760 330.630 ;
        RECT 175.960 330.430 176.220 330.960 ;
        RECT 175.850 329.970 176.220 330.430 ;
        RECT 175.840 329.630 176.220 329.970 ;
        RECT 173.240 329.200 173.560 329.520 ;
        RECT 174.330 329.200 174.650 329.520 ;
        RECT 175.430 329.200 175.750 329.520 ;
        RECT 171.870 328.590 172.410 329.190 ;
        RECT 172.680 328.470 173.000 328.790 ;
        RECT 173.780 328.470 174.100 328.790 ;
        RECT 174.880 328.470 175.200 328.790 ;
        RECT 175.850 328.220 176.220 329.630 ;
        RECT 176.480 330.430 176.740 330.960 ;
        RECT 176.850 330.860 177.090 330.940 ;
        RECT 176.850 330.620 177.260 330.860 ;
        RECT 176.940 330.540 177.260 330.620 ;
        RECT 178.050 330.550 178.370 330.870 ;
        RECT 179.140 330.570 179.460 330.890 ;
        RECT 176.480 329.990 176.850 330.430 ;
        RECT 176.480 329.650 176.860 329.990 ;
        RECT 176.480 328.220 176.850 329.650 ;
        RECT 176.950 329.200 177.270 329.520 ;
        RECT 178.050 329.200 178.370 329.520 ;
        RECT 179.140 329.200 179.460 329.520 ;
        RECT 177.500 328.470 177.820 328.790 ;
        RECT 178.600 328.470 178.920 328.790 ;
        RECT 179.700 328.470 180.020 328.790 ;
        RECT 172.680 327.100 173.000 327.420 ;
        RECT 173.780 327.100 174.100 327.420 ;
        RECT 174.880 327.100 175.200 327.420 ;
        RECT 172.110 326.460 172.430 326.780 ;
        RECT 173.240 326.420 173.560 326.740 ;
        RECT 174.330 326.420 174.650 326.740 ;
        RECT 175.430 326.430 175.750 326.750 ;
        RECT 172.120 325.990 172.440 326.310 ;
        RECT 164.000 323.620 164.650 324.940 ;
        RECT 175.850 324.790 176.850 328.220 ;
        RECT 180.360 328.170 180.700 330.960 ;
        RECT 180.300 327.650 180.760 328.170 ;
        RECT 177.500 327.100 177.820 327.420 ;
        RECT 178.600 327.100 178.920 327.420 ;
        RECT 179.700 327.100 180.020 327.420 ;
        RECT 181.790 327.280 182.130 330.950 ;
        RECT 183.050 330.600 183.370 330.920 ;
        RECT 184.140 330.580 184.460 330.900 ;
        RECT 185.420 330.890 185.660 330.970 ;
        RECT 185.250 330.650 185.660 330.890 ;
        RECT 185.250 330.570 185.570 330.650 ;
        RECT 185.770 330.460 186.030 330.990 ;
        RECT 185.660 329.970 186.030 330.460 ;
        RECT 185.650 329.630 186.030 329.970 ;
        RECT 183.050 329.230 183.370 329.550 ;
        RECT 184.140 329.230 184.460 329.550 ;
        RECT 185.240 329.230 185.560 329.550 ;
        RECT 182.490 328.500 182.810 328.820 ;
        RECT 183.590 328.500 183.910 328.820 ;
        RECT 184.690 328.500 185.010 328.820 ;
        RECT 185.660 328.450 186.030 329.630 ;
        RECT 186.290 330.460 186.550 330.990 ;
        RECT 186.660 330.890 186.900 330.970 ;
        RECT 186.660 330.650 187.070 330.890 ;
        RECT 186.750 330.570 187.070 330.650 ;
        RECT 187.860 330.580 188.180 330.900 ;
        RECT 188.950 330.600 189.270 330.920 ;
        RECT 186.290 328.450 186.660 330.460 ;
        RECT 186.760 329.230 187.080 329.550 ;
        RECT 187.860 329.230 188.180 329.550 ;
        RECT 188.950 329.230 189.270 329.550 ;
        RECT 187.310 328.500 187.630 328.820 ;
        RECT 188.410 328.500 188.730 328.820 ;
        RECT 189.510 328.500 189.830 328.820 ;
        RECT 181.700 326.810 182.220 327.280 ;
        RECT 182.490 327.130 182.810 327.450 ;
        RECT 183.590 327.130 183.910 327.450 ;
        RECT 184.690 327.130 185.010 327.450 ;
        RECT 176.950 326.430 177.270 326.750 ;
        RECT 178.050 326.420 178.370 326.740 ;
        RECT 179.140 326.420 179.460 326.740 ;
        RECT 180.270 326.460 180.590 326.780 ;
        RECT 181.700 326.760 182.240 326.810 ;
        RECT 181.920 326.490 182.240 326.760 ;
        RECT 183.050 326.450 183.370 326.770 ;
        RECT 184.140 326.450 184.460 326.770 ;
        RECT 185.240 326.460 185.560 326.780 ;
        RECT 180.260 325.990 180.580 326.310 ;
        RECT 181.930 326.020 182.250 326.340 ;
        RECT 185.660 324.810 186.660 328.450 ;
        RECT 187.310 327.130 187.630 327.450 ;
        RECT 188.410 327.130 188.730 327.450 ;
        RECT 189.510 327.130 189.830 327.450 ;
        RECT 190.210 326.810 190.480 330.990 ;
        RECT 193.240 330.550 193.560 330.870 ;
        RECT 194.350 330.560 194.670 330.880 ;
        RECT 195.440 330.580 195.760 330.900 ;
        RECT 197.280 330.590 197.530 338.430 ;
        RECT 197.780 331.490 198.030 339.360 ;
        RECT 198.260 332.400 198.510 341.200 ;
        RECT 198.760 333.290 199.010 342.130 ;
        RECT 200.410 341.770 200.810 347.340 ;
        RECT 212.120 346.370 212.490 347.350 ;
        RECT 212.080 345.860 212.570 346.370 ;
        RECT 212.120 345.830 212.490 345.860 ;
        RECT 203.070 343.860 203.470 344.000 ;
        RECT 204.590 343.220 204.910 343.540 ;
        RECT 204.740 342.540 205.060 342.860 ;
        RECT 204.740 341.650 205.060 341.970 ;
        RECT 204.590 340.970 204.910 341.290 ;
        RECT 204.590 340.450 204.910 340.770 ;
        RECT 204.740 339.770 205.060 340.090 ;
        RECT 204.740 338.880 205.060 339.200 ;
        RECT 204.590 338.200 204.910 338.520 ;
        RECT 199.040 337.950 199.420 338.050 ;
        RECT 205.670 337.950 205.900 344.000 ;
        RECT 206.930 339.650 207.160 344.000 ;
        RECT 206.890 339.640 207.170 339.650 ;
        RECT 206.890 339.320 207.190 339.640 ;
        RECT 206.930 337.950 207.160 339.320 ;
        RECT 214.600 334.790 215.100 351.170 ;
        RECT 215.530 340.070 216.030 351.170 ;
        RECT 216.660 345.300 217.160 371.570 ;
        RECT 217.790 359.630 218.290 372.190 ;
        RECT 226.650 370.590 227.930 372.480 ;
        RECT 226.640 369.250 227.930 370.590 ;
        RECT 219.900 365.180 220.320 365.330 ;
        RECT 220.930 365.180 221.350 365.330 ;
        RECT 224.630 365.250 224.860 365.330 ;
        RECT 219.900 365.040 221.350 365.180 ;
        RECT 223.110 362.610 223.580 363.100 ;
        RECT 217.560 359.330 218.290 359.630 ;
        RECT 217.790 359.290 218.290 359.330 ;
        RECT 223.160 359.630 223.560 362.610 ;
        RECT 224.080 362.000 224.500 362.360 ;
        RECT 223.160 359.330 223.680 359.630 ;
        RECT 223.160 359.300 223.560 359.330 ;
        RECT 217.620 359.210 218.290 359.290 ;
        RECT 217.790 356.650 218.290 359.210 ;
        RECT 219.910 359.140 221.350 359.300 ;
        RECT 223.160 359.210 223.640 359.300 ;
        RECT 217.650 356.480 218.290 356.650 ;
        RECT 217.790 356.190 218.290 356.480 ;
        RECT 217.630 355.890 218.290 356.190 ;
        RECT 217.660 355.790 218.290 355.890 ;
        RECT 217.790 350.470 218.290 355.790 ;
        RECT 217.740 349.910 218.290 350.470 ;
        RECT 216.650 344.740 217.170 345.300 ;
        RECT 215.520 339.550 216.040 340.070 ;
        RECT 214.440 334.220 215.100 334.790 ;
        RECT 198.710 332.710 199.080 333.290 ;
        RECT 198.180 331.820 198.550 332.400 ;
        RECT 197.690 330.910 198.060 331.490 ;
        RECT 193.250 329.210 193.570 329.530 ;
        RECT 194.350 329.210 194.670 329.530 ;
        RECT 195.440 329.210 195.760 329.530 ;
        RECT 195.950 328.800 196.280 330.370 ;
        RECT 197.220 330.020 197.570 330.590 ;
        RECT 193.800 328.480 194.120 328.800 ;
        RECT 194.900 328.480 195.220 328.800 ;
        RECT 195.950 328.480 196.320 328.800 ;
        RECT 195.950 327.430 196.280 328.480 ;
        RECT 196.720 327.920 197.000 328.450 ;
        RECT 196.720 327.620 197.180 327.920 ;
        RECT 196.710 327.600 197.180 327.620 ;
        RECT 193.800 327.110 194.120 327.430 ;
        RECT 194.900 327.110 195.220 327.430 ;
        RECT 195.950 327.110 196.320 327.430 ;
        RECT 196.710 327.170 197.000 327.600 ;
        RECT 186.760 326.460 187.080 326.780 ;
        RECT 187.860 326.450 188.180 326.770 ;
        RECT 188.950 326.450 189.270 326.770 ;
        RECT 190.080 326.490 190.480 326.810 ;
        RECT 190.210 326.400 190.480 326.490 ;
        RECT 193.250 326.440 193.570 326.760 ;
        RECT 194.350 326.430 194.670 326.750 ;
        RECT 195.440 326.430 195.760 326.750 ;
        RECT 190.100 326.340 190.590 326.400 ;
        RECT 190.070 326.020 190.590 326.340 ;
        RECT 190.100 325.840 190.590 326.020 ;
        RECT 186.790 324.810 187.680 324.850 ;
        RECT 175.370 324.750 177.300 324.790 ;
        RECT 174.830 323.560 177.300 324.750 ;
        RECT 162.350 319.330 162.720 319.710 ;
        RECT 161.700 318.710 162.090 319.100 ;
        RECT 161.100 318.080 161.480 318.470 ;
        RECT 160.510 317.450 160.860 317.820 ;
        RECT 159.870 316.770 160.230 317.150 ;
        RECT 159.280 316.530 159.620 316.540 ;
        RECT 159.260 316.160 159.640 316.530 ;
        RECT 159.280 316.150 159.610 316.160 ;
        RECT 157.500 314.310 157.850 314.640 ;
        RECT 157.520 314.250 157.850 314.310 ;
        RECT 156.230 313.030 156.580 313.360 ;
        RECT 156.230 312.960 156.560 313.030 ;
        RECT 154.090 312.300 155.330 312.630 ;
        RECT 155.620 312.330 156.060 312.750 ;
        RECT 154.090 312.190 154.670 312.300 ;
        RECT 10.100 312.070 10.870 312.090 ;
        RECT 174.830 312.070 175.770 323.560 ;
        RECT 185.180 323.530 187.680 324.810 ;
        RECT 186.790 313.530 187.680 323.530 ;
        RECT 195.950 320.380 196.280 327.110 ;
        RECT 196.570 326.470 196.890 326.790 ;
        RECT 196.560 326.000 196.880 326.320 ;
        RECT 214.600 325.910 215.100 334.220 ;
        RECT 215.530 326.820 216.030 339.550 ;
        RECT 216.660 327.690 217.160 344.740 ;
        RECT 217.790 329.200 218.290 349.910 ;
        RECT 223.160 356.650 223.560 359.210 ;
        RECT 223.160 356.480 223.610 356.650 ;
        RECT 223.160 356.140 223.560 356.480 ;
        RECT 223.160 355.820 223.650 356.140 ;
        RECT 223.160 355.800 223.610 355.820 ;
        RECT 223.160 353.610 223.560 355.800 ;
        RECT 223.160 353.310 223.650 353.610 ;
        RECT 220.680 336.760 221.260 337.320 ;
        RECT 220.710 336.750 221.220 336.760 ;
        RECT 217.790 328.640 218.350 329.200 ;
        RECT 217.790 328.510 218.290 328.640 ;
        RECT 220.710 324.880 221.210 336.750 ;
        RECT 220.080 323.600 221.210 324.880 ;
        RECT 221.960 324.120 222.190 326.190 ;
        RECT 221.950 323.890 222.240 324.120 ;
        RECT 221.960 322.510 222.190 323.890 ;
        RECT 221.950 322.280 222.240 322.510 ;
        RECT 221.960 320.910 222.190 322.280 ;
        RECT 221.950 320.680 222.240 320.910 ;
        RECT 195.890 319.990 196.320 320.380 ;
        RECT 221.960 319.290 222.190 320.680 ;
        RECT 223.160 319.820 223.560 353.310 ;
        RECT 223.160 319.800 223.690 319.820 ;
        RECT 224.090 319.800 224.480 362.000 ;
        RECT 224.890 360.040 225.310 369.150 ;
        RECT 226.650 368.760 227.930 369.250 ;
        RECT 227.370 366.290 227.600 368.760 ;
        RECT 227.100 365.810 227.600 366.290 ;
        RECT 224.890 359.610 225.450 360.040 ;
        RECT 224.630 359.220 224.860 359.300 ;
        RECT 224.890 357.070 225.410 359.610 ;
        RECT 225.860 359.350 226.240 359.360 ;
        RECT 225.840 359.050 226.260 359.350 ;
        RECT 225.020 319.800 225.410 357.070 ;
        RECT 223.160 319.600 225.680 319.800 ;
        RECT 221.950 319.060 222.240 319.290 ;
        RECT 223.160 319.260 223.560 319.600 ;
        RECT 221.960 317.690 222.190 319.060 ;
        RECT 223.150 318.800 223.620 319.260 ;
        RECT 224.090 318.460 224.480 319.600 ;
        RECT 222.680 318.080 223.000 318.160 ;
        RECT 224.060 318.080 224.520 318.460 ;
        RECT 222.680 317.900 224.770 318.080 ;
        RECT 224.260 317.860 224.770 317.900 ;
        RECT 224.480 317.850 224.770 317.860 ;
        RECT 221.950 317.460 222.240 317.690 ;
        RECT 225.020 317.640 225.410 319.600 ;
        RECT 221.960 316.070 222.190 317.460 ;
        RECT 225.000 317.180 225.470 317.640 ;
        RECT 225.510 316.570 225.680 319.600 ;
        RECT 225.860 316.840 226.240 359.050 ;
        RECT 227.200 357.070 227.600 365.810 ;
        RECT 228.590 367.940 228.820 369.150 ;
        RECT 233.590 368.330 233.900 368.770 ;
        RECT 228.590 367.150 228.850 367.940 ;
        RECT 231.010 367.580 231.210 367.610 ;
        RECT 228.590 365.000 228.820 367.150 ;
        RECT 230.920 367.080 231.230 367.580 ;
        RECT 233.740 367.370 234.060 367.690 ;
        RECT 231.010 365.330 231.210 367.080 ;
        RECT 234.520 366.710 234.710 378.530 ;
        RECT 236.680 376.090 236.870 376.100 ;
        RECT 243.810 376.090 244.530 377.460 ;
        RECT 256.340 376.240 259.570 378.700 ;
        RECT 263.090 378.530 267.040 379.300 ;
        RECT 276.020 378.950 276.580 379.450 ;
        RECT 291.700 379.300 295.610 380.850 ;
        RECT 305.440 380.590 306.060 384.010 ;
        RECT 309.910 381.130 333.260 385.430 ;
        RECT 334.030 384.010 334.600 384.020 ;
        RECT 309.910 380.850 324.200 381.130 ;
        RECT 305.440 380.580 306.010 380.590 ;
        RECT 276.030 378.730 276.580 378.950 ;
        RECT 284.930 376.240 288.160 378.700 ;
        RECT 291.680 378.530 295.630 379.300 ;
        RECT 304.610 378.950 305.170 379.450 ;
        RECT 320.290 379.300 324.200 380.850 ;
        RECT 334.030 380.590 334.650 384.010 ;
        RECT 338.500 381.130 361.850 385.430 ;
        RECT 362.620 384.010 363.190 384.020 ;
        RECT 338.500 380.850 352.790 381.130 ;
        RECT 334.030 380.580 334.600 380.590 ;
        RECT 304.620 378.730 305.170 378.950 ;
        RECT 313.520 376.240 316.750 378.700 ;
        RECT 320.270 378.530 324.220 379.300 ;
        RECT 333.200 378.950 333.760 379.450 ;
        RECT 348.880 379.300 352.790 380.850 ;
        RECT 362.620 380.590 363.240 384.010 ;
        RECT 362.620 380.580 363.190 380.590 ;
        RECT 333.210 378.730 333.760 378.950 ;
        RECT 342.110 376.240 345.340 378.700 ;
        RECT 348.860 378.530 352.810 379.300 ;
        RECT 361.790 378.950 362.350 379.450 ;
        RECT 361.800 378.730 362.350 378.950 ;
        RECT 364.600 378.930 368.020 378.980 ;
        RECT 364.590 378.360 368.030 378.930 ;
        RECT 362.740 377.540 363.460 378.090 ;
        RECT 362.960 377.530 363.460 377.540 ;
        RECT 236.680 375.740 244.530 376.090 ;
        RECT 236.680 373.610 236.870 375.740 ;
        RECT 255.640 375.550 259.590 376.240 ;
        RECT 255.580 375.470 259.590 375.550 ;
        RECT 284.240 375.470 288.190 376.240 ;
        RECT 312.820 375.470 316.770 376.240 ;
        RECT 341.410 375.470 345.360 376.240 ;
        RECT 237.860 375.260 238.680 375.350 ;
        RECT 255.580 375.270 259.570 375.470 ;
        RECT 237.800 374.570 238.680 375.260 ;
        RECT 255.560 375.070 259.570 375.270 ;
        RECT 235.110 367.690 235.300 369.150 ;
        RECT 235.550 368.500 235.830 369.150 ;
        RECT 235.440 367.900 235.830 368.500 ;
        RECT 235.110 367.660 235.330 367.690 ;
        RECT 235.090 367.390 235.340 367.660 ;
        RECT 235.100 367.380 235.340 367.390 ;
        RECT 235.100 367.140 235.330 367.380 ;
        RECT 234.520 366.580 234.950 366.710 ;
        RECT 234.520 366.260 234.970 366.580 ;
        RECT 234.520 365.980 234.710 366.260 ;
        RECT 234.520 365.660 234.970 365.980 ;
        RECT 234.520 365.540 234.950 365.660 ;
        RECT 231.010 365.250 231.340 365.330 ;
        RECT 228.590 364.210 228.850 365.000 ;
        RECT 231.010 364.540 231.210 365.250 ;
        RECT 231.370 364.570 231.570 365.440 ;
        RECT 231.590 365.310 231.870 365.330 ;
        RECT 231.590 365.250 231.930 365.310 ;
        RECT 231.610 365.010 231.930 365.250 ;
        RECT 232.270 365.010 232.590 365.330 ;
        RECT 233.340 365.180 233.660 365.310 ;
        RECT 233.270 364.990 233.660 365.180 ;
        RECT 233.840 365.010 234.160 365.330 ;
        RECT 234.520 365.190 234.710 365.540 ;
        RECT 234.400 365.030 234.710 365.190 ;
        RECT 233.270 364.890 233.500 364.990 ;
        RECT 230.860 364.250 231.210 364.540 ;
        RECT 231.360 364.280 231.590 364.570 ;
        RECT 233.290 364.420 233.480 364.890 ;
        RECT 233.740 364.610 234.060 364.930 ;
        RECT 234.320 364.710 234.710 365.030 ;
        RECT 228.590 361.910 228.820 364.210 ;
        RECT 230.870 364.030 231.210 364.250 ;
        RECT 231.010 363.830 231.210 364.030 ;
        RECT 230.870 363.600 231.210 363.820 ;
        RECT 230.860 363.500 231.210 363.600 ;
        RECT 231.370 363.570 231.570 364.280 ;
        RECT 233.220 364.100 233.480 364.420 ;
        RECT 233.490 364.160 233.810 364.480 ;
        RECT 234.400 364.410 234.710 364.710 ;
        RECT 234.880 364.570 235.070 365.440 ;
        RECT 235.140 365.330 235.300 367.140 ;
        RECT 235.550 366.300 235.830 367.900 ;
        RECT 235.550 365.980 235.910 366.300 ;
        RECT 235.550 365.330 235.830 365.980 ;
        RECT 235.140 365.110 235.830 365.330 ;
        RECT 235.940 365.180 236.220 365.330 ;
        RECT 235.100 364.860 235.830 365.110 ;
        RECT 235.090 364.590 235.830 364.860 ;
        RECT 234.230 364.090 234.710 364.410 ;
        RECT 234.860 364.280 235.090 364.570 ;
        RECT 234.270 364.060 234.710 364.090 ;
        RECT 232.380 363.630 232.700 363.950 ;
        RECT 230.860 363.310 231.090 363.500 ;
        RECT 231.360 363.280 231.590 363.570 ;
        RECT 233.220 363.430 233.480 363.750 ;
        RECT 233.590 363.480 233.900 363.920 ;
        RECT 234.520 363.840 234.710 364.060 ;
        RECT 234.230 363.690 234.490 363.760 ;
        RECT 233.600 363.470 233.810 363.480 ;
        RECT 228.590 361.120 228.850 361.910 ;
        RECT 231.370 361.550 231.570 363.280 ;
        RECT 233.290 362.960 233.480 363.430 ;
        RECT 233.580 363.150 233.840 363.470 ;
        RECT 234.230 363.440 234.590 363.690 ;
        RECT 234.880 363.570 235.070 364.280 ;
        RECT 234.270 363.230 234.590 363.440 ;
        RECT 234.860 363.280 235.090 363.570 ;
        RECT 232.270 362.520 232.590 362.840 ;
        RECT 233.270 362.670 233.500 362.960 ;
        RECT 233.600 362.740 233.810 363.150 ;
        RECT 234.400 362.950 234.590 363.230 ;
        RECT 234.400 362.900 234.630 362.950 ;
        RECT 233.840 362.740 234.160 362.840 ;
        RECT 233.110 362.350 233.430 362.670 ;
        RECT 233.590 362.520 234.160 362.740 ;
        RECT 234.320 362.580 234.640 362.900 ;
        RECT 233.590 362.310 233.900 362.520 ;
        RECT 232.270 361.990 232.590 362.310 ;
        RECT 233.590 362.300 234.160 362.310 ;
        RECT 233.270 361.870 233.500 362.160 ;
        RECT 230.860 361.330 231.090 361.520 ;
        RECT 230.860 361.230 231.210 361.330 ;
        RECT 231.360 361.260 231.590 361.550 ;
        RECT 233.290 361.400 233.480 361.870 ;
        RECT 233.600 361.860 233.810 362.300 ;
        RECT 233.840 361.990 234.160 362.300 ;
        RECT 234.400 362.070 234.630 362.170 ;
        RECT 233.580 361.660 233.810 361.860 ;
        RECT 234.320 361.750 234.640 362.070 ;
        RECT 233.580 361.570 234.060 361.660 ;
        RECT 228.590 358.970 228.820 361.120 ;
        RECT 230.870 361.010 231.210 361.230 ;
        RECT 230.870 360.580 231.210 360.800 ;
        RECT 230.860 360.480 231.210 360.580 ;
        RECT 231.370 360.550 231.570 361.260 ;
        RECT 233.220 361.080 233.480 361.400 ;
        RECT 233.740 361.340 234.060 361.570 ;
        RECT 234.400 361.420 234.590 361.750 ;
        RECT 234.880 361.550 235.070 363.280 ;
        RECT 235.110 361.630 235.830 364.590 ;
        RECT 235.090 361.550 235.830 361.630 ;
        RECT 234.270 361.390 234.590 361.420 ;
        RECT 234.230 361.100 234.590 361.390 ;
        RECT 234.860 361.360 235.830 361.550 ;
        RECT 234.860 361.260 235.090 361.360 ;
        RECT 234.230 361.070 234.490 361.100 ;
        RECT 230.860 360.290 231.090 360.480 ;
        RECT 231.360 360.260 231.590 360.550 ;
        RECT 233.220 360.410 233.480 360.730 ;
        RECT 234.230 360.670 234.490 360.740 ;
        RECT 234.880 360.680 235.070 361.260 ;
        RECT 235.100 361.110 235.830 361.360 ;
        RECT 234.230 360.420 234.590 360.670 ;
        RECT 231.370 359.390 231.570 360.260 ;
        RECT 233.290 359.940 233.480 360.410 ;
        RECT 234.270 360.270 234.590 360.420 ;
        RECT 234.400 359.940 234.590 360.270 ;
        RECT 234.710 360.550 235.070 360.680 ;
        RECT 234.710 360.260 235.090 360.550 ;
        RECT 235.140 360.270 235.830 361.110 ;
        RECT 235.950 363.750 236.220 365.180 ;
        RECT 236.570 364.760 236.890 365.080 ;
        RECT 235.950 363.460 236.230 363.750 ;
        RECT 235.950 361.160 236.220 363.460 ;
        RECT 236.620 362.540 236.940 362.860 ;
        RECT 236.610 361.820 236.930 362.140 ;
        RECT 235.950 360.870 236.230 361.160 ;
        RECT 234.710 360.230 235.070 360.260 ;
        RECT 234.880 359.950 235.070 360.230 ;
        RECT 232.270 359.500 232.590 359.820 ;
        RECT 233.270 359.650 233.500 359.940 ;
        RECT 233.840 359.780 234.160 359.820 ;
        RECT 233.750 359.500 234.160 359.780 ;
        RECT 234.320 359.620 234.640 359.940 ;
        RECT 234.710 359.510 235.070 359.950 ;
        RECT 233.750 359.480 234.070 359.500 ;
        RECT 234.880 359.480 235.070 359.510 ;
        RECT 235.140 359.950 235.910 360.270 ;
        RECT 235.140 359.480 235.830 359.950 ;
        RECT 233.750 359.420 235.830 359.480 ;
        RECT 233.800 359.340 235.830 359.420 ;
        RECT 231.150 359.220 231.340 359.330 ;
        RECT 231.590 359.250 231.870 359.330 ;
        RECT 228.590 358.180 228.850 358.970 ;
        RECT 231.590 358.950 231.910 359.250 ;
        RECT 233.340 358.960 233.660 359.280 ;
        RECT 235.140 359.080 235.830 359.340 ;
        RECT 235.950 359.300 236.220 360.870 ;
        RECT 236.530 359.570 236.850 359.890 ;
        RECT 235.940 359.150 236.220 359.300 ;
        RECT 233.740 358.580 234.060 358.900 ;
        RECT 234.320 358.680 234.640 359.000 ;
        RECT 235.100 358.830 235.830 359.080 ;
        RECT 235.090 358.560 235.830 358.830 ;
        RECT 228.590 357.070 228.820 358.180 ;
        RECT 233.490 358.130 233.810 358.450 ;
        RECT 234.270 358.030 234.590 358.350 ;
        RECT 232.380 357.600 232.700 357.920 ;
        RECT 233.590 357.450 233.900 357.890 ;
        RECT 233.600 357.440 233.810 357.450 ;
        RECT 233.580 357.120 233.840 357.440 ;
        RECT 234.270 357.200 234.590 357.520 ;
        RECT 227.200 335.820 227.430 357.070 ;
        RECT 233.110 356.320 233.430 356.640 ;
        RECT 233.600 355.830 233.810 357.120 ;
        RECT 235.110 357.070 235.830 358.560 ;
        RECT 235.950 357.720 236.220 359.150 ;
        RECT 236.570 358.730 236.890 359.050 ;
        RECT 235.950 357.430 236.230 357.720 ;
        RECT 234.320 356.550 234.640 356.870 ;
        RECT 233.580 355.540 233.810 355.830 ;
        RECT 234.320 355.720 234.640 356.040 ;
        RECT 234.270 355.070 234.590 355.390 ;
        RECT 234.270 354.240 234.590 354.560 ;
        RECT 233.770 353.450 234.100 353.740 ;
        RECT 234.320 353.590 234.640 353.910 ;
        RECT 235.280 353.450 235.620 357.070 ;
        RECT 233.760 353.310 235.620 353.450 ;
        RECT 231.150 353.250 231.340 353.300 ;
        RECT 231.590 353.250 231.870 353.300 ;
        RECT 235.280 353.250 235.620 353.310 ;
        RECT 235.950 355.130 236.220 357.430 ;
        RECT 236.620 356.510 236.940 356.830 ;
        RECT 236.610 355.790 236.930 356.110 ;
        RECT 237.800 355.570 238.510 374.570 ;
        RECT 255.380 371.370 259.730 375.070 ;
        RECT 284.930 370.890 288.160 375.470 ;
        RECT 284.630 366.840 288.180 370.890 ;
        RECT 313.520 365.260 316.750 375.470 ;
        RECT 313.320 362.730 316.910 365.260 ;
        RECT 342.110 361.770 345.340 375.470 ;
        RECT 362.540 368.530 363.310 368.550 ;
        RECT 365.140 368.530 369.440 377.590 ;
        RECT 362.540 366.780 371.840 368.530 ;
        RECT 362.540 366.770 372.790 366.780 ;
        RECT 362.540 366.420 372.940 366.770 ;
        RECT 362.540 366.410 372.790 366.420 ;
        RECT 362.540 364.630 371.840 366.410 ;
        RECT 362.540 364.620 371.470 364.630 ;
        RECT 362.540 364.600 363.310 364.620 ;
        RECT 341.800 358.150 345.560 361.770 ;
        RECT 356.150 361.120 359.560 361.400 ;
        RECT 356.150 361.080 360.270 361.120 ;
        RECT 356.150 357.850 362.790 361.080 ;
        RECT 235.950 354.840 236.230 355.130 ;
        RECT 235.950 353.250 236.220 354.840 ;
        RECT 237.670 354.780 238.510 355.570 ;
        RECT 236.530 353.540 236.850 353.860 ;
        RECT 233.390 336.740 234.110 337.310 ;
        RECT 227.200 335.590 227.440 335.820 ;
        RECT 227.200 329.780 227.430 335.590 ;
        RECT 233.450 329.730 233.960 336.740 ;
        RECT 233.310 329.680 233.960 329.730 ;
        RECT 233.300 329.500 233.960 329.680 ;
        RECT 233.270 329.490 233.960 329.500 ;
        RECT 233.270 329.120 233.870 329.490 ;
        RECT 233.270 327.250 233.850 329.120 ;
        RECT 264.470 327.690 268.890 357.800 ;
        RECT 356.150 357.360 360.270 357.850 ;
        RECT 359.560 357.160 360.270 357.360 ;
        RECT 364.860 354.910 370.010 364.620 ;
        RECT 372.820 360.070 373.410 363.680 ;
        RECT 371.470 359.780 373.410 360.070 ;
        RECT 364.860 354.240 370.000 354.910 ;
        RECT 364.600 350.340 368.020 350.390 ;
        RECT 364.590 349.770 368.030 350.340 ;
        RECT 362.740 348.950 363.460 349.500 ;
        RECT 362.960 348.940 363.460 348.950 ;
        RECT 362.540 339.940 363.310 339.960 ;
        RECT 365.140 339.940 369.440 349.000 ;
        RECT 362.540 338.190 371.840 339.940 ;
        RECT 362.540 338.180 372.790 338.190 ;
        RECT 362.540 337.830 372.940 338.180 ;
        RECT 362.540 337.820 372.790 337.830 ;
        RECT 362.540 336.040 371.840 337.820 ;
        RECT 362.540 336.030 371.470 336.040 ;
        RECT 362.540 336.010 363.310 336.030 ;
        RECT 347.740 332.490 350.060 332.570 ;
        RECT 359.550 332.490 360.250 332.520 ;
        RECT 347.740 329.260 362.780 332.490 ;
        RECT 347.740 329.200 350.060 329.260 ;
        RECT 359.550 328.560 360.250 329.260 ;
        RECT 232.920 326.260 233.850 327.250 ;
        RECT 264.440 326.370 268.910 327.690 ;
        RECT 233.270 325.480 233.850 326.260 ;
        RECT 233.280 324.870 233.850 325.480 ;
        RECT 233.270 323.870 233.850 324.870 ;
        RECT 227.460 323.110 227.780 323.430 ;
        RECT 233.280 323.270 233.850 323.870 ;
        RECT 227.460 322.440 227.780 322.760 ;
        RECT 227.580 321.470 227.900 321.520 ;
        RECT 227.350 321.240 227.900 321.470 ;
        RECT 227.580 321.200 227.900 321.240 ;
        RECT 227.580 319.860 227.900 319.910 ;
        RECT 227.350 319.630 227.900 319.860 ;
        RECT 227.580 319.590 227.900 319.630 ;
        RECT 227.570 318.250 227.890 318.300 ;
        RECT 227.340 318.020 227.890 318.250 ;
        RECT 227.570 317.980 227.890 318.020 ;
        RECT 225.090 316.350 225.680 316.570 ;
        RECT 225.830 316.380 226.270 316.840 ;
        RECT 227.570 316.630 227.890 316.680 ;
        RECT 227.340 316.400 227.890 316.630 ;
        RECT 227.570 316.360 227.890 316.400 ;
        RECT 225.090 316.340 225.380 316.350 ;
        RECT 221.950 315.840 222.240 316.070 ;
        RECT 221.960 314.470 222.190 315.840 ;
        RECT 233.270 315.830 233.850 323.270 ;
        RECT 233.280 315.230 233.850 315.830 ;
        RECT 227.570 315.020 227.890 315.070 ;
        RECT 227.340 314.790 227.890 315.020 ;
        RECT 227.570 314.750 227.890 314.790 ;
        RECT 221.950 314.240 222.240 314.470 ;
        RECT 233.270 314.410 233.850 315.230 ;
        RECT 233.270 314.400 233.810 314.410 ;
        RECT 186.790 312.800 187.710 313.530 ;
        RECT 221.960 312.850 222.190 314.240 ;
        RECT 227.200 313.150 227.520 313.470 ;
        RECT 227.250 312.920 227.480 313.150 ;
        RECT 186.760 312.070 187.680 312.800 ;
        RECT 221.950 312.620 222.240 312.850 ;
        RECT 1.570 310.320 10.870 312.070 ;
        RECT 227.580 311.820 227.900 311.870 ;
        RECT 227.350 311.590 227.900 311.820 ;
        RECT 227.580 311.550 227.900 311.590 ;
        RECT 0.620 310.310 10.870 310.320 ;
        RECT 0.470 309.960 10.870 310.310 ;
        RECT 227.570 310.230 227.890 310.280 ;
        RECT 224.370 310.150 224.690 310.200 ;
        RECT 225.310 310.150 225.630 310.200 ;
        RECT 0.620 309.950 10.870 309.960 ;
        RECT 1.570 308.170 10.870 309.950 ;
        RECT 224.140 309.920 224.690 310.150 ;
        RECT 225.080 309.920 225.630 310.150 ;
        RECT 226.260 310.090 226.580 310.140 ;
        RECT 224.370 309.880 224.690 309.920 ;
        RECT 225.310 309.880 225.630 309.920 ;
        RECT 226.030 309.860 226.580 310.090 ;
        RECT 227.340 310.000 227.890 310.230 ;
        RECT 227.570 309.960 227.890 310.000 ;
        RECT 226.260 309.820 226.580 309.860 ;
        RECT 1.940 308.160 10.870 308.170 ;
        RECT 0.000 303.610 0.590 307.220 ;
        RECT 0.000 303.320 1.940 303.610 ;
        RECT 3.400 298.450 8.550 308.160 ;
        RECT 10.100 308.140 10.870 308.160 ;
        RECT 27.840 304.620 30.070 304.700 ;
        RECT 10.570 301.390 30.070 304.620 ;
        RECT 13.160 300.680 13.800 301.390 ;
        RECT 27.840 301.240 30.070 301.390 ;
        RECT 3.410 297.780 8.550 298.450 ;
        RECT 5.390 293.880 8.810 293.930 ;
        RECT 5.380 293.310 8.820 293.880 ;
        RECT 3.970 283.480 8.270 292.540 ;
        RECT 9.950 292.490 10.670 293.040 ;
        RECT 9.950 292.480 10.450 292.490 ;
        RECT 10.100 283.480 10.870 283.500 ;
        RECT 1.570 281.730 10.870 283.480 ;
        RECT 0.620 281.720 10.870 281.730 ;
        RECT 0.470 281.370 10.870 281.720 ;
        RECT 0.620 281.360 10.870 281.370 ;
        RECT 1.570 279.580 10.870 281.360 ;
        RECT 1.940 279.570 10.870 279.580 ;
        RECT 0.000 275.020 0.590 278.630 ;
        RECT 0.000 274.730 1.940 275.020 ;
        RECT 3.400 269.860 8.550 279.570 ;
        RECT 10.100 279.550 10.870 279.570 ;
        RECT 13.150 276.030 13.790 276.040 ;
        RECT 32.350 276.030 34.760 276.130 ;
        RECT 10.560 272.800 34.760 276.030 ;
        RECT 13.150 272.100 13.790 272.800 ;
        RECT 32.350 272.700 34.760 272.800 ;
        RECT 3.410 269.190 8.550 269.860 ;
        RECT 5.390 265.290 8.810 265.340 ;
        RECT 5.380 264.720 8.820 265.290 ;
        RECT 3.970 254.890 8.270 263.950 ;
        RECT 9.950 263.900 10.670 264.450 ;
        RECT 9.950 263.890 10.450 263.900 ;
        RECT 10.100 254.890 10.870 254.910 ;
        RECT 1.570 253.140 10.870 254.890 ;
        RECT 0.620 253.130 10.870 253.140 ;
        RECT 0.470 252.780 10.870 253.130 ;
        RECT 0.620 252.770 10.870 252.780 ;
        RECT 1.570 250.990 10.870 252.770 ;
        RECT 1.940 250.980 10.870 250.990 ;
        RECT 0.000 246.430 0.590 250.040 ;
        RECT 0.000 246.140 1.940 246.430 ;
        RECT 3.400 241.270 8.550 250.980 ;
        RECT 10.100 250.960 10.870 250.980 ;
        RECT 13.160 247.440 13.800 247.460 ;
        RECT 36.910 247.440 39.180 247.510 ;
        RECT 10.570 244.210 39.180 247.440 ;
        RECT 13.160 243.520 13.800 244.210 ;
        RECT 36.910 244.110 39.180 244.210 ;
        RECT 3.410 240.600 8.550 241.270 ;
        RECT 5.390 236.700 8.810 236.750 ;
        RECT 5.380 236.130 8.820 236.700 ;
        RECT 3.970 226.300 8.270 235.360 ;
        RECT 9.950 235.310 10.670 235.860 ;
        RECT 9.950 235.300 10.450 235.310 ;
        RECT 10.100 226.300 10.870 226.320 ;
        RECT 1.570 224.550 10.870 226.300 ;
        RECT 0.620 224.540 10.870 224.550 ;
        RECT 0.470 224.190 10.870 224.540 ;
        RECT 0.620 224.180 10.870 224.190 ;
        RECT 1.570 222.400 10.870 224.180 ;
        RECT 1.940 222.390 10.870 222.400 ;
        RECT 0.000 217.840 0.590 221.450 ;
        RECT 0.000 217.550 1.940 217.840 ;
        RECT 3.400 212.680 8.550 222.390 ;
        RECT 10.100 222.370 10.870 222.390 ;
        RECT 13.150 218.850 13.790 218.870 ;
        RECT 41.270 218.850 43.520 218.910 ;
        RECT 10.560 215.620 43.520 218.850 ;
        RECT 13.150 214.930 13.790 215.620 ;
        RECT 41.270 215.540 43.520 215.620 ;
        RECT 3.410 212.010 8.550 212.680 ;
        RECT 5.390 208.110 8.810 208.160 ;
        RECT 5.380 207.540 8.820 208.110 ;
        RECT 3.970 197.710 8.270 206.770 ;
        RECT 9.950 206.720 10.670 207.270 ;
        RECT 9.950 206.710 10.450 206.720 ;
        RECT 10.100 197.710 10.870 197.730 ;
        RECT 1.570 195.960 10.870 197.710 ;
        RECT 0.620 195.950 10.870 195.960 ;
        RECT 0.470 195.600 10.870 195.950 ;
        RECT 0.620 195.590 10.870 195.600 ;
        RECT 1.570 193.810 10.870 195.590 ;
        RECT 1.940 193.800 10.870 193.810 ;
        RECT 0.000 189.250 0.590 192.860 ;
        RECT 0.000 188.960 1.940 189.250 ;
        RECT 3.400 184.090 8.550 193.800 ;
        RECT 10.100 193.780 10.870 193.800 ;
        RECT 13.150 190.260 13.790 190.280 ;
        RECT 45.590 190.260 47.840 190.370 ;
        RECT 10.560 187.030 47.990 190.260 ;
        RECT 13.150 186.340 13.790 187.030 ;
        RECT 45.590 186.920 47.840 187.030 ;
        RECT 3.410 183.420 8.550 184.090 ;
        RECT 5.390 179.520 8.810 179.570 ;
        RECT 5.380 178.950 8.820 179.520 ;
        RECT 3.970 169.120 8.270 178.180 ;
        RECT 9.950 178.130 10.670 178.680 ;
        RECT 9.950 178.120 10.450 178.130 ;
        RECT 10.100 169.120 10.870 169.140 ;
        RECT 1.570 167.370 10.870 169.120 ;
        RECT 0.620 167.360 10.870 167.370 ;
        RECT 0.470 167.010 10.870 167.360 ;
        RECT 0.620 167.000 10.870 167.010 ;
        RECT 1.570 165.220 10.870 167.000 ;
        RECT 1.940 165.210 10.870 165.220 ;
        RECT 0.000 160.660 0.590 164.270 ;
        RECT 0.000 160.370 1.940 160.660 ;
        RECT 3.400 155.500 8.550 165.210 ;
        RECT 10.100 165.190 10.870 165.210 ;
        RECT 264.470 165.070 268.890 326.370 ;
        RECT 364.860 326.320 370.010 336.030 ;
        RECT 372.820 331.480 373.410 335.090 ;
        RECT 371.470 331.190 373.410 331.480 ;
        RECT 364.860 325.650 370.000 326.320 ;
        RECT 364.600 321.750 368.020 321.800 ;
        RECT 364.590 321.180 368.030 321.750 ;
        RECT 362.740 320.360 363.460 320.910 ;
        RECT 362.960 320.350 363.460 320.360 ;
        RECT 362.540 311.350 363.310 311.370 ;
        RECT 365.140 311.350 369.440 320.410 ;
        RECT 362.540 309.600 371.840 311.350 ;
        RECT 362.540 309.590 372.790 309.600 ;
        RECT 362.540 309.240 372.940 309.590 ;
        RECT 362.540 309.230 372.790 309.240 ;
        RECT 362.540 307.450 371.840 309.230 ;
        RECT 362.540 307.440 371.470 307.450 ;
        RECT 362.540 307.420 363.310 307.440 ;
        RECT 343.570 303.900 345.930 304.030 ;
        RECT 359.570 303.900 360.270 303.930 ;
        RECT 343.570 300.670 362.800 303.900 ;
        RECT 343.570 300.570 345.930 300.670 ;
        RECT 359.570 299.970 360.270 300.670 ;
        RECT 364.860 297.730 370.010 307.440 ;
        RECT 372.820 302.890 373.410 306.500 ;
        RECT 371.470 302.600 373.410 302.890 ;
        RECT 364.860 297.060 370.000 297.730 ;
        RECT 364.600 293.160 368.020 293.210 ;
        RECT 364.590 292.590 368.030 293.160 ;
        RECT 362.740 291.770 363.460 292.320 ;
        RECT 362.960 291.760 363.460 291.770 ;
        RECT 362.540 282.760 363.310 282.780 ;
        RECT 365.140 282.760 369.440 291.820 ;
        RECT 362.540 281.010 371.840 282.760 ;
        RECT 362.540 281.000 372.790 281.010 ;
        RECT 362.540 280.650 372.940 281.000 ;
        RECT 362.540 280.640 372.790 280.650 ;
        RECT 362.540 278.860 371.840 280.640 ;
        RECT 362.540 278.850 371.470 278.860 ;
        RECT 362.540 278.830 363.310 278.850 ;
        RECT 339.560 275.310 341.840 275.470 ;
        RECT 359.550 275.310 360.250 275.340 ;
        RECT 339.560 272.080 362.780 275.310 ;
        RECT 339.560 271.970 341.840 272.080 ;
        RECT 359.550 271.380 360.250 272.080 ;
        RECT 364.860 269.140 370.010 278.850 ;
        RECT 372.820 274.300 373.410 277.910 ;
        RECT 371.470 274.010 373.410 274.300 ;
        RECT 364.860 268.470 370.000 269.140 ;
        RECT 364.600 264.570 368.020 264.620 ;
        RECT 364.590 264.000 368.030 264.570 ;
        RECT 362.740 263.180 363.460 263.730 ;
        RECT 362.960 263.170 363.460 263.180 ;
        RECT 362.540 254.170 363.310 254.190 ;
        RECT 365.140 254.170 369.440 263.230 ;
        RECT 362.540 252.420 371.840 254.170 ;
        RECT 362.540 252.410 372.790 252.420 ;
        RECT 362.540 252.060 372.940 252.410 ;
        RECT 362.540 252.050 372.790 252.060 ;
        RECT 362.540 250.270 371.840 252.050 ;
        RECT 362.540 250.260 371.470 250.270 ;
        RECT 362.540 250.240 363.310 250.260 ;
        RECT 335.260 246.720 337.680 246.840 ;
        RECT 359.550 246.720 360.250 246.740 ;
        RECT 335.260 243.490 362.780 246.720 ;
        RECT 335.260 243.330 337.680 243.490 ;
        RECT 359.550 242.780 360.250 243.490 ;
        RECT 364.860 240.550 370.010 250.260 ;
        RECT 372.820 245.710 373.410 249.320 ;
        RECT 371.470 245.420 373.410 245.710 ;
        RECT 364.860 239.880 370.000 240.550 ;
        RECT 369.830 237.030 370.820 237.040 ;
        RECT 369.830 236.510 371.220 237.030 ;
        RECT 364.600 235.980 368.020 236.030 ;
        RECT 364.590 235.410 368.030 235.980 ;
        RECT 362.740 234.590 363.460 235.140 ;
        RECT 362.960 234.580 363.460 234.590 ;
        RECT 362.540 225.580 363.310 225.600 ;
        RECT 365.140 225.580 369.440 234.640 ;
        RECT 370.730 232.900 371.220 236.510 ;
        RECT 362.540 223.830 371.840 225.580 ;
        RECT 362.540 223.820 372.790 223.830 ;
        RECT 362.540 223.470 372.940 223.820 ;
        RECT 362.540 223.460 372.790 223.470 ;
        RECT 362.540 221.680 371.840 223.460 ;
        RECT 362.540 221.670 371.470 221.680 ;
        RECT 362.540 221.650 363.310 221.670 ;
        RECT 331.370 218.130 333.640 218.240 ;
        RECT 359.560 218.130 360.260 218.160 ;
        RECT 331.370 214.900 362.790 218.130 ;
        RECT 331.370 214.770 333.640 214.900 ;
        RECT 359.560 214.200 360.260 214.900 ;
        RECT 364.860 211.960 370.010 221.670 ;
        RECT 372.820 217.120 373.410 220.730 ;
        RECT 371.470 216.830 373.410 217.120 ;
        RECT 371.830 213.280 373.080 213.290 ;
        RECT 364.860 211.290 370.000 211.960 ;
        RECT 371.110 211.930 373.080 213.280 ;
        RECT 370.670 211.870 373.080 211.930 ;
        RECT 370.650 211.290 373.080 211.870 ;
        RECT 370.670 210.540 373.080 211.290 ;
        RECT 363.040 209.820 373.080 210.540 ;
        RECT 368.710 209.590 373.080 209.820 ;
        RECT 370.670 209.560 373.080 209.590 ;
        RECT 371.110 209.400 373.080 209.560 ;
        RECT 371.110 209.390 371.830 209.400 ;
        RECT 369.830 208.440 370.820 208.450 ;
        RECT 369.830 207.920 371.220 208.440 ;
        RECT 364.600 207.390 368.020 207.440 ;
        RECT 364.590 206.820 368.030 207.390 ;
        RECT 362.740 206.000 363.460 206.550 ;
        RECT 362.960 205.990 363.460 206.000 ;
        RECT 362.540 196.990 363.310 197.010 ;
        RECT 365.140 196.990 369.440 206.050 ;
        RECT 370.730 204.310 371.220 207.920 ;
        RECT 362.540 195.240 371.840 196.990 ;
        RECT 362.540 195.230 372.790 195.240 ;
        RECT 362.540 194.880 372.940 195.230 ;
        RECT 362.540 194.870 372.790 194.880 ;
        RECT 362.540 193.090 371.840 194.870 ;
        RECT 362.540 193.080 371.470 193.090 ;
        RECT 362.540 193.060 363.310 193.080 ;
        RECT 326.970 189.540 329.270 189.620 ;
        RECT 359.560 189.540 360.260 189.560 ;
        RECT 326.970 186.310 362.790 189.540 ;
        RECT 326.970 186.210 329.270 186.310 ;
        RECT 359.560 185.600 360.260 186.310 ;
        RECT 364.860 183.370 370.010 193.080 ;
        RECT 372.820 188.530 373.410 192.140 ;
        RECT 371.470 188.240 373.410 188.530 ;
        RECT 364.860 182.700 370.000 183.370 ;
        RECT 371.110 183.340 373.080 184.680 ;
        RECT 370.670 183.280 373.080 183.340 ;
        RECT 370.650 182.700 373.080 183.280 ;
        RECT 370.670 181.950 373.080 182.700 ;
        RECT 363.040 181.230 373.080 181.950 ;
        RECT 368.710 181.000 373.080 181.230 ;
        RECT 370.670 180.970 373.080 181.000 ;
        RECT 371.110 180.790 373.080 180.970 ;
        RECT 13.150 161.670 13.790 161.680 ;
        RECT 49.650 161.670 52.060 161.770 ;
        RECT 10.560 158.440 52.060 161.670 ;
        RECT 263.550 161.330 268.890 165.070 ;
        RECT 263.550 160.370 268.310 161.330 ;
        RECT 13.150 157.740 13.790 158.440 ;
        RECT 49.650 158.260 52.060 158.440 ;
        RECT 3.410 154.830 8.550 155.500 ;
        RECT 5.390 150.930 8.810 150.980 ;
        RECT 5.380 150.360 8.820 150.930 ;
        RECT 3.970 140.530 8.270 149.590 ;
        RECT 9.950 149.540 10.670 150.090 ;
        RECT 9.950 149.530 10.450 149.540 ;
        RECT 10.100 140.530 10.870 140.550 ;
        RECT 1.570 138.780 10.870 140.530 ;
        RECT 0.620 138.770 10.870 138.780 ;
        RECT 0.470 138.420 10.870 138.770 ;
        RECT 0.620 138.410 10.870 138.420 ;
        RECT 1.570 136.630 10.870 138.410 ;
        RECT 1.940 136.620 10.870 136.630 ;
        RECT 0.000 132.070 0.590 135.680 ;
        RECT 0.000 131.780 1.940 132.070 ;
        RECT 3.400 126.910 8.550 136.620 ;
        RECT 10.100 136.600 10.870 136.620 ;
        RECT 13.150 133.080 13.790 133.090 ;
        RECT 53.930 133.080 56.390 133.150 ;
        RECT 10.560 129.850 56.390 133.080 ;
        RECT 13.150 129.150 13.790 129.850 ;
        RECT 53.930 129.800 56.390 129.850 ;
        RECT 3.410 126.240 8.550 126.910 ;
        RECT 5.390 122.340 8.810 122.390 ;
        RECT 5.380 121.770 8.820 122.340 ;
        RECT 3.970 111.940 8.270 121.000 ;
        RECT 9.950 120.950 10.670 121.500 ;
        RECT 9.950 120.940 10.450 120.950 ;
        RECT 10.100 111.940 10.870 111.960 ;
        RECT 1.570 110.190 10.870 111.940 ;
        RECT 0.620 110.180 10.870 110.190 ;
        RECT 0.470 109.830 10.870 110.180 ;
        RECT 0.620 109.820 10.870 109.830 ;
        RECT 1.570 108.040 10.870 109.820 ;
        RECT 1.940 108.030 10.870 108.040 ;
        RECT 0.000 103.480 0.590 107.090 ;
        RECT 0.000 103.190 1.940 103.480 ;
        RECT 3.400 98.320 8.550 108.030 ;
        RECT 10.100 108.010 10.870 108.030 ;
        RECT 13.140 104.490 13.780 104.520 ;
        RECT 58.300 104.490 60.700 104.630 ;
        RECT 10.550 101.260 60.700 104.490 ;
        RECT 13.140 100.580 13.780 101.260 ;
        RECT 58.300 101.160 60.700 101.260 ;
        RECT 3.410 97.650 8.550 98.320 ;
        RECT 5.390 93.750 8.810 93.800 ;
        RECT 5.380 93.180 8.820 93.750 ;
        RECT 3.970 83.350 8.270 92.410 ;
        RECT 9.950 92.360 10.670 92.910 ;
        RECT 9.950 92.350 10.450 92.360 ;
        RECT 10.100 83.350 10.870 83.370 ;
        RECT 1.570 81.600 10.870 83.350 ;
        RECT 0.620 81.590 10.870 81.600 ;
        RECT 0.470 81.240 10.870 81.590 ;
        RECT 0.620 81.230 10.870 81.240 ;
        RECT 1.570 79.450 10.870 81.230 ;
        RECT 1.940 79.440 10.870 79.450 ;
        RECT 0.000 74.890 0.590 78.500 ;
        RECT 0.000 74.600 1.940 74.890 ;
        RECT 3.400 69.730 8.550 79.440 ;
        RECT 10.100 79.420 10.870 79.440 ;
        RECT 13.140 75.900 13.780 75.920 ;
        RECT 62.240 75.900 64.730 75.980 ;
        RECT 10.550 72.670 64.730 75.900 ;
        RECT 13.140 71.980 13.780 72.670 ;
        RECT 62.240 72.480 64.730 72.670 ;
        RECT 3.410 69.060 8.550 69.730 ;
        RECT 5.390 65.160 8.810 65.210 ;
        RECT 5.380 64.590 8.820 65.160 ;
        RECT 3.970 54.760 8.270 63.820 ;
        RECT 9.950 63.770 10.670 64.320 ;
        RECT 9.950 63.760 10.450 63.770 ;
        RECT 10.100 54.760 10.870 54.780 ;
        RECT 1.570 53.010 10.870 54.760 ;
        RECT 0.620 53.000 10.870 53.010 ;
        RECT 0.470 52.650 10.870 53.000 ;
        RECT 0.620 52.640 10.870 52.650 ;
        RECT 1.570 50.860 10.870 52.640 ;
        RECT 1.940 50.850 10.870 50.860 ;
        RECT 0.000 46.300 0.590 49.910 ;
        RECT 0.000 46.010 1.940 46.300 ;
        RECT 3.400 41.140 8.550 50.850 ;
        RECT 10.100 50.830 10.870 50.850 ;
        RECT 13.160 47.310 13.800 47.320 ;
        RECT 66.710 47.310 69.060 47.410 ;
        RECT 10.570 44.080 69.060 47.310 ;
        RECT 13.160 43.380 13.800 44.080 ;
        RECT 66.710 43.950 69.060 44.080 ;
        RECT 3.410 40.470 8.550 41.140 ;
        RECT 5.390 36.570 8.810 36.620 ;
        RECT 5.380 36.000 8.820 36.570 ;
        RECT 3.970 26.170 8.270 35.230 ;
        RECT 9.950 35.180 10.670 35.730 ;
        RECT 9.950 35.170 10.450 35.180 ;
        RECT 10.100 26.170 10.870 26.190 ;
        RECT 1.570 24.420 10.870 26.170 ;
        RECT 0.620 24.410 10.870 24.420 ;
        RECT 0.470 24.060 10.870 24.410 ;
        RECT 0.620 24.050 10.870 24.060 ;
        RECT 1.570 22.270 10.870 24.050 ;
        RECT 1.940 22.260 10.870 22.270 ;
        RECT 0.000 17.710 0.590 21.320 ;
        RECT 0.000 17.420 1.940 17.710 ;
        RECT 3.400 12.550 8.550 22.260 ;
        RECT 10.100 22.240 10.870 22.260 ;
        RECT 13.160 18.720 13.800 18.750 ;
        RECT 70.710 18.720 73.420 18.780 ;
        RECT 10.570 15.490 73.420 18.720 ;
        RECT 13.160 14.810 13.800 15.490 ;
        RECT 70.710 15.370 73.420 15.490 ;
        RECT 3.410 11.880 8.550 12.550 ;
      LAYER via ;
        RECT 24.250 386.810 26.280 387.140 ;
        RECT 24.190 385.950 24.890 386.570 ;
        RECT 47.640 386.810 50.630 387.160 ;
        RECT 2.630 380.270 3.390 380.620 ;
        RECT 2.240 376.840 2.590 379.830 ;
        RECT 5.510 379.240 8.680 379.660 ;
        RECT 51.070 386.010 51.420 386.770 ;
        RECT 50.040 380.720 50.460 383.890 ;
        RECT 9.980 378.270 10.500 378.790 ;
        RECT 49.070 378.900 49.590 379.420 ;
        RECT 78.630 380.720 79.050 383.890 ;
        RECT 77.660 378.900 78.180 379.420 ;
        RECT 107.220 380.720 107.640 383.890 ;
        RECT 127.040 382.070 127.430 382.460 ;
        RECT 106.250 378.900 106.770 379.420 ;
        RECT 132.320 381.200 132.580 381.460 ;
        RECT 209.690 381.440 210.060 381.810 ;
        RECT 145.560 379.350 145.820 379.610 ;
        RECT 146.920 379.430 147.180 379.690 ;
        RECT 147.610 379.420 147.870 379.680 ;
        RECT 190.270 379.160 190.790 379.420 ;
        RECT 127.120 378.620 127.510 379.010 ;
        RECT 86.550 370.730 89.780 372.980 ;
        RECT 98.740 369.450 99.260 369.820 ;
        RECT 57.960 366.240 61.190 368.490 ;
        RECT 27.540 361.970 29.790 365.200 ;
        RECT 16.010 358.570 17.870 361.800 ;
        RECT 102.080 365.070 102.490 365.480 ;
        RECT 98.600 361.130 99.120 361.650 ;
        RECT 2.260 353.450 2.590 355.480 ;
        RECT 2.830 353.390 3.450 354.090 ;
        RECT 5.510 350.650 8.680 351.070 ;
        RECT 9.980 349.680 10.500 350.200 ;
        RECT 24.060 329.980 26.140 333.210 ;
        RECT 102.130 360.280 102.540 360.690 ;
        RECT 98.700 325.110 99.220 325.630 ;
        RECT 102.130 324.170 102.540 324.610 ;
        RECT 5.510 322.060 8.680 322.480 ;
        RECT 9.980 321.090 10.500 321.610 ;
        RECT 189.800 378.740 191.150 379.160 ;
        RECT 171.700 377.130 172.140 377.570 ;
        RECT 167.280 376.110 167.720 376.550 ;
        RECT 177.420 377.130 177.860 377.570 ;
        RECT 172.990 376.110 173.430 376.550 ;
        RECT 144.840 375.690 145.100 375.950 ;
        RECT 154.700 375.710 154.960 375.970 ;
        RECT 164.520 373.090 164.780 373.350 ;
        RECT 140.840 367.950 141.100 368.210 ;
        RECT 141.930 367.960 142.190 368.220 ;
        RECT 140.370 367.540 140.630 367.800 ;
        RECT 140.840 367.030 141.100 367.290 ;
        RECT 141.930 367.040 142.190 367.300 ;
        RECT 140.370 366.620 140.630 366.880 ;
        RECT 140.840 366.110 141.100 366.370 ;
        RECT 140.370 365.700 140.630 365.960 ;
        RECT 141.580 366.040 141.840 366.300 ;
        RECT 141.930 366.120 142.190 366.380 ;
        RECT 140.650 365.130 140.910 365.390 ;
        RECT 141.550 365.120 141.810 365.380 ;
        RECT 140.650 364.670 140.910 364.930 ;
        RECT 141.950 365.030 142.210 365.290 ;
        RECT 140.650 364.170 140.910 364.430 ;
        RECT 141.560 364.200 141.820 364.460 ;
        RECT 140.650 363.710 140.910 363.970 ;
        RECT 140.650 363.440 140.910 363.470 ;
        RECT 140.650 363.210 141.170 363.440 ;
        RECT 140.910 363.180 141.170 363.210 ;
        RECT 140.650 362.750 140.910 363.010 ;
        RECT 140.870 362.220 141.130 362.480 ;
        RECT 140.910 361.260 141.170 361.520 ;
        RECT 141.950 364.070 142.210 364.330 ;
        RECT 141.950 363.110 142.210 363.370 ;
        RECT 144.950 370.630 145.300 370.980 ;
        RECT 163.470 369.340 163.730 369.600 ;
        RECT 145.970 368.390 146.230 368.780 ;
        RECT 162.370 368.400 162.700 368.660 ;
        RECT 145.330 367.570 145.590 367.970 ;
        RECT 145.350 366.460 145.610 366.720 ;
        RECT 145.350 365.540 145.610 365.800 ;
        RECT 145.320 364.620 145.580 364.880 ;
        RECT 140.870 345.980 141.130 346.450 ;
        RECT 141.510 345.980 141.770 346.450 ;
        RECT 139.510 344.950 139.770 345.210 ;
        RECT 138.990 344.550 139.250 344.810 ;
        RECT 129.710 343.300 130.370 343.960 ;
        RECT 141.590 344.930 141.850 345.190 ;
        RECT 143.350 344.940 143.620 345.210 ;
        RECT 140.930 344.570 141.190 344.830 ;
        RECT 141.680 343.970 141.940 344.230 ;
        RECT 142.330 343.970 142.590 344.230 ;
        RECT 140.460 343.530 140.720 343.790 ;
        RECT 141.160 343.530 141.420 343.790 ;
        RECT 142.840 342.800 143.100 343.060 ;
        RECT 140.010 342.180 140.270 342.440 ;
        RECT 139.010 340.640 139.270 340.900 ;
        RECT 134.920 338.780 135.290 339.150 ;
        RECT 129.750 337.440 130.410 338.100 ;
        RECT 139.010 337.550 139.270 337.810 ;
        RECT 142.760 341.670 143.020 341.930 ;
        RECT 143.850 344.550 144.110 344.810 ;
        RECT 142.770 341.130 143.030 341.390 ;
        RECT 140.010 340.630 140.270 340.890 ;
        RECT 142.820 340.180 143.080 340.440 ;
        RECT 140.490 339.650 140.750 339.910 ;
        RECT 141.180 339.640 141.440 339.900 ;
        RECT 141.660 338.870 141.920 339.130 ;
        RECT 142.370 338.810 142.630 339.070 ;
        RECT 142.320 337.990 142.580 338.250 ;
        RECT 140.110 337.560 140.370 337.820 ;
        RECT 141.200 337.560 141.460 337.820 ;
        RECT 142.330 337.520 142.590 337.780 ;
        RECT 139.560 336.880 139.820 337.140 ;
        RECT 140.660 336.880 140.920 337.140 ;
        RECT 141.760 336.880 142.020 337.140 ;
        RECT 139.560 335.510 139.820 335.770 ;
        RECT 140.660 335.510 140.920 335.770 ;
        RECT 141.760 335.510 142.020 335.770 ;
        RECT 139.010 334.780 139.270 335.040 ;
        RECT 140.110 334.780 140.370 335.040 ;
        RECT 141.200 334.780 141.460 335.040 ;
        RECT 139.000 333.440 139.260 333.700 ;
        RECT 140.110 333.430 140.370 333.690 ;
        RECT 141.200 333.410 141.460 333.670 ;
        RECT 134.910 332.540 135.280 332.910 ;
        RECT 139.560 332.740 139.820 333.000 ;
        RECT 140.660 332.730 140.920 332.990 ;
        RECT 141.750 332.730 142.010 332.990 ;
        RECT 142.450 332.120 142.710 332.480 ;
        RECT 141.610 330.430 141.870 330.690 ;
        RECT 138.300 329.990 138.560 330.250 ;
        RECT 139.400 330.000 139.660 330.260 ;
        RECT 140.490 330.000 140.750 330.260 ;
        RECT 141.620 329.960 141.880 330.220 ;
        RECT 138.850 329.320 139.110 329.580 ;
        RECT 139.950 329.320 140.210 329.580 ;
        RECT 141.050 329.320 141.310 329.580 ;
        RECT 138.850 327.950 139.110 328.210 ;
        RECT 139.950 327.950 140.210 328.210 ;
        RECT 141.050 327.950 141.310 328.210 ;
        RECT 138.300 327.220 138.560 327.480 ;
        RECT 139.400 327.220 139.660 327.480 ;
        RECT 140.490 327.220 140.750 327.480 ;
        RECT 137.900 326.880 138.190 327.170 ;
        RECT 161.740 366.680 162.070 367.010 ;
        RECT 161.170 365.200 161.500 365.530 ;
        RECT 145.960 363.530 146.220 363.790 ;
        RECT 160.530 363.600 160.860 363.930 ;
        RECT 159.890 363.030 160.220 363.360 ;
        RECT 145.970 362.570 146.230 362.830 ;
        RECT 145.960 361.610 146.220 361.870 ;
        RECT 145.320 343.950 145.580 344.210 ;
        RECT 144.700 342.800 144.960 343.060 ;
        RECT 144.280 340.190 144.540 340.450 ;
        RECT 144.720 334.500 144.980 334.920 ;
        RECT 144.680 332.120 144.940 332.480 ;
        RECT 159.280 361.460 159.610 361.790 ;
        RECT 158.650 359.930 158.980 360.260 ;
        RECT 158.090 358.360 158.420 358.690 ;
        RECT 157.470 352.890 157.800 353.220 ;
        RECT 156.840 351.300 157.170 351.630 ;
        RECT 156.220 349.750 156.550 350.080 ;
        RECT 155.620 348.270 155.950 348.600 ;
        RECT 154.980 343.100 155.310 343.430 ;
        RECT 154.310 341.530 154.640 341.860 ;
        RECT 145.960 339.620 146.220 339.880 ;
        RECT 153.690 339.890 154.020 340.220 ;
        RECT 145.300 328.490 145.560 328.820 ;
        RECT 144.270 326.870 144.560 327.160 ;
        RECT 138.290 325.880 138.550 326.140 ;
        RECT 139.400 325.870 139.660 326.130 ;
        RECT 140.490 325.850 140.750 326.110 ;
        RECT 143.110 325.860 143.710 326.460 ;
        RECT 138.850 325.180 139.110 325.440 ;
        RECT 139.950 325.170 140.210 325.430 ;
        RECT 141.040 325.170 141.300 325.430 ;
        RECT 153.010 338.450 153.340 338.780 ;
        RECT 148.970 334.090 149.550 334.800 ;
        RECT 145.890 320.930 146.150 321.270 ;
        RECT 126.980 319.990 127.370 320.380 ;
        RECT 152.980 314.620 153.410 315.050 ;
        RECT 153.630 313.830 154.060 314.260 ;
        RECT 154.300 313.150 154.700 313.550 ;
        RECT 154.130 312.210 154.640 312.720 ;
        RECT 163.470 367.790 163.730 368.050 ;
        RECT 163.470 366.240 163.730 366.500 ;
        RECT 165.570 370.180 165.830 370.440 ;
        RECT 170.430 370.280 170.690 370.540 ;
        RECT 165.570 368.630 165.830 368.890 ;
        RECT 165.570 367.080 165.830 367.340 ;
        RECT 165.570 365.530 165.830 365.790 ;
        RECT 167.610 369.460 167.870 369.720 ;
        RECT 170.430 368.730 170.690 368.990 ;
        RECT 167.610 367.910 167.870 368.170 ;
        RECT 170.430 367.180 170.690 367.440 ;
        RECT 167.610 366.360 167.870 366.620 ;
        RECT 170.430 365.630 170.690 365.890 ;
        RECT 163.470 364.690 163.730 364.950 ;
        RECT 167.610 364.810 167.870 365.070 ;
        RECT 187.390 376.110 187.830 376.550 ;
        RECT 181.640 372.330 181.900 372.590 ;
        RECT 179.760 368.800 180.020 369.060 ;
        RECT 185.230 371.420 185.490 371.680 ;
        RECT 182.100 370.400 182.360 370.660 ;
        RECT 182.520 368.310 182.780 368.570 ;
        RECT 183.580 367.830 183.840 368.090 ;
        RECT 188.400 372.340 188.660 372.600 ;
        RECT 187.960 371.430 188.220 371.690 ;
        RECT 184.390 362.750 184.650 363.010 ;
        RECT 163.470 362.070 163.730 362.330 ;
        RECT 163.470 360.520 163.730 360.780 ;
        RECT 163.470 358.970 163.730 359.230 ;
        RECT 163.470 357.420 163.730 357.680 ;
        RECT 165.570 361.230 165.830 361.490 ;
        RECT 165.570 359.680 165.830 359.940 ;
        RECT 165.570 358.130 165.830 358.390 ;
        RECT 167.610 361.950 167.870 362.210 ;
        RECT 183.300 362.230 183.560 362.490 ;
        RECT 170.430 361.130 170.690 361.390 ;
        RECT 167.610 360.400 167.870 360.660 ;
        RECT 170.430 359.580 170.690 359.840 ;
        RECT 167.610 358.850 167.870 359.110 ;
        RECT 170.430 358.030 170.690 358.290 ;
        RECT 167.610 357.300 167.870 357.560 ;
        RECT 165.570 356.580 165.830 356.840 ;
        RECT 170.430 356.480 170.690 356.740 ;
        RECT 183.300 361.130 183.560 361.390 ;
        RECT 193.190 376.070 193.630 376.510 ;
        RECT 201.520 377.100 201.800 377.540 ;
        RECT 197.740 370.440 198.960 370.700 ;
        RECT 194.500 369.790 194.760 370.050 ;
        RECT 200.830 369.250 201.090 369.510 ;
        RECT 203.170 372.340 203.430 372.600 ;
        RECT 202.280 371.470 202.540 371.730 ;
        RECT 219.830 380.720 220.250 383.890 ;
        RECT 218.860 378.900 219.380 379.420 ;
        RECT 205.840 373.050 206.100 373.320 ;
        RECT 202.280 367.260 202.540 367.520 ;
        RECT 203.300 367.270 203.560 367.530 ;
        RECT 207.380 368.360 207.640 368.620 ;
        RECT 206.050 367.150 206.480 367.580 ;
        RECT 206.990 366.830 207.250 367.090 ;
        RECT 206.280 366.000 206.540 366.260 ;
        RECT 206.980 365.140 207.240 365.400 ;
        RECT 186.800 362.750 187.060 363.010 ;
        RECT 184.390 360.610 184.650 360.870 ;
        RECT 185.220 360.730 185.490 361.000 ;
        RECT 184.390 359.820 184.650 360.080 ;
        RECT 183.300 359.300 183.560 359.560 ;
        RECT 183.300 358.200 183.560 358.460 ;
        RECT 184.390 357.680 184.650 357.940 ;
        RECT 186.800 360.610 187.060 360.870 ;
        RECT 186.800 359.820 187.060 360.080 ;
        RECT 186.800 357.680 187.060 357.940 ;
        RECT 207.380 363.630 207.640 363.890 ;
        RECT 248.420 380.720 248.840 383.890 ;
        RECT 210.510 377.980 210.880 378.350 ;
        RECT 209.370 365.030 209.630 365.290 ;
        RECT 207.380 362.330 207.640 362.590 ;
        RECT 207.230 361.370 207.490 361.630 ;
        RECT 206.290 360.260 206.550 360.520 ;
        RECT 206.290 359.660 206.550 359.920 ;
        RECT 209.420 358.980 209.680 359.240 ;
        RECT 207.230 358.610 207.490 358.870 ;
        RECT 192.690 356.550 192.950 356.810 ;
        RECT 192.690 356.000 192.950 356.260 ;
        RECT 181.860 354.090 182.140 354.370 ;
        RECT 192.690 355.120 192.950 355.380 ;
        RECT 184.390 352.680 184.650 352.940 ;
        RECT 163.470 351.940 163.730 352.200 ;
        RECT 163.470 350.390 163.730 350.650 ;
        RECT 163.470 348.840 163.730 349.100 ;
        RECT 163.470 347.290 163.730 347.550 ;
        RECT 165.570 351.100 165.830 351.360 ;
        RECT 165.570 349.550 165.830 349.810 ;
        RECT 165.570 348.000 165.830 348.260 ;
        RECT 167.610 351.820 167.870 352.080 ;
        RECT 183.300 352.160 183.560 352.420 ;
        RECT 170.430 351.000 170.690 351.260 ;
        RECT 167.610 350.270 167.870 350.530 ;
        RECT 170.430 349.450 170.690 349.710 ;
        RECT 167.610 348.720 167.870 348.980 ;
        RECT 170.430 347.900 170.690 348.160 ;
        RECT 167.610 347.170 167.870 347.430 ;
        RECT 165.570 346.450 165.830 346.710 ;
        RECT 170.430 346.350 170.690 346.610 ;
        RECT 183.300 351.060 183.560 351.320 ;
        RECT 184.390 350.540 184.650 350.800 ;
        RECT 184.390 349.750 184.650 350.010 ;
        RECT 183.300 349.230 183.560 349.490 ;
        RECT 183.300 348.130 183.560 348.390 ;
        RECT 184.390 347.610 184.650 347.870 ;
        RECT 174.490 345.900 174.750 346.310 ;
        RECT 186.800 352.680 187.060 352.940 ;
        RECT 192.690 354.570 192.950 354.830 ;
        RECT 192.690 353.540 192.950 353.800 ;
        RECT 192.690 352.990 192.950 353.250 ;
        RECT 193.380 353.070 193.640 353.330 ;
        RECT 193.610 352.510 193.870 352.770 ;
        RECT 186.800 350.540 187.060 350.800 ;
        RECT 192.690 352.120 192.950 352.380 ;
        RECT 192.690 351.570 192.950 351.830 ;
        RECT 207.380 357.600 207.640 357.860 ;
        RECT 199.210 353.520 199.470 353.780 ;
        RECT 197.540 352.470 197.800 352.730 ;
        RECT 247.450 378.900 247.970 379.420 ;
        RECT 277.010 380.720 277.430 383.890 ;
        RECT 211.280 373.270 211.650 373.640 ;
        RECT 209.700 354.070 210.070 354.440 ;
        RECT 210.470 353.480 210.840 353.850 ;
        RECT 208.620 352.470 208.880 352.730 ;
        RECT 217.830 372.220 218.330 372.720 ;
        RECT 214.610 370.660 215.110 371.160 ;
        RECT 215.560 371.150 216.060 371.650 ;
        RECT 216.640 371.620 217.140 372.120 ;
        RECT 212.160 368.200 212.530 368.570 ;
        RECT 214.490 361.780 214.750 362.040 ;
        RECT 214.520 358.090 214.780 358.350 ;
        RECT 213.470 356.550 213.730 356.810 ;
        RECT 213.470 356.000 213.730 356.260 ;
        RECT 213.470 355.120 213.730 355.380 ;
        RECT 213.470 354.570 213.730 354.830 ;
        RECT 213.470 353.540 213.730 353.800 ;
        RECT 211.210 351.150 211.580 351.520 ;
        RECT 186.800 349.750 187.060 350.010 ;
        RECT 184.390 342.920 184.650 343.180 ;
        RECT 163.470 342.170 163.730 342.430 ;
        RECT 163.470 340.620 163.730 340.880 ;
        RECT 163.470 339.070 163.730 339.330 ;
        RECT 163.470 337.520 163.730 337.780 ;
        RECT 165.570 341.330 165.830 341.590 ;
        RECT 165.570 339.780 165.830 340.040 ;
        RECT 165.570 338.230 165.830 338.490 ;
        RECT 167.610 342.050 167.870 342.310 ;
        RECT 178.890 342.180 179.150 342.440 ;
        RECT 183.300 342.400 183.560 342.660 ;
        RECT 170.430 341.230 170.690 341.490 ;
        RECT 167.610 340.500 167.870 340.760 ;
        RECT 170.430 339.680 170.690 339.940 ;
        RECT 167.610 338.950 167.870 339.210 ;
        RECT 170.430 338.130 170.690 338.390 ;
        RECT 167.610 337.400 167.870 337.660 ;
        RECT 165.570 336.680 165.830 336.940 ;
        RECT 172.310 337.050 172.570 337.310 ;
        RECT 170.430 336.580 170.690 336.840 ;
        RECT 171.770 336.680 172.060 336.970 ;
        RECT 167.330 336.170 167.640 336.480 ;
        RECT 183.300 341.300 183.560 341.560 ;
        RECT 184.390 340.780 184.650 341.040 ;
        RECT 179.520 339.400 179.780 339.660 ;
        RECT 178.920 337.090 179.180 337.350 ;
        RECT 179.950 337.080 180.210 337.340 ;
        RECT 177.520 336.680 177.780 336.940 ;
        RECT 179.490 336.760 179.750 337.020 ;
        RECT 171.140 335.460 171.560 335.880 ;
        RECT 167.290 334.500 167.710 334.920 ;
        RECT 173.200 336.140 173.460 336.400 ;
        RECT 184.390 339.990 184.650 340.250 ;
        RECT 183.300 339.470 183.560 339.730 ;
        RECT 183.300 338.370 183.560 338.630 ;
        RECT 184.390 337.850 184.650 338.110 ;
        RECT 181.730 336.700 181.990 336.960 ;
        RECT 180.530 335.450 180.860 335.780 ;
        RECT 186.800 347.610 187.060 347.870 ;
        RECT 186.800 342.920 187.060 343.180 ;
        RECT 193.270 347.160 193.530 347.420 ;
        RECT 193.270 346.610 193.530 346.870 ;
        RECT 193.270 345.730 193.530 345.990 ;
        RECT 193.270 345.180 193.530 345.440 ;
        RECT 193.270 344.150 193.530 344.410 ;
        RECT 193.270 343.600 193.530 343.860 ;
        RECT 212.780 353.070 213.040 353.330 ;
        RECT 213.470 352.990 213.730 353.250 ;
        RECT 212.550 352.510 212.810 352.770 ;
        RECT 213.470 352.120 213.730 352.380 ;
        RECT 213.470 351.570 213.730 351.830 ;
        RECT 196.540 343.450 196.800 343.710 ;
        RECT 194.310 343.080 194.570 343.340 ;
        RECT 193.270 342.730 193.530 342.990 ;
        RECT 193.270 342.180 193.530 342.440 ;
        RECT 193.250 341.900 193.510 342.160 ;
        RECT 186.800 340.780 187.060 341.040 ;
        RECT 198.330 343.060 198.600 343.320 ;
        RECT 196.520 342.400 196.780 342.660 ;
        RECT 198.770 342.160 199.030 342.420 ;
        RECT 198.250 341.230 198.510 341.490 ;
        RECT 193.230 340.890 193.490 341.150 ;
        RECT 196.520 340.520 196.780 340.780 ;
        RECT 186.800 339.990 187.060 340.250 ;
        RECT 196.360 339.340 196.620 339.600 ;
        RECT 197.780 339.390 198.040 339.650 ;
        RECT 193.180 338.850 193.440 339.110 ;
        RECT 186.800 337.850 187.060 338.110 ;
        RECT 197.280 338.460 197.540 338.720 ;
        RECT 193.230 338.000 193.490 338.260 ;
        RECT 190.570 337.010 190.920 337.360 ;
        RECT 183.720 336.280 183.980 336.540 ;
        RECT 187.760 336.250 188.030 336.520 ;
        RECT 181.680 335.380 182.020 335.720 ;
        RECT 190.610 335.240 190.870 335.560 ;
        RECT 196.600 335.460 196.860 335.800 ;
        RECT 171.820 334.410 172.140 334.730 ;
        RECT 192.030 334.530 192.410 334.910 ;
        RECT 172.720 331.280 172.980 331.540 ;
        RECT 173.810 331.280 174.070 331.540 ;
        RECT 174.910 331.270 175.170 331.530 ;
        RECT 177.530 331.270 177.790 331.530 ;
        RECT 178.630 331.280 178.890 331.540 ;
        RECT 179.720 331.280 179.980 331.540 ;
        RECT 182.530 331.310 182.790 331.570 ;
        RECT 183.620 331.310 183.880 331.570 ;
        RECT 184.720 331.300 184.980 331.560 ;
        RECT 187.340 331.300 187.600 331.560 ;
        RECT 188.440 331.310 188.700 331.570 ;
        RECT 189.530 331.310 189.790 331.570 ;
        RECT 193.830 331.280 194.090 331.540 ;
        RECT 194.930 331.290 195.190 331.550 ;
        RECT 196.020 331.290 196.280 331.550 ;
        RECT 173.270 330.600 173.530 330.860 ;
        RECT 174.360 330.580 174.620 330.840 ;
        RECT 175.470 330.570 175.730 330.830 ;
        RECT 175.840 329.660 176.120 329.940 ;
        RECT 173.270 329.230 173.530 329.490 ;
        RECT 174.360 329.230 174.620 329.490 ;
        RECT 175.460 329.230 175.720 329.490 ;
        RECT 171.920 328.630 172.380 329.090 ;
        RECT 172.710 328.500 172.970 328.760 ;
        RECT 173.810 328.500 174.070 328.760 ;
        RECT 174.910 328.500 175.170 328.760 ;
        RECT 176.970 330.570 177.230 330.830 ;
        RECT 178.080 330.580 178.340 330.840 ;
        RECT 179.170 330.600 179.430 330.860 ;
        RECT 176.580 329.680 176.860 329.960 ;
        RECT 176.980 329.230 177.240 329.490 ;
        RECT 178.080 329.230 178.340 329.490 ;
        RECT 179.170 329.230 179.430 329.490 ;
        RECT 177.530 328.500 177.790 328.760 ;
        RECT 178.630 328.500 178.890 328.760 ;
        RECT 179.730 328.500 179.990 328.760 ;
        RECT 172.710 327.130 172.970 327.390 ;
        RECT 173.810 327.130 174.070 327.390 ;
        RECT 174.910 327.130 175.170 327.390 ;
        RECT 172.140 326.490 172.400 326.750 ;
        RECT 173.270 326.450 173.530 326.710 ;
        RECT 174.360 326.450 174.620 326.710 ;
        RECT 175.460 326.460 175.720 326.720 ;
        RECT 172.150 326.020 172.410 326.280 ;
        RECT 180.300 327.680 180.760 328.140 ;
        RECT 177.530 327.130 177.790 327.390 ;
        RECT 178.630 327.130 178.890 327.390 ;
        RECT 179.730 327.130 179.990 327.390 ;
        RECT 183.080 330.630 183.340 330.890 ;
        RECT 184.170 330.610 184.430 330.870 ;
        RECT 185.280 330.600 185.540 330.860 ;
        RECT 185.650 329.660 185.930 329.940 ;
        RECT 183.080 329.260 183.340 329.520 ;
        RECT 184.170 329.260 184.430 329.520 ;
        RECT 185.270 329.260 185.530 329.520 ;
        RECT 182.520 328.530 182.780 328.790 ;
        RECT 183.620 328.530 183.880 328.790 ;
        RECT 184.720 328.530 184.980 328.790 ;
        RECT 186.780 330.600 187.040 330.860 ;
        RECT 187.890 330.610 188.150 330.870 ;
        RECT 188.980 330.630 189.240 330.890 ;
        RECT 186.790 329.260 187.050 329.520 ;
        RECT 187.890 329.260 188.150 329.520 ;
        RECT 188.980 329.260 189.240 329.520 ;
        RECT 187.340 328.530 187.600 328.790 ;
        RECT 188.440 328.530 188.700 328.790 ;
        RECT 189.540 328.530 189.800 328.790 ;
        RECT 181.730 326.790 182.190 327.250 ;
        RECT 182.520 327.160 182.780 327.420 ;
        RECT 183.620 327.160 183.880 327.420 ;
        RECT 184.720 327.160 184.980 327.420 ;
        RECT 176.980 326.460 177.240 326.720 ;
        RECT 178.080 326.450 178.340 326.710 ;
        RECT 179.170 326.450 179.430 326.710 ;
        RECT 180.300 326.490 180.560 326.750 ;
        RECT 181.950 326.520 182.210 326.780 ;
        RECT 183.080 326.480 183.340 326.740 ;
        RECT 184.170 326.480 184.430 326.740 ;
        RECT 185.270 326.490 185.530 326.750 ;
        RECT 180.290 326.020 180.550 326.280 ;
        RECT 181.960 326.050 182.220 326.310 ;
        RECT 187.340 327.160 187.600 327.420 ;
        RECT 188.440 327.160 188.700 327.420 ;
        RECT 189.540 327.160 189.800 327.420 ;
        RECT 193.270 330.580 193.530 330.840 ;
        RECT 194.380 330.590 194.640 330.850 ;
        RECT 195.470 330.610 195.730 330.870 ;
        RECT 212.140 345.900 212.510 346.310 ;
        RECT 204.620 343.250 204.880 343.510 ;
        RECT 204.770 342.570 205.030 342.830 ;
        RECT 204.770 341.680 205.030 341.940 ;
        RECT 204.620 341.000 204.880 341.260 ;
        RECT 204.620 340.480 204.880 340.740 ;
        RECT 204.770 339.800 205.030 340.060 ;
        RECT 204.770 338.910 205.030 339.170 ;
        RECT 204.620 338.230 204.880 338.490 ;
        RECT 206.900 339.350 207.170 339.620 ;
        RECT 226.640 369.280 227.920 370.560 ;
        RECT 223.130 362.640 223.530 363.040 ;
        RECT 217.590 359.350 217.850 359.610 ;
        RECT 224.110 362.000 224.470 362.360 ;
        RECT 223.390 359.350 223.650 359.610 ;
        RECT 217.660 355.910 217.920 356.170 ;
        RECT 217.740 349.940 218.240 350.440 ;
        RECT 216.660 344.750 217.160 345.220 ;
        RECT 215.530 339.560 216.030 340.060 ;
        RECT 214.480 334.260 214.980 334.760 ;
        RECT 198.750 332.750 199.010 333.250 ;
        RECT 198.210 331.850 198.470 332.350 ;
        RECT 197.740 330.950 198.000 331.450 ;
        RECT 193.280 329.240 193.540 329.500 ;
        RECT 194.380 329.240 194.640 329.500 ;
        RECT 195.470 329.240 195.730 329.500 ;
        RECT 197.260 330.050 197.520 330.550 ;
        RECT 193.830 328.510 194.090 328.770 ;
        RECT 194.930 328.510 195.190 328.770 ;
        RECT 196.030 328.510 196.290 328.770 ;
        RECT 193.830 327.140 194.090 327.400 ;
        RECT 194.930 327.140 195.190 327.400 ;
        RECT 196.030 327.140 196.290 327.400 ;
        RECT 186.790 326.490 187.050 326.750 ;
        RECT 187.890 326.480 188.150 326.740 ;
        RECT 188.980 326.480 189.240 326.740 ;
        RECT 190.110 326.520 190.370 326.780 ;
        RECT 193.280 326.470 193.540 326.730 ;
        RECT 194.380 326.460 194.640 326.720 ;
        RECT 195.470 326.460 195.730 326.720 ;
        RECT 190.120 326.310 190.580 326.340 ;
        RECT 190.100 326.050 190.580 326.310 ;
        RECT 190.120 325.880 190.580 326.050 ;
        RECT 164.050 323.650 164.310 324.770 ;
        RECT 176.160 324.710 177.280 324.730 ;
        RECT 175.420 323.610 177.280 324.710 ;
        RECT 175.420 323.590 176.540 323.610 ;
        RECT 185.230 323.560 187.090 324.750 ;
        RECT 162.370 319.360 162.700 319.690 ;
        RECT 161.750 318.740 162.080 319.070 ;
        RECT 161.120 318.110 161.450 318.440 ;
        RECT 160.520 317.480 160.850 317.810 ;
        RECT 159.880 316.800 160.210 317.130 ;
        RECT 159.280 316.180 159.610 316.510 ;
        RECT 158.680 315.540 159.010 315.870 ;
        RECT 158.100 314.970 158.430 315.300 ;
        RECT 157.520 314.280 157.850 314.610 ;
        RECT 156.870 313.640 157.200 313.970 ;
        RECT 156.230 312.990 156.560 313.330 ;
        RECT 155.650 312.350 156.020 312.720 ;
        RECT 196.600 326.500 196.860 326.760 ;
        RECT 223.360 355.850 223.620 356.110 ;
        RECT 223.360 353.330 223.620 353.590 ;
        RECT 220.720 336.780 221.220 337.280 ;
        RECT 217.850 328.670 218.350 329.170 ;
        RECT 216.660 327.720 217.160 328.180 ;
        RECT 215.530 326.850 216.030 327.310 ;
        RECT 196.590 326.030 196.850 326.290 ;
        RECT 214.600 325.940 215.100 326.400 ;
        RECT 220.140 323.650 221.080 324.770 ;
        RECT 195.930 320.020 196.260 320.350 ;
        RECT 227.130 365.840 227.390 366.260 ;
        RECT 225.030 359.630 225.420 360.020 ;
        RECT 225.860 359.070 226.240 359.330 ;
        RECT 223.190 318.830 223.590 319.230 ;
        RECT 222.710 317.900 222.970 318.160 ;
        RECT 224.100 318.030 224.490 318.420 ;
        RECT 225.030 317.210 225.420 317.600 ;
        RECT 233.620 368.360 233.880 368.620 ;
        RECT 230.960 367.120 231.220 367.550 ;
        RECT 233.770 367.400 234.030 367.660 ;
        RECT 276.040 378.900 276.560 379.420 ;
        RECT 305.600 380.720 306.020 383.890 ;
        RECT 304.630 378.900 305.150 379.420 ;
        RECT 334.190 380.720 334.610 383.890 ;
        RECT 333.220 378.900 333.740 379.420 ;
        RECT 362.780 380.720 363.200 383.890 ;
        RECT 361.810 378.900 362.330 379.420 ;
        RECT 364.730 378.520 367.900 378.940 ;
        RECT 362.910 377.550 363.430 378.070 ;
        RECT 237.910 374.610 238.620 375.320 ;
        RECT 234.710 366.290 234.970 366.550 ;
        RECT 234.710 365.690 234.970 365.950 ;
        RECT 231.640 365.030 231.900 365.290 ;
        RECT 232.300 365.040 232.560 365.300 ;
        RECT 233.370 365.020 233.630 365.280 ;
        RECT 233.870 365.040 234.130 365.300 ;
        RECT 230.950 364.060 231.210 364.320 ;
        RECT 233.770 364.640 234.030 364.900 ;
        RECT 234.350 364.740 234.610 365.000 ;
        RECT 230.950 363.530 231.210 363.790 ;
        RECT 233.220 364.130 233.480 364.390 ;
        RECT 233.520 364.190 233.780 364.450 ;
        RECT 235.650 366.010 235.910 366.270 ;
        RECT 234.230 364.350 234.490 364.380 ;
        RECT 234.230 364.120 234.560 364.350 ;
        RECT 234.300 364.090 234.560 364.120 ;
        RECT 232.410 363.660 232.670 363.920 ;
        RECT 233.220 363.460 233.480 363.720 ;
        RECT 233.620 363.630 233.880 363.890 ;
        RECT 234.230 363.520 234.490 363.730 ;
        RECT 234.230 363.470 234.560 363.520 ;
        RECT 233.580 363.180 233.840 363.440 ;
        RECT 234.300 363.260 234.560 363.470 ;
        RECT 232.300 362.550 232.560 362.810 ;
        RECT 233.140 362.380 233.400 362.640 ;
        RECT 233.870 362.590 234.130 362.810 ;
        RECT 233.620 362.550 234.130 362.590 ;
        RECT 234.350 362.610 234.610 362.870 ;
        RECT 233.620 362.330 233.880 362.550 ;
        RECT 232.300 362.020 232.560 362.280 ;
        RECT 230.950 361.040 231.210 361.300 ;
        RECT 233.870 362.020 234.130 362.280 ;
        RECT 234.350 361.780 234.610 362.040 ;
        RECT 230.950 360.510 231.210 360.770 ;
        RECT 233.220 361.110 233.480 361.370 ;
        RECT 233.770 361.370 234.030 361.630 ;
        RECT 234.300 361.360 234.560 361.390 ;
        RECT 234.230 361.130 234.560 361.360 ;
        RECT 233.220 360.440 233.480 360.700 ;
        RECT 234.230 360.560 234.490 360.710 ;
        RECT 234.230 360.450 234.560 360.560 ;
        RECT 234.300 360.300 234.560 360.450 ;
        RECT 236.600 364.790 236.860 365.050 ;
        RECT 236.650 362.570 236.910 362.830 ;
        RECT 236.640 361.850 236.900 362.110 ;
        RECT 232.300 359.530 232.560 359.790 ;
        RECT 233.870 359.760 234.130 359.790 ;
        RECT 233.780 359.530 234.130 359.760 ;
        RECT 234.350 359.650 234.610 359.910 ;
        RECT 234.710 359.660 234.970 359.920 ;
        RECT 233.780 359.500 234.040 359.530 ;
        RECT 235.650 359.980 235.910 360.240 ;
        RECT 231.620 358.970 231.880 359.230 ;
        RECT 233.370 358.990 233.630 359.250 ;
        RECT 236.560 359.600 236.820 359.860 ;
        RECT 233.770 358.610 234.030 358.870 ;
        RECT 234.350 358.710 234.610 358.970 ;
        RECT 233.520 358.160 233.780 358.420 ;
        RECT 234.300 358.060 234.560 358.320 ;
        RECT 232.410 357.630 232.670 357.890 ;
        RECT 233.620 357.600 233.880 357.860 ;
        RECT 233.580 357.150 233.840 357.410 ;
        RECT 234.300 357.230 234.560 357.490 ;
        RECT 233.140 356.350 233.400 356.610 ;
        RECT 236.600 358.760 236.860 359.020 ;
        RECT 234.350 356.580 234.610 356.840 ;
        RECT 234.350 355.750 234.610 356.010 ;
        RECT 234.300 355.100 234.560 355.360 ;
        RECT 234.300 354.270 234.560 354.530 ;
        RECT 233.800 353.460 234.070 353.720 ;
        RECT 234.350 353.620 234.610 353.880 ;
        RECT 236.650 356.540 236.910 356.800 ;
        RECT 236.640 355.820 236.900 356.080 ;
        RECT 256.340 372.040 259.570 374.100 ;
        RECT 284.930 367.150 286.990 370.450 ;
        RECT 313.520 362.900 316.750 364.960 ;
        RECT 342.110 358.490 345.340 360.540 ;
        RECT 356.450 357.850 358.440 361.080 ;
        RECT 237.720 354.820 238.430 355.530 ;
        RECT 264.710 356.870 266.930 357.190 ;
        RECT 236.560 353.570 236.820 353.830 ;
        RECT 233.520 336.770 234.030 337.280 ;
        RECT 364.730 349.930 367.900 350.350 ;
        RECT 362.910 348.960 363.430 349.480 ;
        RECT 347.900 329.260 349.990 332.490 ;
        RECT 264.550 326.480 268.830 327.570 ;
        RECT 227.490 323.140 227.750 323.400 ;
        RECT 227.490 322.470 227.750 322.730 ;
        RECT 227.610 321.230 227.870 321.490 ;
        RECT 227.610 319.620 227.870 319.880 ;
        RECT 227.600 318.010 227.860 318.270 ;
        RECT 225.850 316.420 226.230 316.800 ;
        RECT 227.600 316.390 227.860 316.650 ;
        RECT 227.600 314.780 227.860 315.040 ;
        RECT 227.230 313.180 227.490 313.440 ;
        RECT 227.610 311.580 227.870 311.840 ;
        RECT 224.400 309.910 224.660 310.170 ;
        RECT 225.340 309.910 225.600 310.170 ;
        RECT 226.290 309.850 226.550 310.110 ;
        RECT 227.600 309.990 227.860 310.250 ;
        RECT 27.960 301.390 30.040 304.620 ;
        RECT 5.510 293.470 8.680 293.890 ;
        RECT 9.980 292.500 10.500 293.020 ;
        RECT 32.590 272.800 34.670 276.030 ;
        RECT 5.510 264.880 8.680 265.300 ;
        RECT 9.980 263.910 10.500 264.430 ;
        RECT 37.000 244.210 39.080 247.440 ;
        RECT 5.510 236.290 8.680 236.710 ;
        RECT 9.980 235.320 10.500 235.840 ;
        RECT 41.340 215.620 43.420 218.850 ;
        RECT 5.510 207.700 8.680 208.120 ;
        RECT 9.980 206.730 10.500 207.250 ;
        RECT 5.510 179.110 8.680 179.530 ;
        RECT 9.980 178.140 10.500 178.660 ;
        RECT 364.730 321.340 367.900 321.760 ;
        RECT 362.910 320.370 363.430 320.890 ;
        RECT 343.650 300.670 345.740 303.900 ;
        RECT 364.730 292.750 367.900 293.170 ;
        RECT 362.910 291.780 363.430 292.300 ;
        RECT 339.670 272.080 341.760 275.310 ;
        RECT 364.730 264.160 367.900 264.580 ;
        RECT 362.910 263.190 363.430 263.710 ;
        RECT 335.420 243.490 337.510 246.720 ;
        RECT 370.020 236.600 370.780 236.950 ;
        RECT 364.730 235.570 367.900 235.990 ;
        RECT 362.910 234.600 363.430 235.120 ;
        RECT 370.820 233.170 371.170 236.160 ;
        RECT 331.480 214.900 333.570 218.130 ;
        RECT 369.960 209.720 370.580 210.420 ;
        RECT 370.820 209.780 371.150 211.810 ;
        RECT 370.020 208.010 370.780 208.360 ;
        RECT 364.730 206.980 367.900 207.400 ;
        RECT 362.910 206.010 363.430 206.530 ;
        RECT 370.820 204.580 371.170 207.570 ;
        RECT 369.960 181.130 370.580 181.830 ;
        RECT 370.820 181.190 371.150 183.220 ;
        RECT 49.880 158.440 51.960 161.670 ;
        RECT 263.730 160.540 268.150 164.960 ;
        RECT 5.510 150.520 8.680 150.940 ;
        RECT 9.980 149.550 10.500 150.070 ;
        RECT 5.510 121.930 8.680 122.350 ;
        RECT 9.980 120.960 10.500 121.480 ;
        RECT 58.500 101.260 60.580 104.490 ;
        RECT 5.510 93.340 8.680 93.760 ;
        RECT 9.980 92.370 10.500 92.890 ;
        RECT 62.470 72.670 64.550 75.900 ;
        RECT 5.510 64.750 8.680 65.170 ;
        RECT 9.980 63.780 10.500 64.300 ;
        RECT 66.910 44.080 68.990 47.310 ;
        RECT 5.510 36.160 8.680 36.580 ;
        RECT 9.980 35.190 10.500 35.710 ;
        RECT 71.210 15.490 73.290 18.720 ;
      LAYER met2 ;
        RECT 49.930 381.010 50.570 384.020 ;
        RECT 78.520 381.010 79.160 384.020 ;
        RECT 107.110 381.010 107.750 384.020 ;
        RECT 23.590 379.610 109.360 381.010 ;
        RECT 49.030 379.480 51.660 379.610 ;
        RECT 77.620 379.480 80.250 379.610 ;
        RECT 106.210 379.480 108.840 379.610 ;
        RECT 49.030 378.970 51.580 379.480 ;
        RECT 77.620 378.970 80.170 379.480 ;
        RECT 106.210 378.970 108.760 379.480 ;
        RECT 49.030 378.900 49.650 378.970 ;
        RECT 77.620 378.900 78.240 378.970 ;
        RECT 106.210 378.900 106.830 378.970 ;
        RECT 10.680 377.250 16.430 378.650 ;
        RECT 210.460 378.350 210.900 378.370 ;
        RECT 240.500 378.350 241.360 379.030 ;
        RECT 210.460 377.980 241.360 378.350 ;
        RECT 210.460 377.960 210.900 377.980 ;
        RECT 10.680 372.530 12.080 377.250 ;
        RECT 240.500 376.930 241.360 377.980 ;
        RECT 356.070 377.320 362.740 378.720 ;
        RECT 211.240 373.640 211.660 373.660 ;
        RECT 240.470 373.640 241.330 374.940 ;
        RECT 211.240 373.270 241.330 373.640 ;
        RECT 211.240 373.250 211.660 373.270 ;
        RECT 240.470 372.840 241.330 373.270 ;
        RECT 255.190 372.810 259.990 374.900 ;
        RECT 171.800 370.690 171.910 370.890 ;
        RECT 243.490 370.750 260.040 372.810 ;
        RECT 361.330 371.810 362.730 377.320 ;
        RECT 170.400 370.490 170.720 370.540 ;
        RECT 170.400 370.290 172.030 370.490 ;
        RECT 170.400 370.280 170.720 370.290 ;
        RECT 98.690 369.880 99.310 369.900 ;
        RECT 125.010 369.880 126.280 370.240 ;
        RECT 98.690 369.510 127.840 369.880 ;
        RECT 163.110 369.710 163.200 370.030 ;
        RECT 98.690 369.440 99.310 369.510 ;
        RECT 57.870 368.750 61.250 368.860 ;
        RECT 125.010 368.780 126.280 369.510 ;
        RECT 163.300 369.310 163.760 369.630 ;
        RECT 200.800 369.480 201.110 369.540 ;
        RECT 172.500 369.470 201.110 369.480 ;
        RECT 171.800 369.140 171.910 369.340 ;
        RECT 172.170 369.280 201.110 369.470 ;
        RECT 172.170 369.270 172.750 369.280 ;
        RECT 200.800 369.220 201.110 369.280 ;
        RECT 179.730 369.010 180.050 369.060 ;
        RECT 170.400 368.940 170.720 368.990 ;
        RECT 136.360 368.780 136.660 368.790 ;
        RECT 145.950 368.780 146.240 368.800 ;
        RECT 125.010 368.750 146.270 368.780 ;
        RECT 57.460 368.390 146.270 368.750 ;
        RECT 162.340 368.570 162.730 368.660 ;
        RECT 162.340 368.400 164.070 368.570 ;
        RECT 57.460 366.500 127.960 368.390 ;
        RECT 145.950 368.370 146.240 368.390 ;
        RECT 163.110 368.160 163.200 368.400 ;
        RECT 165.570 368.120 165.830 368.920 ;
        RECT 170.400 368.740 172.030 368.940 ;
        RECT 174.730 368.810 180.100 369.010 ;
        RECT 170.400 368.730 170.720 368.740 ;
        RECT 167.570 368.120 167.910 368.180 ;
        RECT 163.300 367.760 163.760 368.080 ;
        RECT 165.470 367.900 167.910 368.120 ;
        RECT 174.730 367.930 174.930 368.810 ;
        RECT 179.730 368.800 180.050 368.810 ;
        RECT 284.780 368.680 288.090 370.740 ;
        RECT 182.490 368.570 182.800 368.580 ;
        RECT 182.490 368.540 182.810 368.570 ;
        RECT 172.490 367.920 174.930 367.930 ;
        RECT 171.800 367.590 171.910 367.790 ;
        RECT 172.200 367.730 174.930 367.920 ;
        RECT 175.240 368.340 182.810 368.540 ;
        RECT 172.200 367.720 172.690 367.730 ;
        RECT 170.400 367.390 170.720 367.440 ;
        RECT 140.810 367.240 141.120 367.330 ;
        RECT 140.210 367.070 141.120 367.240 ;
        RECT 140.810 367.000 141.120 367.070 ;
        RECT 141.900 367.250 142.210 367.340 ;
        RECT 141.900 367.080 143.010 367.250 ;
        RECT 141.900 367.010 142.210 367.080 ;
        RECT 161.740 367.030 162.070 367.040 ;
        RECT 161.720 366.930 162.090 367.030 ;
        RECT 161.720 366.760 164.070 366.930 ;
        RECT 161.720 366.650 162.090 366.760 ;
        RECT 163.110 366.610 163.200 366.760 ;
        RECT 165.570 366.570 165.830 367.370 ;
        RECT 170.400 367.190 172.030 367.390 ;
        RECT 170.400 367.180 170.720 367.190 ;
        RECT 167.570 366.570 167.910 366.630 ;
        RECT 57.870 366.180 61.250 366.500 ;
        RECT 163.300 366.210 163.760 366.530 ;
        RECT 165.470 366.350 167.910 366.570 ;
        RECT 175.240 366.380 175.440 368.340 ;
        RECT 182.490 368.310 182.810 368.340 ;
        RECT 182.490 368.300 182.800 368.310 ;
        RECT 183.550 368.060 183.870 368.100 ;
        RECT 172.490 366.370 175.440 366.380 ;
        RECT 171.800 366.040 171.910 366.240 ;
        RECT 172.200 366.180 175.440 366.370 ;
        RECT 175.790 367.860 183.950 368.060 ;
        RECT 172.200 366.170 172.700 366.180 ;
        RECT 170.400 365.840 170.720 365.890 ;
        RECT 161.140 365.450 161.530 365.550 ;
        RECT 161.140 365.280 164.070 365.450 ;
        RECT 161.140 365.180 161.530 365.280 ;
        RECT 163.110 365.060 163.200 365.280 ;
        RECT 165.570 365.020 165.830 365.820 ;
        RECT 170.400 365.640 172.030 365.840 ;
        RECT 170.400 365.630 170.720 365.640 ;
        RECT 167.570 365.020 167.910 365.080 ;
        RECT 163.300 364.660 163.760 364.980 ;
        RECT 165.470 364.800 167.910 365.020 ;
        RECT 175.790 364.830 175.990 367.860 ;
        RECT 183.550 367.820 183.870 367.860 ;
        RECT 243.490 366.620 288.410 368.680 ;
        RECT 172.500 364.820 175.990 364.830 ;
        RECT 172.200 364.630 175.990 364.820 ;
        RECT 178.940 366.060 179.230 366.240 ;
        RECT 172.200 364.620 172.660 364.630 ;
        RECT 160.500 363.850 160.890 363.940 ;
        RECT 145.930 363.760 146.250 363.790 ;
        RECT 144.720 363.560 146.350 363.760 ;
        RECT 160.500 363.680 164.070 363.850 ;
        RECT 160.500 363.590 160.890 363.680 ;
        RECT 145.930 363.530 146.250 363.560 ;
        RECT 159.860 363.280 160.250 363.390 ;
        RECT 159.860 363.110 164.070 363.280 ;
        RECT 159.860 363.010 160.250 363.110 ;
        RECT 145.940 362.800 146.260 362.830 ;
        RECT 178.940 362.800 179.120 366.060 ;
        RECT 209.140 364.650 209.220 364.830 ;
        RECT 313.170 364.600 317.100 365.050 ;
        RECT 203.290 363.630 203.890 364.190 ;
        RECT 206.890 364.020 212.120 364.250 ;
        RECT 207.360 363.780 207.670 363.920 ;
        RECT 205.190 363.770 207.670 363.780 ;
        RECT 205.190 363.620 216.710 363.770 ;
        RECT 205.190 363.600 207.670 363.620 ;
        RECT 207.360 363.590 207.670 363.600 ;
        RECT 206.900 363.200 212.120 363.420 ;
        RECT 144.720 362.600 146.350 362.800 ;
        RECT 178.110 362.620 179.120 362.800 ;
        RECT 184.360 362.990 184.680 363.040 ;
        RECT 186.770 362.990 187.090 363.010 ;
        RECT 184.360 362.850 187.090 362.990 ;
        RECT 184.360 362.800 188.790 362.850 ;
        RECT 184.360 362.720 184.680 362.800 ;
        RECT 186.770 362.750 188.790 362.800 ;
        RECT 186.810 362.680 188.790 362.750 ;
        RECT 188.270 362.670 188.790 362.680 ;
        RECT 207.360 362.620 207.670 362.630 ;
        RECT 145.940 362.570 146.260 362.600 ;
        RECT 172.500 362.410 172.800 362.440 ;
        RECT 172.500 362.400 172.890 362.410 ;
        RECT 163.300 362.040 163.760 362.360 ;
        RECT 165.470 362.000 167.910 362.220 ;
        RECT 172.200 362.200 172.890 362.400 ;
        RECT 183.120 362.280 183.600 362.510 ;
        RECT 205.190 362.440 216.720 362.620 ;
        RECT 243.490 362.540 317.100 364.600 ;
        RECT 313.170 362.530 317.100 362.540 ;
        RECT 207.360 362.300 207.670 362.440 ;
        RECT 183.260 362.210 183.600 362.280 ;
        RECT 136.660 361.710 142.310 361.900 ;
        RECT 145.930 361.840 146.250 361.870 ;
        RECT 98.570 361.590 99.190 361.680 ;
        RECT 98.570 361.180 127.510 361.590 ;
        RECT 98.570 361.090 99.190 361.180 ;
        RECT 125.730 350.600 127.000 351.250 ;
        RECT 28.120 350.340 127.960 350.600 ;
        RECT 136.660 350.340 137.030 361.710 ;
        RECT 144.720 361.640 146.350 361.840 ;
        RECT 159.250 361.710 159.640 361.810 ;
        RECT 163.110 361.710 163.200 361.960 ;
        RECT 145.930 361.610 146.250 361.640 ;
        RECT 159.250 361.540 164.070 361.710 ;
        RECT 159.250 361.440 159.640 361.540 ;
        RECT 165.570 361.200 165.830 362.000 ;
        RECT 167.570 361.940 167.910 362.000 ;
        RECT 207.210 361.600 207.520 361.670 ;
        RECT 205.190 361.590 207.520 361.600 ;
        RECT 170.400 361.380 170.720 361.390 ;
        RECT 170.400 361.180 172.030 361.380 ;
        RECT 170.400 361.130 170.720 361.180 ;
        RECT 172.470 361.090 172.800 361.290 ;
        RECT 178.500 361.170 179.230 361.350 ;
        RECT 183.260 361.340 183.600 361.410 ;
        RECT 205.190 361.380 216.720 361.590 ;
        RECT 206.500 361.370 216.720 361.380 ;
        RECT 207.210 361.340 207.520 361.370 ;
        RECT 163.300 360.490 163.760 360.810 ;
        RECT 171.800 360.780 171.910 360.980 ;
        RECT 172.470 360.870 172.650 361.090 ;
        RECT 178.500 360.960 178.680 361.170 ;
        RECT 183.120 361.110 183.600 361.340 ;
        RECT 172.450 360.850 172.650 360.870 ;
        RECT 165.470 360.450 167.910 360.670 ;
        RECT 172.200 360.650 172.650 360.850 ;
        RECT 178.110 360.780 178.680 360.960 ;
        RECT 207.670 360.740 212.120 360.900 ;
        RECT 207.640 360.700 212.120 360.740 ;
        RECT 158.620 360.180 159.040 360.270 ;
        RECT 163.110 360.180 163.200 360.410 ;
        RECT 158.620 360.010 164.070 360.180 ;
        RECT 158.620 359.920 159.040 360.010 ;
        RECT 165.570 359.650 165.830 360.450 ;
        RECT 167.570 360.390 167.910 360.450 ;
        RECT 178.600 360.020 179.150 360.200 ;
        RECT 202.230 360.160 202.790 360.700 ;
        RECT 207.640 360.620 207.870 360.700 ;
        RECT 206.260 360.400 216.720 360.620 ;
        RECT 206.260 360.260 206.580 360.400 ;
        RECT 184.360 360.060 184.680 360.110 ;
        RECT 186.770 360.060 187.090 360.080 ;
        RECT 170.400 359.830 170.720 359.840 ;
        RECT 170.400 359.630 172.030 359.830 ;
        RECT 178.600 359.810 178.780 360.020 ;
        RECT 178.110 359.630 178.780 359.810 ;
        RECT 184.360 359.870 187.090 360.060 ;
        RECT 206.280 359.920 206.540 360.260 ;
        RECT 184.360 359.790 184.680 359.870 ;
        RECT 186.770 359.860 187.090 359.870 ;
        RECT 186.770 359.820 188.790 359.860 ;
        RECT 186.880 359.700 188.790 359.820 ;
        RECT 187.600 359.680 188.790 359.700 ;
        RECT 206.260 359.660 206.580 359.920 ;
        RECT 170.400 359.580 170.720 359.630 ;
        RECT 172.450 359.460 172.800 359.530 ;
        RECT 163.300 358.940 163.760 359.260 ;
        RECT 171.800 359.230 171.910 359.430 ;
        RECT 172.450 359.300 172.840 359.460 ;
        RECT 183.120 359.350 183.600 359.580 ;
        RECT 172.260 359.230 172.840 359.300 ;
        RECT 183.260 359.280 183.600 359.350 ;
        RECT 165.470 358.900 167.910 359.120 ;
        RECT 172.260 359.100 172.650 359.230 ;
        RECT 158.060 358.610 158.450 358.700 ;
        RECT 163.110 358.610 163.200 358.860 ;
        RECT 158.060 358.440 164.070 358.610 ;
        RECT 158.060 358.350 158.450 358.440 ;
        RECT 165.570 358.100 165.830 358.900 ;
        RECT 167.570 358.840 167.910 358.900 ;
        RECT 207.210 358.840 207.520 358.910 ;
        RECT 207.640 358.840 207.870 360.400 ;
        RECT 341.970 360.260 345.470 360.800 ;
        RECT 209.140 359.780 209.220 359.960 ;
        RECT 205.190 358.630 216.720 358.840 ;
        RECT 206.500 358.620 216.720 358.630 ;
        RECT 207.210 358.580 207.520 358.620 ;
        RECT 183.260 358.410 183.600 358.480 ;
        RECT 170.400 358.280 170.720 358.290 ;
        RECT 170.400 358.080 172.030 358.280 ;
        RECT 172.540 358.150 172.800 358.360 ;
        RECT 183.120 358.180 183.600 358.410 ;
        RECT 207.640 358.220 207.870 358.620 ;
        RECT 170.400 358.030 170.720 358.080 ;
        RECT 163.300 357.390 163.760 357.710 ;
        RECT 171.800 357.680 171.910 357.880 ;
        RECT 172.540 357.750 172.740 358.150 ;
        RECT 187.540 357.990 188.790 358.000 ;
        RECT 178.110 357.770 178.880 357.950 ;
        RECT 165.470 357.350 167.910 357.570 ;
        RECT 172.400 357.550 172.740 357.750 ;
        RECT 172.540 357.540 172.740 357.550 ;
        RECT 163.110 356.990 163.200 357.310 ;
        RECT 165.570 356.550 165.830 357.350 ;
        RECT 167.570 357.290 167.910 357.350 ;
        RECT 170.400 356.730 170.720 356.740 ;
        RECT 170.400 356.530 172.030 356.730 ;
        RECT 170.400 356.480 170.720 356.530 ;
        RECT 171.800 356.130 171.910 356.330 ;
        RECT 178.700 355.330 178.880 357.770 ;
        RECT 184.360 357.890 184.680 357.970 ;
        RECT 186.850 357.940 188.790 357.990 ;
        RECT 186.770 357.890 188.790 357.940 ;
        RECT 184.360 357.830 188.790 357.890 ;
        RECT 184.360 357.700 187.090 357.830 ;
        RECT 187.540 357.820 188.790 357.830 ;
        RECT 184.360 357.650 184.680 357.700 ;
        RECT 186.770 357.680 187.090 357.700 ;
        RECT 203.270 357.610 203.890 358.140 ;
        RECT 206.890 357.990 207.870 358.220 ;
        RECT 208.480 358.090 212.120 358.290 ;
        RECT 243.490 358.210 345.560 360.260 ;
        RECT 207.360 357.750 207.670 357.890 ;
        RECT 205.190 357.740 207.670 357.750 ;
        RECT 208.480 357.740 208.680 358.090 ;
        RECT 205.190 357.590 216.720 357.740 ;
        RECT 205.190 357.570 207.670 357.590 ;
        RECT 207.360 357.560 207.670 357.570 ;
        RECT 208.480 357.390 208.680 357.590 ;
        RECT 206.900 357.240 208.680 357.390 ;
        RECT 206.900 357.170 208.650 357.240 ;
        RECT 192.670 356.710 192.980 356.850 ;
        RECT 213.440 356.710 213.750 356.850 ;
        RECT 234.320 356.820 234.630 356.870 ;
        RECT 236.620 356.820 236.930 356.840 ;
        RECT 190.510 356.530 200.580 356.710 ;
        RECT 205.840 356.530 215.910 356.710 ;
        RECT 218.450 356.580 227.460 356.800 ;
        RECT 233.110 356.600 233.420 356.640 ;
        RECT 192.670 356.520 192.980 356.530 ;
        RECT 213.440 356.520 213.750 356.530 ;
        RECT 192.670 356.280 192.980 356.300 ;
        RECT 213.440 356.280 213.750 356.300 ;
        RECT 190.510 356.100 200.580 356.280 ;
        RECT 205.840 356.100 215.910 356.280 ;
        RECT 192.670 355.970 192.980 356.100 ;
        RECT 213.440 355.970 213.750 356.100 ;
        RECT 178.700 355.150 179.240 355.330 ;
        RECT 192.670 355.280 192.980 355.410 ;
        RECT 213.440 355.280 213.750 355.410 ;
        RECT 190.510 355.100 200.590 355.280 ;
        RECT 205.830 355.100 215.910 355.280 ;
        RECT 192.670 355.080 192.980 355.100 ;
        RECT 213.440 355.080 213.750 355.100 ;
        RECT 192.670 354.850 192.980 354.860 ;
        RECT 213.440 354.850 213.750 354.860 ;
        RECT 190.510 354.670 200.590 354.850 ;
        RECT 205.830 354.670 215.910 354.850 ;
        RECT 218.500 354.800 224.160 355.020 ;
        RECT 192.670 354.530 192.980 354.670 ;
        RECT 213.440 354.530 213.750 354.670 ;
        RECT 218.000 354.500 218.480 354.510 ;
        RECT 218.000 354.260 218.890 354.500 ;
        RECT 223.940 354.470 224.160 354.800 ;
        RECT 227.240 354.970 227.460 356.580 ;
        RECT 232.790 356.590 233.450 356.600 ;
        RECT 234.320 356.590 237.240 356.820 ;
        RECT 232.790 356.360 233.890 356.590 ;
        RECT 234.320 356.540 234.630 356.590 ;
        RECT 236.620 356.510 236.930 356.590 ;
        RECT 233.110 356.310 233.420 356.360 ;
        RECT 353.670 356.190 359.380 361.830 ;
        RECT 353.230 356.150 359.380 356.190 ;
        RECT 234.320 355.990 234.630 356.050 ;
        RECT 236.610 355.990 236.920 356.120 ;
        RECT 234.320 355.770 237.240 355.990 ;
        RECT 234.320 355.720 234.630 355.770 ;
        RECT 243.490 355.690 359.380 356.150 ;
        RECT 227.240 354.750 230.090 354.970 ;
        RECT 234.270 354.520 234.580 354.560 ;
        RECT 228.310 354.470 234.580 354.520 ;
        RECT 223.940 354.310 234.580 354.470 ;
        RECT 223.940 354.250 228.700 354.310 ;
        RECT 234.270 354.230 234.580 354.310 ;
        RECT 192.670 353.700 192.980 353.840 ;
        RECT 209.150 353.790 209.230 353.930 ;
        RECT 210.440 353.790 210.870 353.870 ;
        RECT 190.510 353.690 192.980 353.700 ;
        RECT 199.180 353.690 210.870 353.790 ;
        RECT 213.440 353.700 213.750 353.840 ;
        RECT 234.320 353.830 234.630 353.910 ;
        RECT 236.530 353.830 236.840 353.870 ;
        RECT 213.440 353.690 215.910 353.700 ;
        RECT 190.510 353.530 215.910 353.690 ;
        RECT 234.320 353.600 237.030 353.830 ;
        RECT 243.490 353.790 359.220 355.690 ;
        RECT 234.320 353.580 234.630 353.600 ;
        RECT 236.530 353.540 236.840 353.600 ;
        RECT 190.510 353.520 200.570 353.530 ;
        RECT 205.850 353.520 215.910 353.530 ;
        RECT 192.670 353.510 192.980 353.520 ;
        RECT 210.440 353.460 210.870 353.520 ;
        RECT 213.440 353.510 213.750 353.520 ;
        RECT 157.450 353.140 157.820 353.260 ;
        RECT 157.450 352.970 163.770 353.140 ;
        RECT 157.450 352.860 157.820 352.970 ;
        RECT 184.360 352.920 184.680 352.970 ;
        RECT 186.770 352.920 187.090 352.940 ;
        RECT 178.870 352.730 180.650 352.850 ;
        RECT 178.280 352.670 180.650 352.730 ;
        RECT 184.360 352.780 187.090 352.920 ;
        RECT 184.360 352.730 188.790 352.780 ;
        RECT 178.280 352.550 179.120 352.670 ;
        RECT 184.360 352.650 184.680 352.730 ;
        RECT 186.770 352.680 188.790 352.730 ;
        RECT 193.150 352.710 193.290 352.900 ;
        RECT 213.180 352.710 213.270 352.890 ;
        RECT 186.810 352.610 188.790 352.680 ;
        RECT 188.270 352.600 188.790 352.610 ;
        RECT 172.540 352.370 172.790 352.390 ;
        RECT 172.540 352.270 172.800 352.370 ;
        RECT 163.300 351.910 163.760 352.230 ;
        RECT 165.470 351.870 167.910 352.090 ;
        RECT 172.200 352.070 172.800 352.270 ;
        RECT 183.120 352.210 183.600 352.440 ;
        RECT 192.670 352.290 192.980 352.410 ;
        RECT 193.150 352.290 193.290 352.470 ;
        RECT 200.410 352.290 200.970 352.420 ;
        RECT 213.180 352.290 213.270 352.460 ;
        RECT 213.440 352.290 213.750 352.410 ;
        RECT 192.670 352.280 200.970 352.290 ;
        RECT 183.260 352.140 183.600 352.210 ;
        RECT 190.510 352.240 200.970 352.280 ;
        RECT 205.850 352.280 213.750 352.290 ;
        RECT 190.510 352.120 200.570 352.240 ;
        RECT 205.850 352.120 215.910 352.280 ;
        RECT 190.510 352.100 193.070 352.120 ;
        RECT 192.670 352.080 192.980 352.100 ;
        RECT 198.250 352.030 199.790 352.120 ;
        RECT 206.630 352.030 208.170 352.120 ;
        RECT 213.350 352.100 215.910 352.120 ;
        RECT 213.440 352.080 213.750 352.100 ;
        RECT 156.810 351.550 157.200 351.640 ;
        RECT 163.110 351.550 163.200 351.830 ;
        RECT 156.810 351.380 163.770 351.550 ;
        RECT 156.810 351.290 157.200 351.380 ;
        RECT 165.570 351.070 165.830 351.870 ;
        RECT 167.570 351.810 167.910 351.870 ;
        RECT 192.670 351.850 192.980 351.860 ;
        RECT 213.440 351.850 213.750 351.860 ;
        RECT 190.510 351.680 200.570 351.850 ;
        RECT 205.850 351.680 215.910 351.850 ;
        RECT 190.510 351.670 192.980 351.680 ;
        RECT 192.670 351.530 192.980 351.670 ;
        RECT 213.440 351.670 215.910 351.680 ;
        RECT 183.260 351.270 183.600 351.340 ;
        RECT 193.150 351.280 193.300 351.470 ;
        RECT 211.180 351.420 211.620 351.540 ;
        RECT 213.440 351.530 213.750 351.670 ;
        RECT 170.400 351.250 170.720 351.260 ;
        RECT 170.400 351.050 172.030 351.250 ;
        RECT 170.400 351.000 170.720 351.050 ;
        RECT 172.390 351.020 172.770 351.220 ;
        RECT 183.120 351.040 183.600 351.270 ;
        RECT 200.420 351.240 211.620 351.420 ;
        RECT 213.150 351.280 213.280 351.460 ;
        RECT 347.890 351.410 349.980 351.590 ;
        RECT 211.180 351.140 211.620 351.240 ;
        RECT 172.390 350.990 172.760 351.020 ;
        RECT 163.300 350.360 163.760 350.680 ;
        RECT 171.800 350.650 171.910 350.850 ;
        RECT 172.390 350.720 172.590 350.990 ;
        RECT 178.890 350.890 180.650 350.990 ;
        RECT 28.120 349.970 137.030 350.340 ;
        RECT 165.470 350.320 167.910 350.540 ;
        RECT 172.200 350.520 172.590 350.720 ;
        RECT 178.290 350.810 180.650 350.890 ;
        RECT 178.290 350.710 179.170 350.810 ;
        RECT 184.360 350.750 184.680 350.830 ;
        RECT 186.840 350.800 188.790 350.940 ;
        RECT 193.150 350.850 193.280 351.030 ;
        RECT 213.140 350.850 213.280 351.030 ;
        RECT 186.770 350.780 188.790 350.800 ;
        RECT 186.770 350.750 187.090 350.780 ;
        RECT 187.570 350.770 188.790 350.780 ;
        RECT 188.270 350.760 188.790 350.770 ;
        RECT 184.360 350.560 187.090 350.750 ;
        RECT 184.360 350.510 184.680 350.560 ;
        RECT 186.770 350.540 187.090 350.560 ;
        RECT 156.190 350.000 156.580 350.080 ;
        RECT 163.110 350.000 163.200 350.280 ;
        RECT 28.120 348.520 127.960 349.970 ;
        RECT 156.190 349.830 163.770 350.000 ;
        RECT 156.190 349.750 156.580 349.830 ;
        RECT 165.570 349.520 165.830 350.320 ;
        RECT 167.570 350.260 167.910 350.320 ;
        RECT 184.360 349.990 184.680 350.040 ;
        RECT 186.770 349.990 187.090 350.010 ;
        RECT 178.900 349.740 180.650 349.840 ;
        RECT 170.400 349.700 170.720 349.710 ;
        RECT 170.400 349.500 172.030 349.700 ;
        RECT 178.290 349.660 180.650 349.740 ;
        RECT 184.360 349.800 187.090 349.990 ;
        RECT 184.360 349.720 184.680 349.800 ;
        RECT 186.770 349.790 187.090 349.800 ;
        RECT 186.770 349.750 188.790 349.790 ;
        RECT 178.290 349.560 179.170 349.660 ;
        RECT 186.880 349.630 188.790 349.750 ;
        RECT 193.150 349.700 193.220 349.880 ;
        RECT 213.190 349.700 213.280 349.880 ;
        RECT 187.600 349.610 188.790 349.630 ;
        RECT 170.400 349.450 170.720 349.500 ;
        RECT 163.300 348.810 163.760 349.130 ;
        RECT 171.800 349.100 171.910 349.300 ;
        RECT 172.600 349.170 172.800 349.450 ;
        RECT 183.120 349.280 183.600 349.510 ;
        RECT 183.260 349.210 183.600 349.280 ;
        RECT 193.150 349.270 193.220 349.450 ;
        RECT 213.190 349.270 213.280 349.450 ;
        RECT 243.490 349.320 349.980 351.410 ;
        RECT 165.470 348.770 167.910 348.990 ;
        RECT 172.200 348.970 172.800 349.170 ;
        RECT 155.580 348.520 156.000 348.610 ;
        RECT 163.110 348.520 163.200 348.730 ;
        RECT 28.120 304.690 30.200 348.520 ;
        RECT 155.580 348.350 163.770 348.520 ;
        RECT 155.580 348.250 156.000 348.350 ;
        RECT 165.570 347.970 165.830 348.770 ;
        RECT 167.570 348.710 167.910 348.770 ;
        RECT 199.850 348.720 206.610 348.900 ;
        RECT 183.260 348.340 183.600 348.410 ;
        RECT 170.400 348.150 170.720 348.160 ;
        RECT 170.400 347.950 172.030 348.150 ;
        RECT 170.400 347.900 170.720 347.950 ;
        RECT 163.300 347.260 163.760 347.580 ;
        RECT 171.800 347.550 171.910 347.750 ;
        RECT 172.600 347.620 172.800 348.290 ;
        RECT 183.120 348.110 183.600 348.340 ;
        RECT 193.150 348.280 193.220 348.460 ;
        RECT 213.190 348.280 213.280 348.460 ;
        RECT 178.870 347.880 180.650 347.990 ;
        RECT 187.540 347.920 188.790 347.930 ;
        RECT 178.290 347.810 180.650 347.880 ;
        RECT 184.360 347.820 184.680 347.900 ;
        RECT 186.850 347.870 188.790 347.920 ;
        RECT 186.770 347.820 188.790 347.870 ;
        RECT 193.150 347.850 193.220 348.030 ;
        RECT 213.190 347.850 213.280 348.030 ;
        RECT 178.290 347.700 179.170 347.810 ;
        RECT 184.360 347.760 188.790 347.820 ;
        RECT 165.470 347.220 167.910 347.440 ;
        RECT 172.200 347.420 172.800 347.620 ;
        RECT 184.360 347.630 187.090 347.760 ;
        RECT 187.540 347.750 188.790 347.760 ;
        RECT 184.360 347.580 184.680 347.630 ;
        RECT 186.770 347.610 187.090 347.630 ;
        RECT 125.670 346.190 126.940 347.030 ;
        RECT 163.110 346.860 163.200 347.180 ;
        RECT 165.570 346.420 165.830 347.220 ;
        RECT 167.570 347.160 167.910 347.220 ;
        RECT 170.400 346.600 170.720 346.610 ;
        RECT 170.400 346.400 172.030 346.600 ;
        RECT 170.400 346.350 170.720 346.400 ;
        RECT 125.670 345.820 135.370 346.190 ;
        RECT 171.800 346.000 171.910 346.200 ;
        RECT 125.670 345.780 126.940 345.820 ;
        RECT 27.900 301.280 30.200 304.690 ;
        RECT 28.120 300.950 30.200 301.280 ;
        RECT 32.460 343.700 127.960 345.780 ;
        RECT 135.000 344.470 135.370 345.820 ;
        RECT 135.000 344.460 137.030 344.470 ;
        RECT 135.000 344.280 137.250 344.460 ;
        RECT 193.250 344.310 193.560 344.450 ;
        RECT 191.080 344.300 193.560 344.310 ;
        RECT 135.000 344.220 138.650 344.280 ;
        RECT 141.650 344.220 141.960 344.260 ;
        RECT 135.000 344.100 141.960 344.220 ;
        RECT 191.080 344.130 193.680 344.300 ;
        RECT 193.250 344.120 193.560 344.130 ;
        RECT 136.660 344.060 141.960 344.100 ;
        RECT 137.030 344.000 141.960 344.060 ;
        RECT 129.660 343.810 130.430 344.000 ;
        RECT 141.650 343.930 141.960 344.000 ;
        RECT 243.490 343.920 345.840 346.010 ;
        RECT 136.660 343.810 137.050 343.830 ;
        RECT 129.660 343.770 137.050 343.810 ;
        RECT 140.430 343.770 140.740 343.820 ;
        RECT 32.460 276.210 34.540 343.700 ;
        RECT 129.660 343.560 140.740 343.770 ;
        RECT 129.660 343.440 137.040 343.560 ;
        RECT 140.430 343.490 140.740 343.560 ;
        RECT 129.660 343.260 130.430 343.440 ;
        RECT 136.660 343.420 137.030 343.440 ;
        RECT 154.940 343.350 155.350 343.450 ;
        RECT 154.940 343.180 163.770 343.350 ;
        RECT 193.200 343.320 193.750 343.500 ;
        RECT 194.280 343.290 194.600 343.350 ;
        RECT 198.300 343.290 198.630 343.320 ;
        RECT 154.940 343.090 155.350 343.180 ;
        RECT 184.360 343.160 184.680 343.210 ;
        RECT 186.770 343.160 187.090 343.180 ;
        RECT 125.730 342.160 127.000 342.930 ;
        RECT 178.140 342.890 180.100 343.070 ;
        RECT 184.360 343.020 187.090 343.160 ;
        RECT 194.280 343.120 198.630 343.290 ;
        RECT 194.280 343.070 194.600 343.120 ;
        RECT 198.300 343.060 198.630 343.120 ;
        RECT 184.360 342.970 188.790 343.020 ;
        RECT 184.360 342.890 184.680 342.970 ;
        RECT 186.770 342.920 188.790 342.970 ;
        RECT 203.820 342.950 203.860 343.040 ;
        RECT 186.810 342.850 188.790 342.920 ;
        RECT 188.270 342.840 188.790 342.850 ;
        RECT 203.710 342.860 204.920 342.950 ;
        RECT 203.710 342.800 205.050 342.860 ;
        RECT 203.710 342.750 207.320 342.800 ;
        RECT 125.730 341.790 131.720 342.160 ;
        RECT 163.300 342.140 163.760 342.460 ;
        RECT 165.470 342.100 167.910 342.320 ;
        RECT 172.180 342.300 172.830 342.500 ;
        RECT 178.940 342.480 180.110 342.630 ;
        RECT 178.880 342.150 179.160 342.480 ;
        RECT 183.120 342.450 183.600 342.680 ;
        RECT 204.740 342.640 207.320 342.750 ;
        RECT 204.740 342.530 205.050 342.640 ;
        RECT 183.260 342.380 183.600 342.450 ;
        RECT 125.730 341.080 127.000 341.790 ;
        RECT 37.000 339.000 127.960 341.080 ;
        RECT 131.350 340.130 131.720 341.790 ;
        RECT 154.280 341.780 154.670 341.890 ;
        RECT 163.110 341.780 163.200 342.060 ;
        RECT 154.280 341.610 163.770 341.780 ;
        RECT 154.280 341.510 154.670 341.610 ;
        RECT 165.570 341.300 165.830 342.100 ;
        RECT 167.570 342.040 167.910 342.100 ;
        RECT 203.810 341.980 205.020 342.090 ;
        RECT 203.810 341.890 205.050 341.980 ;
        RECT 204.740 341.870 205.050 341.890 ;
        RECT 204.740 341.710 207.320 341.870 ;
        RECT 204.740 341.650 205.050 341.710 ;
        RECT 183.260 341.510 183.600 341.580 ;
        RECT 170.400 341.480 170.720 341.490 ;
        RECT 170.400 341.280 172.030 341.480 ;
        RECT 170.400 341.230 170.720 341.280 ;
        RECT 172.560 341.250 172.810 341.480 ;
        RECT 183.120 341.280 183.600 341.510 ;
        RECT 193.180 341.460 193.750 341.640 ;
        RECT 163.300 340.590 163.760 340.910 ;
        RECT 171.800 340.880 171.910 341.080 ;
        RECT 172.560 340.950 172.760 341.250 ;
        RECT 165.470 340.550 167.910 340.770 ;
        RECT 172.200 340.750 172.760 340.950 ;
        RECT 178.140 341.030 180.480 341.210 ;
        RECT 178.140 340.930 178.320 341.030 ;
        RECT 184.360 340.990 184.680 341.070 ;
        RECT 186.840 341.040 188.790 341.180 ;
        RECT 186.770 341.020 188.790 341.040 ;
        RECT 186.770 340.990 187.090 341.020 ;
        RECT 187.570 341.010 188.790 341.020 ;
        RECT 188.270 341.000 188.790 341.010 ;
        RECT 184.360 340.800 187.090 340.990 ;
        RECT 184.360 340.750 184.680 340.800 ;
        RECT 186.770 340.780 187.090 340.800 ;
        RECT 153.670 340.240 154.040 340.250 ;
        RECT 163.110 340.240 163.200 340.510 ;
        RECT 131.350 339.950 137.300 340.130 ;
        RECT 153.670 340.070 163.770 340.240 ;
        RECT 131.350 339.880 137.370 339.950 ;
        RECT 138.760 339.880 140.030 339.890 ;
        RECT 140.460 339.880 140.770 339.940 ;
        RECT 131.350 339.760 140.770 339.880 ;
        RECT 136.660 339.720 140.770 339.760 ;
        RECT 137.020 339.670 140.770 339.720 ;
        RECT 140.460 339.610 140.770 339.670 ;
        RECT 141.150 339.860 141.460 339.930 ;
        RECT 145.940 339.880 146.230 339.900 ;
        RECT 141.150 339.850 143.290 339.860 ;
        RECT 145.930 339.850 146.250 339.880 ;
        RECT 153.670 339.860 154.040 340.070 ;
        RECT 141.150 339.650 146.250 339.850 ;
        RECT 165.570 339.750 165.830 340.550 ;
        RECT 167.570 340.490 167.910 340.550 ;
        RECT 193.200 340.310 193.750 340.490 ;
        RECT 193.200 340.300 193.360 340.310 ;
        RECT 184.360 340.230 184.680 340.280 ;
        RECT 186.770 340.230 187.090 340.250 ;
        RECT 170.400 339.930 170.720 339.940 ;
        RECT 170.400 339.730 172.030 339.930 ;
        RECT 178.150 339.880 180.110 340.060 ;
        RECT 184.360 340.040 187.090 340.230 ;
        RECT 204.740 340.060 205.050 340.090 ;
        RECT 184.360 339.960 184.680 340.040 ;
        RECT 186.770 340.030 187.090 340.040 ;
        RECT 203.800 340.030 205.050 340.060 ;
        RECT 186.770 339.990 188.790 340.030 ;
        RECT 186.880 339.870 188.790 339.990 ;
        RECT 203.800 339.900 207.320 340.030 ;
        RECT 187.600 339.850 188.790 339.870 ;
        RECT 204.740 339.870 207.320 339.900 ;
        RECT 204.740 339.760 205.050 339.870 ;
        RECT 170.400 339.680 170.720 339.730 ;
        RECT 172.570 339.690 172.770 339.700 ;
        RECT 141.150 339.600 141.460 339.650 ;
        RECT 143.080 339.640 146.250 339.650 ;
        RECT 134.890 339.150 135.300 339.170 ;
        RECT 136.660 339.150 138.650 339.170 ;
        RECT 134.890 339.110 138.650 339.150 ;
        RECT 141.630 339.110 141.940 339.160 ;
        RECT 32.250 272.610 34.820 276.210 ;
        RECT 32.460 272.570 34.540 272.610 ;
        RECT 37.000 247.590 39.080 339.000 ;
        RECT 134.890 338.890 141.940 339.110 ;
        RECT 125.730 338.020 127.000 338.840 ;
        RECT 134.890 338.780 137.040 338.890 ;
        RECT 141.630 338.830 141.940 338.890 ;
        RECT 142.340 339.030 142.650 339.100 ;
        RECT 143.080 339.030 143.290 339.640 ;
        RECT 145.930 339.620 146.250 339.640 ;
        RECT 145.940 339.600 146.230 339.620 ;
        RECT 163.300 339.040 163.760 339.360 ;
        RECT 171.800 339.330 171.910 339.530 ;
        RECT 172.570 339.420 172.860 339.690 ;
        RECT 179.490 339.630 179.810 339.680 ;
        RECT 179.490 339.430 180.100 339.630 ;
        RECT 183.120 339.520 183.600 339.750 ;
        RECT 206.870 339.540 207.200 339.630 ;
        RECT 183.260 339.450 183.600 339.520 ;
        RECT 172.570 339.400 172.770 339.420 ;
        RECT 142.340 338.820 143.290 339.030 ;
        RECT 165.470 339.000 167.910 339.220 ;
        RECT 172.160 339.200 172.770 339.400 ;
        RECT 179.490 339.360 179.950 339.430 ;
        RECT 200.520 339.370 207.200 339.540 ;
        RECT 206.870 339.340 207.200 339.370 ;
        RECT 134.890 338.760 135.300 338.780 ;
        RECT 136.660 338.760 137.030 338.780 ;
        RECT 142.340 338.770 142.650 338.820 ;
        RECT 152.980 338.700 153.370 338.800 ;
        RECT 163.110 338.700 163.200 338.960 ;
        RECT 152.980 338.530 163.770 338.700 ;
        RECT 152.980 338.430 153.370 338.530 ;
        RECT 129.660 338.020 130.460 338.160 ;
        RECT 125.730 337.520 130.460 338.020 ;
        RECT 142.300 337.950 142.910 338.280 ;
        RECT 165.570 338.200 165.830 339.000 ;
        RECT 167.570 338.940 167.910 339.000 ;
        RECT 193.150 338.820 193.460 339.150 ;
        RECT 204.740 339.100 205.050 339.210 ;
        RECT 204.740 339.090 207.320 339.100 ;
        RECT 203.810 338.940 207.320 339.090 ;
        RECT 243.490 339.040 341.760 341.130 ;
        RECT 203.810 338.910 205.050 338.940 ;
        RECT 204.740 338.880 205.050 338.910 ;
        RECT 197.250 338.670 197.570 338.720 ;
        RECT 183.260 338.580 183.600 338.650 ;
        RECT 172.550 338.540 172.850 338.580 ;
        RECT 170.400 338.380 170.720 338.390 ;
        RECT 170.400 338.180 172.030 338.380 ;
        RECT 172.540 338.300 172.850 338.540 ;
        RECT 183.120 338.350 183.600 338.580 ;
        RECT 192.730 338.510 197.570 338.670 ;
        RECT 193.220 338.460 193.750 338.510 ;
        RECT 197.250 338.460 197.570 338.510 ;
        RECT 204.590 338.470 204.900 338.530 ;
        RECT 204.040 338.460 204.900 338.470 ;
        RECT 170.400 338.130 170.720 338.180 ;
        RECT 125.730 336.960 127.000 337.520 ;
        RECT 129.660 337.390 130.460 337.520 ;
        RECT 142.310 337.460 142.910 337.950 ;
        RECT 163.300 337.490 163.760 337.810 ;
        RECT 171.800 337.780 171.910 337.980 ;
        RECT 172.540 337.850 172.740 338.300 ;
        RECT 178.150 338.030 180.440 338.210 ;
        RECT 193.200 338.180 193.510 338.300 ;
        RECT 196.460 338.240 204.900 338.460 ;
        RECT 196.460 338.230 204.050 338.240 ;
        RECT 196.460 338.220 197.230 338.230 ;
        RECT 196.460 338.180 196.700 338.220 ;
        RECT 204.590 338.200 204.900 338.240 ;
        RECT 187.540 338.160 188.790 338.170 ;
        RECT 184.360 338.060 184.680 338.140 ;
        RECT 186.850 338.110 188.790 338.160 ;
        RECT 186.770 338.060 188.790 338.110 ;
        RECT 172.190 337.650 172.740 337.850 ;
        RECT 184.360 338.000 188.790 338.060 ;
        RECT 184.360 337.870 187.090 338.000 ;
        RECT 187.540 337.990 188.790 338.000 ;
        RECT 193.200 337.980 196.700 338.180 ;
        RECT 193.200 337.970 195.890 337.980 ;
        RECT 184.360 337.820 184.680 337.870 ;
        RECT 186.770 337.850 187.090 337.870 ;
        RECT 163.110 337.090 163.200 337.410 ;
        RECT 172.280 337.260 172.600 337.310 ;
        RECT 178.890 337.260 179.210 337.360 ;
        RECT 172.280 337.100 179.210 337.260 ;
        RECT 172.280 337.050 172.600 337.100 ;
        RECT 178.890 337.080 179.210 337.100 ;
        RECT 179.920 337.260 180.240 337.350 ;
        RECT 190.540 337.260 190.950 337.370 ;
        RECT 179.920 337.100 190.950 337.260 ;
        RECT 179.920 337.070 180.240 337.100 ;
        RECT 179.480 337.020 179.760 337.030 ;
        RECT 179.460 336.930 179.780 337.020 ;
        RECT 190.540 337.000 190.950 337.100 ;
        RECT 181.700 336.930 182.020 336.960 ;
        RECT 179.430 336.770 182.020 336.930 ;
        RECT 179.460 336.760 179.780 336.770 ;
        RECT 179.480 336.750 179.760 336.760 ;
        RECT 181.700 336.700 182.020 336.770 ;
        RECT 181.720 336.690 182.000 336.700 ;
        RECT 180.500 335.420 180.880 335.810 ;
        RECT 196.580 335.800 196.880 335.820 ;
        RECT 181.650 335.380 182.050 335.720 ;
        RECT 190.240 335.220 190.900 335.580 ;
        RECT 195.870 335.460 196.890 335.800 ;
        RECT 196.580 335.440 196.890 335.460 ;
        RECT 171.800 334.380 172.180 334.760 ;
        RECT 191.990 334.500 192.440 334.930 ;
        RECT 243.490 333.840 337.670 335.930 ;
        RECT 125.670 332.910 126.940 333.690 ;
        RECT 134.900 332.910 135.310 332.930 ;
        RECT 125.670 332.750 135.310 332.910 ;
        RECT 45.690 332.540 135.310 332.750 ;
        RECT 45.690 330.670 127.960 332.540 ;
        RECT 134.900 332.520 135.310 332.540 ;
        RECT 240.740 330.720 240.750 330.730 ;
        RECT 36.840 244.020 39.230 247.590 ;
        RECT 37.000 243.490 39.080 244.020 ;
        RECT 45.690 190.470 47.770 330.670 ;
        RECT 141.590 330.390 142.200 330.720 ;
        RECT 141.600 329.900 142.200 330.390 ;
        RECT 197.230 330.540 243.020 330.550 ;
        RECT 197.230 330.050 243.230 330.540 ;
        RECT 171.820 326.320 172.420 326.810 ;
        RECT 180.280 326.320 180.880 326.810 ;
        RECT 171.820 325.990 172.430 326.320 ;
        RECT 180.270 325.990 180.880 326.320 ;
        RECT 98.670 325.590 99.270 325.640 ;
        RECT 98.670 325.150 128.010 325.590 ;
        RECT 98.670 325.080 99.270 325.150 ;
        RECT 227.630 323.420 227.920 323.480 ;
        RECT 227.460 323.110 227.920 323.420 ;
        RECT 227.630 323.070 227.920 323.110 ;
        RECT 227.640 322.750 227.920 323.070 ;
        RECT 227.460 322.440 227.920 322.750 ;
        RECT 227.640 322.320 227.920 322.440 ;
        RECT 145.870 321.270 146.180 321.290 ;
        RECT 141.640 320.930 146.180 321.270 ;
        RECT 145.870 320.910 146.180 320.930 ;
        RECT 162.320 319.690 162.740 319.700 ;
        RECT 162.320 319.440 202.590 319.690 ;
        RECT 162.320 319.360 202.600 319.440 ;
        RECT 162.320 319.350 162.740 319.360 ;
        RECT 196.560 319.340 202.600 319.360 ;
        RECT 58.360 317.110 127.960 319.190 ;
        RECT 161.720 319.070 162.100 319.080 ;
        RECT 161.720 318.740 198.520 319.070 ;
        RECT 161.720 318.730 162.100 318.740 ;
        RECT 192.450 318.730 198.520 318.740 ;
        RECT 161.080 318.440 161.500 318.450 ;
        RECT 161.080 318.110 194.440 318.440 ;
        RECT 161.080 318.100 161.500 318.110 ;
        RECT 160.490 317.800 160.890 317.820 ;
        RECT 160.490 317.470 190.430 317.800 ;
        RECT 160.490 317.460 160.890 317.470 ;
        RECT 159.830 317.130 160.240 317.140 ;
        RECT 45.440 186.740 48.040 190.470 ;
        RECT 45.690 186.410 47.770 186.740 ;
        RECT 58.360 104.930 60.440 317.110 ;
        RECT 125.600 316.960 126.870 317.110 ;
        RECT 159.820 316.800 186.340 317.130 ;
        RECT 159.830 316.780 160.240 316.800 ;
        RECT 159.250 316.510 159.660 316.520 ;
        RECT 159.250 316.490 182.320 316.510 ;
        RECT 159.250 316.180 182.330 316.490 ;
        RECT 159.250 316.170 159.660 316.180 ;
        RECT 158.650 315.860 159.040 315.870 ;
        RECT 158.650 315.540 178.340 315.860 ;
        RECT 158.750 315.530 178.340 315.540 ;
        RECT 158.070 315.250 158.460 315.300 ;
        RECT 152.930 315.040 153.470 315.080 ;
        RECT 140.100 315.000 153.470 315.040 ;
        RECT 140.050 314.610 153.470 315.000 ;
        RECT 158.070 314.970 174.430 315.250 ;
        RECT 158.330 314.920 174.430 314.970 ;
        RECT 62.510 312.070 127.960 314.150 ;
        RECT 140.050 312.730 142.060 314.610 ;
        RECT 152.930 314.580 153.470 314.610 ;
        RECT 157.490 314.280 170.230 314.610 ;
        RECT 153.580 314.200 154.120 314.270 ;
        RECT 144.150 313.770 154.120 314.200 ;
        RECT 164.100 313.980 166.120 314.000 ;
        RECT 156.940 313.970 166.120 313.980 ;
        RECT 144.150 312.760 146.130 313.770 ;
        RECT 156.840 313.650 166.120 313.970 ;
        RECT 156.840 313.640 157.230 313.650 ;
        RECT 154.260 313.390 154.750 313.590 ;
        RECT 148.650 313.370 154.750 313.390 ;
        RECT 148.080 313.090 154.750 313.370 ;
        RECT 148.080 312.990 154.660 313.090 ;
        RECT 156.200 312.990 162.180 313.330 ;
        RECT 148.080 312.760 150.060 312.990 ;
        RECT 154.090 312.760 154.740 312.770 ;
        RECT 140.030 312.070 142.060 312.730 ;
        RECT 144.100 312.100 146.130 312.760 ;
        RECT 148.060 312.100 150.090 312.760 ;
        RECT 152.060 312.130 154.740 312.760 ;
        RECT 155.590 312.740 156.140 312.760 ;
        RECT 160.170 312.740 162.180 312.990 ;
        RECT 155.590 312.310 158.140 312.740 ;
        RECT 161.840 312.730 162.180 312.740 ;
        RECT 152.060 312.100 154.090 312.130 ;
        RECT 156.110 312.080 158.140 312.310 ;
        RECT 160.140 312.550 162.180 312.730 ;
        RECT 164.080 312.770 166.120 313.650 ;
        RECT 164.080 312.760 166.100 312.770 ;
        RECT 164.080 312.690 166.130 312.760 ;
        RECT 168.180 312.750 170.210 314.280 ;
        RECT 168.180 312.740 170.200 312.750 ;
        RECT 168.180 312.690 170.220 312.740 ;
        RECT 160.140 312.070 162.170 312.550 ;
        RECT 164.100 312.100 166.130 312.690 ;
        RECT 168.190 312.080 170.220 312.690 ;
        RECT 172.360 312.100 174.390 314.920 ;
        RECT 176.350 312.820 178.340 315.530 ;
        RECT 176.340 312.070 178.370 312.820 ;
        RECT 180.330 312.800 182.330 316.180 ;
        RECT 180.300 312.100 182.330 312.800 ;
        RECT 184.430 312.730 186.340 316.800 ;
        RECT 188.470 312.750 190.420 317.470 ;
        RECT 192.450 312.750 194.440 318.110 ;
        RECT 196.560 318.410 198.520 318.730 ;
        RECT 200.660 318.840 202.600 319.340 ;
        RECT 196.560 312.750 198.510 318.410 ;
        RECT 200.660 312.770 202.590 318.840 ;
        RECT 184.350 312.080 186.380 312.730 ;
        RECT 188.420 312.100 190.450 312.750 ;
        RECT 192.450 312.100 194.480 312.750 ;
        RECT 196.500 312.100 198.530 312.750 ;
        RECT 58.140 100.880 60.930 104.930 ;
        RECT 58.360 100.600 60.440 100.880 ;
        RECT 62.510 76.150 64.590 312.070 ;
        RECT 200.570 311.990 202.600 312.770 ;
        RECT 230.070 312.750 230.280 313.640 ;
        RECT 228.950 312.100 230.980 312.750 ;
        RECT 232.000 312.660 232.210 313.640 ;
        RECT 232.970 313.450 233.160 313.620 ;
        RECT 232.970 313.260 237.970 313.450 ;
        RECT 233.130 312.660 235.160 312.750 ;
        RECT 237.780 312.730 237.970 313.260 ;
        RECT 238.620 312.730 238.810 312.800 ;
        RECT 241.220 312.750 243.230 330.050 ;
        RECT 232.000 312.450 235.160 312.660 ;
        RECT 233.130 312.100 235.160 312.450 ;
        RECT 237.110 312.080 239.140 312.730 ;
        RECT 241.160 312.230 243.230 312.750 ;
        RECT 241.160 312.100 243.190 312.230 ;
        RECT 224.370 309.880 224.690 310.200 ;
        RECT 225.310 309.880 225.630 310.200 ;
        RECT 66.860 306.460 127.960 308.540 ;
        RECT 62.020 72.370 64.850 76.150 ;
        RECT 62.510 71.810 64.590 72.370 ;
        RECT 66.860 47.570 68.940 306.460 ;
        RECT 71.020 301.760 127.960 303.840 ;
        RECT 66.510 43.850 69.160 47.570 ;
        RECT 66.860 43.840 68.940 43.850 ;
        RECT 71.020 18.870 73.100 301.760 ;
        RECT 70.830 15.340 73.500 18.870 ;
        RECT 132.560 9.510 135.900 301.900 ;
        RECT 335.580 246.810 337.670 333.840 ;
        RECT 339.670 275.580 341.760 339.040 ;
        RECT 343.750 304.080 345.840 343.920 ;
        RECT 347.890 332.640 349.980 349.320 ;
        RECT 347.690 329.100 350.120 332.640 ;
        RECT 347.890 328.430 349.980 329.100 ;
        RECT 343.510 300.510 346.020 304.080 ;
        RECT 339.470 271.870 341.990 275.580 ;
        RECT 339.670 271.840 341.760 271.870 ;
        RECT 335.310 243.390 337.670 246.810 ;
        RECT 335.580 242.680 337.670 243.390 ;
      LAYER via2 ;
        RECT 203.420 363.740 203.760 364.080 ;
        RECT 202.350 360.260 202.680 360.610 ;
        RECT 203.440 357.690 203.780 358.050 ;
  END
END sky130_hilas_TopProtectStructure

MACRO sky130_hilas_nFETLarge
  CLASS CORE ;
  FOREIGN sky130_hilas_nFETLarge ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.370 BY 5.830 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    USE ANALOG ;
    ANTENNAGATEAREA 6.396000 ;
    PORT
      LAYER met2 ;
        RECT 0.000 0.330 0.600 0.820 ;
        RECT 0.000 0.000 0.610 0.330 ;
    END
  END GATE
  PIN SOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 4.231200 ;
    PORT
      LAYER met2 ;
        RECT 0.330 5.590 3.390 5.600 ;
        RECT 0.240 5.260 3.390 5.590 ;
        RECT 0.240 2.810 0.560 5.260 ;
        RECT 3.060 5.250 3.370 5.260 ;
        RECT 0.240 2.480 3.400 2.810 ;
        RECT 0.240 1.440 0.560 2.480 ;
        RECT 0.240 1.120 3.400 1.440 ;
        RECT 0.860 1.110 1.170 1.120 ;
        RECT 1.960 1.110 2.270 1.120 ;
        RECT 3.060 1.110 3.370 1.120 ;
    END
  END SOURCE
  PIN DRAIN
    USE ANALOG ;
    ANTENNADIFFAREA 4.231200 ;
    PORT
      LAYER met2 ;
        RECT 1.420 4.880 1.730 4.910 ;
        RECT 2.510 4.880 2.820 4.890 ;
        RECT 1.420 4.580 4.370 4.880 ;
        RECT 2.510 4.560 2.820 4.580 ;
        RECT 3.620 4.540 4.370 4.580 ;
        RECT 3.990 4.410 4.370 4.540 ;
        RECT 4.020 3.540 4.370 4.410 ;
        RECT 1.420 3.210 4.370 3.540 ;
        RECT 4.020 0.770 4.370 3.210 ;
        RECT 1.430 0.760 4.370 0.770 ;
        RECT 1.420 0.450 4.370 0.760 ;
        RECT 1.420 0.440 4.140 0.450 ;
        RECT 1.420 0.430 1.730 0.440 ;
        RECT 2.510 0.430 2.820 0.440 ;
    END
  END DRAIN
  PIN VGND
    ANTENNADIFFAREA 1.444000 ;
    PORT
      LAYER met1 ;
        RECT 0.180 1.920 0.460 2.450 ;
        RECT 0.000 1.620 0.460 1.920 ;
        RECT 0.000 1.600 0.470 1.620 ;
        RECT 0.180 1.170 0.470 1.600 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.950 5.550 1.120 5.580 ;
        RECT 0.880 5.510 1.200 5.550 ;
        RECT 0.880 5.320 1.210 5.510 ;
        RECT 0.880 5.290 1.200 5.320 ;
        RECT 0.950 2.770 1.120 5.290 ;
        RECT 1.500 4.870 1.670 5.580 ;
        RECT 2.050 5.550 2.220 5.580 ;
        RECT 1.970 5.510 2.290 5.550 ;
        RECT 1.970 5.320 2.300 5.510 ;
        RECT 1.970 5.290 2.290 5.320 ;
        RECT 1.430 4.830 1.750 4.870 ;
        RECT 1.430 4.640 1.760 4.830 ;
        RECT 1.430 4.610 1.750 4.640 ;
        RECT 1.500 3.500 1.670 4.610 ;
        RECT 1.430 3.460 1.750 3.500 ;
        RECT 1.430 3.270 1.760 3.460 ;
        RECT 1.430 3.240 1.750 3.270 ;
        RECT 0.870 2.730 1.190 2.770 ;
        RECT 0.870 2.540 1.200 2.730 ;
        RECT 0.870 2.510 1.190 2.540 ;
        RECT 0.240 1.200 0.410 2.390 ;
        RECT 0.950 1.400 1.120 2.510 ;
        RECT 0.870 1.360 1.190 1.400 ;
        RECT 0.870 1.170 1.200 1.360 ;
        RECT 0.870 1.140 1.190 1.170 ;
        RECT 0.190 0.750 0.700 1.010 ;
        RECT 0.190 0.680 0.710 0.750 ;
        RECT 0.200 0.000 0.710 0.680 ;
        RECT 0.950 0.400 1.120 1.140 ;
        RECT 1.500 0.720 1.670 3.240 ;
        RECT 2.050 2.770 2.220 5.290 ;
        RECT 2.600 4.850 2.770 5.580 ;
        RECT 3.150 5.540 3.320 5.580 ;
        RECT 3.070 5.500 3.390 5.540 ;
        RECT 3.070 5.310 3.400 5.500 ;
        RECT 3.070 5.280 3.390 5.310 ;
        RECT 2.520 4.810 2.840 4.850 ;
        RECT 2.520 4.620 2.850 4.810 ;
        RECT 2.520 4.590 2.840 4.620 ;
        RECT 2.600 3.500 2.770 4.590 ;
        RECT 2.520 3.460 2.840 3.500 ;
        RECT 2.520 3.270 2.850 3.460 ;
        RECT 2.520 3.240 2.840 3.270 ;
        RECT 1.970 2.730 2.290 2.770 ;
        RECT 1.970 2.540 2.300 2.730 ;
        RECT 1.970 2.510 2.290 2.540 ;
        RECT 2.050 1.400 2.220 2.510 ;
        RECT 1.970 1.360 2.290 1.400 ;
        RECT 1.970 1.170 2.300 1.360 ;
        RECT 1.970 1.140 2.290 1.170 ;
        RECT 1.430 0.680 1.750 0.720 ;
        RECT 1.430 0.490 1.760 0.680 ;
        RECT 1.430 0.460 1.750 0.490 ;
        RECT 1.500 0.400 1.670 0.460 ;
        RECT 2.050 0.400 2.220 1.140 ;
        RECT 2.600 0.720 2.770 3.240 ;
        RECT 3.150 2.770 3.320 5.280 ;
        RECT 3.700 4.840 3.870 5.580 ;
        RECT 3.630 4.800 3.950 4.840 ;
        RECT 3.630 4.610 3.960 4.800 ;
        RECT 3.630 4.580 3.950 4.610 ;
        RECT 3.700 3.500 3.870 4.580 ;
        RECT 3.620 3.460 3.940 3.500 ;
        RECT 3.620 3.270 3.950 3.460 ;
        RECT 3.620 3.240 3.940 3.270 ;
        RECT 3.070 2.730 3.390 2.770 ;
        RECT 3.070 2.540 3.400 2.730 ;
        RECT 3.070 2.510 3.390 2.540 ;
        RECT 3.150 1.400 3.320 2.510 ;
        RECT 3.070 1.360 3.390 1.400 ;
        RECT 3.070 1.170 3.400 1.360 ;
        RECT 3.070 1.140 3.390 1.170 ;
        RECT 2.520 0.680 2.840 0.720 ;
        RECT 2.520 0.490 2.850 0.680 ;
        RECT 2.520 0.460 2.840 0.490 ;
        RECT 2.600 0.400 2.770 0.460 ;
        RECT 3.150 0.400 3.320 1.140 ;
        RECT 3.700 0.730 3.870 3.240 ;
        RECT 3.620 0.690 3.940 0.730 ;
        RECT 3.620 0.500 3.950 0.690 ;
        RECT 3.620 0.470 3.940 0.500 ;
        RECT 3.700 0.400 3.870 0.470 ;
      LAYER mcon ;
        RECT 0.940 5.330 1.110 5.500 ;
        RECT 2.030 5.330 2.200 5.500 ;
        RECT 1.490 4.650 1.660 4.820 ;
        RECT 1.490 3.280 1.660 3.450 ;
        RECT 0.930 2.550 1.100 2.720 ;
        RECT 0.240 2.220 0.410 2.390 ;
        RECT 0.240 1.880 0.410 2.050 ;
        RECT 0.240 1.540 0.410 1.710 ;
        RECT 0.930 1.180 1.100 1.350 ;
        RECT 0.360 0.540 0.530 0.710 ;
        RECT 3.130 5.320 3.300 5.490 ;
        RECT 2.580 4.630 2.750 4.800 ;
        RECT 2.580 3.280 2.750 3.450 ;
        RECT 2.030 2.550 2.200 2.720 ;
        RECT 2.030 1.180 2.200 1.350 ;
        RECT 1.490 0.500 1.660 0.670 ;
        RECT 3.690 4.620 3.860 4.790 ;
        RECT 3.680 3.280 3.850 3.450 ;
        RECT 3.130 2.550 3.300 2.720 ;
        RECT 3.130 1.180 3.300 1.350 ;
        RECT 2.580 0.500 2.750 0.670 ;
        RECT 3.680 0.510 3.850 0.680 ;
        RECT 0.370 0.070 0.540 0.240 ;
      LAYER met1 ;
        RECT 0.870 5.260 1.190 5.580 ;
        RECT 1.960 5.260 2.280 5.580 ;
        RECT 3.060 5.250 3.380 5.570 ;
        RECT 1.420 4.580 1.740 4.900 ;
        RECT 2.510 4.560 2.830 4.880 ;
        RECT 3.620 4.550 3.940 4.870 ;
        RECT 1.420 3.210 1.740 3.530 ;
        RECT 2.510 3.210 2.830 3.530 ;
        RECT 3.610 3.210 3.930 3.530 ;
        RECT 0.860 2.480 1.180 2.800 ;
        RECT 1.960 2.480 2.280 2.800 ;
        RECT 3.060 2.480 3.380 2.800 ;
        RECT 0.860 1.110 1.180 1.430 ;
        RECT 1.960 1.110 2.280 1.430 ;
        RECT 3.060 1.110 3.380 1.430 ;
        RECT 0.290 0.470 0.610 0.790 ;
        RECT 1.420 0.430 1.740 0.750 ;
        RECT 2.510 0.430 2.830 0.750 ;
        RECT 3.610 0.440 3.930 0.760 ;
        RECT 0.300 0.000 0.620 0.320 ;
      LAYER via ;
        RECT 0.900 5.290 1.160 5.550 ;
        RECT 1.990 5.290 2.250 5.550 ;
        RECT 3.090 5.280 3.350 5.540 ;
        RECT 1.450 4.610 1.710 4.870 ;
        RECT 2.540 4.590 2.800 4.850 ;
        RECT 3.650 4.580 3.910 4.840 ;
        RECT 1.450 3.240 1.710 3.500 ;
        RECT 2.540 3.240 2.800 3.500 ;
        RECT 3.640 3.240 3.900 3.500 ;
        RECT 0.890 2.510 1.150 2.770 ;
        RECT 1.990 2.510 2.250 2.770 ;
        RECT 3.090 2.510 3.350 2.770 ;
        RECT 0.890 1.140 1.150 1.400 ;
        RECT 1.990 1.140 2.250 1.400 ;
        RECT 3.090 1.140 3.350 1.400 ;
        RECT 0.320 0.500 0.580 0.760 ;
        RECT 1.450 0.460 1.710 0.720 ;
        RECT 2.540 0.460 2.800 0.720 ;
        RECT 3.640 0.470 3.900 0.730 ;
        RECT 0.330 0.030 0.590 0.290 ;
  END
END sky130_hilas_nFETLarge

END LIBRARY