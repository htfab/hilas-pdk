magic
tech sky130A
timestamp 1632255311
<< error_s >>
rect 63 122 103 129
rect 130 94 137 111
rect 147 98 154 121
rect 166 110 172 115
rect 63 80 103 87
rect 89 61 93 72
rect 108 62 113 67
rect 63 55 103 61
rect 32 31 40 39
rect 43 31 47 40
rect 75 39 79 55
rect 89 53 93 55
rect 101 31 106 36
rect 40 23 48 26
rect 109 23 117 31
rect 63 13 103 19
<< nmos >>
rect 63 87 103 122
rect 63 19 103 55
<< ndiff >>
rect 34 111 63 122
rect 34 94 39 111
rect 56 94 63 111
rect 34 87 63 94
rect 103 111 134 122
rect 103 94 110 111
rect 127 94 134 111
rect 103 87 134 94
rect 34 48 63 55
rect 34 31 40 48
rect 57 31 63 48
rect 34 19 63 31
rect 103 48 133 55
rect 103 31 109 48
rect 126 31 133 48
rect 103 19 133 31
<< ndiffc >>
rect 39 94 56 111
rect 110 94 127 111
rect 40 31 57 48
rect 109 31 126 48
<< psubdiff >>
rect 160 47 183 59
rect 160 30 163 47
rect 180 30 183 47
rect 160 18 183 30
<< psubdiffcont >>
rect 163 30 180 47
<< poly >>
rect 0 130 103 145
rect 63 122 103 130
rect 63 55 103 87
rect 63 6 103 19
<< locali >>
rect 0 94 39 111
rect 56 94 64 111
rect 102 94 110 111
rect 127 94 137 111
rect 0 93 64 94
rect 155 90 180 110
rect 40 48 57 56
rect 106 31 109 48
rect 126 31 135 48
rect 163 47 180 90
rect 40 26 57 31
rect 163 22 180 30
<< metal1 >>
rect 71 128 98 135
rect 71 103 108 128
rect 89 53 108 103
rect 137 0 156 152
<< metal2 >>
rect 0 109 188 129
rect 0 11 57 31
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1632251356
transform 1 0 47 0 1 26
box 0 0 34 33
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1632251332
transform 1 0 145 0 1 95
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_5
timestamp 1632251332
transform 1 0 99 0 1 33
box 0 0 23 29
use sky130_hilas_m12m2  sky130_hilas_m12m2_3
timestamp 1632251372
transform 1 0 78 0 1 113
box 0 0 32 32
<< labels >>
rlabel metal2 182 109 188 129 0 output
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
