magic
tech sky130A
timestamp 1634057788
<< checkpaint >>
rect -575 780 932 937
rect -575 -352 948 780
rect -560 -507 948 -352
rect -560 -600 939 -507
<< nwell >>
rect 0 165 404 302
<< mvnmos >>
rect 62 57 273 118
<< mvpmos >>
rect 62 199 272 261
<< mvndiff >>
rect 33 114 62 118
rect 33 97 39 114
rect 56 97 62 114
rect 33 80 62 97
rect 33 63 39 80
rect 56 63 62 80
rect 33 57 62 63
rect 273 114 302 118
rect 273 97 279 114
rect 296 97 302 114
rect 273 80 302 97
rect 273 63 279 80
rect 296 63 302 80
rect 273 57 302 63
<< mvpdiff >>
rect 33 256 62 261
rect 33 239 39 256
rect 56 239 62 256
rect 33 222 62 239
rect 33 205 39 222
rect 56 205 62 222
rect 33 199 62 205
rect 272 256 302 261
rect 272 239 278 256
rect 295 239 302 256
rect 272 222 302 239
rect 272 205 278 222
rect 295 205 302 222
rect 272 199 302 205
<< mvndiffc >>
rect 39 97 56 114
rect 39 63 56 80
rect 279 97 296 114
rect 279 63 296 80
<< mvpdiffc >>
rect 39 239 56 256
rect 39 205 56 222
rect 278 239 295 256
rect 278 205 295 222
<< psubdiff >>
rect 321 111 390 123
rect 321 94 331 111
rect 348 94 365 111
rect 382 94 390 111
rect 321 77 390 94
rect 321 60 331 77
rect 348 60 365 77
rect 382 60 390 77
rect 321 43 390 60
rect 314 26 331 43
rect 348 26 365 43
rect 382 26 390 43
rect 321 14 390 26
<< mvnsubdiff >>
rect 329 257 371 269
rect 329 240 341 257
rect 358 240 371 257
rect 329 223 371 240
rect 329 206 341 223
rect 358 206 371 223
rect 329 199 371 206
<< psubdiffcont >>
rect 331 94 348 111
rect 365 94 382 111
rect 331 60 348 77
rect 365 60 382 77
rect 331 26 348 43
rect 365 26 382 43
<< mvnsubdiffcont >>
rect 341 240 358 257
rect 341 206 358 223
<< poly >>
rect 62 261 273 276
rect 62 198 272 199
rect 62 181 273 198
rect 62 180 163 181
rect 95 153 96 180
rect 129 153 130 180
rect 236 133 237 159
rect 270 133 271 159
rect 203 132 273 133
rect 62 118 273 132
rect 62 44 273 57
<< locali >>
rect 31 296 361 302
rect 31 295 90 296
rect 98 295 197 296
rect 207 295 361 296
rect 31 292 361 295
rect 31 275 309 292
rect 326 275 344 292
rect 31 257 361 275
rect 31 256 341 257
rect 31 239 39 256
rect 56 239 278 256
rect 295 240 341 256
rect 358 240 361 257
rect 295 239 361 240
rect 31 223 360 239
rect 31 222 341 223
rect 31 205 39 222
rect 56 205 278 222
rect 295 206 341 222
rect 358 206 360 223
rect 295 205 360 206
rect 31 198 360 205
rect 31 114 163 180
rect 203 137 360 198
rect 299 117 382 119
rect 293 114 382 117
rect 31 97 39 114
rect 56 97 279 114
rect 296 111 382 114
rect 296 97 331 111
rect 31 94 331 97
rect 348 94 365 111
rect 31 80 382 94
rect 31 63 39 80
rect 56 63 279 80
rect 296 77 382 80
rect 296 63 331 77
rect 31 60 331 63
rect 348 60 365 77
rect 31 43 382 60
rect 31 26 314 43
rect 31 25 382 26
rect 307 18 382 25
<< viali >>
rect 309 275 326 292
rect 344 275 361 292
rect 314 26 331 43
rect 348 26 365 43
<< metal1 >>
rect 0 292 405 302
rect 0 275 309 292
rect 326 275 344 292
rect 361 275 405 292
rect 0 255 405 275
rect 31 254 405 255
rect 0 49 305 63
rect 0 43 405 49
rect 0 26 314 43
rect 331 26 348 43
rect 365 26 405 43
rect 0 0 405 26
use sky130_hilas_poly2li  sky130_hilas_poly2li_2
timestamp 1634057707
transform 0 1 110 -1 0 171
box 0 0 27 33
use sky130_hilas_poly2li  sky130_hilas_poly2li_1
timestamp 1634057707
transform 0 1 76 -1 0 171
box 0 0 27 33
use sky130_hilas_poly2li  sky130_hilas_poly2li_5
timestamp 1634057707
transform 0 1 144 -1 0 171
box 0 0 27 33
use sky130_hilas_poly2li  sky130_hilas_poly2li_4
timestamp 1634057707
transform 0 1 217 -1 0 150
box 0 0 27 33
use sky130_hilas_poly2li  sky130_hilas_poly2li_0
timestamp 1634057707
transform 0 1 251 -1 0 150
box 0 0 27 33
use sky130_hilas_poly2li  sky130_hilas_poly2li_3
timestamp 1634057707
transform 0 1 285 -1 0 150
box 0 0 27 33
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1634057708
transform 1 0 70 0 1 30
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1634057708
transform 1 0 106 0 1 30
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_3
timestamp 1634057708
transform 1 0 142 0 1 30
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_5
timestamp 1634057708
transform 1 0 178 0 1 30
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_2
timestamp 1634057708
transform 1 0 214 0 1 30
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_4
timestamp 1634057708
transform 1 0 250 0 1 30
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_7
timestamp 1634057708
transform 1 0 286 0 1 30
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_9
timestamp 1634057708
transform 1 0 55 0 1 278
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_10
timestamp 1634057708
transform 1 0 91 0 1 278
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_11
timestamp 1634057708
transform 1 0 127 0 1 278
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_12
timestamp 1634057708
transform 1 0 163 0 1 278
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_13
timestamp 1634057708
transform 1 0 199 0 1 278
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_14
timestamp 1634057708
transform 1 0 235 0 1 278
box 0 0 23 29
use sky130_hilas_li2m1  sky130_hilas_li2m1_15
timestamp 1634057708
transform 1 0 279 0 1 278
box 0 0 23 29
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
