magic
tech sky130A
timestamp 1629137252
<< checkpaint >>
rect -1650 2475 -217 2508
rect -1650 2079 -215 2475
rect -1650 2046 807 2079
rect -1650 1726 809 2046
rect 990 1750 3904 2079
rect 990 1726 3982 1750
rect -1650 644 3982 1726
rect -1081 540 3982 644
rect -630 -233 3982 540
rect 2142 -256 3982 -233
rect 2142 -630 3951 -256
<< error_s >>
rect 543 1021 593 1027
rect 615 1021 665 1027
rect 2584 1021 2634 1027
rect 2656 1021 2706 1027
rect 3044 1025 3071 1031
rect 543 979 593 985
rect 615 979 665 985
rect 2584 979 2634 985
rect 2656 979 2706 985
rect 3044 983 3071 989
rect 3044 958 3071 964
rect 728 877 731 927
rect 770 877 773 927
rect 864 877 866 927
rect 906 877 908 927
rect 3044 916 3071 922
rect 3044 875 3071 881
rect 728 798 731 848
rect 770 798 773 848
rect 864 798 866 848
rect 906 798 908 848
rect 3044 833 3071 839
rect 3044 808 3071 814
rect 3044 766 3071 772
rect 3044 725 3071 731
rect 728 645 731 695
rect 770 645 773 695
rect 864 645 866 695
rect 906 645 908 695
rect 3044 683 3071 689
rect 3044 658 3071 664
rect 3044 616 3071 622
rect 728 566 731 616
rect 770 566 773 616
rect 864 566 866 616
rect 906 566 908 616
rect 3044 575 3071 581
rect 3044 533 3071 539
rect 543 508 593 514
rect 615 508 665 514
rect 2584 508 2634 514
rect 2656 508 2706 514
rect 3044 508 3071 514
rect 543 466 593 472
rect 615 466 665 472
rect 2584 466 2634 472
rect 2656 466 2706 472
rect 3044 466 3071 472
<< nwell >>
rect 476 1048 807 1049
rect 2773 1048 2907 1049
rect 496 1017 528 1047
rect 2723 1017 2755 1047
rect 3158 1031 3286 1049
rect 3158 444 3286 463
<< metal1 >>
rect 512 1047 528 1049
rect 496 1045 528 1047
rect 496 1019 499 1045
rect 525 1019 528 1045
rect 553 1043 572 1049
rect 740 1038 761 1049
rect 787 1041 806 1049
rect 828 1043 849 1049
rect 936 1042 954 1049
rect 1552 1034 1594 1049
rect 1655 1034 1697 1049
rect 2025 1041 2048 1049
rect 2677 1041 2696 1049
rect 2721 1047 2749 1049
rect 2721 1045 2755 1047
rect 2721 1041 2726 1045
rect 1552 1020 1697 1034
rect 496 1017 528 1019
rect 2723 1019 2726 1041
rect 2752 1019 2755 1045
rect 3090 1035 3124 1049
rect 3156 1034 3184 1049
rect 2723 1017 2755 1019
rect 2937 492 2969 494
rect 1318 477 1350 479
rect 741 445 764 457
rect 1318 451 1321 477
rect 1347 451 1350 477
rect 1318 449 1350 451
rect 1898 477 1930 479
rect 1898 451 1901 477
rect 1927 451 1930 477
rect 2937 466 2940 492
rect 2966 466 2969 492
rect 2937 464 2969 466
rect 2937 461 2980 464
rect 3040 463 3091 464
rect 3040 461 3124 463
rect 2937 458 3124 461
rect 2952 453 3124 458
rect 1898 449 1930 451
rect 2955 450 3124 453
rect 2677 444 2696 449
rect 2721 444 2749 449
rect 2958 448 3124 450
rect 2965 447 3061 448
rect 3090 444 3124 448
rect 3157 444 3184 465
<< via1 >>
rect 499 1019 525 1045
rect 2726 1019 2752 1045
rect 1321 451 1347 477
rect 1901 451 1927 477
rect 2940 466 2966 492
<< metal2 >>
rect 496 1045 528 1047
rect 496 1019 499 1045
rect 525 1035 528 1045
rect 2723 1045 2755 1047
rect 2723 1035 2726 1045
rect 525 1019 2726 1035
rect 2752 1019 2755 1045
rect 2833 1022 2864 1046
rect 496 1017 2755 1019
rect 476 981 484 999
rect 2944 959 2966 961
rect 2939 925 2966 959
rect 2765 875 2800 897
rect 2946 868 2966 869
rect 1627 826 2426 846
rect 2946 835 2968 868
rect 2948 834 2968 835
rect 2286 758 2308 759
rect 1628 733 2311 758
rect 2404 754 2426 826
rect 2841 755 2873 779
rect 3275 778 3286 801
rect 1628 641 1979 660
rect 1956 581 1979 641
rect 2282 616 2311 733
rect 2401 750 2426 754
rect 2401 686 2427 750
rect 3275 696 3286 718
rect 2401 665 2814 686
rect 2793 651 2814 665
rect 2793 630 2994 651
rect 2282 594 2571 616
rect 2282 593 2311 594
rect 1956 566 1978 581
rect 2393 566 2993 571
rect 1956 551 2993 566
rect 1956 550 2980 551
rect 1956 544 2432 550
rect 476 494 484 512
rect 2937 492 2969 494
rect 2937 479 2940 492
rect 1318 477 2940 479
rect 1318 451 1321 477
rect 1347 464 1901 477
rect 1347 451 1350 464
rect 1318 449 1350 451
rect 1898 451 1901 464
rect 1927 466 2940 477
rect 2966 466 2969 492
rect 1927 464 2969 466
rect 1927 451 1930 464
rect 1898 449 1930 451
use sky130_hilas_FGBias2x1cell  sky130_hilas_FGBias2x1cell_0
timestamp 1628285143
transform 1 0 2016 0 1 826
box -396 -429 1258 623
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1628285143
transform 1 0 2639 0 -1 609
box 133 -454 682 609
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1629137248
transform 1 0 3131 0 1 485
box 0 0 393 746
use sky130_hilas_FGtrans2x1cell  sky130_hilas_FGtrans2x1cell_0
timestamp 1629137238
transform -1 0 1233 0 1 826
box 0 0 2257 1052
<< labels >>
rlabel metal1 3090 1043 3124 1049 0 VGND
port 11 nsew
rlabel metal1 3156 1043 3184 1049 0 VPWR
port 10 nsew
rlabel metal1 3157 444 3184 450 0 VPWR
port 10 nsew
rlabel metal1 3090 444 3124 450 0 VGND
port 11 nsew
rlabel metal2 2841 755 2873 779 0 VIN21
port 9 nsew
rlabel metal2 2833 1022 2864 1046 1 VIN22
port 8 n
rlabel metal1 741 445 764 457 0 VIN12
port 18 nsew
rlabel metal1 740 1038 761 1049 0 VIN11
port 5 nsew
rlabel metal1 1655 1042 1697 1049 0 VTUN
port 1 nsew
rlabel metal1 1552 1042 1594 1049 0 VTUN
rlabel metal1 828 1043 849 1049 0 PROG
port 3 nsew
rlabel metal1 512 1043 528 1049 0 VINJ
port 6 nsew
rlabel metal1 2721 1041 2749 1049 0 VINJ
port 6 nsew
rlabel metal2 3275 778 3286 801 0 OUTPUT1
port 13 nsew
rlabel metal2 3275 696 3286 718 0 OUTPUT2
port 12 nsew
rlabel metal1 553 1043 572 1049 0 GATESEL1
port 14 nsew
rlabel metal1 2677 444 2696 449 0 GATESEL2
port 15 nsew
rlabel metal1 2721 444 2749 449 0 VINJ
port 6 nsew
rlabel metal1 2677 1041 2696 1049 0 GATESEL2
port 15 nsew
rlabel metal2 476 981 484 999 0 DRAIN1
port 16 nsew
rlabel metal2 476 494 484 512 0 DRAIN2
port 17 nsew
rlabel metal1 2025 1041 2048 1049 0 GATE1
port 4 nsew
rlabel metal1 787 1041 806 1049 0 GATE2
port 19 nsew
rlabel metal1 936 1042 954 1049 0 RUN
port 20 nsew
<< end >>
