magic
tech sky130A
timestamp 1627061426
<< metal1 >>
rect 58 598 83 605
rect 357 598 380 605
rect 492 600 511 605
rect 357 0 380 8
rect 492 0 511 7
<< metal2 >>
rect 5 554 130 555
rect 5 538 199 554
rect 5 537 130 538
rect 564 496 572 519
rect 561 379 572 402
rect 5 367 124 369
rect 5 351 196 367
rect 5 253 57 254
rect 5 252 127 253
rect 5 236 200 252
rect 564 203 572 226
rect 563 86 572 109
rect 5 69 57 70
rect 5 52 203 69
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_0
timestamp 1625970418
transform 1 0 232 0 1 333
box -232 -40 336 119
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_3
timestamp 1625970418
transform 1 0 232 0 -1 272
box -232 -40 336 119
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_1
timestamp 1625970418
transform 1 0 232 0 -1 565
box -232 -40 336 119
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_2
timestamp 1625970418
transform 1 0 232 0 1 40
box -232 -40 336 119
<< labels >>
rlabel metal2 57 537 62 555 0 DRAIN1
port 4 nsew analog default
rlabel metal2 57 351 62 369 0 DRAIN2
port 3 nsew analog default
rlabel metal2 57 236 62 253 0 DRAIN3
port 2 nsew
rlabel metal2 57 52 62 69 0 DRAIN4
port 1 nsew
rlabel metal1 58 598 83 605 0 VINJ
port 9 nsew power default
rlabel metal1 357 598 380 605 0 DRAIN_MUX
port 10 nsew analog default
rlabel metal1 357 0 380 8 0 DRAIN_MUX
port 10 nsew analog default
rlabel metal1 492 0 511 7 0 VGND
port 11 nsew ground default
rlabel metal1 492 600 511 605 0 VGND
port 11 nsew ground default
rlabel metal2 563 86 568 109 0 SELECT4
port 12 nsew
rlabel metal2 564 203 572 226 0 SELECT3
port 13 nsew
rlabel metal2 561 379 572 402 0 SELECT2
port 14 nsew
rlabel metal2 564 496 572 519 0 SELECT1
port 15 nsew
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
