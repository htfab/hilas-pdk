magic
tech sky130A
timestamp 1629420194
<< error_s >>
rect 165 453 205 459
rect 315 453 355 459
rect 165 411 205 417
rect 315 411 355 417
rect 89 387 129 392
rect 315 385 355 392
rect 89 345 129 350
rect 315 343 355 350
rect 89 283 129 288
rect 315 283 355 290
rect 89 241 129 246
rect 315 241 355 248
rect 165 216 205 222
rect 315 216 355 222
rect 165 174 205 180
rect 315 174 355 180
rect 165 133 205 139
rect 315 133 355 139
rect 165 91 205 97
rect 315 91 355 97
rect 89 67 129 72
rect 315 65 355 72
rect 89 25 129 30
rect 315 23 355 30
rect 89 -37 129 -32
rect 315 -37 355 -30
rect 89 -79 129 -74
rect 315 -79 355 -72
rect 165 -104 205 -98
rect 315 -104 355 -98
rect 165 -146 205 -140
rect 315 -146 355 -140
<< nwell >>
rect -24 385 -23 423
<< metal1 >>
rect 38 460 58 464
rect 389 458 408 464
rect 38 -141 58 -137
rect 389 -141 408 -135
<< metal2 >>
rect -36 441 -31 461
rect -36 343 -30 363
rect 433 343 440 363
rect -36 270 -30 290
rect 433 270 440 290
rect -36 172 -31 192
rect -36 121 -31 141
rect -36 23 -30 43
rect 433 23 440 43
rect -36 -50 -30 -30
rect 433 -50 440 -30
rect -36 -148 -31 -128
use sky130_hilas_TgateSingle01  sky130_hilas_TgateSingle01_3
timestamp 1629420194
transform 1 0 227 0 1 342
box -263 -186 213 -25
use sky130_hilas_TgateSingle01  sky130_hilas_TgateSingle01_0
timestamp 1629420194
transform 1 0 227 0 -1 291
box -263 -186 213 -25
use sky130_hilas_TgateSingle01  sky130_hilas_TgateSingle01_2
timestamp 1629420194
transform 1 0 227 0 -1 -29
box -263 -186 213 -25
use sky130_hilas_TgateSingle01  sky130_hilas_TgateSingle01_1
timestamp 1629420194
transform 1 0 227 0 1 22
box -263 -186 213 -25
<< labels >>
rlabel metal2 -36 270 -30 290 0 SELECT2
port 7 nsew analog default
rlabel metal1 38 -141 58 -137 0 VPWR
port 2 nsew analog default
rlabel metal2 -36 172 -31 192 0 INPUT1_2
port 6 nsew analog default
rlabel metal1 389 458 408 464 0 VGND
port 10 nsew ground default
rlabel metal1 389 -141 408 -135 0 VGND
port 10 nsew ground default
rlabel metal2 433 270 440 290 0 OUTPUT2
port 12 nsew analog default
rlabel metal1 38 460 58 464 0 VPWR
port 2 nsew power default
rlabel metal2 433 -50 440 -30 0 OUTPUT4
port 14 nsew
rlabel metal2 433 23 440 43 0 OUTPUT3
port 15 nsew
rlabel metal2 433 343 440 363 0 OUTPUT1
port 16 nsew
rlabel metal2 -36 -148 -31 -128 0 INPUT1_4
port 17 nsew
rlabel metal2 -36 -50 -30 -30 0 SELECT4
port 18 nsew
rlabel metal2 -36 23 -30 43 0 SELECT3
port 19 nsew
rlabel metal2 -36 121 -31 141 0 INPUT1_3
port 20 nsew
rlabel metal2 -36 343 -30 363 0 SELECT1
port 21 nsew
rlabel metal2 -36 441 -31 461 0 INPUT1_1
port 22 nsew
<< end >>
