* NGSPICE file created from /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_nFETmirrorPairs.ext - technology: sky130A


* Top level circuit /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_nFETmirrorPairs

X0 VSUBS a_n66_n378# a_n66_n378# VSUBS sky130_fd_pr__nfet_01v8 w=330000u l=290000u
X1 a_n16_80# a_n66_n378# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=330000u l=290000u
X2 a_154_80# a_124_n238# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=330000u l=290000u
X3 VSUBS a_124_n238# a_124_n238# VSUBS sky130_fd_pr__nfet_01v8 w=330000u l=290000u
.end

