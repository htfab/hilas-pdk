magic
tech sky130A
timestamp 1629420194
<< nwell >>
rect -363 -444 -177 -145
<< mvpmos >>
rect -298 -396 -248 -193
<< mvpdiff >>
rect -329 -200 -298 -193
rect -329 -217 -322 -200
rect -305 -217 -298 -200
rect -329 -234 -298 -217
rect -329 -251 -322 -234
rect -305 -251 -298 -234
rect -329 -268 -298 -251
rect -329 -285 -322 -268
rect -305 -285 -298 -268
rect -329 -302 -298 -285
rect -329 -319 -322 -302
rect -305 -319 -298 -302
rect -329 -336 -298 -319
rect -329 -353 -322 -336
rect -305 -353 -298 -336
rect -329 -370 -298 -353
rect -329 -387 -322 -370
rect -305 -387 -298 -370
rect -329 -396 -298 -387
rect -248 -201 -210 -193
rect -248 -218 -241 -201
rect -224 -218 -210 -201
rect -248 -235 -210 -218
rect -248 -252 -241 -235
rect -224 -252 -210 -235
rect -248 -269 -210 -252
rect -248 -286 -241 -269
rect -224 -286 -210 -269
rect -248 -303 -210 -286
rect -248 -320 -241 -303
rect -224 -320 -210 -303
rect -248 -337 -210 -320
rect -248 -354 -241 -337
rect -224 -354 -210 -337
rect -248 -371 -210 -354
rect -248 -388 -241 -371
rect -224 -388 -210 -371
rect -248 -396 -210 -388
<< mvpdiffc >>
rect -322 -217 -305 -200
rect -322 -251 -305 -234
rect -322 -285 -305 -268
rect -322 -319 -305 -302
rect -322 -353 -305 -336
rect -322 -387 -305 -370
rect -241 -218 -224 -201
rect -241 -252 -224 -235
rect -241 -286 -224 -269
rect -241 -320 -224 -303
rect -241 -354 -224 -337
rect -241 -388 -224 -371
<< poly >>
rect -298 -193 -248 -175
rect -298 -411 -248 -396
<< locali >>
rect -322 -200 -304 -192
rect -305 -217 -304 -200
rect -322 -234 -304 -217
rect -305 -251 -304 -234
rect -322 -268 -304 -251
rect -305 -285 -304 -268
rect -322 -302 -304 -285
rect -305 -319 -304 -302
rect -322 -336 -304 -319
rect -305 -353 -304 -336
rect -322 -370 -304 -353
rect -305 -387 -304 -370
rect -241 -201 -224 -193
rect -241 -235 -224 -218
rect -241 -269 -224 -252
rect -241 -303 -224 -286
rect -241 -337 -224 -320
rect -241 -371 -224 -354
rect -322 -397 -304 -387
rect -249 -388 -241 -371
rect -224 -388 -216 -371
<< end >>
