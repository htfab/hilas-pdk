magic
tech sky130A
timestamp 1628616750
<< nwell >>
rect 0 0 119 287
<< pmos >>
rect 47 18 73 269
<< pdiff >>
rect 18 245 47 269
rect 18 228 24 245
rect 41 228 47 245
rect 18 211 47 228
rect 18 194 24 211
rect 41 194 47 211
rect 18 177 47 194
rect 18 160 24 177
rect 41 160 47 177
rect 18 143 47 160
rect 18 126 24 143
rect 41 126 47 143
rect 18 109 47 126
rect 18 92 24 109
rect 41 92 47 109
rect 18 75 47 92
rect 18 58 24 75
rect 41 58 47 75
rect 18 41 47 58
rect 18 24 24 41
rect 41 24 47 41
rect 18 18 47 24
rect 73 245 101 269
rect 73 228 79 245
rect 96 228 101 245
rect 73 211 101 228
rect 73 194 79 211
rect 96 194 101 211
rect 73 177 101 194
rect 73 160 79 177
rect 96 160 101 177
rect 73 143 101 160
rect 73 126 79 143
rect 96 126 101 143
rect 73 109 101 126
rect 73 92 79 109
rect 96 92 101 109
rect 73 75 101 92
rect 73 58 79 75
rect 96 58 101 75
rect 73 41 101 58
rect 73 24 79 41
rect 96 24 101 41
rect 73 18 101 24
<< pdiffc >>
rect 24 228 41 245
rect 24 194 41 211
rect 24 160 41 177
rect 24 126 41 143
rect 24 92 41 109
rect 24 58 41 75
rect 24 24 41 41
rect 79 228 96 245
rect 79 194 96 211
rect 79 160 96 177
rect 79 126 96 143
rect 79 92 96 109
rect 79 58 96 75
rect 79 24 96 41
<< poly >>
rect 47 269 73 282
rect 47 5 73 18
<< locali >>
rect 24 245 41 264
rect 24 211 41 228
rect 24 177 41 194
rect 24 143 41 160
rect 24 109 41 126
rect 24 75 41 92
rect 24 41 41 58
rect 24 15 41 24
rect 79 245 96 264
rect 79 211 96 228
rect 79 177 96 194
rect 79 143 96 160
rect 79 109 96 126
rect 79 75 96 92
rect 79 41 96 58
rect 79 14 96 24
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
