magic
tech sky130A
timestamp 1632488964
<< nwell >>
rect -173 126 244 333
<< pmos >>
rect -116 243 137 314
rect -116 144 137 214
<< pdiff >>
rect -154 308 -116 314
rect -154 249 -145 308
rect -127 249 -116 308
rect -154 243 -116 249
rect 137 306 182 314
rect 137 243 155 306
rect 146 214 155 243
rect -152 208 -116 214
rect -152 149 -145 208
rect -127 149 -116 208
rect -152 144 -116 149
rect 137 149 155 214
rect 173 149 182 306
rect 137 144 182 149
<< pdiffc >>
rect -145 249 -127 308
rect -145 149 -127 208
rect 155 149 173 306
<< nsubdiff >>
rect 182 304 224 314
rect 182 149 194 304
rect 212 149 224 304
rect 182 144 224 149
<< nsubdiffcont >>
rect 194 149 212 304
<< poly >>
rect -116 314 137 330
rect -116 214 137 243
rect -116 120 137 144
rect -116 103 -108 120
rect 129 103 137 120
rect -116 98 137 103
<< polycont >>
rect -108 103 129 120
<< locali >>
rect -145 308 -127 316
rect -145 241 -127 249
rect 146 306 216 318
rect -145 208 -127 216
rect -145 141 -127 149
rect 146 149 155 306
rect 173 304 216 306
rect 173 287 175 304
rect 192 287 194 304
rect 173 267 194 287
rect 173 250 175 267
rect 192 250 194 267
rect 173 231 194 250
rect 173 214 175 231
rect 192 214 194 231
rect 173 195 194 214
rect 173 178 175 195
rect 192 178 194 195
rect 173 159 194 178
rect 173 149 175 159
rect 146 142 175 149
rect 192 149 194 159
rect 212 149 216 304
rect 192 142 216 149
rect -145 120 -128 141
rect 146 138 216 142
rect -145 103 -108 120
rect 129 103 137 120
<< viali >>
rect 175 287 192 304
rect 175 250 192 267
rect 175 214 192 231
rect 175 178 192 195
rect 175 142 192 159
<< metal1 >>
rect 161 304 204 321
rect 161 287 175 304
rect 192 287 204 304
rect 161 267 204 287
rect 161 250 175 267
rect 192 250 204 267
rect 161 231 204 250
rect 161 214 175 231
rect 192 214 204 231
rect 161 195 204 214
rect 161 178 175 195
rect 192 178 204 195
rect 161 159 204 178
rect 161 142 175 159
rect 192 142 204 159
rect 161 132 204 142
<< end >>
