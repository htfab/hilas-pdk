magic
tech sky130A
timestamp 1627400756
<< error_s >>
rect 514 572 543 588
rect 593 572 622 588
rect 672 572 701 588
rect 751 572 780 588
rect 997 574 1026 592
rect 1153 574 1182 592
rect 1399 572 1428 588
rect 1478 572 1507 588
rect 1557 572 1586 588
rect 1636 572 1665 588
rect 997 542 998 543
rect 1025 542 1026 543
rect 1153 542 1154 543
rect 1181 542 1182 543
rect 514 538 515 539
rect 542 538 543 539
rect 593 538 594 539
rect 621 538 622 539
rect 672 538 673 539
rect 700 538 701 539
rect 751 538 752 539
rect 779 538 780 539
rect 464 509 481 538
rect 513 537 544 538
rect 592 537 623 538
rect 671 537 702 538
rect 750 537 781 538
rect 514 530 543 537
rect 593 530 622 537
rect 672 530 701 537
rect 751 530 780 537
rect 514 516 523 530
rect 770 516 780 530
rect 514 510 543 516
rect 593 510 622 516
rect 672 510 701 516
rect 751 510 780 516
rect 513 509 544 510
rect 592 509 623 510
rect 671 509 702 510
rect 750 509 781 510
rect 812 509 830 538
rect 947 513 965 542
rect 996 541 1027 542
rect 997 532 1026 541
rect 997 523 1007 532
rect 1016 523 1026 532
rect 997 514 1026 523
rect 996 513 1027 514
rect 1058 513 1076 542
rect 1103 513 1121 542
rect 1152 541 1183 542
rect 1153 532 1182 541
rect 1153 523 1163 532
rect 1172 523 1182 532
rect 1153 514 1182 523
rect 1152 513 1183 514
rect 1214 513 1232 542
rect 1399 538 1400 539
rect 1427 538 1428 539
rect 1478 538 1479 539
rect 1506 538 1507 539
rect 1557 538 1558 539
rect 1585 538 1586 539
rect 1636 538 1637 539
rect 1664 538 1665 539
rect 997 512 998 513
rect 1025 512 1026 513
rect 1153 512 1154 513
rect 1181 512 1182 513
rect 1349 509 1367 538
rect 1398 537 1429 538
rect 1477 537 1508 538
rect 1556 537 1587 538
rect 1635 537 1666 538
rect 1399 530 1428 537
rect 1478 530 1507 537
rect 1557 530 1586 537
rect 1636 530 1665 537
rect 1399 516 1409 530
rect 1656 516 1665 530
rect 1399 510 1428 516
rect 1478 510 1507 516
rect 1557 510 1586 516
rect 1636 510 1665 516
rect 1398 509 1429 510
rect 1477 509 1508 510
rect 1556 509 1587 510
rect 1635 509 1666 510
rect 1698 509 1715 538
rect 1732 516 1734 517
rect 514 508 515 509
rect 542 508 543 509
rect 593 508 594 509
rect 621 508 622 509
rect 672 508 673 509
rect 700 508 701 509
rect 751 508 752 509
rect 779 508 780 509
rect 1399 508 1400 509
rect 1427 508 1428 509
rect 1478 508 1479 509
rect 1506 508 1507 509
rect 1557 508 1558 509
rect 1585 508 1586 509
rect 1636 508 1637 509
rect 1664 508 1665 509
rect 514 459 543 474
rect 593 459 622 474
rect 672 459 701 474
rect 751 459 780 474
rect 997 463 1026 481
rect 1153 463 1182 481
rect 1399 459 1428 474
rect 1478 459 1507 474
rect 1557 459 1586 474
rect 1636 459 1665 474
rect 514 425 543 441
rect 593 425 622 441
rect 672 425 701 441
rect 751 425 780 441
rect 997 422 1026 440
rect 1153 422 1182 440
rect 1399 425 1428 441
rect 1478 425 1507 441
rect 1557 425 1586 441
rect 1636 425 1665 441
rect 514 391 515 392
rect 542 391 543 392
rect 593 391 594 392
rect 621 391 622 392
rect 672 391 673 392
rect 700 391 701 392
rect 751 391 752 392
rect 779 391 780 392
rect 1399 391 1400 392
rect 1427 391 1428 392
rect 1478 391 1479 392
rect 1506 391 1507 392
rect 1557 391 1558 392
rect 1585 391 1586 392
rect 1636 391 1637 392
rect 1664 391 1665 392
rect 464 362 481 391
rect 513 390 544 391
rect 592 390 623 391
rect 671 390 702 391
rect 750 390 781 391
rect 514 383 543 390
rect 593 383 622 390
rect 672 383 701 390
rect 751 383 780 390
rect 514 369 523 383
rect 770 369 780 383
rect 514 363 543 369
rect 593 363 622 369
rect 672 363 701 369
rect 751 363 780 369
rect 513 362 544 363
rect 592 362 623 363
rect 671 362 702 363
rect 750 362 781 363
rect 812 362 830 391
rect 997 390 998 391
rect 1025 390 1026 391
rect 1153 390 1154 391
rect 1181 390 1182 391
rect 514 361 515 362
rect 542 361 543 362
rect 593 361 594 362
rect 621 361 622 362
rect 672 361 673 362
rect 700 361 701 362
rect 751 361 752 362
rect 779 361 780 362
rect 947 361 965 390
rect 996 389 1027 390
rect 997 380 1026 389
rect 997 371 1007 380
rect 1016 371 1026 380
rect 997 362 1026 371
rect 996 361 1027 362
rect 1058 361 1076 390
rect 1103 361 1121 390
rect 1152 389 1183 390
rect 1153 380 1182 389
rect 1153 371 1163 380
rect 1172 371 1182 380
rect 1153 362 1182 371
rect 1152 361 1183 362
rect 1214 361 1232 390
rect 1349 362 1367 391
rect 1398 390 1429 391
rect 1477 390 1508 391
rect 1556 390 1587 391
rect 1635 390 1666 391
rect 1399 383 1428 390
rect 1478 383 1507 390
rect 1557 383 1586 390
rect 1636 383 1665 390
rect 1399 369 1409 383
rect 1656 369 1665 383
rect 1399 363 1428 369
rect 1478 363 1507 369
rect 1557 363 1586 369
rect 1636 363 1665 369
rect 1398 362 1429 363
rect 1477 362 1508 363
rect 1556 362 1587 363
rect 1635 362 1666 363
rect 1698 362 1715 391
rect 1399 361 1400 362
rect 1427 361 1428 362
rect 1478 361 1479 362
rect 1506 361 1507 362
rect 1557 361 1558 362
rect 1585 361 1586 362
rect 1636 361 1637 362
rect 1664 361 1665 362
rect 997 360 998 361
rect 1025 360 1026 361
rect 1153 360 1154 361
rect 1181 360 1182 361
rect 514 312 543 327
rect 593 312 622 327
rect 672 312 701 327
rect 751 312 780 327
rect 997 311 1026 329
rect 1153 311 1182 329
rect 1399 312 1428 327
rect 1478 312 1507 327
rect 1557 312 1586 327
rect 1636 312 1665 327
rect 514 278 543 294
rect 593 278 622 294
rect 672 278 701 294
rect 751 278 780 294
rect 997 277 1026 295
rect 1153 277 1182 295
rect 1399 278 1428 294
rect 1478 278 1507 294
rect 1557 278 1586 294
rect 1636 278 1665 294
rect 997 245 998 246
rect 1025 245 1026 246
rect 1153 245 1154 246
rect 1181 245 1182 246
rect 514 244 515 245
rect 542 244 543 245
rect 593 244 594 245
rect 621 244 622 245
rect 672 244 673 245
rect 700 244 701 245
rect 751 244 752 245
rect 779 244 780 245
rect 464 215 481 244
rect 513 243 544 244
rect 592 243 623 244
rect 671 243 702 244
rect 750 243 781 244
rect 514 236 543 243
rect 593 236 622 243
rect 672 236 701 243
rect 751 236 780 243
rect 514 222 523 236
rect 770 222 780 236
rect 514 216 543 222
rect 593 216 622 222
rect 672 216 701 222
rect 751 216 780 222
rect 513 215 544 216
rect 592 215 623 216
rect 671 215 702 216
rect 750 215 781 216
rect 812 215 830 244
rect 947 216 965 245
rect 996 244 1027 245
rect 997 235 1026 244
rect 997 226 1007 235
rect 1016 226 1026 235
rect 997 217 1026 226
rect 996 216 1027 217
rect 1058 216 1076 245
rect 1103 216 1121 245
rect 1152 244 1183 245
rect 1153 235 1182 244
rect 1153 226 1163 235
rect 1172 226 1182 235
rect 1153 217 1182 226
rect 1152 216 1183 217
rect 1214 216 1232 245
rect 1399 244 1400 245
rect 1427 244 1428 245
rect 1478 244 1479 245
rect 1506 244 1507 245
rect 1557 244 1558 245
rect 1585 244 1586 245
rect 1636 244 1637 245
rect 1664 244 1665 245
rect 997 215 998 216
rect 1025 215 1026 216
rect 1153 215 1154 216
rect 1181 215 1182 216
rect 1349 215 1367 244
rect 1398 243 1429 244
rect 1477 243 1508 244
rect 1556 243 1587 244
rect 1635 243 1666 244
rect 1399 236 1428 243
rect 1478 236 1507 243
rect 1557 236 1586 243
rect 1636 236 1665 243
rect 1399 222 1409 236
rect 1656 222 1665 236
rect 1399 216 1428 222
rect 1478 216 1507 222
rect 1557 216 1586 222
rect 1636 216 1665 222
rect 1398 215 1429 216
rect 1477 215 1508 216
rect 1556 215 1587 216
rect 1635 215 1666 216
rect 1698 215 1715 244
rect 514 214 515 215
rect 542 214 543 215
rect 593 214 594 215
rect 621 214 622 215
rect 672 214 673 215
rect 700 214 701 215
rect 751 214 752 215
rect 779 214 780 215
rect 1399 214 1400 215
rect 1427 214 1428 215
rect 1478 214 1479 215
rect 1506 214 1507 215
rect 1557 214 1558 215
rect 1585 214 1586 215
rect 1636 214 1637 215
rect 1664 214 1665 215
rect 514 165 543 180
rect 593 165 622 180
rect 672 165 701 180
rect 751 165 780 180
rect 997 166 1026 184
rect 1153 166 1182 184
rect 1399 165 1428 180
rect 1478 165 1507 180
rect 1557 165 1586 180
rect 1636 165 1665 180
rect 514 131 543 147
rect 593 131 622 147
rect 672 131 701 147
rect 751 131 780 147
rect 997 123 1026 141
rect 1153 123 1182 141
rect 1399 131 1428 147
rect 1478 131 1507 147
rect 1557 131 1586 147
rect 1636 131 1665 147
rect 514 97 515 98
rect 542 97 543 98
rect 593 97 594 98
rect 621 97 622 98
rect 672 97 673 98
rect 700 97 701 98
rect 751 97 752 98
rect 779 97 780 98
rect 1399 97 1400 98
rect 1427 97 1428 98
rect 1478 97 1479 98
rect 1506 97 1507 98
rect 1557 97 1558 98
rect 1585 97 1586 98
rect 1636 97 1637 98
rect 1664 97 1665 98
rect 464 68 481 97
rect 513 96 544 97
rect 592 96 623 97
rect 671 96 702 97
rect 750 96 781 97
rect 514 89 543 96
rect 593 89 622 96
rect 672 89 701 96
rect 751 89 780 96
rect 514 75 523 89
rect 770 75 780 89
rect 514 69 543 75
rect 593 69 622 75
rect 672 69 701 75
rect 751 69 780 75
rect 513 68 544 69
rect 592 68 623 69
rect 671 68 702 69
rect 750 68 781 69
rect 812 68 830 97
rect 997 91 998 92
rect 1025 91 1026 92
rect 1153 91 1154 92
rect 1181 91 1182 92
rect 514 67 515 68
rect 542 67 543 68
rect 593 67 594 68
rect 621 67 622 68
rect 672 67 673 68
rect 700 67 701 68
rect 751 67 752 68
rect 779 67 780 68
rect 947 62 965 91
rect 996 90 1027 91
rect 997 81 1026 90
rect 997 72 1007 81
rect 1016 72 1026 81
rect 997 63 1026 72
rect 996 62 1027 63
rect 1058 62 1076 91
rect 1103 62 1121 91
rect 1152 90 1183 91
rect 1153 81 1182 90
rect 1153 72 1163 81
rect 1172 72 1182 81
rect 1153 63 1182 72
rect 1152 62 1183 63
rect 1214 62 1232 91
rect 1349 68 1367 97
rect 1398 96 1429 97
rect 1477 96 1508 97
rect 1556 96 1587 97
rect 1635 96 1666 97
rect 1399 89 1428 96
rect 1478 89 1507 96
rect 1557 89 1586 96
rect 1636 89 1665 96
rect 1399 75 1409 89
rect 1656 75 1665 89
rect 1399 69 1428 75
rect 1478 69 1507 75
rect 1557 69 1586 75
rect 1636 69 1665 75
rect 1398 68 1429 69
rect 1477 68 1508 69
rect 1556 68 1587 69
rect 1635 68 1666 69
rect 1698 68 1715 97
rect 1399 67 1400 68
rect 1427 67 1428 68
rect 1478 67 1479 68
rect 1506 67 1507 68
rect 1557 67 1558 68
rect 1585 67 1586 68
rect 1636 67 1637 68
rect 1664 67 1665 68
rect 997 61 998 62
rect 1025 61 1026 62
rect 1153 61 1154 62
rect 1181 61 1182 62
rect 514 18 543 33
rect 593 18 622 33
rect 672 18 701 33
rect 751 18 780 33
rect 997 12 1026 30
rect 1153 12 1182 30
rect 1399 18 1428 33
rect 1478 18 1507 33
rect 1557 18 1586 33
rect 1636 18 1665 33
<< metal1 >>
rect 227 599 243 605
rect 268 599 287 605
rect 308 599 324 605
rect 227 1 243 8
rect 268 1 287 8
rect 308 1 324 8
rect 635 0 660 605
rect 996 0 1026 605
rect 1154 0 1184 605
rect 1520 0 1544 605
rect 1855 598 1871 605
rect 1892 598 1911 605
rect 1936 598 1952 605
rect 1855 1 1871 8
rect 1892 1 1911 8
rect 1936 1 1952 8
<< metal2 >>
rect 191 537 199 555
rect 1977 537 1988 555
rect 191 494 199 512
rect 1978 494 1989 512
rect 191 394 199 412
rect 1978 394 1989 412
rect 191 351 199 369
rect 431 361 443 369
rect 1740 355 1752 369
rect 1978 351 1989 369
rect 191 236 198 254
rect 1977 236 1988 254
rect 191 193 198 211
rect 1977 193 1988 211
rect 191 94 198 112
rect 1977 94 1988 112
rect 191 51 198 69
rect 1977 51 1988 69
use sky130_hilas_swc4x1cellOverlap2  sky130_hilas_swc4x1cellOverlap2_1
timestamp 1607392100
transform -1 0 935 0 1 382
box -191 -382 744 223
use sky130_hilas_swc4x1cellOverlap2  sky130_hilas_swc4x1cellOverlap2_0
timestamp 1607392100
transform 1 0 1244 0 1 382
box -191 -382 744 223
<< labels >>
rlabel metal1 308 599 324 605 0 VERT1
port 1 nsew analog default
rlabel metal1 227 599 243 605 0 VINJ
port 10 nsew
rlabel metal1 268 599 287 605 0 GATESELECT1
port 11 nsew analog default
rlabel metal2 191 537 199 555 0 DRAIN1
port 3 nsew analog default
rlabel metal2 191 494 199 512 0 HORIZ1
port 2 nsew analog default
rlabel metal2 191 394 199 412 0 HORIZ2
port 4 nsew analog default
rlabel metal2 191 351 199 369 0 DRAIN2
port 5 nsew analog default
rlabel metal2 191 236 198 254 0 DRAIN3
port 6 nsew analog default
rlabel metal2 191 193 198 211 0 HORIZ3
port 7 nsew analog default
rlabel metal2 191 94 198 112 0 HORIZ4
port 8 nsew analog default
rlabel metal2 191 51 198 69 0 DRAIN4
port 9 nsew analog default
rlabel metal1 227 1 243 8 0 VINJ
port 10 nsew power default
rlabel metal1 308 1 324 8 0 VERT1
port 1 nsew analog default
rlabel metal1 268 1 287 8 0 GATESELECT1
port 11 nsew analog default
rlabel metal1 1936 1 1952 8 0 VINJ
port 10 nsew power default
rlabel metal1 1855 598 1871 605 0 VERT2
port 12 nsew analog default
rlabel metal1 1892 598 1911 605 0 GATESELECT2
port 13 nsew analog default
rlabel metal1 1936 598 1952 605 0 VINJ
port 10 nsew power default
rlabel metal1 1855 1 1871 8 0 VERT2
port 12 nsew analog default
rlabel metal1 1892 1 1911 8 0 GATESELECT2
port 13 nsew analog default
rlabel metal2 1977 537 1988 555 0 DRAIN1
port 3 nsew analog default
rlabel metal2 1978 494 1989 512 0 HORIZ1
port 2 nsew analog default
rlabel metal2 1978 394 1989 412 0 HORIZ2
port 4 nsew analog default
rlabel metal2 1978 351 1989 369 0 DRAIN2
port 5 nsew analog default
rlabel metal2 1977 236 1988 254 0 DRAIN3
port 6 nsew analog default
rlabel metal2 1977 193 1988 211 0 HORIZ3
port 7 nsew analog default
rlabel metal2 1977 94 1988 112 0 HORIZ4
port 8 nsew analog default
rlabel metal2 1977 51 1988 69 0 DRAIN
port 14 nsew analog default
rlabel metal1 1520 600 1544 605 0 GATE2
port 15 nsew analog default
rlabel metal1 1520 0 1544 6 0 GATE2
port 15 nsew analog default
rlabel metal1 635 599 660 605 0 GATE1
port 16 nsew analog default
rlabel metal1 635 0 660 6 0 GATE1
port 16 nsew analog default
rlabel metal1 996 597 1026 605 0 VTUN
port 17 nsew analog default
rlabel metal1 1154 597 1184 605 0 VTUN
rlabel metal1 996 0 1026 8 0 VTUN
port 17 nsew analog default
rlabel metal1 1154 0 1184 8 0 VTUN
port 17 nsew analog default
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
