* Copyright 2020 The Hilas PDK Authors
* 
* This file is part of HILAS.
* 
* HILAS is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published by
* the Free Software Foundation, version 3 of the License.
* 
* HILAS is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
* 
* You should have received a copy of the GNU Lesser General Public License
* along with HILAS.  If not, see <https://www.gnu.org/licenses/>.
* 
* Licensed under the Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
* https://www.gnu.org/licenses/lgpl-3.0.en.html
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
* SPDX-License-Identifier: LGPL-3.0
* 
* 

* NGSPICE file created from sky130_hilas_FGtrans2x1cell.ext - technology: sky130A

.subckt sky130_hilas_TunCap01 VSUBS a_n2872_n666# w_n2902_n800#
X0 a_n2872_n666# w_n2902_n800# w_n2902_n800# sky130_fd_pr__cap_var w=590000u l=500000u
.ends

.subckt sky130_hilas_horizTransCell01 VSUBS a_n512_284# a_n952_238# a_n346_284# a_n654_284#
+ a_n926_284# a_n952_338# a_n952_496# a_n654_438# a_n926_438# a_n300_130# a_n512_162#
+ w_n728_96# a_n654_596# a_n926_596#
X0 a_n654_438# a_n952_338# a_n654_284# w_n728_96# sky130_fd_pr__pfet_g5v0d10v5 w=390000u l=500000u
X1 w_n728_96# a_n300_130# a_n344_162# w_n728_96# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
X2 a_n346_284# a_n952_238# a_n512_284# w_n728_96# sky130_fd_pr__pfet_g5v0d10v5 w=1.84e+06u l=510000u
X3 a_n344_162# a_n952_238# a_n512_162# w_n728_96# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
X4 a_n926_596# a_n952_496# a_n926_438# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=400000u l=500000u
X5 a_n926_438# a_n952_338# a_n926_284# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=400000u l=500000u
X6 a_n654_596# a_n952_496# a_n654_438# w_n728_96# sky130_fd_pr__pfet_g5v0d10v5 w=390000u l=500000u
.ends

.subckt sky130_hilas_FGVaractorCapacitor02 VSUBS a_n1882_n644# w_n2010_n760#
X0 a_n1882_n644# w_n2010_n760# w_n2010_n760# sky130_fd_pr__cap_var w=1.11e+06u l=500000u
.ends

.subckt sky130_hilas_FGtrans2x1cell GATESELECT VINJ FGDRAINPROGRAM1 DRAIN4 PROG RUN
+ GATE1 GATE2 PROGGATE VGND VTUN DRAIN VS
Xsky130_hilas_TunCap01_1 VGND a_n560_n620# VTUN sky130_hilas_TunCap01
Xsky130_hilas_horizTransCell01_0 VGND DRAIN a_n560_n620# VS PROGGATE GATE1 RUN PROG
+ li_724_n408# li_724_n408# GATESELECT DRAIN4 VINJ GATE1 PROGGATE sky130_hilas_horizTransCell01
Xsky130_hilas_TunCap01_3 VGND a_n474_252# VTUN sky130_hilas_TunCap01
Xsky130_hilas_horizTransCell01_1 VGND FGDRAINPROGRAM1 a_n474_252# VS PROGGATE GATE2
+ RUN PROG li_724_56# li_724_56# GATESELECT FGDRAINPROGRAM1 VINJ GATE2 PROGGATE sky130_hilas_horizTransCell01
Xsky130_hilas_FGVaractorCapacitor02_0 VGND a_n560_n620# li_724_n408# sky130_hilas_FGVaractorCapacitor02
Xsky130_hilas_FGVaractorCapacitor02_2 VGND a_n474_252# li_724_56# sky130_hilas_FGVaractorCapacitor02
.ends

