VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO swc4x2cell
  CLASS BLOCK ;
  FOREIGN swc4x2cell ;
  ORIGIN 10.040 0.040 ;
  SIZE 20.120 BY 6.050 ;
  OBS
      LAYER li1 ;
        RECT -9.640 5.330 -9.440 5.680 ;
        RECT -8.160 5.430 -7.630 5.600 ;
        RECT 7.670 5.430 8.200 5.600 ;
        RECT -9.650 5.300 -9.440 5.330 ;
        RECT 9.480 5.330 9.680 5.680 ;
        RECT -9.650 4.710 -9.430 5.300 ;
        RECT -8.910 4.740 -8.710 5.310 ;
        RECT -8.160 4.810 -7.630 4.980 ;
        RECT 7.670 4.810 8.200 4.980 ;
        RECT 8.750 4.740 8.950 5.310 ;
        RECT 9.480 5.300 9.690 5.330 ;
        RECT 9.470 4.710 9.690 5.300 ;
        RECT -9.650 3.680 -9.430 4.270 ;
        RECT -9.650 3.650 -9.440 3.680 ;
        RECT -8.910 3.670 -8.710 4.240 ;
        RECT -8.160 4.000 -7.630 4.170 ;
        RECT 7.670 4.000 8.200 4.170 ;
        RECT 8.750 3.670 8.950 4.240 ;
        RECT 9.470 3.680 9.690 4.270 ;
        RECT -9.640 3.300 -9.440 3.650 ;
        RECT 9.480 3.650 9.690 3.680 ;
        RECT -8.160 3.380 -7.630 3.550 ;
        RECT 7.670 3.380 8.200 3.550 ;
        RECT 9.480 3.300 9.680 3.650 ;
        RECT -9.270 2.900 -8.830 3.070 ;
        RECT -4.970 2.690 -4.420 3.120 ;
        RECT -0.940 2.760 -0.390 3.190 ;
        RECT 0.430 2.760 0.980 3.190 ;
        RECT 4.460 2.690 5.010 3.120 ;
        RECT 8.870 2.900 9.310 3.070 ;
        RECT -9.640 2.320 -9.440 2.670 ;
        RECT -8.160 2.420 -7.630 2.590 ;
        RECT 7.670 2.420 8.200 2.590 ;
        RECT -9.650 2.290 -9.440 2.320 ;
        RECT 9.480 2.320 9.680 2.670 ;
        RECT -9.650 1.700 -9.430 2.290 ;
        RECT -8.910 1.730 -8.710 2.300 ;
        RECT -8.160 1.800 -7.630 1.970 ;
        RECT 7.670 1.800 8.200 1.970 ;
        RECT 8.750 1.730 8.950 2.300 ;
        RECT 9.480 2.290 9.690 2.320 ;
        RECT 9.470 1.700 9.690 2.290 ;
        RECT -9.650 0.680 -9.430 1.270 ;
        RECT -9.650 0.650 -9.440 0.680 ;
        RECT -8.910 0.670 -8.710 1.240 ;
        RECT -8.160 1.000 -7.630 1.170 ;
        RECT 7.670 1.000 8.200 1.170 ;
        RECT 8.750 0.670 8.950 1.240 ;
        RECT 9.470 0.680 9.690 1.270 ;
        RECT -9.640 0.300 -9.440 0.650 ;
        RECT 9.480 0.650 9.690 0.680 ;
        RECT -8.160 0.380 -7.630 0.550 ;
        RECT 7.670 0.380 8.200 0.550 ;
        RECT 9.480 0.300 9.680 0.650 ;
      LAYER mcon ;
        RECT -7.810 5.430 -7.630 5.600 ;
        RECT -9.620 5.130 -9.450 5.300 ;
        RECT -8.890 5.100 -8.720 5.270 ;
        RECT 8.760 5.100 8.930 5.270 ;
        RECT -7.810 4.810 -7.630 4.980 ;
        RECT 9.490 5.130 9.660 5.300 ;
        RECT -9.620 3.680 -9.450 3.850 ;
        RECT -7.810 4.000 -7.630 4.170 ;
        RECT -8.890 3.710 -8.720 3.880 ;
        RECT 8.760 3.710 8.930 3.880 ;
        RECT 9.490 3.680 9.660 3.850 ;
        RECT -7.810 3.380 -7.630 3.550 ;
        RECT -4.690 2.770 -4.420 3.040 ;
        RECT -0.660 2.840 -0.390 3.110 ;
        RECT 0.430 2.840 0.700 3.110 ;
        RECT 4.460 2.770 4.730 3.040 ;
        RECT 9.130 2.900 9.310 3.070 ;
        RECT -7.810 2.420 -7.630 2.590 ;
        RECT -9.620 2.120 -9.450 2.290 ;
        RECT -8.890 2.090 -8.720 2.260 ;
        RECT 8.760 2.090 8.930 2.260 ;
        RECT -7.810 1.800 -7.630 1.970 ;
        RECT 9.490 2.120 9.660 2.290 ;
        RECT -9.620 0.680 -9.450 0.850 ;
        RECT -7.810 1.000 -7.630 1.170 ;
        RECT -8.890 0.710 -8.720 0.880 ;
        RECT 8.760 0.710 8.930 0.880 ;
        RECT 9.490 0.680 9.660 0.850 ;
        RECT -7.810 0.380 -7.630 0.550 ;
      LAYER met1 ;
        RECT -9.680 5.360 -9.520 6.010 ;
        RECT -9.680 4.810 -9.410 5.360 ;
        RECT -9.690 4.760 -9.410 4.810 ;
        RECT -9.270 5.020 -9.080 6.010 ;
        RECT -8.870 5.330 -8.710 6.010 ;
        RECT -7.860 5.330 -7.560 5.710 ;
        RECT -8.910 5.310 -8.710 5.330 ;
        RECT -8.920 5.070 -8.690 5.310 ;
        RECT -9.270 4.900 -9.100 5.020 ;
        RECT -9.690 4.670 -9.520 4.760 ;
        RECT -9.680 4.310 -9.520 4.670 ;
        RECT -9.690 4.220 -9.520 4.310 ;
        RECT -9.690 4.170 -9.410 4.220 ;
        RECT -9.680 3.620 -9.410 4.170 ;
        RECT -9.270 4.080 -9.110 4.900 ;
        RECT -8.910 4.850 -8.710 5.070 ;
        RECT -8.870 4.130 -8.710 4.850 ;
        RECT -7.870 4.710 -7.570 5.080 ;
        RECT -9.270 3.960 -9.100 4.080 ;
        RECT -9.680 2.350 -9.520 3.620 ;
        RECT -9.270 3.100 -9.080 3.960 ;
        RECT -8.910 3.910 -8.710 4.130 ;
        RECT -8.920 3.670 -8.690 3.910 ;
        RECT -7.870 3.900 -7.570 4.270 ;
        RECT -4.750 4.090 -4.370 6.010 ;
        RECT -8.910 3.650 -8.710 3.670 ;
        RECT -9.300 2.870 -9.060 3.100 ;
        RECT -9.680 1.800 -9.410 2.350 ;
        RECT -9.690 1.750 -9.410 1.800 ;
        RECT -9.270 2.010 -9.080 2.870 ;
        RECT -8.870 2.320 -8.710 3.650 ;
        RECT -7.860 3.270 -7.560 3.650 ;
        RECT -7.860 2.320 -7.560 2.700 ;
        RECT -8.910 2.300 -8.710 2.320 ;
        RECT -8.920 2.060 -8.690 2.300 ;
        RECT -4.750 2.230 -4.360 4.090 ;
        RECT -9.270 1.890 -9.100 2.010 ;
        RECT -9.690 1.660 -9.520 1.750 ;
        RECT -9.680 1.310 -9.520 1.660 ;
        RECT -9.690 1.220 -9.520 1.310 ;
        RECT -9.690 1.170 -9.410 1.220 ;
        RECT -9.680 0.620 -9.410 1.170 ;
        RECT -9.270 1.080 -9.110 1.890 ;
        RECT -8.910 1.840 -8.710 2.060 ;
        RECT -8.870 1.130 -8.710 1.840 ;
        RECT -7.870 1.700 -7.570 2.070 ;
        RECT -9.270 0.960 -9.100 1.080 ;
        RECT -9.680 -0.030 -9.520 0.620 ;
        RECT -9.270 -0.030 -9.080 0.960 ;
        RECT -8.910 0.910 -8.710 1.130 ;
        RECT -8.920 0.670 -8.690 0.910 ;
        RECT -7.870 0.900 -7.570 1.270 ;
        RECT -8.910 0.650 -8.710 0.670 ;
        RECT -8.870 -0.030 -8.710 0.650 ;
        RECT -7.860 0.270 -7.560 0.650 ;
        RECT -4.750 -0.030 -4.370 2.230 ;
        RECT -0.720 -0.040 -0.320 5.950 ;
        RECT 0.360 -0.040 0.760 5.950 ;
        RECT 4.410 4.090 4.790 6.010 ;
        RECT 7.600 5.330 7.900 5.710 ;
        RECT 8.750 5.330 8.910 6.010 ;
        RECT 8.750 5.310 8.950 5.330 ;
        RECT 7.610 4.710 7.910 5.080 ;
        RECT 8.730 5.070 8.960 5.310 ;
        RECT 8.750 4.850 8.950 5.070 ;
        RECT 9.120 5.020 9.310 6.010 ;
        RECT 9.560 5.360 9.720 6.010 ;
        RECT 9.140 4.900 9.310 5.020 ;
        RECT 4.400 2.230 4.790 4.090 ;
        RECT 7.610 3.900 7.910 4.270 ;
        RECT 8.750 4.130 8.910 4.850 ;
        RECT 8.750 3.910 8.950 4.130 ;
        RECT 9.150 4.080 9.310 4.900 ;
        RECT 9.450 4.810 9.720 5.360 ;
        RECT 9.450 4.760 9.730 4.810 ;
        RECT 9.560 4.670 9.730 4.760 ;
        RECT 9.560 4.310 9.720 4.670 ;
        RECT 9.560 4.220 9.730 4.310 ;
        RECT 9.140 3.960 9.310 4.080 ;
        RECT 8.730 3.670 8.960 3.910 ;
        RECT 8.750 3.650 8.950 3.670 ;
        RECT 7.600 3.270 7.900 3.650 ;
        RECT 7.600 2.320 7.900 2.700 ;
        RECT 8.750 2.320 8.910 3.650 ;
        RECT 9.120 3.100 9.310 3.960 ;
        RECT 9.450 4.170 9.730 4.220 ;
        RECT 9.450 3.620 9.720 4.170 ;
        RECT 9.100 2.870 9.340 3.100 ;
        RECT 8.750 2.300 8.950 2.320 ;
        RECT 4.410 -0.030 4.790 2.230 ;
        RECT 7.610 1.700 7.910 2.070 ;
        RECT 8.730 2.060 8.960 2.300 ;
        RECT 8.750 1.840 8.950 2.060 ;
        RECT 9.120 2.010 9.310 2.870 ;
        RECT 9.560 2.350 9.720 3.620 ;
        RECT 9.140 1.890 9.310 2.010 ;
        RECT 7.610 0.900 7.910 1.270 ;
        RECT 8.750 1.130 8.910 1.840 ;
        RECT 8.750 0.910 8.950 1.130 ;
        RECT 9.150 1.080 9.310 1.890 ;
        RECT 9.450 1.800 9.720 2.350 ;
        RECT 9.450 1.750 9.730 1.800 ;
        RECT 9.560 1.660 9.730 1.750 ;
        RECT 9.560 1.310 9.720 1.660 ;
        RECT 9.560 1.220 9.730 1.310 ;
        RECT 9.140 0.960 9.310 1.080 ;
        RECT 8.730 0.670 8.960 0.910 ;
        RECT 8.750 0.650 8.950 0.670 ;
        RECT 7.600 0.270 7.900 0.650 ;
        RECT 8.750 -0.030 8.910 0.650 ;
        RECT 9.120 -0.030 9.310 0.960 ;
        RECT 9.450 1.170 9.730 1.220 ;
        RECT 9.450 0.620 9.720 1.170 ;
        RECT 9.560 -0.030 9.720 0.620 ;
      LAYER via ;
        RECT -7.840 5.390 -7.580 5.660 ;
        RECT -7.870 4.740 -7.570 5.050 ;
        RECT -7.870 3.930 -7.570 4.240 ;
        RECT -7.840 3.320 -7.580 3.590 ;
        RECT -7.840 2.380 -7.580 2.650 ;
        RECT -7.870 1.730 -7.570 2.040 ;
        RECT -7.870 0.930 -7.570 1.240 ;
        RECT -7.840 0.320 -7.580 0.590 ;
        RECT 7.620 5.390 7.880 5.660 ;
        RECT 7.610 4.740 7.910 5.050 ;
        RECT 7.610 3.930 7.910 4.240 ;
        RECT 7.620 3.320 7.880 3.590 ;
        RECT 7.620 2.380 7.880 2.650 ;
        RECT 7.610 1.730 7.910 2.040 ;
        RECT 7.610 0.930 7.910 1.240 ;
        RECT 7.620 0.320 7.880 0.590 ;
      LAYER met2 ;
        RECT -7.860 5.510 -7.560 5.710 ;
        RECT 7.600 5.510 7.900 5.710 ;
        RECT -10.040 5.330 10.080 5.510 ;
        RECT -10.040 4.900 10.080 5.080 ;
        RECT -7.870 4.710 -7.570 4.900 ;
        RECT 7.610 4.710 7.910 4.900 ;
        RECT -7.870 4.080 -7.570 4.270 ;
        RECT 7.610 4.080 7.910 4.270 ;
        RECT -10.040 3.900 10.080 4.080 ;
        RECT -10.040 3.470 10.080 3.650 ;
        RECT -7.860 3.270 -7.560 3.470 ;
        RECT 7.600 3.270 7.900 3.470 ;
        RECT -7.860 2.500 -7.560 2.700 ;
        RECT 7.600 2.500 7.900 2.700 ;
        RECT -10.040 2.490 -7.480 2.500 ;
        RECT 7.520 2.490 10.080 2.500 ;
        RECT -10.040 2.320 10.080 2.490 ;
        RECT -10.040 1.900 10.080 2.070 ;
        RECT -10.040 1.890 -7.480 1.900 ;
        RECT 7.520 1.890 10.080 1.900 ;
        RECT -7.870 1.700 -7.570 1.890 ;
        RECT 7.610 1.700 7.910 1.890 ;
        RECT -7.870 1.090 -7.570 1.270 ;
        RECT 7.610 1.090 7.910 1.270 ;
        RECT -7.870 1.080 7.910 1.090 ;
        RECT -10.040 0.920 10.080 1.080 ;
        RECT -10.040 0.900 -7.480 0.920 ;
        RECT -2.300 0.830 -0.760 0.920 ;
        RECT 0.800 0.830 2.340 0.920 ;
        RECT 7.520 0.900 10.080 0.920 ;
        RECT -10.040 0.480 10.080 0.650 ;
        RECT -10.040 0.470 -7.480 0.480 ;
        RECT 7.520 0.470 10.080 0.480 ;
        RECT -7.860 0.270 -7.560 0.470 ;
        RECT 7.600 0.270 7.900 0.470 ;
  END
END swc4x2cell
END LIBRARY

