magic
tech sky130A
timestamp 1628616986
<< checkpaint >>
rect -630 1246 1925 1390
rect -630 -336 2262 1246
rect -294 -480 2262 -336
rect -23 -486 2262 -480
rect 314 -630 2262 -486
<< error_s >>
rect 307 684 308 687
rect 307 533 308 536
rect 307 382 308 385
rect 839 315 891 316
rect 1049 315 1099 316
<< nwell >>
rect 669 749 691 755
rect 669 154 691 159
<< metal1 >>
rect 61 748 83 756
rect 318 747 341 756
rect 367 721 394 750
rect 669 749 691 755
rect 1166 751 1193 756
rect 363 694 366 721
rect 393 694 396 721
rect 459 702 486 707
rect 367 616 394 694
rect 366 613 394 616
rect 393 586 394 613
rect 366 583 394 586
rect 367 580 394 583
rect 413 653 440 660
rect 413 448 440 626
rect 459 561 486 675
rect 554 657 583 662
rect 552 654 583 657
rect 581 625 583 654
rect 552 622 583 625
rect 454 534 457 561
rect 484 534 487 561
rect 412 445 440 448
rect 439 418 440 445
rect 412 415 440 418
rect 413 298 440 415
rect 459 403 486 534
rect 457 400 486 403
rect 484 373 486 400
rect 457 370 486 373
rect 459 368 486 370
rect 506 507 533 513
rect 506 504 534 507
rect 506 477 507 504
rect 506 474 534 477
rect 554 500 583 622
rect 554 474 556 500
rect 582 474 583 500
rect 413 295 443 298
rect 413 268 416 295
rect 413 265 443 268
rect 413 260 440 265
rect 506 253 533 474
rect 504 250 533 253
rect 531 223 533 250
rect 504 220 533 223
rect 506 217 533 220
rect 554 357 583 474
rect 554 354 584 357
rect 554 325 555 354
rect 554 322 584 325
rect 554 200 583 322
rect 554 168 583 171
rect 669 154 691 159
rect 1166 154 1193 159
<< via1 >>
rect 366 694 393 721
rect 459 675 486 702
rect 366 586 393 613
rect 413 626 440 653
rect 552 625 581 654
rect 457 534 484 561
rect 412 418 439 445
rect 457 373 484 400
rect 507 477 534 504
rect 556 474 582 500
rect 416 268 443 295
rect 504 223 531 250
rect 555 325 584 354
rect 554 171 583 200
<< metal2 >>
rect 371 740 608 741
rect 369 725 608 740
rect 369 724 396 725
rect 366 721 396 724
rect 0 699 11 717
rect 343 699 366 717
rect 393 699 396 721
rect 366 691 393 694
rect 456 675 459 702
rect 486 696 489 702
rect 486 680 608 696
rect 486 675 489 680
rect 410 650 413 653
rect 343 632 413 650
rect 410 626 413 632
rect 440 650 443 653
rect 440 631 445 650
rect 440 626 443 631
rect 549 625 552 654
rect 581 647 584 654
rect 581 631 608 647
rect 581 625 584 631
rect 1282 627 1295 644
rect 363 586 366 613
rect 393 607 396 613
rect 393 591 527 607
rect 393 586 396 591
rect 511 590 527 591
rect 511 574 607 590
rect 0 548 11 566
rect 343 564 479 566
rect 343 561 484 564
rect 343 548 457 561
rect 484 534 485 545
rect 457 531 485 534
rect 462 529 485 531
rect 512 529 608 545
rect 512 504 528 529
rect 504 499 507 504
rect 343 481 507 499
rect 504 477 507 481
rect 534 477 537 504
rect 553 474 556 500
rect 582 496 585 500
rect 582 480 608 496
rect 582 474 585 480
rect 1282 476 1295 493
rect 409 418 412 445
rect 439 439 442 445
rect 439 423 608 439
rect 439 418 442 423
rect 0 397 11 415
rect 454 373 457 400
rect 484 394 487 400
rect 484 378 608 394
rect 484 373 487 378
rect 552 348 555 354
rect 343 330 555 348
rect 552 325 555 330
rect 584 348 587 354
rect 584 345 601 348
rect 584 329 608 345
rect 584 325 587 329
rect 1282 325 1295 342
rect 413 268 416 295
rect 443 289 446 295
rect 443 273 608 289
rect 443 268 446 273
rect 501 223 504 250
rect 531 244 534 250
rect 531 228 608 244
rect 531 223 534 228
rect 551 171 554 200
rect 583 195 586 200
rect 583 179 608 195
rect 583 171 586 179
rect 1282 175 1295 192
use sky130_hilas_VinjInv2  VinjInv2_0
timestamp 1628616709
transform 1 0 336 0 1 452
box 0 0 361 164
use sky130_hilas_VinjInv2  VinjInv2_1
timestamp 1628616709
transform 1 0 336 0 1 301
box 0 0 361 164
use sky130_hilas_VinjInv2  VinjInv2_2
timestamp 1628616709
transform 1 0 336 0 1 150
box 0 0 361 164
use sky130_hilas_VinjNOR3  VinjNOR3_2
timestamp 1628616728
transform 1 0 944 0 1 301
box 0 0 688 164
use sky130_hilas_VinjNOR3  VinjNOR3_1
timestamp 1628616728
transform 1 0 944 0 1 150
box 0 0 688 164
use sky130_hilas_VinjNOR3  VinjNOR3_3
timestamp 1628616728
transform 1 0 944 0 1 452
box 0 0 688 164
use sky130_hilas_VinjNOR3  VinjNOR3_0
timestamp 1628616728
transform 1 0 944 0 1 0
box 0 0 688 164
<< labels >>
rlabel metal2 1282 627 1295 644 0 OUTPUT00
port 1 nsew
rlabel metal2 1282 476 1295 493 0 OUTPUT01
port 2 nsew
rlabel metal2 1282 325 1295 342 0 OUTPUT10
port 3 nsew
rlabel metal2 1282 175 1295 192 0 OUTPUT11
port 4 nsew
rlabel metal1 1166 751 1193 756 0 VGND
port 5 nsew
rlabel metal1 1166 154 1193 159 0 VGND
port 5 nsew
rlabel metal1 669 154 691 159 0 VINJ
port 6 nsew
rlabel metal1 669 749 691 755 0 VINJ
port 6 nsew
rlabel metal2 0 699 11 717 0 IN1
port 8 nsew
rlabel metal2 0 548 11 566 0 IN2
port 7 nsew
rlabel metal2 0 397 11 415 0 ENABLE
port 9 nsew
rlabel metal1 61 748 83 756 0 VINJ
port 6 nsew
rlabel metal1 318 747 341 756 0 VGND
port 5 nsew
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
