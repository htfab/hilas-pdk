magic
tech sky130A
timestamp 1628704444
<< checkpaint >>
rect -396 827 897 917
rect -475 -394 897 827
rect -475 -484 818 -394
<< error_s >>
rect 62 542 101 545
rect 62 500 101 503
rect 61 446 100 449
rect 61 404 100 407
rect 61 350 100 353
rect 61 308 100 311
rect 61 254 100 257
rect 61 212 100 215
rect 61 158 100 161
rect 61 116 100 119
rect 62 62 101 65
rect 62 20 101 23
use sky130_hilas_pFETdevice01b  sky130_hilas_pFETdevice01b_1
timestamp 1628704389
transform 1 0 79 0 1 234
box 0 0 188 133
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_0
timestamp 1628704441
transform 1 0 79 0 1 138
box 0 0 161 121
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_3
timestamp 1628704441
transform 1 0 79 0 1 330
box 0 0 161 121
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_6
timestamp 1628704441
transform 1 0 79 0 1 426
box 0 0 161 121
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_0
timestamp 1628704221
transform 1 0 80 0 1 522
box 0 0 172 121
use sky130_hilas_pFETdevice01a  sky130_hilas_pFETdevice01a_0
timestamp 1628704413
transform 1 0 80 0 1 42
box 0 0 161 85
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
