magic
tech sky130A
timestamp 1628616964
<< error_p >>
rect 0 668 85 701
rect 597 603 603 609
rect 646 603 652 609
rect 73 577 79 583
rect 125 577 131 583
rect 67 519 73 525
rect 131 519 137 525
rect 73 467 79 473
rect 125 467 131 473
rect 591 419 597 425
rect 652 419 658 425
rect 661 419 697 420
rect 67 410 73 416
rect 131 410 137 416
rect 593 391 594 395
rect 593 370 599 376
rect 646 370 652 376
rect 73 359 79 365
rect 125 359 131 365
rect 66 309 73 315
rect 131 309 137 315
rect 587 295 593 301
rect 652 295 658 301
rect 932 267 953 268
rect 72 259 78 265
rect 125 259 131 265
rect 66 209 72 215
rect 131 209 137 215
rect 566 198 591 219
rect 566 194 597 198
rect 660 194 666 200
rect 566 167 591 194
rect 72 159 78 165
rect 125 159 131 165
rect 66 109 72 115
rect 131 109 137 115
rect 582 80 591 98
rect 600 80 601 81
rect 666 80 672 86
rect 688 80 691 192
rect 550 78 591 80
rect 599 79 691 80
rect 600 78 691 79
rect 575 55 591 78
rect 945 34 975 35
rect 912 1 959 2
rect 1041 0 1043 86
<< nwell >>
rect 0 617 191 668
rect 1 2 191 617
rect 474 468 753 666
rect 472 189 754 468
rect 476 2 754 189
rect 894 2 1041 668
rect 959 0 1041 2
<< mvpmos >>
rect 945 558 975 608
rect 945 421 975 472
rect 945 348 975 400
rect 945 267 975 319
rect 945 196 975 246
rect 945 61 975 111
<< mvvaractor >>
rect 73 519 131 577
rect 73 410 131 467
rect 597 419 652 603
rect 73 309 131 359
rect 593 295 652 370
rect 72 209 131 259
rect 72 109 131 159
rect 591 80 666 194
rect 591 78 600 80
<< mvpdiff >>
rect 945 631 975 635
rect 945 614 951 631
rect 969 614 975 631
rect 945 608 975 614
rect 945 552 975 558
rect 945 535 951 552
rect 969 535 975 552
rect 945 530 975 535
rect 945 495 975 500
rect 945 478 951 495
rect 969 478 975 495
rect 945 472 975 478
rect 945 400 975 421
rect 945 342 975 348
rect 945 325 951 342
rect 969 325 975 342
rect 945 319 975 325
rect 945 246 975 267
rect 945 190 975 196
rect 945 173 951 190
rect 969 173 975 190
rect 945 169 975 173
rect 945 134 975 138
rect 945 117 951 134
rect 969 117 975 134
rect 945 111 975 117
rect 945 55 975 61
rect 945 38 951 55
rect 969 38 975 55
rect 945 34 975 38
<< mvpdiffc >>
rect 951 614 969 631
rect 951 535 969 552
rect 951 478 969 495
rect 951 325 969 342
rect 951 173 969 190
rect 951 117 969 134
rect 951 38 969 55
<< psubdiff >>
rect 810 81 836 93
rect 810 64 814 81
rect 832 64 836 81
rect 810 52 836 64
<< mvnsubdiff >>
rect 73 577 131 624
rect 597 603 652 633
rect 73 467 131 519
rect 73 359 131 410
rect 597 399 652 419
rect 594 391 652 399
rect 593 370 652 391
rect 72 259 131 309
rect 593 252 652 295
rect 72 159 131 209
rect 591 194 666 252
rect 72 82 131 109
rect 72 55 87 82
rect 115 55 131 82
rect 600 78 666 80
rect 72 45 131 55
rect 591 39 666 78
<< psubdiffcont >>
rect 814 64 832 81
<< mvnsubdiffcont >>
rect 87 55 115 82
<< poly >>
rect 551 602 597 603
rect 30 519 73 577
rect 131 519 174 577
rect 549 496 597 602
rect 515 469 597 496
rect 31 410 73 467
rect 131 410 174 467
rect 549 419 597 469
rect 652 496 697 603
rect 911 558 945 608
rect 975 558 988 608
rect 652 469 723 496
rect 911 472 932 558
rect 652 420 697 469
rect 911 421 945 472
rect 975 421 990 472
rect 652 419 661 420
rect 31 309 73 359
rect 131 309 175 359
rect 551 295 593 370
rect 652 295 695 370
rect 931 348 945 400
rect 975 348 1001 400
rect 978 319 1001 348
rect 30 209 72 259
rect 131 209 174 259
rect 932 267 945 319
rect 975 267 1001 319
rect 916 246 932 247
rect 916 196 945 246
rect 975 196 994 246
rect 30 109 72 159
rect 131 109 174 159
rect 539 78 591 192
rect 666 80 688 194
rect 916 111 932 196
rect 916 61 945 111
rect 975 61 991 111
rect 916 60 932 61
<< locali >>
rect 943 614 951 631
rect 969 614 977 631
rect 943 535 951 552
rect 969 535 977 552
rect 943 478 951 495
rect 969 478 977 495
rect 942 325 951 342
rect 969 325 977 342
rect 943 173 951 190
rect 969 173 977 190
rect 943 117 951 134
rect 969 117 977 134
rect 87 82 115 90
rect 806 64 814 81
rect 832 64 840 81
rect 87 47 115 55
rect 943 38 951 55
rect 969 38 977 55
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
