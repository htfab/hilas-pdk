magic
tech sky130A
timestamp 1628704215
use sky130_hilas_nFETmed  sky130_hilas_nFETmed_3
timestamp 1628285143
transform 1 0 232 0 1 44
box -12 -44 70 228
use sky130_hilas_nFETmed  sky130_hilas_nFETmed_4
timestamp 1628285143
transform 1 0 12 0 1 44
box -12 -44 70 228
use sky130_hilas_nFETmed  sky130_hilas_nFETmed_0
timestamp 1628285143
transform 1 0 67 0 1 44
box -12 -44 70 228
use sky130_hilas_nFETmed  sky130_hilas_nFETmed_1
timestamp 1628285143
transform 1 0 122 0 1 44
box -12 -44 70 228
use sky130_hilas_nFETmed  sky130_hilas_nFETmed_2
timestamp 1628285143
transform 1 0 177 0 1 44
box -12 -44 70 228
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
