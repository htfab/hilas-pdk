magic
tech sky130A
timestamp 1628707326
<< checkpaint >>
rect -472 1020 811 1028
rect -482 994 811 1020
rect -529 980 811 994
rect -538 872 811 980
rect -538 830 816 872
rect -588 815 816 830
rect -602 -420 816 815
rect -602 -430 807 -420
rect -602 -478 801 -430
rect -536 -532 801 -478
rect -536 -547 787 -532
rect -536 -615 786 -547
rect -536 -616 772 -615
rect -522 -630 772 -616
<< nwell >>
rect 0 314 186 321
rect 134 285 179 308
<< poly >>
rect 92 350 115 354
rect 94 47 115 48
<< locali >>
rect 146 384 168 393
rect 146 376 154 384
rect 41 262 59 368
rect 114 321 119 334
rect 102 308 119 321
rect 139 102 146 104
rect 139 88 147 102
rect 116 19 123 45
<< metal1 >>
rect 150 189 171 366
<< metal2 >>
rect 92 285 179 308
rect 92 284 135 285
rect 140 205 187 230
rect 122 102 177 127
rect 68 16 156 41
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628707307
transform 1 0 42 0 1 167
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1628707307
transform -1 0 142 0 -1 33
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628707307
transform 1 0 115 0 1 295
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1628707307
transform -1 0 157 0 -1 116
box 0 0 34 33
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1628707321
transform 1 0 154 0 1 210
box 0 0 32 32
use sky130_hilas_poly2li  sky130_hilas_poly2li_1
timestamp 1628707323
transform 1 0 103 0 1 28
box 0 0 27 33
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1628707287
transform 1 0 158 0 1 369
box 0 0 23 29
use sky130_hilas_poly2li  sky130_hilas_poly2li_0
timestamp 1628707323
transform 1 0 101 0 1 331
box 0 0 27 33
use sky130_hilas_pTransistorVert01  sky130_hilas_pTransistorVert01_1
timestamp 1628707271
transform 1 0 363 0 1 459
box 0 0 186 299
use sky130_hilas_pTransistorVert01  sky130_hilas_pTransistorVert01_0
timestamp 1628707271
transform 1 0 363 0 1 764
box 0 0 186 299
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
