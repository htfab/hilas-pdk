magic
tech sky130A
timestamp 1628616673
<< error_p >>
rect 0 669 85 701
rect 73 577 79 583
rect 125 577 131 583
rect 67 519 73 525
rect 131 519 137 525
rect 597 519 603 525
rect 646 519 652 525
rect 694 496 697 519
rect 73 467 79 473
rect 125 467 131 473
rect 591 446 597 452
rect 652 446 658 452
rect 694 446 697 469
rect 1142 458 1168 680
rect 67 410 73 416
rect 131 410 137 416
rect 593 391 594 395
rect 593 370 599 376
rect 646 370 652 376
rect 73 359 79 365
rect 125 359 131 365
rect 66 309 73 315
rect 131 309 137 315
rect 587 295 593 301
rect 652 295 658 301
rect 995 267 1015 275
rect 72 259 78 265
rect 125 259 131 265
rect 66 209 72 215
rect 131 209 137 215
rect 566 198 591 219
rect 566 194 597 198
rect 660 194 666 200
rect 566 167 591 194
rect 72 159 78 165
rect 125 159 131 165
rect 66 109 72 115
rect 131 109 137 115
rect 582 80 591 98
rect 600 80 601 81
rect 666 80 672 86
rect 688 80 691 192
rect 550 78 591 80
rect 599 79 691 80
rect 600 78 691 79
rect 575 55 591 78
rect 945 34 975 35
rect 912 1 959 2
rect 1041 0 1043 86
<< nwell >>
rect 0 617 191 669
rect 1 2 191 617
rect 474 468 753 666
rect 472 189 754 468
rect 476 2 754 189
rect 894 2 1041 668
rect 1142 459 1468 680
rect 1142 458 1464 459
rect 959 0 1041 2
<< mvpmos >>
rect 945 558 975 608
rect 1244 585 1294 615
rect 1244 523 1294 554
rect 1316 523 1366 554
rect 945 421 975 472
rect 945 348 975 400
rect 945 267 975 319
rect 945 196 975 246
rect 945 61 975 111
<< mvvaractor >>
rect 73 519 131 577
rect 73 410 131 467
rect 597 446 652 519
rect 73 309 131 359
rect 593 295 652 370
rect 72 209 131 259
rect 72 109 131 159
rect 591 80 666 194
rect 591 78 600 80
<< mvpdiff >>
rect 945 631 975 635
rect 945 614 951 631
rect 969 614 975 631
rect 945 608 975 614
rect 1210 609 1244 615
rect 1210 592 1219 609
rect 1237 592 1244 609
rect 1210 585 1244 592
rect 1294 608 1325 615
rect 1294 591 1301 608
rect 1320 591 1325 608
rect 1294 585 1325 591
rect 945 552 975 558
rect 945 535 951 552
rect 969 535 975 552
rect 945 530 975 535
rect 1210 547 1244 554
rect 1210 530 1219 547
rect 1237 530 1244 547
rect 1210 523 1244 530
rect 1294 523 1316 554
rect 1366 547 1400 554
rect 1366 530 1373 547
rect 1393 530 1400 547
rect 1366 523 1400 530
rect 945 495 975 500
rect 945 478 951 495
rect 969 478 975 495
rect 945 472 975 478
rect 945 400 975 421
rect 945 342 975 348
rect 945 325 951 342
rect 969 325 975 342
rect 945 319 975 325
rect 945 246 975 267
rect 945 190 975 196
rect 945 173 951 190
rect 969 173 975 190
rect 945 169 975 173
rect 945 134 975 138
rect 945 117 951 134
rect 969 117 975 134
rect 945 111 975 117
rect 945 55 975 61
rect 945 38 951 55
rect 969 38 975 55
rect 945 34 975 38
<< mvpdiffc >>
rect 951 614 969 631
rect 1219 592 1237 609
rect 1301 591 1320 608
rect 951 535 969 552
rect 1219 530 1237 547
rect 1373 530 1393 547
rect 951 478 969 495
rect 951 325 969 342
rect 951 173 969 190
rect 951 117 969 134
rect 951 38 969 55
<< psubdiff >>
rect 810 81 836 93
rect 810 64 814 81
rect 832 64 836 81
rect 810 52 836 64
<< mvnsubdiff >>
rect 73 577 131 624
rect 597 519 652 633
rect 73 467 131 519
rect 1366 625 1399 629
rect 1366 611 1400 625
rect 1366 593 1373 611
rect 1393 593 1400 611
rect 1366 581 1400 593
rect 73 359 131 410
rect 597 399 652 446
rect 594 391 652 399
rect 593 370 652 391
rect 72 259 131 309
rect 593 252 652 295
rect 72 159 131 209
rect 591 194 666 252
rect 72 82 131 109
rect 72 55 87 82
rect 115 55 131 82
rect 600 78 666 80
rect 72 45 131 55
rect 591 39 666 78
<< psubdiffcont >>
rect 814 64 832 81
<< mvnsubdiffcont >>
rect 1373 593 1393 611
rect 87 55 115 82
<< poly >>
rect 30 519 73 577
rect 131 519 174 577
rect 1244 615 1294 629
rect 911 608 932 610
rect 911 558 945 608
rect 975 558 988 608
rect 551 496 597 519
rect 515 469 597 496
rect 31 410 73 467
rect 131 410 174 467
rect 551 446 597 469
rect 652 496 694 519
rect 652 469 723 496
rect 911 472 932 558
rect 1244 554 1294 585
rect 1329 569 1349 629
rect 1316 554 1366 569
rect 1244 508 1294 523
rect 1316 509 1366 523
rect 652 446 694 469
rect 911 421 945 472
rect 975 421 990 472
rect 31 309 73 359
rect 131 309 175 359
rect 551 295 593 370
rect 652 295 695 370
rect 931 348 945 400
rect 975 348 1019 400
rect 995 319 1019 348
rect 30 209 72 259
rect 131 209 174 259
rect 932 267 945 319
rect 975 275 1019 319
rect 975 267 994 275
rect 995 267 1019 275
rect 932 196 945 246
rect 975 196 994 246
rect 30 109 72 159
rect 131 109 174 159
rect 539 78 591 192
rect 666 80 688 194
rect 929 61 945 111
rect 975 61 991 111
<< locali >>
rect 943 614 951 631
rect 969 614 977 631
rect 1210 592 1219 609
rect 1237 592 1245 609
rect 1300 608 1320 617
rect 1300 591 1301 608
rect 1300 583 1320 591
rect 1373 611 1393 622
rect 943 535 951 552
rect 969 535 977 552
rect 1373 547 1393 593
rect 1210 530 1219 547
rect 1237 530 1245 547
rect 1373 522 1393 530
rect 943 478 951 495
rect 969 478 977 495
rect 942 325 951 342
rect 969 325 977 342
rect 943 173 951 190
rect 969 173 977 190
rect 943 117 951 134
rect 969 117 977 134
rect 87 82 115 90
rect 806 64 814 81
rect 832 64 840 81
rect 87 47 115 55
rect 943 38 951 55
rect 969 38 977 55
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
