magic
tech sky130A
timestamp 1632400811
<< error_s >>
rect -509 717 -459 723
rect -437 717 -387 723
rect -509 675 -459 681
rect -437 675 -387 681
rect -1187 462 -1170 464
rect -1187 443 -1170 445
rect -1187 428 -1170 429
rect 77 421 104 427
rect -1187 409 -1170 410
rect 77 379 104 385
rect 77 354 104 360
rect 77 312 104 318
rect 77 271 104 277
rect 77 229 104 235
rect -509 204 -459 210
rect -437 204 -387 210
rect 77 204 104 210
rect -509 162 -459 168
rect -437 162 -387 168
rect 77 162 104 168
<< nwell >>
rect -328 571 -162 593
rect 191 140 319 159
<< locali >>
rect -1190 479 -1144 488
rect -1190 462 -1187 479
rect -1170 462 -1144 479
rect -149 470 -131 493
rect -1190 410 -1144 462
rect -237 435 -131 470
rect -217 418 -211 435
rect -1190 393 -1187 410
rect -1170 393 -1144 410
rect -1190 387 -1144 393
<< viali >>
rect -1187 462 -1170 479
rect -1187 393 -1170 410
<< metal1 >>
rect -1438 738 -1396 745
rect -1068 737 -1045 745
rect -416 737 -397 745
rect -372 737 -344 745
rect 123 731 157 745
rect 190 730 217 745
rect 127 579 153 605
rect 122 532 165 535
rect 122 498 127 532
rect 161 498 165 532
rect 122 496 165 498
rect 127 495 161 496
rect -1194 484 -1156 488
rect -1194 391 -1190 484
rect -1161 391 -1156 484
rect -1194 387 -1156 391
rect 123 140 157 159
rect 190 140 217 161
<< via1 >>
rect 127 498 161 532
rect -1190 479 -1161 484
rect -1190 462 -1187 479
rect -1187 462 -1170 479
rect -1170 462 -1161 479
rect -1190 410 -1161 462
rect -1190 393 -1187 410
rect -1187 393 -1170 410
rect -1170 393 -1161 410
rect -1190 391 -1161 393
<< metal2 >>
rect -1473 677 -1466 695
rect -328 571 -150 593
rect 124 532 164 533
rect 124 524 127 532
rect -1191 505 127 524
rect -1191 487 -1172 505
rect -42 491 -3 505
rect 124 498 127 505
rect 161 498 164 532
rect 124 497 164 498
rect -1193 484 -1158 487
rect -1193 391 -1190 484
rect -1161 391 -1158 484
rect -62 392 35 434
rect 304 392 319 414
rect -1193 388 -1158 391
rect -177 327 0 347
rect -334 278 -318 318
rect -206 246 0 267
rect -1473 192 -1465 207
rect -286 142 -260 167
use sky130_hilas_pTransistorSingle  sky130_hilas_pTransistorSingle_0
timestamp 1632400113
transform 1 0 -323 0 1 580
box 133 -174 320 165
use sky130_hilas_SingleTACore01  sky130_hilas_SingleTACore01_0
timestamp 1632398358
transform 1 0 164 0 1 181
box -172 -26 155 550
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_0
timestamp 1629420194
transform 1 0 -484 0 1 580
box 133 -440 320 165
use sky130_hilas_FGBias2x1cell  sky130_hilas_FGBias2x1cell_0
timestamp 1631881676
transform 1 0 -1077 0 1 522
box -396 -387 757 228
<< labels >>
rlabel metal1 123 140 157 146 0 VGND
port 7 nsew ground default
rlabel metal1 190 140 217 146 0 VPWR
port 8 nsew power default
rlabel metal1 123 740 157 745 0 VGND
port 7 nsew ground default
rlabel metal1 190 740 217 745 0 VPWR
port 8 nsew power default
rlabel metal2 -286 142 -263 167 0 VIN12
port 2 nsew analog default
rlabel metal2 304 392 319 414 0 OUTPUT1
port 5 nsew
rlabel metal1 -416 737 -397 745 0 COLSEL1
port 1 nsew
rlabel metal2 -1473 677 -1466 695 0 DRAIN1
port 9 nsew
rlabel metal2 -1473 192 -1465 207 0 DRAIN2
port 10 nsew
rlabel metal1 -1438 738 -1396 745 0 VTUN
port 11 nsew
rlabel metal1 -1068 737 -1045 745 0 GATE1
port 12 nsew
rlabel metal1 -372 737 -344 745 0 VINJ
port 13 nsew
<< end >>
