magic
tech sky130A
magscale 1 2
timestamp 1632255311
<< error_s >>
rect 4780 77564 4814 78648
rect 4828 77612 4838 77614
rect 4828 77608 4874 77612
rect 4828 77564 4890 77608
rect 4904 77580 4924 77596
rect 4904 77564 4938 77580
rect 4952 77564 5012 77608
rect 5072 77564 5132 77608
rect 4780 77528 5178 77564
rect 4780 77490 4814 77528
rect 4828 77490 4890 77528
rect 4904 77490 4938 77528
rect 4780 77466 4938 77490
rect 4952 77482 5012 77528
rect 5028 77494 5062 77528
rect 5072 77482 5132 77528
rect 4786 77342 4938 77466
rect 4990 77412 5012 77472
rect 4780 77110 4938 77342
rect 4828 77108 4938 77110
rect 4828 76436 4890 77108
rect 4904 76452 4938 77108
rect 5050 77402 5072 77412
rect 5086 77402 5120 77482
rect 5144 77402 5178 77528
rect 5192 77482 5250 77608
rect 5204 77402 5238 77482
rect 5262 77402 5296 78656
rect 5310 77482 5368 77608
rect 5322 77402 5356 77482
rect 5382 77402 5416 78656
rect 5428 77482 5488 77608
rect 5440 77402 5474 77482
rect 5502 77402 5536 78646
rect 5550 77482 5610 77608
rect 5562 77402 5596 77482
rect 5624 77402 5658 78648
rect 5672 77482 5732 77608
rect 5686 77402 5720 77482
rect 5744 77402 5778 78646
rect 5792 77596 5852 77608
rect 5924 77596 5958 79292
rect 5992 77596 6026 79292
rect 5792 77562 10098 77596
rect 5792 77528 5852 77562
rect 5924 77528 5958 77562
rect 5992 77528 6026 77562
rect 5792 77494 10098 77528
rect 5792 77482 5852 77494
rect 5808 77402 5842 77482
rect 5924 77412 5958 77494
rect 5992 77412 6026 77494
rect 5912 77402 6038 77412
rect 5050 77368 6038 77402
rect 5050 77274 5072 77368
rect 5086 77274 5120 77368
rect 5144 77336 5178 77368
rect 5204 77336 5238 77368
rect 5262 77336 5296 77368
rect 5322 77336 5356 77368
rect 5382 77336 5416 77368
rect 5440 77336 5474 77368
rect 5502 77336 5536 77368
rect 5562 77336 5596 77368
rect 5624 77336 5658 77368
rect 5686 77336 5720 77368
rect 5744 77336 5778 77368
rect 5808 77336 5842 77368
rect 5912 77350 6038 77368
rect 5128 77302 7324 77336
rect 5144 77274 5178 77302
rect 5204 77274 5238 77302
rect 5262 77274 5296 77302
rect 5322 77274 5356 77302
rect 5382 77274 5416 77302
rect 5440 77274 5474 77302
rect 5502 77274 5536 77302
rect 5562 77274 5596 77302
rect 5624 77274 5658 77302
rect 5686 77274 5720 77302
rect 5744 77274 5778 77302
rect 5808 77274 5842 77302
rect 5912 77274 6038 77288
rect 5050 77240 6038 77274
rect 33026 77260 33060 77482
rect 33094 77260 33128 77456
rect 33290 77260 35604 77268
rect 35708 77260 35742 77456
rect 35776 77260 35810 77452
rect 36008 77306 36594 77322
rect 36758 77306 36914 77322
rect 35890 77268 35952 77294
rect 36008 77268 36566 77294
rect 36786 77268 36886 77294
rect 35952 77260 36566 77268
rect 36812 77260 36886 77268
rect 5050 77150 5072 77240
rect 5086 77150 5120 77240
rect 5144 77212 5178 77240
rect 5204 77212 5238 77240
rect 5262 77212 5296 77240
rect 5322 77212 5356 77240
rect 5382 77212 5416 77240
rect 5440 77212 5474 77240
rect 5502 77212 5536 77240
rect 5562 77212 5596 77240
rect 5624 77212 5658 77240
rect 5686 77212 5720 77240
rect 5744 77212 5778 77240
rect 5808 77212 5842 77240
rect 5912 77226 6038 77240
rect 25974 77226 36540 77260
rect 36541 77252 36811 77260
rect 36555 77245 36811 77252
rect 33026 77218 33086 77226
rect 33094 77218 33128 77226
rect 33130 77218 33166 77226
rect 33290 77220 33352 77226
rect 33290 77218 33305 77219
rect 33337 77218 33352 77219
rect 35708 77218 35742 77226
rect 35776 77218 35810 77226
rect 35952 77221 36540 77226
rect 35890 77220 36540 77221
rect 36570 77242 36811 77245
rect 35952 77218 35962 77220
rect 36070 77218 36085 77219
rect 36570 77218 36782 77242
rect 32530 77213 36782 77218
rect 5128 77178 7324 77212
rect 32530 77198 36797 77213
rect 36812 77198 36860 77260
rect 32530 77184 36764 77198
rect 36812 77184 36813 77198
rect 36860 77184 36886 77198
rect 5144 77150 5178 77178
rect 5204 77150 5238 77178
rect 5262 77150 5296 77178
rect 5322 77150 5356 77178
rect 5382 77150 5416 77178
rect 5440 77150 5474 77178
rect 5502 77150 5536 77178
rect 5562 77150 5596 77178
rect 5624 77150 5658 77178
rect 5686 77150 5720 77178
rect 5744 77150 5778 77178
rect 5808 77150 5842 77178
rect 33010 77172 33166 77184
rect 5912 77150 6038 77164
rect 33010 77161 33021 77172
rect 5050 77116 6038 77150
rect 5050 77030 5072 77116
rect 5086 77030 5120 77116
rect 5144 77088 5178 77116
rect 5204 77088 5238 77116
rect 5262 77088 5296 77116
rect 5322 77088 5356 77116
rect 5382 77088 5416 77116
rect 5440 77088 5474 77116
rect 5502 77088 5536 77116
rect 5562 77088 5596 77116
rect 5624 77088 5658 77116
rect 5686 77088 5720 77116
rect 5744 77088 5778 77116
rect 5808 77088 5842 77116
rect 5912 77104 6038 77116
rect 33010 77120 33021 77131
rect 33050 77120 33086 77172
rect 33130 77120 33166 77172
rect 33290 77172 33352 77184
rect 33368 77178 35564 77184
rect 33290 77157 33305 77172
rect 33337 77164 33352 77172
rect 35698 77172 35824 77184
rect 33337 77157 35604 77164
rect 35698 77161 35709 77172
rect 35813 77161 35824 77172
rect 35952 77172 36008 77184
rect 35952 77161 35963 77172
rect 35997 77161 36008 77172
rect 36114 77150 38004 77184
rect 33010 77108 33166 77120
rect 33290 77120 33305 77135
rect 35589 77120 35604 77135
rect 33010 77088 33144 77108
rect 5130 77054 7326 77088
rect 33010 77077 33021 77088
rect 33133 77077 33144 77088
rect 33290 77104 35604 77120
rect 35698 77120 35709 77131
rect 35813 77120 35824 77131
rect 33290 77088 33352 77104
rect 33290 77073 33305 77088
rect 33337 77073 33352 77088
rect 35698 77088 35824 77120
rect 35698 77077 35709 77088
rect 35813 77077 35824 77088
rect 35952 77120 35963 77131
rect 35997 77120 36008 77131
rect 36812 77124 36813 77150
rect 36860 77124 36886 77150
rect 35952 77088 36008 77120
rect 35952 77077 35963 77088
rect 35997 77077 36008 77088
rect 36078 77120 36093 77124
rect 36078 77088 36788 77120
rect 36078 77073 36093 77088
rect 36756 77075 36788 77088
rect 36741 77060 36803 77075
rect 36812 77060 36860 77124
rect 5144 77030 5178 77054
rect 5204 77030 5238 77054
rect 5262 77030 5296 77054
rect 5322 77030 5356 77054
rect 5382 77030 5416 77054
rect 5440 77030 5474 77054
rect 5502 77030 5536 77054
rect 5562 77030 5596 77054
rect 5624 77030 5658 77054
rect 5686 77030 5720 77054
rect 5744 77030 5778 77054
rect 5808 77030 5842 77054
rect 5912 77030 6038 77044
rect 5050 76996 6038 77030
rect 5050 76912 5072 76996
rect 5086 76912 5120 76996
rect 5144 76972 5178 76996
rect 5204 76972 5238 76996
rect 5262 76972 5296 76996
rect 5322 76972 5356 76996
rect 5382 76972 5416 76996
rect 5440 76972 5474 76996
rect 5502 76972 5536 76996
rect 5562 76972 5596 76996
rect 5624 76972 5658 76996
rect 5686 76972 5720 76996
rect 5744 76972 5778 76996
rect 5808 76972 5842 76996
rect 5912 76984 6038 76996
rect 5134 76938 7330 76972
rect 5144 76912 5178 76938
rect 5204 76912 5238 76938
rect 5262 76912 5296 76938
rect 5322 76912 5356 76938
rect 5382 76912 5416 76938
rect 5440 76912 5474 76938
rect 5502 76912 5536 76938
rect 5562 76912 5596 76938
rect 5624 76912 5658 76938
rect 5686 76912 5720 76938
rect 5744 76912 5778 76938
rect 5808 76912 5842 76938
rect 5912 76912 6038 76924
rect 5050 76878 6038 76912
rect 5050 76794 5072 76878
rect 5086 76794 5120 76878
rect 5144 76854 5178 76878
rect 5204 76854 5238 76878
rect 5262 76854 5296 76878
rect 5322 76854 5356 76878
rect 5382 76854 5416 76878
rect 5440 76854 5474 76878
rect 5502 76854 5536 76878
rect 5562 76854 5596 76878
rect 5624 76854 5658 76878
rect 5686 76854 5720 76878
rect 5744 76854 5778 76878
rect 5808 76854 5842 76878
rect 5912 76866 6038 76878
rect 5136 76820 7332 76854
rect 5144 76794 5178 76820
rect 5204 76794 5238 76820
rect 5262 76794 5296 76820
rect 5322 76794 5356 76820
rect 5382 76794 5416 76820
rect 5440 76794 5474 76820
rect 5502 76794 5536 76820
rect 5562 76794 5596 76820
rect 5624 76794 5658 76820
rect 5686 76794 5720 76820
rect 5744 76794 5778 76820
rect 5808 76794 5842 76820
rect 5912 76794 6038 76806
rect 5050 76760 6038 76794
rect 5050 76676 5072 76760
rect 5086 76676 5120 76760
rect 5144 76734 5178 76760
rect 5204 76734 5238 76760
rect 5262 76734 5296 76760
rect 5322 76734 5356 76760
rect 5382 76734 5416 76760
rect 5440 76734 5474 76760
rect 5502 76734 5536 76760
rect 5562 76734 5596 76760
rect 5624 76734 5658 76760
rect 5686 76734 5720 76760
rect 5744 76734 5778 76760
rect 5808 76734 5842 76760
rect 5912 76748 6038 76760
rect 5136 76700 7332 76734
rect 5144 76676 5178 76700
rect 5204 76676 5238 76700
rect 5262 76676 5296 76700
rect 5322 76676 5356 76700
rect 5382 76676 5416 76700
rect 5440 76676 5474 76700
rect 5502 76676 5536 76700
rect 5562 76676 5596 76700
rect 5624 76676 5658 76700
rect 5686 76676 5720 76700
rect 5744 76676 5778 76700
rect 5808 76676 5842 76700
rect 5912 76676 6038 76688
rect 5050 76642 6038 76676
rect 5050 76554 5072 76642
rect 5086 76554 5120 76642
rect 5144 76614 5178 76642
rect 5204 76614 5238 76642
rect 5262 76614 5296 76642
rect 5322 76614 5356 76642
rect 5382 76614 5416 76642
rect 5440 76614 5474 76642
rect 5502 76614 5536 76642
rect 5562 76614 5596 76642
rect 5624 76614 5658 76642
rect 5686 76614 5720 76642
rect 5744 76614 5778 76642
rect 5808 76614 5842 76642
rect 5912 76628 6038 76642
rect 5126 76580 7322 76614
rect 5144 76554 5178 76580
rect 5204 76554 5238 76580
rect 5262 76554 5296 76580
rect 5322 76554 5356 76580
rect 5382 76554 5416 76580
rect 5440 76554 5474 76580
rect 5502 76554 5536 76580
rect 5562 76554 5596 76580
rect 5624 76554 5658 76580
rect 5686 76554 5720 76580
rect 5744 76554 5778 76580
rect 5808 76554 5842 76580
rect 5912 76554 6038 76566
rect 5050 76520 6038 76554
rect 5050 76436 5072 76520
rect 4770 76374 4904 76436
rect 5086 76430 5120 76520
rect 5144 76492 5178 76520
rect 5204 76492 5238 76520
rect 5262 76492 5296 76520
rect 5322 76492 5356 76520
rect 5382 76492 5416 76520
rect 5440 76492 5474 76520
rect 5502 76492 5536 76520
rect 5562 76492 5596 76520
rect 5624 76492 5658 76520
rect 5686 76492 5720 76520
rect 5744 76492 5778 76520
rect 5808 76492 5842 76520
rect 5912 76506 6038 76520
rect 5128 76458 7324 76492
rect 5204 76430 5238 76458
rect 5322 76430 5356 76458
rect 5440 76430 5474 76458
rect 5502 76450 5536 76458
rect 5562 76430 5596 76458
rect 5624 76452 5658 76458
rect 5686 76430 5720 76458
rect 5744 76450 5778 76458
rect 5808 76430 5842 76458
rect 5912 76430 6038 76444
rect 5064 76396 6038 76430
rect 5086 76386 5120 76396
rect 5204 76386 5238 76396
rect 5322 76386 5356 76396
rect 5440 76386 5474 76396
rect 5562 76386 5596 76396
rect 5686 76388 5720 76396
rect 5808 76386 5842 76396
rect 5912 76384 6038 76396
rect 4988 76374 5050 76384
rect 5112 76374 5852 76384
rect 4786 76212 4820 76374
rect 5792 76372 5852 76374
rect 5912 76288 6038 76324
rect 5912 76284 6064 76288
rect 5054 76266 6158 76284
rect 5912 76264 6038 76266
rect 4854 76238 4888 76246
rect 6026 76240 6030 76254
rect 4660 76192 5878 76212
rect 4660 76178 10120 76192
rect 4918 76158 10120 76178
rect 4634 76124 5910 76144
rect 4634 76110 10120 76124
rect 4918 76090 10120 76110
rect 25898 75826 25902 77044
rect 33010 77036 33021 77047
rect 33133 77036 33144 77047
rect 33010 77004 33144 77036
rect 33010 76993 33021 77004
rect 33133 76993 33144 77004
rect 33290 77036 33305 77051
rect 35589 77036 35604 77044
rect 33290 77004 35604 77036
rect 33290 76989 33305 77004
rect 35589 76989 35604 77004
rect 35698 77036 35709 77047
rect 35813 77036 35824 77047
rect 35698 77004 35824 77036
rect 35698 76993 35709 77004
rect 35813 76993 35824 77004
rect 35952 77036 35963 77047
rect 35997 77036 36008 77047
rect 35952 77004 36008 77036
rect 35952 76993 35963 77004
rect 35997 76993 36008 77004
rect 33010 76958 33021 76969
rect 33133 76958 33144 76969
rect 33010 76926 33144 76958
rect 33010 76915 33021 76926
rect 33133 76915 33144 76926
rect 33290 76958 33305 76973
rect 33337 76958 33352 76973
rect 35952 76969 35962 76993
rect 36812 76976 36813 77060
rect 36860 76976 36886 77060
rect 33290 76926 33352 76958
rect 33290 76912 33305 76926
rect 33337 76924 33352 76926
rect 35698 76958 35709 76969
rect 35813 76958 35824 76969
rect 35698 76926 35824 76958
rect 33290 76911 33302 76912
rect 33337 76911 35604 76924
rect 35698 76915 35709 76926
rect 35813 76915 35824 76926
rect 35952 76958 35963 76969
rect 35997 76958 36008 76969
rect 35952 76926 36008 76958
rect 35952 76915 35963 76926
rect 35997 76915 36008 76926
rect 36088 76958 36103 76973
rect 36088 76927 36788 76958
rect 36088 76926 36803 76927
rect 33010 76876 33021 76887
rect 33133 76876 33144 76887
rect 33010 76844 33144 76876
rect 33010 76833 33021 76844
rect 33133 76833 33144 76844
rect 33290 76876 33305 76891
rect 35589 76876 35604 76891
rect 35952 76887 35962 76915
rect 36088 76912 36103 76926
rect 36741 76912 36803 76926
rect 36812 76912 36860 76976
rect 33290 76866 35604 76876
rect 35698 76876 35709 76887
rect 35813 76876 35824 76887
rect 33290 76844 33352 76866
rect 33290 76829 33305 76844
rect 33337 76829 33352 76844
rect 35698 76844 35824 76876
rect 35698 76833 35709 76844
rect 35813 76833 35824 76844
rect 35952 76876 35963 76887
rect 35997 76876 36008 76887
rect 35952 76844 36008 76876
rect 35952 76833 35963 76844
rect 35997 76833 36008 76844
rect 36812 76838 36813 76912
rect 36860 76838 36886 76912
rect 33010 76800 33021 76811
rect 33133 76800 33144 76811
rect 33010 76768 33144 76800
rect 33010 76757 33021 76768
rect 33133 76757 33144 76768
rect 33290 76800 33305 76815
rect 35952 76811 35962 76833
rect 36088 76829 36803 76838
rect 35589 76800 35604 76806
rect 33290 76768 35604 76800
rect 33290 76753 33305 76768
rect 35589 76753 35604 76768
rect 35698 76800 35709 76811
rect 35813 76800 35824 76811
rect 35698 76768 35824 76800
rect 35698 76757 35709 76768
rect 35813 76757 35824 76768
rect 35952 76800 35963 76811
rect 35997 76800 36008 76811
rect 35952 76768 36008 76800
rect 36088 76800 36103 76815
rect 36088 76789 36788 76800
rect 36088 76774 36803 76789
rect 36812 76774 36860 76838
rect 35952 76757 35963 76768
rect 35997 76757 36008 76768
rect 33010 76722 33021 76733
rect 33133 76722 33144 76733
rect 33010 76690 33144 76722
rect 33010 76679 33021 76690
rect 33133 76679 33144 76690
rect 33290 76722 33305 76737
rect 33337 76722 33352 76737
rect 35952 76733 35962 76757
rect 33290 76690 33352 76722
rect 33290 76676 33305 76690
rect 33337 76688 33352 76690
rect 35698 76722 35709 76733
rect 35813 76722 35824 76733
rect 35698 76690 35824 76722
rect 33290 76675 33302 76676
rect 33337 76675 35604 76688
rect 35698 76679 35709 76690
rect 35813 76679 35824 76690
rect 35952 76722 35963 76733
rect 35997 76722 36008 76733
rect 35952 76690 36008 76722
rect 36812 76708 36813 76774
rect 36860 76708 36886 76774
rect 35952 76679 35963 76690
rect 35997 76679 36008 76690
rect 36080 76693 36803 76708
rect 36080 76690 36788 76693
rect 33010 76642 33021 76653
rect 33133 76642 33144 76653
rect 33010 76610 33144 76642
rect 33010 76599 33021 76610
rect 33133 76599 33144 76610
rect 33290 76642 33305 76657
rect 35589 76642 35604 76657
rect 35952 76653 35962 76679
rect 36080 76675 36095 76690
rect 33290 76628 35604 76642
rect 33290 76610 33352 76628
rect 35542 76626 35604 76628
rect 35698 76642 35709 76653
rect 35813 76642 35824 76653
rect 33290 76595 33305 76610
rect 33337 76595 33352 76610
rect 35698 76610 35824 76642
rect 35698 76599 35709 76610
rect 35813 76599 35824 76610
rect 35952 76642 35963 76653
rect 35997 76642 36008 76653
rect 36080 76642 36803 76657
rect 36812 76642 36860 76708
rect 35952 76610 36008 76642
rect 35952 76599 35963 76610
rect 35997 76599 36008 76610
rect 33010 76566 33021 76577
rect 33133 76566 33144 76577
rect 33010 76534 33144 76566
rect 33010 76523 33021 76534
rect 33133 76523 33144 76534
rect 33290 76566 33305 76581
rect 35952 76577 35962 76599
rect 36812 76580 36813 76642
rect 36860 76580 36886 76642
rect 35698 76566 35709 76577
rect 35813 76566 35824 76577
rect 33290 76534 35604 76566
rect 33290 76519 33305 76534
rect 35589 76519 35604 76534
rect 35698 76534 35824 76566
rect 35698 76523 35709 76534
rect 35813 76523 35824 76534
rect 35952 76566 35963 76577
rect 35997 76566 36008 76577
rect 35952 76534 36008 76566
rect 35952 76523 35963 76534
rect 35997 76523 36008 76534
rect 36080 76566 36095 76580
rect 36741 76566 36803 76580
rect 36080 76565 36803 76566
rect 36080 76534 36788 76565
rect 36080 76519 36095 76534
rect 36812 76514 36860 76580
rect 33010 76482 33021 76493
rect 33133 76482 33144 76493
rect 33010 76450 33144 76482
rect 33010 76439 33021 76450
rect 33133 76439 33144 76450
rect 33290 76482 33305 76497
rect 33337 76482 33352 76497
rect 33290 76450 33352 76482
rect 33290 76435 33305 76450
rect 33337 76444 33352 76450
rect 35698 76482 35709 76493
rect 35813 76482 35824 76493
rect 35698 76450 35824 76482
rect 33337 76435 35604 76444
rect 35698 76439 35709 76450
rect 35813 76439 35824 76450
rect 35952 76482 35963 76493
rect 35997 76482 36008 76493
rect 35952 76450 36008 76482
rect 36812 76454 36813 76514
rect 36860 76454 36886 76514
rect 35952 76439 35963 76450
rect 35997 76439 36008 76450
rect 36080 76450 36803 76454
rect 33010 76400 33021 76411
rect 33133 76400 33144 76411
rect 33010 76368 33144 76400
rect 33010 76357 33021 76368
rect 33133 76357 33144 76368
rect 33290 76400 33305 76415
rect 35589 76400 35604 76415
rect 35952 76411 35962 76439
rect 36080 76435 36095 76450
rect 36756 76439 36803 76450
rect 33290 76384 35604 76400
rect 35698 76400 35709 76411
rect 35813 76400 35824 76411
rect 33290 76368 33352 76384
rect 33290 76353 33305 76368
rect 33337 76353 33352 76368
rect 35698 76368 35824 76400
rect 35698 76357 35709 76368
rect 35813 76357 35824 76368
rect 35952 76400 35963 76411
rect 35997 76400 36008 76411
rect 35952 76368 36008 76400
rect 36080 76400 36095 76415
rect 36756 76407 36788 76439
rect 36756 76400 36803 76407
rect 36080 76392 36803 76400
rect 36812 76392 36860 76454
rect 35952 76357 35963 76368
rect 35997 76357 36008 76368
rect 33010 76326 33021 76337
rect 33133 76326 33144 76337
rect 33010 76294 33144 76326
rect 33290 76326 33305 76341
rect 33337 76326 33352 76341
rect 36812 76338 36820 76392
rect 36860 76338 36886 76392
rect 33290 76324 33352 76326
rect 33606 76324 34300 76330
rect 35698 76326 35709 76337
rect 35813 76326 35824 76337
rect 33010 76283 33021 76294
rect 33133 76283 33144 76294
rect 33288 76294 35604 76324
rect 33288 76279 33303 76294
rect 33634 76266 34272 76294
rect 35589 76279 35604 76294
rect 35698 76294 35824 76326
rect 35698 76283 35709 76294
rect 35813 76283 35824 76294
rect 35940 76326 35951 76337
rect 35940 76294 36788 76326
rect 35940 76283 35951 76294
rect 36756 76293 36788 76294
rect 36745 76282 36799 76293
rect 36812 76282 36860 76338
rect 39324 76322 40018 76328
rect 45038 76322 45732 76334
rect 33288 76264 35604 76265
rect 33010 76250 33021 76261
rect 33133 76250 33144 76261
rect 33010 76218 33144 76250
rect 33010 76207 33021 76218
rect 33133 76207 33144 76218
rect 35698 76250 35709 76261
rect 35813 76250 35824 76261
rect 35698 76218 35824 76250
rect 36812 76240 36813 76282
rect 35698 76207 35709 76218
rect 35813 76212 35824 76218
rect 35813 76207 36799 76212
rect 36820 76192 36854 76282
rect 36860 76240 36886 76282
rect 39352 76266 39990 76300
rect 45066 76266 45704 76306
rect 33010 76174 33021 76185
rect 33158 76174 38360 76192
rect 33010 76158 38360 76174
rect 33010 76142 36788 76158
rect 33010 76131 33021 76142
rect 36756 76124 36788 76142
rect 36820 76124 36854 76158
rect 33010 76102 33023 76107
rect 33012 76096 33023 76102
rect 33158 76096 38360 76124
rect 33012 76090 38360 76096
rect 33012 76085 36788 76090
rect 33012 76078 36799 76085
rect 33012 76070 33144 76078
rect 35476 76074 36799 76078
rect 33012 76068 33114 76070
rect 26504 76010 26868 76020
rect 26380 75988 26868 76010
rect 27544 76000 27808 76010
rect 27422 75988 27808 76000
rect 26504 75977 26515 75988
rect 26857 75977 26868 75988
rect 27544 75977 27555 75988
rect 27797 75977 27808 75988
rect 26824 75944 26835 75955
rect 26857 75944 26868 75955
rect 26824 75912 26868 75944
rect 26824 75904 26835 75912
rect 26857 75904 26868 75912
rect 26504 75838 26726 75868
rect 26824 75838 26868 75904
rect 27764 75944 27775 75955
rect 27797 75944 27808 75955
rect 27764 75912 27808 75944
rect 27764 75901 27775 75912
rect 27797 75901 27808 75912
rect 27764 75894 27772 75901
rect 27544 75838 27666 75858
rect 26504 75827 26515 75838
rect 26715 75827 26726 75838
rect 27544 75827 27555 75838
rect 27655 75827 27666 75838
rect 27764 75828 27808 75894
rect 36820 75798 36854 76090
rect 34012 75514 34038 75798
rect 34012 75430 34048 75514
rect 33954 75418 34048 75430
rect 26382 75364 26422 75396
rect 26504 75392 26515 75403
rect 26726 75392 26824 75418
rect 26857 75396 26868 75403
rect 26857 75392 26914 75396
rect 26504 75384 26914 75392
rect 26504 75370 26726 75384
rect 26824 75364 26914 75384
rect 23894 75276 23932 75310
rect 23882 75262 23932 75276
rect 23936 75240 23970 75268
rect 24046 75256 24062 75308
rect 24074 75240 24090 75288
rect 24178 75278 24212 75310
rect 26382 75296 26383 75297
rect 26504 75296 26726 75364
rect 26824 75296 26868 75364
rect 26913 75296 26914 75297
rect 24158 75268 24212 75278
rect 24158 75262 24250 75268
rect 23914 75234 23966 75240
rect 24212 75238 24250 75262
rect 26282 75238 26316 75296
rect 26381 75295 26440 75296
rect 26382 75280 26440 75295
rect 26382 75252 26400 75280
rect 26422 75270 26440 75280
rect 26504 75270 26756 75296
rect 26824 75295 26915 75296
rect 26824 75280 26914 75295
rect 26504 75252 26726 75270
rect 26824 75252 26868 75280
rect 26894 75252 26914 75280
rect 26382 75239 26440 75252
rect 26504 75239 26756 75252
rect 26824 75240 26914 75252
rect 26868 75239 26914 75240
rect 26381 75238 26441 75239
rect 26504 75238 26757 75239
rect 26855 75238 26856 75239
rect 26868 75238 26915 75239
rect 26978 75238 27014 75296
rect 24194 75236 24250 75238
rect 26382 75237 26383 75238
rect 26439 75237 26440 75238
rect 23914 75228 23956 75234
rect 24194 75228 24236 75236
rect 26504 75220 26726 75238
rect 26755 75237 26756 75238
rect 26856 75237 26857 75238
rect 26913 75237 26914 75238
rect 26504 75182 26868 75220
rect 24438 75108 24462 75176
rect 26504 75168 26726 75182
rect 26824 75168 26868 75182
rect 26382 75138 26440 75168
rect 26726 75138 26756 75168
rect 26824 75140 26914 75168
rect 27036 75158 27048 75412
rect 34068 75402 34076 75542
rect 33932 75390 34076 75402
rect 39730 75400 39752 75796
rect 26824 75129 26835 75140
rect 26856 75138 26914 75140
rect 26857 75129 26868 75138
rect 24506 75108 24558 75110
rect 24506 75076 24530 75108
rect 24632 75084 24684 75108
rect 26248 75102 27048 75124
rect 27290 75102 27302 75158
rect 23996 75050 24060 75070
rect 24132 75062 24194 75070
rect 24002 75044 24024 75050
rect 24130 75048 24194 75062
rect 24278 75052 24342 75070
rect 24284 75046 24306 75052
rect 23968 75022 24088 75042
rect 24104 75034 24222 75042
rect 24012 75018 24024 75022
rect 24102 75020 24222 75034
rect 24250 75024 24370 75042
rect 24256 75018 24306 75024
rect 24002 75016 24024 75018
rect 24002 74954 24012 74962
rect 24094 74952 24226 74972
rect 24480 74956 24498 75076
rect 24506 75074 24600 75076
rect 24502 75062 24600 75074
rect 24506 75052 24600 75062
rect 24508 75028 24572 75048
rect 24582 75044 24600 75052
rect 24508 75008 24526 75028
rect 24554 75016 24572 75028
rect 24508 74984 24572 75008
rect 24002 74926 24012 74934
rect 24128 74930 24192 74938
rect 24126 74918 24192 74930
rect 24490 74910 24498 74956
rect 24518 74938 24526 74984
rect 24530 74956 24584 74980
rect 26390 74952 26934 75102
rect 27270 75034 27330 75054
rect 27376 75034 27412 75036
rect 27458 75034 27612 75158
rect 27362 75014 27412 75028
rect 27290 75000 27612 75014
rect 27712 75000 28052 75034
rect 27260 74906 27270 74958
rect 24558 74822 24586 74840
rect 24620 74822 24684 74840
rect 24506 74807 24545 74822
rect 24506 74790 24530 74807
rect 24632 74800 24684 74822
rect 26382 74804 26440 74836
rect 26540 74804 26598 74836
rect 26698 74804 26756 74836
rect 26856 74804 26914 74836
rect 24532 74790 24558 74792
rect 24506 74776 24563 74790
rect 24586 74776 24631 74790
rect 24506 74766 24558 74776
rect 26382 74736 26383 74737
rect 26439 74736 26440 74737
rect 26540 74736 26541 74737
rect 26597 74736 26598 74737
rect 26698 74736 26699 74737
rect 26755 74736 26756 74737
rect 26856 74736 26857 74737
rect 26913 74736 26914 74737
rect 23968 74676 24088 74686
rect 24474 74678 24496 74694
rect 26282 74678 26316 74736
rect 26381 74735 26441 74736
rect 26539 74735 26599 74736
rect 26697 74735 26757 74736
rect 26855 74735 26915 74736
rect 26382 74720 26440 74735
rect 26540 74720 26598 74735
rect 26698 74720 26756 74735
rect 26856 74720 26914 74735
rect 26382 74692 26400 74720
rect 26894 74692 26914 74720
rect 26382 74679 26440 74692
rect 26540 74679 26598 74692
rect 26698 74679 26756 74692
rect 26856 74679 26914 74692
rect 26381 74678 26441 74679
rect 26539 74678 26599 74679
rect 26697 74678 26757 74679
rect 26855 74678 26915 74679
rect 26978 74678 27014 74736
rect 26382 74677 26383 74678
rect 26439 74677 26440 74678
rect 26540 74677 26541 74678
rect 26597 74677 26598 74678
rect 26698 74677 26699 74678
rect 26755 74677 26756 74678
rect 26856 74677 26857 74678
rect 26913 74677 26914 74678
rect 23996 74648 24060 74658
rect 26382 74578 26440 74608
rect 26540 74578 26598 74608
rect 26698 74578 26756 74608
rect 26856 74578 26914 74608
rect 24522 74552 24536 74558
rect 24186 74508 24208 74546
rect 24522 74514 24538 74552
rect 24556 74522 24572 74556
rect 24164 74486 24218 74508
rect 24220 74478 24242 74512
rect 24450 74500 24468 74508
rect 24522 74506 24536 74514
rect 26382 74494 26440 74526
rect 26540 74494 26598 74526
rect 26698 74494 26756 74526
rect 26856 74494 26914 74526
rect 26382 74426 26383 74427
rect 26439 74426 26440 74427
rect 26540 74426 26541 74427
rect 26597 74426 26598 74427
rect 26698 74426 26699 74427
rect 26755 74426 26756 74427
rect 26856 74426 26857 74427
rect 26913 74426 26914 74427
rect 26282 74368 26316 74426
rect 26381 74425 26441 74426
rect 26539 74425 26599 74426
rect 26697 74425 26757 74426
rect 26855 74425 26915 74426
rect 26382 74410 26440 74425
rect 26540 74410 26598 74425
rect 26698 74410 26756 74425
rect 26856 74410 26914 74425
rect 26382 74382 26400 74410
rect 26894 74382 26914 74410
rect 26382 74369 26440 74382
rect 26540 74369 26598 74382
rect 26698 74369 26756 74382
rect 26856 74369 26914 74382
rect 26381 74368 26441 74369
rect 26539 74368 26599 74369
rect 26697 74368 26757 74369
rect 26855 74368 26915 74369
rect 26978 74368 27014 74426
rect 26382 74367 26383 74368
rect 26439 74367 26440 74368
rect 26540 74367 26541 74368
rect 26597 74367 26598 74368
rect 26698 74367 26699 74368
rect 26755 74367 26756 74368
rect 26856 74367 26857 74368
rect 26913 74367 26914 74368
rect 27086 74298 27130 74878
rect 27290 74870 27756 75000
rect 27280 74764 27756 74870
rect 27290 74760 27504 74764
rect 27646 74762 27756 74764
rect 27290 74728 27448 74760
rect 27502 74724 27616 74760
rect 27712 74724 27756 74762
rect 27814 74724 28052 74762
rect 27814 74722 27880 74724
rect 37404 74720 37424 74868
rect 37432 74740 37452 74840
rect 29536 74678 29572 74682
rect 28834 74548 28878 74628
rect 29492 74618 29550 74654
rect 29492 74554 29493 74555
rect 29549 74554 29550 74555
rect 28768 74482 28944 74548
rect 29392 74496 29428 74554
rect 29491 74553 29551 74554
rect 29492 74534 29550 74553
rect 29492 74516 29512 74534
rect 29530 74516 29550 74534
rect 29492 74497 29550 74516
rect 29491 74496 29551 74497
rect 29614 74496 29650 74554
rect 29492 74495 29493 74496
rect 29549 74495 29550 74496
rect 28768 74460 29002 74482
rect 28768 74394 28944 74460
rect 39730 74440 39752 75246
rect 29492 74396 29550 74432
rect 26382 74268 26440 74298
rect 26540 74268 26598 74298
rect 26698 74268 26756 74298
rect 26856 74268 26914 74298
rect 24150 74216 24152 74244
rect 24290 74216 24292 74244
rect 24438 74216 24440 74244
rect 24116 74182 24152 74210
rect 24256 74182 24292 74210
rect 24404 74182 24440 74210
rect 24448 74198 24534 74208
rect 24622 74198 25020 74208
rect 25164 74194 26898 74208
rect 26804 74190 26898 74194
rect 24476 74170 24534 74180
rect 24622 74170 25020 74180
rect 25164 74166 26926 74180
rect 26776 74162 26926 74166
rect 25020 73980 25156 74004
rect 24992 73952 25184 73976
rect 32784 73948 33138 74102
rect 33340 73936 33392 74032
rect 33538 73968 33594 73980
rect 33658 73948 33694 74032
rect 33822 73966 33878 73980
rect 34092 73968 34192 73980
rect 34030 73966 34248 73968
rect 33844 73948 34248 73966
rect 40434 73948 40444 73956
rect 25122 73902 25522 73908
rect 25122 73874 25550 73880
rect 32794 73860 32834 73878
rect 33340 73824 33694 73936
rect 33912 73928 34056 73948
rect 34248 73929 34316 73948
rect 34233 73928 34316 73929
rect 40316 73928 40444 73948
rect 33912 73914 34316 73928
rect 40433 73917 40444 73928
rect 48024 73948 48034 73956
rect 48024 73928 48152 73948
rect 48024 73917 48035 73928
rect 33912 73896 34248 73914
rect 33822 73882 33878 73896
rect 33912 73892 33948 73896
rect 33982 73892 34018 73896
rect 33878 73866 33890 73878
rect 33860 73832 33868 73848
rect 33912 73832 34018 73892
rect 34042 73884 34242 73896
rect 34042 73864 34092 73884
rect 34114 73853 34182 73868
rect 34192 73864 34242 73884
rect 34248 73860 34286 73870
rect 34282 73842 34336 73852
rect 34344 73842 34412 73892
rect 34032 73832 34038 73842
rect 34066 73832 34172 73842
rect 33200 73812 33694 73824
rect 33734 73824 34172 73832
rect 34282 73824 34412 73842
rect 33734 73812 34344 73824
rect 33228 73784 33320 73796
rect 32784 73616 33138 73752
rect 33340 73714 33694 73812
rect 33826 73806 33948 73812
rect 33976 73809 34038 73812
rect 33982 73806 34038 73809
rect 34114 73808 34344 73812
rect 34096 73806 34378 73808
rect 33826 73804 33877 73806
rect 33896 73804 33948 73806
rect 34019 73804 34378 73806
rect 33734 73796 34378 73804
rect 33734 73784 34138 73796
rect 33836 73782 33976 73784
rect 33838 73778 33976 73782
rect 33988 73780 34138 73784
rect 33896 73767 33976 73778
rect 33881 73753 33976 73767
rect 33986 73778 34138 73780
rect 33986 73758 34134 73778
rect 33986 73753 34102 73758
rect 34172 73756 34173 73796
rect 34182 73766 34234 73796
rect 33881 73752 34102 73753
rect 34140 73753 34173 73756
rect 34298 73753 34330 73796
rect 34332 73790 34378 73796
rect 34332 73774 34386 73790
rect 34336 73753 34396 73774
rect 34400 73753 34412 73824
rect 34140 73752 34412 73753
rect 33912 73740 33976 73752
rect 34104 73748 34138 73752
rect 34140 73748 34190 73752
rect 33388 73696 33422 73710
rect 33880 73700 33882 73710
rect 33912 73704 33948 73740
rect 34040 73736 34190 73748
rect 34298 73740 34330 73752
rect 33978 73712 34342 73736
rect 33896 73690 33948 73704
rect 33976 73706 34342 73712
rect 33976 73696 34182 73706
rect 34202 73698 34342 73706
rect 33912 73684 33948 73690
rect 33978 73686 34182 73696
rect 33962 73684 34316 73686
rect 33340 73668 33422 73682
rect 32634 73546 32662 73610
rect 32832 73598 32834 73612
rect 33340 73586 33392 73668
rect 33538 73618 33594 73630
rect 33822 73616 33878 73630
rect 33912 73618 34316 73684
rect 33912 73603 34092 73618
rect 34202 73610 34316 73618
rect 25210 73300 25546 73308
rect 25210 73272 25574 73280
rect 28550 73226 28558 73276
rect 28584 73248 28592 73300
rect 32784 73266 33138 73402
rect 33340 73364 33694 73586
rect 33912 73578 34056 73603
rect 34248 73579 34316 73610
rect 34233 73578 34316 73579
rect 33912 73564 34316 73578
rect 33912 73546 34248 73564
rect 33822 73532 33878 73546
rect 33912 73542 33948 73546
rect 33982 73542 34018 73546
rect 33878 73516 33890 73528
rect 33860 73482 33868 73498
rect 33912 73482 34018 73542
rect 34042 73534 34242 73546
rect 34042 73514 34092 73534
rect 34114 73503 34182 73518
rect 34192 73514 34242 73534
rect 34344 73538 34412 73542
rect 34344 73520 34426 73538
rect 34032 73482 34038 73492
rect 34054 73482 34178 73494
rect 33860 73474 34178 73482
rect 34282 73492 34336 73502
rect 34344 73492 34412 73520
rect 34282 73474 34412 73492
rect 33860 73472 34344 73474
rect 33862 73470 34344 73472
rect 33862 73464 33948 73470
rect 33826 73456 33948 73464
rect 33976 73459 34038 73470
rect 34066 73462 34344 73470
rect 33982 73456 34038 73459
rect 34082 73458 34344 73462
rect 34082 73456 34378 73458
rect 33826 73454 33877 73456
rect 33896 73454 33948 73456
rect 34019 73454 34378 73456
rect 33826 73446 34378 73454
rect 33826 73442 34150 73446
rect 33826 73440 33958 73442
rect 34019 73441 34150 73442
rect 34032 73440 34150 73441
rect 33826 73438 33976 73440
rect 33836 73432 33976 73438
rect 33838 73428 33976 73432
rect 33988 73430 34138 73440
rect 33896 73417 33976 73428
rect 33881 73403 33976 73417
rect 33986 73428 34138 73430
rect 33986 73408 34134 73428
rect 33986 73403 34102 73408
rect 34172 73406 34173 73446
rect 34182 73416 34234 73446
rect 33881 73402 34102 73403
rect 34140 73403 34173 73406
rect 34298 73403 34330 73446
rect 34332 73440 34378 73446
rect 34332 73424 34386 73440
rect 34336 73403 34396 73424
rect 34400 73403 34412 73474
rect 34140 73402 34412 73403
rect 33912 73390 33976 73402
rect 34104 73398 34138 73402
rect 34140 73398 34190 73402
rect 33388 73346 33436 73360
rect 33880 73350 33882 73360
rect 33912 73354 33948 73390
rect 34040 73386 34190 73398
rect 34298 73390 34330 73402
rect 34340 73386 34374 73402
rect 33978 73382 34374 73386
rect 33978 73362 34342 73382
rect 40166 73368 40176 73386
rect 33896 73340 33948 73354
rect 33976 73356 34342 73362
rect 33976 73346 34182 73356
rect 34202 73348 34342 73356
rect 33912 73334 33948 73340
rect 33978 73336 34182 73346
rect 40194 73340 40260 73366
rect 40374 73362 40386 73456
rect 40402 73390 40414 73484
rect 40640 73340 40856 73366
rect 41218 73364 41250 73392
rect 41300 73362 41338 73390
rect 46660 73374 47322 73540
rect 48054 73414 48066 73484
rect 48082 73414 48094 73456
rect 47896 73402 47996 73414
rect 48040 73402 48140 73414
rect 48054 73390 48066 73402
rect 47130 73372 47168 73374
rect 47130 73366 47298 73372
rect 33962 73334 34316 73336
rect 33340 73318 33436 73332
rect 32832 73234 32880 73262
rect 33340 73236 33392 73318
rect 33538 73268 33594 73280
rect 33822 73266 33878 73280
rect 33912 73268 34316 73334
rect 40260 73330 40640 73340
rect 40328 73302 40428 73330
rect 40472 73314 40572 73330
rect 40856 73314 40882 73340
rect 47828 73330 47896 73374
rect 47996 73330 48040 73374
rect 48082 73362 48094 73402
rect 48140 73330 48208 73374
rect 47840 73320 47864 73322
rect 47896 73320 47996 73330
rect 48040 73320 48140 73330
rect 40328 73298 40386 73302
rect 33436 73248 33482 73264
rect 33912 73253 34092 73268
rect 34202 73260 34316 73268
rect 27968 73202 28038 73204
rect 32654 73196 32662 73232
rect 27996 73122 28024 73176
rect 28392 73124 28556 73146
rect 28432 73118 28458 73124
rect 27968 73094 28052 73118
rect 28364 73108 28584 73118
rect 28364 73102 28604 73108
rect 28364 73100 28606 73102
rect 28372 73096 28606 73100
rect 28402 73088 28458 73096
rect 28584 73092 28606 73096
rect 28402 73078 28468 73088
rect 28556 73086 28576 73092
rect 28404 73076 28430 73078
rect 28432 73076 28458 73078
rect 28404 73042 28496 73076
rect 28408 73014 28496 73042
rect 28552 73034 28576 73086
rect 28584 73058 28608 73092
rect 28584 73050 28606 73058
rect 28584 73044 28604 73050
rect 28552 73028 28560 73034
rect 27996 72938 28024 72972
rect 28024 72856 28030 72890
rect 28052 72884 28058 72918
rect 28114 72884 28116 72932
rect 28052 72874 28116 72884
rect 28142 72856 28144 72914
rect 28338 72856 28352 72862
rect 28366 72856 28380 72890
rect 28024 72846 28144 72856
rect 28404 72844 28430 72908
rect 28432 72824 28458 72936
rect 32784 72916 33138 73052
rect 33340 73014 33694 73236
rect 33912 73228 34056 73253
rect 34248 73229 34316 73260
rect 34233 73228 34316 73229
rect 33912 73214 34316 73228
rect 40260 73272 40328 73274
rect 40340 73272 40386 73298
rect 40472 73284 41080 73314
rect 41656 73304 41694 73310
rect 47840 73304 48210 73320
rect 40260 73268 40434 73272
rect 40474 73268 40576 73284
rect 40812 73280 40944 73284
rect 33912 73196 34248 73214
rect 40260 73200 40640 73268
rect 40704 73214 40782 73268
rect 40856 73214 40882 73280
rect 40974 73214 41054 73268
rect 41146 73238 41174 73274
rect 41656 73270 41658 73304
rect 41678 73270 41694 73304
rect 41656 73264 41694 73270
rect 41712 73254 41728 73288
rect 47846 73282 48210 73304
rect 47846 73268 47890 73282
rect 47988 73276 48210 73282
rect 47988 73268 47994 73276
rect 48082 73268 48128 73276
rect 47846 73228 47892 73268
rect 33822 73182 33878 73196
rect 33912 73192 33948 73196
rect 33982 73192 34018 73196
rect 33878 73166 33890 73178
rect 33860 73132 33868 73148
rect 33912 73132 34018 73192
rect 34042 73184 34242 73196
rect 34042 73164 34092 73184
rect 34114 73153 34182 73168
rect 34192 73164 34242 73184
rect 34344 73188 34412 73192
rect 34344 73170 34426 73188
rect 34032 73132 34038 73142
rect 34054 73132 34178 73144
rect 33860 73124 34178 73132
rect 34282 73142 34336 73152
rect 34344 73142 34412 73170
rect 40232 73169 40640 73200
rect 40678 73169 41080 73214
rect 41738 73176 41750 73186
rect 40221 73159 40640 73169
rect 40667 73159 41091 73169
rect 40194 73158 41091 73159
rect 34282 73124 34412 73142
rect 33860 73122 34344 73124
rect 33862 73120 34344 73122
rect 33862 73114 33948 73120
rect 33826 73106 33948 73114
rect 33976 73109 34038 73120
rect 34066 73112 34344 73120
rect 33982 73106 34038 73109
rect 34082 73108 34344 73112
rect 34082 73106 34378 73108
rect 33826 73104 33877 73106
rect 33896 73104 33948 73106
rect 34019 73104 34378 73106
rect 33826 73096 34378 73104
rect 33826 73092 34150 73096
rect 33826 73090 33958 73092
rect 34019 73091 34150 73092
rect 34032 73090 34150 73091
rect 33826 73088 33976 73090
rect 33836 73082 33976 73088
rect 33838 73078 33976 73082
rect 33988 73080 34138 73090
rect 33896 73067 33976 73078
rect 33881 73053 33976 73067
rect 33986 73078 34138 73080
rect 33986 73058 34134 73078
rect 33986 73053 34102 73058
rect 34172 73056 34173 73096
rect 34182 73066 34234 73096
rect 33881 73052 34102 73053
rect 34140 73053 34173 73056
rect 34298 73053 34330 73096
rect 34332 73090 34378 73096
rect 34332 73074 34386 73090
rect 34336 73053 34396 73074
rect 34400 73053 34412 73124
rect 40388 73106 40390 73158
rect 40416 73100 40516 73158
rect 40698 73114 40704 73158
rect 40782 73114 40788 73158
rect 40970 73114 40974 73158
rect 41054 73114 41058 73158
rect 47846 73138 47890 73228
rect 47988 73118 48050 73268
rect 48104 73250 48210 73268
rect 48154 73214 48210 73250
rect 48082 73166 48128 73168
rect 48074 73118 48128 73166
rect 48152 73118 48210 73168
rect 34140 73052 34412 73053
rect 40316 73084 40408 73100
rect 40316 73068 40410 73084
rect 40416 73078 40434 73100
rect 33912 73040 33976 73052
rect 34104 73048 34138 73052
rect 34140 73048 34190 73052
rect 33388 72996 33436 73010
rect 33880 73000 33882 73010
rect 33912 73004 33948 73040
rect 34040 73036 34190 73048
rect 34298 73040 34330 73052
rect 34336 73036 34374 73052
rect 33978 73032 34374 73036
rect 40316 73040 40408 73068
rect 40418 73040 40434 73078
rect 46860 73070 46884 73076
rect 46890 73072 46894 73082
rect 40316 73032 40434 73040
rect 33978 73012 34342 73032
rect 33896 72990 33948 73004
rect 33976 73006 34342 73012
rect 33976 72996 34182 73006
rect 34202 72998 34342 73006
rect 33912 72984 33948 72990
rect 33978 72986 34182 72996
rect 33962 72984 34316 72986
rect 33340 72968 33436 72982
rect 28552 72830 28560 72880
rect 28586 72852 28594 72904
rect 32654 72846 32662 72902
rect 32832 72884 32880 72912
rect 33340 72884 33392 72968
rect 33538 72918 33594 72930
rect 33822 72916 33878 72930
rect 33912 72918 34316 72984
rect 33436 72898 33482 72914
rect 33912 72903 34092 72918
rect 34202 72910 34316 72918
rect 33912 72878 34056 72903
rect 34248 72879 34316 72910
rect 34233 72878 34316 72879
rect 33912 72864 34316 72878
rect 33912 72846 34248 72864
rect 33538 72834 33594 72846
rect 33822 72832 33878 72846
rect 33912 72842 33948 72846
rect 33982 72842 34018 72846
rect 28392 72812 28570 72824
rect 27996 72782 28024 72788
rect 27996 72754 28038 72782
rect 28316 72752 28358 72778
rect 28384 72774 28392 72784
rect 28416 72766 28508 72782
rect 28048 72726 28066 72742
rect 28320 72740 28322 72752
rect 28348 72744 28350 72750
rect 28320 72732 28328 72740
rect 28320 72726 28322 72732
rect 28020 72672 28028 72706
rect 28048 72700 28056 72726
rect 28348 72718 28392 72744
rect 28348 72704 28356 72718
rect 28348 72700 28354 72704
rect 28404 72700 28412 72750
rect 28416 72702 28418 72724
rect 28048 72676 28110 72700
rect 28320 72672 28326 72700
rect 28348 72686 28412 72700
rect 28380 72672 28384 72686
rect 28020 72648 28138 72672
rect 28320 72658 28412 72672
rect 28432 72658 28440 72766
rect 28576 72652 28582 72702
rect 28610 72672 28616 72724
rect 28224 72638 28356 72644
rect 28402 72638 28453 72643
rect 28402 72630 28458 72638
rect 28252 72610 28328 72616
rect 27996 72550 28024 72588
rect 28320 72580 28366 72582
rect 28404 72580 28430 72610
rect 28320 72558 28430 72580
rect 28320 72556 28366 72558
rect 28320 72548 28322 72556
rect 28348 72546 28366 72554
rect 28372 72552 28430 72558
rect 28404 72546 28430 72552
rect 28348 72538 28414 72546
rect 28348 72526 28416 72538
rect 28348 72524 28418 72526
rect 28348 72502 28354 72524
rect 28320 72488 28326 72502
rect 28348 72494 28384 72502
rect 28348 72488 28354 72494
rect 28380 72464 28384 72494
rect 28404 72488 28412 72524
rect 28416 72504 28418 72524
rect 28432 72518 28458 72630
rect 32606 72580 32642 72588
rect 32784 72566 33138 72716
rect 33340 72664 33392 72820
rect 33878 72816 33890 72828
rect 33440 72774 33496 72786
rect 33860 72782 33868 72798
rect 33912 72782 34018 72842
rect 34042 72834 34242 72846
rect 34042 72814 34092 72834
rect 34114 72803 34182 72818
rect 34192 72814 34242 72834
rect 34344 72838 34412 72842
rect 34344 72820 34426 72838
rect 40194 72834 40200 72958
rect 40354 72902 40380 73032
rect 40382 72930 40408 73032
rect 40698 72958 40704 73056
rect 40782 72958 40788 73056
rect 40418 72944 40460 72948
rect 40474 72944 40486 72948
rect 40372 72894 40380 72902
rect 40400 72894 40408 72902
rect 40418 72900 40486 72944
rect 40364 72846 40432 72894
rect 40400 72824 40408 72846
rect 40550 72834 40856 72958
rect 40970 72956 40974 73056
rect 41054 72956 41058 73056
rect 46888 73048 46916 73072
rect 46928 73060 46952 73062
rect 46928 73054 46950 73060
rect 46794 73030 46874 73044
rect 46888 73020 46916 73044
rect 46962 73026 46986 73028
rect 46962 73022 46984 73026
rect 41656 72906 41694 72912
rect 41656 72872 41658 72906
rect 41682 72872 41694 72894
rect 41656 72866 41694 72872
rect 41716 72826 41750 72860
rect 34032 72782 34038 72792
rect 34054 72782 34178 72794
rect 33860 72774 34178 72782
rect 34282 72792 34336 72802
rect 34344 72792 34412 72820
rect 41390 72810 41404 72816
rect 34282 72774 34412 72792
rect 33860 72772 34344 72774
rect 33862 72770 34344 72772
rect 33862 72764 33948 72770
rect 33826 72756 33948 72764
rect 33976 72759 34038 72770
rect 34066 72762 34344 72770
rect 33982 72756 34038 72759
rect 34082 72758 34344 72762
rect 34082 72756 34378 72758
rect 33826 72754 33877 72756
rect 33896 72754 33948 72756
rect 34019 72754 34378 72756
rect 33826 72746 34378 72754
rect 33826 72742 34150 72746
rect 33826 72740 33958 72742
rect 34019 72741 34150 72742
rect 34032 72740 34150 72741
rect 33826 72738 33976 72740
rect 33836 72732 33976 72738
rect 33838 72728 33976 72732
rect 33988 72730 34138 72740
rect 33896 72717 33976 72728
rect 33881 72703 33976 72717
rect 33986 72728 34138 72730
rect 33986 72708 34134 72728
rect 33986 72703 34102 72708
rect 34172 72706 34173 72746
rect 34182 72716 34234 72746
rect 33881 72702 34102 72703
rect 34140 72703 34173 72706
rect 34298 72703 34330 72746
rect 34332 72740 34378 72746
rect 34332 72724 34386 72740
rect 34336 72703 34396 72724
rect 34400 72703 34412 72774
rect 41388 72764 41404 72810
rect 41418 72782 41432 72790
rect 40432 72742 40442 72750
rect 41416 72744 41432 72782
rect 41798 72752 41806 72910
rect 41826 72780 41834 72882
rect 40314 72722 40442 72742
rect 34140 72702 34412 72703
rect 33440 72690 33496 72702
rect 33912 72690 33976 72702
rect 34104 72698 34138 72702
rect 34140 72698 34190 72702
rect 33912 72664 33948 72690
rect 34040 72686 34190 72698
rect 34298 72690 34330 72702
rect 34342 72686 34374 72702
rect 33880 72650 33882 72660
rect 33978 72641 33991 72686
rect 34140 72682 34374 72686
rect 34140 72668 34342 72682
rect 34138 72658 34342 72668
rect 34140 72656 34342 72658
rect 34202 72648 34342 72656
rect 34040 72602 34140 72614
rect 28432 72460 28440 72518
rect 28576 72454 28582 72504
rect 28610 72474 28616 72526
rect 32634 72496 32662 72560
rect 32794 72460 32842 72488
rect 33382 72460 33444 72488
rect 34248 72460 34306 72488
rect 40372 72482 40380 72686
rect 40400 72510 40408 72714
rect 40431 72711 40442 72722
rect 41750 72728 41788 72734
rect 41750 72724 41766 72728
rect 41772 72724 41788 72728
rect 41750 72712 41788 72724
rect 41658 72692 41696 72698
rect 40420 72670 40442 72692
rect 40412 72638 40466 72670
rect 41658 72658 41660 72692
rect 41688 72658 41696 72692
rect 41722 72688 41788 72712
rect 41936 72708 42598 72766
rect 41806 72706 41840 72708
rect 41932 72706 42598 72708
rect 41806 72700 41822 72706
rect 41722 72678 41756 72688
rect 41798 72666 41822 72700
rect 41916 72678 42598 72706
rect 41658 72652 41696 72658
rect 40418 72632 40442 72638
rect 40418 72602 40460 72632
rect 40424 72600 40460 72602
rect 41478 72596 41534 72622
rect 41936 72600 42598 72678
rect 41936 72598 42294 72600
rect 28402 72440 28453 72445
rect 28402 72432 28458 72440
rect 27982 72392 28024 72420
rect 28404 72406 28430 72412
rect 27996 72358 28024 72392
rect 28252 72348 28430 72406
rect 27982 72312 28024 72336
rect 27982 72308 27996 72312
rect 28010 72288 28024 72312
rect 28252 72328 28416 72348
rect 28252 72306 28418 72328
rect 28432 72320 28458 72432
rect 40372 72432 40388 72482
rect 40400 72460 40416 72510
rect 40698 72482 40704 72582
rect 40782 72482 40788 72582
rect 40970 72482 40974 72582
rect 41054 72482 41058 72582
rect 41506 72568 41562 72594
rect 41948 72508 41960 72598
rect 41976 72596 42040 72598
rect 42048 72596 42068 72598
rect 41976 72536 41988 72596
rect 42020 72536 42144 72596
rect 42436 72550 42452 72600
rect 42464 72578 42506 72600
rect 42558 72584 42596 72600
rect 42640 72588 42682 72616
rect 42048 72508 42068 72536
rect 41936 72464 41964 72500
rect 40372 72404 40390 72432
rect 40400 72404 40418 72460
rect 28252 72290 28416 72306
rect 28432 72290 28440 72320
rect 28010 72280 28052 72288
rect 28252 72266 28488 72290
rect 28252 72236 28496 72266
rect 28252 72234 28458 72236
rect 27982 72194 28024 72222
rect 28252 72214 28416 72234
rect 28252 72194 28430 72214
rect 27996 72166 28430 72194
rect 28010 72152 28430 72166
rect 28010 72062 28380 72152
rect 28404 72150 28430 72152
rect 28432 72122 28458 72234
rect 28484 72220 28496 72236
rect 28512 72192 28524 72294
rect 28576 72256 28582 72306
rect 28610 72276 28616 72328
rect 32806 72248 33160 72394
rect 32854 72226 32902 72248
rect 33442 72226 33504 72254
rect 33934 72248 34434 72394
rect 40329 72393 40442 72404
rect 40340 72372 40394 72393
rect 40400 72380 40442 72393
rect 40340 72362 40386 72372
rect 40400 72362 40446 72380
rect 35590 72256 35764 72362
rect 40340 72356 40446 72362
rect 40340 72346 40442 72356
rect 40340 72338 40414 72346
rect 35590 72254 35926 72256
rect 34308 72218 34366 72248
rect 35590 72194 35622 72254
rect 35758 72186 35790 72254
rect 40272 72216 40274 72220
rect 40318 72210 40320 72278
rect 40340 72267 40386 72338
rect 40392 72322 40414 72338
rect 40329 72262 40397 72267
rect 40400 72262 40414 72322
rect 40418 72322 40442 72346
rect 40698 72324 40704 72424
rect 40782 72324 40788 72424
rect 40970 72324 40974 72424
rect 41054 72324 41058 72424
rect 41736 72396 41748 72406
rect 41898 72396 41934 72398
rect 41932 72394 41934 72396
rect 43156 72378 43400 72994
rect 45068 72612 45312 72994
rect 46922 72974 46942 73008
rect 46962 72982 46976 73022
rect 47248 73014 47274 73102
rect 47952 73100 48050 73118
rect 47276 73014 47302 73074
rect 47000 73006 47012 73008
rect 46922 72960 46936 72974
rect 46794 72946 46874 72960
rect 47088 72954 47316 72990
rect 46846 72908 46854 72930
rect 46794 72896 46874 72908
rect 46732 72848 46748 72864
rect 46754 72848 46762 72866
rect 46818 72864 46826 72896
rect 46846 72892 46854 72896
rect 46870 72848 46880 72858
rect 46748 72832 46764 72838
rect 46886 72832 46902 72848
rect 46794 72812 46874 72824
rect 46990 72786 47316 72954
rect 47612 72834 47914 73048
rect 48034 73032 48050 73100
rect 48062 73090 48152 73100
rect 48074 73056 48152 73090
rect 48074 73040 48144 73056
rect 47978 72944 47994 72948
rect 48008 72944 48050 72948
rect 47978 72900 48050 72944
rect 48060 72894 48064 72902
rect 48088 72894 48092 72930
rect 48032 72846 48104 72894
rect 48032 72822 48054 72838
rect 48060 72824 48064 72846
rect 48264 72834 48274 72958
rect 47052 72780 47250 72786
rect 47052 72778 47062 72780
rect 46530 72736 46798 72766
rect 46860 72736 47182 72750
rect 46104 72652 46106 72668
rect 46080 72612 46108 72652
rect 46228 72650 46268 72678
rect 46430 72612 46494 72704
rect 45034 72584 45312 72612
rect 45068 72378 45312 72584
rect 46104 72576 46106 72612
rect 46338 72584 46376 72612
rect 46426 72600 46494 72612
rect 46430 72596 46494 72600
rect 46530 72598 46748 72736
rect 46754 72644 46768 72736
rect 47046 72686 47182 72736
rect 47456 72732 47494 72756
rect 47514 72732 47522 72764
rect 46754 72634 46776 72644
rect 46760 72620 46776 72634
rect 45830 72534 45876 72568
rect 46106 72500 46272 72576
rect 46494 72536 46598 72596
rect 46630 72568 46748 72598
rect 46834 72582 47182 72686
rect 47300 72710 47556 72732
rect 47300 72692 47586 72710
rect 47766 72704 47810 72794
rect 47966 72782 47978 72800
rect 47932 72748 47944 72782
rect 47966 72766 47982 72782
rect 47932 72732 47950 72748
rect 48022 72742 48032 72750
rect 48022 72722 48150 72742
rect 48022 72711 48033 72722
rect 47300 72682 47556 72692
rect 47300 72652 47572 72682
rect 47612 72666 47810 72704
rect 47584 72660 47810 72666
rect 47922 72664 47944 72692
rect 48022 72670 48048 72692
rect 47892 72660 47944 72664
rect 47584 72658 47944 72660
rect 47584 72652 47810 72658
rect 46834 72568 47256 72582
rect 46630 72462 47256 72568
rect 47268 72542 47274 72628
rect 47300 72626 47810 72652
rect 47892 72644 47944 72658
rect 47922 72638 47944 72644
rect 47998 72638 48052 72670
rect 47828 72626 47944 72638
rect 48022 72632 48050 72638
rect 47300 72624 47944 72626
rect 47300 72604 47810 72624
rect 47828 72604 47944 72624
rect 47300 72600 47944 72604
rect 48008 72602 48050 72632
rect 48008 72600 48044 72602
rect 47296 72582 47944 72600
rect 47296 72570 47556 72582
rect 47300 72564 47556 72570
rect 47584 72574 47944 72582
rect 47584 72570 47810 72574
rect 47828 72570 47944 72574
rect 47584 72564 47944 72570
rect 47596 72556 47780 72564
rect 47612 72548 47780 72556
rect 47600 72546 47780 72548
rect 47318 72538 47350 72546
rect 47424 72538 47542 72540
rect 47596 72520 47780 72546
rect 47808 72540 47944 72564
rect 47824 72536 47944 72540
rect 47828 72524 47944 72536
rect 47290 72510 47322 72518
rect 47452 72510 47514 72512
rect 47420 72494 47452 72510
rect 47534 72508 47596 72520
rect 47454 72494 47486 72504
rect 47420 72462 47486 72494
rect 47510 72496 47518 72504
rect 47510 72462 47520 72496
rect 47534 72483 47554 72508
rect 47544 72466 47554 72483
rect 47566 72466 47584 72508
rect 47588 72505 47596 72508
rect 47600 72480 47618 72520
rect 47650 72519 47780 72520
rect 47662 72482 47702 72498
rect 47712 72482 47780 72519
rect 47808 72500 47944 72524
rect 48060 72510 48064 72714
rect 47808 72494 47824 72500
rect 47828 72494 47944 72500
rect 47650 72480 47712 72482
rect 47612 72472 47718 72480
rect 47596 72466 47718 72472
rect 47534 72462 47718 72466
rect 46080 72416 46108 72456
rect 46630 72432 47274 72462
rect 47420 72446 47718 72462
rect 47420 72444 47452 72446
rect 47276 72432 47302 72434
rect 46630 72424 47302 72432
rect 47424 72424 47430 72444
rect 47484 72442 47718 72446
rect 46630 72414 47088 72424
rect 46810 72404 46822 72414
rect 46794 72390 46874 72404
rect 46810 72386 46822 72390
rect 46990 72388 47044 72404
rect 47248 72398 47274 72424
rect 47276 72398 47302 72424
rect 47456 72414 47718 72442
rect 47472 72412 47718 72414
rect 47508 72410 47522 72412
rect 47534 72411 47718 72412
rect 47732 72411 47758 72482
rect 47808 72442 47944 72494
rect 48052 72460 48064 72510
rect 48088 72482 48092 72686
rect 47828 72426 47944 72442
rect 47534 72410 47758 72411
rect 46736 72368 46936 72380
rect 46736 72334 46942 72368
rect 46962 72342 46976 72388
rect 47000 72366 47012 72368
rect 47088 72334 47316 72398
rect 47484 72360 47638 72410
rect 47824 72394 47944 72426
rect 48050 72404 48064 72460
rect 48080 72432 48092 72482
rect 48078 72404 48092 72432
rect 48022 72400 48139 72404
rect 47534 72342 47588 72346
rect 47612 72342 47718 72360
rect 41580 72328 41668 72330
rect 40418 72292 40446 72322
rect 41608 72300 41660 72316
rect 40418 72270 40442 72292
rect 40324 72256 40326 72262
rect 40328 72256 40442 72262
rect 40270 72202 40340 72208
rect 40311 72196 40328 72202
rect 40274 72193 40326 72196
rect 40274 72186 40314 72193
rect 28524 72152 28584 72162
rect 28524 72062 28548 72152
rect 32634 71914 32662 71978
rect 32784 71926 33138 72076
rect 33382 72002 33444 72030
rect 34248 71990 34306 72018
rect 33086 71908 33138 71926
rect 33912 71858 33948 71926
rect 34040 71860 34140 71872
rect 33880 71848 33948 71858
rect 33912 71840 33948 71848
rect 33912 71813 34102 71840
rect 34104 71813 34412 71840
rect 32634 71564 32662 71628
rect 32784 71590 33138 71726
rect 32832 71576 32880 71590
rect 32606 71536 32658 71560
rect 33086 71558 33138 71590
rect 33340 71714 33392 71810
rect 33440 71772 33496 71784
rect 33912 71776 34412 71813
rect 33912 71772 34102 71776
rect 34104 71772 34412 71776
rect 33881 71757 33948 71772
rect 33896 71746 33948 71757
rect 34025 71746 34102 71772
rect 34140 71768 34173 71772
rect 33838 71742 33958 71746
rect 34025 71745 34138 71746
rect 34034 71744 34138 71745
rect 33836 71736 33958 71742
rect 34032 71736 34138 71744
rect 33826 71734 34138 71736
rect 33826 71728 34150 71734
rect 34172 71728 34173 71768
rect 34182 71728 34234 71758
rect 34298 71728 34330 71772
rect 34336 71750 34396 71772
rect 34332 71734 34386 71750
rect 34332 71728 34378 71734
rect 33826 71720 34159 71728
rect 33340 71492 33694 71714
rect 33826 71710 33948 71720
rect 33862 71704 33948 71710
rect 33954 71718 34159 71720
rect 33954 71704 34038 71718
rect 34082 71713 34159 71718
rect 34172 71716 34378 71728
rect 34082 71712 34150 71713
rect 34172 71712 34344 71716
rect 34066 71704 34344 71712
rect 33862 71702 34344 71704
rect 33860 71701 34344 71702
rect 34400 71701 34412 71772
rect 33860 71700 34412 71701
rect 33860 71696 34178 71700
rect 33860 71692 34192 71696
rect 33860 71688 33868 71692
rect 33848 71676 33868 71688
rect 33912 71664 34018 71692
rect 34032 71682 34038 71692
rect 34054 71680 34192 71692
rect 33822 71628 33878 71642
rect 33912 71628 34014 71664
rect 34092 71660 34192 71680
rect 34282 71682 34344 71700
rect 34282 71672 34336 71682
rect 34352 71664 34398 71682
rect 34042 71628 34242 71660
rect 34380 71636 34426 71654
rect 33912 71610 34092 71628
rect 34192 71610 34248 71628
rect 33912 71571 34056 71610
rect 34233 71595 34316 71610
rect 33912 71570 34092 71571
rect 34248 71570 34316 71595
rect 33912 71558 34316 71570
rect 33822 71544 33878 71558
rect 33912 71526 33948 71558
rect 34030 71556 34316 71558
rect 34092 71544 34192 71556
rect 33854 71512 33948 71526
rect 33912 71508 33948 71512
rect 33984 71510 34002 71512
rect 34040 71510 34140 71522
rect 33880 71498 33948 71508
rect 33978 71506 34040 71510
rect 33912 71490 33948 71498
rect 33976 71495 34040 71506
rect 34140 71502 34302 71510
rect 34140 71501 34203 71502
rect 34140 71497 34202 71501
rect 33976 71490 34038 71495
rect 33388 71464 33436 71478
rect 33912 71463 34102 71490
rect 34104 71463 34412 71490
rect 32654 71246 32662 71278
rect 32784 71240 33138 71376
rect 32832 71226 32880 71240
rect 32640 71214 32654 71218
rect 33086 71208 33138 71240
rect 33340 71364 33392 71460
rect 33440 71422 33496 71434
rect 33912 71426 34412 71463
rect 33912 71422 34102 71426
rect 34104 71422 34412 71426
rect 33881 71407 33948 71422
rect 33896 71396 33948 71407
rect 34025 71396 34102 71422
rect 34140 71418 34173 71422
rect 33838 71392 33958 71396
rect 34025 71395 34138 71396
rect 34034 71394 34138 71395
rect 33836 71386 33958 71392
rect 34032 71386 34138 71394
rect 33826 71384 34138 71386
rect 33826 71378 34150 71384
rect 34172 71378 34173 71418
rect 34182 71378 34234 71408
rect 34298 71378 34330 71422
rect 34336 71400 34396 71422
rect 34332 71384 34386 71400
rect 34332 71378 34378 71384
rect 33826 71370 34159 71378
rect 32640 71186 32642 71190
rect 33340 71142 33694 71364
rect 33826 71360 33948 71370
rect 33862 71354 33948 71360
rect 33954 71368 34159 71370
rect 33954 71354 34038 71368
rect 34082 71363 34159 71368
rect 34172 71366 34378 71378
rect 34082 71362 34150 71363
rect 34172 71362 34344 71366
rect 34066 71354 34344 71362
rect 33862 71352 34344 71354
rect 33860 71351 34344 71352
rect 34400 71351 34412 71422
rect 33860 71350 34412 71351
rect 33860 71346 34178 71350
rect 33860 71342 34192 71346
rect 33860 71338 33868 71342
rect 33848 71326 33868 71338
rect 33912 71314 34018 71342
rect 34032 71332 34038 71342
rect 34054 71330 34192 71342
rect 33822 71278 33878 71292
rect 33912 71278 34014 71314
rect 34092 71310 34192 71330
rect 34282 71332 34344 71350
rect 34282 71322 34336 71332
rect 34352 71314 34398 71332
rect 34042 71278 34242 71310
rect 34380 71286 34426 71304
rect 33912 71260 34092 71278
rect 34192 71260 34248 71278
rect 33912 71221 34056 71260
rect 34233 71245 34316 71260
rect 33912 71220 34092 71221
rect 34248 71220 34316 71245
rect 33912 71208 34316 71220
rect 33822 71194 33878 71208
rect 33912 71176 33948 71208
rect 34030 71206 34316 71208
rect 34092 71194 34192 71206
rect 33854 71162 33948 71176
rect 33912 71158 33948 71162
rect 33984 71160 34002 71162
rect 34040 71160 34140 71172
rect 33880 71148 33948 71158
rect 33978 71156 34040 71160
rect 33912 71140 33948 71148
rect 33976 71145 34040 71156
rect 34140 71152 34302 71160
rect 34140 71151 34203 71152
rect 34140 71147 34202 71151
rect 33976 71140 34038 71145
rect 35760 71144 35788 72186
rect 40272 72182 40314 72186
rect 40346 72182 40348 72250
rect 40372 72208 40386 72256
rect 40400 72208 40414 72256
rect 40612 72250 40718 72272
rect 41146 72264 41174 72300
rect 41640 72298 41660 72300
rect 41700 72294 41720 72304
rect 41614 72266 41616 72292
rect 41614 72264 41642 72266
rect 40628 72222 40690 72244
rect 40372 72202 40472 72208
rect 40274 72170 40314 72182
rect 40272 72168 40314 72170
rect 36700 72118 36738 72146
rect 36962 72132 37006 72144
rect 40258 72124 40326 72168
rect 40372 72156 40386 72202
rect 40400 72184 40414 72202
rect 40455 72196 40472 72202
rect 40455 72193 40470 72196
rect 40586 72182 40622 72196
rect 40640 72182 40676 72196
rect 40586 72180 40690 72182
rect 40586 72170 40622 72180
rect 40628 72178 40690 72180
rect 40640 72170 40676 72178
rect 41220 72174 41250 72192
rect 41308 72184 41338 72192
rect 40584 72168 40622 72170
rect 40638 72168 40676 72170
rect 40428 72136 40470 72168
rect 40572 72162 40676 72168
rect 41298 72164 41338 72184
rect 43298 72180 43382 72334
rect 46736 72320 46936 72334
rect 46794 72312 46874 72320
rect 47088 72314 47320 72334
rect 47484 72330 47718 72342
rect 46092 72298 46108 72310
rect 46742 72290 47002 72312
rect 47028 72310 47320 72314
rect 47018 72290 47320 72310
rect 47456 72318 47718 72330
rect 47456 72302 47758 72318
rect 47472 72292 47758 72302
rect 47508 72290 47522 72292
rect 47534 72290 47758 72292
rect 46578 72252 46584 72268
rect 46606 72240 46612 72268
rect 46742 72264 47320 72290
rect 46742 72256 47004 72264
rect 46714 72200 46726 72256
rect 46736 72224 46742 72256
rect 46748 72234 46760 72256
rect 46748 72226 46768 72234
rect 46748 72224 46772 72226
rect 46818 72224 46826 72256
rect 46846 72252 46854 72256
rect 46934 72242 47004 72256
rect 46732 72222 46772 72224
rect 46732 72218 46776 72222
rect 46732 72210 46782 72218
rect 46732 72208 46794 72210
rect 46870 72208 46880 72218
rect 46714 72192 46734 72200
rect 46736 72192 46742 72208
rect 46748 72204 46824 72208
rect 46748 72198 46782 72204
rect 46748 72192 46764 72198
rect 46886 72192 46902 72208
rect 46714 72188 46742 72192
rect 46934 72191 47002 72242
rect 46714 72186 46744 72188
rect 46874 72187 47002 72191
rect 47028 72187 47320 72264
rect 47424 72258 47430 72278
rect 47484 72258 47758 72290
rect 47828 72280 47944 72394
rect 47808 72264 47944 72280
rect 47988 72393 48139 72400
rect 47988 72362 48064 72393
rect 48074 72372 48128 72393
rect 48082 72362 48128 72372
rect 47988 72350 48128 72362
rect 47988 72346 48210 72350
rect 47988 72270 48050 72346
rect 48052 72324 48210 72346
rect 48052 72292 48108 72324
rect 48054 72278 48064 72292
rect 47388 72224 47408 72258
rect 47420 72256 47452 72258
rect 47420 72250 47458 72256
rect 47484 72250 47732 72258
rect 47420 72230 47732 72250
rect 47846 72236 47890 72264
rect 47946 72236 47996 72250
rect 48052 72236 48064 72278
rect 48082 72250 48092 72292
rect 48154 72288 48210 72324
rect 48080 72240 48128 72250
rect 48080 72236 48140 72240
rect 47846 72230 47996 72236
rect 47420 72224 47596 72230
rect 47650 72224 47732 72230
rect 47840 72224 47996 72230
rect 47420 72208 47486 72224
rect 47420 72192 47452 72208
rect 47454 72198 47486 72208
rect 47510 72206 47520 72224
rect 47510 72198 47518 72206
rect 47534 72204 47554 72224
rect 47566 72204 47584 72224
rect 47600 72212 47618 72222
rect 47650 72220 47758 72224
rect 47712 72212 47780 72220
rect 47846 72216 47996 72224
rect 48040 72222 48140 72236
rect 47840 72214 47996 72216
rect 47534 72197 47588 72204
rect 47596 72197 47780 72212
rect 47846 72208 47996 72214
rect 48038 72208 48140 72222
rect 46874 72186 47320 72187
rect 46714 72184 47320 72186
rect 43382 72166 43466 72180
rect 46714 72174 46760 72184
rect 46794 72182 46874 72184
rect 46988 72182 47320 72184
rect 47534 72184 47780 72197
rect 47828 72198 48208 72208
rect 47828 72196 47884 72198
rect 47894 72196 47896 72198
rect 48038 72196 48040 72198
rect 47792 72190 47898 72196
rect 47792 72184 47884 72190
rect 48052 72184 48064 72198
rect 47534 72182 47928 72184
rect 46794 72176 46886 72182
rect 40572 72154 40674 72162
rect 41298 72156 41336 72164
rect 44546 72154 44694 72166
rect 46714 72164 46790 72174
rect 46794 72172 46874 72176
rect 47028 72166 47320 72182
rect 47554 72174 47588 72182
rect 40572 72150 40688 72154
rect 46700 72150 46748 72152
rect 40572 72136 40674 72150
rect 46726 72140 46748 72150
rect 47028 72146 47316 72166
rect 47596 72157 47758 72182
rect 47778 72180 47928 72182
rect 47778 72178 47884 72180
rect 47792 72170 47884 72178
rect 47596 72156 47661 72157
rect 47674 72156 47758 72157
rect 47782 72168 47884 72170
rect 47782 72156 47894 72168
rect 47600 72154 47672 72156
rect 40426 72124 40470 72136
rect 40570 72124 40638 72136
rect 44574 72126 44666 72138
rect 46672 72116 46714 72118
rect 46794 72116 46810 72140
rect 46856 72132 46936 72142
rect 40602 72114 40626 72116
rect 40256 72106 40626 72114
rect 40256 72070 40426 72106
rect 40428 72098 40626 72106
rect 40428 72076 40620 72098
rect 40428 72070 40478 72076
rect 40338 72062 40384 72070
rect 40472 72062 40478 72070
rect 40576 72062 40620 72076
rect 44986 72072 45792 72096
rect 45836 72088 46048 72096
rect 45836 72072 45890 72088
rect 46080 72074 46108 72114
rect 46692 72106 46714 72116
rect 46726 72084 46740 72086
rect 46660 72074 46740 72084
rect 46754 72074 46768 72112
rect 46798 72074 46813 72089
rect 46856 72074 46936 72082
rect 46977 72074 46992 72089
rect 47028 72074 47182 72144
rect 47506 72124 47584 72132
rect 47610 72124 47672 72154
rect 47674 72152 47900 72156
rect 47674 72150 47894 72152
rect 47674 72124 47758 72150
rect 47506 72120 47596 72124
rect 47610 72120 47758 72124
rect 47456 72096 47462 72116
rect 47506 72112 47584 72120
rect 47506 72110 47586 72112
rect 47506 72088 47530 72110
rect 47534 72108 47564 72110
rect 47650 72108 47758 72120
rect 47782 72124 47894 72150
rect 47996 72136 48038 72168
rect 48080 72156 48092 72198
rect 48154 72170 48194 72196
rect 48152 72168 48194 72170
rect 47994 72124 48038 72136
rect 47534 72088 47596 72108
rect 47650 72088 47732 72108
rect 47782 72094 47834 72124
rect 47838 72114 47862 72116
rect 48118 72114 48120 72150
rect 48140 72136 48208 72168
rect 48138 72124 48206 72136
rect 48146 72114 48148 72122
rect 48192 72114 48194 72116
rect 47838 72110 48208 72114
rect 47838 72096 47994 72110
rect 47472 72086 47584 72088
rect 47588 72086 47732 72088
rect 36348 72042 36448 72052
rect 36708 72042 36808 72054
rect 36988 72042 37088 72052
rect 40256 72044 40384 72062
rect 37258 72006 37882 72026
rect 40272 72008 40384 72044
rect 36596 71970 36606 71984
rect 36348 71958 36448 71968
rect 36708 71958 36808 71970
rect 36988 71958 37088 71968
rect 36202 71914 36208 71916
rect 36184 71892 36208 71914
rect 36298 71908 36348 71948
rect 36292 71898 36348 71908
rect 36448 71908 36498 71948
rect 36938 71908 36988 71948
rect 36448 71898 36504 71908
rect 36292 71894 36307 71898
rect 36172 71880 36208 71892
rect 36278 71892 36307 71894
rect 36489 71892 36504 71898
rect 36928 71898 36988 71908
rect 36928 71892 36943 71898
rect 36216 71882 36236 71888
rect 36142 71866 36210 71880
rect 36216 71876 36258 71882
rect 36172 71852 36206 71866
rect 36142 71838 36210 71852
rect 36216 71842 36240 71876
rect 36244 71842 36258 71876
rect 36278 71860 36352 71892
rect 36444 71860 36994 71892
rect 37100 71862 37134 71890
rect 37180 71864 37214 71892
rect 37258 71862 37714 72006
rect 37270 71858 37714 71862
rect 36172 71826 36208 71838
rect 36216 71836 36258 71842
rect 36216 71830 36236 71836
rect 36184 71804 36208 71826
rect 36278 71826 36352 71858
rect 36444 71826 36994 71858
rect 37180 71826 37214 71854
rect 36278 71824 36307 71826
rect 36292 71820 36307 71824
rect 36489 71820 36504 71826
rect 36292 71810 36348 71820
rect 36202 71802 36208 71804
rect 36298 71770 36348 71810
rect 36448 71810 36504 71820
rect 36928 71820 36943 71826
rect 36928 71810 36988 71820
rect 37716 71818 37882 72006
rect 40338 71994 40384 72008
rect 40258 71980 40314 71994
rect 40256 71912 40314 71962
rect 40416 71912 40478 72062
rect 40574 72022 40620 72062
rect 45014 72044 45792 72068
rect 45836 72060 46118 72068
rect 45836 72044 45918 72060
rect 46052 72046 46118 72060
rect 46660 72052 47182 72074
rect 47506 72076 47530 72086
rect 47506 72070 47528 72076
rect 47462 72068 47528 72070
rect 47534 72074 47596 72086
rect 47650 72074 47712 72086
rect 47844 72076 47994 72096
rect 47462 72066 47524 72068
rect 47534 72066 47584 72074
rect 47462 72062 47584 72066
rect 47462 72060 47588 72062
rect 46664 72048 47182 72052
rect 46664 72044 46856 72048
rect 45014 72032 45634 72044
rect 45758 72032 45792 72038
rect 46052 72032 46118 72040
rect 46676 72024 46740 72044
rect 40576 71932 40620 72022
rect 45556 72018 45600 72020
rect 42962 71930 42966 71950
rect 40416 71894 40514 71912
rect 42996 71900 43000 71930
rect 43032 71924 43034 71988
rect 43060 71896 43062 72016
rect 44986 72004 45606 72018
rect 45786 72004 45792 72010
rect 46080 71972 46108 72012
rect 46688 72006 46740 72024
rect 46726 72000 46740 72006
rect 46754 72004 46768 72044
rect 46806 72038 46856 72044
rect 46936 72044 47182 72048
rect 47484 72058 47584 72060
rect 47662 72059 47780 72074
rect 47844 72062 47888 72076
rect 47986 72070 47994 72076
rect 47996 72070 48138 72110
rect 48140 72070 48208 72110
rect 47986 72062 47992 72070
rect 48080 72062 48126 72070
rect 48146 72062 48148 72070
rect 47484 72044 47534 72058
rect 47544 72052 47584 72058
rect 47544 72050 47572 72052
rect 47544 72044 47584 72050
rect 46936 72038 46986 72044
rect 46806 72034 46986 72038
rect 47028 72034 47182 72044
rect 47472 72042 47588 72044
rect 46806 72032 47182 72034
rect 47462 72032 47588 72042
rect 46794 72028 47182 72032
rect 46794 72026 46856 72028
rect 46798 72012 46856 72026
rect 46936 72012 47182 72028
rect 47472 72018 47588 72032
rect 46754 71980 46776 72004
rect 46798 71997 46813 72012
rect 46977 71997 46992 72012
rect 46692 71970 46714 71980
rect 46754 71974 46768 71980
rect 46672 71968 46714 71970
rect 46742 71948 47002 71970
rect 47028 71948 47182 72012
rect 47456 71998 47462 72018
rect 47472 72016 47572 72018
rect 47584 72016 47588 72018
rect 47510 72014 47530 72016
rect 47544 72014 47584 72016
rect 47596 72014 47630 72058
rect 47662 72052 47702 72059
rect 47662 72016 47702 72050
rect 47712 72016 47780 72059
rect 47826 72028 47890 72062
rect 47816 72022 47890 72028
rect 47484 71990 47534 72014
rect 47544 72002 47572 72014
rect 47544 71990 47564 72002
rect 47484 71982 47586 71990
rect 47650 71988 47712 72016
rect 47732 71988 47758 72016
rect 47816 71994 47888 72022
rect 47596 71982 47780 71988
rect 47484 71974 47780 71982
rect 47484 71966 47544 71974
rect 47584 71966 47780 71974
rect 47484 71964 47780 71966
rect 46742 71946 47182 71948
rect 47506 71946 47584 71964
rect 47596 71956 47780 71964
rect 47610 71948 47780 71956
rect 47600 71946 47780 71948
rect 46726 71942 47222 71946
rect 46726 71936 47002 71942
rect 46700 71934 47002 71936
rect 46742 71930 47002 71934
rect 46742 71926 47060 71930
rect 46630 71918 47088 71926
rect 47534 71920 47562 71938
rect 47596 71920 47780 71946
rect 46630 71914 47222 71918
rect 40314 71850 40404 71894
rect 40314 71834 40392 71850
rect 40416 71834 40432 71894
rect 46630 71892 47088 71914
rect 47142 71902 47222 71914
rect 47420 71894 47452 71910
rect 47506 71904 47514 71912
rect 47534 71908 47596 71920
rect 47454 71894 47486 71904
rect 47096 71892 47112 71894
rect 46630 71888 47112 71892
rect 46630 71850 47096 71888
rect 47158 71878 47222 71892
rect 47262 71878 47316 71892
rect 47294 71866 47326 71876
rect 47158 71850 47222 71864
rect 47262 71850 47320 71864
rect 47420 71862 47486 71894
rect 47506 71896 47518 71904
rect 47506 71866 47520 71896
rect 47534 71894 47562 71908
rect 47534 71883 47554 71894
rect 47544 71866 47554 71883
rect 47566 71866 47584 71908
rect 47588 71905 47596 71908
rect 47600 71880 47618 71920
rect 47650 71919 47780 71920
rect 47662 71882 47702 71898
rect 47712 71882 47780 71919
rect 47826 71932 47888 71994
rect 47650 71880 47712 71882
rect 47610 71872 47718 71880
rect 47596 71866 47718 71872
rect 47510 71862 47520 71866
rect 47534 71862 47718 71866
rect 47420 71852 47718 71862
rect 40314 71826 40432 71834
rect 46052 71832 46120 71844
rect 46630 71832 47088 71850
rect 47420 71846 47458 71852
rect 47420 71844 47452 71846
rect 36448 71770 36498 71810
rect 36938 71770 36988 71810
rect 44878 71788 45068 71818
rect 36348 71750 36448 71760
rect 36708 71748 36808 71760
rect 36988 71750 37088 71760
rect 36594 71734 36606 71748
rect 36894 71724 36908 71742
rect 36348 71666 36448 71676
rect 36574 71610 37258 71724
rect 37720 71684 37756 71744
rect 37774 71684 37810 71740
rect 37498 71642 37526 71674
rect 37692 71672 37756 71684
rect 37774 71572 37816 71672
rect 40192 71628 40854 71752
rect 37692 71556 37756 71572
rect 40400 71556 40568 71628
rect 41340 71616 41404 71624
rect 41362 71588 41414 71596
rect 37720 71536 37756 71556
rect 37638 71504 37756 71536
rect 37774 71514 37810 71556
rect 37774 71506 37996 71514
rect 37638 71450 37756 71482
rect 36348 71402 36448 71412
rect 36708 71402 36808 71414
rect 36892 71382 36912 71392
rect 36920 71382 36940 71420
rect 36988 71402 37088 71412
rect 37720 71410 37756 71450
rect 37774 71452 37996 71460
rect 37774 71410 37810 71452
rect 37774 71404 37840 71410
rect 36790 71330 36868 71374
rect 36928 71336 37016 71374
rect 36348 71318 36448 71328
rect 36708 71318 36808 71330
rect 36892 71328 36912 71336
rect 36920 71328 37016 71336
rect 36920 71320 36940 71328
rect 36844 71308 36962 71320
rect 36988 71318 37088 71328
rect 36202 71274 36208 71276
rect 36184 71252 36208 71274
rect 36298 71268 36348 71308
rect 36292 71258 36348 71268
rect 36448 71268 36498 71308
rect 36448 71258 36504 71268
rect 36292 71254 36307 71258
rect 36172 71240 36208 71252
rect 36278 71252 36307 71254
rect 36489 71252 36504 71258
rect 36844 71258 36988 71308
rect 36844 71252 36896 71258
rect 36908 71254 36962 71258
rect 36928 71252 36966 71254
rect 36216 71242 36236 71248
rect 36142 71226 36210 71240
rect 36216 71236 36258 71242
rect 36172 71212 36206 71226
rect 36142 71198 36210 71212
rect 36216 71202 36240 71236
rect 36244 71202 36258 71236
rect 36278 71220 36352 71252
rect 36444 71236 36896 71252
rect 36444 71228 36876 71236
rect 36908 71228 36976 71252
rect 36444 71220 36976 71228
rect 36986 71220 36994 71252
rect 37100 71222 37134 71250
rect 37180 71224 37214 71252
rect 37258 71220 37524 71386
rect 37774 71334 37816 71404
rect 41936 71394 42332 71560
rect 41936 71392 42204 71394
rect 37692 71326 37768 71334
rect 37638 71310 37768 71326
rect 37692 71276 37768 71310
rect 37594 71220 37606 71246
rect 36844 71218 36962 71220
rect 36172 71186 36208 71198
rect 36216 71196 36258 71202
rect 36216 71190 36236 71196
rect 36184 71164 36208 71186
rect 36278 71186 36352 71218
rect 36444 71186 36918 71218
rect 36278 71184 36307 71186
rect 36292 71180 36307 71184
rect 36489 71180 36504 71186
rect 36292 71170 36348 71180
rect 36202 71162 36208 71164
rect 33388 71114 33436 71128
rect 33912 71113 34102 71140
rect 34104 71113 34412 71140
rect 32634 70864 32662 70928
rect 32784 70890 33138 71026
rect 33086 70858 33138 70890
rect 33340 71014 33392 71110
rect 33440 71072 33496 71084
rect 33912 71076 34412 71113
rect 33912 71072 34102 71076
rect 34104 71072 34412 71076
rect 33881 71057 33948 71072
rect 33896 71046 33948 71057
rect 34025 71046 34102 71072
rect 34140 71068 34173 71072
rect 33838 71042 33958 71046
rect 34025 71045 34138 71046
rect 34034 71044 34138 71045
rect 33836 71036 33958 71042
rect 34032 71036 34138 71044
rect 33826 71034 34138 71036
rect 33826 71028 34150 71034
rect 34172 71028 34173 71068
rect 34182 71028 34234 71058
rect 34298 71028 34330 71072
rect 34336 71050 34396 71072
rect 34332 71034 34386 71050
rect 34332 71028 34378 71034
rect 33826 71020 34159 71028
rect 33340 70792 33694 71014
rect 33826 71010 33948 71020
rect 33862 71004 33948 71010
rect 33954 71018 34159 71020
rect 33954 71004 34038 71018
rect 34082 71013 34159 71018
rect 34172 71016 34378 71028
rect 34082 71012 34150 71013
rect 34172 71012 34344 71016
rect 34066 71004 34344 71012
rect 33862 71002 34344 71004
rect 33860 71001 34344 71002
rect 34400 71001 34412 71072
rect 33860 71000 34412 71001
rect 33860 70996 34178 71000
rect 33860 70992 34192 70996
rect 33860 70988 33868 70992
rect 33848 70976 33868 70988
rect 33912 70964 34018 70992
rect 34032 70982 34038 70992
rect 34054 70980 34192 70992
rect 33822 70928 33878 70942
rect 33912 70928 34014 70964
rect 34092 70960 34192 70980
rect 34282 70982 34344 71000
rect 34282 70972 34336 70982
rect 34352 70964 34398 70982
rect 34042 70928 34242 70960
rect 34380 70936 34426 70954
rect 35760 70936 35790 71144
rect 36298 71130 36348 71170
rect 36448 71170 36504 71180
rect 36844 71180 36918 71186
rect 36928 71208 36966 71218
rect 36928 71180 36962 71208
rect 36986 71186 36994 71218
rect 37180 71186 37214 71214
rect 37720 71186 37768 71276
rect 37774 71276 37788 71326
rect 37774 71226 37822 71276
rect 36844 71172 36988 71180
rect 36928 71170 36988 71172
rect 36448 71130 36498 71170
rect 36938 71138 36988 71170
rect 36920 71130 36988 71138
rect 36348 71110 36448 71120
rect 36708 71108 36808 71120
rect 36594 71094 36606 71108
rect 36892 71102 36912 71110
rect 36920 71102 36940 71130
rect 36988 71110 37088 71120
rect 36348 71026 36448 71036
rect 36708 71024 36808 71036
rect 36988 71026 37088 71036
rect 37720 71034 37756 71104
rect 37926 71102 38108 71356
rect 41936 71294 41950 71392
rect 41956 71312 41960 71392
rect 41984 71340 41988 71392
rect 42020 71384 42040 71392
rect 42048 71384 42068 71392
rect 42438 71364 42452 71444
rect 42466 71392 42512 71420
rect 43154 71404 43398 71788
rect 44782 71684 44818 71740
rect 44836 71684 44872 71744
rect 44878 71722 45310 71788
rect 46080 71776 46108 71816
rect 46612 71806 47088 71832
rect 47142 71818 47222 71830
rect 47424 71824 47430 71844
rect 47484 71842 47718 71852
rect 47732 71842 47758 71882
rect 47484 71840 47766 71842
rect 47472 71812 47766 71840
rect 47508 71810 47522 71812
rect 47534 71810 47766 71812
rect 46630 71804 47088 71806
rect 46612 71792 47088 71804
rect 47484 71802 47766 71810
rect 47826 71832 47884 71932
rect 47986 71912 48048 72062
rect 48102 72044 48208 72062
rect 48152 72008 48208 72044
rect 48080 71960 48126 71962
rect 48072 71912 48126 71960
rect 48150 71912 48208 71962
rect 47950 71894 48048 71912
rect 47826 71804 47944 71832
rect 48032 71826 48048 71894
rect 48060 71884 48150 71894
rect 48072 71850 48150 71884
rect 48072 71834 48142 71850
rect 46612 71778 47282 71792
rect 46630 71774 47282 71778
rect 47456 71774 47766 71802
rect 47822 71786 47944 71804
rect 46794 71766 47282 71774
rect 45606 71746 46048 71762
rect 46858 71758 47282 71766
rect 47484 71760 47766 71774
rect 46858 71740 47316 71758
rect 47508 71746 47522 71760
rect 47534 71742 47588 71746
rect 47610 71742 47766 71760
rect 44836 71672 44900 71684
rect 44836 71572 44878 71672
rect 44836 71556 44900 71572
rect 44782 71514 44818 71556
rect 44596 71506 44818 71514
rect 44836 71536 44872 71556
rect 44836 71504 44954 71536
rect 45068 71488 45310 71722
rect 45606 71718 46076 71734
rect 45890 71698 46076 71712
rect 45890 71690 46120 71698
rect 45742 71664 45830 71672
rect 45890 71662 46048 71684
rect 46080 71662 46108 71670
rect 46092 71644 46108 71662
rect 45770 71636 45830 71644
rect 46450 71626 46468 71654
rect 46478 71632 46480 71698
rect 46736 71696 47316 71740
rect 47484 71720 47766 71742
rect 46794 71682 47316 71696
rect 47472 71692 47766 71720
rect 47826 71708 47944 71786
rect 47992 71709 47994 71774
rect 47992 71708 48009 71709
rect 47826 71702 48009 71708
rect 47480 71690 47766 71692
rect 46782 71642 46794 71672
rect 46810 71670 46822 71682
rect 46858 71672 47316 71682
rect 46824 71656 46888 71672
rect 47026 71670 47316 71672
rect 47018 71662 47316 71670
rect 47456 71682 47766 71690
rect 47808 71694 48009 71702
rect 47808 71686 47944 71694
rect 47456 71662 47810 71682
rect 47890 71668 47944 71686
rect 46796 71628 46916 71644
rect 46990 71602 47004 71642
rect 47018 71630 47046 71662
rect 47060 71654 47072 71662
rect 47088 71654 47316 71662
rect 47420 71656 47452 71658
rect 47484 71656 47810 71662
rect 47248 71624 47272 71654
rect 47276 71652 47300 71654
rect 47420 71652 47810 71656
rect 47929 71654 47944 71668
rect 47420 71640 47534 71652
rect 47420 71634 47522 71640
rect 47060 71616 47124 71624
rect 47420 71608 47486 71634
rect 47050 71588 47152 71596
rect 47420 71592 47452 71608
rect 47454 71598 47486 71608
rect 47510 71606 47520 71634
rect 47544 71619 47554 71650
rect 47510 71598 47518 71606
rect 47534 71604 47554 71619
rect 47566 71604 47584 71650
rect 47596 71630 47810 71652
rect 47610 71628 47810 71630
rect 47942 71628 47944 71630
rect 48022 71628 48272 71752
rect 47600 71612 47618 71622
rect 47650 71620 47712 71628
rect 47696 71612 47712 71620
rect 47534 71597 47588 71604
rect 47596 71597 47712 71612
rect 47288 71560 47312 71586
rect 47534 71582 47712 71597
rect 47766 71588 47780 71620
rect 47554 71574 47588 71582
rect 45616 71488 45666 71496
rect 46528 71488 46630 71560
rect 47596 71558 47650 71582
rect 43154 71392 43432 71404
rect 42590 71340 42636 71362
rect 43154 71340 43398 71392
rect 43592 71372 43612 71488
rect 43620 71420 43640 71460
rect 44596 71452 44818 71460
rect 43620 71400 43684 71420
rect 44782 71410 44818 71452
rect 44836 71450 44954 71482
rect 45040 71468 45844 71488
rect 45068 71460 45310 71468
rect 45616 71460 45617 71468
rect 45666 71460 45692 71468
rect 46090 71460 46108 71474
rect 44836 71410 44872 71450
rect 45040 71440 45844 71460
rect 46228 71448 46268 71476
rect 46506 71466 46630 71488
rect 46528 71460 46630 71466
rect 46736 71538 47026 71554
rect 46736 71518 47028 71538
rect 47050 71526 47060 71536
rect 47124 71526 47222 71536
rect 47316 71532 47340 71558
rect 47386 71526 47556 71558
rect 47596 71557 47712 71558
rect 47596 71556 47661 71557
rect 47600 71554 47638 71556
rect 47298 71520 47556 71526
rect 47584 71534 47638 71538
rect 47640 71536 47672 71556
rect 47640 71534 47708 71536
rect 47584 71524 47708 71534
rect 47584 71520 47732 71524
rect 46736 71508 47182 71518
rect 46736 71498 47222 71508
rect 47298 71498 47732 71520
rect 47764 71498 47810 71588
rect 47930 71526 47948 71628
rect 47964 71560 47991 71594
rect 47943 71512 47944 71526
rect 44752 71404 44818 71410
rect 45068 71406 45310 71440
rect 43630 71376 43676 71400
rect 43602 71348 43612 71372
rect 41984 71324 43478 71340
rect 43154 71312 43398 71324
rect 41956 71296 43450 71312
rect 41950 71258 42104 71294
rect 42950 71278 43068 71280
rect 42948 71268 43068 71278
rect 40327 71183 40403 71194
rect 40338 71166 40392 71183
rect 40338 71144 40384 71166
rect 40256 71118 40362 71144
rect 37774 71034 37810 71090
rect 38180 71046 38362 71102
rect 40272 71082 40362 71118
rect 40416 71064 40478 71194
rect 42948 71182 42974 71268
rect 42978 71250 43040 71252
rect 42976 71240 43040 71250
rect 42976 71210 43002 71240
rect 43032 71210 43040 71240
rect 42976 71186 43040 71210
rect 43002 71182 43032 71186
rect 43060 71182 43068 71268
rect 40576 71066 40620 71174
rect 42948 71158 43068 71182
rect 43154 71172 43398 71296
rect 41650 71110 41666 71124
rect 41606 71096 41666 71110
rect 41622 71092 41666 71096
rect 40576 71062 40710 71066
rect 40576 71046 40716 71062
rect 38180 71034 38414 71046
rect 38458 71034 38558 71046
rect 40338 71034 40384 71044
rect 37692 71032 37756 71034
rect 33912 70910 34092 70928
rect 34192 70910 34248 70928
rect 36700 70922 36738 70950
rect 36962 70922 37008 70950
rect 37594 70936 37606 70950
rect 37774 70932 37816 71032
rect 38180 70962 38362 71034
rect 40326 71030 40384 71034
rect 40470 71042 40520 71044
rect 40576 71042 40620 71046
rect 40326 71002 40426 71030
rect 40470 71002 40854 71042
rect 38556 70962 38616 70966
rect 38830 70964 38862 70992
rect 38912 70964 38950 70992
rect 38992 70966 39024 70994
rect 40258 70992 40854 71002
rect 38180 70950 38414 70962
rect 38458 70954 38616 70962
rect 40504 70958 40854 70992
rect 41298 70958 41336 70986
rect 38458 70950 38558 70954
rect 33912 70871 34056 70910
rect 34233 70895 34316 70910
rect 37692 70906 37756 70932
rect 38180 70920 38362 70950
rect 38584 70930 38644 70938
rect 38584 70926 38640 70930
rect 33912 70870 34092 70871
rect 34248 70870 34316 70895
rect 37720 70880 37756 70906
rect 33912 70858 34316 70870
rect 37638 70864 37756 70880
rect 37774 70866 37810 70906
rect 37926 70866 38108 70920
rect 33822 70844 33878 70858
rect 33912 70826 33948 70858
rect 34030 70856 34316 70858
rect 37774 70856 38108 70866
rect 34092 70844 34192 70856
rect 33854 70812 33948 70826
rect 33912 70808 33948 70812
rect 33984 70810 34002 70812
rect 34040 70810 34140 70822
rect 37638 70810 37756 70826
rect 37926 70812 38108 70856
rect 33880 70798 33948 70808
rect 33978 70806 34040 70810
rect 33912 70790 33948 70798
rect 33976 70795 34040 70806
rect 34140 70802 34302 70810
rect 34140 70801 34203 70802
rect 34140 70797 34202 70801
rect 33976 70790 34038 70795
rect 33388 70764 33422 70778
rect 33912 70763 34102 70790
rect 34104 70763 34412 70790
rect 32784 70540 33138 70694
rect 33340 70526 33392 70760
rect 33440 70722 33496 70734
rect 33912 70726 34412 70763
rect 37720 70756 37756 70810
rect 37774 70802 38108 70812
rect 37774 70756 37810 70802
rect 37692 70754 37756 70756
rect 33912 70722 34102 70726
rect 34104 70722 34412 70726
rect 33881 70707 33948 70722
rect 33896 70696 33948 70707
rect 34025 70696 34102 70722
rect 34140 70718 34173 70722
rect 33838 70692 33958 70696
rect 34025 70695 34138 70696
rect 34034 70694 34138 70695
rect 33836 70686 33958 70692
rect 34032 70686 34138 70694
rect 33826 70684 34138 70686
rect 33826 70678 34150 70684
rect 34172 70678 34173 70718
rect 34182 70678 34234 70708
rect 34298 70678 34330 70722
rect 34336 70700 34396 70722
rect 34332 70684 34386 70700
rect 34332 70678 34378 70684
rect 33826 70670 34159 70678
rect 33826 70660 33948 70670
rect 33862 70654 33948 70660
rect 33954 70668 34159 70670
rect 33954 70654 34038 70668
rect 34082 70663 34159 70668
rect 34172 70666 34378 70678
rect 34082 70662 34150 70663
rect 34172 70662 34344 70666
rect 34066 70654 34344 70662
rect 33862 70652 34344 70654
rect 33860 70651 34344 70652
rect 34400 70651 34412 70722
rect 37774 70654 37816 70754
rect 37926 70666 38108 70802
rect 38180 70904 38692 70920
rect 38180 70868 38702 70904
rect 38180 70720 38692 70868
rect 40320 70864 40854 70958
rect 39688 70782 39910 70838
rect 33860 70650 34412 70651
rect 33440 70638 33496 70650
rect 33860 70646 34178 70650
rect 33860 70642 34192 70646
rect 34282 70642 34344 70650
rect 33860 70638 33868 70642
rect 33848 70626 33868 70638
rect 33912 70614 34018 70642
rect 34032 70632 34038 70642
rect 34054 70630 34192 70642
rect 34248 70632 34344 70642
rect 33538 70578 33594 70590
rect 33822 70578 33878 70592
rect 33912 70578 34014 70614
rect 34092 70610 34192 70630
rect 34282 70622 34336 70632
rect 37692 70628 37756 70654
rect 34042 70578 34242 70610
rect 37720 70586 37756 70628
rect 37774 70578 37810 70628
rect 33912 70560 34092 70578
rect 34192 70560 34248 70578
rect 33912 70526 34014 70560
rect 34030 70526 34056 70560
rect 34233 70545 34316 70560
rect 34248 70526 34316 70545
rect 38180 70510 38362 70666
rect 38458 70562 38558 70574
rect 38658 70518 38692 70640
rect 39622 70604 39976 70782
rect 40540 70770 40658 70850
rect 40758 70788 40772 70864
rect 41820 70788 41834 70920
rect 41934 70788 42052 70850
rect 40474 70616 40724 70770
rect 40758 70752 40926 70788
rect 41820 70770 42052 70788
rect 42682 70782 42904 70838
rect 41820 70752 42118 70770
rect 41868 70616 42118 70752
rect 42616 70604 42970 70782
rect 43136 70742 43160 71048
rect 44034 71034 44134 71046
rect 44178 71034 44278 71046
rect 43164 70742 43188 71020
rect 43642 70964 43680 70992
rect 43730 70964 43762 70992
rect 43976 70962 44036 70966
rect 43976 70954 44134 70962
rect 44034 70950 44134 70954
rect 44178 70950 44278 70962
rect 43948 70930 44008 70938
rect 43952 70926 44008 70930
rect 43608 70866 43612 70894
rect 43658 70872 43670 70878
rect 43630 70866 43676 70872
rect 43624 70860 43682 70866
rect 43624 70854 43642 70860
rect 43636 70844 43642 70854
rect 43624 70836 43642 70844
rect 43664 70854 43682 70860
rect 43664 70844 43676 70854
rect 43664 70836 43682 70844
rect 43624 70832 43682 70836
rect 43608 70802 43612 70832
rect 43636 70830 43670 70832
rect 43658 70820 43670 70830
rect 43604 70662 43612 70800
rect 43632 70696 43640 70772
rect 43900 70720 44412 70920
rect 44484 70866 44666 71356
rect 44836 71334 44878 71404
rect 45036 71394 45310 71406
rect 45056 71378 45310 71394
rect 44824 71326 44900 71334
rect 44804 71276 44818 71326
rect 44770 71226 44818 71276
rect 44824 71310 44954 71326
rect 44824 71276 44900 71310
rect 44824 71186 44872 71276
rect 45068 71172 45310 71378
rect 45616 71161 45617 71440
rect 45666 71320 45692 71440
rect 46478 71438 46644 71460
rect 46736 71446 47182 71498
rect 47298 71480 47810 71498
rect 47858 71486 47869 71497
rect 47883 71486 47941 71497
rect 47822 71480 47869 71486
rect 47298 71472 47890 71480
rect 47894 71472 47941 71486
rect 46346 71406 46376 71418
rect 46336 71400 46376 71406
rect 46452 71400 46482 71418
rect 46336 71394 46338 71400
rect 46374 71390 46376 71400
rect 46426 71394 46438 71400
rect 46374 71362 46410 71386
rect 45828 71328 45874 71362
rect 46396 71322 46410 71362
rect 46424 71324 46438 71394
rect 46480 71390 46482 71400
rect 46528 71416 46630 71438
rect 46728 71430 47182 71446
rect 46736 71424 47182 71430
rect 46528 71404 46682 71416
rect 46726 71404 47182 71424
rect 47270 71418 47272 71460
rect 46528 71392 47182 71404
rect 46480 71362 46488 71384
rect 46630 71350 47182 71392
rect 45630 71172 45666 71320
rect 46946 71300 46970 71318
rect 47260 71314 47262 71340
rect 47266 71336 47272 71418
rect 47298 71452 47948 71472
rect 47298 71438 47821 71452
rect 47890 71438 47944 71452
rect 47298 71418 47950 71438
rect 47298 71398 47810 71418
rect 47824 71404 47944 71418
rect 47826 71398 47944 71404
rect 47298 71396 47944 71398
rect 47992 71417 48009 71432
rect 47298 71394 47942 71396
rect 47294 71376 47942 71394
rect 47294 71364 47554 71376
rect 47298 71358 47554 71364
rect 47582 71368 47942 71376
rect 47582 71364 47808 71368
rect 47826 71364 47942 71368
rect 47582 71358 47950 71364
rect 47456 71350 47494 71358
rect 47316 71332 47348 71340
rect 47506 71334 47522 71358
rect 47594 71350 47778 71358
rect 47610 71342 47778 71350
rect 47598 71340 47778 71342
rect 47422 71332 47540 71334
rect 47506 71322 47522 71332
rect 47594 71314 47778 71340
rect 47806 71348 47950 71358
rect 47992 71348 47994 71417
rect 47806 71334 47946 71348
rect 48006 71340 48048 71377
rect 47822 71330 47946 71334
rect 47992 71330 48048 71340
rect 47826 71318 47946 71330
rect 47260 71304 47320 71312
rect 47450 71304 47512 71306
rect 46990 71290 47002 71300
rect 46530 71246 46620 71272
rect 46748 71248 46764 71254
rect 46782 71248 46790 71266
rect 46794 71262 46874 71274
rect 46990 71264 47060 71290
rect 47260 71286 47290 71304
rect 47418 71288 47450 71304
rect 47532 71302 47594 71314
rect 47452 71288 47484 71298
rect 45666 71161 45692 71172
rect 45616 71160 45692 71161
rect 46262 71150 46634 71246
rect 46886 71238 46902 71254
rect 46732 71222 46748 71238
rect 46870 71228 46880 71238
rect 46818 71190 46826 71222
rect 46856 71194 46866 71204
rect 46990 71194 47002 71264
rect 47030 71262 47060 71264
rect 47142 71262 47222 71274
rect 46846 71190 46854 71194
rect 46794 71178 46874 71190
rect 46990 71183 47004 71194
rect 47034 71183 47060 71262
rect 47084 71238 47088 71262
rect 47418 71256 47484 71288
rect 47508 71290 47516 71298
rect 47508 71256 47518 71290
rect 47532 71277 47552 71302
rect 47542 71260 47552 71277
rect 47564 71260 47582 71302
rect 47586 71299 47594 71302
rect 47598 71274 47616 71314
rect 47648 71313 47778 71314
rect 47660 71276 47700 71292
rect 47710 71276 47778 71313
rect 47806 71294 47946 71318
rect 47966 71320 48048 71330
rect 47966 71314 48032 71320
rect 47966 71296 47980 71314
rect 47982 71296 48032 71314
rect 47806 71288 47822 71294
rect 47826 71288 47946 71294
rect 47648 71274 47710 71276
rect 47610 71266 47716 71274
rect 47594 71260 47716 71266
rect 47532 71256 47716 71260
rect 47096 71248 47112 71254
rect 47418 71246 47716 71256
rect 47418 71240 47456 71246
rect 47418 71238 47450 71240
rect 47080 71222 47096 71238
rect 47294 71226 47326 71236
rect 47084 71190 47088 71222
rect 47422 71218 47428 71238
rect 47482 71234 47716 71246
rect 47470 71206 47716 71234
rect 47532 71205 47716 71206
rect 47730 71205 47756 71276
rect 47806 71262 47946 71288
rect 47992 71286 48032 71296
rect 47806 71236 47942 71262
rect 47826 71220 47942 71236
rect 47532 71204 47756 71205
rect 46990 71182 47060 71183
rect 46846 71156 46854 71178
rect 45838 71106 46048 71120
rect 46262 71104 46698 71150
rect 46794 71126 46874 71140
rect 46990 71132 47004 71182
rect 47142 71178 47222 71190
rect 47482 71154 47636 71204
rect 47822 71188 47942 71220
rect 47532 71136 47586 71140
rect 47610 71136 47716 71154
rect 47482 71114 47716 71136
rect 47470 71112 47716 71114
rect 44782 71034 44818 71090
rect 44836 71034 44872 71104
rect 46262 71092 46634 71104
rect 45810 71078 46076 71092
rect 46418 71076 46492 71092
rect 46500 71076 46648 71092
rect 46928 71078 46942 71112
rect 46966 71104 46978 71112
rect 46466 71072 46490 71076
rect 46500 71072 46556 71076
rect 46500 71058 46524 71072
rect 46534 71066 46556 71072
rect 46474 71044 46490 71058
rect 44836 71032 44900 71034
rect 44836 70932 44878 71032
rect 46446 71020 46464 71042
rect 46500 71038 46508 71058
rect 46562 71038 46584 71076
rect 46888 71060 46942 71062
rect 46794 71042 46874 71056
rect 46888 71042 46946 71060
rect 46962 71058 46976 71104
rect 47470 71086 47756 71112
rect 47532 71084 47756 71086
rect 47482 71082 47673 71084
rect 47674 71082 47756 71084
rect 47248 71056 47272 71072
rect 47276 71056 47300 71072
rect 46888 71034 46902 71042
rect 46888 71032 46914 71034
rect 46888 71014 46918 71032
rect 47088 71014 47316 71056
rect 47422 71052 47428 71072
rect 47482 71052 47756 71082
rect 47826 71074 47942 71188
rect 47806 71058 47942 71074
rect 47986 71064 48048 71194
rect 48061 71183 48137 71194
rect 48072 71166 48126 71183
rect 48080 71144 48126 71166
rect 48102 71118 48208 71144
rect 48152 71082 48208 71118
rect 47386 71018 47406 71052
rect 47418 71050 47450 71052
rect 47418 71044 47456 71050
rect 47482 71044 47730 71052
rect 47418 71024 47730 71044
rect 47844 71030 47888 71058
rect 47944 71030 47994 71044
rect 48080 71034 48126 71044
rect 48080 71030 48138 71034
rect 47844 71024 47994 71030
rect 47418 71018 47594 71024
rect 47648 71018 47730 71024
rect 47838 71018 47994 71024
rect 46562 70988 46604 71010
rect 46578 70968 46624 70982
rect 46554 70960 46624 70968
rect 46554 70952 46604 70960
rect 47128 70958 47166 70986
rect 47248 70984 47272 71014
rect 47276 71012 47300 71014
rect 47418 71002 47484 71018
rect 47418 70986 47450 71002
rect 47452 70992 47484 71002
rect 47508 71000 47518 71018
rect 47508 70992 47516 71000
rect 47532 70998 47552 71018
rect 47564 70998 47582 71018
rect 47598 71006 47616 71016
rect 47648 71014 47756 71018
rect 47710 71006 47778 71014
rect 47844 71010 47994 71018
rect 47838 71008 47994 71010
rect 47532 70991 47586 70998
rect 47594 70991 47778 71006
rect 47844 71002 47994 71008
rect 48038 71002 48138 71030
rect 47532 70978 47778 70991
rect 47826 70992 48206 71002
rect 47826 70990 47882 70992
rect 47790 70984 47896 70990
rect 47790 70978 47882 70984
rect 47532 70976 47926 70978
rect 47552 70968 47586 70976
rect 47594 70952 47756 70976
rect 47776 70974 47926 70976
rect 47776 70972 47882 70974
rect 47790 70956 47882 70972
rect 46578 70936 46584 70952
rect 47594 70951 47710 70952
rect 47594 70950 47659 70951
rect 47730 70950 47756 70952
rect 47816 70950 47882 70956
rect 47598 70948 47670 70950
rect 44836 70906 44900 70932
rect 46578 70924 46624 70936
rect 47610 70932 47670 70948
rect 47482 70926 47542 70932
rect 47582 70930 47670 70932
rect 47730 70944 47802 70950
rect 47816 70946 47898 70950
rect 47582 70926 47706 70930
rect 47482 70918 47706 70926
rect 47730 70918 47756 70944
rect 47816 70932 47882 70946
rect 47826 70930 47882 70932
rect 47482 70914 48272 70918
rect 47482 70910 47582 70914
rect 44782 70866 44818 70906
rect 44484 70856 44818 70866
rect 44836 70880 44872 70906
rect 47470 70904 47586 70910
rect 47470 70882 47562 70904
rect 47582 70882 47586 70904
rect 47504 70880 47528 70882
rect 47532 70880 47582 70882
rect 47594 70880 48272 70914
rect 44836 70864 44954 70880
rect 47482 70878 47562 70880
rect 47482 70864 47582 70878
rect 47610 70864 48272 70880
rect 47460 70856 47582 70864
rect 44484 70812 44666 70856
rect 47460 70854 47586 70856
rect 47482 70852 47582 70854
rect 47482 70838 47532 70852
rect 47542 70846 47582 70852
rect 47542 70838 47582 70844
rect 47470 70836 47586 70838
rect 47460 70826 47586 70836
rect 44484 70802 44818 70812
rect 43632 70694 43644 70696
rect 43666 70694 43672 70696
rect 43632 70690 43672 70694
rect 43680 70690 43704 70712
rect 43638 70688 43704 70690
rect 43638 70678 43650 70688
rect 43660 70682 43704 70688
rect 43660 70676 43672 70682
rect 43676 70678 43704 70682
rect 33538 70494 33594 70506
rect 33822 70494 33878 70508
rect 34092 70494 34192 70506
rect 38458 70478 38558 70490
rect 38658 70482 38702 70518
rect 38584 70456 38640 70460
rect 38584 70448 38644 70456
rect 38556 70420 38616 70432
rect 38588 70394 38640 70398
rect 38260 70378 38300 70394
rect 38556 70378 38640 70394
rect 38658 70386 38692 70482
rect 38746 70386 39116 70552
rect 38746 70384 38946 70386
rect 38948 70384 39116 70386
rect 38152 70346 38584 70370
rect 38556 70344 38578 70346
rect 38180 70318 38584 70342
rect 38588 70340 38640 70378
rect 38878 70374 39116 70384
rect 38878 70322 38902 70374
rect 38906 70352 39116 70374
rect 38906 70350 38930 70352
rect 38906 70346 38954 70350
rect 38912 70338 38940 70346
rect 38966 70342 38992 70352
rect 41936 70348 41952 70452
rect 38966 70336 38982 70342
rect 41908 70334 41976 70348
rect 38878 70318 38982 70322
rect 41936 70320 41952 70334
rect 38556 70306 38616 70318
rect 38884 70310 38962 70318
rect 38584 70282 38644 70290
rect 41936 70284 42104 70320
rect 38584 70278 38640 70282
rect 38180 70256 38692 70274
rect 41908 70256 41980 70282
rect 38180 70220 38702 70256
rect 38180 70072 38692 70220
rect 42042 70216 42128 70220
rect 39410 70128 39428 70194
rect 39438 70156 39476 70184
rect 39518 70156 39550 70184
rect 39688 70142 39910 70190
rect 39912 70176 39918 70194
rect 39912 70148 39954 70176
rect 39962 70142 39982 70194
rect 40342 70146 40418 70174
rect 39622 70126 39982 70142
rect 40540 70130 40658 70194
rect 41934 70192 42052 70194
rect 41934 70188 42156 70192
rect 40702 70166 40740 70182
rect 41148 70140 41228 70168
rect 41364 70146 41444 70174
rect 41852 70166 41890 70184
rect 39284 70064 39312 70100
rect 39356 70098 39380 70120
rect 39378 70070 39380 70092
rect 32634 69888 32662 69952
rect 32784 69900 33138 70050
rect 36696 70024 36734 70052
rect 36958 70022 37004 70050
rect 38180 70004 38242 70020
rect 33382 69976 33444 70004
rect 34248 69964 34306 69992
rect 39284 69978 39312 70014
rect 36344 69948 36444 69958
rect 36704 69948 36804 69960
rect 36984 69948 37084 69958
rect 39622 69956 39976 70126
rect 40474 69960 40724 70130
rect 41228 70112 41256 70138
rect 41336 70118 41364 70138
rect 41934 70130 42052 70188
rect 42682 70180 42904 70190
rect 42174 70166 42202 70174
rect 42638 70152 42904 70180
rect 43042 70166 43060 70184
rect 42682 70142 42904 70152
rect 41868 69960 42118 70130
rect 42616 69956 42970 70142
rect 43136 70120 43160 70610
rect 43134 70000 43160 70120
rect 43164 70092 43188 70610
rect 43476 70386 43846 70552
rect 43476 70384 43644 70386
rect 43680 70384 43846 70386
rect 43594 70376 43846 70384
rect 43594 70370 43620 70376
rect 43610 70362 43620 70370
rect 43634 70362 43846 70376
rect 43610 70352 43846 70362
rect 43900 70352 43934 70640
rect 44034 70562 44134 70574
rect 44484 70510 44666 70802
rect 44782 70756 44818 70802
rect 44836 70810 44954 70826
rect 47470 70812 47586 70826
rect 47470 70810 47562 70812
rect 47582 70810 47586 70812
rect 44836 70756 44872 70810
rect 47508 70808 47528 70810
rect 47542 70808 47582 70810
rect 47594 70808 47628 70852
rect 47660 70846 47700 70864
rect 47660 70810 47700 70844
rect 47482 70776 47532 70808
rect 47542 70778 47562 70808
rect 47648 70782 47710 70810
rect 47594 70776 47710 70782
rect 47482 70760 47542 70776
rect 47582 70768 47698 70776
rect 47582 70760 47730 70768
rect 47482 70758 47730 70760
rect 44836 70754 44900 70756
rect 44836 70654 44878 70754
rect 47504 70740 47582 70758
rect 47594 70750 47730 70758
rect 47598 70740 47636 70742
rect 47638 70740 47730 70750
rect 47532 70714 47560 70732
rect 47594 70728 47628 70740
rect 47648 70738 47730 70740
rect 47594 70714 47648 70728
rect 47418 70688 47450 70704
rect 47504 70698 47512 70706
rect 47532 70702 47594 70714
rect 47452 70688 47484 70698
rect 47418 70666 47484 70688
rect 47504 70690 47516 70698
rect 47504 70666 47518 70690
rect 47532 70688 47560 70702
rect 47532 70677 47552 70688
rect 47418 70656 47518 70666
rect 47542 70660 47552 70677
rect 47564 70660 47582 70702
rect 47586 70699 47594 70702
rect 47598 70674 47616 70714
rect 47648 70713 47710 70714
rect 47696 70692 47710 70713
rect 47660 70676 47710 70692
rect 47648 70666 47710 70676
rect 47594 70660 47710 70666
rect 47532 70656 47710 70660
rect 44836 70628 44900 70654
rect 47418 70646 47710 70656
rect 47418 70640 47456 70646
rect 47460 70644 47710 70646
rect 47460 70640 47698 70644
rect 47418 70638 47450 70640
rect 44782 70578 44818 70628
rect 44836 70586 44872 70628
rect 47422 70618 47428 70638
rect 47482 70634 47698 70640
rect 47470 70626 47698 70634
rect 47470 70624 47672 70626
rect 47470 70606 47673 70624
rect 47532 70604 47648 70606
rect 47482 70554 47636 70604
rect 47532 70536 47586 70540
rect 47482 70514 47636 70536
rect 44034 70478 44134 70490
rect 43952 70456 44008 70460
rect 43948 70448 44008 70456
rect 43976 70420 44036 70432
rect 46448 70420 46466 70448
rect 46476 70426 46478 70492
rect 47470 70486 47678 70514
rect 47478 70484 47648 70486
rect 47422 70452 47428 70472
rect 47482 70460 47636 70484
rect 47648 70466 47673 70484
rect 47648 70464 47672 70466
rect 47648 70462 47698 70464
rect 47648 70460 47706 70462
rect 47418 70450 47450 70452
rect 43952 70394 44004 70398
rect 43952 70378 44036 70394
rect 44292 70378 44332 70394
rect 43610 70318 43612 70350
rect 43628 70342 43654 70352
rect 43628 70336 43644 70342
rect 43680 70338 43686 70346
rect 43952 70340 44004 70378
rect 44014 70344 44036 70360
rect 43976 70306 44036 70318
rect 43252 70190 43270 70298
rect 43948 70282 44008 70290
rect 43952 70278 44008 70282
rect 43286 70190 43298 70216
rect 43270 70188 43420 70190
rect 43258 70132 43420 70188
rect 43270 70130 43420 70132
rect 43212 70098 43236 70120
rect 43286 70104 43298 70130
rect 43162 70028 43188 70092
rect 43212 70070 43214 70092
rect 43290 70064 43318 70100
rect 43900 70072 44412 70274
rect 46504 70260 46614 70282
rect 46476 70232 46642 70254
rect 46988 70226 47298 70446
rect 47418 70444 47456 70450
rect 47482 70446 47706 70460
rect 47482 70444 47532 70446
rect 47418 70434 47532 70444
rect 47418 70402 47484 70434
rect 47418 70386 47450 70402
rect 47452 70392 47484 70402
rect 47508 70400 47518 70434
rect 47542 70413 47552 70444
rect 47508 70392 47516 70400
rect 47532 70398 47552 70413
rect 47564 70398 47582 70444
rect 47594 70424 47710 70446
rect 47598 70406 47616 70416
rect 47648 70414 47710 70424
rect 47532 70391 47586 70398
rect 47594 70391 47710 70406
rect 47532 70376 47710 70391
rect 47360 70352 47466 70372
rect 47552 70368 47586 70376
rect 47594 70352 47648 70376
rect 47360 70312 47554 70352
rect 47594 70351 47710 70352
rect 47594 70350 47659 70351
rect 47598 70348 47636 70350
rect 47582 70328 47636 70332
rect 47638 70330 47670 70350
rect 47638 70328 47706 70330
rect 47582 70314 47706 70328
rect 47360 70290 47562 70312
rect 47582 70290 47586 70310
rect 47594 70290 47628 70314
rect 47360 70280 47628 70290
rect 47648 70280 47710 70314
rect 47360 70244 47622 70280
rect 46336 70184 46374 70212
rect 46424 70184 46480 70212
rect 46988 70204 47350 70226
rect 47360 70222 47554 70244
rect 47582 70230 47648 70244
rect 47192 70192 47350 70204
rect 47296 70184 47350 70192
rect 47764 70184 47808 70476
rect 46344 70156 46408 70180
rect 47930 70142 47948 70158
rect 47958 70142 47992 70176
rect 47930 70108 47942 70142
rect 47964 70108 47980 70124
rect 47964 70090 47976 70108
rect 46528 70040 46618 70066
rect 39256 69950 39326 69954
rect 33086 69882 33138 69900
rect 33912 69832 33948 69900
rect 36592 69876 36602 69890
rect 36344 69864 36444 69874
rect 36704 69864 36804 69876
rect 36984 69864 37084 69874
rect 34040 69834 34140 69846
rect 33880 69822 33948 69832
rect 33912 69814 33948 69822
rect 36198 69820 36204 69822
rect 33912 69787 34102 69814
rect 34104 69787 34412 69814
rect 36180 69798 36204 69820
rect 36294 69814 36344 69854
rect 36288 69804 36344 69814
rect 36444 69814 36494 69854
rect 36934 69814 36984 69854
rect 36444 69804 36500 69814
rect 36288 69800 36303 69804
rect 32634 69538 32662 69602
rect 32784 69564 33138 69700
rect 32832 69550 32880 69564
rect 33086 69532 33138 69564
rect 33340 69688 33392 69784
rect 33440 69746 33496 69758
rect 33912 69750 34412 69787
rect 36168 69786 36204 69798
rect 36274 69798 36303 69800
rect 36485 69798 36500 69804
rect 36924 69804 36984 69814
rect 36924 69798 36939 69804
rect 36212 69788 36232 69794
rect 36138 69772 36206 69786
rect 36212 69782 36254 69788
rect 36168 69758 36202 69772
rect 33912 69746 34102 69750
rect 34104 69746 34412 69750
rect 33881 69731 33948 69746
rect 33896 69720 33948 69731
rect 34025 69720 34102 69746
rect 34140 69742 34173 69746
rect 33838 69716 33958 69720
rect 34025 69719 34138 69720
rect 34034 69718 34138 69719
rect 33836 69710 33958 69716
rect 34032 69710 34138 69718
rect 33826 69708 34138 69710
rect 33826 69702 34150 69708
rect 34172 69702 34173 69742
rect 34182 69702 34234 69732
rect 34298 69702 34330 69746
rect 34336 69724 34396 69746
rect 34332 69708 34386 69724
rect 34332 69702 34378 69708
rect 33826 69694 34159 69702
rect 32606 69510 32628 69524
rect 33340 69466 33694 69688
rect 33826 69684 33948 69694
rect 33862 69678 33948 69684
rect 33954 69692 34159 69694
rect 33954 69678 34038 69692
rect 34082 69687 34159 69692
rect 34172 69690 34378 69702
rect 34082 69686 34150 69687
rect 34172 69686 34344 69690
rect 34066 69678 34344 69686
rect 33862 69676 34344 69678
rect 33860 69675 34344 69676
rect 34400 69675 34412 69746
rect 36138 69744 36206 69758
rect 36212 69748 36236 69782
rect 36240 69748 36254 69782
rect 36274 69766 36348 69798
rect 36440 69766 36990 69798
rect 37096 69768 37130 69796
rect 37176 69770 37210 69798
rect 37254 69768 37642 69932
rect 37838 69880 37874 69942
rect 37892 69880 37928 69936
rect 38458 69916 38558 69928
rect 37810 69870 37874 69880
rect 37892 69770 37934 69870
rect 38458 69832 38558 69844
rect 38674 69836 38702 69872
rect 38584 69810 38640 69814
rect 38584 69802 38644 69810
rect 39130 69792 39310 69862
rect 42162 69836 42306 69860
rect 42136 69834 42306 69836
rect 42190 69808 42278 69832
rect 42164 69806 42278 69808
rect 38314 69778 38414 69790
rect 38458 69786 38558 69790
rect 38458 69778 38616 69786
rect 38556 69774 38616 69778
rect 37552 69764 37602 69768
rect 36168 69732 36204 69744
rect 36212 69742 36254 69748
rect 36212 69736 36232 69742
rect 36180 69710 36204 69732
rect 36274 69732 36348 69764
rect 36440 69732 36990 69764
rect 37176 69732 37210 69760
rect 37810 69752 37874 69770
rect 39130 69756 39312 69792
rect 36274 69730 36303 69732
rect 36288 69726 36303 69730
rect 36485 69726 36500 69732
rect 36288 69716 36344 69726
rect 36198 69708 36204 69710
rect 36294 69676 36344 69716
rect 36444 69716 36500 69726
rect 36924 69726 36939 69732
rect 36924 69716 36984 69726
rect 37838 69724 37874 69752
rect 36444 69676 36494 69716
rect 36934 69676 36984 69716
rect 37756 69702 37874 69724
rect 37892 69702 37928 69752
rect 39130 69706 39310 69756
rect 38314 69694 38414 69706
rect 38458 69694 38558 69706
rect 39130 69694 39452 69706
rect 33860 69674 34412 69675
rect 33860 69670 34178 69674
rect 33860 69666 34192 69670
rect 33860 69662 33868 69666
rect 33848 69650 33868 69662
rect 33912 69638 34018 69666
rect 34032 69656 34038 69666
rect 34054 69654 34192 69666
rect 33822 69602 33878 69616
rect 33912 69602 34014 69638
rect 34092 69634 34192 69654
rect 34282 69656 34344 69674
rect 39284 69670 39452 69694
rect 43136 69692 43160 70000
rect 43164 69720 43188 70028
rect 43290 69978 43318 70014
rect 43262 69950 43336 69954
rect 46260 69944 46632 70040
rect 44034 69916 44134 69928
rect 46260 69898 46696 69944
rect 46260 69886 46632 69898
rect 43900 69836 43928 69872
rect 46464 69866 46488 69886
rect 46498 69866 46554 69886
rect 46498 69852 46522 69866
rect 46532 69860 46554 69866
rect 44034 69832 44134 69844
rect 46472 69838 46488 69852
rect 46444 69814 46462 69836
rect 46498 69832 46506 69852
rect 46560 69832 46582 69886
rect 43952 69810 44008 69814
rect 43948 69802 44008 69810
rect 43296 69756 43324 69792
rect 44034 69786 44134 69790
rect 43976 69778 44134 69786
rect 44178 69778 44278 69790
rect 46560 69782 46602 69804
rect 43976 69774 44036 69778
rect 46576 69762 46622 69776
rect 46552 69754 46622 69762
rect 46552 69746 46602 69754
rect 46576 69730 46582 69746
rect 46576 69718 46622 69730
rect 43296 69670 43324 69706
rect 44034 69694 44134 69706
rect 44178 69694 44278 69706
rect 36344 69656 36444 69666
rect 34282 69646 34336 69656
rect 34352 69638 34398 69656
rect 36704 69654 36804 69666
rect 36984 69656 37084 69666
rect 36590 69640 36602 69654
rect 37756 69648 37874 69670
rect 34042 69602 34242 69634
rect 34380 69610 34426 69628
rect 33912 69584 34092 69602
rect 34192 69584 34248 69602
rect 33912 69545 34056 69584
rect 34233 69569 34316 69584
rect 36344 69572 36444 69582
rect 33912 69544 34092 69545
rect 34248 69544 34316 69569
rect 33912 69532 34316 69544
rect 33822 69518 33878 69532
rect 33912 69500 33948 69532
rect 34030 69530 34316 69532
rect 34092 69518 34192 69530
rect 36570 69516 36842 69628
rect 36984 69572 37084 69582
rect 37188 69516 37254 69628
rect 37838 69598 37874 69648
rect 37892 69598 37928 69648
rect 37892 69592 37958 69598
rect 37892 69522 37934 69592
rect 37810 69514 37886 69522
rect 33854 69486 33948 69500
rect 37756 69498 37886 69514
rect 33912 69482 33948 69486
rect 33984 69484 34002 69486
rect 34040 69484 34140 69496
rect 33880 69472 33948 69482
rect 33978 69480 34040 69484
rect 33912 69464 33948 69472
rect 33976 69469 34040 69480
rect 34140 69476 34302 69484
rect 34140 69475 34203 69476
rect 34140 69471 34202 69475
rect 33976 69464 34038 69469
rect 37810 69464 37886 69498
rect 33388 69438 33436 69452
rect 33912 69437 34102 69464
rect 34104 69437 34412 69464
rect 32606 69160 32632 69228
rect 32634 69188 32662 69252
rect 32784 69214 33138 69350
rect 32832 69200 32880 69214
rect 33086 69182 33138 69214
rect 33340 69338 33392 69434
rect 33440 69396 33496 69408
rect 33912 69400 34412 69437
rect 33912 69396 34102 69400
rect 34104 69396 34412 69400
rect 33881 69381 33948 69396
rect 33896 69370 33948 69381
rect 34025 69370 34102 69396
rect 34140 69392 34173 69396
rect 33838 69366 33958 69370
rect 34025 69369 34138 69370
rect 34034 69368 34138 69369
rect 33836 69360 33958 69366
rect 34032 69360 34138 69368
rect 33826 69358 34138 69360
rect 33826 69352 34150 69358
rect 34172 69352 34173 69392
rect 34182 69352 34234 69382
rect 34298 69352 34330 69396
rect 34336 69374 34396 69396
rect 34332 69358 34386 69374
rect 34332 69352 34378 69358
rect 33826 69344 34159 69352
rect 33340 69116 33694 69338
rect 33826 69334 33948 69344
rect 33862 69328 33948 69334
rect 33954 69342 34159 69344
rect 33954 69328 34038 69342
rect 34082 69337 34159 69342
rect 34172 69340 34378 69352
rect 34082 69336 34150 69337
rect 34172 69336 34344 69340
rect 34066 69328 34344 69336
rect 33862 69326 34344 69328
rect 33860 69325 34344 69326
rect 34392 69325 34398 69328
rect 34400 69325 34412 69396
rect 37838 69374 37886 69464
rect 37892 69464 37906 69514
rect 37892 69414 37940 69464
rect 36962 69360 37080 69362
rect 33860 69324 34412 69325
rect 33860 69320 34178 69324
rect 33860 69316 34192 69320
rect 33860 69312 33868 69316
rect 33848 69300 33868 69312
rect 33912 69288 34018 69316
rect 34032 69306 34038 69316
rect 34054 69304 34192 69316
rect 33822 69252 33878 69266
rect 33912 69252 34014 69288
rect 34092 69284 34192 69304
rect 34282 69306 34344 69324
rect 34392 69306 34398 69324
rect 34282 69296 34336 69306
rect 34352 69288 34398 69306
rect 34042 69252 34242 69284
rect 34420 69278 34426 69334
rect 36344 69308 36444 69318
rect 36704 69308 36804 69320
rect 36984 69308 37084 69318
rect 36924 69306 37134 69308
rect 38044 69298 38226 69552
rect 39284 69416 39312 69452
rect 43290 69416 43318 69452
rect 39284 69330 39312 69366
rect 43290 69330 43318 69366
rect 34380 69260 34426 69278
rect 33912 69234 34092 69252
rect 34192 69234 34248 69252
rect 33912 69195 34056 69234
rect 34233 69219 34316 69234
rect 36344 69224 36444 69234
rect 36704 69224 36804 69236
rect 36984 69224 37084 69234
rect 33912 69194 34092 69195
rect 34248 69194 34316 69219
rect 33912 69182 34316 69194
rect 33822 69168 33878 69182
rect 33912 69150 33948 69182
rect 34030 69180 34316 69182
rect 36198 69180 36204 69182
rect 34092 69168 34192 69180
rect 36180 69158 36204 69180
rect 36294 69174 36344 69214
rect 36288 69164 36344 69174
rect 36444 69174 36494 69214
rect 36934 69174 36984 69214
rect 36444 69164 36500 69174
rect 36288 69160 36303 69164
rect 33854 69136 33948 69150
rect 36168 69146 36204 69158
rect 36274 69158 36303 69160
rect 36485 69158 36500 69164
rect 36924 69164 36984 69174
rect 36924 69158 36939 69164
rect 36212 69148 36232 69154
rect 33912 69132 33948 69136
rect 33984 69134 34002 69136
rect 34040 69134 34140 69146
rect 33880 69122 33948 69132
rect 33978 69130 34040 69134
rect 33912 69114 33948 69122
rect 33976 69119 34040 69130
rect 34140 69126 34302 69134
rect 36138 69132 36206 69146
rect 36212 69142 36254 69148
rect 34140 69125 34203 69126
rect 34140 69121 34202 69125
rect 33976 69114 34038 69119
rect 36168 69118 36202 69132
rect 33388 69088 33436 69102
rect 33912 69087 34102 69114
rect 34104 69087 34412 69114
rect 36138 69104 36206 69118
rect 36212 69108 36236 69142
rect 36240 69108 36254 69142
rect 36274 69126 36348 69158
rect 36440 69126 36990 69158
rect 37096 69128 37130 69156
rect 37176 69130 37210 69158
rect 37254 69126 37642 69292
rect 37838 69222 37874 69292
rect 37892 69222 37928 69278
rect 38298 69242 38480 69298
rect 38298 69230 38532 69242
rect 38576 69230 38676 69242
rect 37810 69220 37874 69222
rect 37552 69124 37602 69126
rect 36168 69092 36204 69104
rect 36212 69102 36254 69108
rect 36212 69096 36232 69102
rect 32634 68838 32662 68902
rect 32784 68864 33138 69000
rect 33086 68832 33138 68864
rect 33340 68988 33392 69084
rect 33440 69046 33496 69058
rect 33912 69050 34412 69087
rect 36180 69070 36204 69092
rect 36274 69092 36348 69124
rect 36440 69092 36990 69124
rect 37892 69120 37934 69220
rect 38298 69158 38480 69230
rect 38674 69158 38734 69162
rect 38298 69146 38532 69158
rect 38576 69150 38734 69158
rect 38576 69146 38676 69150
rect 38948 69148 38980 69176
rect 39030 69148 39068 69176
rect 39110 69148 39142 69176
rect 38298 69120 38480 69146
rect 38702 69126 38762 69134
rect 38702 69122 38758 69126
rect 37176 69092 37210 69120
rect 37810 69094 37874 69120
rect 36274 69090 36303 69092
rect 36288 69086 36303 69090
rect 36485 69086 36500 69092
rect 36288 69076 36344 69086
rect 36198 69068 36204 69070
rect 33912 69046 34102 69050
rect 34104 69046 34412 69050
rect 33881 69031 33948 69046
rect 33896 69020 33948 69031
rect 34025 69020 34102 69046
rect 34140 69042 34173 69046
rect 33838 69016 33958 69020
rect 34025 69019 34138 69020
rect 34034 69018 34138 69019
rect 33836 69010 33958 69016
rect 34032 69010 34138 69018
rect 33826 69008 34138 69010
rect 33826 69002 34150 69008
rect 34172 69002 34173 69042
rect 34182 69002 34234 69032
rect 34298 69002 34330 69046
rect 34336 69024 34396 69046
rect 34332 69008 34386 69024
rect 34332 69002 34378 69008
rect 33826 68994 34159 69002
rect 33340 68766 33694 68988
rect 33826 68984 33948 68994
rect 33862 68978 33948 68984
rect 33954 68992 34159 68994
rect 33954 68978 34038 68992
rect 34082 68987 34159 68992
rect 34172 68990 34378 69002
rect 34082 68986 34150 68987
rect 34172 68986 34344 68990
rect 34066 68978 34344 68986
rect 33862 68976 34344 68978
rect 33860 68975 34344 68976
rect 34400 68975 34412 69046
rect 36294 69036 36344 69076
rect 36444 69076 36500 69086
rect 36924 69086 36939 69092
rect 36924 69076 36984 69086
rect 37838 69076 37874 69094
rect 36444 69036 36494 69076
rect 36934 69036 36984 69076
rect 37756 69052 37874 69076
rect 37892 69062 37928 69094
rect 38044 69062 38226 69120
rect 37892 69044 38226 69062
rect 33860 68974 34412 68975
rect 33860 68970 34178 68974
rect 33860 68966 34192 68970
rect 33860 68962 33868 68966
rect 33848 68950 33868 68962
rect 33912 68938 34018 68966
rect 34032 68956 34038 68966
rect 34054 68954 34192 68966
rect 33822 68902 33878 68916
rect 33912 68902 34014 68938
rect 34092 68934 34192 68954
rect 34282 68956 34344 68974
rect 34282 68946 34336 68956
rect 34352 68938 34398 68956
rect 34042 68902 34242 68934
rect 34380 68910 34426 68928
rect 36148 68902 36152 69016
rect 36176 68930 36180 69028
rect 36344 69016 36444 69026
rect 36704 69014 36804 69026
rect 36984 69016 37084 69026
rect 36590 69000 36602 69014
rect 37756 68998 37874 69022
rect 38044 69008 38226 69044
rect 37838 68952 37874 68998
rect 37892 68990 38226 69008
rect 37892 68952 37928 68990
rect 37810 68950 37874 68952
rect 36344 68932 36444 68942
rect 36704 68930 36804 68942
rect 36984 68932 37084 68942
rect 33912 68884 34092 68902
rect 34192 68884 34248 68902
rect 33912 68845 34056 68884
rect 34233 68869 34316 68884
rect 33912 68844 34092 68845
rect 34248 68844 34316 68869
rect 33912 68832 34316 68844
rect 36718 68838 36734 68856
rect 33822 68818 33878 68832
rect 33912 68800 33948 68832
rect 34030 68830 34316 68832
rect 34092 68818 34192 68830
rect 36958 68828 37004 68856
rect 37552 68828 37602 68856
rect 37892 68850 37934 68950
rect 38044 68866 38226 68990
rect 38298 69100 38810 69120
rect 39284 69110 39312 69146
rect 43290 69110 43318 69146
rect 38298 69064 38820 69100
rect 38876 69068 38904 69104
rect 38298 68916 38810 69064
rect 39284 69024 39312 69060
rect 38876 68982 38904 69018
rect 39356 68956 39388 68984
rect 39438 68958 39476 68986
rect 39518 68970 39522 68986
rect 39806 68978 40028 69026
rect 37810 68824 37874 68850
rect 33854 68786 33948 68800
rect 33912 68782 33948 68786
rect 33984 68784 34002 68786
rect 34040 68784 34140 68796
rect 33880 68772 33948 68782
rect 33978 68780 34040 68784
rect 33912 68764 33948 68772
rect 33976 68769 34040 68780
rect 34140 68776 34302 68784
rect 37838 68782 37874 68824
rect 34140 68775 34203 68776
rect 34140 68771 34202 68775
rect 37892 68774 37928 68824
rect 33976 68764 34038 68769
rect 33388 68738 33422 68752
rect 33912 68737 34102 68764
rect 34104 68737 34412 68764
rect 32784 68514 33138 68668
rect 33340 68500 33392 68734
rect 33440 68696 33496 68708
rect 33912 68700 34412 68737
rect 38298 68706 38480 68866
rect 38576 68762 38676 68774
rect 33912 68696 34102 68700
rect 34104 68696 34412 68700
rect 33881 68681 33948 68696
rect 33896 68670 33948 68681
rect 34025 68670 34102 68696
rect 34140 68692 34173 68696
rect 33838 68666 33958 68670
rect 34025 68669 34138 68670
rect 34034 68668 34138 68669
rect 33836 68660 33958 68666
rect 34032 68660 34138 68668
rect 33826 68658 34138 68660
rect 33826 68652 34150 68658
rect 34172 68652 34173 68692
rect 34182 68652 34234 68682
rect 34298 68652 34330 68696
rect 34336 68674 34396 68696
rect 34332 68658 34386 68674
rect 34332 68652 34378 68658
rect 33826 68644 34159 68652
rect 33826 68634 33948 68644
rect 33862 68628 33948 68634
rect 33954 68642 34159 68644
rect 33954 68628 34038 68642
rect 34082 68637 34159 68642
rect 34172 68640 34378 68652
rect 34082 68636 34150 68637
rect 34172 68636 34344 68640
rect 34066 68628 34344 68636
rect 33862 68626 34344 68628
rect 33860 68625 34344 68626
rect 34400 68625 34412 68696
rect 38776 68704 38810 68828
rect 38894 68786 38904 68800
rect 38576 68678 38676 68690
rect 38776 68682 38820 68704
rect 38702 68656 38758 68660
rect 38702 68648 38762 68656
rect 33860 68624 34412 68625
rect 33440 68612 33496 68624
rect 33860 68620 34178 68624
rect 33860 68616 34192 68620
rect 34282 68616 34344 68624
rect 38674 68620 38734 68632
rect 33860 68612 33868 68616
rect 33848 68600 33868 68612
rect 33912 68612 34018 68616
rect 34032 68612 34038 68616
rect 34054 68612 34192 68616
rect 34248 68612 34344 68616
rect 33912 68604 34398 68612
rect 33864 68586 33866 68600
rect 33912 68588 34072 68604
rect 34092 68588 34398 68604
rect 38298 68596 38702 68612
rect 38706 68590 38758 68598
rect 33912 68584 34014 68588
rect 34092 68584 34192 68588
rect 38378 68584 38418 68590
rect 38674 68584 38758 68590
rect 33836 68566 33866 68584
rect 33538 68552 33594 68564
rect 33822 68552 33878 68566
rect 33912 68560 34426 68584
rect 38270 68578 38758 68584
rect 38270 68568 38702 68578
rect 33912 68552 34014 68560
rect 34042 68552 34242 68560
rect 33912 68534 34092 68552
rect 34192 68534 34248 68552
rect 38674 68544 38696 68556
rect 38706 68536 38758 68578
rect 38776 68574 38810 68682
rect 38864 68576 39234 68740
rect 39370 68710 39388 68842
rect 39740 68792 40094 68978
rect 40378 68974 40418 68984
rect 40658 68968 40776 69038
rect 43290 69024 43318 69060
rect 46986 68998 47358 69240
rect 40592 68804 40842 68968
rect 41148 68956 41228 68984
rect 41364 68956 41444 68984
rect 41852 68956 41900 68984
rect 42174 68956 42250 68986
rect 42638 68956 42686 68984
rect 43042 68970 43060 68986
rect 43204 68958 43236 68986
rect 39342 68704 39416 68710
rect 39370 68690 39388 68704
rect 39388 68682 39538 68690
rect 39364 68674 39538 68682
rect 39364 68654 39392 68674
rect 38864 68572 39076 68576
rect 39090 68572 39234 68576
rect 38948 68566 38980 68572
rect 39004 68568 39234 68572
rect 39004 68566 39010 68568
rect 39030 68552 39234 68568
rect 33912 68500 34014 68534
rect 34030 68500 34056 68534
rect 34233 68519 34316 68534
rect 39052 68526 39058 68546
rect 39084 68542 39110 68552
rect 39084 68536 39100 68542
rect 34248 68500 34316 68519
rect 38674 68490 38792 68514
rect 33538 68468 33594 68480
rect 33822 68468 33878 68482
rect 34092 68468 34192 68480
rect 38702 68470 38764 68486
rect 38298 68452 38810 68470
rect 38298 68416 38820 68452
rect 38876 68420 38904 68456
rect 38298 68268 38810 68416
rect 39238 68386 39916 68528
rect 38876 68334 38904 68370
rect 39238 68362 40028 68386
rect 39238 68328 39324 68362
rect 39406 68360 40028 68362
rect 39406 68348 39508 68360
rect 39406 68330 39492 68348
rect 39442 68328 39492 68330
rect 28518 68198 28576 68226
rect 32598 68160 32674 68168
rect 32636 68158 32670 68160
rect 28638 68090 28890 68110
rect 28888 68084 28890 68090
rect 28948 68084 28952 68110
rect 28666 68062 28890 68082
rect 28860 68056 28890 68062
rect 28948 68056 28980 68082
rect 28800 67950 28808 67992
rect 28828 67922 28836 67972
rect 28866 67908 28892 67972
rect 28894 67880 28920 68000
rect 29044 67988 29068 68088
rect 29072 68016 29096 68060
rect 29114 68016 29136 68060
rect 29072 67996 29136 68016
rect 29072 67994 29134 67996
rect 29142 67988 29164 68088
rect 29044 67968 29164 67988
rect 29174 67988 29194 68088
rect 32626 68076 32654 68140
rect 32776 68088 33130 68238
rect 33374 68164 33436 68192
rect 33442 68184 33464 68204
rect 36694 68188 36744 68212
rect 34240 68152 34298 68180
rect 36702 68170 36740 68188
rect 36964 68168 37010 68196
rect 37106 68162 37172 68178
rect 37094 68134 37144 68150
rect 38576 68112 38676 68124
rect 38876 68114 38904 68150
rect 39406 68106 39492 68328
rect 39522 68320 39536 68360
rect 39638 68348 39670 68360
rect 39806 68352 40028 68360
rect 40462 68362 40538 68510
rect 39806 68336 40066 68352
rect 40462 68342 40630 68362
rect 39806 68324 40028 68336
rect 39806 68322 40038 68324
rect 39740 68284 40094 68322
rect 40658 68318 40776 68390
rect 41268 68362 41348 68502
rect 41348 68334 41436 68362
rect 39740 68258 40318 68284
rect 39740 68256 40094 68258
rect 39740 68230 40318 68256
rect 39740 68152 40094 68230
rect 40592 68156 40842 68318
rect 41930 68114 42012 68130
rect 36350 68094 36450 68104
rect 36710 68094 36810 68106
rect 36990 68094 37090 68104
rect 33078 68070 33130 68088
rect 29202 68016 29222 68060
rect 33904 68020 33940 68088
rect 34032 68022 34132 68034
rect 36598 68022 36608 68036
rect 29202 67994 29264 68016
rect 33872 68010 33940 68020
rect 36350 68010 36450 68020
rect 36710 68010 36810 68022
rect 36990 68010 37090 68020
rect 33904 68002 33940 68010
rect 29044 67966 29162 67968
rect 29174 67966 29292 67988
rect 33904 67975 34094 68002
rect 34096 67975 34404 68002
rect 29224 67904 29248 67950
rect 28666 67678 28716 67722
rect 29278 67718 29302 67904
rect 32626 67726 32654 67790
rect 32776 67752 33130 67888
rect 32824 67738 32872 67752
rect 33078 67720 33130 67752
rect 33332 67876 33384 67972
rect 33432 67934 33488 67946
rect 33904 67938 34404 67975
rect 36204 67966 36210 67968
rect 36186 67944 36210 67966
rect 36300 67960 36350 68000
rect 36294 67950 36350 67960
rect 36450 67960 36500 68000
rect 36940 67960 36990 68000
rect 36450 67950 36506 67960
rect 36294 67946 36309 67950
rect 33904 67934 34094 67938
rect 34096 67934 34404 67938
rect 33873 67919 33940 67934
rect 33888 67908 33940 67919
rect 34017 67908 34094 67934
rect 34132 67930 34165 67934
rect 33830 67904 33950 67908
rect 34017 67907 34130 67908
rect 34026 67906 34130 67907
rect 33828 67898 33950 67904
rect 34024 67898 34130 67906
rect 33818 67896 34130 67898
rect 33818 67890 34142 67896
rect 34164 67890 34165 67930
rect 34174 67890 34226 67920
rect 34290 67890 34322 67934
rect 34328 67912 34388 67934
rect 34324 67896 34378 67912
rect 34324 67890 34370 67896
rect 33818 67882 34151 67890
rect 28728 67654 28744 67706
rect 33332 67654 33686 67876
rect 33818 67872 33940 67882
rect 33854 67866 33940 67872
rect 33946 67880 34151 67882
rect 33946 67866 34030 67880
rect 34074 67875 34151 67880
rect 34164 67878 34370 67890
rect 34074 67874 34142 67875
rect 34164 67874 34336 67878
rect 34058 67866 34336 67874
rect 33854 67864 34336 67866
rect 33852 67863 34336 67864
rect 34392 67863 34404 67934
rect 36174 67932 36210 67944
rect 36280 67944 36309 67946
rect 36491 67944 36506 67950
rect 36930 67950 36990 67960
rect 36930 67944 36945 67950
rect 36218 67934 36238 67940
rect 36144 67918 36212 67932
rect 36218 67928 36260 67934
rect 36174 67904 36208 67918
rect 36144 67890 36212 67904
rect 36218 67894 36242 67928
rect 36246 67894 36260 67928
rect 36280 67912 36354 67944
rect 36446 67912 36996 67944
rect 37102 67914 37136 67942
rect 37182 67916 37216 67944
rect 37260 67914 37724 68078
rect 38576 68028 38676 68040
rect 38792 68032 38820 68068
rect 38876 68028 38904 68064
rect 38702 68006 38758 68010
rect 38702 67998 38762 68006
rect 38764 67998 38774 68026
rect 38432 67974 38532 67986
rect 38576 67982 38676 67986
rect 38746 67982 38762 67998
rect 38576 67974 38734 67982
rect 38674 67970 38734 67974
rect 38718 67954 38734 67970
rect 38746 67966 38792 67982
rect 38948 67954 38980 67982
rect 39030 67954 39068 67982
rect 39110 67954 39142 67982
rect 39236 67976 39324 68060
rect 39404 67976 39492 68106
rect 39942 68074 39956 68092
rect 39970 68090 39984 68114
rect 39960 68074 39984 68090
rect 41896 68108 42012 68114
rect 42016 68108 42118 68114
rect 41896 68090 42118 68108
rect 41896 68066 41904 68090
rect 41930 68086 42056 68090
rect 41924 68078 42146 68086
rect 41924 68062 41982 68078
rect 41924 68038 41928 68062
rect 41930 68036 41982 68062
rect 41998 68062 42146 68078
rect 41998 68050 42056 68062
rect 41998 68036 42013 68050
rect 41930 68030 41990 68036
rect 41924 68028 41990 68030
rect 41992 68032 42024 68036
rect 41924 68022 41988 68028
rect 41924 68020 41986 68022
rect 41924 68000 41986 68002
rect 41924 67994 41988 68000
rect 41992 67994 42044 68032
rect 41924 67992 42044 67994
rect 41416 67980 41418 67992
rect 41930 67990 42044 67992
rect 42110 67990 42144 68032
rect 42222 67990 42256 68032
rect 42336 67990 42370 68032
rect 42404 67990 42438 68032
rect 41930 67986 42024 67990
rect 38718 67938 38764 67954
rect 37558 67910 37608 67914
rect 36174 67878 36210 67890
rect 36218 67888 36260 67894
rect 36218 67882 36238 67888
rect 33852 67862 34404 67863
rect 33852 67858 34170 67862
rect 33852 67854 34184 67858
rect 33852 67850 33860 67854
rect 33840 67838 33860 67850
rect 33904 67826 34010 67854
rect 34024 67844 34030 67854
rect 34046 67842 34184 67854
rect 33814 67790 33870 67804
rect 33904 67790 34006 67826
rect 34084 67822 34184 67842
rect 34274 67844 34336 67862
rect 36186 67856 36210 67878
rect 36280 67878 36354 67910
rect 36446 67878 36996 67910
rect 37182 67878 37216 67906
rect 38432 67890 38532 67902
rect 38576 67890 38676 67902
rect 39236 67892 39302 67976
rect 39404 67914 39470 67976
rect 41580 67940 41602 67964
rect 41608 67936 41630 67940
rect 41896 67936 41904 67956
rect 41924 67936 41928 67984
rect 41930 67972 42013 67986
rect 41930 67942 42056 67972
rect 41960 67914 42056 67942
rect 36280 67876 36309 67878
rect 36294 67872 36309 67876
rect 36491 67872 36506 67878
rect 36294 67862 36350 67872
rect 36204 67854 36210 67856
rect 34274 67834 34328 67844
rect 34344 67826 34390 67844
rect 36300 67822 36350 67862
rect 36450 67862 36506 67872
rect 36930 67872 36945 67878
rect 36930 67862 36990 67872
rect 36450 67822 36500 67862
rect 36940 67822 36990 67862
rect 39404 67852 39492 67914
rect 41960 67892 42012 67914
rect 34034 67790 34234 67822
rect 34372 67798 34418 67816
rect 36350 67802 36450 67812
rect 36710 67800 36810 67812
rect 36990 67802 37090 67812
rect 33904 67772 34084 67790
rect 34184 67772 34240 67790
rect 36596 67786 36608 67800
rect 33904 67733 34048 67772
rect 34225 67757 34308 67772
rect 33904 67732 34084 67733
rect 34240 67732 34308 67757
rect 33904 67720 34308 67732
rect 33814 67706 33870 67720
rect 33904 67688 33940 67720
rect 34022 67718 34308 67720
rect 36350 67718 36450 67728
rect 34084 67706 34184 67718
rect 33846 67674 33940 67688
rect 33904 67670 33940 67674
rect 33976 67672 33994 67674
rect 34032 67672 34132 67684
rect 33872 67660 33940 67670
rect 33970 67668 34032 67672
rect 33904 67652 33940 67660
rect 33968 67657 34032 67668
rect 34132 67664 34294 67672
rect 34132 67663 34195 67664
rect 34132 67659 34194 67663
rect 36576 67662 37260 67774
rect 33968 67652 34030 67657
rect 29180 67636 29194 67640
rect 28846 67610 28856 67611
rect 28764 67576 28798 67596
rect 28710 67560 28740 67564
rect 28744 67530 28774 67560
rect 28778 67528 28784 67576
rect 28806 67556 28812 67604
rect 28846 67596 28861 67610
rect 29180 67598 29248 67636
rect 33380 67626 33428 67640
rect 33904 67625 34094 67652
rect 34096 67625 34404 67652
rect 29180 67596 29194 67598
rect 29208 67596 29248 67598
rect 28846 67566 28902 67596
rect 29116 67566 29140 67596
rect 29180 67566 29248 67596
rect 29370 67576 29398 67622
rect 28846 67551 28861 67566
rect 29180 67542 29194 67566
rect 29208 67548 29282 67566
rect 29233 67542 29248 67548
rect 28794 67524 28804 67540
rect 28846 67538 28902 67539
rect 28846 67524 29010 67538
rect 29101 67524 29140 67539
rect 29180 67526 29248 67542
rect 29180 67520 29262 67526
rect 29182 67506 29194 67520
rect 28780 67494 28916 67502
rect 29182 67484 29202 67506
rect 29210 67494 29230 67504
rect 29210 67492 29272 67494
rect 29210 67484 29230 67492
rect 29182 67448 29204 67484
rect 29182 67442 29202 67448
rect 28666 67370 28716 67414
rect 29182 67412 29194 67442
rect 29210 67440 29232 67484
rect 28728 67344 28744 67396
rect 28802 67214 28810 67218
rect 28528 67184 28540 67211
rect 28528 67130 28543 67184
rect 28802 67172 28816 67214
rect 28528 67116 28540 67130
rect 28802 67116 28810 67172
rect 28834 67144 28844 67196
rect 29244 67188 29260 67444
rect 29280 67224 29296 67408
rect 28836 67138 28844 67144
rect 28528 67075 28543 67116
rect 29372 67080 29428 67474
rect 32626 67376 32654 67440
rect 32776 67402 33130 67538
rect 32824 67388 32872 67402
rect 33078 67370 33130 67402
rect 33332 67526 33384 67622
rect 33432 67584 33488 67596
rect 33904 67588 34404 67625
rect 33904 67584 34094 67588
rect 34096 67584 34404 67588
rect 33873 67569 33940 67584
rect 33888 67558 33940 67569
rect 34017 67558 34094 67584
rect 34132 67580 34165 67584
rect 33830 67554 33950 67558
rect 34017 67557 34130 67558
rect 34026 67556 34130 67557
rect 33828 67548 33950 67554
rect 34024 67548 34130 67556
rect 33818 67546 34130 67548
rect 33818 67540 34142 67546
rect 34164 67540 34165 67580
rect 34174 67540 34226 67570
rect 34290 67540 34322 67584
rect 34328 67562 34388 67584
rect 34324 67546 34378 67562
rect 34324 67540 34370 67546
rect 33818 67532 34151 67540
rect 33332 67304 33686 67526
rect 33818 67522 33940 67532
rect 33854 67516 33940 67522
rect 33946 67530 34151 67532
rect 33946 67516 34030 67530
rect 34074 67525 34151 67530
rect 34164 67528 34370 67540
rect 34074 67524 34142 67525
rect 34164 67524 34336 67528
rect 34058 67516 34336 67524
rect 33854 67514 34336 67516
rect 33852 67513 34336 67514
rect 34392 67513 34404 67584
rect 33852 67512 34404 67513
rect 33852 67508 34170 67512
rect 33852 67504 34184 67508
rect 33852 67500 33860 67504
rect 33840 67488 33860 67500
rect 33904 67476 34010 67504
rect 34024 67494 34030 67504
rect 34046 67492 34184 67504
rect 33814 67440 33870 67454
rect 33904 67440 34006 67476
rect 34084 67472 34184 67492
rect 34274 67494 34336 67512
rect 34274 67484 34328 67494
rect 34344 67476 34390 67494
rect 34034 67440 34234 67472
rect 34372 67448 34418 67466
rect 36350 67454 36450 67464
rect 36710 67454 36810 67466
rect 36990 67454 37090 67464
rect 33904 67422 34084 67440
rect 34184 67422 34240 67440
rect 33904 67383 34048 67422
rect 34225 67407 34308 67422
rect 33904 67382 34084 67383
rect 34240 67382 34308 67407
rect 33904 67370 34308 67382
rect 36350 67370 36450 67380
rect 36710 67370 36810 67382
rect 36990 67370 37090 67380
rect 33814 67356 33870 67370
rect 33904 67338 33940 67370
rect 34022 67368 34308 67370
rect 34084 67356 34184 67368
rect 33846 67324 33940 67338
rect 33904 67320 33940 67324
rect 33976 67322 33994 67324
rect 34032 67322 34132 67334
rect 36204 67326 36210 67328
rect 33872 67310 33940 67320
rect 33970 67318 34032 67322
rect 33904 67302 33940 67310
rect 33968 67307 34032 67318
rect 34132 67314 34294 67322
rect 34132 67313 34195 67314
rect 34132 67309 34194 67313
rect 33968 67302 34030 67307
rect 36186 67304 36210 67326
rect 36300 67320 36350 67360
rect 36294 67310 36350 67320
rect 36450 67320 36500 67360
rect 36940 67320 36990 67360
rect 36450 67310 36506 67320
rect 36294 67306 36309 67310
rect 33380 67276 33428 67290
rect 33904 67275 34094 67302
rect 34096 67275 34404 67302
rect 36174 67292 36210 67304
rect 36280 67304 36309 67306
rect 36491 67304 36506 67310
rect 36930 67310 36990 67320
rect 36930 67304 36945 67310
rect 36218 67294 36238 67300
rect 36144 67278 36212 67292
rect 36218 67288 36260 67294
rect 28528 67000 28545 67075
rect 29040 67016 29058 67060
rect 28528 66972 28564 67000
rect 29068 66988 29086 67040
rect 29114 66976 29132 67040
rect 28492 66946 28564 66972
rect 29142 66948 29160 67068
rect 28510 66932 28564 66946
rect 29182 66936 29194 67056
rect 29210 66964 29222 67028
rect 32626 67026 32654 67090
rect 32776 67052 33130 67188
rect 33078 67020 33130 67052
rect 33332 67176 33384 67272
rect 33432 67234 33488 67246
rect 33904 67238 34404 67275
rect 36174 67264 36208 67278
rect 36144 67250 36212 67264
rect 36218 67254 36242 67288
rect 36246 67254 36260 67288
rect 36280 67272 36354 67304
rect 36446 67272 36996 67304
rect 37102 67274 37136 67302
rect 37182 67276 37216 67304
rect 37260 67272 37724 67438
rect 39260 67412 39312 67414
rect 39298 67386 39314 67396
rect 39288 67384 39314 67386
rect 39298 67372 39314 67384
rect 37558 67270 37608 67272
rect 36174 67238 36210 67250
rect 36218 67248 36260 67254
rect 36218 67242 36238 67248
rect 33904 67234 34094 67238
rect 34096 67234 34404 67238
rect 33873 67219 33940 67234
rect 33888 67208 33940 67219
rect 34017 67208 34094 67234
rect 34132 67230 34165 67234
rect 33830 67204 33950 67208
rect 34017 67207 34130 67208
rect 34026 67206 34130 67207
rect 33828 67198 33950 67204
rect 34024 67198 34130 67206
rect 33818 67196 34130 67198
rect 33818 67190 34142 67196
rect 34164 67190 34165 67230
rect 34174 67190 34226 67220
rect 34290 67190 34322 67234
rect 34328 67212 34388 67234
rect 34324 67196 34378 67212
rect 34324 67190 34370 67196
rect 33818 67182 34151 67190
rect 33332 66954 33686 67176
rect 33818 67172 33940 67182
rect 33854 67166 33940 67172
rect 33946 67180 34151 67182
rect 33946 67166 34030 67180
rect 34074 67175 34151 67180
rect 34164 67178 34370 67190
rect 34074 67174 34142 67175
rect 34164 67174 34336 67178
rect 34058 67166 34336 67174
rect 33854 67164 34336 67166
rect 33852 67163 34336 67164
rect 34392 67163 34404 67234
rect 36186 67216 36210 67238
rect 36280 67238 36354 67270
rect 36446 67238 36996 67270
rect 37182 67238 37216 67266
rect 36280 67236 36309 67238
rect 36294 67232 36309 67236
rect 36491 67232 36506 67238
rect 36294 67222 36350 67232
rect 36204 67214 36210 67216
rect 33852 67162 34404 67163
rect 35970 67162 36216 67194
rect 36300 67182 36350 67222
rect 36450 67222 36506 67232
rect 36930 67232 36945 67238
rect 36930 67222 36990 67232
rect 39382 67226 39386 67228
rect 39406 67226 39492 67852
rect 39942 67750 39992 67766
rect 39942 67746 39976 67750
rect 39970 67722 40020 67738
rect 39970 67718 40004 67722
rect 41896 67714 41942 67754
rect 42148 67714 42194 67756
rect 41930 67560 42012 67576
rect 41896 67554 42012 67560
rect 42016 67554 42118 67560
rect 41896 67536 42118 67554
rect 41896 67512 41904 67536
rect 41930 67532 42056 67536
rect 41924 67524 42146 67532
rect 41924 67508 41982 67524
rect 41924 67484 41928 67508
rect 41930 67482 41982 67508
rect 41998 67508 42146 67524
rect 41998 67500 42122 67508
rect 41998 67496 42056 67500
rect 41998 67482 42013 67496
rect 42040 67492 42046 67496
rect 42084 67492 42086 67500
rect 42084 67490 42088 67492
rect 42084 67488 42092 67490
rect 41930 67474 41990 67482
rect 41992 67478 42024 67482
rect 42028 67478 42094 67488
rect 42112 67478 42120 67500
rect 41924 67468 41988 67474
rect 41992 67472 42094 67478
rect 41924 67442 41988 67446
rect 41992 67442 42044 67472
rect 42084 67442 42092 67472
rect 41924 67440 42094 67442
rect 41930 67436 42094 67440
rect 42110 67436 42144 67478
rect 42222 67436 42256 67478
rect 42336 67436 42370 67478
rect 42404 67436 42438 67478
rect 41930 67432 42024 67436
rect 41896 67382 41904 67402
rect 41924 67382 41928 67430
rect 41930 67418 42013 67432
rect 42028 67430 42094 67436
rect 42084 67426 42092 67430
rect 41930 67414 42056 67418
rect 42112 67414 42120 67436
rect 41930 67402 42122 67414
rect 41930 67388 42056 67402
rect 42112 67398 42120 67402
rect 41960 67360 42056 67388
rect 41960 67338 42012 67360
rect 36450 67182 36500 67222
rect 36940 67182 36990 67222
rect 39376 67188 39386 67226
rect 39404 67216 39492 67226
rect 36350 67162 36450 67172
rect 33852 67158 34170 67162
rect 33852 67154 34184 67158
rect 33852 67150 33860 67154
rect 33840 67138 33860 67150
rect 33904 67126 34010 67154
rect 34024 67144 34030 67154
rect 34046 67142 34184 67154
rect 33814 67090 33870 67104
rect 33904 67090 34006 67126
rect 34084 67122 34184 67142
rect 34274 67144 34336 67162
rect 34274 67134 34328 67144
rect 34344 67126 34390 67144
rect 34034 67090 34234 67122
rect 34372 67098 34418 67116
rect 33904 67072 34084 67090
rect 34184 67072 34240 67090
rect 33904 67033 34048 67072
rect 34225 67057 34308 67072
rect 33904 67032 34084 67033
rect 34240 67032 34308 67057
rect 35970 67032 36224 67162
rect 36710 67160 36810 67172
rect 36990 67162 37090 67172
rect 39382 67164 39386 67188
rect 36596 67146 36608 67160
rect 39406 67154 39492 67216
rect 39410 67136 39414 67154
rect 40462 67152 40538 67180
rect 41788 67152 41834 67202
rect 42040 67152 42086 67202
rect 36350 67078 36450 67088
rect 36710 67076 36810 67088
rect 36990 67078 37090 67088
rect 33904 67020 34308 67032
rect 33814 67006 33870 67020
rect 33904 66988 33940 67020
rect 34022 67018 34308 67020
rect 34084 67006 34184 67018
rect 33846 66974 33940 66988
rect 33904 66970 33940 66974
rect 33976 66972 33994 66974
rect 34032 66972 34132 66984
rect 36964 66974 37010 67002
rect 33872 66960 33940 66970
rect 33970 66968 34032 66972
rect 33904 66952 33940 66960
rect 33968 66957 34032 66968
rect 34132 66964 34294 66972
rect 34132 66963 34195 66964
rect 34132 66959 34194 66963
rect 33968 66952 34030 66957
rect 28510 66896 28536 66932
rect 33380 66926 33422 66940
rect 33904 66925 34094 66952
rect 34096 66925 34404 66952
rect 37530 66946 37550 67016
rect 37558 66974 37608 67002
rect 32776 66702 33130 66856
rect 33332 66688 33384 66922
rect 33432 66884 33488 66896
rect 33904 66888 34404 66925
rect 33904 66884 34094 66888
rect 34096 66884 34404 66888
rect 33873 66869 33940 66884
rect 33888 66858 33940 66869
rect 34017 66858 34094 66884
rect 34132 66880 34165 66884
rect 33830 66854 33950 66858
rect 34017 66857 34130 66858
rect 34026 66856 34130 66857
rect 33828 66848 33950 66854
rect 34024 66848 34130 66856
rect 33818 66846 34130 66848
rect 33818 66840 34142 66846
rect 34164 66840 34165 66880
rect 34174 66840 34226 66870
rect 34290 66840 34322 66884
rect 34328 66862 34388 66884
rect 34324 66846 34378 66862
rect 34324 66840 34370 66846
rect 33818 66832 34151 66840
rect 33818 66822 33940 66832
rect 33854 66816 33940 66822
rect 33946 66830 34151 66832
rect 33946 66816 34030 66830
rect 34074 66825 34151 66830
rect 34164 66828 34370 66840
rect 34074 66824 34142 66825
rect 34164 66824 34336 66828
rect 34058 66816 34336 66824
rect 33854 66814 34336 66816
rect 33852 66813 34336 66814
rect 34392 66813 34404 66884
rect 33852 66812 34404 66813
rect 33432 66800 33488 66812
rect 33852 66808 34170 66812
rect 33852 66804 34184 66808
rect 34274 66804 34336 66812
rect 33852 66800 33860 66804
rect 33840 66788 33860 66800
rect 33904 66776 34010 66804
rect 34024 66794 34030 66804
rect 34046 66792 34184 66804
rect 34240 66794 34336 66804
rect 33530 66740 33586 66752
rect 33814 66740 33870 66754
rect 33904 66740 34006 66776
rect 34084 66772 34184 66792
rect 34274 66790 34328 66794
rect 34240 66784 34328 66790
rect 34240 66776 34278 66784
rect 34034 66762 34234 66772
rect 34034 66748 34278 66762
rect 34034 66740 34234 66748
rect 33904 66722 34084 66740
rect 34184 66722 34240 66740
rect 33904 66688 34006 66722
rect 34022 66688 34048 66722
rect 34225 66707 34308 66722
rect 34240 66688 34308 66707
rect 33530 66656 33586 66668
rect 33814 66656 33870 66670
rect 34084 66656 34184 66668
rect 34250 66660 34270 66688
rect 27794 66588 27796 66620
rect 27828 66604 27830 66642
rect 27987 66600 28002 66615
rect 27836 66570 27894 66600
rect 27946 66570 28002 66600
rect 28014 66588 28016 66620
rect 28048 66604 28050 66640
rect 28114 66620 28126 66630
rect 28234 66570 28236 66620
rect 28268 66604 28270 66640
rect 28334 66620 28346 66630
rect 27987 66555 28002 66570
rect 37092 66540 37114 66568
rect 37258 66540 37280 66568
rect 35076 66472 35124 66536
rect 35324 66472 35372 66536
rect 37038 66476 37086 66540
rect 37286 66476 37334 66540
rect 27454 66442 27506 66472
rect 27564 66442 27616 66472
rect 27674 66442 27726 66472
rect 27784 66442 27836 66472
rect 27894 66442 27946 66472
rect 35076 66204 35124 66268
rect 35324 66202 35372 66266
rect 37038 66208 37086 66272
rect 37286 66206 37334 66270
rect 27987 66044 28002 66059
rect 27836 66014 27894 66044
rect 27946 66014 28002 66044
rect 27987 65999 28002 66014
rect 38252 65964 38448 65992
rect 38252 65954 38267 65964
rect 36120 65948 36138 65954
rect 36230 65948 36248 65954
rect 38252 65952 38286 65954
rect 34294 65922 34344 65934
rect 34396 65922 34454 65934
rect 34506 65922 34564 65934
rect 34616 65922 34666 65934
rect 35782 65922 35832 65934
rect 35884 65922 35942 65934
rect 35994 65928 36044 65934
rect 36162 65928 36180 65948
rect 36272 65928 36290 65948
rect 36358 65928 36416 65940
rect 36468 65928 36526 65940
rect 36578 65928 36628 65940
rect 37744 65928 37794 65940
rect 37846 65928 37904 65940
rect 37956 65928 38014 65940
rect 38066 65928 38116 65940
rect 38252 65928 38296 65952
rect 35994 65922 36028 65928
rect 36037 65922 36086 65928
rect 36147 65922 36196 65928
rect 36257 65924 36306 65928
rect 36619 65924 36634 65928
rect 34657 65918 34672 65922
rect 34292 65884 34344 65918
rect 34396 65884 34454 65918
rect 34506 65884 34564 65918
rect 34616 65884 34672 65918
rect 35776 65918 35791 65922
rect 36037 65918 36052 65922
rect 36147 65918 36180 65922
rect 27702 65458 27716 65578
rect 27740 65550 27784 65634
rect 27730 65486 27784 65550
rect 28380 65536 28410 65604
rect 28470 65550 28478 65583
rect 28494 65562 28516 65604
rect 28536 65536 28558 65562
rect 28368 65521 28531 65536
rect 27740 65312 27784 65486
rect 28380 65516 28516 65521
rect 28380 65462 28426 65516
rect 28472 65490 28516 65516
rect 28472 65482 28553 65490
rect 28478 65462 28516 65482
rect 27616 65058 27784 65312
rect 27802 65106 27804 65108
rect 27702 64904 27716 65024
rect 27740 64996 27784 65058
rect 27802 65032 27804 65070
rect 27814 65058 27816 65218
rect 27902 65108 27912 65118
rect 28004 65084 28070 65312
rect 28122 65108 28132 65118
rect 28004 65080 28084 65084
rect 27912 65058 27914 65074
rect 27814 65050 27982 65058
rect 28004 65050 28096 65080
rect 27912 65032 27914 65050
rect 28016 65032 28024 65050
rect 28040 65044 28056 65050
rect 28064 65044 28084 65050
rect 28040 65035 28055 65044
rect 28098 65038 28118 65084
rect 28126 65038 28132 65108
rect 28160 65080 28166 65142
rect 28176 65140 28194 65142
rect 28174 65080 28194 65140
rect 28210 65106 28228 65108
rect 28148 65050 28206 65080
rect 28160 65044 28166 65050
rect 28174 65044 28194 65050
rect 28208 65040 28228 65106
rect 28210 65038 28228 65040
rect 28236 65106 28244 65108
rect 28236 65074 28242 65106
rect 28270 65080 28276 65128
rect 28342 65108 28352 65118
rect 28284 65080 28304 65084
rect 28236 65038 28244 65074
rect 28258 65050 28316 65080
rect 28270 65044 28276 65050
rect 28284 65044 28304 65050
rect 28318 65038 28338 65084
rect 28346 65072 28352 65108
rect 28380 65080 28420 65462
rect 34292 65435 34330 65884
rect 34657 65869 34672 65884
rect 34968 65720 34984 65726
rect 34968 65712 34986 65720
rect 34968 65676 34988 65712
rect 34968 65662 34984 65676
rect 34996 65634 35012 65754
rect 35018 65746 35020 65750
rect 35018 65704 35022 65746
rect 35048 65716 35058 65742
rect 35096 65714 35140 65896
rect 35428 65746 35430 65750
rect 35390 65716 35400 65740
rect 35076 65650 35140 65714
rect 35096 65594 35140 65650
rect 35324 65648 35372 65712
rect 35426 65704 35430 65746
rect 35436 65634 35452 65754
rect 35476 65726 35520 65896
rect 35776 65884 35832 65918
rect 35884 65884 35942 65918
rect 35994 65884 36086 65918
rect 36138 65913 36162 65918
rect 36138 65885 36156 65913
rect 35776 65869 35791 65884
rect 36052 65880 36074 65884
rect 36006 65862 36074 65880
rect 36105 65880 36156 65885
rect 36162 65880 36184 65891
rect 36254 65890 36306 65924
rect 36358 65890 36416 65924
rect 36468 65890 36526 65924
rect 36578 65890 36634 65924
rect 37738 65924 37753 65928
rect 36105 65874 36184 65880
rect 36215 65880 36248 65885
rect 36254 65880 36294 65890
rect 36215 65874 36294 65880
rect 36325 65880 36358 65885
rect 36325 65874 36404 65880
rect 36619 65875 36634 65890
rect 36006 65846 36085 65862
rect 36116 65846 36184 65874
rect 36226 65846 36294 65874
rect 36336 65846 36404 65874
rect 36006 65840 36040 65846
rect 36116 65840 36156 65846
rect 36226 65840 36292 65846
rect 36336 65840 36370 65846
rect 36052 65812 36085 65823
rect 36138 65817 36156 65840
rect 36254 65823 36292 65840
rect 36006 65810 36085 65812
rect 36105 65812 36156 65817
rect 36162 65812 36184 65823
rect 36006 65778 36074 65810
rect 36105 65806 36184 65812
rect 36215 65812 36248 65817
rect 36254 65812 36294 65823
rect 36215 65806 36294 65812
rect 36325 65812 36358 65817
rect 36325 65806 36404 65812
rect 36116 65778 36184 65806
rect 36226 65778 36294 65806
rect 36336 65778 36404 65806
rect 36006 65772 36040 65778
rect 36116 65772 36156 65778
rect 36226 65772 36292 65778
rect 36336 65772 36370 65778
rect 36052 65744 36074 65755
rect 36138 65749 36156 65772
rect 36254 65755 36292 65772
rect 35464 65720 35520 65726
rect 35462 65712 35520 65720
rect 35460 65676 35520 65712
rect 36006 65710 36074 65744
rect 36105 65744 36156 65749
rect 36162 65744 36184 65755
rect 36105 65738 36184 65744
rect 36215 65744 36248 65749
rect 36254 65744 36294 65755
rect 36215 65738 36294 65744
rect 36325 65744 36358 65749
rect 36325 65738 36404 65744
rect 36116 65710 36184 65738
rect 36226 65710 36294 65738
rect 36336 65710 36404 65738
rect 36930 65726 36946 65732
rect 36930 65718 36948 65726
rect 36006 65704 36040 65710
rect 36116 65704 36156 65710
rect 36226 65704 36292 65710
rect 36336 65704 36370 65710
rect 36052 65676 36074 65687
rect 36138 65681 36156 65704
rect 36254 65687 36292 65704
rect 35464 65662 35520 65676
rect 35476 65594 35520 65662
rect 36006 65642 36074 65676
rect 36105 65676 36156 65681
rect 36162 65676 36184 65687
rect 36105 65670 36184 65676
rect 36215 65676 36248 65681
rect 36254 65676 36294 65687
rect 36930 65682 36950 65718
rect 36215 65670 36294 65676
rect 36325 65676 36358 65681
rect 36325 65670 36404 65676
rect 36116 65642 36184 65670
rect 36226 65642 36294 65670
rect 36336 65642 36404 65670
rect 36930 65668 36946 65682
rect 36006 65636 36040 65642
rect 36116 65636 36156 65642
rect 36226 65636 36292 65642
rect 36336 65636 36370 65642
rect 36958 65640 36974 65760
rect 36980 65752 36982 65756
rect 36980 65710 36984 65752
rect 37010 65722 37020 65746
rect 37058 65718 37102 65902
rect 37390 65752 37392 65756
rect 37352 65722 37362 65746
rect 37038 65654 37102 65718
rect 37286 65654 37334 65718
rect 37388 65710 37392 65752
rect 36052 65608 36074 65619
rect 36138 65613 36156 65636
rect 36254 65619 36292 65636
rect 34286 65424 34344 65435
rect 34124 65394 34176 65424
rect 34234 65420 34396 65424
rect 34234 65394 34286 65420
rect 34292 65382 34330 65420
rect 34344 65394 34396 65420
rect 34454 65394 34506 65424
rect 34564 65394 34616 65424
rect 34452 65382 34460 65384
rect 34642 65382 34708 65594
rect 34896 65382 34898 65500
rect 34972 65458 35140 65594
rect 34968 65394 35140 65458
rect 34972 65382 35140 65394
rect 34292 65360 34328 65382
rect 34344 65360 34372 65382
rect 34452 65364 35140 65382
rect 34292 65356 34372 65360
rect 34286 65342 34344 65356
rect 34360 65342 34366 65356
rect 34374 65342 34394 65358
rect 34396 65356 34454 65360
rect 34424 65354 34432 65356
rect 34470 65354 34476 65358
rect 34484 65354 34504 65358
rect 34506 65356 34564 65360
rect 34580 65354 34586 65364
rect 34594 65354 34614 65364
rect 34642 65360 34708 65364
rect 34616 65356 34708 65360
rect 34642 65354 34708 65356
rect 34722 65354 34724 65358
rect 34832 65354 34834 65358
rect 34896 65354 34898 65364
rect 34942 65354 34944 65358
rect 34972 65354 35140 65364
rect 34424 65346 35140 65354
rect 34408 65342 35140 65346
rect 34286 65341 35140 65342
rect 28346 65038 28354 65072
rect 28368 65050 28420 65080
rect 28380 65049 28420 65050
rect 34292 65340 34332 65341
rect 34338 65340 35140 65341
rect 35352 65488 35520 65594
rect 35550 65488 35552 65500
rect 35740 65488 35806 65594
rect 36006 65574 36074 65608
rect 36105 65608 36156 65613
rect 36162 65608 36184 65619
rect 36105 65602 36184 65608
rect 36215 65608 36248 65613
rect 36254 65608 36294 65619
rect 36215 65602 36294 65608
rect 36325 65608 36358 65613
rect 36325 65602 36404 65608
rect 36116 65574 36184 65602
rect 36226 65574 36294 65602
rect 36336 65574 36404 65602
rect 37058 65600 37102 65654
rect 37398 65640 37414 65760
rect 37438 65732 37482 65902
rect 37738 65890 37794 65924
rect 37846 65890 37904 65924
rect 37956 65890 38014 65924
rect 38066 65890 38118 65924
rect 38252 65917 38344 65928
rect 38251 65906 38344 65917
rect 37738 65875 37753 65890
rect 37426 65726 37482 65732
rect 37424 65718 37482 65726
rect 37422 65682 37482 65718
rect 37426 65668 37482 65682
rect 37438 65600 37482 65668
rect 36006 65568 36040 65574
rect 36116 65568 36156 65574
rect 36226 65568 36292 65574
rect 36336 65568 36370 65574
rect 36052 65540 36074 65551
rect 36138 65545 36156 65568
rect 36254 65551 36292 65568
rect 36006 65506 36074 65540
rect 36105 65540 36156 65545
rect 36162 65540 36184 65551
rect 36105 65534 36184 65540
rect 36215 65540 36248 65545
rect 36254 65540 36294 65551
rect 36215 65534 36294 65540
rect 36325 65540 36358 65545
rect 36325 65534 36404 65540
rect 36116 65506 36184 65534
rect 36226 65506 36294 65534
rect 36336 65506 36404 65534
rect 36006 65500 36040 65506
rect 36116 65500 36156 65506
rect 36226 65500 36292 65506
rect 36336 65500 36370 65506
rect 35352 65462 35558 65488
rect 35660 65462 35806 65488
rect 35878 65462 35996 65488
rect 36052 65472 36074 65483
rect 36138 65477 36156 65500
rect 36254 65483 36292 65500
rect 35352 65460 35520 65462
rect 35352 65434 35530 65460
rect 35352 65382 35520 65434
rect 35550 65382 35552 65462
rect 35740 65460 35806 65462
rect 35688 65434 35806 65460
rect 35906 65434 35968 65460
rect 36006 65438 36074 65472
rect 36105 65472 36156 65477
rect 36162 65472 36184 65483
rect 36105 65466 36184 65472
rect 36215 65472 36248 65477
rect 36254 65472 36294 65483
rect 36215 65466 36294 65472
rect 36325 65472 36358 65477
rect 36325 65466 36404 65472
rect 36116 65438 36184 65466
rect 36226 65438 36294 65466
rect 36336 65464 36404 65466
rect 36604 65464 36670 65600
rect 36858 65464 36860 65506
rect 36934 65464 37102 65600
rect 36336 65462 36442 65464
rect 36504 65462 36670 65464
rect 36722 65462 36880 65464
rect 36336 65438 36404 65462
rect 35740 65382 35806 65434
rect 36006 65432 36040 65438
rect 36116 65435 36156 65438
rect 36116 65432 36162 65435
rect 36226 65432 36292 65438
rect 36336 65432 36370 65438
rect 36604 65436 36670 65462
rect 36858 65436 36860 65462
rect 36414 65434 36442 65436
rect 36504 65434 36670 65436
rect 36722 65434 36880 65436
rect 36138 65430 36162 65432
rect 36248 65430 36292 65432
rect 36358 65430 36373 65432
rect 36052 65426 36118 65430
rect 36138 65426 36373 65430
rect 35832 65394 35884 65424
rect 35942 65394 35994 65424
rect 36052 65420 36373 65426
rect 36052 65400 36118 65420
rect 36120 65400 36156 65420
rect 36052 65394 36104 65400
rect 36118 65394 36156 65400
rect 36162 65400 36248 65420
rect 36254 65400 36358 65420
rect 36416 65400 36468 65430
rect 36526 65400 36578 65430
rect 36162 65394 36214 65400
rect 36254 65394 36324 65400
rect 36120 65382 36156 65394
rect 36254 65388 36292 65394
rect 36196 65382 36198 65388
rect 35352 65364 35996 65382
rect 35352 65354 35520 65364
rect 35538 65354 35540 65358
rect 35550 65354 35552 65364
rect 35740 65360 35806 65364
rect 35648 65354 35650 65358
rect 35740 65356 35832 65360
rect 35740 65354 35806 65356
rect 35834 65354 35854 65364
rect 35862 65354 35868 65364
rect 36162 65362 36198 65382
rect 36254 65362 36290 65388
rect 36306 65382 36334 65388
rect 36604 65382 36670 65434
rect 36858 65382 36860 65434
rect 36930 65400 37102 65464
rect 36934 65382 37102 65400
rect 36414 65370 37102 65382
rect 35884 65356 35942 65360
rect 35946 65354 35964 65358
rect 35972 65354 35980 65358
rect 35994 65356 36028 65360
rect 36037 65358 36086 65362
rect 36037 65356 36090 65358
rect 35352 65340 36024 65354
rect 36037 65347 36052 65356
rect 36082 65352 36090 65356
rect 36138 65356 36196 65362
rect 36248 65356 36306 65362
rect 36082 65340 36088 65352
rect 36138 65347 36162 65356
rect 36248 65352 36292 65356
rect 36248 65347 36294 65352
rect 34292 65336 35140 65340
rect 34292 65310 34454 65336
rect 34470 65318 34476 65336
rect 28368 65038 28426 65049
rect 28096 65034 28148 65038
rect 28206 65034 28258 65038
rect 28316 65034 28478 65038
rect 28046 65030 28420 65034
rect 28096 65008 28148 65030
rect 28206 65008 28258 65030
rect 28316 65008 28368 65030
rect 27730 64932 27784 64996
rect 28382 64996 28420 65030
rect 28426 65008 28478 65034
rect 28536 65008 28588 65038
rect 27794 64960 27952 64980
rect 28014 64960 28170 64980
rect 28232 64960 28260 64980
rect 28382 64970 28410 64996
rect 28426 64970 28462 64996
rect 28368 64955 28426 64970
rect 27794 64932 27952 64952
rect 28014 64932 28170 64952
rect 28232 64932 28288 64952
rect 27690 64644 27694 64686
rect 27692 64640 27694 64644
rect 27700 64636 27716 64756
rect 27740 64728 27784 64932
rect 27728 64714 27784 64728
rect 27724 64678 27784 64714
rect 27726 64670 27784 64678
rect 27728 64664 27784 64670
rect 27740 64494 27784 64664
rect 28040 64506 28055 64521
rect 28382 64506 28420 64955
rect 34159 64928 34286 64955
rect 34292 64928 34332 65310
rect 34338 65250 34430 65310
rect 34436 65262 34442 65310
rect 34468 65284 34476 65318
rect 34470 65282 34476 65284
rect 34484 65282 34504 65336
rect 34506 65310 34564 65336
rect 34518 65250 34538 65310
rect 34518 65248 34536 65250
rect 34546 65248 34552 65310
rect 34580 65282 34586 65336
rect 34594 65316 34614 65336
rect 34616 65316 34672 65336
rect 34690 65318 34696 65336
rect 34896 65332 35140 65336
rect 34594 65310 34672 65316
rect 34594 65306 34624 65310
rect 34628 65306 34648 65310
rect 34656 65295 34672 65310
rect 34656 65262 34662 65295
rect 34688 65284 34696 65318
rect 34834 65306 34844 65316
rect 34908 65284 34910 65298
rect 34690 65282 34696 65284
rect 34722 65282 34724 65284
rect 34942 65282 34944 65284
rect 34159 64908 34332 64928
rect 34196 64887 34332 64908
rect 34161 64869 34332 64887
rect 34161 64854 34344 64869
rect 34196 64828 34218 64854
rect 34344 64828 34374 64854
rect 34968 64840 34982 64904
rect 34996 64812 35010 64932
rect 35096 64756 35140 65332
rect 35476 65336 36088 65340
rect 35438 64812 35452 64932
rect 35476 64904 35520 65336
rect 35550 65332 35718 65336
rect 35740 65332 35832 65336
rect 35752 65318 35758 65332
rect 35604 65306 35614 65316
rect 35538 65282 35540 65298
rect 35752 65282 35760 65318
rect 35776 65316 35832 65332
rect 35834 65316 35854 65336
rect 35776 65310 35854 65316
rect 35776 65295 35792 65310
rect 35800 65306 35820 65310
rect 35824 65306 35854 65310
rect 35786 65262 35792 65295
rect 35862 65282 35868 65336
rect 35884 65310 35942 65336
rect 35896 65248 35902 65310
rect 35910 65250 35930 65310
rect 35944 65284 35964 65336
rect 35946 65282 35964 65284
rect 35972 65318 35978 65336
rect 35972 65282 35980 65318
rect 35994 65310 36088 65336
rect 36116 65319 36122 65346
rect 36138 65319 36156 65347
rect 36254 65346 36294 65347
rect 36006 65282 36088 65310
rect 36105 65314 36156 65319
rect 36162 65314 36184 65325
rect 36105 65308 36184 65314
rect 36215 65314 36248 65319
rect 36254 65316 36306 65346
rect 36322 65319 36328 65364
rect 36336 65346 36356 65364
rect 36358 65362 36416 65366
rect 36432 65354 36438 65364
rect 36446 65354 36466 65364
rect 36468 65362 36526 65366
rect 36542 65354 36548 65370
rect 36556 65354 36576 65370
rect 36604 65366 36670 65370
rect 36578 65362 36670 65366
rect 36604 65354 36670 65362
rect 36684 65356 36686 65364
rect 36794 65356 36796 65364
rect 36858 65354 36860 65370
rect 36904 65360 36906 65364
rect 36934 65354 37102 65370
rect 36386 65352 37102 65354
rect 36370 65346 37102 65352
rect 37314 65382 37482 65600
rect 37512 65382 37514 65506
rect 37702 65382 37768 65600
rect 38080 65441 38118 65890
rect 38252 65849 38344 65906
rect 38251 65838 38344 65849
rect 38252 65781 38344 65838
rect 38251 65770 38344 65781
rect 38252 65713 38344 65770
rect 38251 65702 38344 65713
rect 38252 65645 38344 65702
rect 38251 65634 38344 65645
rect 38252 65577 38344 65634
rect 38251 65566 38344 65577
rect 38252 65504 38344 65566
rect 38380 65504 38448 65964
rect 38841 65890 38856 65905
rect 38690 65860 38748 65890
rect 38800 65860 38856 65890
rect 38841 65845 38856 65860
rect 38252 65500 38470 65504
rect 38298 65476 38380 65500
rect 38308 65474 38380 65476
rect 38418 65474 38470 65500
rect 38528 65474 38580 65504
rect 38638 65474 38690 65504
rect 38748 65474 38800 65504
rect 38329 65468 38380 65474
rect 38066 65430 38124 65441
rect 38298 65436 38380 65468
rect 38252 65430 38344 65436
rect 37794 65400 37846 65430
rect 37904 65400 37956 65430
rect 38014 65426 38176 65430
rect 38014 65400 38066 65426
rect 38080 65388 38118 65426
rect 38124 65400 38176 65426
rect 38234 65426 38344 65430
rect 38234 65400 38296 65426
rect 38298 65420 38330 65426
rect 37314 65370 37958 65382
rect 37314 65354 37482 65370
rect 37500 65360 37502 65364
rect 37512 65354 37514 65370
rect 37702 65366 37768 65370
rect 37610 65356 37612 65364
rect 37702 65362 37794 65366
rect 37702 65354 37768 65362
rect 37796 65354 37816 65370
rect 37824 65354 37830 65370
rect 38080 65366 38108 65388
rect 37846 65362 37904 65366
rect 37908 65356 37926 65364
rect 37906 65354 37926 65356
rect 37934 65356 37942 65364
rect 37956 65362 38014 65366
rect 38018 65358 38036 65364
rect 37934 65354 37940 65356
rect 37314 65352 37986 65354
rect 37314 65346 38002 65352
rect 36358 65342 37102 65346
rect 36358 65319 36416 65342
rect 36432 65324 36438 65342
rect 36322 65316 36416 65319
rect 36254 65314 36294 65316
rect 36215 65308 36294 65314
rect 36006 65280 36085 65282
rect 36116 65280 36184 65308
rect 36006 65274 36040 65280
rect 36116 65274 36156 65280
rect 36226 65274 36294 65308
rect 36322 65314 36358 65316
rect 36398 65314 36404 65316
rect 36322 65308 36404 65314
rect 36322 65288 36328 65308
rect 36336 65280 36404 65308
rect 36430 65290 36438 65324
rect 36432 65288 36438 65290
rect 36446 65288 36466 65342
rect 36468 65316 36526 65342
rect 36336 65274 36370 65280
rect 36006 65262 36012 65274
rect 35912 65248 35930 65250
rect 36052 65246 36074 65257
rect 36116 65251 36122 65274
rect 36138 65251 36156 65274
rect 36006 65212 36074 65246
rect 36105 65246 36156 65251
rect 36162 65246 36184 65257
rect 36105 65240 36184 65246
rect 36215 65246 36248 65251
rect 36254 65246 36294 65274
rect 36398 65268 36404 65280
rect 36480 65256 36500 65316
rect 36480 65254 36498 65256
rect 36508 65254 36514 65316
rect 36542 65288 36548 65342
rect 36556 65322 36576 65342
rect 36578 65322 36634 65342
rect 36652 65324 36658 65342
rect 36858 65338 37102 65342
rect 36556 65316 36634 65322
rect 36556 65312 36586 65316
rect 36590 65312 36610 65316
rect 36618 65301 36634 65316
rect 36618 65268 36624 65301
rect 36650 65290 36658 65324
rect 36796 65312 36806 65322
rect 36870 65290 36872 65304
rect 36652 65288 36658 65290
rect 36684 65288 36686 65290
rect 36904 65288 36906 65290
rect 36215 65240 36294 65246
rect 36325 65246 36358 65251
rect 36325 65240 36404 65246
rect 36116 65212 36184 65240
rect 36006 65206 36040 65212
rect 36116 65206 36156 65212
rect 36226 65206 36294 65240
rect 36336 65212 36404 65240
rect 36336 65206 36370 65212
rect 36052 65178 36074 65189
rect 36138 65183 36156 65206
rect 36006 65144 36074 65178
rect 36105 65178 36156 65183
rect 36162 65178 36184 65189
rect 36105 65172 36184 65178
rect 36215 65178 36248 65183
rect 36254 65178 36294 65206
rect 36215 65172 36294 65178
rect 36325 65178 36358 65183
rect 36325 65172 36404 65178
rect 36116 65144 36184 65172
rect 36006 65138 36040 65144
rect 36116 65138 36156 65144
rect 36226 65138 36294 65172
rect 36336 65144 36404 65172
rect 36336 65138 36370 65144
rect 36052 65110 36074 65121
rect 36138 65115 36156 65138
rect 36006 65076 36074 65110
rect 36105 65110 36156 65115
rect 36162 65110 36184 65121
rect 36105 65104 36184 65110
rect 36215 65110 36248 65115
rect 36254 65110 36294 65138
rect 36215 65104 36294 65110
rect 36325 65110 36358 65115
rect 36325 65104 36404 65110
rect 36116 65076 36184 65104
rect 36006 65070 36040 65076
rect 36116 65070 36156 65076
rect 36226 65070 36294 65104
rect 36336 65076 36404 65104
rect 36336 65070 36370 65076
rect 36008 65060 36106 65068
rect 36014 65054 36106 65060
rect 36052 65042 36074 65053
rect 36138 65047 36156 65070
rect 36006 65040 36074 65042
rect 36105 65042 36156 65047
rect 36162 65042 36184 65053
rect 36006 65032 36080 65040
rect 36105 65036 36184 65042
rect 36215 65042 36248 65047
rect 36254 65042 36294 65070
rect 36215 65036 36294 65042
rect 36325 65042 36358 65047
rect 36325 65036 36404 65042
rect 36006 65008 36085 65032
rect 36116 65008 36184 65036
rect 36006 65002 36040 65008
rect 36116 65002 36156 65008
rect 36226 65002 36294 65036
rect 36336 65008 36404 65036
rect 36336 65002 36370 65008
rect 36052 64974 36074 64985
rect 36138 64979 36156 65002
rect 36006 64940 36074 64974
rect 36105 64974 36156 64979
rect 36162 64974 36184 64985
rect 36105 64968 36184 64974
rect 36215 64974 36248 64979
rect 36254 64974 36294 65002
rect 36215 64968 36294 64974
rect 36325 64974 36358 64979
rect 36325 64968 36404 64974
rect 36116 64961 36184 64968
rect 36226 64961 36294 64968
rect 36116 64946 36294 64961
rect 36116 64944 36306 64946
rect 36006 64934 36040 64940
rect 36116 64934 36308 64944
rect 36336 64940 36404 64968
rect 36336 64934 36370 64940
rect 36052 64906 36074 64917
rect 36121 64914 36308 64934
rect 36138 64911 36308 64914
rect 35466 64840 35520 64904
rect 36006 64872 36074 64906
rect 36105 64900 36308 64911
rect 36325 64906 36358 64911
rect 36388 64906 36442 64910
rect 36325 64900 36442 64906
rect 36116 64876 36308 64900
rect 36336 64898 36442 64900
rect 36504 64898 36660 64910
rect 36722 64898 36880 64910
rect 36006 64866 36040 64872
rect 36116 64866 36294 64876
rect 36336 64872 36410 64898
rect 36336 64866 36370 64872
rect 36416 64870 36442 64882
rect 36504 64870 36660 64882
rect 36722 64870 36880 64882
rect 36123 64860 36294 64866
rect 36358 64860 36373 64866
rect 36104 64854 36287 64860
rect 36324 64854 36373 64860
rect 36188 64846 36194 64854
rect 36216 64852 36222 64854
rect 36266 64852 36280 64854
rect 36170 64844 36204 64846
rect 36416 64844 36438 64870
rect 36930 64846 36944 64910
rect 36172 64840 36204 64844
rect 35476 64756 35520 64840
rect 36116 64828 36146 64834
rect 36190 64778 36192 64816
rect 36206 64806 36238 64840
rect 36958 64818 36972 64938
rect 36172 64772 36204 64778
rect 36218 64772 36220 64806
rect 36190 64752 36192 64772
rect 36206 64744 36238 64772
rect 37058 64762 37102 65338
rect 37438 65342 38014 65346
rect 37400 64818 37414 64938
rect 37438 64910 37482 65342
rect 37512 65338 37680 65342
rect 37702 65338 37794 65342
rect 37714 65324 37720 65338
rect 37566 65312 37576 65322
rect 37500 65288 37502 65304
rect 37714 65288 37722 65324
rect 37738 65322 37794 65338
rect 37796 65322 37816 65342
rect 37738 65316 37816 65322
rect 37738 65301 37754 65316
rect 37762 65312 37782 65316
rect 37786 65312 37816 65316
rect 37748 65268 37754 65301
rect 37824 65288 37830 65342
rect 37846 65316 37904 65342
rect 37858 65254 37864 65316
rect 37872 65256 37892 65316
rect 37906 65290 37926 65342
rect 37908 65288 37926 65290
rect 37934 65324 37940 65342
rect 37934 65288 37942 65324
rect 37956 65322 38014 65342
rect 38016 65322 38036 65358
rect 37956 65316 38036 65322
rect 37968 65268 37974 65316
rect 37982 65312 38002 65316
rect 38006 65312 38036 65316
rect 38044 65358 38052 65364
rect 38066 65362 38116 65366
rect 38124 65362 38160 65388
rect 38252 65362 38296 65400
rect 38044 65288 38050 65358
rect 38066 65347 38124 65362
rect 38252 65361 38344 65362
rect 38251 65350 38344 65361
rect 38078 65346 38118 65347
rect 38066 65316 38118 65346
rect 37874 65254 37892 65256
rect 38078 64934 38118 65316
rect 38252 65293 38344 65350
rect 38251 65282 38344 65293
rect 38252 65225 38344 65282
rect 38251 65214 38344 65225
rect 38252 65157 38344 65214
rect 38251 65146 38344 65157
rect 38252 65089 38344 65146
rect 38251 65078 38344 65089
rect 38252 65021 38344 65078
rect 38251 65010 38344 65021
rect 38124 64934 38251 64961
rect 38252 64945 38344 65010
rect 38380 64945 38448 65436
rect 38586 65366 39106 65382
rect 38586 65338 39134 65354
rect 38841 65334 38856 65338
rect 38648 65284 38650 65316
rect 38690 65304 38748 65334
rect 38800 65304 38856 65334
rect 38682 65262 38684 65300
rect 38841 65289 38856 65304
rect 38868 65284 38870 65316
rect 38934 65308 38946 65318
rect 38902 65264 38904 65300
rect 39088 65284 39090 65334
rect 39154 65308 39166 65318
rect 39122 65264 39124 65300
rect 38252 64944 38448 64945
rect 38078 64920 38251 64934
rect 38298 64920 38344 64944
rect 38078 64914 38270 64920
rect 38308 64918 38344 64920
rect 37428 64846 37482 64910
rect 37492 64898 37650 64910
rect 37712 64898 37868 64910
rect 37930 64898 37984 64910
rect 38078 64893 38124 64914
rect 38156 64898 38270 64914
rect 38329 64906 38344 64918
rect 38332 64903 38344 64906
rect 38640 64898 38798 64906
rect 38860 64898 39016 64906
rect 39078 64898 39132 64906
rect 39304 64898 39418 64916
rect 38170 64893 38214 64898
rect 37492 64870 37650 64882
rect 37712 64870 37868 64882
rect 37930 64870 37956 64882
rect 38078 64875 38249 64893
rect 38066 64860 38249 64875
rect 38640 64870 38798 64878
rect 38860 64870 39016 64878
rect 39078 64870 39104 64878
rect 39304 64870 39390 64888
rect 37438 64762 37482 64846
rect 38078 64834 38108 64860
rect 38234 64834 38256 64860
rect 37942 64816 37956 64834
rect 38092 64822 38102 64824
rect 37970 64792 37984 64806
rect 38064 64804 38074 64806
rect 38062 64802 38074 64804
rect 38090 64802 38102 64822
rect 38516 64814 39104 64830
rect 38562 64812 39104 64814
rect 37970 64788 37978 64792
rect 38062 64730 38072 64802
rect 38090 64758 38100 64802
rect 38488 64786 39132 64802
rect 38534 64784 39132 64786
rect 44972 64774 45204 64844
rect 28604 64584 28634 64600
rect 28646 64584 28682 64610
rect 28040 64472 28096 64506
rect 28148 64472 28206 64506
rect 28258 64472 28316 64506
rect 28368 64472 28420 64506
rect 28582 64566 28646 64584
rect 28582 64516 28668 64566
rect 28582 64482 28646 64516
rect 28040 64468 28055 64472
rect 28584 64468 28646 64482
rect 28046 64456 28096 64468
rect 28148 64456 28206 64468
rect 28258 64456 28316 64468
rect 28368 64456 28418 64468
rect 28584 64442 28588 64468
rect 28584 64431 28595 64442
rect 28682 64432 28708 64584
rect 44780 64520 44950 64774
rect 44972 64522 45740 64774
rect 45744 64646 45750 64724
rect 45852 64646 45858 64724
rect 45936 64646 45942 64724
rect 44820 64324 44826 64402
rect 44904 64324 44910 64402
rect 44820 64002 44826 64080
rect 44904 64002 44910 64080
rect 44820 63680 44826 63758
rect 44904 63680 44910 63758
rect 44658 63416 44666 63512
rect 44686 63444 44694 63484
rect 44820 63358 44826 63436
rect 44904 63358 44910 63436
rect 44780 63256 44852 63268
rect 44742 63236 44764 63240
rect 44740 63206 44764 63236
rect 44770 63208 44792 63212
rect 44768 63206 44792 63208
rect 44780 63130 44950 63166
rect 44742 63098 44764 63130
rect 44770 63126 44950 63130
rect 44780 62924 44950 63126
rect 44972 63164 45204 64520
rect 45276 64342 45282 64398
rect 45254 64320 45282 64342
rect 45360 64320 45366 64398
rect 45468 64320 45474 64398
rect 45552 64320 45558 64398
rect 45660 64320 45666 64398
rect 45744 64320 45750 64398
rect 45852 64324 45858 64402
rect 45936 64324 45942 64402
rect 45254 64308 45276 64320
rect 45288 64274 45310 64308
rect 45480 64274 45546 64276
rect 45486 64240 45524 64242
rect 45450 64204 45480 64210
rect 45348 64088 45354 64112
rect 45276 63998 45282 64076
rect 45348 64054 45388 64078
rect 45360 63998 45366 64054
rect 45468 63998 45474 64076
rect 45552 63998 45558 64076
rect 45660 63998 45666 64076
rect 45744 63998 45750 64076
rect 45852 64002 45858 64080
rect 45936 64002 45942 64080
rect 45500 63808 45512 63818
rect 45528 63808 45540 63846
rect 45458 63774 45466 63796
rect 45474 63759 45481 63808
rect 45500 63796 45552 63808
rect 45500 63793 45584 63796
rect 45500 63788 45512 63793
rect 45518 63780 45584 63793
rect 45620 63780 45626 63824
rect 45537 63765 45552 63780
rect 45276 63676 45282 63754
rect 45360 63676 45366 63754
rect 45468 63676 45474 63754
rect 45552 63676 45558 63754
rect 45660 63676 45666 63754
rect 45744 63676 45750 63754
rect 45852 63680 45858 63758
rect 45936 63680 45942 63758
rect 45282 63622 45301 63630
rect 45268 63574 45270 63596
rect 45218 63542 45270 63574
rect 45302 63562 45304 63630
rect 45300 63354 45306 63432
rect 45384 63354 45390 63432
rect 45428 63354 45452 63474
rect 45458 63452 45468 63474
rect 45474 63437 45483 63486
rect 45503 63474 45552 63486
rect 45503 63471 45584 63474
rect 45518 63458 45584 63471
rect 45620 63458 45626 63502
rect 45537 63443 45552 63458
rect 45468 63354 45474 63432
rect 45552 63354 45558 63432
rect 45660 63354 45666 63432
rect 45744 63354 45750 63432
rect 45852 63358 45858 63436
rect 45936 63358 45942 63436
rect 45325 63326 45384 63335
rect 45322 63300 45384 63326
rect 45322 63216 45348 63300
rect 45356 63250 45382 63292
rect 45428 63284 45458 63346
rect 45428 63280 45464 63284
rect 45428 63278 45536 63280
rect 45406 63254 45422 63262
rect 45428 63254 45548 63278
rect 45620 63254 45692 63264
rect 45812 63256 45884 63268
rect 45402 63238 45422 63254
rect 45444 63236 45472 63238
rect 45474 63236 45502 63238
rect 45444 63232 45460 63236
rect 45474 63232 45528 63236
rect 45444 63208 45660 63232
rect 45456 63176 45660 63208
rect 45456 63166 45706 63176
rect 44972 62952 45334 63164
rect 45348 63090 45406 63164
rect 45456 63090 45982 63166
rect 45348 62952 45982 63090
rect 44972 62944 45982 62952
rect 44972 62922 45334 62944
rect 45348 62934 45982 62944
rect 44780 62910 44950 62912
rect 45348 62910 45502 62934
rect 45548 62924 45982 62934
rect 45548 62922 45790 62924
rect 44820 62714 44826 62792
rect 44904 62714 44910 62792
rect 44820 62392 44826 62470
rect 44904 62392 44910 62470
rect 44820 62070 44826 62148
rect 44904 62070 44910 62148
rect 44820 61748 44826 61826
rect 44904 61748 44910 61826
rect 44972 61624 45204 62910
rect 45458 62808 45466 62830
rect 45474 62793 45481 62842
rect 45503 62830 45552 62842
rect 45503 62827 45584 62830
rect 45518 62812 45584 62827
rect 45620 62812 45626 62858
rect 45537 62797 45552 62812
rect 45276 62710 45282 62788
rect 45360 62710 45366 62788
rect 45468 62710 45474 62788
rect 45552 62710 45558 62788
rect 45660 62710 45666 62788
rect 45744 62710 45750 62788
rect 45852 62714 45858 62792
rect 45936 62714 45942 62792
rect 45458 62486 45464 62508
rect 45474 62471 45479 62520
rect 45501 62508 45552 62520
rect 45501 62505 45582 62508
rect 45516 62490 45582 62505
rect 45620 62490 45624 62536
rect 45537 62475 45552 62490
rect 45276 62388 45282 62466
rect 45360 62388 45366 62466
rect 45468 62388 45474 62466
rect 45552 62388 45558 62466
rect 45660 62388 45666 62466
rect 45744 62388 45750 62466
rect 45852 62392 45858 62470
rect 45936 62392 45942 62470
rect 46526 62376 46528 62450
rect 45428 62288 45482 62294
rect 45390 62214 45407 62236
rect 45334 62210 45454 62214
rect 45352 62186 45354 62190
rect 45359 62186 45360 62198
rect 45374 62196 45438 62210
rect 45386 62186 45388 62196
rect 45334 62182 45426 62186
rect 45346 62168 45426 62182
rect 45352 62156 45354 62168
rect 45386 62166 45388 62168
rect 45276 62066 45282 62144
rect 45360 62066 45366 62144
rect 45468 62066 45474 62144
rect 45552 62066 45558 62144
rect 45660 62066 45666 62144
rect 45744 62066 45750 62144
rect 45852 62070 45858 62148
rect 45936 62070 45942 62148
rect 45236 61966 45308 61968
rect 45428 61966 45500 61968
rect 45620 61966 45692 61968
rect 45458 61842 45464 61868
rect 45474 61827 45479 61878
rect 45501 61868 45552 61878
rect 45501 61863 45582 61868
rect 45516 61850 45582 61863
rect 45620 61850 45624 61896
rect 45537 61835 45552 61850
rect 45276 61748 45282 61826
rect 45360 61748 45366 61826
rect 45468 61748 45474 61826
rect 45552 61748 45558 61826
rect 45660 61748 45666 61826
rect 45744 61748 45750 61826
rect 45852 61748 45858 61826
rect 45936 61748 45942 61826
<< metal1 >>
rect 4724 77582 5502 77816
rect 10442 77580 11220 77814
rect 16160 77580 16938 77814
rect 24540 77586 25318 77820
rect 32964 77582 33742 77816
rect 38682 77582 39460 77816
rect 44402 77582 45180 77816
rect 50120 77582 50898 77816
rect 55838 77582 56616 77816
rect 61556 77580 62334 77814
rect 67274 77580 68052 77814
rect 5828 73118 6474 75740
rect 11546 73800 12192 75740
rect 17264 74658 17910 75740
rect 19772 75298 19806 75322
rect 17178 74596 17944 74658
rect 17178 74146 17264 74596
rect 17910 74146 17944 74596
rect 17178 74110 17944 74146
rect 19702 73986 19806 75298
rect 19690 73964 19820 73986
rect 19690 73890 19702 73964
rect 19806 73890 19820 73964
rect 19690 73884 19820 73890
rect 11514 73698 12214 73800
rect 11514 73248 11546 73698
rect 12192 73248 12214 73698
rect 11514 73222 12214 73248
rect 5394 73040 6474 73118
rect 5394 72394 5462 73040
rect 5912 72394 6474 73040
rect 2906 72378 3584 72392
rect 2712 72360 3584 72378
rect 2066 71714 3156 72360
rect 3528 71714 3584 72360
rect 5394 72358 5982 72394
rect 19702 72348 19806 73884
rect 20382 73102 20464 75344
rect 25804 74944 26036 75326
rect 25804 74718 31276 74944
rect 25804 74678 31314 74718
rect 31010 74398 31276 74678
rect 34068 74496 34714 75742
rect 36396 75326 36518 75354
rect 36392 74934 36628 75326
rect 36232 74752 36628 74934
rect 36232 74716 36594 74752
rect 37280 74720 37424 75492
rect 36232 74578 36378 74716
rect 39786 74496 40432 75740
rect 45504 74496 46150 75740
rect 47290 75218 47328 75220
rect 48716 75218 48860 75492
rect 47290 75148 48860 75218
rect 47290 74722 47328 75148
rect 51222 75110 51868 75740
rect 51070 75054 51868 75110
rect 51066 75014 51868 75054
rect 51030 74820 51900 75014
rect 51030 74408 51222 74820
rect 51868 74408 51900 74820
rect 51030 74274 51900 74408
rect 56940 74178 57586 75740
rect 56880 74090 57590 74178
rect 56880 73430 56940 74090
rect 57352 73430 57590 74090
rect 56880 73368 57590 73430
rect 20358 73096 20464 73102
rect 20358 73014 20370 73096
rect 20452 73014 20464 73096
rect 62658 73052 63304 75740
rect 20358 73008 20464 73014
rect 19662 72330 19806 72348
rect 19662 72226 19674 72330
rect 19778 72226 19806 72330
rect 19662 72202 19806 72226
rect 2712 71578 3584 71714
rect 0 70610 250 71388
rect 4740 66642 5192 66650
rect 2066 65996 4766 66642
rect 5182 65996 5192 66642
rect 4740 65988 5192 65996
rect 2 64894 252 65672
rect 19702 65132 19806 72202
rect 20382 72158 20464 73008
rect 62618 72992 63336 73052
rect 62618 72580 62658 72992
rect 63304 72580 63336 72992
rect 62618 72546 63336 72580
rect 68376 72354 69022 75740
rect 20354 72138 20478 72158
rect 20354 72056 20380 72138
rect 20462 72056 20478 72138
rect 20354 72040 20478 72056
rect 68314 72108 69066 72354
rect 19686 65126 19812 65132
rect 19686 65022 19694 65126
rect 19798 65022 19812 65126
rect 19686 65012 19812 65022
rect 20382 64928 20464 72040
rect 68314 71698 68376 72108
rect 69022 71698 69066 72108
rect 68314 71630 69066 71698
rect 71184 72216 71866 72280
rect 71184 71570 71244 72216
rect 71642 71570 72512 72216
rect 52848 71438 53732 71560
rect 71184 71472 71866 71570
rect 52848 71374 52896 71438
rect 53340 71374 53732 71438
rect 52848 65538 53732 71374
rect 74320 70470 74570 71248
rect 69502 66498 69966 66514
rect 69502 65852 69534 66498
rect 69952 65852 72510 66498
rect 69502 65840 69966 65852
rect 52842 65514 53736 65538
rect 52842 65296 52864 65514
rect 53720 65296 53736 65514
rect 52842 65274 53736 65296
rect 20372 64922 20468 64928
rect 20372 64834 20380 64922
rect 20462 64834 20468 64922
rect 20372 64828 20468 64834
rect 5522 60924 5968 60940
rect 2068 60278 5546 60924
rect 5962 60278 5968 60924
rect 5522 60248 5968 60278
rect 0 59174 250 59952
rect 6424 55206 6906 55226
rect 2066 54560 6472 55206
rect 6888 54560 6906 55206
rect 6424 54540 6906 54560
rect 4 53456 254 54234
rect 7336 49488 7790 49502
rect 2068 48842 7354 49488
rect 7770 48842 7790 49488
rect 7336 48822 7790 48842
rect 2 47740 252 48518
rect 8208 43770 8658 43782
rect 2066 43124 8222 43770
rect 8638 43124 8658 43770
rect 8208 43108 8658 43124
rect 0 42020 250 42798
rect 9072 38052 9522 38074
rect 2066 37406 9552 38052
rect 9072 37384 9522 37406
rect 2 36304 252 37082
rect 52848 33014 53732 65274
rect 74318 64750 74568 65528
rect 68668 60780 69140 60806
rect 68668 60134 68684 60780
rect 69102 60134 72514 60780
rect 68668 60114 69140 60134
rect 74318 59030 74568 59808
rect 67866 55062 68322 55094
rect 67866 54416 67888 55062
rect 68306 54416 72510 55062
rect 67866 54394 68322 54416
rect 74320 53318 74570 54096
rect 67006 49344 67490 49368
rect 67006 48698 67038 49344
rect 67456 48698 72510 49344
rect 67006 48666 67490 48698
rect 74316 47596 74566 48374
rect 66228 43626 66682 43648
rect 66228 42980 66250 43626
rect 66668 42980 72512 43626
rect 66228 42954 66682 42980
rect 74320 41880 74570 42658
rect 65348 37908 65808 37924
rect 65348 37262 72512 37908
rect 65348 37242 65808 37262
rect 74320 36158 74570 36936
rect 52664 32992 53732 33014
rect 9884 32334 10366 32354
rect 2066 31688 9930 32334
rect 10346 31688 10366 32334
rect 52664 32108 52700 32992
rect 53584 32266 53732 32992
rect 53584 32108 53616 32266
rect 52664 32074 53616 32108
rect 9884 31652 10366 31688
rect 8 30588 258 31366
rect 10740 26616 11232 26630
rect 2066 25970 11232 26616
rect 10740 25960 11232 25970
rect 4 24866 254 25644
rect 11614 20898 12094 20926
rect 2064 20252 11654 20898
rect 12070 20252 12094 20898
rect 11614 20232 12094 20252
rect 2 19148 252 19926
rect 12402 15180 12900 15196
rect 2064 14534 12448 15180
rect 12864 14534 12900 15180
rect 12402 14496 12900 14534
rect 2 13430 252 14208
rect 13296 9462 13766 9482
rect 2068 8816 13336 9462
rect 13752 8816 13766 9462
rect 13296 8790 13766 8816
rect 4 7712 254 8490
rect 14096 3744 14638 3756
rect 2068 3098 14196 3744
rect 14612 3098 14638 3744
rect 14096 3074 14638 3098
rect 4 1996 254 2774
<< via1 >>
rect 17264 74146 17910 74596
rect 19702 73890 19806 73964
rect 11546 73248 12192 73698
rect 5462 72394 5912 73040
rect 3156 71714 3528 72360
rect 51222 74408 51868 74820
rect 56940 73430 57352 74090
rect 20370 73014 20452 73096
rect 19674 72226 19778 72330
rect 4766 65996 5182 66642
rect 62658 72580 63304 72992
rect 20380 72056 20462 72138
rect 19694 65022 19798 65126
rect 68376 71698 69022 72108
rect 71244 71570 71642 72216
rect 52896 71374 53340 71438
rect 69534 65852 69952 66498
rect 52864 65296 53720 65514
rect 20380 64834 20462 64922
rect 5546 60278 5962 60924
rect 6472 54560 6888 55206
rect 7354 48842 7770 49488
rect 8222 43124 8638 43770
rect 68684 60134 69102 60780
rect 67888 54416 68306 55062
rect 67038 48698 67456 49344
rect 66250 42980 66668 43626
rect 9930 31688 10346 32334
rect 52700 32108 53584 32992
rect 11654 20252 12070 20898
rect 12448 14534 12864 15180
rect 13336 8816 13752 9462
rect 14196 3098 14612 3744
<< metal2 >>
rect 73698 77004 73936 77006
rect 684 77002 3270 77004
rect 658 76724 3270 77002
rect 71338 76900 73936 77004
rect 71296 76748 73936 76900
rect 658 76420 1116 76724
rect 748 76412 1116 76420
rect 836 74708 1116 76412
rect 73504 76484 73936 76748
rect 2090 75450 3240 75730
rect 71168 75464 72502 75744
rect 2090 74506 2370 75450
rect 50992 74820 51952 74980
rect 17152 74648 17970 74698
rect 17152 74596 25546 74648
rect 17152 74146 17264 74596
rect 17910 74198 25546 74596
rect 50992 74562 51222 74820
rect 48652 74408 51222 74562
rect 51868 74562 51952 74820
rect 51868 74408 51962 74562
rect 17910 74146 17970 74198
rect 48652 74150 51962 74408
rect 72220 74362 72500 75464
rect 73504 74638 73760 76484
rect 73608 74490 73760 74638
rect 17152 74078 17970 74146
rect 56910 74090 57572 74148
rect 19692 73976 19816 73980
rect 19692 73964 25522 73976
rect 19692 73890 19702 73964
rect 19806 73902 25522 73964
rect 19806 73890 19816 73902
rect 19692 73888 19816 73890
rect 11528 73750 12204 73772
rect 11446 73698 25546 73750
rect 56910 73736 56940 74090
rect 11446 73300 11546 73698
rect 11528 73248 11546 73300
rect 12192 73300 25546 73698
rect 48652 73430 56940 73736
rect 57352 73736 57572 74090
rect 57352 73430 57636 73736
rect 48652 73324 57636 73430
rect 12192 73248 12204 73300
rect 11528 73236 12204 73248
rect 20362 73096 20458 73098
rect 5420 73040 5948 73088
rect 5420 72852 5462 73040
rect 5404 72402 5462 72852
rect 5420 72394 5462 72402
rect 5912 72852 5948 73040
rect 20362 73014 20370 73096
rect 20452 73092 20458 73096
rect 20452 73016 25520 73092
rect 20452 73014 20458 73016
rect 20362 73012 20458 73014
rect 62588 72992 63374 73010
rect 62588 72920 62658 72992
rect 5912 72402 25466 72852
rect 48652 72580 62658 72920
rect 63304 72580 63374 72992
rect 48652 72508 63374 72580
rect 62588 72506 63374 72508
rect 5912 72394 5948 72402
rect 2974 72360 3552 72376
rect 5420 72368 5948 72394
rect 2974 71984 3156 72360
rect 2968 71714 3156 71984
rect 3528 71984 3552 72360
rect 19668 72330 19792 72336
rect 19668 72226 19674 72330
rect 19778 72318 19792 72330
rect 19778 72236 25456 72318
rect 19778 72226 19792 72236
rect 19668 72218 19792 72226
rect 70688 72216 71830 72366
rect 20362 72138 20470 72144
rect 20362 72056 20380 72138
rect 20462 72056 25448 72138
rect 68348 72108 69048 72160
rect 20362 72048 20470 72056
rect 68348 72052 68376 72108
rect 3528 71714 25392 71984
rect 2968 71612 25392 71714
rect 48652 71698 68376 72052
rect 69022 72052 69048 72108
rect 69022 71698 69066 72052
rect 48652 71642 69066 71698
rect 70688 71570 71244 72216
rect 71642 71570 71830 72216
rect 48688 71438 53354 71448
rect 48688 71374 52896 71438
rect 53340 71374 53354 71438
rect 48688 71362 53354 71374
rect 70688 71238 71830 71570
rect 70600 71230 71830 71238
rect 48652 71138 71830 71230
rect 4746 70680 25450 71096
rect 48652 70758 71798 71138
rect 4746 66658 5162 70680
rect 69532 70282 69950 70318
rect 5578 69704 25546 70120
rect 48652 69864 69950 70282
rect 4732 66642 5200 66658
rect 4732 65996 4766 66642
rect 5182 65996 5200 66642
rect 4732 65984 5200 65996
rect 4746 65810 5162 65984
rect 5578 60938 5994 69704
rect 5534 60924 5994 60938
rect 5534 60278 5546 60924
rect 5962 60278 5994 60924
rect 5534 60256 5994 60278
rect 5578 60190 5994 60256
rect 6446 68740 25546 69156
rect 48652 68784 69122 69202
rect 6446 55242 6862 68740
rect 7354 67800 25546 68216
rect 48652 67808 68306 68226
rect 6404 55206 6918 55242
rect 6404 54560 6472 55206
rect 6888 54560 6918 55206
rect 6404 54522 6918 54560
rect 6446 54514 6862 54522
rect 7354 49518 7770 67800
rect 8224 66948 25546 67364
rect 7322 49488 7800 49518
rect 7322 48842 7354 49488
rect 7770 48842 7800 49488
rect 7322 48804 7800 48842
rect 7354 48698 7770 48804
rect 8224 43796 8640 66948
rect 48652 66768 67488 67186
rect 9092 66134 25546 66550
rect 8188 43770 8678 43796
rect 8188 43124 8222 43770
rect 8638 43124 8678 43770
rect 8188 43092 8678 43124
rect 8224 43068 8640 43092
rect 9092 38094 9508 66134
rect 48652 65760 66662 66178
rect 9924 65304 25546 65720
rect 52846 65516 53752 65532
rect 48708 65514 53766 65516
rect 9042 37348 9562 38094
rect 9092 37282 9508 37348
rect 9924 32368 10340 65304
rect 48708 65296 52864 65514
rect 53720 65296 53766 65514
rect 48708 65286 53766 65296
rect 52846 65282 53752 65286
rect 19688 65126 19808 65128
rect 19688 65022 19694 65126
rect 19798 65118 19808 65126
rect 19798 65030 25556 65118
rect 19798 65022 19808 65030
rect 19688 65016 19808 65022
rect 20374 64922 20466 64924
rect 20374 64834 20380 64922
rect 20462 64834 25548 64922
rect 20374 64830 20466 64834
rect 10774 64274 25546 64690
rect 48716 64658 65814 65076
rect 9840 32334 10382 32368
rect 9840 31688 9930 32334
rect 10346 31688 10382 32334
rect 9840 31634 10382 31688
rect 9924 31490 10340 31634
rect 10774 26644 11190 64274
rect 11626 63422 25546 63838
rect 10708 25948 11256 26644
rect 10774 25786 11190 25948
rect 11626 20986 12042 63422
rect 12456 62414 25546 62830
rect 11582 20898 12140 20986
rect 11582 20252 11654 20898
rect 12070 20252 12140 20898
rect 11582 20176 12140 20252
rect 11626 20120 12042 20176
rect 12456 15230 12872 62414
rect 13326 61292 25546 61708
rect 12358 15180 12924 15230
rect 12358 14534 12448 15180
rect 12864 14534 12924 15180
rect 12358 14474 12924 14534
rect 12456 14362 12872 14474
rect 13326 9514 13742 61292
rect 14158 60352 25546 60768
rect 13256 9462 13786 9514
rect 13256 8816 13336 9462
rect 13752 8816 13786 9462
rect 13256 8770 13786 8816
rect 13326 8768 13742 8770
rect 14158 3774 14574 60352
rect 14120 3744 14654 3774
rect 14120 3098 14196 3744
rect 14612 3098 14654 3744
rect 14120 3068 14654 3098
rect 26466 1902 27134 60380
rect 28398 1042 28802 60360
rect 29210 1356 29614 60360
rect 29210 1044 29616 1356
rect 30004 1354 30408 60360
rect 30804 1354 31208 60360
rect 29210 1042 29614 1044
rect 30002 1042 30408 1354
rect 30802 1042 31208 1354
rect 31614 1042 32018 60360
rect 32416 1356 32820 60360
rect 32414 1044 32820 1356
rect 32416 1042 32820 1044
rect 33216 1042 33620 60360
rect 34034 1042 34438 60360
rect 34860 1354 35264 60360
rect 35660 1354 36064 60360
rect 36452 1354 36856 60360
rect 34858 1042 35264 1354
rect 35658 1042 36064 1354
rect 36450 1042 36856 1354
rect 37262 1356 37666 60360
rect 37262 1044 37668 1356
rect 37262 1042 37666 1044
rect 38080 1042 38484 60360
rect 38882 1352 39286 60360
rect 39690 1354 40094 60360
rect 38882 1042 39288 1352
rect 39690 1042 40096 1354
rect 40508 1350 40912 60360
rect 40508 1042 40914 1350
rect 41318 1042 41722 60360
rect 42112 1042 42516 60360
rect 42936 1042 43340 60360
rect 38884 1040 39288 1042
rect 40510 1038 40914 1042
rect 43762 1040 44166 60360
rect 44564 1042 44968 60360
rect 45366 1378 45770 60360
rect 45366 1046 45774 1378
rect 46184 1374 46588 60360
rect 46184 1042 46590 1374
rect 47018 1042 47422 60360
rect 47818 1374 48222 60360
rect 48620 1374 49024 60360
rect 49412 1374 49816 60360
rect 47818 1042 48224 1374
rect 48614 1042 49024 1374
rect 49410 1042 49816 1374
rect 50222 1374 50626 60360
rect 51034 1374 51438 60360
rect 65396 38372 65814 64658
rect 66244 43666 66662 65760
rect 67070 49362 67488 66768
rect 67888 55116 68306 67808
rect 68704 60816 69122 68784
rect 69532 66528 69950 69864
rect 69492 66498 69978 66528
rect 69492 65852 69534 66498
rect 69952 65852 69978 66498
rect 69492 65820 69978 65852
rect 69532 65686 69950 65820
rect 68656 60780 69158 60816
rect 68656 60134 68684 60780
rect 69102 60134 69158 60780
rect 68656 60102 69158 60134
rect 67848 55062 68352 55116
rect 67848 54416 67888 55062
rect 68306 54416 68352 55062
rect 67848 54374 68352 54416
rect 67888 54368 68306 54374
rect 67016 49344 67488 49362
rect 67016 48698 67038 49344
rect 67456 48698 67488 49344
rect 67016 48678 67488 48698
rect 67070 48536 67488 48678
rect 66210 43626 66696 43666
rect 66210 42980 66250 43626
rect 66668 42980 66696 43626
rect 66210 42924 66696 42980
rect 65398 37992 65814 38372
rect 65398 37968 65816 37992
rect 65376 37956 65816 37968
rect 65324 37220 65830 37956
rect 65376 37216 65794 37220
rect 73612 34678 73760 34746
rect 72216 34472 72496 34628
rect 73480 34598 73762 34678
rect 72214 34448 72496 34472
rect 73484 34460 73760 34598
rect 72212 34418 72496 34448
rect 72212 34238 72494 34418
rect 73482 34226 73762 34460
rect 52678 32992 53598 33002
rect 52678 32108 52700 32992
rect 53584 32846 53598 32992
rect 53584 32510 72508 32846
rect 53584 32252 72534 32510
rect 53584 32108 53598 32252
rect 52678 32088 53598 32108
rect 50222 1042 50630 1374
rect 51034 1042 51442 1374
rect 830 66 1110 460
rect 2090 0 2370 732
use sky130_hilas_TopProtection  sky130_hilas_TopProtection_0
timestamp 1632255311
transform 1 0 3186 0 1 75246
box 1490 0 69756 2786
use sky130_hilas_LeftProtection  sky130_hilas_LeftProtection_0
timestamp 1632255311
transform 1 0 4380 0 1 17330
box -296 1490 2464 75824
use sky130_hilas_TopLevelTextStructure  sky130_hilas_TopLevelTextStructure_0
timestamp 1632255311
transform 1 0 24956 0 1 61922
box -1152 -476 26050 15156
use sky130_hilas_RightProtection  sky130_hilas_RightProtection_0
timestamp 1632255311
transform 1 0 75972 0 1 17186
box 0 1490 2772 41516
<< labels >>
rlabel metal1 74320 36158 74570 36936 0 IO07
port 1 nsew
rlabel metal1 74320 41880 74570 42658 0 IO08
port 2 nsew
rlabel metal1 74316 47596 74566 48374 0 IO09
port 3 nsew
rlabel metal1 74320 53318 74570 54096 0 IO10
port 4 nsew
rlabel metal1 74318 59030 74568 59808 0 IO11
port 5 nsew
rlabel metal1 74318 64750 74568 65528 0 IO12
port 6 nsew
rlabel metal1 74320 70470 74570 71248 0 IO13
port 7 nsew
rlabel metal1 0 70610 250 71388 0 IO25
port 8 nsew
rlabel metal1 2 64894 252 65672 0 IO26
port 9 nsew
rlabel metal1 0 59174 250 59952 0 IO27
port 10 nsew
rlabel metal1 4 53456 254 54234 0 IO28
port 11 nsew
rlabel metal1 2 47740 252 48518 0 IO29
port 12 nsew
rlabel metal1 0 42020 250 42798 0 IO30
port 13 nsew
rlabel metal1 2 36304 252 37082 0 IO31
port 14 nsew
rlabel metal1 8 30588 258 31366 0 IO32
port 15 nsew
rlabel metal1 4 24866 254 25644 0 IO33
port 16 nsew
rlabel metal1 2 19148 252 19926 0 IO34
port 17 nsew
rlabel metal1 2 13430 252 14208 0 IO35
port 18 nsew
rlabel metal1 4 7712 254 8490 0 IO36
port 19 nsew
rlabel metal1 4 1996 254 2774 0 IO37
port 20 nsew
rlabel metal2 658 76420 994 77002 0 VSSA1
port 21 nsew
rlabel metal1 4724 77582 5502 77816 0 ANALOG10
port 22 nsew
rlabel metal1 10442 77580 11220 77814 0 ANALOG09
port 23 nsew
rlabel metal1 16160 77580 16938 77814 0 ANALOG08
port 24 nsew
rlabel metal1 24540 77586 25318 77820 0 ANALOG07
port 25 nsew
rlabel metal1 32964 77582 33742 77816 0 ANALOG06
port 26 nsew
rlabel metal1 38682 77582 39460 77816 0 ANALOG05
port 27 nsew
rlabel metal1 44402 77582 45180 77816 0 ANALOG04
port 28 nsew
rlabel metal1 50120 77582 50898 77816 0 ANALOG03
port 29 nsew
rlabel metal1 55838 77582 56616 77816 0 ANALOG02
port 30 nsew
rlabel metal1 61556 77580 62334 77814 0 ANALOG01
port 31 nsew
rlabel metal1 67274 77580 68052 77814 0 ANALOG00
port 32 nsew
rlabel metal2 73698 76490 73936 77006 0 VSSA1
port 33 nsew
rlabel metal2 2090 0 2370 280 0 VDDA1
port 34 nsew
rlabel metal2 830 66 1110 346 0 VSSA1
port 33 nsew
rlabel metal2 72214 34238 72494 34472 0 VDDA1
port 34 nsew
rlabel metal2 73482 34226 73762 34460 0 VSSA1
port 33 nsew
rlabel metal2 28398 1042 28802 1354 0 LADATAOUT00
port 36 nsew
rlabel metal2 29212 1044 29616 1356 0 LADATAOUT01
port 35 nsew
rlabel metal2 30002 1042 30406 1354 0 LADATAOUT02
port 37 nsew
rlabel metal2 30802 1042 31206 1354 0 LADATAOUT03
port 38 nsew
rlabel metal2 31614 1042 32018 1354 0 LADATAOUT04
port 39 nsew
rlabel metal2 32414 1044 32818 1356 0 LADATAOUT05
port 40 nsew
rlabel metal2 33216 1042 33620 1354 0 LADATAOUT06
port 41 nsew
rlabel metal2 34034 1042 34438 1354 0 LADATAOUT07
port 42 nsew
rlabel metal2 34858 1042 35262 1354 0 LADATAOUT08
port 43 nsew
rlabel metal2 35658 1042 36062 1354 0 LADATAOUT09
port 44 nsew
rlabel metal2 36450 1042 36854 1354 0 LADATAOUT10
port 45 nsew
rlabel metal2 37264 1044 37668 1356 0 LADATAOUT11
port 46 nsew
rlabel metal2 38080 1042 38484 1354 0 LADATAOUT12
port 47 nsew
rlabel metal2 38884 1040 39288 1352 0 LADATAOUT13
port 48 nsew
rlabel metal2 39692 1042 40096 1354 0 LADATAOUT14
port 49 nsew
rlabel metal2 40510 1038 40914 1350 0 LADATAOUT15
port 50 nsew
rlabel metal2 41318 1042 41722 1354 0 LADATA16
port 51 nsew
rlabel metal2 42112 1042 42516 1354 0 LADATAOUT17
port 52 nsew
rlabel metal2 42936 1044 43340 1356 0 LADATAOUT18
port 53 nsew
rlabel metal2 43762 1040 44166 1352 0 LADATAOUT19
port 54 nsew
rlabel metal2 44564 1042 44968 1354 0 LADATAOUT20
port 55 nsew
rlabel metal2 45366 1046 45774 1378 0 LADATAOUT21
port 56 nsew
rlabel metal2 46184 1042 46590 1374 0 LADATAOUT22
port 57 nsew
rlabel metal2 47014 1042 47420 1374 0 LADATAOUT23
port 58 nsew
rlabel metal2 47818 1042 48224 1374 0 LADATAOUT24
port 59 nsew
rlabel metal2 48614 1042 49020 1374 0 LADATAIN00
port 60 nsew
rlabel metal2 49410 1042 49816 1374 0 LADATAIN01
port 61 nsew
rlabel metal2 50224 1042 50630 1374 0 LADATAIN02
port 62 nsew
rlabel metal2 51036 1042 51442 1374 0 LADATAIN03
port 63 nsew
rlabel metal2 72302 32252 72534 32504 0 VCCA
port 64 nsew
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
