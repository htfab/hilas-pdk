magic
tech sky130A
timestamp 1627061235
<< error_s >>
rect 681 365 683 366
<< nwell >>
rect 237 496 1380 503
<< locali >>
rect 398 503 415 504
rect 1295 503 1316 581
rect 1362 503 1379 571
rect 237 480 1380 503
rect 237 124 254 480
rect 303 1 320 447
rect 398 124 415 480
rect 466 1 483 443
rect 557 124 574 480
rect 626 1 643 451
rect 719 124 736 480
rect 788 1 805 446
rect 881 126 898 480
rect 948 1 965 451
rect 1041 127 1058 480
rect 1110 1 1127 451
rect 1202 126 1219 480
rect 1270 1 1287 449
rect 1363 123 1380 480
rect 1431 1 1448 467
<< metal1 >>
rect 674 356 1019 373
rect 829 103 847 257
rect 999 172 1019 356
rect 304 1 1658 24
<< metal2 >>
rect 0 578 705 597
rect 0 576 15 578
rect 0 496 206 502
rect 348 496 370 542
rect 840 497 865 573
rect 840 496 868 497
rect 0 481 868 496
rect 26 457 46 481
rect 190 466 868 481
rect 1011 309 1031 565
rect 0 288 1031 309
rect 1171 211 1186 585
rect 1271 569 1387 597
rect 1346 568 1387 569
rect 0 191 1187 211
rect 0 190 14 191
rect 0 79 854 99
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_8
timestamp 1607270276
transform 1 0 202 0 1 566
box -9 -26 24 29
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_9
timestamp 1607270276
transform 1 0 43 0 1 565
box -9 -26 24 29
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_10
timestamp 1607270276
transform 1 0 29 0 1 434
box -9 -26 24 29
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_11
timestamp 1607270276
transform 1 0 35 0 1 339
box -9 -26 24 29
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_12
timestamp 1607270276
transform 1 0 35 0 1 245
box -9 -26 24 29
use sky130_hilas_DAC6TransistorStack01a  sky130_hilas_DAC6TransistorStack01a_0
timestamp 1607478455
transform 1 0 9 0 1 177
box 28 -174 200 391
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1607179295
transform 1 0 311 0 1 8
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_6
timestamp 1607179295
transform 1 0 473 0 1 8
box -10 -8 13 21
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_6
timestamp 1607270276
transform 1 0 522 0 1 565
box -9 -26 24 29
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_7
timestamp 1607270276
transform 0 1 357 -1 0 549
box -9 -26 24 29
use sky130_hilas_DAC6TransistorStack01  sky130_hilas_DAC6TransistorStack01_0
array 0 2 161 0 0 566
timestamp 1607480432
transform 1 0 170 0 1 177
box 28 -174 200 391
use sky130_hilas_li2m1  sky130_hilas_li2m1_7
timestamp 1607179295
transform 1 0 633 0 1 8
box -10 -8 13 21
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_5
timestamp 1607270276
transform 1 0 683 0 1 565
box -9 -26 24 29
use sky130_hilas_DAC6TransistorStack01b  sky130_hilas_DAC6TransistorStack01b_0
timestamp 1607480432
transform 1 0 653 0 1 177
box 15 -174 200 391
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1607949437
transform 1 0 835 0 1 83
box -9 -10 23 22
use sky130_hilas_li2m1  sky130_hilas_li2m1_5
timestamp 1607179295
transform 1 0 955 0 1 8
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1607179295
transform 1 0 795 0 1 8
box -10 -8 13 21
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_4
timestamp 1607270276
transform 1 0 845 0 1 565
box -9 -26 24 29
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_3
timestamp 1607270276
transform 1 0 1006 0 1 566
box -9 -26 24 29
use sky130_hilas_DAC6TransistorStack01c  sky130_hilas_DAC6TransistorStack01c_0
timestamp 1607478930
transform 1 0 814 0 1 177
box 28 -174 215 391
use sky130_hilas_DAC6TransistorStack01  sky130_hilas_DAC6TransistorStack01_2
array 0 2 161 0 0 566
timestamp 1607480432
transform 1 0 975 0 1 177
box 28 -174 200 391
use sky130_hilas_DAC6TransistorStack01a  sky130_hilas_DAC6TransistorStack01a_1
timestamp 1607478455
transform 1 0 1458 0 1 177
box 28 -174 200 391
use sky130_hilas_li2m1  sky130_hilas_li2m1_2
timestamp 1607179295
transform 1 0 1117 0 1 8
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_4
timestamp 1607179295
transform 1 0 1438 0 1 8
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_3
timestamp 1607179295
transform 1 0 1277 0 1 8
box -10 -8 13 21
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1607089160
transform 1 0 1364 0 1 566
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1607089160
transform 1 0 1297 0 1 566
box -14 -15 20 18
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_2
timestamp 1607270276
transform 1 0 1167 0 1 566
box -9 -26 24 29
<< labels >>
rlabel metal2 1 576 11 597 0 A4
port 5 nsew analog default
rlabel metal2 0 481 10 502 0 A3
port 4 nsew analog default
rlabel metal2 1 288 11 309 0 A2
port 3 nsew analog default
rlabel metal2 1 190 11 211 0 A1
port 2 nsew analog default
rlabel metal2 0 79 8 99 0 A0
port 1 nsew analog default
rlabel metal2 1271 583 1346 597 0 VPWR
port 6 nsew analog default
rlabel metal1 1646 1 1658 24 0 OUT
port 7 nsew analog default
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
