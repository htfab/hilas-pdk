magic
tech sky130A
timestamp 1627742263
<< error_s >>
rect -18 20 21 23
rect -18 -22 21 -19
<< nwell >>
rect -121 -55 82 44
<< pmos >>
rect -18 -19 21 20
<< pdiff >>
rect -46 9 -18 20
rect -46 -8 -41 9
rect -24 -8 -18 9
rect -46 -19 -18 -8
rect 21 9 48 20
rect 21 -8 27 9
rect 44 -8 48 9
rect 21 -19 48 -8
<< pdiffc >>
rect -41 -8 -24 9
rect 27 -8 44 9
<< poly >>
rect -18 20 21 33
rect -80 -27 -54 -19
rect -18 -27 21 -19
rect -80 -42 21 -27
<< locali >>
rect -55 9 -24 17
rect -55 -1 -41 9
rect -57 -3 -41 -1
rect -41 -16 -24 -8
rect 27 9 44 17
rect 27 -16 44 -8
<< metal2 >>
rect -121 -3 -84 16
rect -121 -45 -83 -26
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_0
timestamp 1627742263
transform 0 1 -87 -1 0 -28
box -9 -26 24 29
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1627742263
transform 1 0 57 0 1 -1
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1627742263
transform 1 0 -73 0 1 9
box -14 -15 20 18
<< end >>
