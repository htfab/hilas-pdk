magic
tech sky130A
timestamp 1631574905
<< nwell >>
rect 310 -168 555 1
rect 310 -169 421 -168
<< nmos >>
rect 334 -548 539 -528
<< pmos >>
rect 336 -102 537 -82
<< ndiff >>
rect 334 -505 539 -501
rect 334 -522 350 -505
rect 524 -522 539 -505
rect 334 -528 539 -522
rect 334 -554 539 -548
rect 334 -571 350 -554
rect 524 -571 539 -554
rect 334 -580 539 -571
<< pdiff >>
rect 336 -58 537 -47
rect 336 -75 348 -58
rect 525 -75 537 -58
rect 336 -82 537 -75
rect 336 -108 537 -102
rect 336 -125 348 -108
rect 525 -125 537 -108
rect 336 -130 537 -125
<< ndiffc >>
rect 350 -522 524 -505
rect 350 -571 524 -554
<< pdiffc >>
rect 348 -75 525 -58
rect 348 -125 525 -108
<< psubdiff >>
rect 334 -591 539 -580
rect 334 -593 388 -591
rect 405 -593 425 -591
rect 442 -593 460 -591
rect 477 -593 496 -591
rect 513 -593 539 -591
rect 334 -610 349 -593
rect 525 -610 539 -593
rect 334 -616 539 -610
<< nsubdiff >>
rect 336 -24 537 -17
rect 336 -41 348 -24
rect 525 -41 537 -24
rect 336 -47 537 -41
<< psubdiffcont >>
rect 388 -593 405 -591
rect 425 -593 442 -591
rect 460 -593 477 -591
rect 496 -593 513 -591
rect 349 -610 525 -593
<< nsubdiffcont >>
rect 348 -41 525 -24
<< poly >>
rect 322 -102 336 -82
rect 537 -102 566 -82
rect 551 -147 566 -102
rect 322 -155 566 -147
rect 322 -172 349 -155
rect 522 -172 566 -155
rect 322 -177 566 -172
rect 321 -465 562 -460
rect 321 -482 351 -465
rect 525 -482 562 -465
rect 321 -489 562 -482
rect 547 -528 562 -489
rect 321 -548 334 -528
rect 539 -548 562 -528
<< polycont >>
rect 349 -172 522 -155
rect 351 -482 525 -465
<< locali >>
rect 340 -24 537 -22
rect 340 -41 348 -24
rect 525 -41 537 -24
rect 340 -42 364 -41
rect 381 -42 429 -41
rect 446 -42 494 -41
rect 511 -42 537 -41
rect 340 -58 537 -42
rect 340 -75 348 -58
rect 525 -75 537 -58
rect 340 -78 396 -75
rect 413 -78 463 -75
rect 480 -78 537 -75
rect 340 -80 537 -78
rect 491 -108 535 -105
rect 340 -125 348 -108
rect 525 -125 535 -108
rect 491 -126 505 -125
rect 522 -126 535 -125
rect 491 -129 535 -126
rect 341 -155 381 -152
rect 341 -172 349 -155
rect 522 -172 530 -155
rect 341 -175 381 -172
rect 343 -482 351 -465
rect 525 -482 534 -465
rect 494 -484 534 -482
rect 342 -505 389 -502
rect 342 -522 350 -505
rect 524 -522 532 -505
rect 342 -523 353 -522
rect 370 -523 389 -522
rect 342 -525 389 -523
rect 341 -554 532 -552
rect 341 -571 350 -554
rect 524 -571 532 -554
rect 341 -572 371 -571
rect 388 -572 407 -571
rect 424 -572 443 -571
rect 460 -572 479 -571
rect 496 -572 532 -571
rect 341 -591 532 -572
rect 341 -593 352 -591
rect 369 -593 388 -591
rect 341 -610 349 -593
rect 405 -593 425 -591
rect 442 -593 460 -591
rect 477 -593 496 -591
rect 513 -593 532 -591
rect 525 -610 533 -593
rect 341 -613 525 -610
<< viali >>
rect 364 -41 381 -25
rect 429 -41 446 -25
rect 494 -41 511 -25
rect 364 -42 381 -41
rect 429 -42 446 -41
rect 494 -42 511 -41
rect 396 -75 413 -61
rect 463 -75 480 -61
rect 396 -78 413 -75
rect 463 -78 480 -75
rect 505 -125 522 -109
rect 505 -126 522 -125
rect 354 -172 371 -155
rect 505 -482 522 -465
rect 353 -522 370 -505
rect 353 -523 370 -522
rect 371 -571 388 -555
rect 407 -571 424 -555
rect 443 -571 460 -555
rect 479 -571 496 -555
rect 371 -572 388 -571
rect 407 -572 424 -571
rect 443 -572 460 -571
rect 479 -572 496 -571
rect 352 -593 369 -591
rect 352 -608 369 -593
rect 388 -608 405 -591
rect 460 -608 477 -591
rect 496 -608 513 -591
<< metal1 >>
rect 357 11 518 13
rect 357 -15 361 11
rect 387 -15 425 11
rect 451 -15 489 11
rect 515 -15 518 11
rect 357 -25 518 -15
rect 357 -42 364 -25
rect 381 -42 429 -25
rect 446 -42 494 -25
rect 511 -42 518 -25
rect 357 -45 518 -42
rect 360 -46 518 -45
rect 360 -61 534 -46
rect 360 -78 396 -61
rect 413 -78 463 -61
rect 480 -78 534 -61
rect 360 -81 534 -78
rect 494 -109 534 -81
rect 494 -126 505 -109
rect 522 -126 534 -109
rect 344 -155 384 -151
rect 344 -172 354 -155
rect 371 -172 384 -155
rect 344 -505 384 -172
rect 494 -465 534 -126
rect 494 -482 505 -465
rect 522 -482 534 -465
rect 494 -485 534 -482
rect 344 -523 353 -505
rect 370 -523 384 -505
rect 344 -552 384 -523
rect 344 -554 519 -552
rect 347 -555 519 -554
rect 347 -572 371 -555
rect 388 -572 407 -555
rect 424 -572 443 -555
rect 460 -572 479 -555
rect 496 -572 519 -555
rect 347 -586 519 -572
rect 346 -591 519 -586
rect 346 -593 352 -591
rect 334 -608 352 -593
rect 369 -599 388 -591
rect 405 -599 460 -591
rect 477 -599 496 -591
rect 405 -608 415 -599
rect 334 -610 363 -608
rect 346 -625 363 -610
rect 389 -625 415 -608
rect 441 -608 460 -599
rect 493 -608 496 -599
rect 513 -608 519 -591
rect 441 -625 467 -608
rect 493 -625 519 -608
rect 346 -629 519 -625
<< via1 >>
rect 361 -15 387 11
rect 425 -15 451 11
rect 489 -15 515 11
rect 363 -608 369 -599
rect 369 -608 388 -599
rect 388 -608 389 -599
rect 363 -625 389 -608
rect 415 -625 441 -599
rect 467 -608 477 -599
rect 477 -608 493 -599
rect 467 -625 493 -608
<< metal2 >>
rect 246 11 619 17
rect 246 -15 361 11
rect 387 -15 425 11
rect 451 -15 489 11
rect 515 -15 619 11
rect 246 -21 619 -15
rect 246 -75 619 -49
rect 246 -139 619 -113
rect 246 -199 619 -173
rect 246 -253 619 -227
rect 246 -307 619 -281
rect 246 -359 619 -333
rect 246 -411 619 -385
rect 246 -463 619 -437
rect 246 -515 619 -489
rect 246 -567 619 -541
rect 246 -599 619 -593
rect 246 -625 363 -599
rect 389 -625 415 -599
rect 441 -625 467 -599
rect 493 -625 619 -599
rect 246 -633 619 -625
<< labels >>
rlabel metal2 608 -21 619 17 0 VPWR
port 1 nsew
rlabel metal2 246 -21 256 17 0 VPWR
port 1 nsew
rlabel metal2 608 -633 619 -593 0 VGND
port 2 nsew
rlabel metal2 246 -633 257 -593 0 VGND
port 2 nsew
<< end >>
