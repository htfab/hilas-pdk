magic
tech sky130A
timestamp 1627737364
<< error_s >>
rect -147 86 -97 97
rect 173 86 223 97
rect -97 80 -67 86
rect 145 80 173 86
rect 223 80 251 86
rect -72 61 -67 80
rect -210 56 -193 58
rect -48 55 -43 61
rect -147 44 -97 55
rect -48 48 -43 49
rect -48 44 -31 48
rect 173 44 223 55
rect -210 37 -193 39
rect -147 25 -97 35
rect -7 24 43 35
rect 173 24 223 35
rect -210 22 -193 24
rect -210 3 -193 5
rect -147 -17 -97 -7
rect -7 -18 43 -7
rect 173 -18 223 -7
<< nwell >>
rect -232 -40 110 119
<< mvnmos >>
rect 173 55 223 86
rect 173 -7 223 24
<< mvpmos >>
rect -147 55 -97 86
rect -147 -7 -97 25
rect -7 -7 43 24
<< mvndiff >>
rect 145 79 173 86
rect 145 62 150 79
rect 167 62 173 79
rect 145 55 173 62
rect 223 79 251 86
rect 223 62 229 79
rect 246 62 251 79
rect 223 55 251 62
rect 145 17 173 24
rect 145 0 150 17
rect 167 0 173 17
rect 145 -7 173 0
rect 223 17 251 24
rect 223 0 229 17
rect 246 0 251 17
rect 223 -7 251 0
<< mvpdiff >>
rect -177 78 -147 86
rect -177 61 -170 78
rect -153 61 -147 78
rect -177 55 -147 61
rect -97 79 -67 86
rect -97 62 -91 79
rect -74 62 -67 79
rect -97 55 -67 62
rect -177 18 -147 25
rect -177 1 -170 18
rect -153 1 -147 18
rect -177 -7 -147 1
rect -97 17 -67 25
rect -97 0 -91 17
rect -73 0 -67 17
rect -97 -7 -67 0
rect -37 17 -7 24
rect -37 0 -30 17
rect -13 0 -7 17
rect -37 -7 -7 0
rect 43 17 73 24
rect 43 0 49 17
rect 66 0 73 17
rect 43 -7 73 0
<< mvndiffc >>
rect 150 62 167 79
rect 229 62 246 79
rect 150 0 167 17
rect 229 0 246 17
<< mvpdiffc >>
rect -170 61 -153 78
rect -91 62 -74 79
rect -170 1 -153 18
rect -91 0 -73 17
rect -30 0 -13 17
rect 49 0 66 17
<< psubdiff >>
rect 283 22 314 34
rect 283 5 287 22
rect 304 5 314 22
rect 283 -7 314 5
<< nsubdiff >>
rect -214 56 -189 86
rect -214 39 -210 56
rect -193 39 -189 56
rect -214 22 -189 39
rect -214 5 -210 22
rect -193 5 -189 22
rect -214 -7 -189 5
<< psubdiffcont >>
rect 287 5 304 22
<< nsubdiffcont >>
rect -210 39 -193 56
rect -210 5 -193 22
<< poly >>
rect -147 96 319 103
rect -147 88 294 96
rect -147 86 -97 88
rect 173 86 223 88
rect -58 61 43 67
rect -147 25 -97 55
rect -58 44 -48 61
rect -31 44 43 61
rect 283 79 294 88
rect 311 79 319 96
rect 283 74 319 79
rect -58 38 43 44
rect -7 24 43 38
rect 173 24 223 55
rect -147 -20 -97 -7
rect -7 -20 43 -7
rect 173 -20 223 -7
<< polycont >>
rect -48 44 -31 61
rect 294 79 311 96
<< locali >>
rect 294 96 311 104
rect -170 78 -153 86
rect -100 62 -91 79
rect -74 62 150 79
rect 167 62 175 79
rect 221 62 229 79
rect 246 62 258 79
rect 294 69 311 79
rect -170 50 -153 61
rect -56 61 -23 62
rect -56 44 -48 61
rect -31 44 -23 61
rect 294 52 300 69
rect 294 48 311 52
rect -170 18 -153 33
rect 287 22 304 30
rect -170 -7 -153 1
rect -100 0 -91 17
rect -73 1 -72 17
rect 199 17 223 21
rect -55 1 -30 17
rect -73 0 -30 1
rect -13 0 -4 17
rect 41 0 49 17
rect 66 0 128 17
rect 145 0 150 17
rect 167 0 175 17
rect 199 0 203 17
rect 220 0 229 17
rect 246 0 256 17
rect 199 -3 223 0
<< viali >>
rect -210 56 -193 73
rect -210 22 -193 39
rect -210 -12 -193 5
rect -170 33 -153 50
rect 300 52 317 69
rect -72 1 -55 18
rect 128 0 145 17
rect 203 0 220 17
rect 287 -12 304 5
<< metal1 >>
rect -174 89 -149 119
rect -213 73 -149 89
rect -213 56 -210 73
rect -193 56 -149 73
rect -213 50 -149 56
rect -213 39 -170 50
rect -213 22 -210 39
rect -193 33 -170 39
rect -153 33 -149 50
rect -193 22 -149 33
rect -213 5 -149 22
rect -59 22 -25 25
rect -59 21 -54 22
rect -213 -12 -210 5
rect -193 -12 -149 5
rect -81 18 -54 21
rect -81 1 -72 18
rect -55 1 -54 18
rect -81 -2 -54 1
rect -59 -4 -54 -2
rect -28 17 -25 22
rect 125 17 148 119
rect 260 31 279 119
rect 293 74 325 75
rect 293 48 296 74
rect 322 48 325 74
rect 293 47 325 48
rect -28 0 -13 17
rect 125 0 128 17
rect 145 0 148 17
rect -28 -4 -25 0
rect -59 -7 -25 -4
rect -213 -18 -149 -12
rect -174 -40 -149 -18
rect 125 -40 148 0
rect 184 22 221 23
rect 184 -4 187 22
rect 213 17 226 22
rect 220 0 226 17
rect 213 -4 226 0
rect 260 5 307 31
rect 184 -6 221 -4
rect 260 -12 287 5
rect 304 -12 307 5
rect 260 -18 307 -12
rect 260 -40 279 -18
<< via1 >>
rect -54 -4 -28 22
rect 296 69 322 74
rect 296 52 300 69
rect 300 52 317 69
rect 317 52 322 69
rect 296 48 322 52
rect 187 17 213 22
rect 187 0 203 17
rect 203 0 213 17
rect 187 -4 213 0
<< metal2 >>
rect 292 74 326 76
rect 292 48 296 74
rect 322 69 326 74
rect 322 48 336 69
rect 292 46 336 48
rect 184 22 216 25
rect -57 -4 -54 22
rect -28 17 -25 22
rect 184 17 187 22
rect -28 -2 187 17
rect -28 -4 -25 -2
rect 184 -4 187 -2
rect 213 -4 216 22
rect 184 -7 216 -4
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1627737364
transform 1 0 266 0 1 65
box -10 -8 13 21
<< end >>
