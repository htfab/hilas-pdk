VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_ptransistorpair
  CLASS BLOCK ;
  FOREIGN sky130_hilas_ptransistorpair ;
  ORIGIN -1.330 4.400 ;
  SIZE 1.870 BY 6.050 ;
  OBS
      LAYER nwell ;
        RECT 1.330 -1.400 3.190 -1.330 ;
        RECT 2.670 -1.690 3.120 -1.460 ;
      LAYER li1 ;
        RECT 2.790 -0.700 3.010 -0.610 ;
        RECT 2.790 -0.780 2.870 -0.700 ;
        RECT 1.740 -1.920 1.920 -0.860 ;
        RECT 2.470 -1.330 2.520 -1.200 ;
        RECT 2.350 -1.460 2.520 -1.330 ;
        RECT 2.720 -3.520 2.790 -3.500 ;
        RECT 2.720 -3.660 2.800 -3.520 ;
        RECT 2.490 -4.350 2.560 -4.090 ;
      LAYER met1 ;
        RECT 2.830 -2.650 3.040 -0.880 ;
      LAYER met2 ;
        RECT 2.250 -1.690 3.120 -1.460 ;
        RECT 2.250 -1.700 2.680 -1.690 ;
        RECT 2.730 -2.490 3.200 -2.240 ;
        RECT 2.550 -3.520 3.100 -3.270 ;
        RECT 2.010 -4.380 2.890 -4.130 ;
  END
END sky130_hilas_ptransistorpair
END LIBRARY

