magic
tech sky130A
timestamp 1628707338
<< checkpaint >>
rect -42 1175 1502 1420
rect -485 952 1502 1175
rect -592 -383 1502 952
rect -485 -427 1502 -383
rect -485 -672 1059 -427
<< metal2 >>
rect 0 485 578 503
rect 0 442 578 460
rect 3 342 578 360
rect 3 299 578 317
rect 2 237 29 265
rect 542 241 579 269
rect 3 184 578 201
rect 3 142 578 159
rect 3 44 578 61
rect 3 0 578 17
<< metal3 >>
rect 145 290 172 291
rect 145 215 559 290
<< metal4 >>
rect 258 278 302 362
rect 116 277 217 278
rect 257 277 303 278
rect 45 227 303 277
rect 45 226 152 227
rect 257 161 303 227
rect 257 111 305 161
rect 302 81 305 111
use sky130_hilas_m22m4  sky130_hilas_m22m4_0
timestamp 1628707333
transform 1 0 38 0 1 247
box 0 0 79 75
use sky130_hilas_m22m4  sky130_hilas_m22m4_1
timestamp 1628707333
transform 1 0 523 0 1 251
box 0 0 79 75
use sky130_hilas_CapModule01  sky130_hilas_CapModule01_0
timestamp 1628705754
transform 1 0 588 0 1 203
box 0 0 284 286
use sky130_hilas_CapModule01  sky130_hilas_CapModule01_1
timestamp 1628705754
transform 1 0 588 0 1 504
box 0 0 284 286
<< labels >>
rlabel metal2 2 237 9 265 0 CAPTERM01
port 2 nsew analog default
rlabel metal2 571 241 579 269 0 CAPTERM02
port 1 nsew analog default
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
