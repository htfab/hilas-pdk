magic
tech sky130A
timestamp 1628704262
<< checkpaint >>
rect 2197 916 3624 1218
rect 2063 -75 3624 916
rect 2063 -373 3481 -75
rect 2069 -428 3481 -373
rect 2194 -463 3481 -428
<< error_s >>
rect 964 566 993 582
rect 1043 566 1072 582
rect 1122 566 1151 582
rect 1201 566 1230 582
rect 964 532 965 533
rect 992 532 993 533
rect 1043 532 1044 533
rect 1071 532 1072 533
rect 1122 532 1123 533
rect 1150 532 1151 533
rect 1201 532 1202 533
rect 1229 532 1230 533
rect 914 503 932 532
rect 963 531 994 532
rect 1042 531 1073 532
rect 1121 531 1152 532
rect 1200 531 1231 532
rect 964 524 993 531
rect 1043 524 1072 531
rect 1122 524 1151 531
rect 1201 524 1230 531
rect 964 510 974 524
rect 1221 510 1230 524
rect 964 504 993 510
rect 1043 504 1072 510
rect 1122 504 1151 510
rect 1201 504 1230 510
rect 963 503 994 504
rect 1042 503 1073 504
rect 1121 503 1152 504
rect 1200 503 1231 504
rect 1263 503 1280 532
rect 964 502 965 503
rect 992 502 993 503
rect 1043 502 1044 503
rect 1071 502 1072 503
rect 1122 502 1123 503
rect 1150 502 1151 503
rect 1201 502 1202 503
rect 1229 502 1230 503
rect 964 453 993 468
rect 1043 453 1072 468
rect 1122 453 1151 468
rect 1201 453 1230 468
rect 964 286 993 302
rect 1043 286 1072 302
rect 1122 286 1151 302
rect 1201 286 1230 302
rect 964 252 965 253
rect 992 252 993 253
rect 1043 252 1044 253
rect 1071 252 1072 253
rect 1122 252 1123 253
rect 1150 252 1151 253
rect 1201 252 1202 253
rect 1229 252 1230 253
rect 914 223 932 252
rect 963 251 994 252
rect 1042 251 1073 252
rect 1121 251 1152 252
rect 1200 251 1231 252
rect 964 244 993 251
rect 1043 244 1072 251
rect 1122 244 1151 251
rect 1201 244 1230 251
rect 964 230 974 244
rect 1221 230 1230 244
rect 964 224 993 230
rect 1043 224 1072 230
rect 1122 224 1151 230
rect 1201 224 1230 230
rect 963 223 994 224
rect 1042 223 1073 224
rect 1121 223 1152 224
rect 1200 223 1231 224
rect 1263 223 1280 252
rect 964 222 965 223
rect 992 222 993 223
rect 1043 222 1044 223
rect 1071 222 1072 223
rect 1122 222 1123 223
rect 1150 222 1151 223
rect 1201 222 1202 223
rect 1229 222 1230 223
rect 105 204 134 222
rect 964 173 993 188
rect 1043 173 1072 188
rect 1122 173 1151 188
rect 1201 173 1230 188
rect 105 172 106 173
rect 133 172 134 173
rect 55 143 73 172
rect 104 171 135 172
rect 105 162 134 171
rect 105 153 115 162
rect 124 153 134 162
rect 105 144 134 153
rect 104 143 135 144
rect 166 143 184 172
rect 105 142 106 143
rect 133 142 134 143
rect 964 131 993 147
rect 1043 131 1072 147
rect 1122 131 1151 147
rect 1201 131 1230 147
rect 105 93 134 111
rect 964 97 965 98
rect 992 97 993 98
rect 1043 97 1044 98
rect 1071 97 1072 98
rect 1122 97 1123 98
rect 1150 97 1151 98
rect 1201 97 1202 98
rect 1229 97 1230 98
rect 914 68 932 97
rect 963 96 994 97
rect 1042 96 1073 97
rect 1121 96 1152 97
rect 1200 96 1231 97
rect 964 89 993 96
rect 1043 89 1072 96
rect 1122 89 1151 96
rect 1201 89 1230 96
rect 964 75 974 89
rect 1221 75 1230 89
rect 964 69 993 75
rect 1043 69 1072 75
rect 1122 69 1151 75
rect 1201 69 1230 75
rect 963 68 994 69
rect 1042 68 1073 69
rect 1121 68 1152 69
rect 1200 68 1231 69
rect 1263 68 1280 97
rect 964 67 965 68
rect 992 67 993 68
rect 1043 67 1044 68
rect 1071 67 1072 68
rect 1122 67 1123 68
rect 1150 67 1151 68
rect 1201 67 1202 68
rect 1229 67 1230 68
rect 964 18 993 33
rect 1043 18 1072 33
rect 1122 18 1151 33
rect 1201 18 1230 33
<< nwell >>
rect 916 438 1031 455
rect 1035 438 1086 455
rect 897 320 1297 438
rect 897 319 1086 320
rect 1218 319 1297 320
rect 916 300 1031 319
rect 1035 299 1086 319
rect 1191 300 1218 318
rect 2711 250 2985 600
rect 503 168 525 179
<< mvnmos >>
rect 2600 505 2663 555
rect 2600 283 2663 333
rect 2600 116 2662 193
rect 2745 116 2809 171
rect 2887 116 2951 171
<< mvpmos >>
rect 2748 479 2808 534
rect 2888 479 2948 534
rect 2748 312 2808 367
rect 2888 312 2948 367
<< mvndiff >>
rect 2600 578 2663 582
rect 2600 561 2606 578
rect 2623 561 2640 578
rect 2657 561 2663 578
rect 2600 555 2663 561
rect 2600 492 2663 505
rect 2600 333 2663 338
rect 2600 277 2663 283
rect 2600 260 2605 277
rect 2622 260 2639 277
rect 2656 260 2663 277
rect 2600 254 2663 260
rect 2600 216 2662 224
rect 2600 199 2605 216
rect 2622 199 2639 216
rect 2656 199 2662 216
rect 2600 193 2662 199
rect 2745 194 2809 201
rect 2745 177 2752 194
rect 2769 177 2786 194
rect 2803 177 2809 194
rect 2745 171 2809 177
rect 2887 194 2951 200
rect 2887 177 2893 194
rect 2910 177 2927 194
rect 2944 177 2951 194
rect 2887 171 2951 177
rect 2600 110 2662 116
rect 2600 93 2604 110
rect 2621 93 2638 110
rect 2655 93 2662 110
rect 2600 86 2662 93
rect 2745 110 2809 116
rect 2745 93 2752 110
rect 2769 93 2786 110
rect 2803 93 2809 110
rect 2745 86 2809 93
rect 2887 110 2951 116
rect 2887 93 2893 110
rect 2910 93 2927 110
rect 2944 93 2951 110
rect 2887 87 2951 93
<< mvpdiff >>
rect 2748 557 2808 563
rect 2748 540 2752 557
rect 2769 540 2786 557
rect 2803 540 2808 557
rect 2748 534 2808 540
rect 2888 557 2948 563
rect 2888 540 2893 557
rect 2910 540 2927 557
rect 2944 540 2948 557
rect 2888 534 2948 540
rect 2748 472 2808 479
rect 2748 455 2752 472
rect 2769 455 2786 472
rect 2803 455 2808 472
rect 2748 438 2808 455
rect 2748 390 2808 408
rect 2748 373 2752 390
rect 2769 373 2786 390
rect 2803 373 2808 390
rect 2748 367 2808 373
rect 2888 472 2948 479
rect 2888 455 2893 472
rect 2910 455 2927 472
rect 2944 455 2948 472
rect 2888 438 2948 455
rect 2888 390 2948 408
rect 2888 373 2893 390
rect 2910 373 2927 390
rect 2944 373 2948 390
rect 2888 367 2948 373
rect 2748 306 2808 312
rect 2748 289 2752 306
rect 2769 289 2786 306
rect 2803 289 2808 306
rect 2748 283 2808 289
rect 2888 306 2948 312
rect 2888 289 2893 306
rect 2910 289 2927 306
rect 2944 289 2948 306
rect 2888 283 2948 289
<< mvndiffc >>
rect 2606 561 2623 578
rect 2640 561 2657 578
rect 2605 260 2622 277
rect 2639 260 2656 277
rect 2605 199 2622 216
rect 2639 199 2656 216
rect 2752 177 2769 194
rect 2786 177 2803 194
rect 2893 177 2910 194
rect 2927 177 2944 194
rect 2604 93 2621 110
rect 2638 93 2655 110
rect 2752 93 2769 110
rect 2786 93 2803 110
rect 2893 93 2910 110
rect 2927 93 2944 110
<< mvpdiffc >>
rect 2752 540 2769 557
rect 2786 540 2803 557
rect 2893 540 2910 557
rect 2927 540 2944 557
rect 2752 455 2769 472
rect 2786 455 2803 472
rect 2752 373 2769 390
rect 2786 373 2803 390
rect 2893 455 2910 472
rect 2927 455 2944 472
rect 2893 373 2910 390
rect 2927 373 2944 390
rect 2752 289 2769 306
rect 2786 289 2803 306
rect 2893 289 2910 306
rect 2927 289 2944 306
<< psubdiff >>
rect 379 378 713 383
rect 379 361 419 378
rect 436 361 453 378
rect 470 361 487 378
rect 504 361 521 378
rect 538 361 555 378
rect 572 361 589 378
rect 606 361 623 378
rect 640 361 657 378
rect 674 361 713 378
rect 379 357 713 361
rect 379 338 408 357
rect 379 321 385 338
rect 402 321 408 338
rect 379 309 408 321
rect 263 304 408 309
rect 263 296 385 304
rect 263 279 283 296
rect 300 279 317 296
rect 334 279 351 296
rect 368 287 385 296
rect 402 287 408 304
rect 368 279 408 287
rect 263 271 408 279
rect 379 270 408 271
rect 379 253 385 270
rect 402 253 408 270
rect 379 236 408 253
rect 379 219 385 236
rect 402 219 408 236
rect 379 202 408 219
rect 379 185 385 202
rect 402 185 408 202
rect 379 168 408 185
rect 1360 344 1399 377
rect 1360 327 1372 344
rect 1389 327 1399 344
rect 1360 298 1399 327
rect 1360 281 1372 298
rect 1389 281 1399 298
rect 1360 260 1399 281
rect 1360 243 1372 260
rect 1389 243 1399 260
rect 1360 217 1399 243
rect 1360 200 1372 217
rect 1389 200 1399 217
rect 379 151 385 168
rect 402 151 408 168
rect 379 134 408 151
rect 379 117 385 134
rect 402 117 408 134
rect 379 100 408 117
rect 379 83 385 100
rect 402 83 408 100
rect 1360 162 1399 200
rect 1360 145 1372 162
rect 1389 145 1399 162
rect 1360 122 1399 145
rect 1360 105 1372 122
rect 1389 105 1399 122
rect 379 71 408 83
rect 1360 86 1399 105
rect 1360 69 1372 86
rect 1389 69 1399 86
rect 1360 48 1399 69
rect 1360 31 1371 48
rect 1388 31 1399 48
rect 1360 15 1399 31
<< mvpsubdiff >>
rect 2601 43 2955 49
rect 2601 42 2681 43
rect 2601 25 2613 42
rect 2630 25 2647 42
rect 2664 26 2681 42
rect 2698 26 2717 43
rect 2734 26 2753 43
rect 2770 26 2787 43
rect 2804 26 2821 43
rect 2838 26 2855 43
rect 2872 26 2889 43
rect 2906 26 2923 43
rect 2940 26 2955 43
rect 2664 25 2955 26
rect 2601 19 2955 25
<< mvnsubdiff >>
rect 1223 429 1264 437
rect 1223 416 1235 429
rect 1209 412 1235 416
rect 1252 412 1264 429
rect 1209 395 1264 412
rect 1209 378 1235 395
rect 1252 378 1264 395
rect 1209 377 1264 378
rect 1223 361 1264 377
rect 1223 344 1235 361
rect 1252 344 1264 361
rect 1223 339 1264 344
rect 1224 335 1264 339
rect 2748 431 2808 438
rect 2748 414 2769 431
rect 2786 414 2808 431
rect 2748 408 2808 414
rect 2888 431 2948 438
rect 2888 414 2909 431
rect 2926 414 2948 431
rect 2888 408 2948 414
rect 503 168 525 179
<< psubdiffcont >>
rect 419 361 436 378
rect 453 361 470 378
rect 487 361 504 378
rect 521 361 538 378
rect 555 361 572 378
rect 589 361 606 378
rect 623 361 640 378
rect 657 361 674 378
rect 385 321 402 338
rect 283 279 300 296
rect 317 279 334 296
rect 351 279 368 296
rect 385 287 402 304
rect 385 253 402 270
rect 385 219 402 236
rect 385 185 402 202
rect 1372 327 1389 344
rect 1372 281 1389 298
rect 1372 243 1389 260
rect 1372 200 1389 217
rect 385 151 402 168
rect 385 117 402 134
rect 385 83 402 100
rect 1372 145 1389 162
rect 1372 105 1389 122
rect 1372 69 1389 86
rect 1371 31 1388 48
<< mvpsubdiffcont >>
rect 2613 25 2630 42
rect 2647 25 2664 42
rect 2681 26 2698 43
rect 2717 26 2734 43
rect 2753 26 2770 43
rect 2787 26 2804 43
rect 2821 26 2838 43
rect 2855 26 2872 43
rect 2889 26 2906 43
rect 2923 26 2940 43
<< mvnsubdiffcont >>
rect 1235 412 1252 429
rect 1235 378 1252 395
rect 1235 344 1252 361
rect 2769 414 2786 431
rect 2909 414 2926 431
<< poly >>
rect 204 487 232 537
rect 207 420 232 487
rect 726 457 775 544
rect 2389 542 2600 555
rect 726 455 920 457
rect 1203 455 1254 456
rect 1277 455 1473 542
rect 2388 505 2600 542
rect 2663 505 2676 555
rect 2824 556 2832 572
rect 2824 534 2844 556
rect 2965 555 2974 572
rect 2962 534 2980 555
rect 2388 491 2442 505
rect 2734 479 2748 534
rect 2808 479 2844 534
rect 2872 479 2888 534
rect 2948 479 2980 534
rect 726 420 1072 455
rect 95 396 1072 420
rect 95 217 133 396
rect 726 300 1072 396
rect 2646 399 2693 433
rect 2677 333 2693 399
rect 2824 367 2844 479
rect 2963 367 2980 479
rect 1203 318 1254 319
rect 1191 300 1254 318
rect 726 299 920 300
rect 1021 299 1072 300
rect 726 174 775 299
rect 2585 283 2600 333
rect 2663 283 2693 333
rect 2734 312 2748 367
rect 2808 312 2844 367
rect 2874 312 2888 367
rect 2948 312 2980 367
rect 2688 236 2726 237
rect 726 145 1015 174
rect 2670 198 2726 236
rect 2670 193 2691 198
rect 726 90 775 145
rect 2585 116 2600 193
rect 2662 178 2691 193
rect 2662 116 2676 178
rect 2729 116 2745 171
rect 2809 116 2887 171
rect 2951 116 2964 171
<< locali >>
rect 2598 561 2606 578
rect 2657 561 2665 578
rect 2828 557 2836 572
rect 2965 558 2974 572
rect 2885 557 2985 558
rect 2744 540 2752 557
rect 2803 540 2845 557
rect 2885 540 2893 557
rect 2944 540 2985 557
rect 2744 455 2752 472
rect 2803 455 2893 472
rect 2944 455 2952 472
rect 1235 429 1252 437
rect 2752 414 2769 431
rect 2803 414 2892 431
rect 2926 414 2934 431
rect 1235 402 1252 412
rect 1235 395 1295 402
rect 385 378 402 380
rect 1252 378 1295 395
rect 385 361 419 378
rect 436 361 453 378
rect 470 361 487 378
rect 504 361 521 378
rect 538 361 555 378
rect 572 361 589 378
rect 606 361 623 378
rect 640 361 657 378
rect 674 361 691 378
rect 1235 376 1295 378
rect 1235 361 1252 376
rect 2744 373 2752 390
rect 2803 373 2893 390
rect 2944 373 2952 390
rect 385 338 402 361
rect 1235 336 1252 344
rect 1372 344 1389 355
rect 385 304 402 321
rect 275 279 283 296
rect 300 279 317 296
rect 334 279 351 296
rect 368 287 385 296
rect 368 279 402 287
rect 385 270 402 279
rect 385 236 402 253
rect 385 202 402 219
rect 385 168 402 185
rect 385 134 402 151
rect 385 100 402 117
rect 1372 298 1389 327
rect 2744 289 2752 306
rect 2803 289 2812 306
rect 2885 289 2893 306
rect 2944 289 2952 306
rect 1372 260 1389 281
rect 2597 260 2605 277
rect 2622 260 2639 277
rect 2656 260 2711 277
rect 1372 217 1389 243
rect 1372 162 1389 200
rect 2597 199 2605 216
rect 2656 199 2664 216
rect 2744 177 2752 194
rect 2803 177 2832 194
rect 2885 177 2893 194
rect 2944 177 2952 194
rect 1372 122 1389 145
rect 1372 90 1389 105
rect 2595 93 2604 110
rect 2621 93 2638 110
rect 2655 93 2752 110
rect 2769 93 2786 110
rect 2803 93 2893 110
rect 2910 93 2927 110
rect 2944 93 2953 110
rect 385 38 402 83
rect 1371 86 1389 90
rect 1371 69 1372 86
rect 1371 48 1389 69
rect 1388 31 1389 48
rect 2622 43 2690 48
rect 2622 42 2681 43
rect 1371 17 1389 31
rect 2605 25 2613 42
rect 2630 25 2647 42
rect 2664 26 2681 42
rect 2698 26 2717 43
rect 2734 26 2753 43
rect 2770 26 2787 43
rect 2804 26 2821 43
rect 2838 26 2855 43
rect 2872 26 2889 43
rect 2906 26 2923 43
rect 2940 26 2948 43
rect 2664 25 2690 26
<< viali >>
rect 2623 561 2640 578
rect 2769 540 2786 557
rect 2910 540 2927 557
rect 2769 455 2786 472
rect 2910 455 2927 472
rect 2786 414 2803 431
rect 2892 414 2909 431
rect 2769 373 2786 390
rect 2910 373 2927 390
rect 2769 289 2786 306
rect 2910 289 2927 306
rect 2622 199 2639 216
rect 2769 177 2786 194
rect 2910 177 2927 194
<< metal1 >>
rect 28 516 54 605
rect 498 480 525 605
rect 1085 564 1109 605
rect 2617 578 2646 581
rect 2617 561 2623 578
rect 2640 561 2646 578
rect 2617 558 2646 561
rect 2693 557 2796 565
rect 2693 540 2769 557
rect 2786 540 2796 557
rect 2693 534 2796 540
rect 2899 557 2937 565
rect 2899 540 2910 557
rect 2927 540 2937 557
rect 2899 534 2937 540
rect 2618 489 2645 502
rect 2609 480 2645 489
rect 2609 460 2651 480
rect 2609 366 2632 460
rect 2609 348 2645 366
rect 107 18 132 205
rect 106 0 132 18
rect 497 0 528 259
rect 2618 219 2645 348
rect 2693 257 2717 534
rect 2766 472 2789 478
rect 2766 455 2769 472
rect 2786 455 2789 472
rect 2906 472 2930 478
rect 2906 455 2910 472
rect 2927 455 2930 472
rect 2761 431 2936 455
rect 2761 414 2786 431
rect 2803 414 2892 431
rect 2909 414 2936 431
rect 2761 390 2936 414
rect 2761 389 2769 390
rect 2766 373 2769 389
rect 2786 389 2910 390
rect 2786 373 2789 389
rect 2766 367 2789 373
rect 2906 373 2910 389
rect 2927 389 2936 390
rect 2927 373 2930 389
rect 2906 367 2930 373
rect 2766 306 2789 312
rect 2766 289 2769 306
rect 2786 289 2789 306
rect 2612 216 2645 219
rect 2612 199 2622 216
rect 2639 199 2645 216
rect 2612 196 2645 199
rect 2766 194 2789 289
rect 1086 0 1110 188
rect 2766 177 2769 194
rect 2786 177 2789 194
rect 2766 171 2789 177
rect 2907 306 2930 312
rect 2907 289 2910 306
rect 2927 289 2930 306
rect 2907 194 2930 289
rect 2907 177 2910 194
rect 2927 177 2930 194
rect 2907 171 2930 177
rect 2417 0 2446 106
<< metal2 >>
rect 2616 558 2905 582
rect 1263 459 2728 472
rect 1263 451 2995 459
rect 1086 381 1116 427
rect 1159 382 1189 428
rect 1297 384 1321 451
rect 2714 434 2995 451
rect 2650 300 2677 428
rect 2728 383 2995 434
rect 2650 299 2929 300
rect 2650 277 2995 299
rect 2702 276 2995 277
rect 2933 228 2995 260
rect 2692 189 2995 212
rect 2607 62 2995 95
rect 2606 53 2995 62
rect 2607 46 2995 53
rect 2631 28 2675 46
rect 381 7 2704 28
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_1
timestamp 1628285143
transform 1 0 1475 0 1 814
box -1005 -380 -733 -211
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_2
timestamp 1628285143
transform 1 0 1475 0 1 515
box -1005 -380 -733 -211
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_0
timestamp 1628285143
transform 1 0 1475 0 1 414
box -1005 -380 -733 -211
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_0
timestamp 1628285143
transform 1 0 117 0 1 136
box -62 -43 67 86
use sky130_hilas_FGVaractorTunnelCap01  sky130_hilas_FGVaractorTunnelCap01_0
timestamp 1628285143
transform 1 0 1005 0 1 809
box -1005 -380 -783 -211
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_0
timestamp 1628285143
transform 1 0 1418 0 1 489
box -521 -54 -121 110
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_2
timestamp 1628285143
transform 1 0 1418 0 1 54
box -521 -54 -121 110
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_1
timestamp 1628285143
transform 1 0 1418 0 1 209
box -521 -54 -121 110
use sky130_hilas_li2m2  sky130_hilas_li2m2_14
timestamp 1628285143
transform 1 0 392 0 1 24
box -14 -15 20 18
use sky130_hilas_FGHugeVaractorCapacitor01  sky130_hilas_FGHugeVaractorCapacitor01_0
timestamp 1628285143
transform 1 0 2011 0 1 818
box -556 -816 473 -217
use sky130_hilas_pFETdevice01w1  sky130_hilas_pFETdevice01w1_0
timestamp 1628285143
transform 1 0 1136 0 1 396
box -79 -78 82 43
use sky130_hilas_li2m2  sky130_hilas_li2m2_11
timestamp 1628285143
transform 1 0 1306 0 1 388
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_12
timestamp 1628285143
transform 1 0 1170 0 1 396
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_13
timestamp 1628285143
transform 1 0 1101 0 1 395
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628285143
transform 1 0 1378 0 1 22
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_9
timestamp 1628285143
transform 1 0 2618 0 1 39
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_4
timestamp 1628285143
transform 1 0 2704 0 1 100
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_5
timestamp 1628285143
transform 1 0 2689 0 1 40
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_6
timestamp 1628285143
transform 1 0 2763 0 1 40
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1628285143
transform 1 0 2847 0 1 98
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_7
timestamp 1628285143
transform 1 0 2833 0 1 40
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_8
timestamp 1628285143
transform 1 0 2926 0 1 40
box -14 -15 20 18
use sky130_hilas_poly2li  sky130_hilas_poly2li_5
timestamp 1628285143
transform -1 0 2717 0 -1 221
box -9 -14 18 19
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1628285143
transform 1 0 2703 0 1 265
box -10 -8 13 21
use sky130_hilas_li2m2  sky130_hilas_li2m2_10
timestamp 1628285143
transform -1 0 2707 0 -1 220
box -14 -15 20 18
use sky130_hilas_poly2li  sky130_hilas_poly2li_3
timestamp 1628285143
transform 1 0 2833 0 1 181
box -9 -14 18 19
use sky130_hilas_m12m2  sky130_hilas_m12m2_9
timestamp 1628285143
transform 1 0 2912 0 1 238
box -9 -10 23 22
use sky130_hilas_nDiffThOxContact  sky130_hilas_nDiffThOxContact_3
timestamp 1628704229
transform 1 0 2624 0 1 321
box 0 0 67 29
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_0
timestamp 1628285143
transform 1 0 2655 0 1 407
box -9 -26 24 29
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1628285143
transform 1 0 2771 0 1 417
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_4
timestamp 1628285143
transform 1 0 2769 0 1 375
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_6
timestamp 1628285143
transform 1 0 2771 0 1 461
box -9 -10 23 22
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628285143
transform 1 0 2845 0 1 378
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1628285143
transform 1 0 2845 0 1 462
box -14 -15 20 18
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1628285143
transform 1 0 2912 0 1 415
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_2
timestamp 1628285143
transform 1 0 2912 0 1 460
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_3
timestamp 1628285143
transform 1 0 2912 0 1 373
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_10
timestamp 1628285143
transform 1 0 2625 0 1 568
box -9 -10 23 22
use sky130_hilas_nDiffThOxContact  sky130_hilas_nDiffThOxContact_0
timestamp 1628704229
transform 1 0 2624 0 1 464
box 0 0 67 29
use sky130_hilas_poly2li  sky130_hilas_poly2li_1
timestamp 1628285143
transform 1 0 2836 0 1 569
box -9 -14 18 19
use sky130_hilas_poly2li  sky130_hilas_poly2li_4
timestamp 1628285143
transform 1 0 2976 0 1 569
box -9 -14 18 19
use sky130_hilas_m12m2  sky130_hilas_m12m2_7
timestamp 1628285143
transform 1 0 2911 0 1 563
box -9 -10 23 22
<< labels >>
rlabel metal2 2989 46 2995 95 0 VGND
port 8 nsew ground default
rlabel metal2 2989 228 2995 260 0 OUTPUT
port 10 nsew analog default
rlabel metal2 2988 383 2995 459 0 VINJ
port 9 nsew power default
rlabel metal2 2989 189 2995 212 0 VBIAS
port 12 nsew analog default
rlabel metal2 2989 276 2995 299 0 VREF
port 11 nsew analog default
rlabel metal1 2417 2 2446 7 0 LARGECAPACITOR
port 7 nsew analog default
rlabel metal1 1085 599 1109 605 0 GATE3
port 3 nsew analog default
rlabel metal1 1086 0 1110 7 0 GATE4
port 6 nsew analog default
rlabel metal1 497 0 528 7 0 GATE2
port 5 nsew analog default
rlabel metal1 498 596 525 605 0 GATE1
port 2 nsew analog default
rlabel metal1 106 0 132 10 0 VTUNOVERLAP01
port 4 nsew analog default
rlabel metal1 28 598 54 605 0 VTUN
port 1 nsew analog default
rlabel metal2 1086 416 1116 427 0 DRAIN1
port 13 nsew
rlabel metal2 1159 417 1188 428 0 SOURCE1
port 14 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
