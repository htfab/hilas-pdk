magic
tech sky130A
timestamp 1627759641
<< error_s >>
rect 35 489 85 500
rect 85 483 119 489
rect 368 486 418 495
rect 418 480 449 486
rect 525 480 553 496
rect 667 480 695 496
rect 35 447 85 458
rect 636 454 641 459
rect 184 446 201 451
rect 368 444 418 453
rect 525 438 553 454
rect 667 438 695 454
rect 106 427 156 438
rect 296 418 347 428
rect 264 413 283 418
rect 476 417 504 434
rect 716 417 744 434
rect 156 396 188 401
rect 106 385 156 396
rect 264 386 269 413
rect 347 386 378 392
rect 296 376 347 386
rect 476 375 504 392
rect 716 375 744 392
rect 35 334 85 345
rect 85 328 119 334
rect 368 331 418 340
rect 418 325 449 331
rect 525 325 553 341
rect 667 325 695 341
rect 35 292 85 303
rect 636 299 641 304
rect 184 291 201 296
rect 368 289 418 298
rect 525 283 553 299
rect 667 283 695 299
rect 106 272 156 283
rect 296 263 347 273
rect 264 258 283 263
rect 476 262 504 279
rect 716 262 744 279
rect 156 241 188 246
rect 106 230 156 241
rect 264 231 269 258
rect 347 231 378 237
rect 296 221 347 231
rect 476 220 504 237
rect 716 220 744 237
rect 35 179 85 190
rect 85 173 119 179
rect 368 176 418 185
rect 418 170 449 176
rect 525 170 553 186
rect 667 170 695 186
rect 35 137 85 148
rect 636 144 641 149
rect 184 136 201 141
rect 368 134 418 143
rect 525 128 553 144
rect 667 128 695 144
rect 106 117 156 128
rect 296 108 347 118
rect 264 103 283 108
rect 476 107 504 124
rect 716 107 744 124
rect 156 86 188 91
rect 106 75 156 86
rect 264 76 269 103
rect 347 76 378 82
rect 296 66 347 76
rect 476 65 504 82
rect 716 65 744 82
rect 35 24 85 35
rect 85 18 119 24
rect 368 21 418 30
rect 418 15 449 21
rect 525 15 553 31
rect 667 15 695 31
rect 35 -18 85 -7
rect 636 -11 641 -6
rect 184 -19 201 -14
rect 368 -21 418 -12
rect 525 -27 553 -11
rect 667 -27 695 -11
rect 106 -38 156 -27
rect 296 -47 347 -37
rect 264 -52 283 -47
rect 476 -48 504 -31
rect 716 -48 744 -31
rect 156 -69 188 -64
rect 106 -80 156 -69
rect 264 -79 269 -52
rect 347 -79 378 -73
rect 296 -89 347 -79
rect 476 -90 504 -73
rect 716 -90 744 -73
use sky130_hilas_StepUpDigital  StepUpDigital_3
timestamp 1627759641
transform 1 0 -49 0 1 -62
box 19 -40 899 119
use sky130_hilas_StepUpDigital  StepUpDigital_0
timestamp 1627759641
transform 1 0 -49 0 1 93
box 19 -40 899 119
use sky130_hilas_StepUpDigital  StepUpDigital_1
timestamp 1627759641
transform 1 0 -49 0 1 248
box 19 -40 899 119
use sky130_hilas_StepUpDigital  StepUpDigital_2
timestamp 1627759641
transform 1 0 -49 0 1 403
box 19 -40 899 119
<< labels >>
rlabel metal2 841 372 850 404 0 INPUT1
port 1 nsew
rlabel metal2 841 217 850 249 0 INPUT2
port 2 nsew
rlabel metal2 841 62 850 94 0 INPUT3
port 3 nsew
rlabel metal2 841 -93 850 -61 0 INPUT4
port 4 nsew
rlabel metal1 746 517 770 522 0 VPWR
port 5 nsew
rlabel metal1 746 -102 770 -97 0 VPWR
port 5 nsew
rlabel metal1 4 517 33 522 0 VINJ
port 6 nsew
rlabel metal1 4 -102 33 -97 0 VINJ
port 6 nsew
rlabel metal2 -30 470 -19 490 0 OUTPUT1
port 7 nsew
rlabel metal2 -30 315 -19 335 0 OUTPUT2
port 8 nsew
rlabel metal2 -30 160 -19 180 0 OUTPUT3
port 9 nsew
rlabel metal2 -30 5 -19 25 0 OUTPUT4
port 10 nsew
rlabel metal1 445 515 476 522 0 VGND
port 11 nsew
rlabel metal1 445 -102 476 -96 0 VGND
port 11 nsew
<< end >>
