magic
tech sky130A
timestamp 1607701799
<< metal2 >>
rect -14 18 23 24
rect -14 -10 -9 18
rect 19 -10 23 18
rect -14 -16 23 -10
<< via2 >>
rect -9 -10 19 18
<< metal3 >>
rect -36 27 43 39
rect -36 -21 -17 27
rect 26 -21 43 27
rect -36 -36 43 -21
<< via3 >>
rect -17 18 26 27
rect -17 -10 -9 18
rect -9 -10 19 18
rect 19 -10 26 18
rect -17 -21 26 -10
<< metal4 >>
rect -27 27 39 36
rect -27 -21 -17 27
rect 26 -21 39 27
rect -27 -30 39 -21
<< end >>
