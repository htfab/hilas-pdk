magic
tech sky130A
timestamp 1628616721
<< checkpaint >>
rect -352 -630 1522 799
<< error_s >>
rect 87 135 137 141
rect 410 136 460 142
rect 567 135 595 142
rect 709 136 737 142
rect 87 93 137 99
rect 410 94 460 100
rect 567 93 595 100
rect 709 94 737 100
rect 158 69 208 75
rect 338 64 389 70
rect 518 64 546 70
rect 758 64 786 70
rect 158 27 208 33
rect 338 22 389 28
rect 518 22 546 28
rect 758 22 786 28
<< nwell >>
rect 22 0 272 175
rect 659 168 836 175
rect 659 0 836 9
<< mvpmos >>
rect 87 99 137 135
rect 158 33 208 69
<< mvpdiff >>
rect 56 123 87 135
rect 56 106 64 123
rect 81 106 87 123
rect 56 99 87 106
rect 137 124 171 135
rect 137 107 143 124
rect 160 107 171 124
rect 137 99 171 107
rect 127 60 158 69
rect 127 43 133 60
rect 151 43 158 60
rect 127 33 158 43
rect 208 62 239 69
rect 208 45 214 62
rect 232 45 239 62
rect 208 33 239 45
<< mvpdiffc >>
rect 64 106 81 123
rect 143 107 160 124
rect 133 43 151 60
rect 214 45 232 62
<< mvnsubdiff >>
rect 57 60 127 69
rect 57 43 83 60
rect 100 43 127 60
rect 57 33 127 43
<< mvnsubdiffcont >>
rect 83 43 100 60
<< poly >>
rect 87 143 237 158
rect 87 135 137 143
rect 210 131 237 143
rect 210 114 215 131
rect 232 114 237 131
rect 210 104 237 114
rect 264 129 298 134
rect 264 112 273 129
rect 290 112 298 129
rect 264 104 298 112
rect 87 84 137 99
rect 158 69 208 83
rect 264 70 280 104
rect 248 46 280 70
rect 158 25 208 33
rect 248 25 264 46
rect 158 10 264 25
<< polycont >>
rect 215 114 232 131
rect 273 112 290 129
<< locali >>
rect 150 131 195 139
rect 150 124 167 131
rect 56 106 64 123
rect 81 106 89 123
rect 135 107 143 124
rect 160 114 167 124
rect 184 114 195 131
rect 160 107 195 114
rect 215 131 232 139
rect 63 97 81 106
rect 80 80 81 97
rect 63 61 81 80
rect 215 63 232 114
rect 265 129 294 132
rect 265 127 273 129
rect 265 110 271 127
rect 290 112 298 129
rect 288 110 294 112
rect 265 108 294 110
rect 215 62 253 63
rect 80 60 81 61
rect 80 44 83 60
rect 63 43 83 44
rect 100 43 133 60
rect 151 43 159 60
rect 206 45 214 62
rect 232 56 253 62
rect 232 51 287 56
rect 232 45 288 51
rect 214 39 288 45
rect 214 34 253 39
<< viali >>
rect 167 114 184 131
rect 63 80 80 97
rect 271 112 273 127
rect 273 112 288 127
rect 271 110 288 112
rect 63 44 80 61
<< metal1 >>
rect 56 97 85 175
rect 487 169 518 175
rect 788 168 812 175
rect 160 136 192 139
rect 160 110 163 136
rect 189 110 192 136
rect 265 132 296 133
rect 160 109 192 110
rect 264 106 267 132
rect 293 106 296 132
rect 264 105 296 106
rect 265 104 294 105
rect 56 80 63 97
rect 80 80 85 97
rect 56 61 85 80
rect 56 44 63 61
rect 80 44 85 61
rect 56 0 85 44
<< via1 >>
rect 163 131 189 136
rect 163 114 167 131
rect 167 114 184 131
rect 184 114 189 131
rect 163 110 189 114
rect 267 127 293 132
rect 267 110 271 127
rect 271 110 288 127
rect 288 110 293 127
rect 267 106 293 110
<< metal2 >>
rect 160 131 163 136
rect 29 111 163 131
rect 160 110 163 111
rect 189 131 192 136
rect 263 132 295 133
rect 263 131 267 132
rect 189 111 267 131
rect 189 110 192 111
rect 263 106 267 111
rect 293 106 296 132
rect 263 104 295 106
use sky130_hilas_StepUpDigitalPart1  StepUpDigitalPart1_0
timestamp 1628616705
transform 1 0 0 0 1 49
box 0 0 614 169
<< labels >>
rlabel metal2 29 111 36 131 0 Output
rlabel metal1 56 155 85 163 0 Vinj
rlabel metal1 56 4 85 12 0 Vinj
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
