VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_swc4x1BiasCell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc4x1BiasCell ;
  ORIGIN 2.660 3.820 ;
  SIZE 10.110 BY 6.050 ;
  PIN bias1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -2.640 1.110 -2.490 1.300 ;
    END
  END bias1
  PIN bias2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -2.660 0.120 -2.520 0.320 ;
    END
  END bias2
  PIN bias3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -2.630 -1.870 5.000 -1.710 ;
    END
  END bias3
  PIN bias4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -2.630 -2.860 5.000 -2.690 ;
    END
  END bias4
  PIN Vtun
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT -2.280 -0.670 -1.880 2.230 ;
    END
    PORT
      LAYER met1 ;
        RECT -2.280 -3.820 -1.880 -0.940 ;
    END
  END Vtun
  PIN Gate
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 1.770 -3.820 2.150 -1.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.770 -0.740 2.150 2.230 ;
    END
  END Gate
  PIN Vinj
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 6.920 1.520 7.080 2.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.920 -3.810 7.080 -3.100 ;
    END
  END Vinj
  PIN Vdd
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 6.110 1.490 6.270 2.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.110 -3.810 6.270 -3.070 ;
    END
  END Vdd
  PIN GateSelect
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 6.480 -3.810 6.670 -2.820 ;
    END
  END GateSelect
  PIN drain1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.260 1.550 7.440 1.730 ;
    END
  END drain1
  PIN Horiz1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.260 1.120 7.440 1.300 ;
    END
  END Horiz1
  PIN Horiz2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.260 0.120 7.450 0.300 ;
    END
  END Horiz2
  PIN drain2
    PORT
      LAYER met2 ;
        RECT 5.260 -0.310 7.440 -0.130 ;
    END
  END drain2
  PIN drain3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.260 -1.460 7.450 -1.280 ;
    END
  END drain3
  PIN Horiz3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.260 -1.890 7.440 -1.710 ;
    END
  END Horiz3
  PIN Horiz4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.260 -2.880 7.440 -2.700 ;
    END
  END Horiz4
  PIN drain4
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 5.260 -3.310 7.440 -3.130 ;
    END
  END drain4
  OBS
      LAYER li1 ;
        RECT -2.210 -3.480 7.050 1.900 ;
      LAYER met1 ;
        RECT -1.600 -3.440 1.490 2.230 ;
        RECT 2.430 1.210 5.830 2.230 ;
        RECT 6.550 1.240 6.640 2.230 ;
        RECT 6.550 1.210 7.090 1.240 ;
        RECT 2.430 -2.540 7.090 1.210 ;
        RECT 2.430 -2.790 6.200 -2.540 ;
        RECT 2.430 -3.440 5.830 -2.790 ;
        RECT 6.950 -2.820 7.090 -2.540 ;
      LAYER met2 ;
        RECT -2.620 1.580 4.980 1.870 ;
        RECT -2.210 0.840 4.980 1.580 ;
        RECT -2.210 0.830 5.280 0.840 ;
        RECT -2.620 0.600 5.280 0.830 ;
        RECT -2.240 0.580 5.280 0.600 ;
        RECT -2.240 -0.160 4.980 0.580 ;
        RECT -2.620 -0.590 4.980 -0.160 ;
        RECT -2.620 -1.000 5.280 -0.590 ;
        RECT -2.620 -1.430 4.980 -1.000 ;
        RECT -2.620 -2.170 4.980 -2.150 ;
        RECT -2.620 -2.410 5.280 -2.170 ;
        RECT -2.620 -3.450 4.980 -3.140 ;
  END
END sky130_hilas_swc4x1BiasCell
END LIBRARY

