magic
tech sky130A
magscale 1 2
timestamp 1632256350
<< checkpaint >>
rect -1260 2404 5310 4234
rect -1260 -468 6644 2404
rect 3558 -1184 6644 -468
<< error_s >>
rect 968 2746 1032 2756
rect 968 2628 1032 2646
rect 1050 2468 1116 2474
rect 1032 2374 1044 2398
rect 968 2340 1044 2374
rect 1202 2174 1384 2428
rect 1456 2118 1638 2174
rect 1456 2106 1690 2118
rect 1734 2106 1834 2118
rect 968 2096 1032 2098
rect 1456 2034 1638 2106
rect 1832 2034 1892 2038
rect 1456 2022 1690 2034
rect 1734 2026 1892 2034
rect 1734 2022 1834 2026
rect 2106 2024 2138 2052
rect 2188 2024 2226 2052
rect 2268 2024 2300 2052
rect 1456 1996 1638 2022
rect 1860 2002 1920 2010
rect 1860 1998 1916 2002
rect 968 1970 1032 1996
rect 1202 1938 1384 1996
rect 1186 1920 1384 1938
rect 1202 1884 1384 1920
rect 1186 1866 1384 1884
rect 968 1826 1032 1828
rect 1202 1742 1384 1866
rect 1456 1976 1968 1996
rect 1456 1940 1978 1976
rect 2034 1944 2062 1980
rect 1456 1792 1968 1940
rect 2034 1858 2062 1894
rect 2964 1854 3186 1902
rect 968 1700 1032 1726
rect 1456 1582 1638 1742
rect 1734 1638 1834 1650
rect 1934 1594 1968 1704
rect 2034 1640 2062 1676
rect 1734 1554 1834 1566
rect 1934 1558 1978 1594
rect 1860 1532 1916 1536
rect 1860 1524 1920 1532
rect 1832 1496 1892 1508
rect 1864 1466 1916 1474
rect 1536 1454 1576 1466
rect 1832 1454 1916 1466
rect 1832 1420 1854 1432
rect 1864 1412 1916 1454
rect 1934 1450 1968 1558
rect 2022 1452 2392 1616
rect 2528 1566 2546 1718
rect 2898 1668 3252 1854
rect 3816 1844 3934 1914
rect 3750 1680 4000 1844
rect 2546 1558 2696 1566
rect 2522 1550 2696 1558
rect 2522 1530 2550 1550
rect 2022 1448 2234 1452
rect 2248 1448 2392 1452
rect 2106 1442 2138 1448
rect 2162 1444 2392 1448
rect 2162 1442 2168 1444
rect 2188 1428 2392 1444
rect 2210 1402 2216 1422
rect 2242 1418 2268 1428
rect 2242 1412 2258 1418
rect 1832 1378 1892 1390
rect 1860 1354 1920 1362
rect 1860 1350 1916 1354
rect 1456 1328 1968 1346
rect 1456 1292 1978 1328
rect 2034 1296 2062 1332
rect 1456 1144 1968 1292
rect 2396 1262 3074 1404
rect 2034 1210 2062 1246
rect 2396 1238 3186 1262
rect 2396 1204 2482 1238
rect 2564 1236 3186 1238
rect 2564 1224 2666 1236
rect 2564 1206 2650 1224
rect 2600 1204 2650 1206
rect 1734 988 1834 1000
rect 2034 990 2062 1026
rect 2564 982 2650 1204
rect 2680 1196 2694 1236
rect 2796 1224 2828 1236
rect 2964 1228 3186 1236
rect 3620 1238 3696 1386
rect 2964 1212 3224 1228
rect 3620 1218 3788 1238
rect 2964 1200 3186 1212
rect 2964 1198 3196 1200
rect 2898 1160 3252 1198
rect 3816 1194 3934 1266
rect 4426 1238 4506 1378
rect 4506 1210 4594 1238
rect 2898 1134 3476 1160
rect 2898 1132 3252 1134
rect 2898 1106 3476 1132
rect 2898 1028 3252 1106
rect 3750 1032 4000 1194
rect 5088 990 5170 1006
rect 1734 904 1834 916
rect 1950 908 1978 944
rect 2034 904 2062 940
rect 1860 882 1916 886
rect 1860 874 1920 882
rect 1590 850 1690 862
rect 1734 858 1834 862
rect 1734 850 1892 858
rect 1832 846 1892 850
rect 2106 830 2138 858
rect 2188 830 2226 858
rect 2268 830 2300 858
rect 2394 852 2482 936
rect 2562 852 2650 982
rect 3100 950 3114 968
rect 3128 966 3142 990
rect 3118 950 3142 966
rect 5054 984 5170 990
rect 5174 984 5276 990
rect 5054 966 5276 984
rect 5054 942 5062 966
rect 5088 962 5214 966
rect 5082 954 5304 962
rect 5082 938 5140 954
rect 5082 914 5086 938
rect 5088 912 5140 938
rect 5156 938 5304 954
rect 5156 926 5214 938
rect 5156 912 5171 926
rect 5088 906 5148 912
rect 5082 904 5148 906
rect 5150 908 5182 912
rect 5082 898 5146 904
rect 5082 896 5144 898
rect 5082 876 5144 878
rect 5082 870 5146 876
rect 5150 870 5202 908
rect 5082 868 5202 870
rect 4574 856 4576 868
rect 5088 866 5202 868
rect 5268 866 5302 908
rect 5380 866 5414 908
rect 5494 866 5528 908
rect 5562 866 5596 908
rect 5088 862 5182 866
rect 1590 766 1690 778
rect 1734 766 1834 778
rect 2394 768 2460 852
rect 2562 790 2628 852
rect 4738 816 4760 840
rect 4766 812 4788 816
rect 5054 812 5062 832
rect 5082 812 5086 860
rect 5088 848 5171 862
rect 5088 818 5214 848
rect 5118 790 5214 818
rect 2562 728 2650 790
rect 5118 768 5170 790
rect 2448 310 2560 326
rect 2470 282 2532 298
rect 2456 248 2472 272
rect 2564 30 2650 728
rect 3100 626 3150 642
rect 3100 622 3134 626
rect 3128 598 3178 614
rect 3128 594 3162 598
rect 5054 590 5100 630
rect 5306 590 5352 632
rect 5088 436 5170 452
rect 5054 430 5170 436
rect 5174 430 5276 436
rect 5054 412 5276 430
rect 5054 388 5062 412
rect 5088 408 5214 412
rect 5082 400 5304 408
rect 5082 384 5140 400
rect 5082 360 5086 384
rect 5088 358 5140 384
rect 5156 384 5304 400
rect 5156 376 5280 384
rect 5156 372 5214 376
rect 5156 358 5171 372
rect 5198 368 5204 372
rect 5242 368 5244 376
rect 5242 366 5246 368
rect 5242 364 5250 366
rect 5088 350 5148 358
rect 5150 354 5182 358
rect 5186 354 5252 364
rect 5270 354 5278 376
rect 5082 344 5146 350
rect 5150 348 5252 354
rect 5082 318 5146 322
rect 5150 318 5202 348
rect 5242 318 5250 348
rect 5082 316 5252 318
rect 5088 312 5252 316
rect 5268 312 5302 354
rect 5380 312 5414 354
rect 5494 312 5528 354
rect 5562 312 5596 354
rect 5088 308 5182 312
rect 5054 258 5062 278
rect 5082 258 5086 306
rect 5088 294 5171 308
rect 5186 306 5252 312
rect 5242 302 5250 306
rect 5088 290 5214 294
rect 5270 290 5278 312
rect 5088 278 5280 290
rect 5088 264 5214 278
rect 5270 274 5278 278
rect 5118 236 5214 264
rect 5118 214 5170 236
rect 3620 28 3696 56
rect 4946 28 4992 78
rect 5198 28 5244 78
<< nwell >>
rect 2482 1236 3074 1238
rect 2482 1206 2564 1236
rect 3620 1218 3696 1238
rect 4426 1210 4506 1238
rect 2482 1204 2600 1206
rect 2482 852 2564 1204
rect 2460 768 2564 852
rect 2460 728 2562 768
rect 2460 622 2564 728
rect 2482 30 2564 622
<< poly >>
rect 5102 1146 5142 1238
rect 5102 28 5142 78
<< locali >>
rect 2454 64 2490 248
<< metal1 >>
rect 2634 1224 2666 1238
rect 2716 1224 2754 1238
rect 2796 1224 2828 1238
rect 3620 1218 3696 1238
rect 4426 1182 4506 1238
rect 4946 1146 4992 1238
rect 5198 1146 5244 1238
rect 3120 974 3162 1122
rect 2460 622 2502 852
rect 3116 300 3148 600
rect 5198 368 5244 378
rect 5190 366 5246 368
rect 5190 362 5250 366
rect 5190 308 5192 362
rect 5246 308 5250 362
rect 5190 302 5250 308
rect 3620 28 3696 48
rect 4946 28 4992 78
rect 5198 28 5244 78
<< via1 >>
rect 5192 308 5246 362
<< metal2 >>
rect 2452 1144 2598 1180
rect 3168 1138 4698 1176
rect 3168 1134 4732 1138
rect 4656 1096 4732 1134
rect 4554 1094 4582 1096
rect 2460 968 2490 1052
rect 4554 1028 4584 1094
rect 4554 988 4796 1028
rect 2460 950 3114 968
rect 5024 966 5276 998
rect 2460 938 3146 950
rect 3086 918 3146 938
rect 2456 818 2520 872
rect 4576 856 4816 876
rect 4574 840 4816 856
rect 4760 816 4816 840
rect 4760 812 4766 816
rect 2446 754 2562 790
rect 5024 780 5276 812
rect 3102 722 3148 724
rect 3102 716 4616 722
rect 3102 682 4628 716
rect 3102 662 3150 682
rect 2460 626 3150 662
rect 4590 642 4732 682
rect 2460 622 3134 626
rect 3130 582 4620 586
rect 3130 542 4732 582
rect 3130 540 3194 542
rect 2452 496 2562 532
rect 2448 350 2488 450
rect 4572 418 4772 450
rect 5024 412 5276 444
rect 5186 362 5252 364
rect 2448 310 3158 350
rect 5186 346 5192 362
rect 3916 312 5192 346
rect 5186 308 5192 312
rect 5246 308 5252 362
rect 5186 306 5252 308
rect 2446 208 2502 262
rect 4574 222 4774 256
rect 5028 226 5276 258
rect 4574 220 4762 222
rect 2448 104 2562 140
rect 4620 130 4730 132
rect 3104 86 4730 130
rect 3104 84 4622 86
rect 3104 82 3258 84
rect 2456 48 2524 74
rect 3104 48 3152 82
rect 2456 32 3152 48
rect 2478 0 3152 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_5
timestamp 1632251372
transform 1 0 3102 0 1 320
box 0 0 64 64
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1632251372
transform 1 0 2470 0 1 630
box 0 0 64 64
use sky130_hilas_m12m2  sky130_hilas_m12m2_3
timestamp 1632251372
transform 1 0 2474 0 1 832
box 0 0 64 64
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1632251372
transform 1 0 3132 0 1 1142
box 0 0 64 64
use sky130_hilas_m12m2  sky130_hilas_m12m2_2
timestamp 1632251372
transform 1 0 3128 0 1 932
box 0 0 64 64
use sky130_hilas_m12m2  sky130_hilas_m12m2_4
timestamp 1632251372
transform 1 0 3128 0 1 556
box 0 0 64 64
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1632251356
transform 1 0 2480 0 1 40
box 0 0 68 66
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1632251356
transform 1 0 2470 0 1 232
box 0 0 68 66
use sky130_hilas_WTA4stage01  sky130_hilas_WTA4stage01_0
timestamp 1632256327
transform 1 0 4818 0 1 76
box 0 0 566 1068
use sky130_hilas_swc4x1BiasCell  sky130_hilas_swc4x1BiasCell_0
timestamp 1632256328
transform -1 0 4050 0 1 792
box 0 0 4050 2182
<< labels >>
rlabel metal2 5262 966 5276 998 0 OUTPUT1
port 4 nsew analog default
rlabel metal2 5266 780 5276 812 0 OUTPUT2
port 5 nsew analog default
rlabel metal2 5266 412 5276 444 0 OUTPUT3
port 6 nsew analog default
rlabel metal2 5266 226 5276 258 0 OUTPUT4
port 7 nsew analog default
rlabel metal1 5198 1226 5244 1238 0 VGND
port 1 nsew ground default
rlabel metal1 5198 28 5244 40 0 VGND
port 1 nsew ground default
rlabel metal2 2460 1012 2490 1052 0 INPUT1
port 8 nsew analog default
rlabel metal2 2460 818 2512 870 0 INPUT2
port 9 nsew analog default
rlabel metal2 2448 416 2488 450 0 INPUT3
port 10 nsew analog default
rlabel metal2 2446 208 2502 262 0 INPUT4
port 11 nsew analog default
rlabel metal1 3622 1218 3694 1238 0 GATE1
port 16 nsew
rlabel metal1 4426 1210 4506 1238 0 VTUN
port 17 nsew
rlabel metal1 4946 28 4992 40 0 WTAMIDDLENODE
port 18 nsew
rlabel metal1 4946 1226 4992 1238 0 WTAMIDDLENODE
port 18 nsew
rlabel metal1 2716 1224 2754 1238 0 COLSEL1
port 19 nsew
rlabel metal1 2634 1224 2666 1238 0 VINJ
port 21 nsew
rlabel metal1 2796 1224 2828 1238 0 VPWR
port 20 nsew
rlabel metal2 2452 1144 2470 1180 0 DRAIN1
port 12 nsew
rlabel metal2 2446 754 2464 790 0 DRAIN2
port 22 nsew
rlabel metal2 2452 496 2470 532 0 DRAIN3
port 23 nsew
rlabel metal2 2448 104 2466 140 0 DRAIN4
port 24 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
