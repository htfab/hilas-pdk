magic
tech sky130A
timestamp 1637974713
<< error_s >>
rect 766 617 818 623
rect 818 616 846 617
rect 1120 616 1170 621
rect 766 575 818 581
rect 1120 574 1170 579
rect 692 550 745 555
rect 839 550 891 555
rect 1049 549 1099 555
rect 1191 549 1241 555
rect 84 542 137 549
rect 263 541 315 549
rect 692 508 745 513
rect 839 508 891 513
rect 1049 507 1099 513
rect 1191 507 1241 513
rect 84 500 137 507
rect 263 499 315 507
rect 766 457 818 463
rect 818 456 846 457
rect 1120 456 1170 461
rect 766 415 818 421
rect 1120 414 1170 419
rect 84 391 137 398
rect 263 390 315 398
rect 692 390 745 395
rect 839 390 891 395
rect 1049 389 1099 395
rect 1191 389 1241 395
rect 84 349 137 356
rect 263 348 315 356
rect 692 348 745 353
rect 839 348 891 353
rect 1049 347 1099 353
rect 1191 347 1241 353
rect 766 297 818 303
rect 818 296 846 297
rect 1120 296 1170 301
rect 766 255 818 261
rect 1120 254 1170 259
rect 84 240 137 247
rect 263 239 315 247
rect 692 230 745 235
rect 839 230 891 235
rect 1049 229 1099 235
rect 1191 229 1241 235
rect 84 198 137 205
rect 263 197 315 205
rect 692 188 745 193
rect 839 188 891 193
rect 1049 187 1099 193
rect 1191 187 1241 193
rect 766 137 818 143
rect 818 136 846 137
rect 1120 136 1170 141
rect 766 95 818 101
rect 1120 94 1170 99
rect 692 70 745 75
rect 839 70 891 75
rect 1049 69 1099 75
rect 1191 69 1241 75
rect 692 28 745 33
rect 839 28 891 33
rect 1049 27 1099 33
rect 1191 27 1241 33
<< metal1 >>
rect -73 452 -51 1641
rect -79 449 -51 452
rect -53 423 -51 449
rect -79 420 -51 423
rect -73 -963 -51 420
rect -27 603 -5 1641
rect 61 611 83 1641
rect 318 615 341 1641
rect 669 624 691 1642
rect 1166 623 1193 1641
rect -27 600 -1 603
rect -27 571 -1 574
rect -27 -963 -5 571
rect 61 -963 83 22
rect 318 -962 341 23
rect 669 -961 691 22
rect 1166 -960 1193 27
<< via1 >>
rect -79 423 -53 449
rect -27 574 -1 600
<< metal2 >>
rect 1311 1268 1462 1286
rect -30 574 -27 600
rect -1 596 2 600
rect -1 578 18 596
rect 1311 589 1331 1268
rect -1 574 2 578
rect 1317 515 1331 589
rect 1348 618 1462 636
rect -82 423 -79 449
rect -53 445 -50 449
rect -53 427 18 445
rect -53 423 -50 427
rect 1348 376 1362 618
rect 1318 369 1362 376
rect 1317 355 1362 369
rect -86 276 18 294
rect 1319 211 1362 213
rect 1317 197 1362 211
rect 1319 195 1362 197
rect 1317 -664 1334 53
rect 1348 -14 1362 195
rect 1348 -32 1462 -14
rect 1317 -682 1462 -664
use sky130_hilas_VinjDecode2to4  sky130_hilas_VinjDecode2to4_0
timestamp 1637953024
transform 1 0 637 0 1 -31
box -637 31 694 681
<< labels >>
rlabel metal2 -86 276 -79 294 0 SELECT
port 1 nsew
rlabel metal1 -73 -963 -51 -956 0 A2
port 2 nsew
rlabel metal1 -27 -963 -5 -956 0 A3
port 3 nsew
<< end >>
