magic
tech sky130A
timestamp 1628616971
<< checkpaint >>
rect 1353 1613 3642 2047
rect 817 1608 3642 1613
rect 347 1233 3642 1608
rect -188 1228 3642 1233
rect -658 188 3642 1228
rect -658 -61 3605 188
rect -658 -75 3596 -61
rect -658 -201 3562 -75
rect -603 -537 3562 -201
rect -280 -590 3562 -537
rect -280 -605 3548 -590
rect -280 -606 3240 -605
rect -280 -621 3086 -606
rect 239 -628 3086 -621
rect 239 -630 1899 -628
<< error_s >>
rect 936 566 965 582
rect 1015 566 1044 582
rect 1094 566 1123 582
rect 1173 566 1202 582
rect 936 532 937 533
rect 964 532 965 533
rect 1015 532 1016 533
rect 1043 532 1044 533
rect 1094 532 1095 533
rect 1122 532 1123 533
rect 1173 532 1174 533
rect 1201 532 1202 533
rect 886 503 904 532
rect 935 531 966 532
rect 1014 531 1045 532
rect 1093 531 1124 532
rect 1172 531 1203 532
rect 936 524 965 531
rect 1015 524 1044 531
rect 1094 524 1123 531
rect 1173 524 1202 531
rect 936 510 946 524
rect 1193 510 1202 524
rect 936 504 965 510
rect 1015 504 1044 510
rect 1094 504 1123 510
rect 1173 504 1202 510
rect 935 503 966 504
rect 1014 503 1045 504
rect 1093 503 1124 504
rect 1172 503 1203 504
rect 1235 503 1252 532
rect 936 502 937 503
rect 964 502 965 503
rect 1015 502 1016 503
rect 1043 502 1044 503
rect 1094 502 1095 503
rect 1122 502 1123 503
rect 1173 502 1174 503
rect 1201 502 1202 503
rect 936 453 965 468
rect 1015 453 1044 468
rect 1094 453 1123 468
rect 1173 453 1202 468
rect 936 286 965 302
rect 1015 286 1044 302
rect 1094 286 1123 302
rect 1173 286 1202 302
rect 936 252 937 253
rect 964 252 965 253
rect 1015 252 1016 253
rect 1043 252 1044 253
rect 1094 252 1095 253
rect 1122 252 1123 253
rect 1173 252 1174 253
rect 1201 252 1202 253
rect 886 223 904 252
rect 935 251 966 252
rect 1014 251 1045 252
rect 1093 251 1124 252
rect 1172 251 1203 252
rect 936 244 965 251
rect 1015 244 1044 251
rect 1094 244 1123 251
rect 1173 244 1202 251
rect 936 230 946 244
rect 1193 230 1202 244
rect 936 224 965 230
rect 1015 224 1044 230
rect 1094 224 1123 230
rect 1173 224 1202 230
rect 935 223 966 224
rect 1014 223 1045 224
rect 1093 223 1124 224
rect 1172 223 1203 224
rect 1235 223 1252 252
rect 936 222 937 223
rect 964 222 965 223
rect 1015 222 1016 223
rect 1043 222 1044 223
rect 1094 222 1095 223
rect 1122 222 1123 223
rect 1173 222 1174 223
rect 1201 222 1202 223
rect 77 204 106 222
rect 936 173 965 188
rect 1015 173 1044 188
rect 1094 173 1123 188
rect 1173 173 1202 188
rect 77 172 78 173
rect 105 172 106 173
rect 27 143 45 172
rect 76 171 107 172
rect 77 162 106 171
rect 77 153 87 162
rect 96 153 106 162
rect 77 144 106 153
rect 76 143 107 144
rect 138 143 156 172
rect 77 142 78 143
rect 105 142 106 143
rect 936 131 965 147
rect 1015 131 1044 147
rect 1094 131 1123 147
rect 1173 131 1202 147
rect 77 93 106 111
rect 936 97 937 98
rect 964 97 965 98
rect 1015 97 1016 98
rect 1043 97 1044 98
rect 1094 97 1095 98
rect 1122 97 1123 98
rect 1173 97 1174 98
rect 1201 97 1202 98
rect 886 68 904 97
rect 935 96 966 97
rect 1014 96 1045 97
rect 1093 96 1124 97
rect 1172 96 1203 97
rect 936 89 965 96
rect 1015 89 1044 96
rect 1094 89 1123 96
rect 1173 89 1202 96
rect 936 75 946 89
rect 1193 75 1202 89
rect 936 69 965 75
rect 1015 69 1044 75
rect 1094 69 1123 75
rect 1173 69 1202 75
rect 935 68 966 69
rect 1014 68 1045 69
rect 1093 68 1124 69
rect 1172 68 1203 69
rect 1235 68 1252 97
rect 936 67 937 68
rect 964 67 965 68
rect 1015 67 1016 68
rect 1043 67 1044 68
rect 1094 67 1095 68
rect 1122 67 1123 68
rect 1173 67 1174 68
rect 1201 67 1202 68
rect 936 18 965 33
rect 1015 18 1044 33
rect 1094 18 1123 33
rect 1173 18 1202 33
<< nwell >>
rect 888 438 1003 455
rect 1007 438 1058 455
rect 869 320 1269 438
rect 869 319 1058 320
rect 1190 319 1269 320
rect 888 300 1003 319
rect 1007 299 1058 319
rect 1163 300 1190 318
rect 2683 250 2957 600
rect 475 168 497 179
<< mvnmos >>
rect 2572 505 2635 555
rect 2572 283 2635 333
rect 2572 116 2634 193
rect 2717 116 2781 171
rect 2859 116 2923 171
<< mvpmos >>
rect 2720 479 2780 534
rect 2860 479 2920 534
rect 2720 312 2780 367
rect 2860 312 2920 367
<< mvndiff >>
rect 2572 578 2635 582
rect 2572 561 2578 578
rect 2595 561 2612 578
rect 2629 561 2635 578
rect 2572 555 2635 561
rect 2572 492 2635 505
rect 2572 333 2635 338
rect 2572 277 2635 283
rect 2572 260 2577 277
rect 2594 260 2611 277
rect 2628 260 2635 277
rect 2572 254 2635 260
rect 2572 216 2634 224
rect 2572 199 2577 216
rect 2594 199 2611 216
rect 2628 199 2634 216
rect 2572 193 2634 199
rect 2717 194 2781 201
rect 2717 177 2724 194
rect 2741 177 2758 194
rect 2775 177 2781 194
rect 2717 171 2781 177
rect 2859 194 2923 200
rect 2859 177 2865 194
rect 2882 177 2899 194
rect 2916 177 2923 194
rect 2859 171 2923 177
rect 2572 110 2634 116
rect 2572 93 2576 110
rect 2593 93 2610 110
rect 2627 93 2634 110
rect 2572 86 2634 93
rect 2717 110 2781 116
rect 2717 93 2724 110
rect 2741 93 2758 110
rect 2775 93 2781 110
rect 2717 86 2781 93
rect 2859 110 2923 116
rect 2859 93 2865 110
rect 2882 93 2899 110
rect 2916 93 2923 110
rect 2859 87 2923 93
<< mvpdiff >>
rect 2720 557 2780 563
rect 2720 540 2724 557
rect 2741 540 2758 557
rect 2775 540 2780 557
rect 2720 534 2780 540
rect 2860 557 2920 563
rect 2860 540 2865 557
rect 2882 540 2899 557
rect 2916 540 2920 557
rect 2860 534 2920 540
rect 2720 472 2780 479
rect 2720 455 2724 472
rect 2741 455 2758 472
rect 2775 455 2780 472
rect 2720 438 2780 455
rect 2720 390 2780 408
rect 2720 373 2724 390
rect 2741 373 2758 390
rect 2775 373 2780 390
rect 2720 367 2780 373
rect 2860 472 2920 479
rect 2860 455 2865 472
rect 2882 455 2899 472
rect 2916 455 2920 472
rect 2860 438 2920 455
rect 2860 390 2920 408
rect 2860 373 2865 390
rect 2882 373 2899 390
rect 2916 373 2920 390
rect 2860 367 2920 373
rect 2720 306 2780 312
rect 2720 289 2724 306
rect 2741 289 2758 306
rect 2775 289 2780 306
rect 2720 283 2780 289
rect 2860 306 2920 312
rect 2860 289 2865 306
rect 2882 289 2899 306
rect 2916 289 2920 306
rect 2860 283 2920 289
<< mvndiffc >>
rect 2578 561 2595 578
rect 2612 561 2629 578
rect 2577 260 2594 277
rect 2611 260 2628 277
rect 2577 199 2594 216
rect 2611 199 2628 216
rect 2724 177 2741 194
rect 2758 177 2775 194
rect 2865 177 2882 194
rect 2899 177 2916 194
rect 2576 93 2593 110
rect 2610 93 2627 110
rect 2724 93 2741 110
rect 2758 93 2775 110
rect 2865 93 2882 110
rect 2899 93 2916 110
<< mvpdiffc >>
rect 2724 540 2741 557
rect 2758 540 2775 557
rect 2865 540 2882 557
rect 2899 540 2916 557
rect 2724 455 2741 472
rect 2758 455 2775 472
rect 2724 373 2741 390
rect 2758 373 2775 390
rect 2865 455 2882 472
rect 2899 455 2916 472
rect 2865 373 2882 390
rect 2899 373 2916 390
rect 2724 289 2741 306
rect 2758 289 2775 306
rect 2865 289 2882 306
rect 2899 289 2916 306
<< psubdiff >>
rect 351 378 685 383
rect 351 361 391 378
rect 408 361 425 378
rect 442 361 459 378
rect 476 361 493 378
rect 510 361 527 378
rect 544 361 561 378
rect 578 361 595 378
rect 612 361 629 378
rect 646 361 685 378
rect 351 357 685 361
rect 351 338 380 357
rect 351 321 357 338
rect 374 321 380 338
rect 351 309 380 321
rect 235 304 380 309
rect 235 296 357 304
rect 235 279 255 296
rect 272 279 289 296
rect 306 279 323 296
rect 340 287 357 296
rect 374 287 380 304
rect 340 279 380 287
rect 235 271 380 279
rect 351 270 380 271
rect 351 253 357 270
rect 374 253 380 270
rect 351 236 380 253
rect 351 219 357 236
rect 374 219 380 236
rect 351 202 380 219
rect 351 185 357 202
rect 374 185 380 202
rect 351 168 380 185
rect 1332 344 1371 377
rect 1332 327 1344 344
rect 1361 327 1371 344
rect 1332 298 1371 327
rect 1332 281 1344 298
rect 1361 281 1371 298
rect 1332 260 1371 281
rect 1332 243 1344 260
rect 1361 243 1371 260
rect 1332 217 1371 243
rect 1332 200 1344 217
rect 1361 200 1371 217
rect 351 151 357 168
rect 374 151 380 168
rect 351 134 380 151
rect 351 117 357 134
rect 374 117 380 134
rect 351 100 380 117
rect 351 83 357 100
rect 374 83 380 100
rect 1332 162 1371 200
rect 1332 145 1344 162
rect 1361 145 1371 162
rect 1332 122 1371 145
rect 1332 105 1344 122
rect 1361 105 1371 122
rect 351 71 380 83
rect 1332 86 1371 105
rect 1332 69 1344 86
rect 1361 69 1371 86
rect 1332 48 1371 69
rect 1332 31 1343 48
rect 1360 31 1371 48
rect 1332 15 1371 31
<< mvpsubdiff >>
rect 2573 43 2927 49
rect 2573 42 2653 43
rect 2573 25 2585 42
rect 2602 25 2619 42
rect 2636 26 2653 42
rect 2670 26 2689 43
rect 2706 26 2725 43
rect 2742 26 2759 43
rect 2776 26 2793 43
rect 2810 26 2827 43
rect 2844 26 2861 43
rect 2878 26 2895 43
rect 2912 26 2927 43
rect 2636 25 2927 26
rect 2573 19 2927 25
<< mvnsubdiff >>
rect 1195 429 1236 437
rect 1195 416 1207 429
rect 1181 412 1207 416
rect 1224 412 1236 429
rect 1181 395 1236 412
rect 1181 378 1207 395
rect 1224 378 1236 395
rect 1181 377 1236 378
rect 1195 361 1236 377
rect 1195 344 1207 361
rect 1224 344 1236 361
rect 1195 339 1236 344
rect 1196 335 1236 339
rect 2720 431 2780 438
rect 2720 414 2741 431
rect 2758 414 2780 431
rect 2720 408 2780 414
rect 2860 431 2920 438
rect 2860 414 2881 431
rect 2898 414 2920 431
rect 2860 408 2920 414
rect 475 168 497 179
<< psubdiffcont >>
rect 391 361 408 378
rect 425 361 442 378
rect 459 361 476 378
rect 493 361 510 378
rect 527 361 544 378
rect 561 361 578 378
rect 595 361 612 378
rect 629 361 646 378
rect 357 321 374 338
rect 255 279 272 296
rect 289 279 306 296
rect 323 279 340 296
rect 357 287 374 304
rect 357 253 374 270
rect 357 219 374 236
rect 357 185 374 202
rect 1344 327 1361 344
rect 1344 281 1361 298
rect 1344 243 1361 260
rect 1344 200 1361 217
rect 357 151 374 168
rect 357 117 374 134
rect 357 83 374 100
rect 1344 145 1361 162
rect 1344 105 1361 122
rect 1344 69 1361 86
rect 1343 31 1360 48
<< mvpsubdiffcont >>
rect 2585 25 2602 42
rect 2619 25 2636 42
rect 2653 26 2670 43
rect 2689 26 2706 43
rect 2725 26 2742 43
rect 2759 26 2776 43
rect 2793 26 2810 43
rect 2827 26 2844 43
rect 2861 26 2878 43
rect 2895 26 2912 43
<< mvnsubdiffcont >>
rect 1207 412 1224 429
rect 1207 378 1224 395
rect 1207 344 1224 361
rect 2741 414 2758 431
rect 2881 414 2898 431
<< poly >>
rect 176 487 204 537
rect 179 420 204 487
rect 698 457 747 544
rect 2361 542 2572 555
rect 698 455 892 457
rect 1175 455 1226 456
rect 1249 455 1445 542
rect 2360 505 2572 542
rect 2635 505 2648 555
rect 2796 556 2804 572
rect 2796 534 2816 556
rect 2937 555 2946 572
rect 2934 534 2952 555
rect 2360 491 2414 505
rect 2706 479 2720 534
rect 2780 479 2816 534
rect 2844 479 2860 534
rect 2920 479 2952 534
rect 698 420 1044 455
rect 67 396 1044 420
rect 67 217 105 396
rect 698 300 1044 396
rect 2618 399 2665 433
rect 2649 333 2665 399
rect 2796 367 2816 479
rect 2935 367 2952 479
rect 1175 318 1226 319
rect 1163 300 1226 318
rect 698 299 892 300
rect 993 299 1044 300
rect 698 174 747 299
rect 2557 283 2572 333
rect 2635 283 2665 333
rect 2706 312 2720 367
rect 2780 312 2816 367
rect 2846 312 2860 367
rect 2920 312 2952 367
rect 2660 236 2698 237
rect 698 145 987 174
rect 2642 198 2698 236
rect 2642 193 2663 198
rect 698 90 747 145
rect 2557 116 2572 193
rect 2634 178 2663 193
rect 2634 116 2648 178
rect 2701 116 2717 171
rect 2781 116 2859 171
rect 2923 116 2936 171
<< locali >>
rect 2570 561 2578 578
rect 2629 561 2637 578
rect 2800 557 2808 572
rect 2937 558 2946 572
rect 2857 557 2957 558
rect 2716 540 2724 557
rect 2775 540 2817 557
rect 2857 540 2865 557
rect 2916 540 2957 557
rect 2716 455 2724 472
rect 2775 455 2865 472
rect 2916 455 2924 472
rect 1207 429 1224 437
rect 2724 414 2741 431
rect 2775 414 2864 431
rect 2898 414 2906 431
rect 1207 402 1224 412
rect 1207 395 1267 402
rect 357 378 374 380
rect 1224 378 1267 395
rect 357 361 391 378
rect 408 361 425 378
rect 442 361 459 378
rect 476 361 493 378
rect 510 361 527 378
rect 544 361 561 378
rect 578 361 595 378
rect 612 361 629 378
rect 646 361 663 378
rect 1207 376 1267 378
rect 1207 361 1224 376
rect 2716 373 2724 390
rect 2775 373 2865 390
rect 2916 373 2924 390
rect 357 338 374 361
rect 1207 336 1224 344
rect 1344 344 1361 355
rect 357 304 374 321
rect 247 279 255 296
rect 272 279 289 296
rect 306 279 323 296
rect 340 287 357 296
rect 340 279 374 287
rect 357 270 374 279
rect 357 236 374 253
rect 357 202 374 219
rect 357 168 374 185
rect 357 134 374 151
rect 357 100 374 117
rect 1344 298 1361 327
rect 2716 289 2724 306
rect 2775 289 2784 306
rect 2857 289 2865 306
rect 2916 289 2924 306
rect 1344 260 1361 281
rect 2569 260 2577 277
rect 2594 260 2611 277
rect 2628 260 2683 277
rect 1344 217 1361 243
rect 1344 162 1361 200
rect 2569 199 2577 216
rect 2628 199 2636 216
rect 2716 177 2724 194
rect 2775 177 2804 194
rect 2857 177 2865 194
rect 2916 177 2924 194
rect 1344 122 1361 145
rect 1344 90 1361 105
rect 2567 93 2576 110
rect 2593 93 2610 110
rect 2627 93 2724 110
rect 2741 93 2758 110
rect 2775 93 2865 110
rect 2882 93 2899 110
rect 2916 93 2925 110
rect 357 38 374 83
rect 1343 86 1361 90
rect 1343 69 1344 86
rect 1343 48 1361 69
rect 1360 31 1361 48
rect 2594 43 2662 48
rect 2594 42 2653 43
rect 1343 17 1361 31
rect 2577 25 2585 42
rect 2602 25 2619 42
rect 2636 26 2653 42
rect 2670 26 2689 43
rect 2706 26 2725 43
rect 2742 26 2759 43
rect 2776 26 2793 43
rect 2810 26 2827 43
rect 2844 26 2861 43
rect 2878 26 2895 43
rect 2912 26 2920 43
rect 2636 25 2662 26
<< viali >>
rect 2595 561 2612 578
rect 2741 540 2758 557
rect 2882 540 2899 557
rect 2741 455 2758 472
rect 2882 455 2899 472
rect 2758 414 2775 431
rect 2864 414 2881 431
rect 2741 373 2758 390
rect 2882 373 2899 390
rect 2741 289 2758 306
rect 2882 289 2899 306
rect 2594 199 2611 216
rect 2741 177 2758 194
rect 2882 177 2899 194
<< metal1 >>
rect 0 516 26 605
rect 470 480 497 605
rect 1057 564 1081 605
rect 2589 578 2618 581
rect 2589 561 2595 578
rect 2612 561 2618 578
rect 2589 558 2618 561
rect 2665 557 2768 565
rect 2665 540 2741 557
rect 2758 540 2768 557
rect 2665 534 2768 540
rect 2871 557 2909 565
rect 2871 540 2882 557
rect 2899 540 2909 557
rect 2871 534 2909 540
rect 2590 489 2617 502
rect 2581 480 2617 489
rect 2581 460 2623 480
rect 2581 366 2604 460
rect 2581 348 2617 366
rect 79 18 104 205
rect 78 0 104 18
rect 469 0 500 259
rect 2590 219 2617 348
rect 2665 257 2689 534
rect 2738 472 2761 478
rect 2738 455 2741 472
rect 2758 455 2761 472
rect 2878 472 2902 478
rect 2878 455 2882 472
rect 2899 455 2902 472
rect 2733 431 2908 455
rect 2733 414 2758 431
rect 2775 414 2864 431
rect 2881 414 2908 431
rect 2733 390 2908 414
rect 2733 389 2741 390
rect 2738 373 2741 389
rect 2758 389 2882 390
rect 2758 373 2761 389
rect 2738 367 2761 373
rect 2878 373 2882 389
rect 2899 389 2908 390
rect 2899 373 2902 389
rect 2878 367 2902 373
rect 2738 306 2761 312
rect 2738 289 2741 306
rect 2758 289 2761 306
rect 2584 216 2617 219
rect 2584 199 2594 216
rect 2611 199 2617 216
rect 2584 196 2617 199
rect 2738 194 2761 289
rect 1058 0 1082 188
rect 2738 177 2741 194
rect 2758 177 2761 194
rect 2738 171 2761 177
rect 2879 306 2902 312
rect 2879 289 2882 306
rect 2899 289 2902 306
rect 2879 194 2902 289
rect 2879 177 2882 194
rect 2899 177 2902 194
rect 2879 171 2902 177
rect 2389 0 2418 106
<< metal2 >>
rect 2588 558 2877 582
rect 1235 459 2700 472
rect 1235 451 2967 459
rect 1058 381 1088 427
rect 1131 382 1161 428
rect 1269 384 1293 451
rect 2686 434 2967 451
rect 2622 300 2649 428
rect 2700 383 2967 434
rect 2622 299 2901 300
rect 2622 277 2967 299
rect 2674 276 2967 277
rect 2905 228 2967 260
rect 2664 189 2967 212
rect 2579 62 2967 95
rect 2578 53 2967 62
rect 2579 46 2967 53
rect 2603 28 2647 46
rect 353 7 2676 28
use sky130_hilas_li2m2  sky130_hilas_li2m2_13
timestamp 1628616688
transform 1 0 1073 0 1 395
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_14
timestamp 1628616688
transform 1 0 364 0 1 24
box 0 0 34 33
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_0
timestamp 1628616694
transform 1 0 89 0 1 136
box 0 0 129 129
use sky130_hilas_pFETdevice01w1  sky130_hilas_pFETdevice01w1_0
timestamp 1628616668
transform 1 0 1108 0 1 396
box 0 0 161 121
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628616688
transform 1 0 1350 0 1 22
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_12
timestamp 1628616688
transform 1 0 1142 0 1 396
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_11
timestamp 1628616688
transform 1 0 1278 0 1 388
box 0 0 34 33
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_0
timestamp 1628616755
transform 1 0 1447 0 1 414
box 0 0 272 169
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_2
timestamp 1628616755
transform 1 0 1447 0 1 515
box 0 0 272 169
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_1
timestamp 1628616674
transform 1 0 1390 0 1 209
box 0 0 400 164
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_2
timestamp 1628616674
transform 1 0 1390 0 1 54
box 0 0 400 164
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_0
timestamp 1628616674
transform 1 0 1390 0 1 489
box 0 0 400 164
use sky130_hilas_li2m2  sky130_hilas_li2m2_9
timestamp 1628616688
transform 1 0 2590 0 1 39
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_4
timestamp 1628616688
transform 1 0 2676 0 1 100
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_5
timestamp 1628616688
transform 1 0 2661 0 1 40
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_6
timestamp 1628616688
transform 1 0 2735 0 1 40
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1628616688
transform 1 0 2819 0 1 98
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_7
timestamp 1628616688
transform 1 0 2805 0 1 40
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_8
timestamp 1628616688
transform 1 0 2898 0 1 40
box 0 0 34 33
use sky130_hilas_nDiffThOxContact  sky130_hilas_nDiffThOxContact_3
timestamp 1628616954
transform 1 0 2596 0 1 321
box 0 0 67 29
use sky130_hilas_poly2li  sky130_hilas_poly2li_5
timestamp 1628616704
transform -1 0 2689 0 -1 221
box 0 0 27 33
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1628616665
transform 1 0 2675 0 1 265
box 0 0 23 29
use sky130_hilas_li2m2  sky130_hilas_li2m2_10
timestamp 1628616688
transform -1 0 2679 0 -1 220
box 0 0 34 33
use sky130_hilas_poly2li  sky130_hilas_poly2li_3
timestamp 1628616704
transform 1 0 2805 0 1 181
box 0 0 27 33
use sky130_hilas_m12m2  sky130_hilas_m12m2_9
timestamp 1628616702
transform 1 0 2884 0 1 238
box 0 0 32 32
use sky130_hilas_nDiffThOxContact  sky130_hilas_nDiffThOxContact_0
timestamp 1628616954
transform 1 0 2596 0 1 464
box 0 0 67 29
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_0
timestamp 1628616734
transform 1 0 2627 0 1 407
box 0 0 33 55
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1628616702
transform 1 0 2743 0 1 417
box 0 0 32 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_4
timestamp 1628616702
transform 1 0 2741 0 1 375
box 0 0 32 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_6
timestamp 1628616702
transform 1 0 2743 0 1 461
box 0 0 32 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1628616702
transform 1 0 2884 0 1 415
box 0 0 32 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_2
timestamp 1628616702
transform 1 0 2884 0 1 460
box 0 0 32 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_3
timestamp 1628616702
transform 1 0 2884 0 1 373
box 0 0 32 32
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628616688
transform 1 0 2817 0 1 378
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1628616688
transform 1 0 2817 0 1 462
box 0 0 34 33
use sky130_hilas_m12m2  sky130_hilas_m12m2_10
timestamp 1628616702
transform 1 0 2597 0 1 568
box 0 0 32 32
use sky130_hilas_poly2li  sky130_hilas_poly2li_1
timestamp 1628616704
transform 1 0 2808 0 1 569
box 0 0 27 33
use sky130_hilas_m12m2  sky130_hilas_m12m2_7
timestamp 1628616702
transform 1 0 2883 0 1 563
box 0 0 32 32
use sky130_hilas_poly2li  sky130_hilas_poly2li_4
timestamp 1628616704
transform 1 0 2948 0 1 569
box 0 0 27 33
use sky130_hilas_FGVaractorTunnelCap01  sky130_hilas_FGVaractorTunnelCap01_0
timestamp 1628616690
transform 1 0 977 0 1 809
box 0 0 222 169
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_1
timestamp 1628616755
transform 1 0 1447 0 1 814
box 0 0 272 169
use sky130_hilas_FGHugeVaractorCapacitor01  sky130_hilas_FGHugeVaractorCapacitor01_0
timestamp 1628616676
transform 1 0 1983 0 1 818
box 0 0 1029 599
<< labels >>
rlabel metal2 2961 46 2967 95 0 VGND
port 8 nsew ground default
rlabel metal2 2961 228 2967 260 0 OUTPUT
port 10 nsew analog default
rlabel metal2 2960 383 2967 459 0 VINJ
port 9 nsew power default
rlabel metal2 2961 189 2967 212 0 VBIAS
port 12 nsew analog default
rlabel metal2 2961 276 2967 299 0 VREF
port 11 nsew analog default
rlabel metal1 2389 2 2418 7 0 LARGECAPACITOR
port 7 nsew analog default
rlabel metal1 1057 599 1081 605 0 GATE3
port 3 nsew analog default
rlabel metal1 1058 0 1082 7 0 GATE4
port 6 nsew analog default
rlabel metal1 469 0 500 7 0 GATE2
port 5 nsew analog default
rlabel metal1 470 596 497 605 0 GATE1
port 2 nsew analog default
rlabel metal1 78 0 104 10 0 VTUNOVERLAP01
port 4 nsew analog default
rlabel metal1 0 598 26 605 0 VTUN
port 1 nsew analog default
rlabel metal2 1058 416 1088 427 0 DRAIN1
port 13 nsew
rlabel metal2 1131 417 1160 428 0 SOURCE1
port 14 nsew
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
