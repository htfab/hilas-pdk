magic
tech sky130A
magscale 1 2
timestamp 1632256331
<< checkpaint >>
rect -810 2666 1976 2758
rect -1212 -1156 1976 2666
rect -810 -1254 1976 -1156
<< error_s >>
rect 650 1494 662 1504
rect 616 1452 628 1486
rect 650 1460 716 1494
rect 616 1436 634 1452
rect 168 1356 228 1370
rect 268 1356 334 1370
rect 168 1348 218 1356
rect 228 1348 248 1354
rect 156 1346 248 1348
rect 268 1346 272 1348
rect 156 1344 272 1346
rect 156 1320 248 1344
rect 268 1320 272 1344
rect 194 1318 214 1320
rect 228 1318 268 1320
rect 280 1318 314 1356
rect 346 1320 386 1334
rect 450 1320 464 1424
rect 492 1362 578 1364
rect 480 1328 544 1330
rect 168 1286 218 1318
rect 228 1288 248 1318
rect 334 1292 396 1320
rect 280 1286 396 1292
rect 168 1268 228 1286
rect 268 1278 384 1286
rect 268 1268 416 1278
rect 280 1260 416 1268
rect 284 1250 322 1252
rect 324 1250 416 1260
rect 108 1242 226 1244
rect 280 1238 314 1250
rect 334 1248 416 1250
rect 280 1224 334 1238
rect 136 1214 198 1216
rect 104 1198 136 1214
rect 218 1212 280 1224
rect 138 1198 170 1208
rect 104 1166 170 1198
rect 194 1200 202 1208
rect 194 1166 204 1200
rect 218 1187 238 1212
rect 228 1170 238 1187
rect 250 1170 268 1212
rect 272 1209 280 1212
rect 284 1184 302 1224
rect 334 1223 396 1224
rect 346 1186 386 1202
rect 450 1186 464 1292
rect 480 1284 546 1308
rect 480 1278 544 1284
rect 492 1250 580 1274
rect 492 1244 578 1250
rect 334 1176 396 1186
rect 280 1170 396 1176
rect 218 1166 396 1170
rect 104 1156 396 1166
rect 104 1150 142 1156
rect 168 1154 396 1156
rect 104 1148 136 1150
rect 108 1128 114 1148
rect 168 1144 384 1154
rect 156 1136 384 1144
rect 156 1134 358 1136
rect 156 1116 359 1134
rect 218 1114 334 1116
rect 168 1064 322 1114
rect 218 1046 272 1050
rect 168 1024 322 1046
rect 360 1044 398 1050
rect 360 1026 362 1044
rect 360 1024 398 1026
rect 156 1004 398 1024
rect 156 996 364 1004
rect 164 994 334 996
rect 108 962 114 982
rect 168 970 322 994
rect 334 992 359 994
rect 326 970 394 992
rect 104 960 136 962
rect 104 954 142 960
rect 168 956 392 970
rect 168 954 218 956
rect 104 944 218 954
rect 104 912 170 944
rect 104 896 136 912
rect 138 902 170 912
rect 194 910 204 944
rect 228 923 238 954
rect 194 902 202 910
rect 218 908 238 923
rect 250 908 268 954
rect 280 934 396 956
rect 284 916 302 926
rect 334 924 396 934
rect 218 901 272 908
rect 280 901 396 916
rect 218 886 396 901
rect 238 878 272 886
rect 280 862 334 886
rect 280 861 396 862
rect 280 860 345 861
rect 284 858 322 860
rect 168 824 228 842
rect 268 824 322 842
rect 324 840 356 860
rect 324 824 392 840
rect 168 820 218 824
rect 228 820 248 822
rect 156 792 248 820
rect 268 792 272 820
rect 194 790 214 792
rect 228 790 268 792
rect 280 790 314 824
rect 334 790 396 824
rect 168 774 218 790
rect 146 766 218 774
rect 228 788 248 790
rect 228 766 268 788
rect 146 764 272 766
rect 168 748 218 764
rect 228 756 268 764
rect 228 748 268 754
rect 156 746 272 748
rect 146 736 272 746
rect 156 722 272 736
rect 156 720 248 722
rect 268 720 272 722
rect 194 718 214 720
rect 228 718 268 720
rect 280 718 314 762
rect 346 756 386 788
rect 346 720 386 754
rect 168 686 218 718
rect 228 688 248 718
rect 334 692 396 720
rect 280 686 396 692
rect 168 668 228 686
rect 268 678 384 686
rect 268 668 416 678
rect 280 660 416 668
rect 284 650 322 652
rect 324 650 416 660
rect 280 638 314 650
rect 334 648 416 650
rect 280 624 334 638
rect 104 598 136 614
rect 218 612 280 624
rect 138 598 170 608
rect 104 566 170 598
rect 194 600 202 608
rect 194 566 204 600
rect 218 587 238 612
rect 228 570 238 587
rect 250 570 268 612
rect 272 609 280 612
rect 284 584 302 624
rect 334 623 396 624
rect 382 602 396 623
rect 346 586 396 602
rect 334 576 396 586
rect 280 570 396 576
rect 218 566 396 570
rect 104 556 396 566
rect 104 550 142 556
rect 168 554 396 556
rect 104 548 136 550
rect 108 528 114 548
rect 168 544 384 554
rect 156 536 384 544
rect 156 534 358 536
rect 156 516 359 534
rect 218 514 334 516
rect 168 464 322 514
rect 218 446 272 450
rect 168 424 322 446
rect 156 396 364 424
rect 164 394 334 396
rect 108 362 114 382
rect 168 370 322 394
rect 334 376 359 394
rect 334 374 358 376
rect 334 372 384 374
rect 334 370 392 372
rect 104 360 136 362
rect 104 354 142 360
rect 168 356 392 370
rect 168 354 218 356
rect 104 344 218 354
rect 104 312 170 344
rect 104 296 136 312
rect 138 302 170 312
rect 194 310 204 344
rect 228 323 238 354
rect 194 302 202 310
rect 218 308 238 323
rect 250 308 268 354
rect 280 334 396 356
rect 284 316 302 326
rect 334 324 396 334
rect 218 301 272 308
rect 280 301 396 316
rect 218 286 396 301
rect 450 286 464 324
rect 238 278 272 286
rect 280 262 334 286
rect 280 261 396 262
rect 280 260 345 261
rect 284 258 322 260
rect 168 224 228 242
rect 268 238 322 242
rect 324 240 356 260
rect 324 238 392 240
rect 268 224 392 238
rect 168 220 218 224
rect 228 220 248 222
rect 156 192 248 220
rect 268 192 272 220
rect 194 190 214 192
rect 228 190 268 192
rect 280 190 314 224
rect 334 190 396 224
rect 168 166 218 190
rect 228 166 248 190
rect 168 164 272 166
rect 168 154 218 164
rect 228 156 248 164
rect 450 154 464 190
rect 168 140 228 154
rect 268 140 334 154
rect 616 52 634 68
rect 644 52 678 86
rect 616 18 628 52
rect 650 18 666 34
rect 650 0 662 18
<< metal1 >>
rect 192 184 260 1328
rect 326 186 380 1326
<< metal2 >>
rect 2 1242 510 1288
rect 54 814 584 860
rect 2 650 584 694
rect 0 216 542 262
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1632251332
transform 1 0 356 0 1 480
box 0 0 46 58
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1632251356
transform 1 0 470 0 1 234
box 0 0 68 66
use sky130_hilas_pFETmirror02  sky130_hilas_pFETmirror02_0
timestamp 1632256314
transform 1 0 450 0 1 6
box 0 0 266 584
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_0
timestamp 1632256312
transform 1 0 48 0 -1 422
box 0 0 368 318
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_1
timestamp 1632256312
transform 1 0 48 0 1 488
box 0 0 368 318
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1632251332
transform 1 0 356 0 1 998
box 0 0 46 58
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1632251356
transform 1 0 488 0 1 828
box 0 0 68 66
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1632251356
transform 1 0 486 0 1 684
box 0 0 68 66
use sky130_hilas_pFETmirror02  sky130_hilas_pFETmirror02_1
timestamp 1632256314
transform 1 0 450 0 -1 1498
box 0 0 266 584
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_2
timestamp 1632256312
transform 1 0 48 0 1 1088
box 0 0 368 318
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_3
timestamp 1632256312
transform 1 0 48 0 -1 1022
box 0 0 368 318
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1632251356
transform 1 0 478 0 1 1272
box 0 0 68 66
<< labels >>
rlabel metal2 562 814 584 860 0 output1
rlabel space 562 650 584 696 0 output2
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
