VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_hilas_TA2Cell_1FG_Strong
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TA2Cell_1FG_Strong ;
  ORIGIN 26.170 -1.350 ;
  SIZE 28.100 BY 6.150 ;
  PIN VTUN
    ANTENNADIFFAREA 5.032200 ;
    PORT
      LAYER nwell ;
        RECT -16.380 6.700 -12.990 7.450 ;
        RECT -16.390 3.130 -12.980 6.700 ;
        RECT -16.380 1.410 -12.990 3.130 ;
      LAYER met1 ;
        RECT -15.410 7.300 -14.990 7.450 ;
        RECT -14.380 7.300 -13.960 7.450 ;
        RECT -15.410 7.160 -13.960 7.300 ;
        RECT -15.410 1.400 -14.990 7.160 ;
        RECT -14.380 1.400 -13.960 7.160 ;
    END
  END VTUN
  PIN PROG
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER met1 ;
        RECT -22.650 4.730 -22.440 7.450 ;
        RECT -22.680 4.220 -22.440 4.730 ;
        RECT -22.650 1.400 -22.440 4.220 ;
    END
  END PROG
  PIN GATE1
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT -10.960 5.060 -8.240 6.710 ;
        RECT -10.960 5.020 -8.250 5.060 ;
        RECT -10.960 3.690 -8.250 3.730 ;
        RECT -10.960 2.040 -8.240 3.690 ;
      LAYER met1 ;
        RECT -10.680 6.240 -10.450 7.450 ;
        RECT -10.680 5.450 -10.420 6.240 ;
        RECT -10.680 3.300 -10.450 5.450 ;
        RECT -10.680 2.510 -10.420 3.300 ;
        RECT -10.680 1.400 -10.450 2.510 ;
    END
  END GATE1
  PIN VIN11
    ANTENNADIFFAREA 0.217200 ;
    PORT
      LAYER met1 ;
        RECT -23.530 7.080 -23.320 7.450 ;
        RECT -23.540 6.790 -23.310 7.080 ;
        RECT -23.530 5.090 -23.320 6.790 ;
        RECT -23.540 4.800 -23.310 5.090 ;
        RECT -23.530 4.660 -23.320 4.800 ;
    END
  END VIN11
  PIN VINJ
    ANTENNADIFFAREA 2.118400 ;
    PORT
      LAYER nwell ;
        RECT -26.170 1.350 -22.860 7.500 ;
        RECT -6.510 7.450 -3.200 7.500 ;
        RECT -6.510 7.440 -1.860 7.450 ;
        RECT -6.510 1.400 -1.350 7.440 ;
        RECT -6.510 1.350 -3.200 1.400 ;
      LAYER met2 ;
        RECT -25.970 7.310 -25.650 7.430 ;
        RECT -3.700 7.310 -3.380 7.430 ;
        RECT -25.970 7.130 -3.380 7.310 ;
        RECT -4.590 4.590 -4.270 4.850 ;
        RECT -4.550 4.570 -3.370 4.590 ;
        RECT -4.550 4.310 -3.330 4.570 ;
        RECT -4.550 4.250 -3.370 4.310 ;
        RECT -4.590 4.240 -3.370 4.250 ;
        RECT -4.590 3.990 -4.270 4.240 ;
    END
    PORT
      LAYER met1 ;
        RECT -3.720 7.430 -3.440 7.450 ;
        RECT -3.720 7.130 -3.380 7.430 ;
        RECT -3.720 6.800 -3.440 7.130 ;
        RECT -3.830 6.200 -3.440 6.800 ;
        RECT -3.720 4.600 -3.440 6.200 ;
        RECT -3.720 4.280 -3.360 4.600 ;
        RECT -3.720 2.650 -3.440 4.280 ;
        RECT -3.830 2.050 -3.440 2.650 ;
        RECT -3.720 1.400 -3.440 2.050 ;
      LAYER via ;
        RECT -3.670 7.150 -3.410 7.410 ;
        RECT -3.620 4.310 -3.360 4.570 ;
    END
  END VINJ
  PIN VIN22
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -1.960 7.430 -1.650 7.440 ;
        RECT -2.530 7.420 -1.650 7.430 ;
        RECT -2.600 7.180 -1.650 7.420 ;
        RECT -1.960 7.110 -1.650 7.180 ;
    END
  END VIN22
  PIN VIN21
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -2.200 4.750 -1.890 4.790 ;
        RECT -2.520 4.740 -1.860 4.750 ;
        RECT -2.520 4.510 -1.420 4.740 ;
        RECT -2.200 4.460 -1.890 4.510 ;
    END
  END VIN21
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.650 1.400 1.930 7.450 ;
      LAYER met1 ;
        RECT 0.630 7.300 0.910 7.450 ;
        RECT 0.640 5.870 0.910 7.300 ;
        RECT 0.640 5.580 0.920 5.870 ;
        RECT 0.640 3.280 0.910 5.580 ;
        RECT 0.640 2.990 0.920 3.280 ;
        RECT 0.640 1.400 0.910 2.990 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT -1.560 1.750 -1.240 1.900 ;
        RECT -17.750 1.600 -1.240 1.750 ;
        RECT -17.750 1.450 -17.430 1.600 ;
        RECT -11.950 1.450 -11.630 1.600 ;
    END
    PORT
      LAYER met1 ;
        RECT -1.560 1.600 -1.240 1.900 ;
        RECT -0.030 1.600 0.310 7.450 ;
        RECT -1.560 1.570 -1.130 1.600 ;
        RECT -0.530 1.570 0.310 1.600 ;
        RECT -1.560 1.540 0.310 1.570 ;
        RECT -1.410 1.490 0.310 1.540 ;
        RECT -1.380 1.460 0.310 1.490 ;
        RECT -1.350 1.440 0.310 1.460 ;
        RECT -1.280 1.430 -0.320 1.440 ;
        RECT -0.030 1.400 0.310 1.440 ;
      LAYER via ;
        RECT -1.530 1.620 -1.270 1.880 ;
    END
  END VGND
  PIN OUTPUT2
    ANTENNADIFFAREA 0.308800 ;
    PORT
      LAYER met2 ;
        RECT -0.990 4.140 -0.680 4.190 ;
        RECT 1.300 4.140 1.610 4.270 ;
        RECT -0.990 3.920 1.930 4.140 ;
        RECT -0.990 3.860 -0.680 3.920 ;
    END
  END OUTPUT2
  PIN OUTPUT1
    ANTENNADIFFAREA 0.308800 ;
    PORT
      LAYER met2 ;
        RECT -0.990 4.970 -0.680 5.030 ;
        RECT 1.310 4.970 1.620 4.990 ;
        RECT -0.990 4.740 1.930 4.970 ;
        RECT -0.990 4.700 -0.680 4.740 ;
        RECT 1.310 4.660 1.620 4.740 ;
    END
  END OUTPUT1
  PIN GATESEL1
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT -25.400 5.990 -25.210 7.450 ;
        RECT -25.430 5.960 -25.210 5.990 ;
        RECT -25.440 5.690 -25.190 5.960 ;
        RECT -25.440 5.680 -25.200 5.690 ;
        RECT -25.430 5.440 -25.200 5.680 ;
        RECT -25.400 3.410 -25.240 5.440 ;
        RECT -25.430 3.170 -25.200 3.410 ;
        RECT -25.440 3.160 -25.200 3.170 ;
        RECT -25.440 2.890 -25.190 3.160 ;
        RECT -25.430 2.860 -25.210 2.890 ;
        RECT -25.400 1.400 -25.210 2.860 ;
    END
  END GATESEL1
  PIN GATESEL2
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT -4.160 5.990 -3.970 7.450 ;
        RECT -4.160 5.960 -3.940 5.990 ;
        RECT -4.180 5.690 -3.930 5.960 ;
        RECT -4.170 5.680 -3.930 5.690 ;
        RECT -4.170 5.440 -3.940 5.680 ;
        RECT -4.130 3.410 -3.970 5.440 ;
        RECT -4.170 3.170 -3.940 3.410 ;
        RECT -4.170 3.160 -3.930 3.170 ;
        RECT -4.180 2.890 -3.930 3.160 ;
        RECT -4.160 2.860 -3.940 2.890 ;
        RECT -4.160 1.400 -3.970 2.860 ;
    END
  END GATESEL2
  PIN DRAIN1
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER met2 ;
        RECT -23.760 6.960 -23.440 6.970 ;
        RECT -24.000 6.950 -23.440 6.960 ;
        RECT -5.680 6.950 -5.370 6.960 ;
        RECT -26.170 6.770 -3.200 6.950 ;
        RECT -24.000 6.630 -23.690 6.770 ;
        RECT -5.680 6.630 -5.370 6.770 ;
    END
  END DRAIN1
  PIN DRAIN2
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER met2 ;
        RECT -24.000 2.080 -23.690 2.220 ;
        RECT -26.170 2.070 -23.690 2.080 ;
        RECT -5.680 2.080 -5.370 2.220 ;
        RECT -5.680 2.070 -3.200 2.080 ;
        RECT -26.170 1.920 -3.200 2.070 ;
        RECT -26.170 1.900 -23.690 1.920 ;
        RECT -24.000 1.890 -23.690 1.900 ;
        RECT -5.680 1.900 -3.200 1.920 ;
        RECT -5.680 1.890 -5.370 1.900 ;
    END
  END DRAIN2
  PIN VIN12
    ANTENNADIFFAREA 0.217200 ;
    PORT
      LAYER met1 ;
        RECT -23.510 4.020 -23.320 4.150 ;
        RECT -23.530 3.730 -23.300 4.020 ;
        RECT -23.510 2.110 -23.320 3.730 ;
        RECT -23.510 1.900 -23.280 2.110 ;
        RECT -23.520 1.820 -23.280 1.900 ;
        RECT -23.520 1.400 -23.290 1.820 ;
    END
  END VIN12
  PIN GATE2
    ANTENNADIFFAREA 0.434600 ;
    PORT
      LAYER met1 ;
        RECT -23.060 6.520 -22.870 7.450 ;
        RECT -23.070 6.230 -22.840 6.520 ;
        RECT -23.060 4.200 -22.870 6.230 ;
        RECT -23.070 3.910 -22.840 4.200 ;
        RECT -23.060 2.620 -22.870 3.910 ;
        RECT -23.080 2.330 -22.850 2.620 ;
        RECT -23.060 1.400 -22.870 2.330 ;
    END
  END GATE2
  PIN RUN
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER met1 ;
        RECT -21.570 2.920 -21.390 7.450 ;
        RECT -21.630 2.580 -21.340 2.920 ;
        RECT -21.570 1.400 -21.390 2.580 ;
    END
  END RUN
  OBS
      LAYER nwell ;
        RECT -21.130 5.060 -18.410 6.710 ;
        RECT -21.130 5.020 -18.420 5.060 ;
        RECT -21.130 3.690 -18.420 3.730 ;
        RECT -21.130 2.040 -18.410 3.690 ;
      LAYER li1 ;
        RECT -2.220 7.400 -2.050 7.450 ;
        RECT -2.220 7.140 -1.660 7.400 ;
        RECT -0.750 7.150 -0.550 7.190 ;
        RECT -2.220 7.120 -2.050 7.140 ;
        RECT -25.770 6.770 -25.570 7.120 ;
        RECT -24.290 6.870 -23.760 7.040 ;
        RECT -23.520 7.020 -23.330 7.050 ;
        RECT -23.520 6.850 -22.460 7.020 ;
        RECT -5.610 6.870 -5.080 7.040 ;
        RECT -23.520 6.820 -23.330 6.850 ;
        RECT -25.780 6.740 -25.570 6.770 ;
        RECT -25.780 6.160 -25.560 6.740 ;
        RECT -25.780 6.150 -25.570 6.160 ;
        RECT -25.400 5.980 -25.210 5.990 ;
        RECT -25.410 5.690 -25.210 5.980 ;
        RECT -25.470 5.360 -25.200 5.690 ;
        RECT -25.010 4.880 -24.840 6.490 ;
        RECT -24.180 5.390 -24.010 6.480 ;
        RECT -23.050 6.460 -22.860 6.490 ;
        RECT -23.590 6.290 -22.860 6.460 ;
        RECT -22.630 6.460 -22.460 6.850 ;
        RECT -3.800 6.770 -3.600 7.120 ;
        RECT -3.800 6.740 -3.590 6.770 ;
        RECT -22.630 6.290 -21.890 6.460 ;
        RECT -23.050 6.260 -22.860 6.290 ;
        RECT -20.830 5.670 -20.600 6.190 ;
        RECT -23.590 5.500 -20.600 5.670 ;
        RECT -24.410 5.350 -24.010 5.390 ;
        RECT -24.420 5.160 -24.010 5.350 ;
        RECT -15.630 5.310 -15.080 5.740 ;
        RECT -14.290 5.310 -13.740 5.740 ;
        RECT -10.660 5.500 -10.430 6.190 ;
        RECT -5.360 5.960 -5.190 6.480 ;
        RECT -5.520 5.700 -5.190 5.960 ;
        RECT -24.410 5.130 -24.010 5.160 ;
        RECT -25.020 4.690 -24.840 4.880 ;
        RECT -24.180 4.790 -24.010 5.130 ;
        RECT -23.520 4.880 -23.330 5.060 ;
        RECT -23.590 4.710 -23.240 4.880 ;
        RECT -22.670 4.300 -22.460 4.730 ;
        RECT -22.240 4.710 -21.900 4.880 ;
        RECT -22.650 4.280 -22.480 4.300 ;
        RECT -25.020 3.970 -24.840 4.160 ;
        RECT -25.470 3.160 -25.200 3.490 ;
        RECT -25.410 2.870 -25.210 3.160 ;
        RECT -25.400 2.860 -25.210 2.870 ;
        RECT -25.780 2.690 -25.570 2.700 ;
        RECT -25.780 2.110 -25.560 2.690 ;
        RECT -25.010 2.360 -24.840 3.970 ;
        RECT -24.180 3.700 -24.010 4.060 ;
        RECT -23.590 3.970 -23.240 4.140 ;
        RECT -23.050 4.120 -22.860 4.170 ;
        RECT -22.150 4.140 -21.980 4.710 ;
        RECT -17.870 4.480 -17.680 4.880 ;
        RECT -11.690 4.480 -11.500 4.880 ;
        RECT -5.360 4.790 -5.190 5.700 ;
        RECT -4.530 4.880 -4.360 6.490 ;
        RECT -3.810 6.160 -3.590 6.740 ;
        RECT -3.800 6.150 -3.590 6.160 ;
        RECT -2.800 6.040 -2.620 6.970 ;
        RECT -0.980 6.890 -0.550 7.150 ;
        RECT -2.070 6.710 -1.740 6.880 ;
        RECT -0.750 6.860 -0.550 6.890 ;
        RECT -1.990 6.570 -1.740 6.710 ;
        RECT -1.990 6.310 -1.510 6.570 ;
        RECT -1.160 6.500 -0.990 6.540 ;
        RECT -0.750 6.500 -0.550 6.530 ;
        RECT -2.920 6.010 -2.600 6.040 ;
        RECT -4.160 5.980 -3.970 5.990 ;
        RECT -4.160 5.690 -3.960 5.980 ;
        RECT -2.920 5.820 -2.590 6.010 ;
        RECT -2.920 5.780 -2.600 5.820 ;
        RECT -4.170 5.360 -3.880 5.690 ;
        RECT -4.530 4.690 -4.350 4.880 ;
        RECT -17.870 4.470 -17.490 4.480 ;
        RECT -21.230 4.290 -17.490 4.470 ;
        RECT -17.870 4.250 -17.490 4.290 ;
        RECT -11.880 4.470 -11.500 4.480 ;
        RECT -11.880 4.290 -8.140 4.470 ;
        RECT -11.880 4.250 -11.500 4.290 ;
        RECT -23.050 4.110 -22.820 4.120 ;
        RECT -22.240 4.110 -21.900 4.140 ;
        RECT -23.050 3.970 -21.900 4.110 ;
        RECT -23.510 3.760 -23.320 3.970 ;
        RECT -23.050 3.940 -22.070 3.970 ;
        RECT -22.910 3.910 -22.070 3.940 ;
        RECT -17.870 3.870 -17.680 4.250 ;
        RECT -24.420 3.660 -24.010 3.700 ;
        RECT -24.430 3.470 -24.010 3.660 ;
        RECT -15.630 3.580 -15.080 4.010 ;
        RECT -14.290 3.580 -13.740 4.010 ;
        RECT -11.690 3.870 -11.500 4.250 ;
        RECT -24.420 3.440 -24.010 3.470 ;
        RECT -24.180 2.370 -24.010 3.440 ;
        RECT -23.590 3.250 -20.660 3.350 ;
        RECT -23.590 3.180 -20.600 3.250 ;
        RECT -21.570 2.860 -21.400 2.920 ;
        RECT -21.590 2.650 -21.380 2.860 ;
        RECT -23.060 2.560 -22.870 2.590 ;
        RECT -21.570 2.580 -21.400 2.650 ;
        RECT -20.830 2.560 -20.600 3.180 ;
        RECT -10.660 2.560 -10.430 3.290 ;
        RECT -5.360 3.200 -5.190 4.060 ;
        RECT -5.520 2.940 -5.190 3.200 ;
        RECT -23.590 2.390 -22.870 2.560 ;
        RECT -23.060 2.360 -22.870 2.390 ;
        RECT -22.700 2.390 -21.890 2.560 ;
        RECT -25.780 2.080 -25.570 2.110 ;
        RECT -25.770 1.730 -25.570 2.080 ;
        RECT -23.490 2.050 -23.300 2.080 ;
        RECT -22.700 2.050 -22.510 2.390 ;
        RECT -5.360 2.370 -5.190 2.940 ;
        RECT -4.530 3.970 -4.350 4.160 ;
        RECT -4.530 2.360 -4.360 3.970 ;
        RECT -4.170 3.160 -3.880 3.490 ;
        RECT -4.160 2.870 -3.960 3.160 ;
        RECT -4.160 2.860 -3.970 2.870 ;
        RECT -3.800 2.690 -3.590 2.700 ;
        RECT -3.810 2.110 -3.590 2.690 ;
        RECT -24.290 1.810 -23.760 1.980 ;
        RECT -23.490 1.870 -22.510 2.050 ;
        RECT -3.800 2.080 -3.590 2.110 ;
        RECT -23.490 1.850 -23.300 1.870 ;
        RECT -5.610 1.810 -5.080 1.980 ;
        RECT -3.800 1.730 -3.600 2.080 ;
        RECT -2.800 1.870 -2.620 5.780 ;
        RECT -1.990 4.930 -1.820 6.310 ;
        RECT -1.160 6.240 -0.550 6.500 ;
        RECT -1.160 6.210 -0.990 6.240 ;
        RECT -0.750 6.200 -0.550 6.240 ;
        RECT -0.160 6.200 0.390 7.190 ;
        RECT 1.210 7.040 1.840 7.210 ;
        RECT 1.210 6.940 1.600 7.040 ;
        RECT 1.210 6.910 1.590 6.940 ;
        RECT 1.210 6.760 1.570 6.910 ;
        RECT 0.860 6.590 1.570 6.760 ;
        RECT 0.860 5.840 1.560 6.150 ;
        RECT -1.160 5.650 -0.990 5.680 ;
        RECT -0.750 5.650 -0.550 5.690 ;
        RECT -1.160 5.390 -0.550 5.650 ;
        RECT -1.160 5.350 -0.990 5.390 ;
        RECT -0.750 5.360 -0.550 5.390 ;
        RECT -0.750 5.000 -0.550 5.030 ;
        RECT -2.190 4.730 -1.870 4.760 ;
        RECT -0.980 4.740 -0.550 5.000 ;
        RECT -2.190 4.540 -1.860 4.730 ;
        RECT -0.750 4.700 -0.550 4.740 ;
        RECT -0.160 4.700 0.390 5.690 ;
        RECT 0.710 5.610 1.560 5.840 ;
        RECT 0.860 5.270 1.560 5.610 ;
        RECT 1.320 4.910 1.640 4.950 ;
        RECT 1.320 4.850 1.650 4.910 ;
        RECT 0.850 4.720 1.650 4.850 ;
        RECT 0.850 4.690 1.640 4.720 ;
        RECT 0.850 4.670 1.550 4.690 ;
        RECT -2.190 4.500 -1.870 4.540 ;
        RECT -2.190 4.420 -2.020 4.500 ;
        RECT -2.240 4.250 -2.020 4.420 ;
        RECT -2.240 4.090 -2.070 4.250 ;
        RECT 1.310 4.190 1.630 4.230 ;
        RECT -0.750 4.150 -0.550 4.190 ;
        RECT -1.710 3.830 -1.520 3.950 ;
        RECT -0.980 3.890 -0.550 4.150 ;
        RECT -0.750 3.860 -0.550 3.890 ;
        RECT -2.070 3.720 -1.520 3.830 ;
        RECT -2.070 3.660 -1.530 3.720 ;
        RECT -1.990 1.880 -1.820 3.660 ;
        RECT -1.160 3.500 -0.990 3.540 ;
        RECT -0.750 3.500 -0.550 3.530 ;
        RECT -1.160 3.240 -0.550 3.500 ;
        RECT -1.160 3.210 -0.990 3.240 ;
        RECT -0.750 3.200 -0.550 3.240 ;
        RECT -0.160 3.200 0.390 4.190 ;
        RECT 0.850 4.010 1.640 4.190 ;
        RECT 1.310 4.000 1.640 4.010 ;
        RECT 1.310 3.970 1.630 4.000 ;
        RECT 0.860 3.250 1.560 3.590 ;
        RECT 0.710 3.020 1.560 3.250 ;
        RECT 0.860 2.710 1.560 3.020 ;
        RECT -1.160 2.650 -0.990 2.680 ;
        RECT -0.750 2.650 -0.550 2.690 ;
        RECT -1.160 2.390 -0.550 2.650 ;
        RECT -1.160 2.350 -0.990 2.390 ;
        RECT -0.750 2.360 -0.550 2.390 ;
        RECT -0.750 2.000 -0.550 2.030 ;
        RECT -0.980 1.740 -0.550 2.000 ;
        RECT -0.750 1.700 -0.550 1.740 ;
        RECT -0.160 1.700 0.390 2.690 ;
        RECT 0.860 2.100 1.570 2.270 ;
        RECT 1.210 1.820 1.570 2.100 ;
        RECT 1.210 1.650 1.840 1.820 ;
      LAYER mcon ;
        RECT -1.890 7.180 -1.720 7.350 ;
        RECT -23.940 6.870 -23.760 7.040 ;
        RECT -23.510 6.850 -23.340 7.020 ;
        RECT -25.750 6.570 -25.580 6.740 ;
        RECT -25.400 5.730 -25.220 5.920 ;
        RECT -23.040 6.290 -22.870 6.460 ;
        RECT -3.790 6.570 -3.620 6.740 ;
        RECT -20.800 5.990 -20.630 6.160 ;
        RECT -10.630 5.990 -10.460 6.160 ;
        RECT -20.800 5.540 -20.630 5.710 ;
        RECT -24.320 5.170 -24.150 5.340 ;
        RECT -15.350 5.390 -15.080 5.660 ;
        RECT -14.290 5.390 -14.020 5.660 ;
        RECT -10.630 5.540 -10.460 5.710 ;
        RECT -5.460 5.740 -5.290 5.910 ;
        RECT -23.510 4.860 -23.340 5.030 ;
        RECT -0.920 6.930 -0.750 7.100 ;
        RECT 0.060 6.610 0.230 6.780 ;
        RECT 1.330 6.950 1.500 7.120 ;
        RECT -1.740 6.350 -1.570 6.520 ;
        RECT -4.150 5.730 -3.970 5.920 ;
        RECT -2.860 5.830 -2.690 6.000 ;
        RECT -17.670 4.280 -17.500 4.450 ;
        RECT -11.870 4.280 -11.700 4.450 ;
        RECT -25.400 2.930 -25.220 3.120 ;
        RECT -23.040 3.970 -22.870 4.140 ;
        RECT -23.500 3.790 -23.330 3.960 ;
        RECT -24.330 3.480 -24.160 3.650 ;
        RECT -15.350 3.660 -15.080 3.930 ;
        RECT -14.290 3.660 -14.020 3.930 ;
        RECT -20.800 3.040 -20.630 3.210 ;
        RECT -20.800 2.590 -20.630 2.760 ;
        RECT -10.630 3.040 -10.460 3.210 ;
        RECT -5.460 2.980 -5.290 3.150 ;
        RECT -10.630 2.590 -10.460 2.760 ;
        RECT -23.050 2.390 -22.880 2.560 ;
        RECT -25.750 2.110 -25.580 2.280 ;
        RECT -4.150 2.930 -3.970 3.120 ;
        RECT -3.790 2.110 -3.620 2.280 ;
        RECT -23.940 1.810 -23.760 1.980 ;
        RECT -23.480 1.880 -23.310 2.050 ;
        RECT -0.970 6.280 -0.800 6.450 ;
        RECT -0.970 5.440 -0.800 5.610 ;
        RECT 0.720 5.640 0.890 5.810 ;
        RECT 0.060 5.110 0.230 5.280 ;
        RECT -0.920 4.790 -0.750 4.960 ;
        RECT -2.130 4.550 -1.960 4.720 ;
        RECT 1.380 4.730 1.550 4.900 ;
        RECT -1.700 3.750 -1.530 3.920 ;
        RECT -0.920 3.930 -0.750 4.100 ;
        RECT 1.370 4.010 1.540 4.180 ;
        RECT 0.060 3.610 0.230 3.780 ;
        RECT -0.970 3.280 -0.800 3.450 ;
        RECT 0.720 3.050 0.890 3.220 ;
        RECT -0.970 2.440 -0.800 2.610 ;
        RECT 0.060 2.110 0.230 2.280 ;
        RECT -0.920 1.790 -0.750 1.960 ;
        RECT 1.290 1.760 1.460 1.930 ;
      LAYER met1 ;
        RECT -25.810 7.430 -25.650 7.450 ;
        RECT -25.970 7.130 -25.650 7.430 ;
        RECT -25.810 6.800 -25.650 7.130 ;
        RECT -25.810 6.250 -25.540 6.800 ;
        RECT -24.000 6.630 -23.690 7.070 ;
        RECT -25.820 6.200 -25.540 6.250 ;
        RECT -25.820 6.110 -25.650 6.200 ;
        RECT -25.810 2.740 -25.650 6.110 ;
        RECT -20.850 5.450 -20.590 6.240 ;
        RECT -24.400 5.100 -24.080 5.420 ;
        RECT -25.050 4.590 -24.810 5.010 ;
        RECT -25.080 4.270 -24.810 4.590 ;
        RECT -25.050 3.840 -24.810 4.270 ;
        RECT -24.410 3.410 -24.090 3.730 ;
        RECT -25.820 2.650 -25.650 2.740 ;
        RECT -25.820 2.600 -25.540 2.650 ;
        RECT -25.810 2.050 -25.540 2.600 ;
        RECT -20.850 2.510 -20.590 3.300 ;
        RECT -25.810 1.400 -25.650 2.050 ;
        RECT -24.000 1.780 -23.690 2.220 ;
        RECT -17.700 1.750 -17.470 7.450 ;
        RECT -11.900 1.750 -11.670 7.450 ;
        RECT -1.970 7.110 -1.650 7.430 ;
        RECT -5.680 6.630 -5.370 7.070 ;
        RECT -0.990 6.860 -0.670 7.180 ;
        RECT 1.260 6.880 1.580 7.200 ;
        RECT -1.820 6.280 -1.500 6.600 ;
        RECT -1.040 6.210 -0.720 6.530 ;
        RECT -5.530 5.670 -5.210 5.990 ;
        RECT -2.930 5.750 -2.610 6.070 ;
        RECT -1.710 5.590 -1.500 5.700 ;
        RECT -1.730 5.270 -1.470 5.590 ;
        RECT -1.040 5.360 -0.720 5.680 ;
        RECT -4.560 4.880 -4.320 5.010 ;
        RECT -4.560 4.560 -4.300 4.880 ;
        RECT -2.200 4.470 -1.880 4.790 ;
        RECT -4.560 3.960 -4.300 4.280 ;
        RECT -1.710 3.980 -1.500 5.270 ;
        RECT -0.990 4.710 -0.670 5.030 ;
        RECT 1.310 4.660 1.630 4.980 ;
        RECT -4.560 3.840 -4.320 3.960 ;
        RECT -1.730 3.690 -1.500 3.980 ;
        RECT -0.990 3.860 -0.670 4.180 ;
        RECT 1.300 3.940 1.620 4.260 ;
        RECT -5.530 2.910 -5.210 3.230 ;
        RECT -1.040 3.210 -0.720 3.530 ;
        RECT -1.040 2.360 -0.720 2.680 ;
        RECT -5.680 1.780 -5.370 2.220 ;
        RECT -17.750 1.450 -17.430 1.750 ;
        RECT -11.950 1.450 -11.630 1.750 ;
        RECT -0.990 1.710 -0.670 2.030 ;
        RECT 1.220 1.690 1.540 2.010 ;
        RECT -17.700 1.400 -17.470 1.450 ;
        RECT -11.900 1.400 -11.670 1.450 ;
      LAYER via ;
        RECT -25.940 7.150 -25.680 7.410 ;
        RECT -23.980 6.660 -23.720 6.920 ;
        RECT -24.370 5.130 -24.110 5.390 ;
        RECT -25.080 4.300 -24.820 4.560 ;
        RECT -24.380 3.440 -24.120 3.700 ;
        RECT -23.980 1.930 -23.720 2.190 ;
        RECT -1.940 7.140 -1.680 7.400 ;
        RECT -5.650 6.660 -5.390 6.920 ;
        RECT -0.960 6.890 -0.700 7.150 ;
        RECT 1.290 6.910 1.550 7.170 ;
        RECT -1.790 6.310 -1.530 6.570 ;
        RECT -1.010 6.240 -0.750 6.500 ;
        RECT -5.500 5.700 -5.240 5.960 ;
        RECT -2.900 5.780 -2.640 6.040 ;
        RECT -1.730 5.300 -1.470 5.560 ;
        RECT -1.010 5.390 -0.750 5.650 ;
        RECT -4.560 4.590 -4.300 4.850 ;
        RECT -2.170 4.500 -1.910 4.760 ;
        RECT -4.560 3.990 -4.300 4.250 ;
        RECT -0.960 4.740 -0.700 5.000 ;
        RECT 1.340 4.690 1.600 4.950 ;
        RECT -0.960 3.890 -0.700 4.150 ;
        RECT 1.330 3.970 1.590 4.230 ;
        RECT -1.010 3.240 -0.750 3.500 ;
        RECT -5.500 2.940 -5.240 3.200 ;
        RECT -1.010 2.390 -0.750 2.650 ;
        RECT -5.650 1.930 -5.390 2.190 ;
        RECT -17.720 1.470 -17.460 1.730 ;
        RECT -11.920 1.470 -11.660 1.730 ;
        RECT -0.960 1.740 -0.700 2.000 ;
        RECT 1.250 1.720 1.510 1.980 ;
      LAYER met2 ;
        RECT -0.990 7.110 -0.680 7.190 ;
        RECT 1.260 7.110 1.570 7.210 ;
        RECT -0.990 6.880 1.570 7.110 ;
        RECT -0.990 6.860 -0.680 6.880 ;
        RECT -1.810 6.570 -1.500 6.610 ;
        RECT -1.990 6.460 -1.270 6.570 ;
        RECT -1.040 6.460 -0.730 6.540 ;
        RECT -1.990 6.320 -0.730 6.460 ;
        RECT -1.810 6.280 -0.730 6.320 ;
        RECT -1.540 6.250 -0.730 6.280 ;
        RECT -1.540 6.210 -1.270 6.250 ;
        RECT -1.040 6.210 -0.730 6.250 ;
        RECT -5.530 5.930 -5.220 6.000 ;
        RECT -2.930 5.930 -2.620 6.070 ;
        RECT -5.530 5.740 -2.620 5.930 ;
        RECT -5.530 5.710 -2.930 5.740 ;
        RECT -5.530 5.670 -5.220 5.710 ;
        RECT -1.470 5.640 -1.270 5.650 ;
        RECT -1.040 5.640 -0.730 5.680 ;
        RECT -1.470 5.560 -0.730 5.640 ;
        RECT -1.760 5.540 -0.730 5.560 ;
        RECT -1.810 5.430 -0.730 5.540 ;
        RECT -24.390 5.410 -24.080 5.430 ;
        RECT -14.660 5.410 -6.670 5.420 ;
        RECT -24.390 5.220 -6.670 5.410 ;
        RECT -1.810 5.300 -1.250 5.430 ;
        RECT -1.040 5.350 -0.730 5.430 ;
        RECT -1.810 5.290 -1.340 5.300 ;
        RECT -24.390 5.100 -24.080 5.220 ;
        RECT -25.110 4.530 -24.790 4.560 ;
        RECT -8.070 4.540 -7.850 4.550 ;
        RECT -14.650 4.530 -7.820 4.540 ;
        RECT -25.110 4.300 -7.820 4.530 ;
        RECT -6.890 4.500 -6.670 5.220 ;
        RECT -14.650 4.290 -7.820 4.300 ;
        RECT -24.400 3.550 -24.090 3.740 ;
        RECT -14.650 3.550 -11.140 3.560 ;
        RECT -24.400 3.410 -11.140 3.550 ;
        RECT -24.370 3.370 -11.140 3.410 ;
        RECT -24.370 3.360 -14.650 3.370 ;
        RECT -11.370 2.770 -11.140 3.370 ;
        RECT -8.110 3.120 -7.820 4.290 ;
        RECT -6.920 4.460 -6.670 4.500 ;
        RECT -6.920 3.820 -6.660 4.460 ;
        RECT -6.920 3.610 -2.790 3.820 ;
        RECT -3.000 3.470 -2.790 3.610 ;
        RECT -1.040 3.470 -0.730 3.540 ;
        RECT -3.000 3.260 -0.730 3.470 ;
        RECT -1.340 3.250 -0.730 3.260 ;
        RECT -5.530 3.170 -5.220 3.240 ;
        RECT -1.040 3.210 -0.730 3.250 ;
        RECT -5.530 3.120 -3.200 3.170 ;
        RECT -8.110 2.960 -3.200 3.120 ;
        RECT -8.110 2.900 -5.220 2.960 ;
        RECT -8.110 2.890 -7.820 2.900 ;
        RECT -11.370 2.620 -11.150 2.770 ;
        RECT -1.040 2.670 -0.730 2.680 ;
        RECT -7.000 2.620 -0.730 2.670 ;
        RECT -11.370 2.460 -0.730 2.620 ;
        RECT -11.370 2.400 -6.610 2.460 ;
        RECT -1.340 2.430 -0.730 2.460 ;
        RECT -1.040 2.350 -0.730 2.430 ;
        RECT -0.990 1.980 -0.680 2.030 ;
        RECT 1.220 1.980 1.530 2.020 ;
        RECT -0.990 1.750 1.720 1.980 ;
        RECT -0.990 1.700 -0.680 1.750 ;
        RECT 1.220 1.690 1.530 1.750 ;
  END
END sky130_hilas_TA2Cell_1FG_Strong

MACRO sky130_hilas_TA2Cell_NoFG
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TA2Cell_NoFG ;
  ORIGIN 14.730 -1.350 ;
  SIZE 17.920 BY 6.150 ;
  PIN COLSEL1
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT -4.160 5.990 -3.970 7.450 ;
        RECT -4.160 5.960 -3.940 5.990 ;
        RECT -4.180 5.690 -3.930 5.960 ;
        RECT -4.170 5.680 -3.930 5.690 ;
        RECT -4.170 5.440 -3.940 5.680 ;
        RECT -4.130 3.410 -3.970 5.440 ;
        RECT -4.170 3.170 -3.940 3.410 ;
        RECT -4.170 3.160 -3.930 3.170 ;
        RECT -4.180 2.890 -3.930 3.160 ;
        RECT -4.160 2.860 -3.940 2.890 ;
        RECT -4.160 1.400 -3.970 2.860 ;
    END
  END COLSEL1
  PIN VIN12
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -2.260 1.670 -1.950 1.740 ;
        RECT -2.860 1.420 -1.950 1.670 ;
        RECT -2.260 1.410 -1.950 1.420 ;
    END
  END VIN12
  PIN VIN21
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -0.940 4.750 -0.630 4.790 ;
        RECT -1.030 4.740 -0.600 4.750 ;
        RECT -1.260 4.510 -0.160 4.740 ;
        RECT -0.940 4.460 -0.630 4.510 ;
    END
  END VIN21
  PIN VIN22
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -1.300 7.430 -1.050 7.440 ;
        RECT -0.700 7.430 -0.390 7.440 ;
        RECT -1.300 7.180 -0.390 7.430 ;
        RECT -0.700 7.110 -0.390 7.180 ;
    END
  END VIN22
  PIN OUTPUT1
    ANTENNADIFFAREA 0.308800 ;
    PORT
      LAYER met2 ;
        RECT 0.270 4.140 0.580 4.190 ;
        RECT 2.560 4.140 2.870 4.270 ;
        RECT 0.270 3.920 3.190 4.140 ;
        RECT 0.270 3.860 0.580 3.920 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    ANTENNADIFFAREA 0.308800 ;
    PORT
      LAYER met2 ;
        RECT 0.270 4.970 0.580 5.030 ;
        RECT 2.570 4.970 2.880 4.990 ;
        RECT 0.270 4.740 3.190 4.970 ;
        RECT 0.270 4.700 0.580 4.740 ;
        RECT 2.570 4.660 2.880 4.740 ;
    END
  END OUTPUT2
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 1.230 6.000 1.570 6.090 ;
        RECT -1.120 5.810 1.570 6.000 ;
        RECT -1.120 5.240 -0.930 5.810 ;
        RECT 1.230 5.760 1.570 5.810 ;
        RECT -11.910 5.050 -0.930 5.240 ;
        RECT -11.910 4.870 -11.720 5.050 ;
        RECT -11.930 3.880 -11.580 4.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.230 1.400 1.570 7.450 ;
      LAYER via ;
        RECT 1.270 5.790 1.530 6.050 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 1.920 7.270 3.190 7.450 ;
        RECT 1.910 1.400 3.190 7.270 ;
      LAYER met1 ;
        RECT 1.900 5.870 2.170 7.450 ;
        RECT 1.900 5.580 2.180 5.870 ;
        RECT 1.900 3.280 2.170 5.580 ;
        RECT 1.900 2.990 2.180 3.280 ;
        RECT 1.900 1.400 2.170 2.990 ;
    END
  END VPWR
  PIN DRAIN1
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT -5.680 6.950 -5.370 6.960 ;
        RECT -14.730 6.770 -3.200 6.950 ;
        RECT -5.680 6.630 -5.370 6.770 ;
    END
  END DRAIN1
  PIN DRAIN2
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT -5.680 2.080 -5.370 2.220 ;
        RECT -5.680 2.070 -3.200 2.080 ;
        RECT -14.730 1.920 -3.200 2.070 ;
        RECT -5.680 1.900 -3.200 1.920 ;
        RECT -5.680 1.890 -5.370 1.900 ;
    END
  END DRAIN2
  PIN VTUN
    ANTENNADIFFAREA 2.516100 ;
    PORT
      LAYER nwell ;
        RECT -14.720 6.700 -12.990 7.450 ;
        RECT -14.720 5.550 -12.980 6.700 ;
        RECT -14.710 3.310 -12.980 5.550 ;
        RECT -14.720 3.130 -12.980 3.310 ;
        RECT -14.720 1.410 -12.990 3.130 ;
      LAYER met1 ;
        RECT -14.380 1.400 -13.960 7.450 ;
    END
  END VTUN
  PIN GATE1
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT -10.960 5.060 -8.240 6.710 ;
        RECT -10.960 5.020 -8.250 5.060 ;
        RECT -10.960 3.690 -8.250 3.730 ;
        RECT -10.960 2.040 -8.240 3.690 ;
      LAYER met1 ;
        RECT -10.680 6.240 -10.450 7.450 ;
        RECT -10.680 5.450 -10.420 6.240 ;
        RECT -10.680 3.300 -10.450 5.450 ;
        RECT -10.680 2.510 -10.420 3.300 ;
        RECT -10.680 1.400 -10.450 2.510 ;
    END
  END GATE1
  PIN VINJ
    ANTENNADIFFAREA 1.574400 ;
    PORT
      LAYER nwell ;
        RECT -6.510 7.450 -3.200 7.500 ;
        RECT -6.510 7.440 -1.650 7.450 ;
        RECT -6.510 1.410 -0.090 7.440 ;
        RECT -6.510 1.350 -3.200 1.410 ;
        RECT -1.950 1.400 -0.090 1.410 ;
      LAYER met2 ;
        RECT -4.590 4.590 -4.270 4.850 ;
        RECT -4.550 4.570 -3.370 4.590 ;
        RECT -4.550 4.310 -3.330 4.570 ;
        RECT -4.550 4.250 -3.370 4.310 ;
        RECT -4.590 4.240 -3.370 4.250 ;
        RECT -4.590 3.990 -4.270 4.240 ;
    END
  END VINJ
  PIN VIN11
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -2.500 4.340 -2.190 4.390 ;
        RECT -2.820 4.110 -1.720 4.340 ;
        RECT -2.820 4.100 -2.160 4.110 ;
        RECT -2.500 4.060 -2.190 4.100 ;
    END
  END VIN11
  OBS
      LAYER li1 ;
        RECT -0.960 7.400 -0.790 7.450 ;
        RECT -0.960 7.140 -0.400 7.400 ;
        RECT 0.510 7.150 0.710 7.190 ;
        RECT -0.960 7.120 -0.790 7.140 ;
        RECT -5.610 6.870 -5.080 7.040 ;
        RECT -3.800 6.770 -3.600 7.120 ;
        RECT -3.800 6.740 -3.590 6.770 ;
        RECT -14.290 5.310 -13.740 5.740 ;
        RECT -10.660 5.500 -10.430 6.190 ;
        RECT -5.360 5.960 -5.190 6.480 ;
        RECT -5.520 5.700 -5.190 5.960 ;
        RECT -11.900 4.470 -11.440 4.880 ;
        RECT -5.360 4.790 -5.190 5.700 ;
        RECT -4.530 4.880 -4.360 6.490 ;
        RECT -3.810 6.160 -3.590 6.740 ;
        RECT -3.800 6.150 -3.590 6.160 ;
        RECT -4.160 5.980 -3.970 5.990 ;
        RECT -4.160 5.690 -3.960 5.980 ;
        RECT -4.170 5.360 -3.880 5.690 ;
        RECT -4.530 4.690 -4.350 4.880 ;
        RECT -11.900 4.290 -8.140 4.470 ;
        RECT -14.290 3.580 -13.740 4.010 ;
        RECT -11.900 3.870 -11.440 4.290 ;
        RECT -10.660 2.560 -10.430 3.290 ;
        RECT -5.360 3.200 -5.190 4.060 ;
        RECT -5.520 2.940 -5.190 3.200 ;
        RECT -5.360 2.370 -5.190 2.940 ;
        RECT -4.530 3.970 -4.350 4.160 ;
        RECT -4.530 2.360 -4.360 3.970 ;
        RECT -4.170 3.160 -3.880 3.490 ;
        RECT -4.160 2.870 -3.960 3.160 ;
        RECT -3.100 3.070 -2.920 6.980 ;
        RECT -2.290 5.190 -2.120 6.970 ;
        RECT -1.540 6.040 -1.360 6.970 ;
        RECT 0.280 6.890 0.710 7.150 ;
        RECT -0.810 6.710 -0.480 6.880 ;
        RECT 0.510 6.860 0.710 6.890 ;
        RECT -0.730 6.570 -0.480 6.710 ;
        RECT -0.730 6.310 -0.250 6.570 ;
        RECT 0.100 6.500 0.270 6.540 ;
        RECT 0.510 6.500 0.710 6.530 ;
        RECT -1.660 6.010 -1.340 6.040 ;
        RECT -1.660 5.820 -1.330 6.010 ;
        RECT -1.660 5.780 -1.340 5.820 ;
        RECT -2.370 5.130 -1.830 5.190 ;
        RECT -2.370 5.020 -1.820 5.130 ;
        RECT -2.010 4.900 -1.820 5.020 ;
        RECT -2.540 4.600 -2.370 4.760 ;
        RECT -2.540 4.430 -2.320 4.600 ;
        RECT -2.490 4.350 -2.320 4.430 ;
        RECT -2.490 4.310 -2.170 4.350 ;
        RECT -2.490 4.120 -2.160 4.310 ;
        RECT -2.490 4.090 -2.170 4.120 ;
        RECT -3.220 3.030 -2.900 3.070 ;
        RECT -4.160 2.860 -3.970 2.870 ;
        RECT -3.220 2.840 -2.890 3.030 ;
        RECT -3.220 2.810 -2.900 2.840 ;
        RECT -3.800 2.690 -3.590 2.700 ;
        RECT -3.810 2.110 -3.590 2.690 ;
        RECT -3.800 2.080 -3.590 2.110 ;
        RECT -5.610 1.810 -5.080 1.980 ;
        RECT -3.800 1.730 -3.600 2.080 ;
        RECT -3.100 1.880 -2.920 2.810 ;
        RECT -2.290 2.540 -2.120 3.920 ;
        RECT -2.290 2.280 -1.810 2.540 ;
        RECT -2.290 2.140 -2.040 2.280 ;
        RECT -2.370 1.970 -2.040 2.140 ;
        RECT -1.540 1.870 -1.360 5.780 ;
        RECT -0.730 4.930 -0.560 6.310 ;
        RECT 0.100 6.240 0.710 6.500 ;
        RECT 0.100 6.210 0.270 6.240 ;
        RECT 0.510 6.200 0.710 6.240 ;
        RECT 1.100 6.200 1.650 7.190 ;
        RECT 2.470 7.040 3.100 7.210 ;
        RECT 2.470 6.940 2.860 7.040 ;
        RECT 2.470 6.910 2.850 6.940 ;
        RECT 2.470 6.760 2.830 6.910 ;
        RECT 2.120 6.590 2.830 6.760 ;
        RECT 2.120 5.840 2.820 6.150 ;
        RECT 0.100 5.650 0.270 5.680 ;
        RECT 0.510 5.650 0.710 5.690 ;
        RECT 0.100 5.390 0.710 5.650 ;
        RECT 0.100 5.350 0.270 5.390 ;
        RECT 0.510 5.360 0.710 5.390 ;
        RECT 0.510 5.000 0.710 5.030 ;
        RECT -0.930 4.730 -0.610 4.760 ;
        RECT 0.280 4.740 0.710 5.000 ;
        RECT -0.930 4.540 -0.600 4.730 ;
        RECT 0.510 4.700 0.710 4.740 ;
        RECT 1.100 4.700 1.650 5.690 ;
        RECT 1.970 5.610 2.820 5.840 ;
        RECT 2.120 5.270 2.820 5.610 ;
        RECT 2.580 4.910 2.900 4.950 ;
        RECT 2.580 4.850 2.910 4.910 ;
        RECT 2.110 4.720 2.910 4.850 ;
        RECT 2.110 4.690 2.900 4.720 ;
        RECT 2.110 4.670 2.810 4.690 ;
        RECT -0.930 4.500 -0.610 4.540 ;
        RECT -0.930 4.420 -0.760 4.500 ;
        RECT -0.980 4.250 -0.760 4.420 ;
        RECT -0.980 4.090 -0.810 4.250 ;
        RECT 2.570 4.190 2.890 4.230 ;
        RECT 0.510 4.150 0.710 4.190 ;
        RECT -0.450 3.830 -0.260 3.950 ;
        RECT 0.280 3.890 0.710 4.150 ;
        RECT 0.510 3.860 0.710 3.890 ;
        RECT -0.810 3.720 -0.260 3.830 ;
        RECT -0.810 3.660 -0.270 3.720 ;
        RECT -0.730 1.880 -0.560 3.660 ;
        RECT 0.100 3.500 0.270 3.540 ;
        RECT 0.510 3.500 0.710 3.530 ;
        RECT 0.100 3.240 0.710 3.500 ;
        RECT 0.100 3.210 0.270 3.240 ;
        RECT 0.510 3.200 0.710 3.240 ;
        RECT 1.100 3.200 1.650 4.190 ;
        RECT 2.110 4.010 2.900 4.190 ;
        RECT 2.570 4.000 2.900 4.010 ;
        RECT 2.570 3.970 2.890 4.000 ;
        RECT 2.120 3.250 2.820 3.590 ;
        RECT 1.970 3.020 2.820 3.250 ;
        RECT 2.120 2.710 2.820 3.020 ;
        RECT 0.100 2.650 0.270 2.680 ;
        RECT 0.510 2.650 0.710 2.690 ;
        RECT 0.100 2.390 0.710 2.650 ;
        RECT 0.100 2.350 0.270 2.390 ;
        RECT 0.510 2.360 0.710 2.390 ;
        RECT 0.510 2.000 0.710 2.030 ;
        RECT 0.280 1.740 0.710 2.000 ;
        RECT -2.520 1.710 -2.350 1.730 ;
        RECT -2.520 1.450 -1.960 1.710 ;
        RECT 0.510 1.700 0.710 1.740 ;
        RECT 1.100 1.700 1.650 2.690 ;
        RECT 2.120 2.100 2.830 2.270 ;
        RECT 2.470 1.820 2.830 2.100 ;
        RECT 2.470 1.650 3.100 1.820 ;
        RECT -2.520 1.400 -2.350 1.450 ;
      LAYER mcon ;
        RECT -0.630 7.180 -0.460 7.350 ;
        RECT -3.790 6.570 -3.620 6.740 ;
        RECT -10.630 5.990 -10.460 6.160 ;
        RECT -14.290 5.390 -14.020 5.660 ;
        RECT -10.630 5.540 -10.460 5.710 ;
        RECT -5.460 5.740 -5.290 5.910 ;
        RECT -4.150 5.730 -3.970 5.920 ;
        RECT -11.870 4.620 -11.700 4.790 ;
        RECT -11.870 4.280 -11.700 4.450 ;
        RECT -14.290 3.660 -14.020 3.930 ;
        RECT -11.870 3.930 -11.700 4.100 ;
        RECT -10.630 3.040 -10.460 3.210 ;
        RECT -5.460 2.980 -5.290 3.150 ;
        RECT -10.630 2.590 -10.460 2.760 ;
        RECT -4.150 2.930 -3.970 3.120 ;
        RECT 0.340 6.930 0.510 7.100 ;
        RECT 1.320 6.610 1.490 6.780 ;
        RECT 2.590 6.950 2.760 7.120 ;
        RECT -0.480 6.350 -0.310 6.520 ;
        RECT -1.600 5.830 -1.430 6.000 ;
        RECT -2.000 4.930 -1.830 5.100 ;
        RECT -2.430 4.130 -2.260 4.300 ;
        RECT -3.160 2.850 -2.990 3.020 ;
        RECT -3.790 2.110 -3.620 2.280 ;
        RECT -2.040 2.330 -1.870 2.500 ;
        RECT 0.290 6.280 0.460 6.450 ;
        RECT 0.290 5.440 0.460 5.610 ;
        RECT 1.980 5.640 2.150 5.810 ;
        RECT 1.320 5.110 1.490 5.280 ;
        RECT 0.340 4.790 0.510 4.960 ;
        RECT -0.870 4.550 -0.700 4.720 ;
        RECT 2.640 4.730 2.810 4.900 ;
        RECT -0.440 3.750 -0.270 3.920 ;
        RECT 0.340 3.930 0.510 4.100 ;
        RECT 2.630 4.010 2.800 4.180 ;
        RECT 1.320 3.610 1.490 3.780 ;
        RECT 0.290 3.280 0.460 3.450 ;
        RECT 1.980 3.050 2.150 3.220 ;
        RECT 0.290 2.440 0.460 2.610 ;
        RECT 1.320 2.110 1.490 2.280 ;
        RECT 0.340 1.790 0.510 1.960 ;
        RECT 2.550 1.760 2.720 1.930 ;
        RECT -2.190 1.500 -2.020 1.670 ;
      LAYER met1 ;
        RECT -11.900 4.880 -11.670 7.450 ;
        RECT -5.680 6.630 -5.370 7.070 ;
        RECT -3.720 6.800 -3.440 7.450 ;
        RECT -0.710 7.110 -0.390 7.430 ;
        RECT 0.270 6.860 0.590 7.180 ;
        RECT 2.520 6.880 2.840 7.200 ;
        RECT -3.830 6.200 -3.440 6.800 ;
        RECT -0.560 6.280 -0.240 6.600 ;
        RECT 0.220 6.210 0.540 6.530 ;
        RECT -5.530 5.670 -5.210 5.990 ;
        RECT -4.560 4.880 -4.320 5.010 ;
        RECT -11.940 3.870 -11.560 4.880 ;
        RECT -4.560 4.560 -4.300 4.880 ;
        RECT -3.720 4.600 -3.440 6.200 ;
        RECT -1.670 5.750 -1.350 6.070 ;
        RECT -0.450 5.590 -0.240 5.700 ;
        RECT -0.470 5.270 -0.210 5.590 ;
        RECT 0.220 5.360 0.540 5.680 ;
        RECT -2.030 4.870 -1.800 5.160 ;
        RECT -3.720 4.280 -3.360 4.600 ;
        RECT -4.560 3.960 -4.300 4.280 ;
        RECT -11.900 1.400 -11.670 3.870 ;
        RECT -4.560 3.840 -4.320 3.960 ;
        RECT -5.530 2.910 -5.210 3.230 ;
        RECT -3.720 2.650 -3.440 4.280 ;
        RECT -2.500 4.060 -2.180 4.380 ;
        RECT -2.010 3.580 -1.800 4.870 ;
        RECT -0.940 4.470 -0.620 4.790 ;
        RECT -0.450 3.980 -0.240 5.270 ;
        RECT 0.270 4.710 0.590 5.030 ;
        RECT 2.570 4.660 2.890 4.980 ;
        RECT -0.470 3.690 -0.240 3.980 ;
        RECT 0.270 3.860 0.590 4.180 ;
        RECT 2.560 3.940 2.880 4.260 ;
        RECT -2.030 3.260 -1.770 3.580 ;
        RECT -2.010 3.150 -1.800 3.260 ;
        RECT 0.220 3.210 0.540 3.530 ;
        RECT -3.230 2.780 -2.910 3.100 ;
        RECT -5.680 1.780 -5.370 2.220 ;
        RECT -3.830 2.050 -3.440 2.650 ;
        RECT -2.120 2.250 -1.800 2.570 ;
        RECT 0.220 2.360 0.540 2.680 ;
        RECT -3.720 1.400 -3.440 2.050 ;
        RECT -2.270 1.420 -1.950 1.740 ;
        RECT 0.270 1.710 0.590 2.030 ;
        RECT 2.480 1.690 2.800 2.010 ;
      LAYER via ;
        RECT -5.650 6.660 -5.390 6.920 ;
        RECT -0.680 7.140 -0.420 7.400 ;
        RECT 0.300 6.890 0.560 7.150 ;
        RECT 2.550 6.910 2.810 7.170 ;
        RECT -0.530 6.310 -0.270 6.570 ;
        RECT 0.250 6.240 0.510 6.500 ;
        RECT -5.500 5.700 -5.240 5.960 ;
        RECT -11.900 3.910 -11.610 4.840 ;
        RECT -4.560 4.590 -4.300 4.850 ;
        RECT -1.640 5.780 -1.380 6.040 ;
        RECT -0.470 5.300 -0.210 5.560 ;
        RECT 0.250 5.390 0.510 5.650 ;
        RECT -3.620 4.310 -3.360 4.570 ;
        RECT -4.560 3.990 -4.300 4.250 ;
        RECT -5.500 2.940 -5.240 3.200 ;
        RECT -2.470 4.090 -2.210 4.350 ;
        RECT -0.910 4.500 -0.650 4.760 ;
        RECT 0.300 4.740 0.560 5.000 ;
        RECT 2.600 4.690 2.860 4.950 ;
        RECT 0.300 3.890 0.560 4.150 ;
        RECT 2.590 3.970 2.850 4.230 ;
        RECT -2.030 3.290 -1.770 3.550 ;
        RECT 0.250 3.240 0.510 3.500 ;
        RECT -3.200 2.810 -2.940 3.070 ;
        RECT -5.650 1.930 -5.390 2.190 ;
        RECT -2.090 2.280 -1.830 2.540 ;
        RECT 0.250 2.390 0.510 2.650 ;
        RECT 0.300 1.740 0.560 2.000 ;
        RECT 2.510 1.720 2.770 1.980 ;
        RECT -2.240 1.450 -1.980 1.710 ;
      LAYER met2 ;
        RECT 0.270 7.110 0.580 7.190 ;
        RECT 2.520 7.110 2.830 7.210 ;
        RECT 0.270 6.880 2.830 7.110 ;
        RECT 0.270 6.860 0.580 6.880 ;
        RECT -0.550 6.570 -0.240 6.610 ;
        RECT -0.730 6.460 0.010 6.570 ;
        RECT 0.220 6.460 0.530 6.540 ;
        RECT -0.730 6.320 0.530 6.460 ;
        RECT -0.550 6.280 0.530 6.320 ;
        RECT -0.240 6.250 0.530 6.280 ;
        RECT -0.240 6.200 0.010 6.250 ;
        RECT 0.220 6.210 0.530 6.250 ;
        RECT -5.530 5.930 -5.220 6.000 ;
        RECT -1.670 5.930 -1.360 6.070 ;
        RECT -5.530 5.740 -1.360 5.930 ;
        RECT -5.530 5.710 -1.620 5.740 ;
        RECT -5.530 5.670 -5.220 5.710 ;
        RECT 0.220 5.640 0.530 5.680 ;
        RECT -0.210 5.560 0.530 5.640 ;
        RECT -0.500 5.540 0.530 5.560 ;
        RECT -0.550 5.430 0.530 5.540 ;
        RECT -0.550 5.350 0.000 5.430 ;
        RECT 0.220 5.350 0.530 5.430 ;
        RECT -0.550 5.290 -0.080 5.350 ;
        RECT -2.110 3.470 -1.640 3.560 ;
        RECT -2.110 3.460 0.000 3.470 ;
        RECT 0.220 3.460 0.530 3.540 ;
        RECT -2.110 3.310 0.530 3.460 ;
        RECT -2.060 3.290 0.530 3.310 ;
        RECT -1.770 3.270 0.530 3.290 ;
        RECT -0.080 3.250 0.530 3.270 ;
        RECT -5.530 3.170 -5.220 3.240 ;
        RECT 0.220 3.210 0.530 3.250 ;
        RECT -3.340 3.170 -3.180 3.180 ;
        RECT -5.530 3.110 -3.180 3.170 ;
        RECT -5.530 2.960 -2.920 3.110 ;
        RECT -5.530 2.910 -5.220 2.960 ;
        RECT -3.340 2.780 -2.920 2.960 ;
        RECT -2.060 2.640 0.000 2.670 ;
        RECT 0.220 2.640 0.530 2.680 ;
        RECT -2.060 2.570 0.530 2.640 ;
        RECT -2.110 2.530 0.530 2.570 ;
        RECT -2.290 2.460 0.530 2.530 ;
        RECT -2.290 2.280 -1.740 2.460 ;
        RECT -0.080 2.430 0.530 2.460 ;
        RECT 0.220 2.350 0.530 2.430 ;
        RECT -2.110 2.240 -1.800 2.280 ;
        RECT 0.270 1.980 0.580 2.030 ;
        RECT 2.480 1.980 2.790 2.020 ;
        RECT 0.270 1.750 2.980 1.980 ;
        RECT 0.270 1.700 0.580 1.750 ;
        RECT 2.480 1.690 2.790 1.750 ;
  END
END sky130_hilas_TA2Cell_NoFG

MACRO sky130_hilas_pFETLarge
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pFETLarge ;
  ORIGIN -0.640 -4.190 ;
  SIZE 4.640 BY 5.990 ;
  PIN GATE
    ANTENNAGATEAREA 6.526000 ;
    PORT
      LAYER met2 ;
        RECT 0.640 4.530 1.240 5.020 ;
        RECT 0.640 4.200 1.250 4.530 ;
    END
  END GATE
  PIN SOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 4.367400 ;
    PORT
      LAYER met2 ;
        RECT 0.970 9.790 4.030 9.800 ;
        RECT 0.880 9.460 4.030 9.790 ;
        RECT 0.880 7.010 1.200 9.460 ;
        RECT 3.700 9.450 4.010 9.460 ;
        RECT 0.880 6.680 4.040 7.010 ;
        RECT 0.880 5.640 1.200 6.680 ;
        RECT 0.880 5.320 4.040 5.640 ;
        RECT 1.500 5.310 1.810 5.320 ;
        RECT 2.600 5.310 2.910 5.320 ;
        RECT 3.700 5.310 4.010 5.320 ;
    END
  END SOURCE
  PIN DRAIN
    USE ANALOG ;
    ANTENNADIFFAREA 4.317200 ;
    PORT
      LAYER met2 ;
        RECT 2.060 9.080 2.370 9.110 ;
        RECT 3.150 9.080 3.460 9.090 ;
        RECT 2.060 8.780 5.010 9.080 ;
        RECT 3.150 8.760 3.460 8.780 ;
        RECT 4.260 8.740 5.010 8.780 ;
        RECT 4.630 8.610 5.010 8.740 ;
        RECT 4.660 7.740 5.010 8.610 ;
        RECT 2.060 7.410 5.010 7.740 ;
        RECT 4.660 4.970 5.010 7.410 ;
        RECT 2.070 4.960 5.010 4.970 ;
        RECT 2.060 4.650 5.010 4.960 ;
        RECT 2.060 4.640 4.780 4.650 ;
        RECT 2.060 4.630 2.370 4.640 ;
        RECT 3.150 4.630 3.460 4.640 ;
    END
  END DRAIN
  PIN WELL
    USE ANALOG ;
    ANTENNADIFFAREA 0.213200 ;
    PORT
      LAYER nwell ;
        RECT 1.360 4.370 5.280 10.070 ;
      LAYER met1 ;
        RECT 4.780 9.980 5.040 10.180 ;
        RECT 4.780 9.170 5.090 9.980 ;
        RECT 4.780 4.190 5.040 9.170 ;
    END
  END WELL
  OBS
      LAYER li1 ;
        RECT 1.600 9.750 1.770 9.840 ;
        RECT 1.520 9.710 1.840 9.750 ;
        RECT 1.520 9.520 1.850 9.710 ;
        RECT 1.520 9.490 1.840 9.520 ;
        RECT 1.600 6.970 1.770 9.490 ;
        RECT 2.150 9.070 2.320 9.840 ;
        RECT 2.700 9.750 2.870 9.840 ;
        RECT 2.610 9.710 2.930 9.750 ;
        RECT 2.610 9.520 2.940 9.710 ;
        RECT 2.610 9.490 2.930 9.520 ;
        RECT 2.070 9.030 2.390 9.070 ;
        RECT 2.070 8.840 2.400 9.030 ;
        RECT 2.070 8.810 2.390 8.840 ;
        RECT 2.150 7.700 2.320 8.810 ;
        RECT 2.070 7.660 2.390 7.700 ;
        RECT 2.070 7.470 2.400 7.660 ;
        RECT 2.070 7.440 2.390 7.470 ;
        RECT 1.510 6.930 1.830 6.970 ;
        RECT 1.510 6.740 1.840 6.930 ;
        RECT 1.510 6.710 1.830 6.740 ;
        RECT 1.600 5.600 1.770 6.710 ;
        RECT 1.510 5.560 1.830 5.600 ;
        RECT 1.510 5.370 1.840 5.560 ;
        RECT 1.510 5.340 1.830 5.370 ;
        RECT 0.830 5.130 1.340 5.210 ;
        RECT 0.830 4.880 1.350 5.130 ;
        RECT 0.840 4.200 1.350 4.880 ;
        RECT 1.600 4.520 1.770 5.340 ;
        RECT 2.150 4.920 2.320 7.440 ;
        RECT 2.700 6.970 2.870 9.490 ;
        RECT 3.250 9.050 3.420 9.840 ;
        RECT 3.800 9.740 3.970 9.840 ;
        RECT 3.710 9.700 4.030 9.740 ;
        RECT 3.710 9.510 4.040 9.700 ;
        RECT 3.710 9.480 4.030 9.510 ;
        RECT 3.160 9.010 3.480 9.050 ;
        RECT 3.160 8.820 3.490 9.010 ;
        RECT 3.160 8.790 3.480 8.820 ;
        RECT 3.250 7.700 3.420 8.790 ;
        RECT 3.160 7.660 3.480 7.700 ;
        RECT 3.160 7.470 3.490 7.660 ;
        RECT 3.160 7.440 3.480 7.470 ;
        RECT 2.610 6.930 2.930 6.970 ;
        RECT 2.610 6.740 2.940 6.930 ;
        RECT 2.610 6.710 2.930 6.740 ;
        RECT 2.700 5.600 2.870 6.710 ;
        RECT 2.610 5.560 2.930 5.600 ;
        RECT 2.610 5.370 2.940 5.560 ;
        RECT 2.610 5.340 2.930 5.370 ;
        RECT 2.070 4.880 2.390 4.920 ;
        RECT 2.070 4.690 2.400 4.880 ;
        RECT 2.070 4.660 2.390 4.690 ;
        RECT 2.150 4.510 2.320 4.660 ;
        RECT 2.700 4.510 2.870 5.340 ;
        RECT 3.250 4.920 3.420 7.440 ;
        RECT 3.800 6.970 3.970 9.480 ;
        RECT 4.350 9.040 4.520 9.840 ;
        RECT 4.890 9.110 5.060 9.870 ;
        RECT 4.270 9.000 4.590 9.040 ;
        RECT 4.270 8.810 4.600 9.000 ;
        RECT 4.270 8.780 4.590 8.810 ;
        RECT 4.350 7.700 4.520 8.780 ;
        RECT 4.260 7.660 4.580 7.700 ;
        RECT 4.260 7.470 4.590 7.660 ;
        RECT 4.260 7.440 4.580 7.470 ;
        RECT 3.710 6.930 4.030 6.970 ;
        RECT 3.710 6.740 4.040 6.930 ;
        RECT 3.710 6.710 4.030 6.740 ;
        RECT 3.800 5.600 3.970 6.710 ;
        RECT 3.710 5.560 4.030 5.600 ;
        RECT 3.710 5.370 4.040 5.560 ;
        RECT 3.710 5.340 4.030 5.370 ;
        RECT 3.160 4.880 3.480 4.920 ;
        RECT 3.160 4.690 3.490 4.880 ;
        RECT 3.160 4.660 3.480 4.690 ;
        RECT 3.250 4.510 3.420 4.660 ;
        RECT 3.800 4.510 3.970 5.340 ;
        RECT 4.350 4.930 4.520 7.440 ;
        RECT 4.260 4.890 4.580 4.930 ;
        RECT 4.260 4.700 4.590 4.890 ;
        RECT 4.260 4.670 4.580 4.700 ;
        RECT 4.350 4.510 4.520 4.670 ;
      LAYER mcon ;
        RECT 1.580 9.530 1.750 9.700 ;
        RECT 2.670 9.530 2.840 9.700 ;
        RECT 2.130 8.850 2.300 9.020 ;
        RECT 2.130 7.480 2.300 7.650 ;
        RECT 1.570 6.750 1.740 6.920 ;
        RECT 1.570 5.380 1.740 5.550 ;
        RECT 1.000 4.740 1.170 4.910 ;
        RECT 3.770 9.520 3.940 9.690 ;
        RECT 3.220 8.830 3.390 9.000 ;
        RECT 3.220 7.480 3.390 7.650 ;
        RECT 2.670 6.750 2.840 6.920 ;
        RECT 2.670 5.380 2.840 5.550 ;
        RECT 2.130 4.700 2.300 4.870 ;
        RECT 4.890 9.700 5.060 9.870 ;
        RECT 4.890 9.340 5.060 9.510 ;
        RECT 4.330 8.820 4.500 8.990 ;
        RECT 4.320 7.480 4.490 7.650 ;
        RECT 3.770 6.750 3.940 6.920 ;
        RECT 3.770 5.380 3.940 5.550 ;
        RECT 3.220 4.700 3.390 4.870 ;
        RECT 4.320 4.710 4.490 4.880 ;
        RECT 1.010 4.270 1.180 4.440 ;
      LAYER met1 ;
        RECT 1.510 9.460 1.830 9.780 ;
        RECT 2.600 9.460 2.920 9.780 ;
        RECT 3.700 9.450 4.020 9.770 ;
        RECT 2.060 8.780 2.380 9.100 ;
        RECT 3.150 8.760 3.470 9.080 ;
        RECT 4.260 8.750 4.580 9.070 ;
        RECT 2.060 7.410 2.380 7.730 ;
        RECT 3.150 7.410 3.470 7.730 ;
        RECT 4.250 7.410 4.570 7.730 ;
        RECT 1.500 6.680 1.820 7.000 ;
        RECT 2.600 6.680 2.920 7.000 ;
        RECT 3.700 6.680 4.020 7.000 ;
        RECT 1.500 5.310 1.820 5.630 ;
        RECT 2.600 5.310 2.920 5.630 ;
        RECT 3.700 5.310 4.020 5.630 ;
        RECT 0.930 4.670 1.250 4.990 ;
        RECT 2.060 4.630 2.380 4.950 ;
        RECT 3.150 4.630 3.470 4.950 ;
        RECT 4.250 4.640 4.570 4.960 ;
        RECT 0.940 4.200 1.260 4.520 ;
      LAYER via ;
        RECT 1.540 9.490 1.800 9.750 ;
        RECT 2.630 9.490 2.890 9.750 ;
        RECT 3.730 9.480 3.990 9.740 ;
        RECT 2.090 8.810 2.350 9.070 ;
        RECT 3.180 8.790 3.440 9.050 ;
        RECT 4.290 8.780 4.550 9.040 ;
        RECT 2.090 7.440 2.350 7.700 ;
        RECT 3.180 7.440 3.440 7.700 ;
        RECT 4.280 7.440 4.540 7.700 ;
        RECT 1.530 6.710 1.790 6.970 ;
        RECT 2.630 6.710 2.890 6.970 ;
        RECT 3.730 6.710 3.990 6.970 ;
        RECT 1.530 5.340 1.790 5.600 ;
        RECT 2.630 5.340 2.890 5.600 ;
        RECT 3.730 5.340 3.990 5.600 ;
        RECT 0.960 4.700 1.220 4.960 ;
        RECT 2.090 4.660 2.350 4.920 ;
        RECT 3.180 4.660 3.440 4.920 ;
        RECT 4.280 4.670 4.540 4.930 ;
        RECT 0.970 4.230 1.230 4.490 ;
  END
END sky130_hilas_pFETLarge

MACRO sky130_hilas_VinjInv2
  CLASS BLOCK ;
  FOREIGN sky130_hilas_VinjInv2 ;
  ORIGIN 3.360 -1.440 ;
  SIZE 3.610 BY 1.640 ;
  OBS
      LAYER nwell ;
        RECT -3.360 1.440 -1.380 3.080 ;
      LAYER li1 ;
        RECT -2.740 2.650 -2.570 2.790 ;
        RECT -2.740 2.480 -2.550 2.650 ;
        RECT -2.740 2.380 -2.570 2.480 ;
        RECT -3.170 2.000 -3.000 2.100 ;
        RECT -3.190 1.830 -3.000 2.000 ;
        RECT -3.170 1.770 -3.000 1.830 ;
        RECT -2.750 2.040 -2.580 2.100 ;
        RECT -2.750 1.770 -2.500 2.040 ;
        RECT -2.010 2.020 -1.760 2.100 ;
        RECT -2.010 1.850 -0.710 2.020 ;
        RECT -0.150 2.010 0.020 2.640 ;
        RECT -2.740 1.750 -2.500 1.770 ;
        RECT -1.930 1.760 -1.760 1.850 ;
        RECT -0.230 1.840 0.100 2.010 ;
      LAYER mcon ;
        RECT -2.720 2.480 -2.550 2.650 ;
        RECT -0.150 2.120 0.020 2.290 ;
        RECT -2.710 1.800 -2.540 1.970 ;
        RECT -1.370 1.850 -1.200 2.020 ;
      LAYER met1 ;
        RECT -2.750 2.700 -2.530 3.040 ;
        RECT -2.750 2.440 -2.520 2.700 ;
        RECT -3.280 1.760 -2.970 2.110 ;
        RECT -2.750 2.040 -2.530 2.440 ;
        RECT -2.750 1.730 -2.500 2.040 ;
        RECT -1.450 1.800 -1.130 2.060 ;
        RECT -2.750 1.530 -2.530 1.730 ;
        RECT -0.180 1.530 0.050 3.040 ;
      LAYER via ;
        RECT -3.250 1.790 -2.990 2.050 ;
        RECT -1.420 1.800 -1.160 2.060 ;
      LAYER met2 ;
        RECT -3.360 2.470 0.250 2.650 ;
        RECT -3.280 1.950 -2.960 2.050 ;
        RECT -3.290 1.790 -2.960 1.950 ;
        RECT -1.450 1.980 -1.130 2.060 ;
        RECT -1.450 1.800 0.250 1.980 ;
  END
END sky130_hilas_VinjInv2

MACRO sky130_hilas_capacitorSize03
  CLASS BLOCK ;
  FOREIGN sky130_hilas_capacitorSize03 ;
  ORIGIN -14.140 0.470 ;
  SIZE 5.790 BY 5.870 ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 19.100 2.160 19.760 2.820 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 16.710 4.060 17.160 4.070 ;
        RECT 16.690 3.570 17.210 4.060 ;
        RECT 14.250 2.720 14.910 2.780 ;
        RECT 16.720 2.730 17.160 3.570 ;
        RECT 15.300 2.720 16.310 2.730 ;
        RECT 16.710 2.720 17.170 2.730 ;
        RECT 14.250 2.220 17.170 2.720 ;
        RECT 14.250 2.210 15.660 2.220 ;
        RECT 14.250 2.120 14.910 2.210 ;
        RECT 16.710 1.560 17.170 2.220 ;
        RECT 16.710 1.050 17.190 1.560 ;
        RECT 16.690 0.560 17.210 1.050 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 14.140 4.800 19.920 4.980 ;
        RECT 14.140 4.370 19.920 4.550 ;
        RECT 14.170 3.370 19.920 3.550 ;
        RECT 14.170 2.940 19.920 3.120 ;
        RECT 14.380 2.600 14.750 2.660 ;
        RECT 14.160 2.320 14.750 2.600 ;
        RECT 14.380 2.260 14.750 2.320 ;
        RECT 19.230 2.640 19.600 2.700 ;
        RECT 19.230 2.360 19.930 2.640 ;
        RECT 19.230 2.300 19.600 2.360 ;
        RECT 14.170 1.790 19.920 1.960 ;
        RECT 14.170 1.370 19.920 1.540 ;
        RECT 14.170 0.390 19.920 0.560 ;
        RECT 14.170 -0.050 19.920 0.120 ;
      LAYER via2 ;
        RECT 14.430 2.320 14.710 2.600 ;
        RECT 19.280 2.360 19.560 2.640 ;
      LAYER met3 ;
        RECT 15.590 2.850 18.430 5.400 ;
        RECT 14.160 2.060 14.950 2.810 ;
        RECT 15.590 2.100 19.800 2.850 ;
        RECT 15.590 -0.470 18.430 2.100 ;
      LAYER via3 ;
        RECT 14.350 2.210 14.780 2.690 ;
        RECT 19.200 2.250 19.630 2.730 ;
  END
END sky130_hilas_capacitorSize03

MACRO sky130_hilas_swc4x1BiasCell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc4x1BiasCell ;
  ORIGIN 2.640 4.000 ;
  SIZE 10.080 BY 6.500 ;
  PIN ROW1
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 4.970 1.510 5.280 1.530 ;
        RECT -2.630 1.330 7.440 1.510 ;
        RECT -2.630 1.320 5.280 1.330 ;
        RECT 4.970 1.200 5.280 1.320 ;
    END
  END ROW1
  PIN ROW2
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 4.970 0.420 5.280 0.550 ;
        RECT -2.630 0.240 7.440 0.420 ;
        RECT 4.970 0.220 5.280 0.240 ;
    END
  END ROW2
  PIN ROW3
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -2.630 -1.870 -2.160 -1.710 ;
        RECT -2.620 -1.880 -2.160 -1.870 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.970 -1.730 5.280 -1.710 ;
        RECT -1.860 -1.900 7.440 -1.730 ;
        RECT 4.880 -1.910 7.440 -1.900 ;
        RECT 4.970 -2.040 5.280 -1.910 ;
    END
  END ROW3
  PIN ROW4
    USE ANALOG ;
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT -2.630 -2.700 5.000 -2.690 ;
        RECT -2.630 -2.830 5.280 -2.700 ;
        RECT -2.630 -2.860 7.440 -2.830 ;
        RECT 4.880 -3.010 7.440 -2.860 ;
        RECT 4.970 -3.030 5.280 -3.010 ;
    END
  END ROW4
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 2.243500 ;
    PORT
      LAYER nwell ;
        RECT -2.630 -4.000 -0.900 2.500 ;
      LAYER met1 ;
        RECT -2.280 -4.000 -1.880 2.500 ;
    END
  END VTUN
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 3.253900 ;
    PORT
      LAYER nwell ;
        RECT 1.120 -4.000 3.350 2.490 ;
      LAYER met1 ;
        RECT 1.770 0.310 2.150 2.500 ;
        RECT 1.760 -1.550 2.150 0.310 ;
        RECT 1.770 -4.000 2.150 -1.550 ;
    END
  END GATE1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 4.880 -4.000 7.440 2.500 ;
      LAYER met1 ;
        RECT 6.920 1.790 7.080 2.490 ;
        RECT 6.810 1.240 7.080 1.790 ;
        RECT 6.810 1.190 7.090 1.240 ;
        RECT 6.920 1.100 7.090 1.190 ;
        RECT 6.920 0.650 7.080 1.100 ;
        RECT 6.920 0.560 7.090 0.650 ;
        RECT 6.810 0.510 7.090 0.560 ;
        RECT 6.810 -0.040 7.080 0.510 ;
        RECT 6.920 -1.450 7.080 -0.040 ;
        RECT 6.810 -2.000 7.080 -1.450 ;
        RECT 6.810 -2.050 7.090 -2.000 ;
        RECT 6.920 -2.140 7.090 -2.050 ;
        RECT 6.920 -2.600 7.080 -2.140 ;
        RECT 6.920 -2.690 7.090 -2.600 ;
        RECT 6.810 -2.740 7.090 -2.690 ;
        RECT 6.810 -3.290 7.080 -2.740 ;
        RECT 6.920 -3.990 7.080 -3.290 ;
    END
  END VINJ
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 6.110 1.760 6.270 2.490 ;
        RECT 6.110 1.740 6.310 1.760 ;
        RECT 6.090 1.500 6.320 1.740 ;
        RECT 6.110 1.450 6.320 1.500 ;
        RECT 6.480 1.450 6.670 2.440 ;
        RECT 6.110 0.300 6.270 1.450 ;
        RECT 6.500 1.330 6.670 1.450 ;
        RECT 6.510 0.420 6.670 1.330 ;
        RECT 6.500 0.300 6.670 0.420 ;
        RECT 6.110 0.250 6.320 0.300 ;
        RECT 6.090 0.010 6.320 0.250 ;
        RECT 6.110 -0.010 6.310 0.010 ;
        RECT 6.110 -0.650 6.270 -0.010 ;
        RECT 6.480 -0.620 6.670 0.300 ;
        RECT 6.460 -0.650 6.700 -0.620 ;
        RECT 6.110 -0.820 6.700 -0.650 ;
        RECT 6.110 -1.480 6.270 -0.820 ;
        RECT 6.460 -0.850 6.700 -0.820 ;
        RECT 6.110 -1.500 6.310 -1.480 ;
        RECT 6.090 -1.740 6.320 -1.500 ;
        RECT 6.110 -1.790 6.320 -1.740 ;
        RECT 6.480 -1.790 6.670 -0.850 ;
        RECT 6.110 -2.950 6.270 -1.790 ;
        RECT 6.500 -1.910 6.670 -1.790 ;
        RECT 6.510 -2.830 6.670 -1.910 ;
        RECT 6.500 -2.950 6.670 -2.830 ;
        RECT 6.110 -3.000 6.320 -2.950 ;
        RECT 6.090 -3.240 6.320 -3.000 ;
        RECT 6.110 -3.260 6.310 -3.240 ;
        RECT 6.110 -3.990 6.270 -3.260 ;
        RECT 6.480 -3.940 6.670 -2.950 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT -0.100 -2.300 0.230 -2.270 ;
        RECT 3.930 -2.300 4.250 -2.240 ;
        RECT -0.100 -2.470 4.250 -2.300 ;
        RECT -0.100 -2.530 0.230 -2.470 ;
        RECT 3.930 -2.520 4.250 -2.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.960 -2.210 4.210 2.500 ;
        RECT 3.950 -2.240 4.230 -2.210 ;
        RECT 3.940 -2.520 4.240 -2.240 ;
        RECT 3.950 -2.540 4.230 -2.520 ;
        RECT 3.960 -4.000 4.210 -2.540 ;
      LAYER via ;
        RECT 3.960 -2.510 4.220 -2.250 ;
    END
    PORT
      LAYER met1 ;
        RECT -0.070 -2.240 0.200 2.500 ;
        RECT -0.090 -2.550 0.220 -2.240 ;
        RECT -0.070 -4.000 0.200 -2.550 ;
      LAYER via ;
        RECT -0.070 -2.530 0.200 -2.270 ;
    END
  END VGND
  PIN DRAIN3
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 4.970 -1.290 5.280 -1.160 ;
        RECT 4.850 -1.300 5.280 -1.290 ;
        RECT 4.850 -1.460 7.440 -1.300 ;
        RECT 4.970 -1.480 7.440 -1.460 ;
        RECT 4.970 -1.490 5.280 -1.480 ;
    END
  END DRAIN3
  PIN DRAIN4
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 4.970 -3.260 5.280 -3.250 ;
        RECT 4.970 -3.440 7.440 -3.260 ;
        RECT 4.970 -3.580 5.280 -3.440 ;
    END
  END DRAIN4
  PIN DRAIN1
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 4.970 1.940 5.280 2.080 ;
        RECT 4.970 1.760 7.440 1.940 ;
        RECT 4.970 1.750 5.280 1.760 ;
    END
  END DRAIN1
  PIN DRAIN2
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 4.970 -0.010 5.280 0.000 ;
        RECT 4.970 -0.170 7.440 -0.010 ;
        RECT 4.880 -0.190 7.440 -0.170 ;
        RECT 4.880 -0.310 5.280 -0.190 ;
        RECT 4.970 -0.330 5.280 -0.310 ;
    END
  END DRAIN2
  OBS
      LAYER li1 ;
        RECT 4.980 2.030 5.300 2.040 ;
        RECT 4.980 1.860 5.560 2.030 ;
        RECT 4.980 1.810 5.310 1.860 ;
        RECT 4.980 1.780 5.300 1.810 ;
        RECT 6.840 1.760 7.040 2.110 ;
        RECT 4.980 1.450 5.300 1.490 ;
        RECT 4.980 1.410 5.310 1.450 ;
        RECT 4.980 1.240 5.560 1.410 ;
        RECT 4.980 1.230 5.300 1.240 ;
        RECT 6.110 1.140 6.310 1.740 ;
        RECT 6.840 1.730 7.050 1.760 ;
        RECT 6.830 1.140 7.050 1.730 ;
        RECT -0.020 0.480 0.150 1.010 ;
        RECT 4.000 0.450 4.170 0.980 ;
        RECT 4.980 0.510 5.300 0.520 ;
        RECT 4.980 0.340 5.560 0.510 ;
        RECT 4.980 0.300 5.310 0.340 ;
        RECT 4.980 0.260 5.300 0.300 ;
        RECT 6.110 0.010 6.310 0.610 ;
        RECT 6.830 0.020 7.050 0.610 ;
        RECT 6.840 -0.010 7.050 0.020 ;
        RECT 4.980 -0.060 5.300 -0.030 ;
        RECT 4.980 -0.110 5.310 -0.060 ;
        RECT -2.210 -1.020 -1.660 -0.590 ;
        RECT -0.010 -1.450 0.160 -0.280 ;
        RECT 1.820 -1.090 2.370 -0.660 ;
        RECT 4.010 -1.410 4.180 -0.220 ;
        RECT 4.980 -0.280 5.560 -0.110 ;
        RECT 4.980 -0.290 5.300 -0.280 ;
        RECT 6.840 -0.360 7.040 -0.010 ;
        RECT 6.230 -0.820 6.670 -0.650 ;
        RECT 4.980 -1.210 5.300 -1.200 ;
        RECT 4.980 -1.380 5.560 -1.210 ;
        RECT 4.980 -1.430 5.310 -1.380 ;
        RECT 4.980 -1.460 5.300 -1.430 ;
        RECT 6.840 -1.480 7.040 -1.130 ;
        RECT 4.980 -1.790 5.300 -1.750 ;
        RECT 4.980 -1.830 5.310 -1.790 ;
        RECT 4.980 -2.000 5.560 -1.830 ;
        RECT 4.980 -2.010 5.300 -2.000 ;
        RECT 6.110 -2.100 6.310 -1.500 ;
        RECT 6.840 -1.510 7.050 -1.480 ;
        RECT 6.830 -2.100 7.050 -1.510 ;
        RECT 4.980 -2.740 5.300 -2.730 ;
        RECT 4.980 -2.910 5.560 -2.740 ;
        RECT 4.980 -2.950 5.310 -2.910 ;
        RECT 4.980 -2.990 5.300 -2.950 ;
        RECT 6.110 -3.240 6.310 -2.640 ;
        RECT 6.830 -3.230 7.050 -2.640 ;
        RECT 6.840 -3.260 7.050 -3.230 ;
        RECT 4.980 -3.310 5.300 -3.280 ;
        RECT 4.980 -3.360 5.310 -3.310 ;
        RECT 4.980 -3.530 5.560 -3.360 ;
        RECT 4.980 -3.540 5.300 -3.530 ;
        RECT 6.840 -3.610 7.040 -3.260 ;
      LAYER mcon ;
        RECT 5.040 1.820 5.210 1.990 ;
        RECT 6.120 1.530 6.290 1.700 ;
        RECT 5.040 1.270 5.210 1.440 ;
        RECT 6.850 1.560 7.020 1.730 ;
        RECT -0.020 0.840 0.150 1.010 ;
        RECT 4.000 0.810 4.170 0.980 ;
        RECT 5.040 0.310 5.210 0.480 ;
        RECT 6.120 0.050 6.290 0.220 ;
        RECT 6.850 0.020 7.020 0.190 ;
        RECT -0.010 -0.450 0.160 -0.280 ;
        RECT -2.210 -0.940 -1.940 -0.670 ;
        RECT 4.010 -0.390 4.180 -0.220 ;
        RECT 5.040 -0.240 5.210 -0.070 ;
        RECT -0.010 -1.090 0.160 -0.920 ;
        RECT 1.820 -1.010 2.090 -0.740 ;
        RECT 6.490 -0.820 6.670 -0.650 ;
        RECT 4.010 -1.050 4.180 -0.880 ;
        RECT 5.040 -1.420 5.210 -1.250 ;
        RECT 6.120 -1.710 6.290 -1.540 ;
        RECT 5.040 -1.970 5.210 -1.800 ;
        RECT 6.850 -1.680 7.020 -1.510 ;
        RECT 5.040 -2.940 5.210 -2.770 ;
        RECT 6.120 -3.200 6.290 -3.030 ;
        RECT 6.850 -3.230 7.020 -3.060 ;
        RECT 5.040 -3.490 5.210 -3.320 ;
      LAYER met1 ;
        RECT 4.970 1.750 5.290 2.070 ;
        RECT 4.970 1.200 5.290 1.520 ;
        RECT 4.970 0.230 5.290 0.550 ;
        RECT 4.970 -0.320 5.290 0.000 ;
        RECT 4.970 -1.490 5.290 -1.170 ;
        RECT 4.970 -2.040 5.290 -1.720 ;
        RECT 4.970 -3.020 5.290 -2.700 ;
        RECT 4.970 -3.570 5.290 -3.250 ;
      LAYER via ;
        RECT 5.000 1.780 5.260 2.040 ;
        RECT 5.000 1.230 5.260 1.490 ;
        RECT 5.000 0.260 5.260 0.520 ;
        RECT 5.000 -0.290 5.260 -0.030 ;
        RECT 5.000 -1.460 5.260 -1.200 ;
        RECT 5.000 -2.010 5.260 -1.750 ;
        RECT 5.000 -2.990 5.260 -2.730 ;
        RECT 5.000 -3.540 5.260 -3.280 ;
  END
END sky130_hilas_swc4x1BiasCell

MACRO sky130_hilas_FGtrans2x1cell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_FGtrans2x1cell ;
  ORIGIN 3.950 3.870 ;
  SIZE 11.520 BY 6.150 ;
  PIN COLSEL1
    USE ANALOG ;
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT 6.610 0.770 6.800 2.230 ;
        RECT 6.610 0.740 6.830 0.770 ;
        RECT 6.590 0.470 6.840 0.740 ;
        RECT 6.600 0.460 6.840 0.470 ;
        RECT 6.600 0.220 6.830 0.460 ;
        RECT 6.640 -1.810 6.800 0.220 ;
        RECT 6.600 -2.050 6.830 -1.810 ;
        RECT 6.600 -2.060 6.840 -2.050 ;
        RECT 6.590 -2.330 6.840 -2.060 ;
        RECT 6.610 -2.360 6.830 -2.330 ;
        RECT 6.610 -3.820 6.800 -2.360 ;
    END
  END COLSEL1
  PIN VINJ
    USE ANALOG ;
    ANTENNADIFFAREA 0.544000 ;
    PORT
      LAYER nwell ;
        RECT 4.260 -3.870 7.570 2.280 ;
      LAYER met1 ;
        RECT 7.050 1.580 7.210 2.230 ;
        RECT 6.940 1.030 7.210 1.580 ;
        RECT 6.940 0.980 7.220 1.030 ;
        RECT 7.050 0.890 7.220 0.980 ;
        RECT 7.050 -2.480 7.210 0.890 ;
        RECT 7.050 -2.570 7.220 -2.480 ;
        RECT 6.940 -2.620 7.220 -2.570 ;
        RECT 6.940 -3.170 7.210 -2.620 ;
        RECT 7.050 -3.820 7.210 -3.170 ;
    END
  END VINJ
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 4.840 1.740 5.160 1.750 ;
        RECT 4.840 1.730 5.400 1.740 ;
        RECT -3.950 1.550 7.570 1.730 ;
        RECT 5.090 1.410 5.400 1.550 ;
    END
  END DRAIN1
  PIN DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 5.090 -3.140 5.400 -3.000 ;
        RECT 5.090 -3.150 7.570 -3.140 ;
        RECT -3.950 -3.300 7.570 -3.150 ;
        RECT 5.090 -3.320 7.570 -3.300 ;
        RECT 5.090 -3.330 5.400 -3.320 ;
    END
  END DRAIN2
  PIN PROG
    USE ANALOG ;
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER met1 ;
        RECT 3.840 -0.490 4.050 2.230 ;
        RECT 3.840 -1.000 4.080 -0.490 ;
        RECT 3.840 -3.820 4.050 -1.000 ;
    END
  END PROG
  PIN RUN
    USE ANALOG ;
    ANTENNAGATEAREA 0.790000 ;
    PORT
      LAYER met1 ;
        RECT 2.790 -2.300 2.970 2.230 ;
        RECT 2.740 -2.640 3.030 -2.300 ;
        RECT 2.790 -3.820 2.970 -2.640 ;
    END
  END RUN
  PIN VIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.217200 ;
    PORT
      LAYER met1 ;
        RECT 4.720 -1.200 4.910 -1.070 ;
        RECT 4.700 -1.490 4.930 -1.200 ;
        RECT 4.720 -3.110 4.910 -1.490 ;
        RECT 4.680 -3.320 4.910 -3.110 ;
        RECT 4.680 -3.400 4.920 -3.320 ;
        RECT 4.690 -3.820 4.920 -3.400 ;
    END
  END VIN2
  PIN VIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.217200 ;
    PORT
      LAYER met1 ;
        RECT 4.720 1.860 4.930 2.230 ;
        RECT 4.710 1.570 4.940 1.860 ;
        RECT 4.720 -0.130 4.930 1.570 ;
        RECT 4.710 -0.420 4.940 -0.130 ;
        RECT 4.720 -0.560 4.930 -0.420 ;
    END
  END VIN1
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 0.434600 ;
    PORT
      LAYER met1 ;
        RECT 4.270 1.300 4.460 2.230 ;
        RECT 4.240 1.010 4.470 1.300 ;
        RECT 4.270 -1.020 4.460 1.010 ;
        RECT 4.240 -1.310 4.470 -1.020 ;
        RECT 4.270 -2.600 4.460 -1.310 ;
        RECT 4.250 -2.890 4.480 -2.600 ;
        RECT 4.270 -3.820 4.460 -2.890 ;
    END
  END GATE1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT -1.130 -3.820 -0.900 2.230 ;
    END
  END VGND
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 2.516100 ;
    PORT
      LAYER nwell ;
        RECT -3.950 1.480 -2.220 2.230 ;
        RECT -3.950 0.330 -2.210 1.480 ;
        RECT -3.940 -1.910 -2.210 0.330 ;
        RECT -3.950 -2.090 -2.210 -1.910 ;
        RECT -3.950 -3.810 -2.220 -2.090 ;
      LAYER met1 ;
        RECT -3.610 -3.820 -3.190 2.230 ;
    END
  END VTUN
  PIN COL1
    ANTENNADIFFAREA 1.030400 ;
    PORT
      LAYER met2 ;
        RECT 6.190 -0.690 6.510 -0.660 ;
        RECT -3.950 -0.920 6.510 -0.690 ;
    END
  END COL1
  PIN ROW1
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 5.480 0.190 5.790 0.210 ;
        RECT -3.950 0.000 5.790 0.190 ;
        RECT 5.480 -0.120 5.790 0.000 ;
    END
  END ROW1
  PIN ROW2
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 5.490 -1.670 5.800 -1.480 ;
        RECT -3.950 -1.810 5.800 -1.670 ;
        RECT -3.950 -1.860 5.770 -1.810 ;
    END
  END ROW2
  OBS
      LAYER nwell ;
        RECT -0.190 -0.160 2.530 1.490 ;
        RECT -0.180 -0.200 2.530 -0.160 ;
        RECT -0.180 -1.530 2.530 -1.490 ;
        RECT -0.190 -3.180 2.530 -1.530 ;
      LAYER li1 ;
        RECT 4.730 1.800 4.920 1.830 ;
        RECT 3.860 1.630 4.920 1.800 ;
        RECT 5.160 1.650 5.690 1.820 ;
        RECT 3.860 1.240 4.030 1.630 ;
        RECT 4.730 1.600 4.920 1.630 ;
        RECT 6.970 1.550 7.170 1.900 ;
        RECT 6.970 1.520 7.180 1.550 ;
        RECT 3.290 1.070 4.030 1.240 ;
        RECT 4.260 1.240 4.450 1.270 ;
        RECT 4.260 1.070 4.990 1.240 ;
        RECT 4.260 1.040 4.450 1.070 ;
        RECT -3.520 0.090 -2.970 0.520 ;
        RECT 2.000 0.450 2.230 0.970 ;
        RECT 2.000 0.280 4.990 0.450 ;
        RECT 5.410 0.170 5.580 1.260 ;
        RECT 5.410 0.130 5.810 0.170 ;
        RECT 5.410 -0.060 5.820 0.130 ;
        RECT 5.410 -0.090 5.810 -0.060 ;
        RECT 4.730 -0.340 4.920 -0.160 ;
        RECT -0.920 -0.740 -0.730 -0.340 ;
        RECT 3.300 -0.510 3.640 -0.340 ;
        RECT -1.110 -0.750 -0.730 -0.740 ;
        RECT -1.110 -0.930 2.630 -0.750 ;
        RECT -1.110 -0.970 -0.730 -0.930 ;
        RECT -3.520 -1.640 -2.970 -1.210 ;
        RECT -0.920 -1.350 -0.730 -0.970 ;
        RECT 3.380 -1.080 3.550 -0.510 ;
        RECT 3.860 -0.920 4.070 -0.490 ;
        RECT 4.640 -0.510 4.990 -0.340 ;
        RECT 5.410 -0.430 5.580 -0.090 ;
        RECT 6.240 -0.340 6.410 1.270 ;
        RECT 6.960 0.940 7.180 1.520 ;
        RECT 6.970 0.930 7.180 0.940 ;
        RECT 6.610 0.760 6.800 0.770 ;
        RECT 6.610 0.470 6.810 0.760 ;
        RECT 6.600 0.140 6.870 0.470 ;
        RECT 6.240 -0.530 6.420 -0.340 ;
        RECT 3.880 -0.940 4.050 -0.920 ;
        RECT 3.300 -1.110 3.640 -1.080 ;
        RECT 4.260 -1.100 4.450 -1.050 ;
        RECT 4.220 -1.110 4.450 -1.100 ;
        RECT 3.300 -1.250 4.450 -1.110 ;
        RECT 4.640 -1.250 4.990 -1.080 ;
        RECT 3.470 -1.280 4.450 -1.250 ;
        RECT 3.470 -1.310 4.310 -1.280 ;
        RECT 4.720 -1.460 4.910 -1.250 ;
        RECT 5.410 -1.520 5.580 -1.160 ;
        RECT 6.240 -1.250 6.420 -1.060 ;
        RECT 5.410 -1.560 5.820 -1.520 ;
        RECT 5.410 -1.750 5.830 -1.560 ;
        RECT 5.410 -1.780 5.820 -1.750 ;
        RECT 2.060 -1.970 4.990 -1.870 ;
        RECT 2.000 -2.040 4.990 -1.970 ;
        RECT 2.000 -2.660 2.230 -2.040 ;
        RECT 2.800 -2.360 2.970 -2.300 ;
        RECT 2.780 -2.570 2.990 -2.360 ;
        RECT 2.800 -2.640 2.970 -2.570 ;
        RECT 4.270 -2.660 4.460 -2.630 ;
        RECT 3.290 -2.830 4.100 -2.660 ;
        RECT 3.910 -3.170 4.100 -2.830 ;
        RECT 4.270 -2.830 4.990 -2.660 ;
        RECT 4.270 -2.860 4.460 -2.830 ;
        RECT 5.410 -2.850 5.580 -1.780 ;
        RECT 6.240 -2.860 6.410 -1.250 ;
        RECT 6.600 -2.060 6.870 -1.730 ;
        RECT 6.610 -2.350 6.810 -2.060 ;
        RECT 6.610 -2.360 6.800 -2.350 ;
        RECT 6.970 -2.530 7.180 -2.520 ;
        RECT 6.960 -3.110 7.180 -2.530 ;
        RECT 6.970 -3.140 7.180 -3.110 ;
        RECT 4.700 -3.170 4.890 -3.140 ;
        RECT 3.910 -3.350 4.890 -3.170 ;
        RECT 4.700 -3.370 4.890 -3.350 ;
        RECT 5.160 -3.410 5.690 -3.240 ;
        RECT 6.970 -3.490 7.170 -3.140 ;
      LAYER mcon ;
        RECT 4.740 1.630 4.910 1.800 ;
        RECT 6.980 1.350 7.150 1.520 ;
        RECT 4.270 1.070 4.440 1.240 ;
        RECT 2.030 0.770 2.200 0.940 ;
        RECT -3.520 0.170 -3.250 0.440 ;
        RECT 2.030 0.320 2.200 0.490 ;
        RECT 5.550 -0.050 5.720 0.120 ;
        RECT 4.740 -0.360 4.910 -0.190 ;
        RECT -1.100 -0.940 -0.930 -0.770 ;
        RECT -3.520 -1.560 -3.250 -1.290 ;
        RECT 6.620 0.510 6.800 0.700 ;
        RECT 4.270 -1.250 4.440 -1.080 ;
        RECT 4.730 -1.430 4.900 -1.260 ;
        RECT 5.560 -1.740 5.730 -1.570 ;
        RECT 2.030 -2.180 2.200 -2.010 ;
        RECT 2.030 -2.630 2.200 -2.460 ;
        RECT 4.280 -2.830 4.450 -2.660 ;
        RECT 6.620 -2.290 6.800 -2.100 ;
        RECT 6.980 -3.110 7.150 -2.940 ;
        RECT 4.710 -3.340 4.880 -3.170 ;
      LAYER met1 ;
        RECT 5.090 1.410 5.400 1.850 ;
        RECT 1.990 0.230 2.250 1.020 ;
        RECT 5.480 -0.120 5.800 0.200 ;
        RECT 6.210 -0.630 6.450 -0.210 ;
        RECT 6.210 -0.950 6.480 -0.630 ;
        RECT 6.210 -1.380 6.450 -0.950 ;
        RECT 5.490 -1.810 5.810 -1.490 ;
        RECT 1.990 -2.710 2.250 -1.920 ;
        RECT 5.090 -3.440 5.400 -3.000 ;
      LAYER via ;
        RECT 5.120 1.440 5.380 1.700 ;
        RECT 5.510 -0.090 5.770 0.170 ;
        RECT 6.220 -0.920 6.480 -0.660 ;
        RECT 5.520 -1.780 5.780 -1.520 ;
        RECT 5.120 -3.290 5.380 -3.030 ;
  END
END sky130_hilas_FGtrans2x1cell

MACRO sky130_hilas_capacitorSize01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_capacitorSize01 ;
  ORIGIN -14.140 0.480 ;
  SIZE 10.420 BY 5.830 ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 23.740 2.130 24.400 2.790 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 14.250 2.720 14.910 2.780 ;
        RECT 15.300 2.720 16.310 2.730 ;
        RECT 14.250 2.220 17.940 2.720 ;
        RECT 14.250 2.210 15.660 2.220 ;
        RECT 14.250 2.120 14.910 2.210 ;
        RECT 17.300 1.100 17.930 2.220 ;
        RECT 17.300 1.090 19.450 1.100 ;
        RECT 16.490 0.620 19.530 1.090 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 14.140 4.800 24.560 4.980 ;
        RECT 14.140 4.370 24.560 4.550 ;
        RECT 14.170 3.370 24.560 3.550 ;
        RECT 22.650 3.120 24.560 3.130 ;
        RECT 14.170 2.940 24.560 3.120 ;
        RECT 14.380 2.600 14.750 2.660 ;
        RECT 14.160 2.320 14.750 2.600 ;
        RECT 14.380 2.260 14.750 2.320 ;
        RECT 23.870 2.610 24.240 2.670 ;
        RECT 23.870 2.330 24.560 2.610 ;
        RECT 23.870 2.270 24.240 2.330 ;
        RECT 14.170 1.790 24.560 1.960 ;
        RECT 14.170 1.370 24.560 1.540 ;
        RECT 14.170 0.390 24.560 0.560 ;
        RECT 14.170 -0.050 24.560 0.120 ;
      LAYER via2 ;
        RECT 14.430 2.320 14.710 2.600 ;
        RECT 23.920 2.330 24.200 2.610 ;
      LAYER met3 ;
        RECT 15.600 5.320 18.420 5.350 ;
        RECT 15.600 2.820 22.800 5.320 ;
        RECT 14.160 2.060 14.950 2.810 ;
        RECT 15.600 2.070 24.440 2.820 ;
        RECT 15.600 -0.460 22.800 2.070 ;
        RECT 18.390 -0.480 22.800 -0.460 ;
      LAYER via3 ;
        RECT 14.350 2.210 14.780 2.690 ;
        RECT 23.840 2.220 24.270 2.700 ;
  END
END sky130_hilas_capacitorSize01

MACRO sky130_hilas_Tgate4Double01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_Tgate4Double01 ;
  ORIGIN 0.360 1.410 ;
  SIZE 7.080 BY 6.050 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER nwell ;
        RECT -0.240 -1.410 3.230 4.640 ;
      LAYER met1 ;
        RECT 0.380 3.770 0.580 4.640 ;
        RECT 0.370 3.480 0.600 3.770 ;
        RECT 0.380 2.770 0.580 3.480 ;
        RECT 0.370 2.480 0.600 2.770 ;
        RECT 0.380 0.750 0.580 2.480 ;
        RECT 0.370 0.460 0.600 0.750 ;
        RECT 0.380 -0.250 0.580 0.460 ;
        RECT 0.370 -0.540 0.600 -0.250 ;
        RECT 0.380 -1.410 0.580 -0.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.210 3.770 6.400 4.640 ;
        RECT 6.190 3.480 6.420 3.770 ;
        RECT 6.210 2.770 6.400 3.480 ;
        RECT 6.190 2.480 6.420 2.770 ;
        RECT 6.210 0.750 6.400 2.480 ;
        RECT 6.190 0.460 6.420 0.750 ;
        RECT 6.210 -0.250 6.400 0.460 ;
        RECT 6.190 -0.540 6.420 -0.250 ;
        RECT 6.210 -1.410 6.400 -0.540 ;
    END
  END VGND
  PIN INPUT1_1
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.090 4.530 2.400 4.540 ;
        RECT -0.360 4.330 5.480 4.530 ;
        RECT 2.090 4.210 2.400 4.330 ;
        RECT 5.170 4.200 5.480 4.330 ;
    END
  END INPUT1_1
  PIN SELECT1
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER met2 ;
        RECT -0.360 3.350 0.250 3.550 ;
        RECT -0.070 3.260 0.250 3.350 ;
    END
  END SELECT1
  PIN SELECT2
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER met2 ;
        RECT -0.070 2.900 0.250 2.990 ;
        RECT -0.360 2.700 0.250 2.900 ;
    END
  END SELECT2
  PIN INPUT2_2
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 0.740 2.400 1.050 2.410 ;
        RECT 3.660 2.400 3.970 2.410 ;
        RECT -0.360 2.200 4.010 2.400 ;
        RECT 0.740 2.080 1.050 2.200 ;
        RECT 3.660 2.080 3.970 2.200 ;
    END
  END INPUT2_2
  PIN INPUT1_2
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.090 1.920 2.400 2.040 ;
        RECT 5.170 1.920 5.480 2.050 ;
        RECT -0.360 1.720 5.480 1.920 ;
        RECT 2.090 1.710 2.400 1.720 ;
    END
  END INPUT1_2
  PIN SELECT3
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER met2 ;
        RECT -0.360 0.330 0.250 0.530 ;
        RECT -0.070 0.240 0.250 0.330 ;
    END
  END SELECT3
  PIN INPUT2_3
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 0.740 1.030 1.050 1.150 ;
        RECT 3.660 1.030 3.970 1.150 ;
        RECT -0.360 0.830 4.010 1.030 ;
        RECT 0.740 0.820 1.050 0.830 ;
        RECT 3.660 0.820 3.970 0.830 ;
    END
  END INPUT2_3
  PIN SELECT4
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER met2 ;
        RECT -0.070 -0.120 0.250 -0.030 ;
        RECT -0.360 -0.320 0.250 -0.120 ;
    END
  END SELECT4
  PIN INPUT2_4
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 0.740 -0.620 1.050 -0.610 ;
        RECT 3.660 -0.620 3.970 -0.610 ;
        RECT -0.360 -0.820 4.010 -0.620 ;
        RECT 0.740 -0.940 1.050 -0.820 ;
        RECT 3.660 -0.940 3.970 -0.820 ;
    END
  END INPUT2_4
  PIN INPUT1_4
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.090 -1.100 2.400 -0.980 ;
        RECT 5.170 -1.100 5.480 -0.970 ;
        RECT -0.360 -1.300 5.480 -1.100 ;
        RECT 2.090 -1.310 2.400 -1.300 ;
    END
  END INPUT1_4
  PIN OUTPUT4
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER met2 ;
        RECT 1.320 -0.120 1.640 -0.110 ;
        RECT 2.740 -0.120 3.060 -0.100 ;
        RECT 4.490 -0.120 4.810 -0.080 ;
        RECT 5.530 -0.120 5.850 -0.090 ;
        RECT 1.320 -0.320 6.720 -0.120 ;
        RECT 1.320 -0.370 1.640 -0.320 ;
        RECT 2.740 -0.360 3.060 -0.320 ;
        RECT 4.490 -0.340 4.810 -0.320 ;
        RECT 5.530 -0.350 5.850 -0.320 ;
    END
  END OUTPUT4
  PIN OUTPUT3
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER met2 ;
        RECT 1.320 0.530 1.640 0.580 ;
        RECT 2.740 0.530 3.060 0.570 ;
        RECT 4.490 0.530 4.810 0.550 ;
        RECT 5.530 0.530 5.850 0.560 ;
        RECT 1.320 0.330 6.720 0.530 ;
        RECT 1.320 0.320 1.640 0.330 ;
        RECT 2.740 0.310 3.060 0.330 ;
        RECT 4.490 0.290 4.810 0.330 ;
        RECT 5.530 0.300 5.850 0.330 ;
    END
  END OUTPUT3
  PIN OUTPUT2
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER met2 ;
        RECT 1.320 2.900 1.640 2.910 ;
        RECT 2.740 2.900 3.060 2.920 ;
        RECT 4.490 2.900 4.810 2.940 ;
        RECT 5.530 2.900 5.850 2.930 ;
        RECT 1.320 2.700 6.720 2.900 ;
        RECT 1.320 2.650 1.640 2.700 ;
        RECT 2.740 2.660 3.060 2.700 ;
        RECT 4.490 2.680 4.810 2.700 ;
        RECT 5.530 2.670 5.850 2.700 ;
    END
  END OUTPUT2
  PIN OUTPUT1
    ANTENNADIFFAREA 0.365800 ;
    PORT
      LAYER met2 ;
        RECT 1.320 3.550 1.640 3.600 ;
        RECT 2.740 3.550 3.060 3.590 ;
        RECT 4.490 3.550 4.810 3.570 ;
        RECT 5.530 3.550 5.850 3.580 ;
        RECT 1.320 3.350 6.720 3.550 ;
        RECT 1.320 3.340 1.640 3.350 ;
        RECT 2.740 3.330 3.060 3.350 ;
        RECT 4.490 3.310 4.810 3.350 ;
        RECT 5.530 3.320 5.850 3.350 ;
    END
  END OUTPUT1
  PIN INPUT2_1
    ANTENNADIFFAREA 0.192200 ;
    PORT
      LAYER met2 ;
        RECT 0.740 4.050 1.050 4.170 ;
        RECT 3.660 4.050 3.970 4.170 ;
        RECT -0.360 3.850 4.010 4.050 ;
        RECT 0.740 3.840 1.050 3.850 ;
        RECT 3.660 3.840 3.970 3.850 ;
    END
  END INPUT2_1
  PIN INPUT1_3
    ANTENNADIFFAREA 0.179800 ;
    PORT
      LAYER met2 ;
        RECT 2.090 1.510 2.400 1.520 ;
        RECT -0.360 1.310 5.480 1.510 ;
        RECT 2.090 1.190 2.400 1.310 ;
        RECT 5.170 1.180 5.480 1.310 ;
    END
  END INPUT1_3
  OBS
      LAYER li1 ;
        RECT 2.100 4.480 2.420 4.510 ;
        RECT 0.070 4.130 0.240 4.410 ;
        RECT 0.580 4.170 0.930 4.340 ;
        RECT 0.750 4.140 0.930 4.170 ;
        RECT 1.350 4.150 1.520 4.420 ;
        RECT 2.100 4.290 2.430 4.480 ;
        RECT 5.180 4.470 5.500 4.500 ;
        RECT 2.100 4.250 2.420 4.290 ;
        RECT 0.070 4.090 0.280 4.130 ;
        RECT 0.750 4.110 1.070 4.140 ;
        RECT 0.070 4.070 0.300 4.090 ;
        RECT 0.070 4.050 0.330 4.070 ;
        RECT 0.070 4.000 0.410 4.050 ;
        RECT 0.070 3.940 0.560 4.000 ;
        RECT 0.070 3.910 0.580 3.940 ;
        RECT 0.110 3.880 0.580 3.910 ;
        RECT 0.750 3.920 1.080 4.110 ;
        RECT 1.350 3.930 1.550 4.150 ;
        RECT 2.130 4.080 2.300 4.250 ;
        RECT 2.820 4.130 2.990 4.420 ;
        RECT 3.780 4.140 3.950 4.420 ;
        RECT 4.520 4.140 4.690 4.430 ;
        RECT 5.180 4.280 5.510 4.470 ;
        RECT 5.750 4.330 5.940 4.360 ;
        RECT 5.180 4.240 5.500 4.280 ;
        RECT 1.360 3.920 1.550 3.930 ;
        RECT 0.750 3.880 1.070 3.920 ;
        RECT 2.810 3.900 3.000 4.130 ;
        RECT 3.670 4.110 3.990 4.140 ;
        RECT 3.670 3.920 4.000 4.110 ;
        RECT 3.670 3.880 3.990 3.920 ;
        RECT 4.520 3.910 4.710 4.140 ;
        RECT 5.240 4.080 5.410 4.240 ;
        RECT 5.750 4.160 6.190 4.330 ;
        RECT 5.750 4.130 5.940 4.160 ;
        RECT 0.240 3.830 0.580 3.880 ;
        RECT 0.360 3.820 0.580 3.830 ;
        RECT 0.370 3.790 0.580 3.820 ;
        RECT 0.390 3.710 0.580 3.790 ;
        RECT 1.750 3.710 2.080 3.830 ;
        RECT 6.470 3.740 6.640 4.420 ;
        RECT -0.100 3.660 0.070 3.680 ;
        RECT -0.120 3.230 0.090 3.660 ;
        RECT 0.390 3.540 0.910 3.710 ;
        RECT 0.390 3.510 0.580 3.540 ;
        RECT 1.260 3.530 5.480 3.710 ;
        RECT 6.210 3.700 6.640 3.740 ;
        RECT 5.860 3.540 6.640 3.700 ;
        RECT 5.860 3.530 6.400 3.540 ;
        RECT 6.210 3.510 6.400 3.530 ;
        RECT -0.120 2.590 0.090 3.020 ;
        RECT 0.390 2.710 0.580 2.740 ;
        RECT 6.210 2.720 6.400 2.740 ;
        RECT -0.100 2.570 0.070 2.590 ;
        RECT 0.390 2.540 0.910 2.710 ;
        RECT 1.260 2.540 5.480 2.720 ;
        RECT 5.860 2.710 6.400 2.720 ;
        RECT 5.860 2.550 6.640 2.710 ;
        RECT 0.390 2.460 0.580 2.540 ;
        RECT 0.370 2.430 0.580 2.460 ;
        RECT 0.360 2.420 0.580 2.430 ;
        RECT 1.750 2.420 2.080 2.540 ;
        RECT 6.210 2.510 6.640 2.550 ;
        RECT 0.240 2.370 0.580 2.420 ;
        RECT 0.110 2.340 0.580 2.370 ;
        RECT 0.070 2.310 0.580 2.340 ;
        RECT 0.750 2.330 1.070 2.370 ;
        RECT 0.070 2.250 0.560 2.310 ;
        RECT 0.070 2.200 0.410 2.250 ;
        RECT 0.070 2.180 0.330 2.200 ;
        RECT 0.070 2.160 0.300 2.180 ;
        RECT 0.070 2.120 0.280 2.160 ;
        RECT 0.750 2.140 1.080 2.330 ;
        RECT 1.360 2.320 1.550 2.330 ;
        RECT 0.070 1.840 0.240 2.120 ;
        RECT 0.750 2.110 1.070 2.140 ;
        RECT 0.750 2.080 0.930 2.110 ;
        RECT 0.580 1.910 0.930 2.080 ;
        RECT 1.350 2.100 1.550 2.320 ;
        RECT 1.350 1.830 1.520 2.100 ;
        RECT 2.130 2.000 2.300 2.170 ;
        RECT 2.810 2.120 3.000 2.350 ;
        RECT 3.670 2.330 3.990 2.370 ;
        RECT 3.670 2.140 4.000 2.330 ;
        RECT 2.100 1.960 2.420 2.000 ;
        RECT 2.100 1.770 2.430 1.960 ;
        RECT 2.820 1.830 2.990 2.120 ;
        RECT 3.670 2.110 3.990 2.140 ;
        RECT 4.520 2.110 4.710 2.340 ;
        RECT 3.780 1.830 3.950 2.110 ;
        RECT 4.520 1.820 4.690 2.110 ;
        RECT 5.240 2.010 5.410 2.170 ;
        RECT 5.750 2.090 5.940 2.120 ;
        RECT 5.180 1.970 5.500 2.010 ;
        RECT 5.180 1.780 5.510 1.970 ;
        RECT 5.750 1.920 6.190 2.090 ;
        RECT 5.750 1.890 5.940 1.920 ;
        RECT 6.470 1.830 6.640 2.510 ;
        RECT 2.100 1.740 2.420 1.770 ;
        RECT 5.180 1.750 5.500 1.780 ;
        RECT 2.100 1.460 2.420 1.490 ;
        RECT 0.070 1.110 0.240 1.390 ;
        RECT 0.580 1.150 0.930 1.320 ;
        RECT 0.750 1.120 0.930 1.150 ;
        RECT 1.350 1.130 1.520 1.400 ;
        RECT 2.100 1.270 2.430 1.460 ;
        RECT 5.180 1.450 5.500 1.480 ;
        RECT 2.100 1.230 2.420 1.270 ;
        RECT 0.070 1.070 0.280 1.110 ;
        RECT 0.750 1.090 1.070 1.120 ;
        RECT 0.070 1.050 0.300 1.070 ;
        RECT 0.070 1.030 0.330 1.050 ;
        RECT 0.070 0.980 0.410 1.030 ;
        RECT 0.070 0.920 0.560 0.980 ;
        RECT 0.070 0.890 0.580 0.920 ;
        RECT 0.110 0.860 0.580 0.890 ;
        RECT 0.750 0.900 1.080 1.090 ;
        RECT 1.350 0.910 1.550 1.130 ;
        RECT 2.130 1.060 2.300 1.230 ;
        RECT 2.820 1.110 2.990 1.400 ;
        RECT 3.780 1.120 3.950 1.400 ;
        RECT 4.520 1.120 4.690 1.410 ;
        RECT 5.180 1.260 5.510 1.450 ;
        RECT 5.750 1.310 5.940 1.340 ;
        RECT 5.180 1.220 5.500 1.260 ;
        RECT 1.360 0.900 1.550 0.910 ;
        RECT 0.750 0.860 1.070 0.900 ;
        RECT 2.810 0.880 3.000 1.110 ;
        RECT 3.670 1.090 3.990 1.120 ;
        RECT 3.670 0.900 4.000 1.090 ;
        RECT 3.670 0.860 3.990 0.900 ;
        RECT 4.520 0.890 4.710 1.120 ;
        RECT 5.240 1.060 5.410 1.220 ;
        RECT 5.750 1.140 6.190 1.310 ;
        RECT 5.750 1.110 5.940 1.140 ;
        RECT 0.240 0.810 0.580 0.860 ;
        RECT 0.360 0.800 0.580 0.810 ;
        RECT 0.370 0.770 0.580 0.800 ;
        RECT 0.390 0.690 0.580 0.770 ;
        RECT 1.750 0.690 2.080 0.810 ;
        RECT 6.470 0.720 6.640 1.400 ;
        RECT -0.100 0.640 0.070 0.660 ;
        RECT -0.120 0.210 0.090 0.640 ;
        RECT 0.390 0.520 0.910 0.690 ;
        RECT 0.390 0.490 0.580 0.520 ;
        RECT 1.260 0.510 5.480 0.690 ;
        RECT 6.210 0.680 6.640 0.720 ;
        RECT 5.860 0.520 6.640 0.680 ;
        RECT 5.860 0.510 6.400 0.520 ;
        RECT 6.210 0.490 6.400 0.510 ;
        RECT -0.120 -0.430 0.090 0.000 ;
        RECT 0.390 -0.310 0.580 -0.280 ;
        RECT 6.210 -0.300 6.400 -0.280 ;
        RECT -0.100 -0.450 0.070 -0.430 ;
        RECT 0.390 -0.480 0.910 -0.310 ;
        RECT 1.260 -0.480 5.480 -0.300 ;
        RECT 5.860 -0.310 6.400 -0.300 ;
        RECT 5.860 -0.470 6.640 -0.310 ;
        RECT 0.390 -0.560 0.580 -0.480 ;
        RECT 0.370 -0.590 0.580 -0.560 ;
        RECT 0.360 -0.600 0.580 -0.590 ;
        RECT 1.750 -0.600 2.080 -0.480 ;
        RECT 6.210 -0.510 6.640 -0.470 ;
        RECT 0.240 -0.650 0.580 -0.600 ;
        RECT 0.110 -0.680 0.580 -0.650 ;
        RECT 0.070 -0.710 0.580 -0.680 ;
        RECT 0.750 -0.690 1.070 -0.650 ;
        RECT 0.070 -0.770 0.560 -0.710 ;
        RECT 0.070 -0.820 0.410 -0.770 ;
        RECT 0.070 -0.840 0.330 -0.820 ;
        RECT 0.070 -0.860 0.300 -0.840 ;
        RECT 0.070 -0.900 0.280 -0.860 ;
        RECT 0.750 -0.880 1.080 -0.690 ;
        RECT 1.360 -0.700 1.550 -0.690 ;
        RECT 0.070 -1.180 0.240 -0.900 ;
        RECT 0.750 -0.910 1.070 -0.880 ;
        RECT 0.750 -0.940 0.930 -0.910 ;
        RECT 0.580 -1.110 0.930 -0.940 ;
        RECT 1.350 -0.920 1.550 -0.700 ;
        RECT 1.350 -1.190 1.520 -0.920 ;
        RECT 2.130 -1.020 2.300 -0.850 ;
        RECT 2.810 -0.900 3.000 -0.670 ;
        RECT 3.670 -0.690 3.990 -0.650 ;
        RECT 3.670 -0.880 4.000 -0.690 ;
        RECT 2.100 -1.060 2.420 -1.020 ;
        RECT 2.100 -1.250 2.430 -1.060 ;
        RECT 2.820 -1.190 2.990 -0.900 ;
        RECT 3.670 -0.910 3.990 -0.880 ;
        RECT 4.520 -0.910 4.710 -0.680 ;
        RECT 3.780 -1.190 3.950 -0.910 ;
        RECT 4.520 -1.200 4.690 -0.910 ;
        RECT 5.240 -1.010 5.410 -0.850 ;
        RECT 5.750 -0.930 5.940 -0.900 ;
        RECT 5.180 -1.050 5.500 -1.010 ;
        RECT 5.180 -1.240 5.510 -1.050 ;
        RECT 5.750 -1.100 6.190 -0.930 ;
        RECT 5.750 -1.130 5.940 -1.100 ;
        RECT 6.470 -1.190 6.640 -0.510 ;
        RECT 2.100 -1.280 2.420 -1.250 ;
        RECT 5.180 -1.270 5.500 -1.240 ;
      LAYER mcon ;
        RECT 2.160 4.300 2.330 4.470 ;
        RECT 0.810 3.930 0.980 4.100 ;
        RECT 1.370 3.950 1.540 4.120 ;
        RECT 5.240 4.290 5.410 4.460 ;
        RECT 2.820 3.930 2.990 4.100 ;
        RECT 3.730 3.930 3.900 4.100 ;
        RECT 4.530 3.940 4.700 4.110 ;
        RECT 5.760 4.160 5.930 4.330 ;
        RECT -0.100 3.510 0.070 3.680 ;
        RECT 0.400 3.540 0.570 3.710 ;
        RECT 6.220 3.540 6.390 3.710 ;
        RECT 0.400 2.540 0.570 2.710 ;
        RECT 6.220 2.540 6.390 2.710 ;
        RECT 0.810 2.150 0.980 2.320 ;
        RECT 1.370 2.130 1.540 2.300 ;
        RECT 2.820 2.150 2.990 2.320 ;
        RECT 3.730 2.150 3.900 2.320 ;
        RECT 4.530 2.140 4.700 2.310 ;
        RECT 2.160 1.780 2.330 1.950 ;
        RECT 5.240 1.790 5.410 1.960 ;
        RECT 5.760 1.920 5.930 2.090 ;
        RECT 2.160 1.280 2.330 1.450 ;
        RECT 0.810 0.910 0.980 1.080 ;
        RECT 1.370 0.930 1.540 1.100 ;
        RECT 5.240 1.270 5.410 1.440 ;
        RECT 2.820 0.910 2.990 1.080 ;
        RECT 3.730 0.910 3.900 1.080 ;
        RECT 4.530 0.920 4.700 1.090 ;
        RECT 5.760 1.140 5.930 1.310 ;
        RECT -0.100 0.490 0.070 0.660 ;
        RECT 0.400 0.520 0.570 0.690 ;
        RECT 6.220 0.520 6.390 0.690 ;
        RECT 0.400 -0.480 0.570 -0.310 ;
        RECT 6.220 -0.480 6.390 -0.310 ;
        RECT 0.810 -0.870 0.980 -0.700 ;
        RECT 1.370 -0.890 1.540 -0.720 ;
        RECT 2.820 -0.870 2.990 -0.700 ;
        RECT 3.730 -0.870 3.900 -0.700 ;
        RECT 4.530 -0.880 4.700 -0.710 ;
        RECT 2.160 -1.240 2.330 -1.070 ;
        RECT 5.240 -1.230 5.410 -1.060 ;
        RECT 5.760 -1.100 5.930 -0.930 ;
      LAYER met1 ;
        RECT 2.090 4.220 2.410 4.540 ;
        RECT 5.170 4.210 5.490 4.530 ;
        RECT 0.740 3.850 1.060 4.170 ;
        RECT 1.340 3.890 1.570 4.180 ;
        RECT -0.130 3.550 0.100 3.740 ;
        RECT 1.360 3.630 1.530 3.890 ;
        RECT 2.790 3.870 3.020 4.160 ;
        RECT -0.130 3.450 0.220 3.550 ;
        RECT -0.120 3.230 0.220 3.450 ;
        RECT 1.350 3.310 1.610 3.630 ;
        RECT 2.810 3.620 2.980 3.870 ;
        RECT 3.660 3.850 3.980 4.170 ;
        RECT 4.500 3.880 4.730 4.170 ;
        RECT 5.730 4.100 5.960 4.390 ;
        RECT 2.770 3.300 3.030 3.620 ;
        RECT 4.530 3.600 4.700 3.880 ;
        RECT 5.730 3.610 5.920 4.100 ;
        RECT 4.520 3.280 4.780 3.600 ;
        RECT 5.560 3.360 5.920 3.610 ;
        RECT 5.560 3.290 5.820 3.360 ;
        RECT -0.120 2.800 0.220 3.020 ;
        RECT -0.130 2.700 0.220 2.800 ;
        RECT -0.130 2.510 0.100 2.700 ;
        RECT 1.350 2.620 1.610 2.940 ;
        RECT 2.770 2.630 3.030 2.950 ;
        RECT 4.520 2.650 4.780 2.970 ;
        RECT 5.560 2.890 5.820 2.960 ;
        RECT 0.740 2.080 1.060 2.400 ;
        RECT 1.360 2.360 1.530 2.620 ;
        RECT 2.810 2.380 2.980 2.630 ;
        RECT 1.340 2.070 1.570 2.360 ;
        RECT 2.790 2.090 3.020 2.380 ;
        RECT 3.660 2.080 3.980 2.400 ;
        RECT 4.530 2.370 4.700 2.650 ;
        RECT 5.560 2.640 5.920 2.890 ;
        RECT 4.500 2.080 4.730 2.370 ;
        RECT 5.730 2.150 5.920 2.640 ;
        RECT 2.090 1.710 2.410 2.030 ;
        RECT 5.170 1.720 5.490 2.040 ;
        RECT 5.730 1.860 5.960 2.150 ;
        RECT 2.090 1.200 2.410 1.520 ;
        RECT 5.170 1.190 5.490 1.510 ;
        RECT 0.740 0.830 1.060 1.150 ;
        RECT 1.340 0.870 1.570 1.160 ;
        RECT -0.130 0.530 0.100 0.720 ;
        RECT 1.360 0.610 1.530 0.870 ;
        RECT 2.790 0.850 3.020 1.140 ;
        RECT -0.130 0.430 0.220 0.530 ;
        RECT -0.120 0.210 0.220 0.430 ;
        RECT 1.350 0.290 1.610 0.610 ;
        RECT 2.810 0.600 2.980 0.850 ;
        RECT 3.660 0.830 3.980 1.150 ;
        RECT 4.500 0.860 4.730 1.150 ;
        RECT 5.730 1.080 5.960 1.370 ;
        RECT 2.770 0.280 3.030 0.600 ;
        RECT 4.530 0.580 4.700 0.860 ;
        RECT 5.730 0.590 5.920 1.080 ;
        RECT 4.520 0.260 4.780 0.580 ;
        RECT 5.560 0.340 5.920 0.590 ;
        RECT 5.560 0.270 5.820 0.340 ;
        RECT -0.120 -0.220 0.220 0.000 ;
        RECT -0.130 -0.320 0.220 -0.220 ;
        RECT -0.130 -0.510 0.100 -0.320 ;
        RECT 1.350 -0.400 1.610 -0.080 ;
        RECT 2.770 -0.390 3.030 -0.070 ;
        RECT 4.520 -0.370 4.780 -0.050 ;
        RECT 5.560 -0.130 5.820 -0.060 ;
        RECT 0.740 -0.940 1.060 -0.620 ;
        RECT 1.360 -0.660 1.530 -0.400 ;
        RECT 2.810 -0.640 2.980 -0.390 ;
        RECT 1.340 -0.950 1.570 -0.660 ;
        RECT 2.790 -0.930 3.020 -0.640 ;
        RECT 3.660 -0.940 3.980 -0.620 ;
        RECT 4.530 -0.650 4.700 -0.370 ;
        RECT 5.560 -0.380 5.920 -0.130 ;
        RECT 4.500 -0.940 4.730 -0.650 ;
        RECT 5.730 -0.870 5.920 -0.380 ;
        RECT 2.090 -1.310 2.410 -0.990 ;
        RECT 5.170 -1.300 5.490 -0.980 ;
        RECT 5.730 -1.160 5.960 -0.870 ;
      LAYER via ;
        RECT 2.120 4.250 2.380 4.510 ;
        RECT 5.200 4.240 5.460 4.500 ;
        RECT 0.770 3.880 1.030 4.140 ;
        RECT 3.690 3.880 3.950 4.140 ;
        RECT -0.040 3.260 0.220 3.520 ;
        RECT 1.350 3.340 1.610 3.600 ;
        RECT 2.770 3.330 3.030 3.590 ;
        RECT 4.520 3.310 4.780 3.570 ;
        RECT 5.560 3.320 5.820 3.580 ;
        RECT -0.040 2.730 0.220 2.990 ;
        RECT 1.350 2.650 1.610 2.910 ;
        RECT 2.770 2.660 3.030 2.920 ;
        RECT 4.520 2.680 4.780 2.940 ;
        RECT 5.560 2.670 5.820 2.930 ;
        RECT 0.770 2.110 1.030 2.370 ;
        RECT 3.690 2.110 3.950 2.370 ;
        RECT 2.120 1.740 2.380 2.000 ;
        RECT 5.200 1.750 5.460 2.010 ;
        RECT 2.120 1.230 2.380 1.490 ;
        RECT 5.200 1.220 5.460 1.480 ;
        RECT 0.770 0.860 1.030 1.120 ;
        RECT 3.690 0.860 3.950 1.120 ;
        RECT -0.040 0.240 0.220 0.500 ;
        RECT 1.350 0.320 1.610 0.580 ;
        RECT 2.770 0.310 3.030 0.570 ;
        RECT 4.520 0.290 4.780 0.550 ;
        RECT 5.560 0.300 5.820 0.560 ;
        RECT -0.040 -0.290 0.220 -0.030 ;
        RECT 1.350 -0.370 1.610 -0.110 ;
        RECT 2.770 -0.360 3.030 -0.100 ;
        RECT 4.520 -0.340 4.780 -0.080 ;
        RECT 5.560 -0.350 5.820 -0.090 ;
        RECT 0.770 -0.910 1.030 -0.650 ;
        RECT 3.690 -0.910 3.950 -0.650 ;
        RECT 2.120 -1.280 2.380 -1.020 ;
        RECT 5.200 -1.270 5.460 -1.010 ;
  END
END sky130_hilas_Tgate4Double01

MACRO sky130_hilas_cellAttempt01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_cellAttempt01 ;
  ORIGIN 2.630 4.040 ;
  SIZE 10.070 BY 6.500 ;
  PIN VTUN
    ANTENNADIFFAREA 2.237600 ;
    PORT
      LAYER nwell ;
        RECT -2.630 -4.040 -0.900 2.450 ;
      LAYER met1 ;
        RECT -2.280 -4.040 -1.880 2.460 ;
    END
  END VTUN
  PIN VINJ
    ANTENNADIFFAREA 1.088000 ;
    PORT
      LAYER nwell ;
        RECT 4.880 -4.040 7.440 2.460 ;
      LAYER met1 ;
        RECT 6.920 1.750 7.080 2.450 ;
        RECT 6.810 1.200 7.080 1.750 ;
        RECT 6.810 1.150 7.090 1.200 ;
        RECT 6.920 1.060 7.090 1.150 ;
        RECT 6.920 0.590 7.080 1.060 ;
        RECT 6.920 0.500 7.090 0.590 ;
        RECT 6.810 0.450 7.090 0.500 ;
        RECT 6.810 -0.100 7.080 0.450 ;
        RECT 6.920 -1.490 7.080 -0.100 ;
        RECT 6.810 -2.040 7.080 -1.490 ;
        RECT 6.810 -2.090 7.090 -2.040 ;
        RECT 6.920 -2.180 7.090 -2.090 ;
        RECT 6.920 -2.640 7.080 -2.180 ;
        RECT 6.920 -2.730 7.090 -2.640 ;
        RECT 6.810 -2.780 7.090 -2.730 ;
        RECT 6.810 -3.330 7.080 -2.780 ;
        RECT 6.920 -4.030 7.080 -3.330 ;
    END
  END VINJ
  PIN COLSEL1
    ANTENNAGATEAREA 0.720000 ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met1 ;
        RECT 6.110 1.720 6.270 2.450 ;
        RECT 6.110 1.700 6.310 1.720 ;
        RECT 6.090 1.460 6.320 1.700 ;
        RECT 6.110 1.410 6.320 1.460 ;
        RECT 6.480 1.410 6.670 2.400 ;
        RECT 6.110 0.240 6.270 1.410 ;
        RECT 6.500 1.290 6.670 1.410 ;
        RECT 6.510 0.360 6.670 1.290 ;
        RECT 6.500 0.240 6.670 0.360 ;
        RECT 6.110 0.190 6.320 0.240 ;
        RECT 6.090 -0.050 6.320 0.190 ;
        RECT 6.110 -0.070 6.310 -0.050 ;
        RECT 6.110 -0.700 6.270 -0.070 ;
        RECT 6.480 -0.680 6.670 0.240 ;
        RECT 6.460 -0.700 6.700 -0.680 ;
        RECT 6.110 -0.890 6.700 -0.700 ;
        RECT 6.110 -1.520 6.270 -0.890 ;
        RECT 6.460 -0.910 6.700 -0.890 ;
        RECT 6.110 -1.540 6.310 -1.520 ;
        RECT 6.090 -1.780 6.320 -1.540 ;
        RECT 6.110 -1.830 6.320 -1.780 ;
        RECT 6.480 -1.830 6.670 -0.910 ;
        RECT 6.110 -2.990 6.270 -1.830 ;
        RECT 6.500 -1.950 6.670 -1.830 ;
        RECT 6.510 -2.870 6.670 -1.950 ;
        RECT 6.500 -2.990 6.670 -2.870 ;
        RECT 6.110 -3.040 6.320 -2.990 ;
        RECT 6.090 -3.280 6.320 -3.040 ;
        RECT 6.110 -3.300 6.310 -3.280 ;
        RECT 6.110 -4.030 6.270 -3.300 ;
        RECT 6.480 -3.980 6.670 -2.990 ;
    END
  END COLSEL1
  PIN GATE1
    ANTENNADIFFAREA 3.253900 ;
    PORT
      LAYER nwell ;
        RECT 1.120 -4.040 3.350 2.450 ;
      LAYER met1 ;
        RECT 1.770 0.310 2.150 2.460 ;
        RECT 1.760 -1.550 2.150 0.310 ;
        RECT 1.770 -4.040 2.150 -1.550 ;
    END
  END GATE1
  PIN ROW4
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 4.970 -2.870 5.280 -2.740 ;
        RECT -2.630 -3.050 7.440 -2.870 ;
        RECT 4.970 -3.070 5.280 -3.050 ;
    END
  END ROW4
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.120 -2.260 0.440 -2.250 ;
        RECT 4.050 -2.260 4.370 -2.200 ;
        RECT 0.120 -2.440 4.370 -2.260 ;
        RECT 0.120 -2.510 0.440 -2.440 ;
        RECT 4.050 -2.490 4.370 -2.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.090 1.070 4.330 2.460 ;
        RECT 4.070 0.410 4.340 1.070 ;
        RECT 4.090 -2.180 4.330 0.410 ;
        RECT 4.080 -2.500 4.340 -2.180 ;
        RECT 4.090 -4.040 4.330 -2.500 ;
      LAYER via ;
        RECT 4.080 -2.470 4.340 -2.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.160 1.050 0.400 2.460 ;
        RECT 0.150 0.390 0.410 1.050 ;
        RECT 0.160 -2.220 0.400 0.390 ;
        RECT 0.150 -2.540 0.410 -2.220 ;
        RECT 0.160 -4.040 0.400 -2.540 ;
      LAYER via ;
        RECT 0.150 -2.510 0.410 -2.250 ;
    END
  END VGND
  PIN DRAIN4
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 4.970 -3.300 5.280 -3.290 ;
        RECT -2.630 -3.470 7.440 -3.300 ;
        RECT 4.970 -3.480 7.440 -3.470 ;
        RECT 4.970 -3.620 5.280 -3.480 ;
    END
  END DRAIN4
  PIN DRAIN1
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 4.970 1.900 5.280 2.040 ;
        RECT -2.630 1.720 7.440 1.900 ;
        RECT 4.970 1.710 5.280 1.720 ;
    END
  END DRAIN1
  PIN ROW1
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 4.970 1.470 5.280 1.490 ;
        RECT 4.880 1.460 7.440 1.470 ;
        RECT -2.630 1.290 7.440 1.460 ;
        RECT -2.630 1.280 5.280 1.290 ;
        RECT 4.970 1.160 5.280 1.280 ;
    END
  END ROW1
  PIN ROW3
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 4.970 -1.770 5.280 -1.750 ;
        RECT -2.630 -1.950 7.440 -1.770 ;
        RECT 4.970 -2.080 5.280 -1.950 ;
    END
  END ROW3
  PIN DRAIN3
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 4.970 -1.340 5.280 -1.200 ;
        RECT -2.630 -1.520 7.440 -1.340 ;
        RECT 4.970 -1.530 5.280 -1.520 ;
    END
  END DRAIN3
  PIN DRAIN2
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT 4.970 -0.070 5.280 -0.060 ;
        RECT -2.630 -0.250 7.440 -0.070 ;
        RECT 4.970 -0.390 5.280 -0.250 ;
    END
  END DRAIN2
  PIN ROW2
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER met2 ;
        RECT 4.970 0.360 5.280 0.490 ;
        RECT -2.630 0.180 7.440 0.360 ;
        RECT 4.970 0.160 5.280 0.180 ;
    END
  END ROW2
  OBS
      LAYER li1 ;
        RECT 4.980 1.990 5.300 2.000 ;
        RECT 4.980 1.820 5.560 1.990 ;
        RECT 4.980 1.770 5.310 1.820 ;
        RECT 4.980 1.740 5.300 1.770 ;
        RECT 6.840 1.720 7.040 2.070 ;
        RECT 4.980 1.410 5.300 1.450 ;
        RECT 4.980 1.370 5.310 1.410 ;
        RECT 4.980 1.200 5.560 1.370 ;
        RECT 4.980 1.190 5.300 1.200 ;
        RECT 6.110 1.100 6.310 1.700 ;
        RECT 6.840 1.690 7.050 1.720 ;
        RECT 6.830 1.100 7.050 1.690 ;
        RECT 0.190 0.480 0.360 1.010 ;
        RECT 4.130 0.470 4.300 1.000 ;
        RECT 4.980 0.450 5.300 0.460 ;
        RECT 4.980 0.280 5.560 0.450 ;
        RECT 4.980 0.240 5.310 0.280 ;
        RECT 4.980 0.200 5.300 0.240 ;
        RECT 6.110 -0.050 6.310 0.550 ;
        RECT 6.830 -0.040 7.050 0.550 ;
        RECT 6.840 -0.070 7.050 -0.040 ;
        RECT 4.980 -0.120 5.300 -0.090 ;
        RECT 4.980 -0.170 5.310 -0.120 ;
        RECT -2.210 -1.020 -1.660 -0.590 ;
        RECT 0.200 -1.230 0.370 -0.220 ;
        RECT 4.980 -0.340 5.560 -0.170 ;
        RECT 4.980 -0.350 5.300 -0.340 ;
        RECT 1.820 -1.090 2.370 -0.660 ;
        RECT 4.130 -1.370 4.300 -0.360 ;
        RECT 6.840 -0.420 7.040 -0.070 ;
        RECT 6.230 -0.880 6.670 -0.710 ;
        RECT 4.980 -1.250 5.300 -1.240 ;
        RECT 4.980 -1.420 5.560 -1.250 ;
        RECT 4.980 -1.470 5.310 -1.420 ;
        RECT 4.980 -1.500 5.300 -1.470 ;
        RECT 6.840 -1.520 7.040 -1.170 ;
        RECT 4.980 -1.830 5.300 -1.790 ;
        RECT 4.980 -1.870 5.310 -1.830 ;
        RECT 4.980 -2.040 5.560 -1.870 ;
        RECT 4.980 -2.050 5.300 -2.040 ;
        RECT 6.110 -2.140 6.310 -1.540 ;
        RECT 6.840 -1.550 7.050 -1.520 ;
        RECT 6.830 -2.140 7.050 -1.550 ;
        RECT 4.980 -2.780 5.300 -2.770 ;
        RECT 4.980 -2.950 5.560 -2.780 ;
        RECT 4.980 -2.990 5.310 -2.950 ;
        RECT 4.980 -3.030 5.300 -2.990 ;
        RECT 6.110 -3.280 6.310 -2.680 ;
        RECT 6.830 -3.270 7.050 -2.680 ;
        RECT 6.840 -3.300 7.050 -3.270 ;
        RECT 4.980 -3.350 5.300 -3.320 ;
        RECT 4.980 -3.400 5.310 -3.350 ;
        RECT 4.980 -3.570 5.560 -3.400 ;
        RECT 4.980 -3.580 5.300 -3.570 ;
        RECT 6.840 -3.650 7.040 -3.300 ;
      LAYER mcon ;
        RECT 5.040 1.780 5.210 1.950 ;
        RECT 6.120 1.490 6.290 1.660 ;
        RECT 5.040 1.230 5.210 1.400 ;
        RECT 6.850 1.520 7.020 1.690 ;
        RECT 0.190 0.840 0.360 1.010 ;
        RECT 4.130 0.830 4.300 1.000 ;
        RECT 5.040 0.250 5.210 0.420 ;
        RECT 6.120 -0.010 6.290 0.160 ;
        RECT 6.850 -0.040 7.020 0.130 ;
        RECT 5.040 -0.300 5.210 -0.130 ;
        RECT -2.210 -0.940 -1.940 -0.670 ;
        RECT 0.200 -0.620 0.370 -0.450 ;
        RECT 0.200 -0.980 0.370 -0.810 ;
        RECT 1.820 -1.010 2.090 -0.740 ;
        RECT 4.130 -0.760 4.300 -0.590 ;
        RECT 6.490 -0.880 6.670 -0.710 ;
        RECT 4.130 -1.120 4.300 -0.950 ;
        RECT 5.040 -1.460 5.210 -1.290 ;
        RECT 6.120 -1.750 6.290 -1.580 ;
        RECT 5.040 -2.010 5.210 -1.840 ;
        RECT 6.850 -1.720 7.020 -1.550 ;
        RECT 5.040 -2.980 5.210 -2.810 ;
        RECT 6.120 -3.240 6.290 -3.070 ;
        RECT 6.850 -3.270 7.020 -3.100 ;
        RECT 5.040 -3.530 5.210 -3.360 ;
      LAYER met1 ;
        RECT 4.970 1.710 5.290 2.030 ;
        RECT 4.970 1.160 5.290 1.480 ;
        RECT 4.970 0.170 5.290 0.490 ;
        RECT 4.970 -0.380 5.290 -0.060 ;
        RECT 4.970 -1.530 5.290 -1.210 ;
        RECT 4.970 -2.080 5.290 -1.760 ;
        RECT 4.970 -3.060 5.290 -2.740 ;
        RECT 4.970 -3.610 5.290 -3.290 ;
      LAYER via ;
        RECT 5.000 1.740 5.260 2.000 ;
        RECT 5.000 1.190 5.260 1.450 ;
        RECT 5.000 0.200 5.260 0.460 ;
        RECT 5.000 -0.350 5.260 -0.090 ;
        RECT 5.000 -1.500 5.260 -1.240 ;
        RECT 5.000 -2.050 5.260 -1.790 ;
        RECT 5.000 -3.030 5.260 -2.770 ;
        RECT 5.000 -3.580 5.260 -3.320 ;
  END
END sky130_hilas_cellAttempt01

MACRO sky130_hilas_StepUpDigital
  CLASS BLOCK ;
  FOREIGN sky130_hilas_StepUpDigital ;
  ORIGIN 0.740 0.440 ;
  SIZE 9.630 BY 1.750 ;
  OBS
      LAYER nwell ;
        RECT 0.190 -0.440 2.690 1.310 ;
        RECT 6.560 -0.440 8.330 1.310 ;
      LAYER li1 ;
        RECT 1.470 0.800 1.920 0.950 ;
        RECT 0.530 0.620 0.860 0.790 ;
        RECT 1.320 0.630 1.920 0.800 ;
        RECT 0.600 0.160 0.780 0.620 ;
        RECT 2.120 0.190 2.290 0.950 ;
        RECT 2.620 0.860 2.910 0.880 ;
        RECT 2.620 0.820 3.080 0.860 ;
        RECT 2.620 0.800 4.060 0.820 ;
        RECT 2.620 0.640 4.100 0.800 ;
        RECT 2.910 0.630 4.100 0.640 ;
        RECT 4.550 0.770 5.010 0.800 ;
        RECT 6.320 0.770 6.670 0.870 ;
        RECT 4.550 0.630 5.660 0.770 ;
        RECT 4.840 0.600 5.660 0.630 ;
        RECT 5.900 0.600 7.070 0.770 ;
        RECT 7.320 0.600 8.080 0.770 ;
        RECT 4.840 0.460 5.100 0.600 ;
        RECT 3.920 0.290 5.100 0.460 ;
        RECT 7.850 0.590 8.080 0.600 ;
        RECT 2.120 0.180 2.500 0.190 ;
        RECT 0.600 -0.010 1.560 0.160 ;
        RECT 2.030 0.120 2.500 0.180 ;
        RECT 2.030 0.010 3.370 0.120 ;
        RECT 2.110 -0.050 3.370 0.010 ;
        RECT 2.110 -0.100 2.500 -0.050 ;
        RECT 3.920 -0.150 4.100 0.290 ;
        RECT 4.840 0.150 5.100 0.290 ;
        RECT 6.310 0.150 6.640 0.410 ;
        RECT 7.850 0.150 8.120 0.590 ;
        RECT 4.340 -0.210 4.550 0.120 ;
        RECT 4.840 -0.020 5.170 0.150 ;
        RECT 5.410 -0.020 7.570 0.150 ;
        RECT 4.840 -0.070 5.010 -0.020 ;
        RECT 7.820 -0.030 8.150 0.150 ;
        RECT 8.500 0.010 8.670 0.070 ;
        RECT 8.480 -0.210 8.700 0.010 ;
        RECT 8.500 -0.260 8.670 -0.210 ;
      LAYER mcon ;
        RECT 1.640 0.700 1.810 0.870 ;
        RECT 0.600 0.360 0.770 0.530 ;
        RECT 2.680 0.660 2.850 0.830 ;
        RECT 6.380 0.640 6.590 0.850 ;
        RECT 0.600 0.000 0.770 0.170 ;
        RECT 7.890 0.270 8.060 0.440 ;
      LAYER met1 ;
        RECT 0.530 -0.440 0.820 1.310 ;
        RECT 1.570 0.650 1.890 0.950 ;
        RECT 2.620 0.880 2.930 0.890 ;
        RECT 2.610 0.610 2.930 0.880 ;
        RECT 2.620 0.600 2.910 0.610 ;
        RECT 4.310 -0.150 4.590 0.180 ;
        RECT 4.840 -0.440 5.150 1.310 ;
        RECT 6.320 0.600 6.670 0.890 ;
        RECT 6.470 0.580 6.670 0.600 ;
        RECT 7.850 -0.440 8.090 1.310 ;
        RECT 8.420 -0.260 8.830 0.070 ;
      LAYER via ;
        RECT 1.600 0.660 1.860 0.920 ;
        RECT 2.640 0.620 2.900 0.880 ;
        RECT 4.320 -0.110 4.580 0.150 ;
        RECT 6.360 0.610 6.620 0.870 ;
        RECT 8.460 -0.230 8.720 0.030 ;
      LAYER met2 ;
        RECT 1.570 0.870 1.890 0.920 ;
        RECT 2.600 0.880 2.920 0.890 ;
        RECT 2.600 0.870 2.930 0.880 ;
        RECT -0.740 0.670 -0.030 0.870 ;
        RECT 0.110 0.670 2.930 0.870 ;
        RECT 1.570 0.660 1.890 0.670 ;
        RECT 2.600 0.620 2.930 0.670 ;
        RECT 2.600 0.600 2.920 0.620 ;
        RECT 4.280 0.100 4.620 0.160 ;
        RECT 6.360 0.100 6.620 0.900 ;
        RECT 4.280 -0.120 6.720 0.100 ;
        RECT 8.430 -0.260 8.890 0.060 ;
  END
END sky130_hilas_StepUpDigital

MACRO sky130_hilas_VinjNOR3
  CLASS BLOCK ;
  FOREIGN sky130_hilas_VinjNOR3 ;
  ORIGIN 3.370 -1.440 ;
  SIZE 6.880 BY 1.640 ;
  OBS
      LAYER nwell ;
        RECT -3.360 1.440 0.080 3.080 ;
      LAYER li1 ;
        RECT -2.740 2.650 -2.570 2.790 ;
        RECT -2.010 2.670 -1.840 2.750 ;
        RECT -1.200 2.670 -1.030 2.750 ;
        RECT 0.340 2.710 0.510 2.830 ;
        RECT -2.740 2.480 -2.550 2.650 ;
        RECT -2.740 2.380 -2.570 2.480 ;
        RECT -2.010 2.100 -1.800 2.670 ;
        RECT -1.240 2.420 -1.030 2.670 ;
        RECT -0.640 2.490 -0.470 2.590 ;
        RECT 0.300 2.540 0.510 2.710 ;
        RECT 2.230 2.640 2.490 2.710 ;
        RECT 3.030 2.640 3.210 2.770 ;
        RECT 0.340 2.500 0.510 2.540 ;
        RECT -1.240 2.100 -1.070 2.420 ;
        RECT -0.670 2.320 -0.470 2.490 ;
        RECT -0.640 2.220 -0.470 2.320 ;
        RECT 0.900 2.460 1.770 2.630 ;
        RECT 2.230 2.460 3.210 2.640 ;
        RECT -3.170 2.000 -3.000 2.100 ;
        RECT -3.190 1.830 -3.000 2.000 ;
        RECT -3.170 1.770 -3.000 1.830 ;
        RECT -2.750 2.040 -2.580 2.100 ;
        RECT -2.750 1.770 -2.500 2.040 ;
        RECT -2.010 1.850 -1.760 2.100 ;
        RECT -2.740 1.750 -2.500 1.770 ;
        RECT -1.930 1.760 -1.760 1.850 ;
        RECT -1.280 1.850 -1.070 2.100 ;
        RECT 0.900 2.020 1.070 2.460 ;
        RECT 2.230 2.020 2.490 2.460 ;
        RECT 3.030 2.350 3.210 2.460 ;
        RECT -0.560 1.850 1.070 2.020 ;
        RECT 1.520 1.850 2.490 2.020 ;
        RECT 2.940 1.850 3.280 2.020 ;
        RECT -1.280 1.770 -1.110 1.850 ;
        RECT 0.210 1.810 0.380 1.850 ;
      LAYER mcon ;
        RECT -2.720 2.480 -2.550 2.650 ;
        RECT -2.710 1.800 -2.540 1.970 ;
        RECT 2.260 2.140 2.440 2.320 ;
      LAYER met1 ;
        RECT -2.750 2.700 -2.530 3.040 ;
        RECT -2.750 2.440 -2.520 2.700 ;
        RECT -3.280 1.760 -2.970 2.110 ;
        RECT -2.750 2.040 -2.530 2.440 ;
        RECT -0.730 2.280 -0.400 2.540 ;
        RECT 0.240 2.500 0.670 2.790 ;
        RECT -2.750 1.730 -2.500 2.040 ;
        RECT 0.110 1.750 0.500 2.020 ;
        RECT -2.750 1.530 -2.530 1.730 ;
        RECT 2.220 1.530 2.490 3.050 ;
        RECT 3.040 1.760 3.350 2.080 ;
      LAYER via ;
        RECT -3.250 1.790 -2.990 2.050 ;
        RECT -0.690 2.280 -0.430 2.540 ;
        RECT 0.300 2.530 0.560 2.790 ;
        RECT 0.170 1.750 0.430 2.010 ;
        RECT 3.070 1.790 3.330 2.050 ;
      LAYER met2 ;
        RECT -3.370 2.730 0.670 2.890 ;
        RECT -0.730 2.460 -0.400 2.540 ;
        RECT 0.250 2.500 0.670 2.730 ;
        RECT -1.000 2.440 -0.400 2.460 ;
        RECT -3.360 2.280 -0.400 2.440 ;
        RECT -3.280 1.950 -2.960 2.050 ;
        RECT -3.360 1.790 -2.960 1.950 ;
        RECT 0.130 1.930 0.500 2.010 ;
        RECT 0.130 1.920 1.160 1.930 ;
        RECT 3.040 1.920 3.350 2.080 ;
        RECT 0.130 1.750 3.510 1.920 ;
  END
END sky130_hilas_VinjNOR3

MACRO sky130_hilas_VinjDiodeProtect01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_VinjDiodeProtect01 ;
  ORIGIN 7.450 2.290 ;
  SIZE 28.590 BY 10.870 ;
  PIN OUTPUT 
    ANTENNADIFFAREA 58.900799 ;
    PORT
      LAYER met1 ;
        RECT 6.900 7.960 7.250 8.120 ;
        RECT 6.890 7.010 7.260 7.960 ;
        RECT 6.540 6.640 9.010 7.010 ;
        RECT 5.100 5.180 9.010 6.640 ;
        RECT -4.610 5.170 9.010 5.180 ;
        RECT -5.280 4.610 9.010 5.170 ;
        RECT -5.280 0.310 18.070 4.610 ;
        RECT -5.280 0.030 9.010 0.310 ;
        RECT 5.100 -1.520 9.010 0.030 ;
        RECT 5.080 -2.290 9.030 -1.520 ;
    END
  END OUTPUT 
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT -7.450 5.090 21.140 6.490 ;
        RECT -6.980 5.080 -6.050 5.090 ;
        RECT -6.730 3.970 -6.560 5.080 ;
    END
    PORT
      LAYER met1 ;
        RECT -7.010 5.840 -4.640 6.470 ;
        RECT 16.330 5.990 20.460 6.390 ;
        RECT 16.330 5.900 20.470 5.990 ;
        RECT -6.980 3.880 -6.030 5.840 ;
        RECT -5.280 5.820 -4.700 5.840 ;
        RECT 19.940 5.000 20.470 5.900 ;
        RECT -6.750 -1.790 -6.030 3.880 ;
      LAYER via ;
        RECT -6.790 5.990 -4.760 6.320 ;
        RECT 16.600 5.990 19.590 6.340 ;
        RECT -6.850 5.130 -6.150 5.750 ;
        RECT 20.030 5.190 20.380 5.950 ;
    END
  END VGND
  PIN VINJ
    ANTENNADIFFAREA 9.088799 ;
    PORT
      LAYER nwell ;
        RECT 7.420 -0.380 19.470 5.560 ;
      LAYER met2 ;
        RECT 18.890 0.190 19.530 3.200 ;
        RECT -7.450 -1.210 21.140 0.190 ;
        RECT 17.990 -1.340 20.620 -1.210 ;
        RECT 17.990 -1.850 20.540 -1.340 ;
        RECT 17.990 -1.920 18.610 -1.850 ;
    END
  END VINJ
  PIN INPUT
    PORT
      LAYER met1 ;
        RECT 0.260 7.990 4.160 8.580 ;
        RECT 0.260 6.640 0.550 7.990 ;
    END
  END INPUT
  OBS
      LAYER li1 ;
        RECT 0.280 6.640 0.530 8.100 ;
        RECT 0.320 6.630 0.490 6.640 ;
        RECT 6.960 6.610 7.210 8.090 ;
        RECT -6.900 5.890 20.480 6.400 ;
        RECT -6.900 3.960 -6.100 5.890 ;
        RECT -5.520 5.440 -5.350 5.520 ;
        RECT 5.720 5.440 5.950 5.530 ;
        RECT -5.520 5.430 5.950 5.440 ;
        RECT -6.900 -0.620 -6.390 3.960 ;
        RECT -5.530 -0.040 5.950 5.430 ;
        RECT -5.600 -0.210 5.950 -0.040 ;
        RECT -5.530 -0.270 -5.340 -0.210 ;
        RECT 5.720 -0.450 5.950 -0.210 ;
        RECT -5.650 -0.620 -3.850 -0.610 ;
        RECT 6.510 -0.620 7.020 5.890 ;
        RECT 7.780 5.000 19.030 5.170 ;
        RECT 7.780 0.130 7.950 5.000 ;
        RECT 8.340 4.670 18.450 4.690 ;
        RECT 8.340 4.630 18.470 4.670 ;
        RECT 8.290 4.460 18.470 4.630 ;
        RECT 8.340 0.440 18.470 4.460 ;
        RECT 18.860 3.240 19.030 5.000 ;
        RECT 8.340 0.360 18.450 0.440 ;
        RECT 7.770 0.060 7.950 0.130 ;
        RECT 18.860 0.060 19.470 3.240 ;
        RECT 7.770 -0.110 19.470 0.060 ;
        RECT 18.930 -0.220 19.470 -0.110 ;
        RECT 19.930 -0.460 20.480 5.890 ;
        RECT 19.920 -0.620 20.480 -0.460 ;
        RECT -6.900 -0.960 20.480 -0.620 ;
        RECT -6.870 -1.130 20.480 -0.960 ;
        RECT -6.870 -1.150 -6.180 -1.130 ;
        RECT -5.670 -1.140 -3.870 -1.130 ;
      LAYER mcon ;
        RECT 0.320 7.580 0.490 7.750 ;
        RECT 0.320 7.220 0.490 7.390 ;
        RECT 0.320 6.850 0.490 7.020 ;
        RECT 7.000 7.900 7.170 8.070 ;
        RECT 7.000 7.540 7.170 7.710 ;
        RECT 7.000 7.180 7.170 7.350 ;
        RECT 7.000 6.820 7.170 6.990 ;
        RECT -6.820 6.230 -4.960 6.240 ;
        RECT -6.820 6.060 -4.950 6.230 ;
        RECT 16.540 6.050 19.700 6.230 ;
        RECT -6.780 3.970 -6.600 5.870 ;
        RECT -6.380 3.960 -6.200 5.870 ;
        RECT -5.190 4.930 5.790 5.100 ;
        RECT -5.190 4.310 5.790 4.480 ;
        RECT -5.180 3.690 5.800 3.860 ;
        RECT -5.160 3.110 5.820 3.280 ;
        RECT -5.150 2.520 5.830 2.690 ;
        RECT -5.150 1.920 5.830 2.090 ;
        RECT -5.200 1.320 5.780 1.490 ;
        RECT -5.190 0.710 5.790 0.880 ;
        RECT -5.200 0.110 5.780 0.280 ;
        RECT 8.540 4.170 17.990 4.340 ;
        RECT 8.530 3.420 17.920 3.590 ;
        RECT 8.560 2.700 17.960 2.870 ;
        RECT 8.570 2.040 17.940 2.210 ;
        RECT 8.560 1.390 18.010 1.560 ;
        RECT 8.570 0.750 17.960 0.920 ;
        RECT 20.110 5.070 20.310 6.000 ;
        RECT 19.040 -0.170 19.390 3.130 ;
      LAYER met1 ;
        RECT 18.840 3.190 19.410 3.200 ;
        RECT 18.840 -0.230 19.460 3.190 ;
        RECT 18.840 -0.240 19.410 -0.230 ;
        RECT 18.010 -1.870 18.570 -1.370 ;
        RECT 18.020 -2.090 18.570 -1.870 ;
      LAYER via ;
        RECT 19.000 -0.100 19.420 3.070 ;
        RECT 18.030 -1.920 18.550 -1.400 ;
  END
END sky130_hilas_VinjDiodeProtect01

MACRO sky130_hilas_LevelShift4InputUp
  CLASS BLOCK ;
  FOREIGN sky130_hilas_LevelShift4InputUp ;
  ORIGIN 1.230 1.060 ;
  SIZE 10.585 BY 7.000 ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 6.070 -1.060 7.840 5.940 ;
      LAYER met1 ;
        RECT 7.360 -1.060 7.600 5.940 ;
    END
  END VPWR
  PIN VINJ
    ANTENNADIFFAREA 1.900800 ;
    PORT
      LAYER nwell ;
        RECT -0.300 -1.060 2.200 5.940 ;
      LAYER met1 ;
        RECT 0.040 -1.060 0.330 5.940 ;
    END
  END VINJ
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 4.350 -1.060 4.660 5.940 ;
    END
  END VGND
  PIN INPUT4
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 7.940 -0.570 8.540 -0.560 ;
        RECT 7.940 -0.880 9.355 -0.570 ;
    END
  END INPUT4
  PIN INPUT3
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 7.940 0.870 9.000 1.190 ;
    END
  END INPUT3
  PIN INPUT2
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 7.940 2.620 8.920 2.940 ;
    END
  END INPUT2
  PIN INPUT1
    ANTENNAGATEAREA 0.201600 ;
    PORT
      LAYER met2 ;
        RECT 7.940 4.370 8.650 4.690 ;
    END
  END INPUT1
  OBS
      LAYER li1 ;
        RECT 0.980 5.430 1.430 5.580 ;
        RECT 0.040 5.250 0.370 5.420 ;
        RECT 0.830 5.260 1.430 5.430 ;
        RECT 0.110 4.790 0.290 5.250 ;
        RECT 1.630 4.820 1.800 5.580 ;
        RECT 2.130 5.490 2.420 5.510 ;
        RECT 2.130 5.450 2.590 5.490 ;
        RECT 2.130 5.430 3.570 5.450 ;
        RECT 2.130 5.270 3.610 5.430 ;
        RECT 2.420 5.260 3.610 5.270 ;
        RECT 4.060 5.400 4.520 5.430 ;
        RECT 5.830 5.400 6.180 5.500 ;
        RECT 4.060 5.260 5.170 5.400 ;
        RECT 4.350 5.230 5.170 5.260 ;
        RECT 5.410 5.230 6.580 5.400 ;
        RECT 6.830 5.230 7.590 5.400 ;
        RECT 4.350 5.090 4.610 5.230 ;
        RECT 3.430 4.920 4.610 5.090 ;
        RECT 7.360 5.220 7.590 5.230 ;
        RECT 1.630 4.810 2.010 4.820 ;
        RECT 0.110 4.620 1.070 4.790 ;
        RECT 1.540 4.750 2.010 4.810 ;
        RECT 1.540 4.640 2.880 4.750 ;
        RECT 1.620 4.580 2.880 4.640 ;
        RECT 1.620 4.530 2.010 4.580 ;
        RECT 3.430 4.480 3.610 4.920 ;
        RECT 4.350 4.780 4.610 4.920 ;
        RECT 5.820 4.780 6.150 5.040 ;
        RECT 7.360 4.780 7.630 5.220 ;
        RECT 3.850 4.420 4.060 4.750 ;
        RECT 4.350 4.610 4.680 4.780 ;
        RECT 4.920 4.610 7.080 4.780 ;
        RECT 4.350 4.560 4.520 4.610 ;
        RECT 7.330 4.600 7.660 4.780 ;
        RECT 8.010 4.640 8.180 4.700 ;
        RECT 7.990 4.420 8.210 4.640 ;
        RECT 8.010 4.370 8.180 4.420 ;
        RECT 0.980 3.680 1.430 3.830 ;
        RECT 0.040 3.500 0.370 3.670 ;
        RECT 0.830 3.510 1.430 3.680 ;
        RECT 0.110 3.040 0.290 3.500 ;
        RECT 1.630 3.070 1.800 3.830 ;
        RECT 2.130 3.740 2.420 3.760 ;
        RECT 2.130 3.700 2.590 3.740 ;
        RECT 2.130 3.680 3.570 3.700 ;
        RECT 2.130 3.520 3.610 3.680 ;
        RECT 2.420 3.510 3.610 3.520 ;
        RECT 4.060 3.650 4.520 3.680 ;
        RECT 5.830 3.650 6.180 3.750 ;
        RECT 4.060 3.510 5.170 3.650 ;
        RECT 4.350 3.480 5.170 3.510 ;
        RECT 5.410 3.480 6.580 3.650 ;
        RECT 6.830 3.480 7.590 3.650 ;
        RECT 4.350 3.340 4.610 3.480 ;
        RECT 3.430 3.170 4.610 3.340 ;
        RECT 7.360 3.470 7.590 3.480 ;
        RECT 1.630 3.060 2.010 3.070 ;
        RECT 0.110 2.870 1.070 3.040 ;
        RECT 1.540 3.000 2.010 3.060 ;
        RECT 1.540 2.890 2.880 3.000 ;
        RECT 1.620 2.830 2.880 2.890 ;
        RECT 1.620 2.780 2.010 2.830 ;
        RECT 3.430 2.730 3.610 3.170 ;
        RECT 4.350 3.030 4.610 3.170 ;
        RECT 5.820 3.030 6.150 3.290 ;
        RECT 7.360 3.030 7.630 3.470 ;
        RECT 3.850 2.670 4.060 3.000 ;
        RECT 4.350 2.860 4.680 3.030 ;
        RECT 4.920 2.860 7.080 3.030 ;
        RECT 4.350 2.810 4.520 2.860 ;
        RECT 7.330 2.850 7.660 3.030 ;
        RECT 8.010 2.890 8.180 2.950 ;
        RECT 7.990 2.670 8.210 2.890 ;
        RECT 8.010 2.620 8.180 2.670 ;
        RECT 0.980 1.930 1.430 2.080 ;
        RECT 0.040 1.750 0.370 1.920 ;
        RECT 0.830 1.760 1.430 1.930 ;
        RECT 0.110 1.290 0.290 1.750 ;
        RECT 1.630 1.320 1.800 2.080 ;
        RECT 2.130 1.990 2.420 2.010 ;
        RECT 2.130 1.950 2.590 1.990 ;
        RECT 2.130 1.930 3.570 1.950 ;
        RECT 2.130 1.770 3.610 1.930 ;
        RECT 2.420 1.760 3.610 1.770 ;
        RECT 4.060 1.900 4.520 1.930 ;
        RECT 5.830 1.900 6.180 2.000 ;
        RECT 4.060 1.760 5.170 1.900 ;
        RECT 4.350 1.730 5.170 1.760 ;
        RECT 5.410 1.730 6.580 1.900 ;
        RECT 6.830 1.730 7.590 1.900 ;
        RECT 4.350 1.590 4.610 1.730 ;
        RECT 3.430 1.420 4.610 1.590 ;
        RECT 7.360 1.720 7.590 1.730 ;
        RECT 1.630 1.310 2.010 1.320 ;
        RECT 0.110 1.120 1.070 1.290 ;
        RECT 1.540 1.250 2.010 1.310 ;
        RECT 1.540 1.140 2.880 1.250 ;
        RECT 1.620 1.080 2.880 1.140 ;
        RECT 1.620 1.030 2.010 1.080 ;
        RECT 3.430 0.980 3.610 1.420 ;
        RECT 4.350 1.280 4.610 1.420 ;
        RECT 5.820 1.280 6.150 1.540 ;
        RECT 7.360 1.280 7.630 1.720 ;
        RECT 3.850 0.920 4.060 1.250 ;
        RECT 4.350 1.110 4.680 1.280 ;
        RECT 4.920 1.110 7.080 1.280 ;
        RECT 4.350 1.060 4.520 1.110 ;
        RECT 7.330 1.100 7.660 1.280 ;
        RECT 8.010 1.140 8.180 1.200 ;
        RECT 7.990 0.920 8.210 1.140 ;
        RECT 8.010 0.870 8.180 0.920 ;
        RECT 0.980 0.180 1.430 0.330 ;
        RECT 0.040 0.000 0.370 0.170 ;
        RECT 0.830 0.010 1.430 0.180 ;
        RECT 0.110 -0.460 0.290 0.000 ;
        RECT 1.630 -0.430 1.800 0.330 ;
        RECT 2.130 0.240 2.420 0.260 ;
        RECT 2.130 0.200 2.590 0.240 ;
        RECT 2.130 0.180 3.570 0.200 ;
        RECT 2.130 0.020 3.610 0.180 ;
        RECT 2.420 0.010 3.610 0.020 ;
        RECT 4.060 0.150 4.520 0.180 ;
        RECT 5.830 0.150 6.180 0.250 ;
        RECT 4.060 0.010 5.170 0.150 ;
        RECT 4.350 -0.020 5.170 0.010 ;
        RECT 5.410 -0.020 6.580 0.150 ;
        RECT 6.830 -0.020 7.590 0.150 ;
        RECT 4.350 -0.160 4.610 -0.020 ;
        RECT 3.430 -0.330 4.610 -0.160 ;
        RECT 7.360 -0.030 7.590 -0.020 ;
        RECT 1.630 -0.440 2.010 -0.430 ;
        RECT 0.110 -0.630 1.070 -0.460 ;
        RECT 1.540 -0.500 2.010 -0.440 ;
        RECT 1.540 -0.610 2.880 -0.500 ;
        RECT 1.620 -0.670 2.880 -0.610 ;
        RECT 1.620 -0.720 2.010 -0.670 ;
        RECT 3.430 -0.770 3.610 -0.330 ;
        RECT 4.350 -0.470 4.610 -0.330 ;
        RECT 5.820 -0.470 6.150 -0.210 ;
        RECT 7.360 -0.470 7.630 -0.030 ;
        RECT 3.850 -0.830 4.060 -0.500 ;
        RECT 4.350 -0.640 4.680 -0.470 ;
        RECT 4.920 -0.640 7.080 -0.470 ;
        RECT 4.350 -0.690 4.520 -0.640 ;
        RECT 7.330 -0.650 7.660 -0.470 ;
        RECT 8.010 -0.610 8.180 -0.550 ;
        RECT 7.990 -0.830 8.210 -0.610 ;
        RECT 8.010 -0.880 8.180 -0.830 ;
      LAYER mcon ;
        RECT 1.150 5.330 1.320 5.500 ;
        RECT 0.110 4.990 0.280 5.160 ;
        RECT 2.190 5.290 2.360 5.460 ;
        RECT 5.890 5.270 6.100 5.480 ;
        RECT 0.110 4.630 0.280 4.800 ;
        RECT 7.400 4.900 7.570 5.070 ;
        RECT 1.150 3.580 1.320 3.750 ;
        RECT 0.110 3.240 0.280 3.410 ;
        RECT 2.190 3.540 2.360 3.710 ;
        RECT 5.890 3.520 6.100 3.730 ;
        RECT 0.110 2.880 0.280 3.050 ;
        RECT 7.400 3.150 7.570 3.320 ;
        RECT 1.150 1.830 1.320 2.000 ;
        RECT 0.110 1.490 0.280 1.660 ;
        RECT 2.190 1.790 2.360 1.960 ;
        RECT 5.890 1.770 6.100 1.980 ;
        RECT 0.110 1.130 0.280 1.300 ;
        RECT 7.400 1.400 7.570 1.570 ;
        RECT 1.150 0.080 1.320 0.250 ;
        RECT 0.110 -0.260 0.280 -0.090 ;
        RECT 2.190 0.040 2.360 0.210 ;
        RECT 5.890 0.020 6.100 0.230 ;
        RECT 0.110 -0.620 0.280 -0.450 ;
        RECT 7.400 -0.350 7.570 -0.180 ;
      LAYER met1 ;
        RECT 1.080 5.280 1.400 5.580 ;
        RECT 2.130 5.510 2.440 5.520 ;
        RECT 2.120 5.240 2.440 5.510 ;
        RECT 2.130 5.230 2.420 5.240 ;
        RECT 5.830 5.230 6.180 5.520 ;
        RECT 5.980 5.210 6.180 5.230 ;
        RECT 3.820 4.480 4.100 4.810 ;
        RECT 7.930 4.370 8.340 4.700 ;
        RECT 1.080 3.530 1.400 3.830 ;
        RECT 2.130 3.760 2.440 3.770 ;
        RECT 2.120 3.490 2.440 3.760 ;
        RECT 2.130 3.480 2.420 3.490 ;
        RECT 5.830 3.480 6.180 3.770 ;
        RECT 5.980 3.460 6.180 3.480 ;
        RECT 3.820 2.730 4.100 3.060 ;
        RECT 7.930 2.620 8.340 2.950 ;
        RECT 1.080 1.780 1.400 2.080 ;
        RECT 2.130 2.010 2.440 2.020 ;
        RECT 2.120 1.740 2.440 2.010 ;
        RECT 2.130 1.730 2.420 1.740 ;
        RECT 5.830 1.730 6.180 2.020 ;
        RECT 5.980 1.710 6.180 1.730 ;
        RECT 3.820 0.980 4.100 1.310 ;
        RECT 7.930 0.870 8.340 1.200 ;
        RECT 1.080 0.030 1.400 0.330 ;
        RECT 2.130 0.260 2.440 0.270 ;
        RECT 2.120 -0.010 2.440 0.260 ;
        RECT 2.130 -0.020 2.420 -0.010 ;
        RECT 5.830 -0.020 6.180 0.270 ;
        RECT 5.980 -0.040 6.180 -0.020 ;
        RECT 3.820 -0.770 4.100 -0.440 ;
        RECT 7.930 -0.880 8.340 -0.550 ;
      LAYER via ;
        RECT 1.110 5.290 1.370 5.550 ;
        RECT 2.150 5.250 2.410 5.510 ;
        RECT 5.870 5.240 6.130 5.500 ;
        RECT 3.830 4.520 4.090 4.780 ;
        RECT 7.970 4.400 8.230 4.660 ;
        RECT 1.110 3.540 1.370 3.800 ;
        RECT 2.150 3.500 2.410 3.760 ;
        RECT 5.870 3.490 6.130 3.750 ;
        RECT 3.830 2.770 4.090 3.030 ;
        RECT 7.970 2.650 8.230 2.910 ;
        RECT 1.110 1.790 1.370 2.050 ;
        RECT 2.150 1.750 2.410 2.010 ;
        RECT 5.870 1.740 6.130 2.000 ;
        RECT 3.830 1.020 4.090 1.280 ;
        RECT 7.970 0.900 8.230 1.160 ;
        RECT 1.110 0.040 1.370 0.300 ;
        RECT 2.150 0.000 2.410 0.260 ;
        RECT 5.870 -0.010 6.130 0.250 ;
        RECT 3.830 -0.730 4.090 -0.470 ;
        RECT 7.970 -0.850 8.230 -0.590 ;
      LAYER met2 ;
        RECT 1.080 5.500 1.400 5.550 ;
        RECT 2.110 5.510 2.430 5.520 ;
        RECT 2.110 5.500 2.440 5.510 ;
        RECT -1.230 5.300 -0.520 5.500 ;
        RECT -0.380 5.300 2.440 5.500 ;
        RECT 1.080 5.290 1.400 5.300 ;
        RECT 2.110 5.250 2.440 5.300 ;
        RECT 2.110 5.230 2.430 5.250 ;
        RECT 3.790 4.730 4.130 4.790 ;
        RECT 5.870 4.730 6.130 5.530 ;
        RECT 3.790 4.510 6.230 4.730 ;
        RECT 1.080 3.750 1.400 3.800 ;
        RECT 2.110 3.760 2.430 3.770 ;
        RECT 2.110 3.750 2.440 3.760 ;
        RECT -1.230 3.550 -0.520 3.750 ;
        RECT -0.380 3.550 2.440 3.750 ;
        RECT 1.080 3.540 1.400 3.550 ;
        RECT 2.110 3.500 2.440 3.550 ;
        RECT 2.110 3.480 2.430 3.500 ;
        RECT 3.790 2.980 4.130 3.040 ;
        RECT 5.870 2.980 6.130 3.780 ;
        RECT 3.790 2.760 6.230 2.980 ;
        RECT 1.080 2.000 1.400 2.050 ;
        RECT 2.110 2.010 2.430 2.020 ;
        RECT 2.110 2.000 2.440 2.010 ;
        RECT -1.230 1.800 -0.520 2.000 ;
        RECT -0.380 1.800 2.440 2.000 ;
        RECT 1.080 1.790 1.400 1.800 ;
        RECT 2.110 1.750 2.440 1.800 ;
        RECT 2.110 1.730 2.430 1.750 ;
        RECT 3.790 1.230 4.130 1.290 ;
        RECT 5.870 1.230 6.130 2.030 ;
        RECT 3.790 1.010 6.230 1.230 ;
        RECT 1.080 0.250 1.400 0.300 ;
        RECT 2.110 0.260 2.430 0.270 ;
        RECT 2.110 0.250 2.440 0.260 ;
        RECT -1.230 0.050 -0.520 0.250 ;
        RECT -0.380 0.050 2.440 0.250 ;
        RECT 1.080 0.040 1.400 0.050 ;
        RECT 2.110 0.000 2.440 0.050 ;
        RECT 2.110 -0.020 2.430 0.000 ;
        RECT 3.790 -0.520 4.130 -0.460 ;
        RECT 5.870 -0.520 6.130 0.280 ;
        RECT 3.790 -0.740 6.230 -0.520 ;
  END
END sky130_hilas_LevelShift4InputUp

MACRO sky130_hilas_WTA4Stage01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_WTA4Stage01 ;
  ORIGIN 11.210 0.610 ;
  SIZE 14.170 BY 6.500 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 2.510 1.160 2.840 1.250 ;
        RECT -7.420 1.090 -7.100 1.150 ;
        RECT -3.840 1.090 2.840 1.160 ;
        RECT -7.420 0.990 2.840 1.090 ;
        RECT -7.420 0.920 -3.070 0.990 ;
        RECT 2.510 0.960 2.840 0.990 ;
        RECT -7.420 0.870 -7.100 0.920 ;
        RECT -3.400 0.860 -3.070 0.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.570 1.270 2.800 5.620 ;
        RECT 2.530 1.260 2.810 1.270 ;
        RECT 2.530 0.940 2.830 1.260 ;
        RECT 2.570 -0.430 2.800 0.940 ;
      LAYER via ;
        RECT 2.540 0.970 2.810 1.240 ;
    END
  END VGND
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT -8.450 4.900 -8.140 4.920 ;
        RECT -0.650 4.900 -0.510 4.910 ;
        RECT -10.610 4.720 -0.500 4.900 ;
        RECT -8.450 4.710 -0.500 4.720 ;
        RECT -8.450 4.590 -8.140 4.710 ;
        RECT -0.650 4.570 -0.500 4.710 ;
        RECT -0.650 4.480 0.560 4.570 ;
        RECT -0.650 4.420 0.690 4.480 ;
        RECT -0.650 4.370 2.960 4.420 ;
        RECT 0.380 4.260 2.960 4.370 ;
        RECT 0.380 4.150 0.690 4.260 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT -8.450 3.810 -8.140 3.940 ;
        RECT -10.610 3.630 0.660 3.810 ;
        RECT -8.450 3.610 -8.140 3.630 ;
        RECT 0.380 3.600 0.660 3.630 ;
        RECT 0.380 3.490 0.690 3.600 ;
        RECT 0.380 3.330 2.960 3.490 ;
        RECT 0.380 3.270 0.690 3.330 ;
    END
  END OUTPUT2
  PIN OUTPUT3
    USE ANALOG ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT 0.380 1.680 0.690 1.710 ;
        RECT -1.010 1.650 0.690 1.680 ;
        RECT -1.010 1.520 2.960 1.650 ;
        RECT -1.010 1.510 -0.550 1.520 ;
        RECT 0.380 1.490 2.960 1.520 ;
        RECT 0.380 1.380 0.690 1.490 ;
    END
  END OUTPUT3
  PIN OUTPUT4
    USE ANALOG ;
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 0.380 0.720 0.690 0.830 ;
        RECT 0.380 0.710 2.960 0.720 ;
        RECT -0.550 0.700 2.960 0.710 ;
        RECT -8.170 0.690 2.960 0.700 ;
        RECT -8.450 0.560 2.960 0.690 ;
        RECT -10.610 0.530 0.690 0.560 ;
        RECT -10.610 0.380 -8.050 0.530 ;
        RECT 0.380 0.500 0.690 0.530 ;
        RECT -8.450 0.360 -8.140 0.380 ;
    END
  END OUTPUT4
  PIN INPUT1
    USE ANALOG ;
    ANTENNAGATEAREA 0.118000 ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT -7.850 5.310 -7.530 5.330 ;
        RECT -7.850 5.120 0.070 5.310 ;
        RECT 0.230 5.120 0.540 5.160 ;
        RECT -7.850 5.100 0.540 5.120 ;
        RECT -7.850 5.070 -7.530 5.100 ;
        RECT -0.140 4.910 0.540 5.100 ;
        RECT 0.230 4.830 0.540 4.910 ;
        RECT -11.120 4.270 -10.970 4.690 ;
        RECT -7.870 4.270 -7.550 4.280 ;
        RECT -11.120 4.120 -7.550 4.270 ;
        RECT -7.990 4.020 -7.550 4.120 ;
    END
  END INPUT1
  PIN INPUT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.118000 ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT -11.140 3.520 -10.820 3.790 ;
        RECT -7.910 3.040 -7.680 3.050 ;
        RECT -7.910 3.010 -0.340 3.040 ;
        RECT -7.910 2.840 -0.280 3.010 ;
        RECT 0.230 2.840 0.540 2.920 ;
        RECT -11.160 2.740 -10.840 2.770 ;
        RECT -7.910 2.740 -7.670 2.840 ;
        RECT -11.160 2.560 -7.670 2.740 ;
        RECT -0.470 2.640 0.540 2.840 ;
        RECT 0.130 2.630 0.540 2.640 ;
        RECT 0.230 2.590 0.540 2.630 ;
        RECT -11.160 2.540 -7.750 2.560 ;
        RECT -11.160 2.510 -10.840 2.540 ;
    END
  END INPUT2
  PIN INPUT3
    USE ANALOG ;
    ANTENNAGATEAREA 0.118000 ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT -7.870 2.360 -7.550 2.400 ;
        RECT -7.870 2.340 -0.320 2.360 ;
        RECT 0.230 2.350 0.540 2.390 ;
        RECT 0.130 2.340 0.540 2.350 ;
        RECT -7.870 2.140 0.540 2.340 ;
        RECT -7.770 2.130 -7.450 2.140 ;
        RECT 0.230 2.060 0.540 2.140 ;
        RECT -11.180 1.180 -10.980 1.680 ;
        RECT -8.000 1.180 -7.680 1.220 ;
        RECT -11.180 0.980 -7.630 1.180 ;
        RECT -8.000 0.960 -7.680 0.980 ;
    END
  END INPUT3
  PIN INPUT4
    USE ANALOG ;
    ANTENNAGATEAREA 0.118000 ;
    ANTENNADIFFAREA 0.171100 ;
    PORT
      LAYER met2 ;
        RECT -11.210 0.440 -10.900 0.770 ;
        RECT 0.230 0.090 0.540 0.150 ;
        RECT -0.320 0.080 0.540 0.090 ;
        RECT -7.900 -0.140 0.540 0.080 ;
        RECT -7.900 -0.150 -0.310 -0.140 ;
        RECT -7.900 -0.160 -7.130 -0.150 ;
        RECT -11.160 -0.200 -10.850 -0.190 ;
        RECT -11.160 -0.330 -10.800 -0.200 ;
        RECT -7.900 -0.330 -7.660 -0.160 ;
        RECT 0.230 -0.180 0.540 -0.140 ;
        RECT -11.160 -0.520 -7.660 -0.330 ;
        RECT -11.030 -0.570 -7.660 -0.520 ;
    END
  END INPUT4
  PIN DRAIN1
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT -8.450 5.330 -8.140 5.470 ;
        RECT -11.160 5.150 -8.140 5.330 ;
        RECT -8.450 5.140 -8.140 5.150 ;
    END
  END DRAIN1
  PIN GATE1
    ANTENNADIFFAREA 3.253900 ;
    PORT
      LAYER nwell ;
        RECT -6.520 -0.610 -4.290 5.880 ;
      LAYER met1 ;
        RECT -5.320 3.700 -4.940 5.890 ;
        RECT -5.320 1.840 -4.930 3.700 ;
        RECT -5.320 -0.610 -4.940 1.840 ;
    END
  END GATE1
  PIN VTUN
    ANTENNADIFFAREA 2.243500 ;
    PORT
      LAYER nwell ;
        RECT -2.270 -0.610 -0.540 5.890 ;
      LAYER met1 ;
        RECT -1.290 -0.610 -0.890 5.890 ;
    END
  END VTUN
  PIN WTAMIDDLENODE
    ANTENNAGATEAREA 0.472000 ;
    ANTENNADIFFAREA 0.708000 ;
    PORT
      LAYER met1 ;
        RECT 1.310 -0.430 1.540 5.620 ;
    END
  END WTAMIDDLENODE
  PIN COLSEL1
    ANTENNAGATEAREA 0.720000 ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met1 ;
        RECT -9.840 4.840 -9.650 5.830 ;
        RECT -9.440 5.150 -9.280 5.880 ;
        RECT -9.480 5.130 -9.280 5.150 ;
        RECT -9.490 4.890 -9.260 5.130 ;
        RECT -9.490 4.840 -9.280 4.890 ;
        RECT -9.840 4.720 -9.670 4.840 ;
        RECT -9.840 3.810 -9.680 4.720 ;
        RECT -9.840 3.690 -9.670 3.810 ;
        RECT -9.440 3.690 -9.280 4.840 ;
        RECT -9.840 2.770 -9.650 3.690 ;
        RECT -9.490 3.640 -9.280 3.690 ;
        RECT -9.490 3.400 -9.260 3.640 ;
        RECT -9.480 3.380 -9.280 3.400 ;
        RECT -9.870 2.740 -9.630 2.770 ;
        RECT -9.440 2.740 -9.280 3.380 ;
        RECT -9.870 2.570 -9.280 2.740 ;
        RECT -9.870 2.540 -9.630 2.570 ;
        RECT -9.840 1.600 -9.650 2.540 ;
        RECT -9.440 1.910 -9.280 2.570 ;
        RECT -9.480 1.890 -9.280 1.910 ;
        RECT -9.490 1.650 -9.260 1.890 ;
        RECT -9.490 1.600 -9.280 1.650 ;
        RECT -9.840 1.480 -9.670 1.600 ;
        RECT -9.840 0.560 -9.680 1.480 ;
        RECT -9.840 0.440 -9.670 0.560 ;
        RECT -9.440 0.440 -9.280 1.600 ;
        RECT -9.840 -0.550 -9.650 0.440 ;
        RECT -9.490 0.390 -9.280 0.440 ;
        RECT -9.490 0.150 -9.260 0.390 ;
        RECT -9.480 0.130 -9.280 0.150 ;
        RECT -9.440 -0.600 -9.280 0.130 ;
    END
  END COLSEL1
  PIN VINJ
    ANTENNADIFFAREA 1.088000 ;
    PORT
      LAYER nwell ;
        RECT -10.610 5.620 -8.050 5.890 ;
        RECT -11.010 3.690 -8.050 5.620 ;
        RECT -11.120 2.540 -8.050 3.690 ;
        RECT -11.010 -0.420 -8.050 2.540 ;
        RECT -10.610 -0.610 -8.050 -0.420 ;
      LAYER met1 ;
        RECT -10.250 5.180 -10.090 5.880 ;
        RECT -10.250 4.630 -9.980 5.180 ;
        RECT -10.260 4.580 -9.980 4.630 ;
        RECT -10.260 4.490 -10.090 4.580 ;
        RECT -10.250 4.040 -10.090 4.490 ;
        RECT -10.260 3.950 -10.090 4.040 ;
        RECT -10.260 3.900 -9.980 3.950 ;
        RECT -10.250 3.350 -9.980 3.900 ;
        RECT -10.250 1.940 -10.090 3.350 ;
        RECT -10.250 1.390 -9.980 1.940 ;
        RECT -10.260 1.340 -9.980 1.390 ;
        RECT -10.260 1.250 -10.090 1.340 ;
        RECT -10.250 0.790 -10.090 1.250 ;
        RECT -10.260 0.700 -10.090 0.790 ;
        RECT -10.260 0.650 -9.980 0.700 ;
        RECT -10.250 0.100 -9.980 0.650 ;
        RECT -10.250 -0.600 -10.090 0.100 ;
    END
  END VINJ
  PIN DRAIN2
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT -8.450 3.380 -8.140 3.390 ;
        RECT -11.190 3.220 -8.140 3.380 ;
        RECT -11.190 3.200 -8.050 3.220 ;
        RECT -8.450 3.080 -8.050 3.200 ;
        RECT -8.450 3.060 -8.140 3.080 ;
    END
  END DRAIN2
  PIN DRAIN3
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT -8.450 2.100 -8.140 2.230 ;
        RECT -8.450 2.090 -8.020 2.100 ;
        RECT -11.160 1.930 -8.020 2.090 ;
        RECT -11.160 1.910 -8.140 1.930 ;
        RECT -8.450 1.900 -8.140 1.910 ;
    END
  END DRAIN3
  PIN DRAIN4
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT -8.450 0.130 -8.140 0.140 ;
        RECT -11.180 -0.050 -8.140 0.130 ;
        RECT -8.450 -0.190 -8.140 -0.050 ;
    END
  END DRAIN4
  OBS
      LAYER li1 ;
        RECT -10.210 5.150 -10.010 5.500 ;
        RECT -8.470 5.420 -8.150 5.430 ;
        RECT -8.730 5.250 -8.150 5.420 ;
        RECT -8.480 5.200 -8.150 5.250 ;
        RECT -8.470 5.170 -8.150 5.200 ;
        RECT -10.220 5.120 -10.010 5.150 ;
        RECT -10.220 4.530 -10.000 5.120 ;
        RECT -9.480 4.530 -9.280 5.130 ;
        RECT 0.240 5.100 0.560 5.130 ;
        RECT 0.240 4.930 2.030 5.100 ;
        RECT 0.240 4.910 0.570 4.930 ;
        RECT -8.470 4.840 -8.150 4.880 ;
        RECT 0.240 4.870 0.560 4.910 ;
        RECT -8.480 4.800 -8.150 4.840 ;
        RECT -8.730 4.630 -8.150 4.800 ;
        RECT 1.860 4.700 2.030 4.930 ;
        RECT -8.470 4.620 -8.150 4.630 ;
        RECT 0.710 4.450 1.050 4.700 ;
        RECT 1.220 4.530 1.550 4.700 ;
        RECT 1.770 4.530 2.110 4.700 ;
        RECT -10.220 3.410 -10.000 4.000 ;
        RECT -10.220 3.380 -10.010 3.410 ;
        RECT -9.480 3.400 -9.280 4.000 ;
        RECT -8.470 3.900 -8.150 3.910 ;
        RECT -8.730 3.730 -8.150 3.900 ;
        RECT -7.340 3.840 -7.170 4.370 ;
        RECT -3.320 3.870 -3.150 4.400 ;
        RECT 0.390 4.190 1.050 4.450 ;
        RECT 1.300 4.360 1.470 4.530 ;
        RECT 1.860 4.360 2.030 4.530 ;
        RECT 1.220 4.190 1.550 4.360 ;
        RECT 1.770 4.190 2.110 4.360 ;
        RECT 1.300 3.960 1.550 4.190 ;
        RECT 2.430 4.110 2.940 4.780 ;
        RECT -8.480 3.690 -8.150 3.730 ;
        RECT -8.470 3.650 -8.150 3.690 ;
        RECT 1.300 3.790 1.970 3.960 ;
        RECT 1.300 3.560 1.550 3.790 ;
        RECT -10.210 3.030 -10.010 3.380 ;
        RECT -8.470 3.330 -8.150 3.360 ;
        RECT -8.480 3.280 -8.150 3.330 ;
        RECT 0.390 3.300 1.050 3.560 ;
        RECT 1.220 3.390 1.550 3.560 ;
        RECT 1.770 3.390 2.110 3.560 ;
        RECT -8.730 3.110 -8.150 3.280 ;
        RECT -8.470 3.100 -8.150 3.110 ;
        RECT -9.840 2.570 -9.400 2.740 ;
        RECT -10.210 1.910 -10.010 2.260 ;
        RECT -8.470 2.180 -8.150 2.190 ;
        RECT -8.730 2.010 -8.150 2.180 ;
        RECT -8.480 1.960 -8.150 2.010 ;
        RECT -7.350 1.980 -7.180 3.170 ;
        RECT -5.540 2.300 -4.990 2.730 ;
        RECT -8.470 1.930 -8.150 1.960 ;
        RECT -3.330 1.940 -3.160 3.110 ;
        RECT 0.710 3.050 1.050 3.300 ;
        RECT 1.300 3.220 1.470 3.390 ;
        RECT 1.860 3.220 2.030 3.390 ;
        RECT 1.220 3.050 1.550 3.220 ;
        RECT 1.770 3.050 2.110 3.220 ;
        RECT 0.240 2.840 0.560 2.880 ;
        RECT 0.240 2.820 0.570 2.840 ;
        RECT 1.860 2.820 2.030 3.050 ;
        RECT 2.430 2.970 2.940 3.640 ;
        RECT -1.510 2.370 -0.960 2.800 ;
        RECT 0.240 2.650 2.030 2.820 ;
        RECT 0.240 2.620 0.560 2.650 ;
        RECT 0.240 2.330 0.560 2.360 ;
        RECT 0.240 2.160 2.030 2.330 ;
        RECT 0.240 2.140 0.570 2.160 ;
        RECT 0.240 2.100 0.560 2.140 ;
        RECT 1.860 1.930 2.030 2.160 ;
        RECT -10.220 1.880 -10.010 1.910 ;
        RECT -10.220 1.290 -10.000 1.880 ;
        RECT -9.480 1.290 -9.280 1.890 ;
        RECT 0.710 1.680 1.050 1.930 ;
        RECT 1.220 1.760 1.550 1.930 ;
        RECT 1.770 1.760 2.110 1.930 ;
        RECT -8.470 1.600 -8.150 1.640 ;
        RECT -8.480 1.560 -8.150 1.600 ;
        RECT -8.730 1.390 -8.150 1.560 ;
        RECT 0.390 1.420 1.050 1.680 ;
        RECT 1.300 1.590 1.470 1.760 ;
        RECT 1.860 1.590 2.030 1.760 ;
        RECT 1.220 1.420 1.550 1.590 ;
        RECT 1.770 1.420 2.110 1.590 ;
        RECT -8.470 1.380 -8.150 1.390 ;
        RECT 1.300 1.190 1.550 1.420 ;
        RECT 2.430 1.340 2.940 2.010 ;
        RECT 1.300 1.020 1.970 1.190 ;
        RECT 1.300 0.790 1.550 1.020 ;
        RECT -11.200 0.690 -10.880 0.730 ;
        RECT -11.200 0.500 -10.870 0.690 ;
        RECT -11.200 0.470 -10.880 0.500 ;
        RECT -11.150 -0.230 -10.970 0.470 ;
        RECT -10.220 0.160 -10.000 0.750 ;
        RECT -10.220 0.130 -10.010 0.160 ;
        RECT -9.480 0.150 -9.280 0.750 ;
        RECT -8.470 0.650 -8.150 0.660 ;
        RECT -8.730 0.480 -8.150 0.650 ;
        RECT 0.390 0.530 1.050 0.790 ;
        RECT 1.220 0.620 1.550 0.790 ;
        RECT 1.770 0.620 2.110 0.790 ;
        RECT -8.480 0.440 -8.150 0.480 ;
        RECT -8.470 0.400 -8.150 0.440 ;
        RECT 0.710 0.280 1.050 0.530 ;
        RECT 1.300 0.450 1.470 0.620 ;
        RECT 1.860 0.450 2.030 0.620 ;
        RECT 1.220 0.280 1.550 0.450 ;
        RECT 1.770 0.280 2.110 0.450 ;
        RECT -10.210 -0.220 -10.010 0.130 ;
        RECT -8.470 0.080 -8.150 0.110 ;
        RECT -8.480 0.030 -8.150 0.080 ;
        RECT -8.730 -0.140 -8.150 0.030 ;
        RECT -8.470 -0.150 -8.150 -0.140 ;
        RECT 0.240 0.070 0.560 0.110 ;
        RECT 0.240 0.050 0.570 0.070 ;
        RECT 1.860 0.050 2.030 0.280 ;
        RECT 2.430 0.200 2.940 0.870 ;
        RECT 0.240 -0.120 2.030 0.050 ;
        RECT 0.240 -0.150 0.560 -0.120 ;
        RECT -11.150 -0.270 -10.830 -0.230 ;
        RECT -11.150 -0.460 -10.820 -0.270 ;
        RECT -11.150 -0.490 -10.830 -0.460 ;
      LAYER mcon ;
        RECT -8.380 5.210 -8.210 5.380 ;
        RECT -10.190 4.950 -10.020 5.120 ;
        RECT -9.460 4.920 -9.290 5.090 ;
        RECT 0.300 4.920 0.470 5.090 ;
        RECT -8.380 4.660 -8.210 4.830 ;
        RECT -7.340 4.200 -7.170 4.370 ;
        RECT -10.190 3.410 -10.020 3.580 ;
        RECT -8.380 3.700 -8.210 3.870 ;
        RECT -3.320 4.230 -3.150 4.400 ;
        RECT 0.450 4.240 0.620 4.410 ;
        RECT 2.600 4.360 2.770 4.530 ;
        RECT 1.340 3.790 1.510 3.960 ;
        RECT -9.460 3.440 -9.290 3.610 ;
        RECT -8.380 3.150 -8.210 3.320 ;
        RECT 0.450 3.340 0.620 3.510 ;
        RECT -7.350 3.000 -7.180 3.170 ;
        RECT -3.330 2.940 -3.160 3.110 ;
        RECT 2.600 3.220 2.770 3.390 ;
        RECT -7.350 2.340 -7.180 2.510 ;
        RECT -8.380 1.970 -8.210 2.140 ;
        RECT -5.260 2.380 -4.990 2.650 ;
        RECT -3.330 2.300 -3.160 2.470 ;
        RECT -1.230 2.450 -0.960 2.720 ;
        RECT 0.300 2.660 0.470 2.830 ;
        RECT 0.300 2.150 0.470 2.320 ;
        RECT -10.190 1.710 -10.020 1.880 ;
        RECT -9.460 1.680 -9.290 1.850 ;
        RECT -8.380 1.420 -8.210 1.590 ;
        RECT 0.450 1.470 0.620 1.640 ;
        RECT 2.600 1.590 2.770 1.760 ;
        RECT 1.340 1.020 1.510 1.190 ;
        RECT -11.140 0.510 -10.970 0.680 ;
        RECT -10.190 0.160 -10.020 0.330 ;
        RECT -8.380 0.450 -8.210 0.620 ;
        RECT 0.450 0.570 0.620 0.740 ;
        RECT -9.460 0.190 -9.290 0.360 ;
        RECT 2.600 0.450 2.770 0.620 ;
        RECT -8.380 -0.100 -8.210 0.070 ;
        RECT 0.300 -0.110 0.470 0.060 ;
        RECT -11.090 -0.450 -10.920 -0.280 ;
      LAYER met1 ;
        RECT -8.460 5.140 -8.140 5.460 ;
        RECT -7.820 5.040 -7.560 5.360 ;
        RECT -8.460 4.590 -8.140 4.910 ;
        RECT -7.820 4.310 -7.610 5.040 ;
        RECT -7.840 3.990 -7.580 4.310 ;
        RECT -11.110 3.690 -10.850 3.810 ;
        RECT -11.120 3.490 -10.850 3.690 ;
        RECT -8.460 3.620 -8.140 3.940 ;
        RECT -11.120 2.800 -10.910 3.490 ;
        RECT -8.460 3.070 -8.140 3.390 ;
        RECT -11.130 2.480 -10.870 2.800 ;
        RECT -8.460 1.900 -8.140 2.220 ;
        RECT -7.840 2.110 -7.580 2.430 ;
        RECT -8.460 1.350 -8.140 1.670 ;
        RECT -7.840 1.250 -7.680 2.110 ;
        RECT -7.970 0.930 -7.680 1.250 ;
        RECT -7.380 1.180 -7.130 5.890 ;
        RECT -7.400 1.150 -7.120 1.180 ;
        RECT -3.370 1.150 -3.100 5.890 ;
        RECT 0.230 4.840 0.550 5.160 ;
        RECT 0.380 4.160 0.700 4.480 ;
        RECT 0.380 3.270 0.700 3.590 ;
        RECT 0.230 2.590 0.550 2.910 ;
        RECT 0.230 2.070 0.550 2.390 ;
        RECT 0.380 1.390 0.700 1.710 ;
        RECT -7.410 0.870 -7.110 1.150 ;
        RECT -7.400 0.850 -7.120 0.870 ;
        RECT -11.210 0.440 -10.890 0.760 ;
        RECT -8.460 0.370 -8.140 0.690 ;
        RECT -8.460 -0.180 -8.140 0.140 ;
        RECT -11.160 -0.520 -10.840 -0.200 ;
        RECT -7.380 -0.610 -7.130 0.850 ;
        RECT -3.390 0.840 -3.080 1.150 ;
        RECT -3.370 -0.610 -3.100 0.840 ;
        RECT 0.380 0.500 0.700 0.820 ;
        RECT 0.230 -0.180 0.550 0.140 ;
      LAYER via ;
        RECT -8.430 5.170 -8.170 5.430 ;
        RECT -7.820 5.070 -7.560 5.330 ;
        RECT -8.430 4.620 -8.170 4.880 ;
        RECT -7.840 4.020 -7.580 4.280 ;
        RECT -11.110 3.520 -10.850 3.780 ;
        RECT -8.430 3.650 -8.170 3.910 ;
        RECT -8.430 3.100 -8.170 3.360 ;
        RECT -11.130 2.510 -10.870 2.770 ;
        RECT -8.430 1.930 -8.170 2.190 ;
        RECT -7.840 2.140 -7.580 2.400 ;
        RECT -8.430 1.380 -8.170 1.640 ;
        RECT -7.970 0.960 -7.710 1.220 ;
        RECT 0.260 4.870 0.520 5.130 ;
        RECT 0.410 4.190 0.670 4.450 ;
        RECT 0.410 3.300 0.670 3.560 ;
        RECT 0.260 2.620 0.520 2.880 ;
        RECT 0.260 2.100 0.520 2.360 ;
        RECT 0.410 1.420 0.670 1.680 ;
        RECT -7.390 0.880 -7.130 1.140 ;
        RECT -3.370 0.860 -3.100 1.120 ;
        RECT -11.180 0.470 -10.920 0.730 ;
        RECT -8.430 0.400 -8.170 0.660 ;
        RECT -8.430 -0.150 -8.170 0.110 ;
        RECT -11.130 -0.490 -10.870 -0.230 ;
        RECT 0.410 0.530 0.670 0.790 ;
        RECT 0.260 -0.150 0.520 0.110 ;
      LAYER met2 ;
        RECT -8.450 1.660 -8.140 1.680 ;
        RECT -10.610 1.490 -1.310 1.660 ;
        RECT -10.610 1.480 -8.050 1.490 ;
        RECT -8.450 1.350 -8.140 1.480 ;
  END
END sky130_hilas_WTA4Stage01

MACRO sky130_hilas_Trans4small
  CLASS BLOCK ;
  FOREIGN sky130_hilas_Trans4small ;
  ORIGIN -1.910 1.500 ;
  SIZE 2.800 BY 6.050 ;
  PIN NFET_SOURCE1
    USE ANALOG ;
    ANTENNADIFFAREA 0.130200 ;
    PORT
      LAYER met2 ;
        RECT 2.500 4.250 2.810 4.340 ;
        RECT 1.910 4.080 2.810 4.250 ;
        RECT 1.910 3.980 2.050 4.080 ;
        RECT 2.500 4.010 2.810 4.080 ;
    END
  END NFET_SOURCE1
  PIN NFET_GATE1
    USE ANALOG ;
    ANTENNAGATEAREA 0.113400 ;
    PORT
      LAYER met2 ;
        RECT 2.070 3.740 2.380 3.840 ;
        RECT 1.910 3.570 2.380 3.740 ;
        RECT 2.070 3.510 2.380 3.570 ;
    END
  END NFET_GATE1
  PIN NFET_SOURCE2
    USE ANALOG ;
    ANTENNADIFFAREA 0.130200 ;
    PORT
      LAYER met2 ;
        RECT 2.510 3.260 2.820 3.350 ;
        RECT 1.980 3.230 2.820 3.260 ;
        RECT 1.910 3.090 2.820 3.230 ;
        RECT 1.910 3.060 2.050 3.090 ;
        RECT 2.510 3.020 2.820 3.090 ;
    END
  END NFET_SOURCE2
  PIN NFET_GATE2
    USE ANALOG ;
    ANTENNAGATEAREA 0.113400 ;
    PORT
      LAYER met2 ;
        RECT 2.050 2.820 2.360 2.920 ;
        RECT 1.910 2.650 2.360 2.820 ;
        RECT 2.050 2.590 2.360 2.650 ;
    END
  END NFET_GATE2
  PIN NFET_SOURCE3
    USE ANALOG ;
    ANTENNADIFFAREA 0.130200 ;
    PORT
      LAYER met2 ;
        RECT 1.910 2.280 2.050 2.310 ;
        RECT 1.910 2.270 2.120 2.280 ;
        RECT 2.510 2.270 2.820 2.360 ;
        RECT 1.910 2.140 2.820 2.270 ;
        RECT 1.980 2.100 2.820 2.140 ;
        RECT 2.510 2.030 2.820 2.100 ;
    END
  END NFET_SOURCE3
  PIN NFET_GATE3
    USE ANALOG ;
    ANTENNAGATEAREA 0.113400 ;
    PORT
      LAYER met2 ;
        RECT 2.030 1.900 2.340 1.930 ;
        RECT 1.910 1.730 2.340 1.900 ;
        RECT 2.030 1.600 2.340 1.730 ;
    END
  END NFET_GATE3
  PIN PFET_SOURCE1
    USE ANALOG ;
    ANTENNADIFFAREA 0.117600 ;
    PORT
      LAYER met2 ;
        RECT 2.320 1.320 2.630 1.430 ;
        RECT 1.980 1.310 2.630 1.320 ;
        RECT 1.910 1.130 2.630 1.310 ;
        RECT 1.910 1.120 2.050 1.130 ;
        RECT 2.320 1.100 2.630 1.130 ;
    END
  END PFET_SOURCE1
  PIN PFET_GATE1
    USE ANALOG ;
    ANTENNAGATEAREA 0.163800 ;
    PORT
      LAYER met2 ;
        RECT 2.290 0.900 2.610 0.960 ;
        RECT 1.980 0.890 2.610 0.900 ;
        RECT 1.910 0.710 2.610 0.890 ;
        RECT 1.910 0.700 2.050 0.710 ;
        RECT 2.290 0.640 2.610 0.710 ;
    END
  END PFET_GATE1
  PIN PFET_SOURCE2
    USE ANALOG ;
    ANTENNADIFFAREA 0.117600 ;
    PORT
      LAYER met2 ;
        RECT 1.910 0.330 2.050 0.350 ;
        RECT 2.320 0.330 2.630 0.440 ;
        RECT 1.910 0.160 2.630 0.330 ;
        RECT 1.980 0.140 2.630 0.160 ;
        RECT 2.320 0.110 2.630 0.140 ;
    END
  END PFET_SOURCE2
  PIN PFET_GATE2
    USE ANALOG ;
    ANTENNAGATEAREA 0.163800 ;
    PORT
      LAYER met2 ;
        RECT 1.910 -0.090 2.050 -0.070 ;
        RECT 2.290 -0.090 2.610 -0.030 ;
        RECT 1.910 -0.260 2.610 -0.090 ;
        RECT 1.980 -0.280 2.610 -0.260 ;
        RECT 2.290 -0.350 2.610 -0.280 ;
    END
  END PFET_GATE2
  PIN PFET_SOURCE3
    USE ANALOG ;
    ANTENNADIFFAREA 0.117600 ;
    PORT
      LAYER met2 ;
        RECT 1.910 -0.660 2.050 -0.610 ;
        RECT 2.320 -0.660 2.630 -0.550 ;
        RECT 1.910 -0.800 2.630 -0.660 ;
        RECT 1.980 -0.850 2.630 -0.800 ;
        RECT 2.320 -0.880 2.630 -0.850 ;
    END
  END PFET_SOURCE3
  PIN PFET_GATE3
    USE ANALOG ;
    ANTENNAGATEAREA 0.163800 ;
    PORT
      LAYER met2 ;
        RECT 1.910 -1.050 2.050 -1.030 ;
        RECT 1.910 -1.080 2.060 -1.050 ;
        RECT 2.290 -1.080 2.610 -1.020 ;
        RECT 1.910 -1.220 2.610 -1.080 ;
        RECT 1.980 -1.270 2.610 -1.220 ;
        RECT 2.290 -1.340 2.610 -1.270 ;
    END
  END PFET_GATE3
  PIN WELL
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 1.980 1.590 4.010 1.600 ;
        RECT 1.980 -1.500 4.550 1.590 ;
      LAYER met1 ;
        RECT 4.090 -0.200 4.310 4.380 ;
        RECT 4.040 -0.430 4.330 -0.200 ;
        RECT 4.090 -1.500 4.310 -0.430 ;
    END
  END WELL
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 4.490 3.750 4.710 4.380 ;
        RECT 4.480 3.460 4.710 3.750 ;
        RECT 4.490 -1.500 4.710 3.460 ;
    END
  END VGND
  PIN PFET_DRAIN3
    USE ANALOG ;
    ANTENNADIFFAREA 0.113400 ;
    PORT
      LAYER met2 ;
        RECT 3.620 -0.670 3.930 -0.650 ;
        RECT 3.620 -0.870 4.710 -0.670 ;
        RECT 3.620 -0.980 3.930 -0.870 ;
    END
  END PFET_DRAIN3
  PIN PFET_DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.113400 ;
    PORT
      LAYER met2 ;
        RECT 3.620 0.290 3.930 0.340 ;
        RECT 3.620 0.090 4.710 0.290 ;
        RECT 3.620 0.010 3.930 0.090 ;
    END
  END PFET_DRAIN2
  PIN PFET_DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.113400 ;
    PORT
      LAYER met2 ;
        RECT 3.620 1.250 3.930 1.330 ;
        RECT 3.620 1.050 4.710 1.250 ;
        RECT 3.620 1.000 3.930 1.050 ;
    END
  END PFET_DRAIN1
  PIN NFET_DRAIN3
    USE ANALOG ;
    ANTENNADIFFAREA 0.130200 ;
    PORT
      LAYER met2 ;
        RECT 3.600 2.320 3.910 2.370 ;
        RECT 3.600 2.150 4.710 2.320 ;
        RECT 3.600 2.110 4.060 2.150 ;
        RECT 3.600 2.040 3.910 2.110 ;
    END
  END NFET_DRAIN3
  PIN NFET_DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.130200 ;
    PORT
      LAYER met2 ;
        RECT 3.600 3.270 3.910 3.360 ;
        RECT 3.600 3.240 4.060 3.270 ;
        RECT 3.600 3.070 4.710 3.240 ;
        RECT 3.600 3.030 3.910 3.070 ;
    END
  END NFET_DRAIN2
  PIN NFET_DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.130200 ;
    PORT
      LAYER met2 ;
        RECT 3.590 4.260 3.900 4.350 ;
        RECT 3.590 4.160 4.050 4.260 ;
        RECT 3.590 4.020 4.710 4.160 ;
        RECT 3.890 3.990 4.710 4.020 ;
    END
  END NFET_DRAIN1
  OBS
      LAYER li1 ;
        RECT 2.820 4.300 3.020 4.340 ;
        RECT 2.510 4.040 3.020 4.300 ;
        RECT 2.820 4.010 3.020 4.040 ;
        RECT 3.410 4.310 3.610 4.340 ;
        RECT 3.410 4.270 3.920 4.310 ;
        RECT 3.410 4.080 3.930 4.270 ;
        RECT 3.410 4.050 3.920 4.080 ;
        RECT 3.410 4.010 3.610 4.050 ;
        RECT 2.240 3.800 2.600 3.870 ;
        RECT 2.080 3.700 2.600 3.800 ;
        RECT 4.110 3.760 4.280 3.810 ;
        RECT 4.100 3.730 4.280 3.760 ;
        RECT 4.100 3.720 4.530 3.730 ;
        RECT 2.080 3.620 2.450 3.700 ;
        RECT 2.080 3.570 2.410 3.620 ;
        RECT 2.080 3.540 2.400 3.570 ;
        RECT 4.100 3.490 4.690 3.720 ;
        RECT 4.100 3.480 4.530 3.490 ;
        RECT 4.100 3.450 4.290 3.480 ;
        RECT 4.110 3.420 4.290 3.450 ;
        RECT 2.830 3.310 3.030 3.350 ;
        RECT 2.520 3.050 3.030 3.310 ;
        RECT 2.830 3.020 3.030 3.050 ;
        RECT 3.420 3.320 3.620 3.350 ;
        RECT 3.420 3.280 3.930 3.320 ;
        RECT 3.420 3.090 3.940 3.280 ;
        RECT 3.420 3.060 3.930 3.090 ;
        RECT 3.420 3.020 3.620 3.060 ;
        RECT 2.060 2.710 2.610 2.880 ;
        RECT 2.060 2.650 2.390 2.710 ;
        RECT 2.060 2.620 2.380 2.650 ;
        RECT 2.830 2.320 3.030 2.360 ;
        RECT 2.520 2.060 3.030 2.320 ;
        RECT 2.830 2.030 3.030 2.060 ;
        RECT 3.420 2.330 3.620 2.360 ;
        RECT 3.420 2.290 3.930 2.330 ;
        RECT 3.420 2.100 3.940 2.290 ;
        RECT 3.420 2.070 3.930 2.100 ;
        RECT 3.420 2.030 3.620 2.070 ;
        RECT 2.040 1.720 2.610 1.890 ;
        RECT 2.040 1.660 2.370 1.720 ;
        RECT 2.040 1.630 2.360 1.660 ;
        RECT 2.330 1.350 2.650 1.390 ;
        RECT 2.330 1.330 2.660 1.350 ;
        RECT 2.330 1.130 2.950 1.330 ;
        RECT 2.780 1.000 2.950 1.130 ;
        RECT 3.460 1.290 3.630 1.330 ;
        RECT 3.460 1.250 3.950 1.290 ;
        RECT 3.460 1.060 3.960 1.250 ;
        RECT 3.460 1.030 3.950 1.060 ;
        RECT 3.460 1.000 3.630 1.030 ;
        RECT 2.140 0.890 2.570 0.910 ;
        RECT 2.120 0.720 2.570 0.890 ;
        RECT 2.140 0.700 2.570 0.720 ;
        RECT 2.330 0.360 2.650 0.400 ;
        RECT 2.330 0.340 2.660 0.360 ;
        RECT 2.330 0.140 2.950 0.340 ;
        RECT 2.780 0.010 2.950 0.140 ;
        RECT 3.460 0.300 3.630 0.340 ;
        RECT 3.460 0.260 3.950 0.300 ;
        RECT 3.460 0.070 3.960 0.260 ;
        RECT 3.460 0.040 3.950 0.070 ;
        RECT 3.460 0.010 3.630 0.040 ;
        RECT 2.140 -0.100 2.570 -0.080 ;
        RECT 2.120 -0.270 2.570 -0.100 ;
        RECT 4.070 -0.230 4.300 -0.220 ;
        RECT 2.140 -0.290 2.570 -0.270 ;
        RECT 3.990 -0.400 4.320 -0.230 ;
        RECT 4.070 -0.410 4.300 -0.400 ;
        RECT 2.330 -0.630 2.650 -0.590 ;
        RECT 2.330 -0.650 2.660 -0.630 ;
        RECT 2.330 -0.850 2.950 -0.650 ;
        RECT 2.780 -0.980 2.950 -0.850 ;
        RECT 3.460 -0.690 3.630 -0.650 ;
        RECT 3.460 -0.730 3.950 -0.690 ;
        RECT 3.460 -0.920 3.960 -0.730 ;
        RECT 3.460 -0.950 3.950 -0.920 ;
        RECT 3.460 -0.980 3.630 -0.950 ;
        RECT 2.140 -1.090 2.570 -1.070 ;
        RECT 2.120 -1.260 2.570 -1.090 ;
        RECT 2.140 -1.280 2.570 -1.260 ;
      LAYER mcon ;
        RECT 2.570 4.080 2.740 4.250 ;
        RECT 3.660 4.090 3.830 4.260 ;
        RECT 2.140 3.580 2.310 3.750 ;
        RECT 4.510 3.520 4.680 3.690 ;
        RECT 2.580 3.090 2.750 3.260 ;
        RECT 3.670 3.100 3.840 3.270 ;
        RECT 2.120 2.660 2.290 2.830 ;
        RECT 2.580 2.100 2.750 2.270 ;
        RECT 3.670 2.110 3.840 2.280 ;
        RECT 2.100 1.670 2.270 1.840 ;
        RECT 2.390 1.170 2.560 1.340 ;
        RECT 3.690 1.070 3.860 1.240 ;
        RECT 2.390 0.180 2.560 0.350 ;
        RECT 3.690 0.080 3.860 0.250 ;
        RECT 4.100 -0.400 4.270 -0.230 ;
        RECT 2.390 -0.810 2.560 -0.640 ;
        RECT 3.690 -0.910 3.860 -0.740 ;
      LAYER met1 ;
        RECT 2.500 4.010 2.820 4.330 ;
        RECT 3.590 4.020 3.910 4.340 ;
        RECT 2.070 3.510 2.390 3.830 ;
        RECT 2.510 3.020 2.830 3.340 ;
        RECT 3.600 3.030 3.920 3.350 ;
        RECT 2.050 2.590 2.370 2.910 ;
        RECT 2.510 2.030 2.830 2.350 ;
        RECT 3.600 2.040 3.920 2.360 ;
        RECT 2.030 1.600 2.350 1.920 ;
        RECT 2.320 1.100 2.640 1.420 ;
        RECT 3.620 1.000 3.940 1.320 ;
        RECT 2.290 0.920 2.610 0.960 ;
        RECT 2.060 0.690 2.610 0.920 ;
        RECT 2.290 0.640 2.610 0.690 ;
        RECT 2.320 0.110 2.640 0.430 ;
        RECT 3.620 0.010 3.940 0.330 ;
        RECT 2.290 -0.070 2.610 -0.030 ;
        RECT 2.060 -0.300 2.610 -0.070 ;
        RECT 2.290 -0.350 2.610 -0.300 ;
        RECT 2.320 -0.880 2.640 -0.560 ;
        RECT 3.620 -0.980 3.940 -0.660 ;
        RECT 2.290 -1.060 2.610 -1.020 ;
        RECT 2.060 -1.290 2.610 -1.060 ;
        RECT 2.290 -1.340 2.610 -1.290 ;
      LAYER via ;
        RECT 2.530 4.040 2.790 4.300 ;
        RECT 3.620 4.050 3.880 4.310 ;
        RECT 2.100 3.540 2.360 3.800 ;
        RECT 2.540 3.050 2.800 3.310 ;
        RECT 3.630 3.060 3.890 3.320 ;
        RECT 2.080 2.620 2.340 2.880 ;
        RECT 2.540 2.060 2.800 2.320 ;
        RECT 3.630 2.070 3.890 2.330 ;
        RECT 2.060 1.630 2.320 1.890 ;
        RECT 2.350 1.130 2.610 1.390 ;
        RECT 3.650 1.030 3.910 1.290 ;
        RECT 2.320 0.670 2.580 0.930 ;
        RECT 2.350 0.140 2.610 0.400 ;
        RECT 3.650 0.040 3.910 0.300 ;
        RECT 2.320 -0.320 2.580 -0.060 ;
        RECT 2.350 -0.850 2.610 -0.590 ;
        RECT 3.650 -0.950 3.910 -0.690 ;
        RECT 2.320 -1.310 2.580 -1.050 ;
  END
END sky130_hilas_Trans4small

MACRO sky130_hilas_FGBiasWeakGate2x1cell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_FGBiasWeakGate2x1cell ;
  ORIGIN 3.960 3.870 ;
  SIZE 11.530 BY 6.150 ;
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 5.090 1.730 5.400 1.740 ;
        RECT -3.960 1.550 7.570 1.730 ;
        RECT 5.090 1.410 5.400 1.550 ;
    END
  END DRAIN1
  PIN VIN11
    PORT
      LAYER met2 ;
        RECT -2.020 1.140 -1.710 1.190 ;
        RECT -2.170 1.130 -1.710 1.140 ;
        RECT -3.960 0.950 -1.710 1.130 ;
        RECT -2.020 0.860 -1.710 0.950 ;
    END
  END VIN11
  PIN ROW1
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 5.240 0.710 5.550 0.780 ;
        RECT 5.240 0.700 7.570 0.710 ;
        RECT -3.960 0.490 7.570 0.700 ;
        RECT -3.960 0.480 6.260 0.490 ;
        RECT 5.240 0.450 5.550 0.480 ;
    END
  END ROW1
  PIN ROW2
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 5.240 -2.050 5.550 -1.980 ;
        RECT -3.960 -2.260 7.570 -2.050 ;
        RECT -3.960 -2.270 6.260 -2.260 ;
        RECT 5.240 -2.310 5.550 -2.270 ;
    END
  END ROW2
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 4.260 -3.870 7.570 2.280 ;
      LAYER met1 ;
        RECT 7.050 1.580 7.330 2.230 ;
        RECT 6.940 0.980 7.330 1.580 ;
        RECT 7.050 -2.570 7.330 0.980 ;
        RECT 6.940 -3.170 7.330 -2.570 ;
        RECT 7.050 -3.820 7.330 -3.170 ;
    END
  END VINJ
  PIN COLSEL1
    USE ANALOG ;
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT 6.610 0.770 6.800 2.230 ;
        RECT 6.610 0.740 6.830 0.770 ;
        RECT 6.590 0.470 6.840 0.740 ;
        RECT 6.600 0.460 6.840 0.470 ;
        RECT 6.600 0.220 6.830 0.460 ;
        RECT 6.640 -1.810 6.800 0.220 ;
        RECT 6.600 -2.050 6.830 -1.810 ;
        RECT 6.600 -2.060 6.840 -2.050 ;
        RECT 6.590 -2.330 6.840 -2.060 ;
        RECT 6.610 -2.360 6.830 -2.330 ;
        RECT 6.610 -3.820 6.800 -2.360 ;
    END
  END COLSEL1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT -1.130 1.260 -0.900 2.230 ;
        RECT -1.130 1.010 -0.890 1.260 ;
        RECT -1.130 -3.820 -0.900 1.010 ;
    END
  END VGND
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT -0.190 -0.160 2.530 1.490 ;
        RECT -0.190 -0.200 2.520 -0.160 ;
        RECT -0.190 -1.530 2.520 -1.490 ;
        RECT -0.190 -3.180 2.530 -1.530 ;
      LAYER met1 ;
        RECT 0.090 1.020 0.320 2.230 ;
        RECT 0.090 0.230 0.350 1.020 ;
        RECT 0.090 -1.920 0.320 0.230 ;
        RECT 0.090 -2.710 0.350 -1.920 ;
        RECT 0.090 -3.820 0.320 -2.710 ;
    END
  END GATE1
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 2.516100 ;
    PORT
      LAYER nwell ;
        RECT -3.950 1.480 -2.220 2.230 ;
        RECT -3.950 0.330 -2.210 1.480 ;
        RECT -3.940 -1.910 -2.210 0.330 ;
        RECT -3.950 -2.090 -2.210 -1.910 ;
        RECT -3.950 -3.810 -2.220 -2.090 ;
      LAYER met1 ;
        RECT -3.610 -3.810 -3.190 2.230 ;
    END
  END VTUN
  PIN DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 5.090 -3.140 5.400 -3.000 ;
        RECT 5.090 -3.150 7.570 -3.140 ;
        RECT -3.960 -3.300 7.570 -3.150 ;
        RECT 5.090 -3.320 7.570 -3.300 ;
        RECT 5.090 -3.330 5.400 -3.320 ;
    END
  END DRAIN2
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -2.050 -2.580 -1.740 -2.500 ;
        RECT -3.960 -2.790 -1.740 -2.580 ;
        RECT -2.050 -2.830 -1.740 -2.790 ;
    END
  END VIN12
  PIN COMMONSOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 1.030400 ;
    PORT
      LAYER met2 ;
        RECT -3.960 -0.490 6.500 -0.270 ;
        RECT 6.180 -0.630 6.500 -0.490 ;
        RECT 6.220 -0.970 6.480 -0.630 ;
        RECT 6.180 -1.230 6.500 -0.970 ;
    END
  END COMMONSOURCE
  OBS
      LAYER li1 ;
        RECT -2.090 1.220 2.970 2.050 ;
        RECT 5.160 1.650 5.690 1.820 ;
        RECT 6.970 1.550 7.170 1.900 ;
        RECT 6.970 1.520 7.180 1.550 ;
        RECT -2.020 1.140 -1.540 1.220 ;
        RECT -2.010 0.890 -1.540 1.140 ;
        RECT -3.520 0.090 -2.970 0.520 ;
        RECT 0.110 0.280 0.340 0.970 ;
        RECT 5.410 0.740 5.580 1.260 ;
        RECT 5.250 0.480 5.580 0.740 ;
        RECT -0.920 -0.740 -0.730 -0.340 ;
        RECT 5.410 -0.430 5.580 0.480 ;
        RECT 6.240 -0.340 6.410 1.270 ;
        RECT 6.960 0.940 7.180 1.520 ;
        RECT 6.970 0.930 7.180 0.940 ;
        RECT 6.610 0.760 6.800 0.770 ;
        RECT 6.610 0.470 6.810 0.760 ;
        RECT 6.600 0.140 6.890 0.470 ;
        RECT 6.240 -0.530 6.420 -0.340 ;
        RECT -1.110 -0.750 -0.730 -0.740 ;
        RECT -1.110 -0.930 2.630 -0.750 ;
        RECT -1.110 -0.970 -0.730 -0.930 ;
        RECT -3.520 -1.640 -2.970 -1.210 ;
        RECT -0.920 -1.350 -0.730 -0.970 ;
        RECT -2.040 -2.790 -1.700 -2.540 ;
        RECT 0.110 -2.660 0.340 -1.930 ;
        RECT 5.410 -2.020 5.580 -1.160 ;
        RECT 5.250 -2.280 5.580 -2.020 ;
        RECT -2.050 -2.870 -1.700 -2.790 ;
        RECT 5.410 -2.850 5.580 -2.280 ;
        RECT 6.240 -1.250 6.420 -1.060 ;
        RECT 6.240 -2.860 6.410 -1.250 ;
        RECT 6.600 -2.060 6.890 -1.730 ;
        RECT 6.610 -2.350 6.810 -2.060 ;
        RECT 6.610 -2.360 6.800 -2.350 ;
        RECT 6.970 -2.530 7.180 -2.520 ;
        RECT -2.050 -3.720 3.000 -2.870 ;
        RECT 6.960 -3.110 7.180 -2.530 ;
        RECT 6.970 -3.140 7.180 -3.110 ;
        RECT 5.160 -3.410 5.690 -3.240 ;
        RECT 6.970 -3.490 7.170 -3.140 ;
      LAYER mcon ;
        RECT 6.980 1.350 7.150 1.520 ;
        RECT -1.950 0.930 -1.780 1.100 ;
        RECT 0.140 0.770 0.310 0.940 ;
        RECT -3.520 0.170 -3.250 0.440 ;
        RECT 0.140 0.320 0.310 0.490 ;
        RECT 5.310 0.520 5.480 0.690 ;
        RECT 6.620 0.510 6.800 0.700 ;
        RECT -1.100 -0.940 -0.930 -0.770 ;
        RECT -3.520 -1.560 -3.250 -1.290 ;
        RECT 0.140 -2.180 0.310 -2.010 ;
        RECT 5.310 -2.240 5.480 -2.070 ;
        RECT -1.980 -2.760 -1.810 -2.590 ;
        RECT 0.140 -2.630 0.310 -2.460 ;
        RECT 6.620 -2.290 6.800 -2.100 ;
        RECT 6.980 -3.110 7.150 -2.940 ;
      LAYER met1 ;
        RECT 5.090 1.410 5.400 1.850 ;
        RECT -2.020 0.860 -1.700 1.180 ;
        RECT 5.240 0.450 5.560 0.770 ;
        RECT 6.210 -0.340 6.450 -0.210 ;
        RECT 6.210 -0.660 6.470 -0.340 ;
        RECT 6.210 -1.260 6.470 -0.940 ;
        RECT 6.210 -1.380 6.450 -1.260 ;
        RECT 5.240 -2.310 5.560 -1.990 ;
        RECT -2.050 -2.830 -1.730 -2.510 ;
        RECT 5.090 -3.440 5.400 -3.000 ;
      LAYER via ;
        RECT 5.120 1.440 5.380 1.700 ;
        RECT -1.990 0.890 -1.730 1.150 ;
        RECT 5.270 0.480 5.530 0.740 ;
        RECT 6.210 -0.630 6.470 -0.370 ;
        RECT 6.210 -1.230 6.470 -0.970 ;
        RECT 5.270 -2.280 5.530 -2.020 ;
        RECT -2.020 -2.800 -1.760 -2.540 ;
        RECT 5.120 -3.290 5.380 -3.030 ;
  END
END sky130_hilas_FGBiasWeakGate2x1cell

MACRO sky130_hilas_swc4x2cell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc4x2cell ;
  ORIGIN 10.040 0.260 ;
  SIZE 20.120 BY 6.500 ;
  PIN GATE2
    USE ANALOG ;
    ANTENNADIFFAREA 3.253900 ;
    PORT
      LAYER nwell ;
        RECT 3.760 -0.260 5.990 6.230 ;
      LAYER met1 ;
        RECT 4.410 4.090 4.790 6.240 ;
        RECT 4.400 2.230 4.790 4.090 ;
        RECT 4.410 -0.260 4.790 2.230 ;
    END
  END GATE2
  PIN VTUN
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -1.700 -0.260 1.740 6.230 ;
      LAYER met1 ;
        RECT -0.720 5.870 -0.320 6.240 ;
        RECT 0.360 5.870 0.760 6.240 ;
        RECT -0.720 5.650 0.760 5.870 ;
        RECT -0.720 -0.260 -0.320 5.650 ;
        RECT 0.360 -0.260 0.760 5.650 ;
    END
  END VTUN
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 3.253900 ;
    PORT
      LAYER nwell ;
        RECT -5.950 -0.260 -3.720 6.230 ;
      LAYER met1 ;
        RECT -4.750 4.090 -4.370 6.240 ;
        RECT -4.750 2.230 -4.360 4.090 ;
        RECT -4.750 -0.260 -4.370 2.230 ;
    END
  END GATE1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -10.040 -0.260 -7.480 6.240 ;
        RECT 7.520 -0.260 10.080 6.240 ;
      LAYER met2 ;
        RECT -9.840 5.960 9.900 6.140 ;
        RECT -9.840 5.820 -9.420 5.960 ;
        RECT 9.560 5.830 9.900 5.960 ;
    END
  END VINJ
  PIN VINJ
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 9.560 6.120 9.720 6.230 ;
        RECT 9.560 5.840 9.890 6.120 ;
        RECT 9.560 5.530 9.720 5.840 ;
        RECT 9.450 4.980 9.720 5.530 ;
        RECT 9.450 4.930 9.730 4.980 ;
        RECT 9.560 4.840 9.730 4.930 ;
        RECT 9.560 4.370 9.720 4.840 ;
        RECT 9.560 4.280 9.730 4.370 ;
        RECT 9.450 4.230 9.730 4.280 ;
        RECT 9.450 3.680 9.720 4.230 ;
        RECT 9.560 2.290 9.720 3.680 ;
        RECT 9.450 1.740 9.720 2.290 ;
        RECT 9.450 1.690 9.730 1.740 ;
        RECT 9.560 1.600 9.730 1.690 ;
        RECT 9.560 1.140 9.720 1.600 ;
        RECT 9.560 1.050 9.730 1.140 ;
        RECT 9.450 1.000 9.730 1.050 ;
        RECT 9.450 0.450 9.720 1.000 ;
        RECT 9.560 -0.250 9.720 0.450 ;
      LAYER via ;
        RECT 9.600 5.850 9.860 6.110 ;
    END
    PORT
      LAYER met1 ;
        RECT -9.680 6.110 -9.520 6.230 ;
        RECT -9.830 5.970 -9.520 6.110 ;
        RECT -9.840 5.820 -9.520 5.970 ;
        RECT -9.680 5.530 -9.520 5.820 ;
        RECT -9.680 4.980 -9.410 5.530 ;
        RECT -9.690 4.930 -9.410 4.980 ;
        RECT -9.690 4.840 -9.520 4.930 ;
        RECT -9.680 4.370 -9.520 4.840 ;
        RECT -9.690 4.280 -9.520 4.370 ;
        RECT -9.690 4.230 -9.410 4.280 ;
        RECT -9.680 3.680 -9.410 4.230 ;
        RECT -9.680 2.290 -9.520 3.680 ;
        RECT -9.680 1.740 -9.410 2.290 ;
        RECT -9.690 1.690 -9.410 1.740 ;
        RECT -9.690 1.600 -9.520 1.690 ;
        RECT -9.680 1.140 -9.520 1.600 ;
        RECT -9.690 1.050 -9.520 1.140 ;
        RECT -9.690 1.000 -9.410 1.050 ;
        RECT -9.680 0.450 -9.410 1.000 ;
        RECT -9.680 -0.250 -9.520 0.450 ;
      LAYER via ;
        RECT -9.800 5.840 -9.540 6.100 ;
    END
  END VINJ
  PIN GATESELECT1
    USE ANALOG ;
    ANTENNAGATEAREA 0.720000 ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met1 ;
        RECT -9.270 5.190 -9.080 6.180 ;
        RECT -8.870 5.500 -8.710 6.230 ;
        RECT -8.910 5.480 -8.710 5.500 ;
        RECT -8.920 5.240 -8.690 5.480 ;
        RECT -8.920 5.190 -8.710 5.240 ;
        RECT -9.270 5.070 -9.100 5.190 ;
        RECT -9.270 4.140 -9.110 5.070 ;
        RECT -9.270 4.020 -9.100 4.140 ;
        RECT -8.870 4.020 -8.710 5.190 ;
        RECT -9.270 3.100 -9.080 4.020 ;
        RECT -8.920 3.970 -8.710 4.020 ;
        RECT -8.920 3.730 -8.690 3.970 ;
        RECT -8.910 3.710 -8.710 3.730 ;
        RECT -9.300 3.080 -9.060 3.100 ;
        RECT -8.870 3.080 -8.710 3.710 ;
        RECT -9.300 2.890 -8.710 3.080 ;
        RECT -9.300 2.870 -9.060 2.890 ;
        RECT -9.270 1.950 -9.080 2.870 ;
        RECT -8.870 2.260 -8.710 2.890 ;
        RECT -8.910 2.240 -8.710 2.260 ;
        RECT -8.920 2.000 -8.690 2.240 ;
        RECT -8.920 1.950 -8.710 2.000 ;
        RECT -9.270 1.830 -9.100 1.950 ;
        RECT -9.270 0.910 -9.110 1.830 ;
        RECT -9.270 0.790 -9.100 0.910 ;
        RECT -8.870 0.790 -8.710 1.950 ;
        RECT -9.270 -0.200 -9.080 0.790 ;
        RECT -8.920 0.740 -8.710 0.790 ;
        RECT -8.920 0.500 -8.690 0.740 ;
        RECT -8.910 0.480 -8.710 0.500 ;
        RECT -8.870 -0.250 -8.710 0.480 ;
    END
  END GATESELECT1
  PIN GATESELECT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.720000 ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met1 ;
        RECT 8.750 5.500 8.910 6.230 ;
        RECT 8.750 5.480 8.950 5.500 ;
        RECT 8.730 5.240 8.960 5.480 ;
        RECT 8.750 5.190 8.960 5.240 ;
        RECT 9.120 5.190 9.310 6.180 ;
        RECT 8.750 4.020 8.910 5.190 ;
        RECT 9.140 5.070 9.310 5.190 ;
        RECT 9.150 4.140 9.310 5.070 ;
        RECT 9.140 4.020 9.310 4.140 ;
        RECT 8.750 3.970 8.960 4.020 ;
        RECT 8.730 3.730 8.960 3.970 ;
        RECT 8.750 3.710 8.950 3.730 ;
        RECT 8.750 3.080 8.910 3.710 ;
        RECT 9.120 3.100 9.310 4.020 ;
        RECT 9.100 3.080 9.340 3.100 ;
        RECT 8.750 2.890 9.340 3.080 ;
        RECT 8.750 2.260 8.910 2.890 ;
        RECT 9.100 2.870 9.340 2.890 ;
        RECT 8.750 2.240 8.950 2.260 ;
        RECT 8.730 2.000 8.960 2.240 ;
        RECT 8.750 1.950 8.960 2.000 ;
        RECT 9.120 1.950 9.310 2.870 ;
        RECT 8.750 0.790 8.910 1.950 ;
        RECT 9.140 1.830 9.310 1.950 ;
        RECT 9.150 0.910 9.310 1.830 ;
        RECT 9.140 0.790 9.310 0.910 ;
        RECT 8.750 0.740 8.960 0.790 ;
        RECT 8.730 0.500 8.960 0.740 ;
        RECT 8.750 0.480 8.950 0.500 ;
        RECT 8.750 -0.250 8.910 0.480 ;
        RECT 9.120 -0.200 9.310 0.790 ;
    END
  END GATESELECT2
  PIN ROW1
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT -7.880 5.250 -7.570 5.270 ;
        RECT 7.610 5.250 7.920 5.270 ;
        RECT -10.040 5.240 -7.480 5.250 ;
        RECT 7.520 5.240 10.080 5.250 ;
        RECT -10.040 5.070 10.080 5.240 ;
        RECT -7.880 5.060 7.920 5.070 ;
        RECT -7.880 4.940 -7.570 5.060 ;
        RECT 7.610 4.940 7.920 5.060 ;
    END
  END ROW1
  PIN ROW2
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT -7.880 4.140 -7.570 4.270 ;
        RECT 7.610 4.140 7.920 4.270 ;
        RECT -10.040 3.960 10.080 4.140 ;
        RECT -7.880 3.940 -7.570 3.960 ;
        RECT 7.610 3.940 7.920 3.960 ;
    END
  END ROW2
  PIN DRAIN1
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT -7.880 5.680 -7.570 5.820 ;
        RECT 7.610 5.680 7.920 5.820 ;
        RECT -10.040 5.500 10.080 5.680 ;
        RECT -7.880 5.490 -7.570 5.500 ;
        RECT 7.610 5.490 7.920 5.500 ;
    END
  END DRAIN1
  PIN DRAIN2
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT -7.880 3.710 -7.570 3.720 ;
        RECT 7.610 3.710 7.920 3.720 ;
        RECT -10.040 3.530 10.080 3.710 ;
        RECT -7.880 3.390 -7.570 3.530 ;
        RECT 7.610 3.390 7.920 3.530 ;
    END
  END DRAIN2
  PIN DRAIN3
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT -7.880 2.440 -7.570 2.580 ;
        RECT 7.610 2.440 7.920 2.580 ;
        RECT -10.040 2.260 10.080 2.440 ;
        RECT -7.880 2.250 -7.570 2.260 ;
        RECT 7.610 2.250 7.920 2.260 ;
    END
  END DRAIN3
  PIN ROW3
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT -7.880 2.010 -7.570 2.030 ;
        RECT 7.610 2.010 7.920 2.030 ;
        RECT -10.040 1.830 10.080 2.010 ;
        RECT -7.880 1.700 -7.570 1.830 ;
        RECT 7.610 1.700 7.920 1.830 ;
    END
  END ROW3
  PIN ROW4
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT -7.880 0.910 -7.570 1.040 ;
        RECT 7.610 0.910 7.920 1.040 ;
        RECT -10.040 0.730 10.080 0.910 ;
        RECT -7.880 0.710 -7.570 0.730 ;
        RECT 7.610 0.710 7.920 0.730 ;
    END
  END ROW4
  PIN DRAIN4
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT -7.880 0.480 -7.570 0.490 ;
        RECT 7.610 0.480 7.920 0.490 ;
        RECT -10.040 0.310 10.080 0.480 ;
        RECT -10.040 0.300 -7.570 0.310 ;
        RECT -7.880 0.160 -7.570 0.300 ;
        RECT 7.610 0.300 10.080 0.310 ;
        RECT 7.610 0.160 7.920 0.300 ;
    END
  END DRAIN4
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT -6.970 1.520 -6.650 1.580 ;
        RECT -3.040 1.520 -2.720 1.530 ;
        RECT 2.760 1.520 3.080 1.530 ;
        RECT 6.690 1.520 7.010 1.580 ;
        RECT -6.970 1.340 7.010 1.520 ;
        RECT -6.970 1.290 -6.650 1.340 ;
        RECT -3.040 1.270 -2.720 1.340 ;
        RECT 2.760 1.270 3.080 1.340 ;
        RECT 6.690 1.290 7.010 1.340 ;
    END
    PORT
      LAYER met1 ;
        RECT -6.930 4.850 -6.690 6.240 ;
        RECT -6.940 4.190 -6.670 4.850 ;
        RECT -6.930 1.600 -6.690 4.190 ;
        RECT -6.940 1.280 -6.680 1.600 ;
        RECT -6.930 -0.260 -6.690 1.280 ;
      LAYER via ;
        RECT -6.940 1.310 -6.680 1.570 ;
    END
    PORT
      LAYER met1 ;
        RECT -3.000 4.830 -2.760 6.240 ;
        RECT -3.010 4.170 -2.750 4.830 ;
        RECT -3.000 1.560 -2.760 4.170 ;
        RECT -3.010 1.240 -2.750 1.560 ;
        RECT -3.000 -0.260 -2.760 1.240 ;
      LAYER via ;
        RECT -3.010 1.270 -2.750 1.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.800 4.830 3.040 6.240 ;
        RECT 2.790 4.170 3.050 4.830 ;
        RECT 2.800 1.560 3.040 4.170 ;
        RECT 2.790 1.240 3.050 1.560 ;
        RECT 2.800 -0.260 3.040 1.240 ;
      LAYER via ;
        RECT 2.790 1.270 3.050 1.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.730 4.850 6.970 6.240 ;
        RECT 6.710 4.190 6.980 4.850 ;
        RECT 6.730 1.600 6.970 4.190 ;
        RECT 6.720 1.280 6.980 1.600 ;
        RECT 6.730 -0.260 6.970 1.280 ;
      LAYER via ;
        RECT 6.720 1.310 6.980 1.570 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT -9.640 5.500 -9.440 5.850 ;
        RECT -7.900 5.770 -7.580 5.780 ;
        RECT -8.160 5.600 -7.580 5.770 ;
        RECT -7.910 5.550 -7.580 5.600 ;
        RECT -7.900 5.520 -7.580 5.550 ;
        RECT 7.620 5.770 7.940 5.780 ;
        RECT 7.620 5.600 8.200 5.770 ;
        RECT 7.620 5.550 7.950 5.600 ;
        RECT 7.620 5.520 7.940 5.550 ;
        RECT -9.650 5.470 -9.440 5.500 ;
        RECT 9.480 5.500 9.680 5.850 ;
        RECT -9.650 4.880 -9.430 5.470 ;
        RECT -8.910 4.880 -8.710 5.480 ;
        RECT -7.900 5.190 -7.580 5.230 ;
        RECT -7.910 5.150 -7.580 5.190 ;
        RECT -8.160 4.980 -7.580 5.150 ;
        RECT -7.900 4.970 -7.580 4.980 ;
        RECT 7.620 5.190 7.940 5.230 ;
        RECT 7.620 5.150 7.950 5.190 ;
        RECT 7.620 4.980 8.200 5.150 ;
        RECT 7.620 4.970 7.940 4.980 ;
        RECT 8.750 4.880 8.950 5.480 ;
        RECT 9.480 5.470 9.690 5.500 ;
        RECT 9.470 4.880 9.690 5.470 ;
        RECT -9.650 3.740 -9.430 4.330 ;
        RECT -9.650 3.710 -9.440 3.740 ;
        RECT -8.910 3.730 -8.710 4.330 ;
        RECT -6.900 4.250 -6.730 4.780 ;
        RECT -2.960 4.260 -2.790 4.790 ;
        RECT 2.830 4.260 3.000 4.790 ;
        RECT 6.770 4.250 6.940 4.780 ;
        RECT -7.900 4.230 -7.580 4.240 ;
        RECT -8.160 4.060 -7.580 4.230 ;
        RECT -7.910 4.020 -7.580 4.060 ;
        RECT -7.900 3.980 -7.580 4.020 ;
        RECT 7.620 4.230 7.940 4.240 ;
        RECT 7.620 4.060 8.200 4.230 ;
        RECT 7.620 4.020 7.950 4.060 ;
        RECT 7.620 3.980 7.940 4.020 ;
        RECT 8.750 3.730 8.950 4.330 ;
        RECT 9.470 3.740 9.690 4.330 ;
        RECT -9.640 3.360 -9.440 3.710 ;
        RECT 9.480 3.710 9.690 3.740 ;
        RECT -7.900 3.660 -7.580 3.690 ;
        RECT -7.910 3.610 -7.580 3.660 ;
        RECT -8.160 3.440 -7.580 3.610 ;
        RECT 7.620 3.660 7.940 3.690 ;
        RECT 7.620 3.610 7.950 3.660 ;
        RECT -7.900 3.430 -7.580 3.440 ;
        RECT -9.270 2.900 -8.830 3.070 ;
        RECT -9.640 2.260 -9.440 2.610 ;
        RECT -7.900 2.530 -7.580 2.540 ;
        RECT -8.160 2.360 -7.580 2.530 ;
        RECT -6.900 2.410 -6.730 3.420 ;
        RECT -4.970 2.690 -4.420 3.120 ;
        RECT -2.970 2.550 -2.800 3.560 ;
        RECT -0.940 2.760 -0.390 3.190 ;
        RECT 0.430 2.760 0.980 3.190 ;
        RECT 2.840 2.550 3.010 3.560 ;
        RECT 7.620 3.440 8.200 3.610 ;
        RECT 7.620 3.430 7.940 3.440 ;
        RECT 4.460 2.690 5.010 3.120 ;
        RECT 6.770 2.410 6.940 3.420 ;
        RECT 9.480 3.360 9.680 3.710 ;
        RECT 8.870 2.900 9.310 3.070 ;
        RECT 7.620 2.530 7.940 2.540 ;
        RECT -7.910 2.310 -7.580 2.360 ;
        RECT -7.900 2.280 -7.580 2.310 ;
        RECT 7.620 2.360 8.200 2.530 ;
        RECT 7.620 2.310 7.950 2.360 ;
        RECT 7.620 2.280 7.940 2.310 ;
        RECT -9.650 2.230 -9.440 2.260 ;
        RECT 9.480 2.260 9.680 2.610 ;
        RECT -9.650 1.640 -9.430 2.230 ;
        RECT -8.910 1.640 -8.710 2.240 ;
        RECT -7.900 1.950 -7.580 1.990 ;
        RECT -7.910 1.910 -7.580 1.950 ;
        RECT -8.160 1.740 -7.580 1.910 ;
        RECT -7.900 1.730 -7.580 1.740 ;
        RECT 7.620 1.950 7.940 1.990 ;
        RECT 7.620 1.910 7.950 1.950 ;
        RECT 7.620 1.740 8.200 1.910 ;
        RECT 7.620 1.730 7.940 1.740 ;
        RECT 8.750 1.640 8.950 2.240 ;
        RECT 9.480 2.230 9.690 2.260 ;
        RECT 9.470 1.640 9.690 2.230 ;
        RECT -9.650 0.510 -9.430 1.100 ;
        RECT -9.650 0.480 -9.440 0.510 ;
        RECT -8.910 0.500 -8.710 1.100 ;
        RECT -7.900 1.000 -7.580 1.010 ;
        RECT -8.160 0.830 -7.580 1.000 ;
        RECT -7.910 0.790 -7.580 0.830 ;
        RECT -7.900 0.750 -7.580 0.790 ;
        RECT 7.620 1.000 7.940 1.010 ;
        RECT 7.620 0.830 8.200 1.000 ;
        RECT 7.620 0.790 7.950 0.830 ;
        RECT 7.620 0.750 7.940 0.790 ;
        RECT 8.750 0.500 8.950 1.100 ;
        RECT 9.470 0.510 9.690 1.100 ;
        RECT -9.640 0.130 -9.440 0.480 ;
        RECT 9.480 0.480 9.690 0.510 ;
        RECT -7.900 0.430 -7.580 0.460 ;
        RECT -7.910 0.380 -7.580 0.430 ;
        RECT -8.160 0.210 -7.580 0.380 ;
        RECT -7.900 0.200 -7.580 0.210 ;
        RECT 7.620 0.430 7.940 0.460 ;
        RECT 7.620 0.380 7.950 0.430 ;
        RECT 7.620 0.210 8.200 0.380 ;
        RECT 7.620 0.200 7.940 0.210 ;
        RECT 9.480 0.130 9.680 0.480 ;
      LAYER mcon ;
        RECT -7.810 5.560 -7.640 5.730 ;
        RECT 7.680 5.560 7.850 5.730 ;
        RECT -9.620 5.300 -9.450 5.470 ;
        RECT -8.890 5.270 -8.720 5.440 ;
        RECT 8.760 5.270 8.930 5.440 ;
        RECT -7.810 5.010 -7.640 5.180 ;
        RECT 7.680 5.010 7.850 5.180 ;
        RECT 9.490 5.300 9.660 5.470 ;
        RECT -6.900 4.610 -6.730 4.780 ;
        RECT -9.620 3.740 -9.450 3.910 ;
        RECT -2.960 4.620 -2.790 4.790 ;
        RECT 2.830 4.620 3.000 4.790 ;
        RECT 6.770 4.610 6.940 4.780 ;
        RECT -7.810 4.030 -7.640 4.200 ;
        RECT 7.680 4.030 7.850 4.200 ;
        RECT -8.890 3.770 -8.720 3.940 ;
        RECT 8.760 3.770 8.930 3.940 ;
        RECT 9.490 3.740 9.660 3.910 ;
        RECT -7.810 3.480 -7.640 3.650 ;
        RECT -6.900 3.020 -6.730 3.190 ;
        RECT -2.970 3.160 -2.800 3.330 ;
        RECT 7.680 3.480 7.850 3.650 ;
        RECT -6.900 2.660 -6.730 2.830 ;
        RECT -4.690 2.770 -4.420 3.040 ;
        RECT -2.970 2.800 -2.800 2.970 ;
        RECT -7.810 2.320 -7.640 2.490 ;
        RECT -0.660 2.840 -0.390 3.110 ;
        RECT 0.430 2.840 0.700 3.110 ;
        RECT 2.840 3.160 3.010 3.330 ;
        RECT 2.840 2.800 3.010 2.970 ;
        RECT 4.460 2.770 4.730 3.040 ;
        RECT 6.770 3.020 6.940 3.190 ;
        RECT 9.130 2.900 9.310 3.070 ;
        RECT 6.770 2.660 6.940 2.830 ;
        RECT 7.680 2.320 7.850 2.490 ;
        RECT -9.620 2.060 -9.450 2.230 ;
        RECT -8.890 2.030 -8.720 2.200 ;
        RECT 8.760 2.030 8.930 2.200 ;
        RECT -7.810 1.770 -7.640 1.940 ;
        RECT 7.680 1.770 7.850 1.940 ;
        RECT 9.490 2.060 9.660 2.230 ;
        RECT -9.620 0.510 -9.450 0.680 ;
        RECT -7.810 0.800 -7.640 0.970 ;
        RECT 7.680 0.800 7.850 0.970 ;
        RECT -8.890 0.540 -8.720 0.710 ;
        RECT 8.760 0.540 8.930 0.710 ;
        RECT 9.490 0.510 9.660 0.680 ;
        RECT -7.810 0.250 -7.640 0.420 ;
        RECT 7.680 0.250 7.850 0.420 ;
      LAYER met1 ;
        RECT -7.890 5.490 -7.570 5.810 ;
        RECT 7.610 5.490 7.930 5.810 ;
        RECT -7.890 4.940 -7.570 5.260 ;
        RECT 7.610 4.940 7.930 5.260 ;
        RECT -7.890 3.950 -7.570 4.270 ;
        RECT 7.610 3.950 7.930 4.270 ;
        RECT -7.890 3.400 -7.570 3.720 ;
        RECT 7.610 3.400 7.930 3.720 ;
        RECT -7.890 2.250 -7.570 2.570 ;
        RECT 7.610 2.250 7.930 2.570 ;
        RECT -7.890 1.700 -7.570 2.020 ;
        RECT 7.610 1.700 7.930 2.020 ;
        RECT -7.890 0.720 -7.570 1.040 ;
        RECT 7.610 0.720 7.930 1.040 ;
        RECT -7.890 0.170 -7.570 0.490 ;
        RECT 7.610 0.170 7.930 0.490 ;
      LAYER via ;
        RECT -7.860 5.520 -7.600 5.780 ;
        RECT 7.640 5.520 7.900 5.780 ;
        RECT -7.860 4.970 -7.600 5.230 ;
        RECT 7.640 4.970 7.900 5.230 ;
        RECT -7.860 3.980 -7.600 4.240 ;
        RECT 7.640 3.980 7.900 4.240 ;
        RECT -7.860 3.430 -7.600 3.690 ;
        RECT 7.640 3.430 7.900 3.690 ;
        RECT -7.860 2.280 -7.600 2.540 ;
        RECT 7.640 2.280 7.900 2.540 ;
        RECT -7.860 1.730 -7.600 1.990 ;
        RECT 7.640 1.730 7.900 1.990 ;
        RECT -7.860 0.750 -7.600 1.010 ;
        RECT 7.640 0.750 7.900 1.010 ;
        RECT -7.860 0.200 -7.600 0.460 ;
        RECT 7.640 0.200 7.900 0.460 ;
  END
END sky130_hilas_swc4x2cell

MACRO sky130_hilas_polyresistorGND
  CLASS BLOCK ;
  FOREIGN sky130_hilas_polyresistorGND ;
  ORIGIN 27.490 0.570 ;
  SIZE 55.470 BY 10.890 ;
  PIN INPUT
    PORT
      LAYER met1 ;
        RECT -6.430 9.680 -4.020 10.320 ;
        RECT -6.410 8.330 -6.000 9.680 ;
    END
  END INPUT
  PIN OUTPUT
    ANTENNADIFFAREA 16.452000 ;
    PORT
      LAYER met2 ;
        RECT -27.490 6.810 27.980 8.200 ;
    END
  END OUTPUT
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.320 9.020 0.730 9.790 ;
        RECT 0.050 8.750 0.730 9.020 ;
        RECT 0.050 8.320 1.740 8.750 ;
        RECT -27.160 8.140 -2.790 8.160 ;
        RECT -27.220 7.750 -2.790 8.140 ;
        RECT -27.220 -0.500 -26.810 7.750 ;
        RECT -0.620 0.250 1.740 8.320 ;
        RECT 6.010 8.150 27.370 8.160 ;
        RECT 5.950 7.760 27.370 8.150 ;
        RECT 5.950 7.750 27.210 7.760 ;
        RECT -0.740 -0.570 1.740 0.250 ;
      LAYER via ;
        RECT -26.670 7.840 -2.870 8.100 ;
        RECT 6.010 7.840 26.870 8.100 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT -6.350 8.550 -6.130 9.670 ;
        RECT -6.400 8.360 -6.070 8.550 ;
        RECT 0.390 8.360 0.630 9.710 ;
        RECT -27.110 7.890 27.630 8.160 ;
        RECT -27.110 7.760 -2.770 7.890 ;
        RECT 5.920 7.760 27.630 7.890 ;
        RECT -27.110 0.160 -26.940 7.760 ;
        RECT 27.460 0.680 27.630 7.760 ;
        RECT -0.670 -0.180 1.690 -0.010 ;
      LAYER mcon ;
        RECT -6.320 9.470 -6.150 9.640 ;
        RECT -6.320 9.110 -6.150 9.280 ;
        RECT -6.320 8.750 -6.150 8.920 ;
        RECT -6.320 8.390 -6.150 8.560 ;
        RECT 0.430 9.300 0.600 9.470 ;
        RECT 0.430 8.940 0.600 9.110 ;
        RECT 0.430 8.580 0.600 8.750 ;
        RECT -26.770 7.780 -2.870 7.950 ;
        RECT 6.010 7.780 27.180 7.950 ;
        RECT -0.300 -0.180 -0.130 -0.010 ;
        RECT 0.070 -0.180 0.240 -0.010 ;
        RECT 0.430 -0.180 0.600 -0.010 ;
        RECT 0.790 -0.180 0.960 -0.010 ;
        RECT 1.150 -0.180 1.330 -0.010 ;
        RECT 1.520 -0.180 1.690 -0.010 ;
      LAYER met2 ;
        RECT -27.490 0.510 27.980 1.910 ;
  END
END sky130_hilas_polyresistorGND

MACRO sky130_hilas_swc4x2cellOverlap
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc4x2cellOverlap ;
  ORIGIN 10.010 -7.230 ;
  SIZE 17.980 BY 6.160 ;
  PIN VERT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met1 ;
        RECT -8.840 12.650 -8.680 13.380 ;
        RECT -8.880 12.630 -8.680 12.650 ;
        RECT -8.890 12.390 -8.660 12.630 ;
        RECT -8.890 12.340 -8.680 12.390 ;
        RECT -8.840 11.280 -8.680 12.340 ;
        RECT -8.890 11.230 -8.680 11.280 ;
        RECT -8.890 10.990 -8.660 11.230 ;
        RECT -8.880 10.970 -8.680 10.990 ;
        RECT -8.840 9.640 -8.680 10.970 ;
        RECT -8.880 9.620 -8.680 9.640 ;
        RECT -8.890 9.380 -8.660 9.620 ;
        RECT -8.890 9.330 -8.680 9.380 ;
        RECT -8.840 8.280 -8.680 9.330 ;
        RECT -8.890 8.230 -8.680 8.280 ;
        RECT -8.890 7.990 -8.660 8.230 ;
        RECT -8.880 7.970 -8.680 7.990 ;
        RECT -8.840 7.240 -8.680 7.970 ;
    END
  END VERT1
  PIN HORIZ1
    USE ANALOG ;
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT -7.850 12.400 -7.540 12.420 ;
        RECT 5.490 12.400 5.800 12.420 ;
        RECT -10.010 12.220 7.970 12.400 ;
        RECT -7.850 12.090 -7.540 12.220 ;
        RECT 5.490 12.090 5.800 12.220 ;
    END
  END HORIZ1
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT -7.850 12.830 -7.540 12.970 ;
        RECT 5.490 12.830 5.800 12.970 ;
        RECT -10.010 12.650 7.960 12.830 ;
        RECT -7.850 12.640 -7.540 12.650 ;
        RECT 5.490 12.640 5.800 12.650 ;
    END
  END DRAIN1
  PIN HORIZ2
    USE ANALOG ;
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT -7.850 11.400 -7.540 11.530 ;
        RECT 5.490 11.400 5.800 11.530 ;
        RECT -10.010 11.220 7.970 11.400 ;
        RECT -7.850 11.200 -7.540 11.220 ;
        RECT 5.490 11.200 5.800 11.220 ;
    END
  END HORIZ2
  PIN DRAIN2
    USE ANALOG ;
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT -7.850 10.970 -7.540 10.980 ;
        RECT 5.490 10.970 5.800 10.980 ;
        RECT -10.010 10.790 7.970 10.970 ;
        RECT -7.850 10.650 -7.540 10.790 ;
        RECT 5.490 10.650 5.800 10.790 ;
    END
  END DRAIN2
  PIN DRAIN3
    USE ANALOG ;
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT -7.850 9.820 -7.540 9.960 ;
        RECT -10.010 9.810 -7.540 9.820 ;
        RECT 5.490 9.820 5.800 9.960 ;
        RECT 5.490 9.810 7.960 9.820 ;
        RECT -10.010 9.640 7.960 9.810 ;
        RECT -7.850 9.630 -7.540 9.640 ;
        RECT 5.490 9.630 5.800 9.640 ;
    END
  END DRAIN3
  PIN HORIZ3
    USE ANALOG ;
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT -7.850 9.390 -7.540 9.410 ;
        RECT 5.490 9.390 5.800 9.410 ;
        RECT -10.010 9.220 7.960 9.390 ;
        RECT -10.010 9.210 -7.450 9.220 ;
        RECT 5.400 9.210 7.960 9.220 ;
        RECT -7.850 9.080 -7.540 9.210 ;
        RECT 5.490 9.080 5.800 9.210 ;
    END
  END HORIZ3
  PIN HORIZ4
    USE ANALOG ;
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT -7.850 8.410 -7.540 8.530 ;
        RECT 5.490 8.410 5.800 8.530 ;
        RECT -7.850 8.400 5.800 8.410 ;
        RECT -10.010 8.240 7.960 8.400 ;
        RECT -10.010 8.220 -7.450 8.240 ;
        RECT 5.400 8.220 7.960 8.240 ;
        RECT -7.850 8.200 -7.540 8.220 ;
        RECT 5.490 8.200 5.800 8.220 ;
    END
  END HORIZ4
  PIN DRAIN4
    USE ANALOG ;
    ANTENNADIFFAREA 0.230400 ;
    PORT
      LAYER met2 ;
        RECT -7.850 7.970 -7.540 7.980 ;
        RECT 5.490 7.970 5.800 7.980 ;
        RECT -10.010 7.800 7.960 7.970 ;
        RECT -10.010 7.790 -7.540 7.800 ;
        RECT -7.850 7.650 -7.540 7.790 ;
        RECT 5.490 7.790 7.960 7.800 ;
        RECT 5.490 7.650 5.800 7.790 ;
    END
  END DRAIN4
  PIN VINJ
    ANTENNADIFFAREA 1.088000 ;
    PORT
      LAYER nwell ;
        RECT -10.010 13.330 -7.450 13.390 ;
        RECT -10.010 7.280 -3.450 13.330 ;
        RECT -10.010 7.230 -7.450 7.280 ;
      LAYER met1 ;
        RECT -9.650 12.680 -9.490 13.380 ;
        RECT -9.650 12.130 -9.380 12.680 ;
        RECT -9.660 12.080 -9.380 12.130 ;
        RECT -9.660 11.990 -9.490 12.080 ;
        RECT -9.650 11.630 -9.490 11.990 ;
        RECT -9.660 11.540 -9.490 11.630 ;
        RECT -9.660 11.490 -9.380 11.540 ;
        RECT -9.650 10.940 -9.380 11.490 ;
        RECT -9.650 9.670 -9.490 10.940 ;
        RECT -9.650 9.120 -9.380 9.670 ;
        RECT -9.660 9.070 -9.380 9.120 ;
        RECT -9.660 8.980 -9.490 9.070 ;
        RECT -9.650 8.630 -9.490 8.980 ;
        RECT -9.660 8.540 -9.490 8.630 ;
        RECT -9.660 8.490 -9.380 8.540 ;
        RECT -9.650 7.940 -9.380 8.490 ;
        RECT -9.650 7.240 -9.490 7.940 ;
    END
    PORT
      LAYER nwell ;
        RECT 5.400 13.330 7.960 13.390 ;
        RECT 1.400 7.280 7.960 13.330 ;
        RECT 5.400 7.230 7.960 7.280 ;
      LAYER met1 ;
        RECT 7.440 12.680 7.600 13.380 ;
        RECT 7.330 12.130 7.600 12.680 ;
        RECT 7.330 12.080 7.610 12.130 ;
        RECT 7.440 11.990 7.610 12.080 ;
        RECT 7.440 11.630 7.600 11.990 ;
        RECT 7.440 11.540 7.610 11.630 ;
        RECT 7.330 11.490 7.610 11.540 ;
        RECT 7.330 10.940 7.600 11.490 ;
        RECT 7.440 9.670 7.600 10.940 ;
        RECT 7.330 9.120 7.600 9.670 ;
        RECT 7.330 9.070 7.610 9.120 ;
        RECT 7.440 8.980 7.610 9.070 ;
        RECT 7.440 8.630 7.600 8.980 ;
        RECT 7.440 8.540 7.610 8.630 ;
        RECT 7.330 8.490 7.610 8.540 ;
        RECT 7.330 7.940 7.600 8.490 ;
        RECT 7.440 7.240 7.600 7.940 ;
    END
  END VINJ
  PIN GATESELECT1
    USE ANALOG ;
    ANTENNAGATEAREA 0.720000 ;
    PORT
      LAYER met1 ;
        RECT -9.240 12.340 -9.050 13.330 ;
        RECT -9.240 12.220 -9.070 12.340 ;
        RECT -9.240 11.400 -9.080 12.220 ;
        RECT -9.240 11.280 -9.070 11.400 ;
        RECT -9.240 10.420 -9.050 11.280 ;
        RECT -9.270 10.190 -9.030 10.420 ;
        RECT -9.240 9.330 -9.050 10.190 ;
        RECT -9.240 9.210 -9.070 9.330 ;
        RECT -9.240 8.400 -9.080 9.210 ;
        RECT -9.240 8.280 -9.070 8.400 ;
        RECT -9.240 7.290 -9.050 8.280 ;
    END
  END GATESELECT1
  PIN VERT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met1 ;
        RECT 6.630 12.650 6.790 13.380 ;
        RECT 6.630 12.630 6.830 12.650 ;
        RECT 6.610 12.390 6.840 12.630 ;
        RECT 6.630 12.340 6.840 12.390 ;
        RECT 6.630 11.280 6.790 12.340 ;
        RECT 6.630 11.230 6.840 11.280 ;
        RECT 6.610 10.990 6.840 11.230 ;
        RECT 6.630 10.970 6.830 10.990 ;
        RECT 6.630 9.640 6.790 10.970 ;
        RECT 6.630 9.620 6.830 9.640 ;
        RECT 6.610 9.380 6.840 9.620 ;
        RECT 6.630 9.330 6.840 9.380 ;
        RECT 6.630 8.280 6.790 9.330 ;
        RECT 6.630 8.230 6.840 8.280 ;
        RECT 6.610 7.990 6.840 8.230 ;
        RECT 6.630 7.970 6.830 7.990 ;
        RECT 6.630 7.240 6.790 7.970 ;
    END
  END VERT2
  PIN GATESELECT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.720000 ;
    PORT
      LAYER met1 ;
        RECT 7.000 12.340 7.190 13.330 ;
        RECT 7.020 12.220 7.190 12.340 ;
        RECT 7.030 11.400 7.190 12.220 ;
        RECT 7.020 11.280 7.190 11.400 ;
        RECT 7.000 10.420 7.190 11.280 ;
        RECT 6.980 10.190 7.220 10.420 ;
        RECT 7.000 9.330 7.190 10.190 ;
        RECT 7.020 9.210 7.190 9.330 ;
        RECT 7.030 8.400 7.190 9.210 ;
        RECT 7.020 8.280 7.190 8.400 ;
        RECT 7.000 7.290 7.190 8.280 ;
    END
  END GATESELECT2
  PIN GATE2
    USE ANALOG ;
    ANTENNADIFFAREA 1.345600 ;
    PORT
      LAYER met1 ;
        RECT 3.280 12.100 3.520 13.330 ;
        RECT 3.280 11.880 3.530 12.100 ;
        RECT 3.280 10.630 3.520 11.880 ;
        RECT 3.280 10.410 3.530 10.630 ;
        RECT 3.280 9.160 3.520 10.410 ;
        RECT 3.280 8.940 3.530 9.160 ;
        RECT 3.280 7.690 3.520 8.940 ;
        RECT 3.280 7.470 3.530 7.690 ;
        RECT 3.280 7.280 3.520 7.470 ;
    END
  END GATE2
  PIN GATE1
    USE ANALOG ;
    ANTENNADIFFAREA 1.345600 ;
    PORT
      LAYER met1 ;
        RECT -5.570 12.100 -5.320 13.330 ;
        RECT -5.580 11.880 -5.320 12.100 ;
        RECT -5.570 10.630 -5.320 11.880 ;
        RECT -5.580 10.410 -5.320 10.630 ;
        RECT -5.570 9.160 -5.320 10.410 ;
        RECT -5.580 8.940 -5.320 9.160 ;
        RECT -5.570 7.690 -5.320 8.940 ;
        RECT -5.580 7.470 -5.320 7.690 ;
        RECT -5.570 7.280 -5.320 7.470 ;
    END
  END GATE1
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 0.336400 ;
    PORT
      LAYER met1 ;
        RECT -1.960 7.280 -1.660 13.330 ;
    END
    PORT
      LAYER met1 ;
        RECT -0.380 7.280 -0.080 13.330 ;
    END
  END VTUN
  OBS
      LAYER li1 ;
        RECT -9.610 12.650 -9.410 13.000 ;
        RECT -7.870 12.920 -7.550 12.930 ;
        RECT -8.130 12.750 -7.550 12.920 ;
        RECT -7.880 12.700 -7.550 12.750 ;
        RECT -7.870 12.670 -7.550 12.700 ;
        RECT -9.620 12.620 -9.410 12.650 ;
        RECT -9.620 12.030 -9.400 12.620 ;
        RECT -8.880 12.030 -8.680 12.630 ;
        RECT -7.870 12.340 -7.550 12.380 ;
        RECT -7.880 12.300 -7.550 12.340 ;
        RECT -8.130 12.130 -7.550 12.300 ;
        RECT -7.870 12.120 -7.550 12.130 ;
        RECT -7.110 12.020 -3.800 13.000 ;
        RECT -1.890 12.120 -1.720 13.010 ;
        RECT -0.330 12.120 -0.160 13.010 ;
        RECT 1.750 12.020 5.060 13.000 ;
        RECT 5.500 12.920 5.820 12.930 ;
        RECT 5.500 12.750 6.080 12.920 ;
        RECT 5.500 12.700 5.830 12.750 ;
        RECT 5.500 12.670 5.820 12.700 ;
        RECT 7.360 12.650 7.560 13.000 ;
        RECT 5.500 12.340 5.820 12.380 ;
        RECT 5.500 12.300 5.830 12.340 ;
        RECT 5.500 12.130 6.080 12.300 ;
        RECT 5.500 12.120 5.820 12.130 ;
        RECT 6.630 12.030 6.830 12.630 ;
        RECT 7.360 12.620 7.570 12.650 ;
        RECT 7.350 12.030 7.570 12.620 ;
        RECT -9.620 11.000 -9.400 11.590 ;
        RECT -9.620 10.970 -9.410 11.000 ;
        RECT -8.880 10.990 -8.680 11.590 ;
        RECT -7.870 11.490 -7.550 11.500 ;
        RECT -8.130 11.320 -7.550 11.490 ;
        RECT -7.880 11.280 -7.550 11.320 ;
        RECT -7.870 11.240 -7.550 11.280 ;
        RECT -9.610 10.620 -9.410 10.970 ;
        RECT -7.870 10.920 -7.550 10.950 ;
        RECT -7.880 10.870 -7.550 10.920 ;
        RECT -8.130 10.700 -7.550 10.870 ;
        RECT -7.870 10.690 -7.550 10.700 ;
        RECT -7.110 10.550 -3.800 11.530 ;
        RECT -1.890 10.600 -1.720 11.490 ;
        RECT -0.330 10.600 -0.160 11.490 ;
        RECT 1.750 10.550 5.060 11.530 ;
        RECT 5.500 11.490 5.820 11.500 ;
        RECT 5.500 11.320 6.080 11.490 ;
        RECT 5.500 11.280 5.830 11.320 ;
        RECT 5.500 11.240 5.820 11.280 ;
        RECT 6.630 10.990 6.830 11.590 ;
        RECT 7.350 11.000 7.570 11.590 ;
        RECT 7.360 10.970 7.570 11.000 ;
        RECT 5.500 10.920 5.820 10.950 ;
        RECT 5.500 10.870 5.830 10.920 ;
        RECT 5.500 10.700 6.080 10.870 ;
        RECT 5.500 10.690 5.820 10.700 ;
        RECT 7.360 10.620 7.560 10.970 ;
        RECT -9.240 10.220 -8.800 10.390 ;
        RECT 6.750 10.220 7.190 10.390 ;
        RECT -9.610 9.640 -9.410 9.990 ;
        RECT -7.870 9.910 -7.550 9.920 ;
        RECT -8.130 9.740 -7.550 9.910 ;
        RECT -7.880 9.690 -7.550 9.740 ;
        RECT -7.870 9.660 -7.550 9.690 ;
        RECT -9.620 9.610 -9.410 9.640 ;
        RECT -9.620 9.020 -9.400 9.610 ;
        RECT -8.880 9.020 -8.680 9.620 ;
        RECT -7.870 9.330 -7.550 9.370 ;
        RECT -7.880 9.290 -7.550 9.330 ;
        RECT -8.130 9.120 -7.550 9.290 ;
        RECT -7.870 9.110 -7.550 9.120 ;
        RECT -7.110 9.080 -3.800 10.060 ;
        RECT -1.890 9.150 -1.720 10.040 ;
        RECT -0.330 9.150 -0.160 10.040 ;
        RECT 1.750 9.080 5.060 10.060 ;
        RECT 5.500 9.910 5.820 9.920 ;
        RECT 5.500 9.740 6.080 9.910 ;
        RECT 5.500 9.690 5.830 9.740 ;
        RECT 5.500 9.660 5.820 9.690 ;
        RECT 7.360 9.640 7.560 9.990 ;
        RECT 5.500 9.330 5.820 9.370 ;
        RECT 5.500 9.290 5.830 9.330 ;
        RECT 5.500 9.120 6.080 9.290 ;
        RECT 5.500 9.110 5.820 9.120 ;
        RECT 6.630 9.020 6.830 9.620 ;
        RECT 7.360 9.610 7.570 9.640 ;
        RECT 7.350 9.020 7.570 9.610 ;
        RECT -9.620 8.000 -9.400 8.590 ;
        RECT -9.620 7.970 -9.410 8.000 ;
        RECT -8.880 7.990 -8.680 8.590 ;
        RECT -7.870 8.490 -7.550 8.500 ;
        RECT -8.130 8.320 -7.550 8.490 ;
        RECT -7.880 8.280 -7.550 8.320 ;
        RECT -7.870 8.240 -7.550 8.280 ;
        RECT -9.610 7.620 -9.410 7.970 ;
        RECT -7.870 7.920 -7.550 7.950 ;
        RECT -7.880 7.870 -7.550 7.920 ;
        RECT -8.130 7.700 -7.550 7.870 ;
        RECT -7.870 7.690 -7.550 7.700 ;
        RECT -7.110 7.610 -3.800 8.590 ;
        RECT -1.890 7.610 -1.720 8.500 ;
        RECT -0.330 7.610 -0.160 8.500 ;
        RECT 1.750 7.610 5.060 8.590 ;
        RECT 5.500 8.490 5.820 8.500 ;
        RECT 5.500 8.320 6.080 8.490 ;
        RECT 5.500 8.280 5.830 8.320 ;
        RECT 5.500 8.240 5.820 8.280 ;
        RECT 6.630 7.990 6.830 8.590 ;
        RECT 7.350 8.000 7.570 8.590 ;
        RECT 7.360 7.970 7.570 8.000 ;
        RECT 5.500 7.920 5.820 7.950 ;
        RECT 5.500 7.870 5.830 7.920 ;
        RECT 5.500 7.700 6.080 7.870 ;
        RECT 5.500 7.690 5.820 7.700 ;
        RECT 7.360 7.620 7.560 7.970 ;
      LAYER mcon ;
        RECT -7.780 12.710 -7.610 12.880 ;
        RECT -5.540 12.770 -5.370 12.940 ;
        RECT -9.590 12.450 -9.420 12.620 ;
        RECT -8.860 12.420 -8.690 12.590 ;
        RECT -7.780 12.160 -7.610 12.330 ;
        RECT -5.540 12.080 -5.370 12.250 ;
        RECT -1.890 12.810 -1.720 12.980 ;
        RECT -0.330 12.810 -0.160 12.980 ;
        RECT 3.320 12.770 3.490 12.940 ;
        RECT 5.560 12.710 5.730 12.880 ;
        RECT 6.640 12.420 6.810 12.590 ;
        RECT 3.320 12.080 3.490 12.250 ;
        RECT 5.560 12.160 5.730 12.330 ;
        RECT 7.370 12.450 7.540 12.620 ;
        RECT -9.590 11.000 -9.420 11.170 ;
        RECT -7.780 11.290 -7.610 11.460 ;
        RECT -5.540 11.300 -5.370 11.470 ;
        RECT -8.860 11.030 -8.690 11.200 ;
        RECT -7.780 10.740 -7.610 10.910 ;
        RECT -5.540 10.610 -5.370 10.780 ;
        RECT -1.890 11.290 -1.720 11.460 ;
        RECT -0.330 11.290 -0.160 11.460 ;
        RECT 3.320 11.300 3.490 11.470 ;
        RECT 5.560 11.290 5.730 11.460 ;
        RECT 6.640 11.030 6.810 11.200 ;
        RECT 7.370 11.000 7.540 11.170 ;
        RECT 3.320 10.610 3.490 10.780 ;
        RECT 5.560 10.740 5.730 10.910 ;
        RECT 7.010 10.220 7.190 10.390 ;
        RECT -7.780 9.700 -7.610 9.870 ;
        RECT -5.540 9.830 -5.370 10.000 ;
        RECT -9.590 9.440 -9.420 9.610 ;
        RECT -8.860 9.410 -8.690 9.580 ;
        RECT -7.780 9.150 -7.610 9.320 ;
        RECT -5.540 9.140 -5.370 9.310 ;
        RECT -1.890 9.840 -1.720 10.010 ;
        RECT -0.330 9.840 -0.160 10.010 ;
        RECT 3.320 9.830 3.490 10.000 ;
        RECT 5.560 9.700 5.730 9.870 ;
        RECT 6.640 9.410 6.810 9.580 ;
        RECT 3.320 9.140 3.490 9.310 ;
        RECT 5.560 9.150 5.730 9.320 ;
        RECT 7.370 9.440 7.540 9.610 ;
        RECT -9.590 8.000 -9.420 8.170 ;
        RECT -7.780 8.290 -7.610 8.460 ;
        RECT -5.540 8.360 -5.370 8.530 ;
        RECT -8.860 8.030 -8.690 8.200 ;
        RECT -7.780 7.740 -7.610 7.910 ;
        RECT -5.540 7.670 -5.370 7.840 ;
        RECT -1.890 8.300 -1.720 8.470 ;
        RECT -0.330 8.300 -0.160 8.470 ;
        RECT 3.320 8.360 3.490 8.530 ;
        RECT 5.560 8.290 5.730 8.460 ;
        RECT 6.640 8.030 6.810 8.200 ;
        RECT 7.370 8.000 7.540 8.170 ;
        RECT 3.320 7.670 3.490 7.840 ;
        RECT 5.560 7.740 5.730 7.910 ;
      LAYER met1 ;
        RECT -7.860 12.640 -7.540 12.960 ;
        RECT 5.490 12.640 5.810 12.960 ;
        RECT -7.860 12.090 -7.540 12.410 ;
        RECT 5.490 12.090 5.810 12.410 ;
        RECT -7.860 11.210 -7.540 11.530 ;
        RECT 5.490 11.210 5.810 11.530 ;
        RECT -7.860 10.660 -7.540 10.980 ;
        RECT 5.490 10.660 5.810 10.980 ;
        RECT -7.860 9.630 -7.540 9.950 ;
        RECT 5.490 9.630 5.810 9.950 ;
        RECT -7.860 9.080 -7.540 9.400 ;
        RECT 5.490 9.080 5.810 9.400 ;
        RECT -7.860 8.210 -7.540 8.530 ;
        RECT 5.490 8.210 5.810 8.530 ;
        RECT -7.860 7.660 -7.540 7.980 ;
        RECT 5.490 7.660 5.810 7.980 ;
      LAYER via ;
        RECT -7.830 12.670 -7.570 12.930 ;
        RECT 5.520 12.670 5.780 12.930 ;
        RECT -7.830 12.120 -7.570 12.380 ;
        RECT 5.520 12.120 5.780 12.380 ;
        RECT -7.830 11.240 -7.570 11.500 ;
        RECT 5.520 11.240 5.780 11.500 ;
        RECT -7.830 10.690 -7.570 10.950 ;
        RECT 5.520 10.690 5.780 10.950 ;
        RECT -7.830 9.660 -7.570 9.920 ;
        RECT 5.520 9.660 5.780 9.920 ;
        RECT -7.830 9.110 -7.570 9.370 ;
        RECT 5.520 9.110 5.780 9.370 ;
        RECT -7.830 8.240 -7.570 8.500 ;
        RECT 5.520 8.240 5.780 8.500 ;
        RECT -7.830 7.690 -7.570 7.950 ;
        RECT 5.520 7.690 5.780 7.950 ;
  END
END sky130_hilas_swc4x2cellOverlap

MACRO sky130_hilas_FGBias2x1cell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_FGBias2x1cell ;
  ORIGIN 3.960 3.870 ;
  SIZE 11.530 BY 6.150 ;
  PIN VTUN
    USE ANALOG ;
    ANTENNADIFFAREA 2.516100 ;
    PORT
      LAYER nwell ;
        RECT -3.950 1.480 -2.220 2.230 ;
        RECT -3.950 0.330 -2.210 1.480 ;
        RECT -3.940 -1.910 -2.210 0.330 ;
        RECT -3.950 -2.090 -2.210 -1.910 ;
        RECT -3.950 -3.810 -2.220 -2.090 ;
      LAYER met1 ;
        RECT -3.610 -3.820 -3.190 2.230 ;
    END
  END VTUN
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT -1.130 -3.820 -0.900 2.230 ;
    END
  END VGND
  PIN GATE_CONTROL
    USE ANALOG ;
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT -0.190 -0.160 2.530 1.490 ;
        RECT -0.190 -0.200 2.520 -0.160 ;
        RECT -0.190 -1.530 2.520 -1.490 ;
        RECT -0.190 -3.180 2.530 -1.530 ;
      LAYER met1 ;
        RECT 0.090 1.020 0.320 2.230 ;
        RECT 0.090 0.230 0.350 1.020 ;
        RECT 0.090 -1.920 0.320 0.230 ;
        RECT 0.090 -2.710 0.350 -1.920 ;
        RECT 0.090 -3.820 0.320 -2.710 ;
    END
  END GATE_CONTROL
  PIN DRAIN1
    USE ANALOG ;
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 5.090 1.730 5.400 1.740 ;
        RECT -3.960 1.550 7.570 1.730 ;
        RECT 5.090 1.410 5.400 1.550 ;
    END
  END DRAIN1
  PIN DRAIN4
    USE ANALOG ;
    ANTENNADIFFAREA 0.122400 ;
    PORT
      LAYER met2 ;
        RECT 5.090 -3.140 5.400 -3.000 ;
        RECT 5.090 -3.150 7.570 -3.140 ;
        RECT -3.960 -3.300 7.570 -3.150 ;
        RECT 5.090 -3.320 7.570 -3.300 ;
        RECT 5.090 -3.330 5.400 -3.320 ;
    END
  END DRAIN4
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 4.260 -3.870 7.570 2.280 ;
      LAYER met2 ;
        RECT 6.180 -0.630 6.500 -0.370 ;
        RECT 6.220 -0.650 7.400 -0.630 ;
        RECT 6.220 -0.910 7.440 -0.650 ;
        RECT 6.220 -0.970 7.400 -0.910 ;
        RECT 6.180 -0.980 7.400 -0.970 ;
        RECT 6.180 -1.230 6.500 -0.980 ;
    END
  END VINJ
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 5.240 0.710 5.550 0.780 ;
        RECT 5.240 0.490 7.570 0.710 ;
        RECT 5.240 0.450 5.550 0.490 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.588800 ;
    PORT
      LAYER met2 ;
        RECT 5.240 -2.050 5.550 -1.980 ;
        RECT 5.240 -2.260 7.570 -2.050 ;
        RECT 5.240 -2.310 5.550 -2.260 ;
    END
  END OUTPUT2
  PIN GATECOL
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT 6.610 0.770 6.800 2.230 ;
        RECT 6.610 0.740 6.830 0.770 ;
        RECT 6.590 0.470 6.840 0.740 ;
        RECT 6.600 0.460 6.840 0.470 ;
        RECT 6.600 0.220 6.830 0.460 ;
        RECT 6.640 -1.810 6.800 0.220 ;
        RECT 6.600 -2.050 6.830 -1.810 ;
        RECT 6.600 -2.060 6.840 -2.050 ;
        RECT 6.590 -2.330 6.840 -2.060 ;
        RECT 6.610 -2.360 6.830 -2.330 ;
        RECT 6.610 -3.820 6.800 -2.360 ;
    END
  END GATECOL
  PIN VINJ
    ANTENNADIFFAREA 0.544000 ;
    PORT
      LAYER met1 ;
        RECT 7.050 1.580 7.330 2.230 ;
        RECT 6.940 0.980 7.330 1.580 ;
        RECT 7.050 -0.620 7.330 0.980 ;
        RECT 7.050 -0.940 7.410 -0.620 ;
        RECT 7.050 -2.570 7.330 -0.940 ;
        RECT 6.940 -3.170 7.330 -2.570 ;
        RECT 7.050 -3.820 7.330 -3.170 ;
      LAYER via ;
        RECT 7.150 -0.910 7.410 -0.650 ;
    END
  END VINJ
  OBS
      LAYER li1 ;
        RECT 5.160 1.650 5.690 1.820 ;
        RECT 6.970 1.550 7.170 1.900 ;
        RECT 6.970 1.520 7.180 1.550 ;
        RECT -3.520 0.090 -2.970 0.520 ;
        RECT 0.110 0.280 0.340 0.970 ;
        RECT 5.410 0.740 5.580 1.260 ;
        RECT 5.250 0.480 5.580 0.740 ;
        RECT -0.920 -0.740 -0.730 -0.340 ;
        RECT 5.410 -0.430 5.580 0.480 ;
        RECT 6.240 -0.340 6.410 1.270 ;
        RECT 6.960 0.940 7.180 1.520 ;
        RECT 6.970 0.930 7.180 0.940 ;
        RECT 6.610 0.760 6.800 0.770 ;
        RECT 6.610 0.470 6.810 0.760 ;
        RECT 6.600 0.140 6.890 0.470 ;
        RECT 6.240 -0.530 6.420 -0.340 ;
        RECT -1.110 -0.750 -0.730 -0.740 ;
        RECT -1.110 -0.930 2.630 -0.750 ;
        RECT -1.110 -0.970 -0.730 -0.930 ;
        RECT -3.520 -1.640 -2.970 -1.210 ;
        RECT -0.920 -1.350 -0.730 -0.970 ;
        RECT 0.110 -2.660 0.340 -1.930 ;
        RECT 5.410 -2.020 5.580 -1.160 ;
        RECT 5.250 -2.280 5.580 -2.020 ;
        RECT 5.410 -2.850 5.580 -2.280 ;
        RECT 6.240 -1.250 6.420 -1.060 ;
        RECT 6.240 -2.860 6.410 -1.250 ;
        RECT 6.600 -2.060 6.890 -1.730 ;
        RECT 6.610 -2.350 6.810 -2.060 ;
        RECT 6.610 -2.360 6.800 -2.350 ;
        RECT 6.970 -2.530 7.180 -2.520 ;
        RECT 6.960 -3.110 7.180 -2.530 ;
        RECT 6.970 -3.140 7.180 -3.110 ;
        RECT 5.160 -3.410 5.690 -3.240 ;
        RECT 6.970 -3.490 7.170 -3.140 ;
      LAYER mcon ;
        RECT 6.980 1.350 7.150 1.520 ;
        RECT 0.140 0.770 0.310 0.940 ;
        RECT -3.520 0.170 -3.250 0.440 ;
        RECT 0.140 0.320 0.310 0.490 ;
        RECT 5.310 0.520 5.480 0.690 ;
        RECT 6.620 0.510 6.800 0.700 ;
        RECT -1.100 -0.940 -0.930 -0.770 ;
        RECT -3.520 -1.560 -3.250 -1.290 ;
        RECT 0.140 -2.180 0.310 -2.010 ;
        RECT 5.310 -2.240 5.480 -2.070 ;
        RECT 0.140 -2.630 0.310 -2.460 ;
        RECT 6.620 -2.290 6.800 -2.100 ;
        RECT 6.980 -3.110 7.150 -2.940 ;
      LAYER met1 ;
        RECT 5.090 1.410 5.400 1.850 ;
        RECT 5.240 0.450 5.560 0.770 ;
        RECT 6.210 -0.340 6.450 -0.210 ;
        RECT 6.210 -0.660 6.470 -0.340 ;
        RECT 6.210 -1.260 6.470 -0.940 ;
        RECT 6.210 -1.380 6.450 -1.260 ;
        RECT 5.240 -2.310 5.560 -1.990 ;
        RECT 5.090 -3.440 5.400 -3.000 ;
      LAYER via ;
        RECT 5.120 1.440 5.380 1.700 ;
        RECT 5.270 0.480 5.530 0.740 ;
        RECT 6.210 -0.630 6.470 -0.370 ;
        RECT 6.210 -1.230 6.470 -0.970 ;
        RECT 5.270 -2.280 5.530 -2.020 ;
        RECT 5.120 -3.290 5.380 -3.030 ;
  END
END sky130_hilas_FGBias2x1cell

MACRO sky130_hilas_drainSelect01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_drainSelect01 ;
  ORIGIN -10.500 0.280 ;
  SIZE 5.720 BY 6.590 ;
  PIN DRAIN3
    ANTENNADIFFAREA 0.322600 ;
    PORT
      LAYER met2 ;
        RECT 12.250 2.680 12.570 2.700 ;
        RECT 14.660 2.680 14.980 2.730 ;
        RECT 10.500 2.580 11.070 2.590 ;
        RECT 10.500 2.570 11.770 2.580 ;
        RECT 12.250 2.570 14.980 2.680 ;
        RECT 10.500 2.490 14.980 2.570 ;
        RECT 10.500 2.440 12.570 2.490 ;
        RECT 10.500 2.410 12.500 2.440 ;
        RECT 14.660 2.410 14.980 2.490 ;
    END
  END DRAIN3
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 10.500 -0.280 13.920 6.310 ;
      LAYER met1 ;
        RECT 11.080 6.040 11.330 6.260 ;
        RECT 10.690 4.970 11.330 6.040 ;
        RECT 11.080 4.260 11.330 4.970 ;
        RECT 10.690 3.190 11.330 4.260 ;
        RECT 11.080 2.840 11.330 3.190 ;
        RECT 10.690 1.770 11.330 2.840 ;
        RECT 11.080 1.060 11.330 1.770 ;
        RECT 10.690 -0.010 11.330 1.060 ;
        RECT 11.080 -0.230 11.330 -0.010 ;
    END
  END VINJ
  PIN DRAIN_MUX
    USE ANALOG ;
    ANTENNADIFFAREA 0.846400 ;
    PORT
      LAYER met1 ;
        RECT 14.070 -0.230 14.300 6.260 ;
    END
  END DRAIN_MUX
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 15.420 6.040 15.610 6.260 ;
        RECT 15.420 5.550 15.890 6.040 ;
        RECT 15.420 5.290 15.610 5.550 ;
        RECT 15.380 5.000 15.610 5.290 ;
        RECT 15.420 4.230 15.610 5.000 ;
        RECT 15.380 3.940 15.610 4.230 ;
        RECT 15.420 3.680 15.610 3.940 ;
        RECT 15.420 3.190 15.890 3.680 ;
        RECT 15.420 2.840 15.610 3.190 ;
        RECT 15.420 2.350 15.890 2.840 ;
        RECT 15.420 2.090 15.610 2.350 ;
        RECT 15.380 1.800 15.610 2.090 ;
        RECT 15.420 1.030 15.610 1.800 ;
        RECT 15.380 0.740 15.610 1.030 ;
        RECT 15.420 0.480 15.610 0.740 ;
        RECT 15.420 -0.010 15.890 0.480 ;
        RECT 15.420 -0.230 15.610 -0.010 ;
    END
  END VGND
  PIN SELECT2
    ANTENNAGATEAREA 0.730000 ;
    PORT
      LAYER met2 ;
        RECT 15.740 4.070 16.080 4.130 ;
        RECT 15.740 3.830 16.220 4.070 ;
    END
  END SELECT2
  PIN SELECT1
    ANTENNAGATEAREA 0.730000 ;
    PORT
      LAYER met2 ;
        RECT 15.740 5.170 16.220 5.400 ;
        RECT 15.740 5.100 16.080 5.170 ;
    END
  END SELECT1
  PIN SELECT3
    ANTENNAGATEAREA 0.730000 ;
    PORT
      LAYER met2 ;
        RECT 15.740 1.970 16.220 2.200 ;
        RECT 15.740 1.900 16.080 1.970 ;
    END
  END SELECT3
  PIN SELECT4
    ANTENNAGATEAREA 0.730000 ;
    PORT
      LAYER met2 ;
        RECT 15.740 0.860 16.080 0.930 ;
        RECT 15.740 0.630 16.220 0.860 ;
    END
  END SELECT4
  OBS
      LAYER li1 ;
        RECT 10.720 5.090 10.890 5.980 ;
        RECT 11.120 5.000 11.290 5.930 ;
        RECT 14.810 5.860 15.050 5.890 ;
        RECT 11.820 5.690 12.780 5.860 ;
        RECT 13.230 5.690 14.570 5.860 ;
        RECT 14.810 5.690 15.380 5.860 ;
        RECT 12.100 5.680 12.270 5.690 ;
        RECT 14.810 5.650 15.050 5.690 ;
        RECT 15.690 5.560 15.860 5.980 ;
        RECT 12.300 5.240 12.640 5.420 ;
        RECT 15.760 5.340 15.930 5.380 ;
        RECT 15.400 5.240 15.590 5.260 ;
        RECT 11.820 5.070 14.570 5.240 ;
        RECT 15.030 5.070 15.590 5.240 ;
        RECT 15.400 5.030 15.590 5.070 ;
        RECT 15.760 5.170 15.990 5.340 ;
        RECT 15.760 4.820 15.930 5.170 ;
        RECT 10.720 3.250 10.890 4.140 ;
        RECT 11.120 3.300 11.290 4.230 ;
        RECT 15.400 4.160 15.590 4.200 ;
        RECT 11.820 3.990 14.570 4.160 ;
        RECT 15.030 3.990 15.590 4.160 ;
        RECT 12.300 3.810 12.640 3.990 ;
        RECT 15.400 3.970 15.590 3.990 ;
        RECT 15.760 4.060 15.930 4.410 ;
        RECT 15.760 3.890 15.990 4.060 ;
        RECT 15.760 3.850 15.930 3.890 ;
        RECT 12.100 3.540 12.270 3.550 ;
        RECT 14.810 3.540 15.050 3.580 ;
        RECT 11.820 3.370 12.780 3.540 ;
        RECT 13.230 3.370 14.570 3.540 ;
        RECT 14.810 3.370 15.380 3.540 ;
        RECT 14.810 3.340 15.050 3.370 ;
        RECT 15.690 3.250 15.860 3.670 ;
        RECT 10.720 1.890 10.890 2.780 ;
        RECT 11.120 1.800 11.290 2.730 ;
        RECT 14.810 2.660 15.050 2.690 ;
        RECT 11.820 2.490 12.780 2.660 ;
        RECT 13.230 2.490 14.570 2.660 ;
        RECT 14.810 2.490 15.380 2.660 ;
        RECT 12.100 2.480 12.270 2.490 ;
        RECT 14.810 2.450 15.050 2.490 ;
        RECT 15.690 2.360 15.860 2.780 ;
        RECT 12.300 2.040 12.640 2.220 ;
        RECT 15.760 2.140 15.930 2.180 ;
        RECT 15.400 2.040 15.590 2.060 ;
        RECT 11.820 1.870 14.570 2.040 ;
        RECT 15.030 1.870 15.590 2.040 ;
        RECT 15.400 1.830 15.590 1.870 ;
        RECT 15.760 1.970 15.990 2.140 ;
        RECT 15.760 1.620 15.930 1.970 ;
        RECT 10.720 0.050 10.890 0.940 ;
        RECT 11.120 0.100 11.290 1.030 ;
        RECT 15.400 0.960 15.590 1.000 ;
        RECT 11.820 0.790 14.570 0.960 ;
        RECT 15.030 0.790 15.590 0.960 ;
        RECT 12.300 0.610 12.640 0.790 ;
        RECT 15.400 0.770 15.590 0.790 ;
        RECT 15.760 0.860 15.930 1.210 ;
        RECT 15.760 0.690 15.990 0.860 ;
        RECT 15.760 0.650 15.930 0.690 ;
        RECT 12.100 0.340 12.270 0.350 ;
        RECT 14.810 0.340 15.050 0.380 ;
        RECT 11.820 0.170 12.780 0.340 ;
        RECT 13.230 0.170 14.570 0.340 ;
        RECT 14.810 0.170 15.380 0.340 ;
        RECT 14.810 0.140 15.050 0.170 ;
        RECT 15.690 0.050 15.860 0.470 ;
      LAYER mcon ;
        RECT 10.720 5.810 10.890 5.980 ;
        RECT 10.720 5.450 10.890 5.620 ;
        RECT 14.100 5.690 14.270 5.860 ;
        RECT 14.850 5.690 15.020 5.860 ;
        RECT 15.690 5.810 15.860 5.980 ;
        RECT 11.120 5.360 11.290 5.530 ;
        RECT 15.410 5.060 15.580 5.230 ;
        RECT 15.820 5.170 15.990 5.340 ;
        RECT 10.720 3.970 10.890 4.140 ;
        RECT 10.720 3.610 10.890 3.780 ;
        RECT 15.410 4.000 15.580 4.170 ;
        RECT 11.120 3.700 11.290 3.870 ;
        RECT 15.820 3.890 15.990 4.060 ;
        RECT 12.100 3.380 12.270 3.550 ;
        RECT 14.100 3.370 14.270 3.540 ;
        RECT 14.850 3.370 15.020 3.540 ;
        RECT 10.720 2.610 10.890 2.780 ;
        RECT 10.720 2.250 10.890 2.420 ;
        RECT 14.100 2.490 14.270 2.660 ;
        RECT 14.850 2.490 15.020 2.660 ;
        RECT 15.690 2.610 15.860 2.780 ;
        RECT 11.120 2.160 11.290 2.330 ;
        RECT 15.410 1.860 15.580 2.030 ;
        RECT 15.820 1.970 15.990 2.140 ;
        RECT 10.720 0.770 10.890 0.940 ;
        RECT 10.720 0.410 10.890 0.580 ;
        RECT 15.410 0.800 15.580 0.970 ;
        RECT 11.120 0.500 11.290 0.670 ;
        RECT 15.820 0.690 15.990 0.860 ;
        RECT 12.100 0.180 12.270 0.350 ;
        RECT 14.100 0.170 14.270 0.340 ;
        RECT 14.850 0.170 15.020 0.340 ;
      LAYER met1 ;
        RECT 12.230 5.880 12.570 5.930 ;
        RECT 12.010 5.860 12.570 5.880 ;
        RECT 14.660 5.900 15.030 5.920 ;
        RECT 12.010 5.690 12.690 5.860 ;
        RECT 12.010 5.650 12.570 5.690 ;
        RECT 12.230 5.610 12.570 5.650 ;
        RECT 14.660 5.640 15.080 5.900 ;
        RECT 14.660 5.630 15.030 5.640 ;
        RECT 15.750 5.110 16.070 5.390 ;
        RECT 15.750 3.840 16.070 4.120 ;
        RECT 12.230 3.580 12.570 3.620 ;
        RECT 12.010 3.540 12.570 3.580 ;
        RECT 14.660 3.590 15.030 3.600 ;
        RECT 12.010 3.370 12.690 3.540 ;
        RECT 12.010 3.350 12.570 3.370 ;
        RECT 12.230 3.300 12.570 3.350 ;
        RECT 14.660 3.330 15.080 3.590 ;
        RECT 14.660 3.310 15.030 3.330 ;
        RECT 12.230 2.680 12.570 2.730 ;
        RECT 12.010 2.660 12.570 2.680 ;
        RECT 14.660 2.700 15.030 2.720 ;
        RECT 12.010 2.490 12.690 2.660 ;
        RECT 12.010 2.450 12.570 2.490 ;
        RECT 12.230 2.410 12.570 2.450 ;
        RECT 14.660 2.440 15.080 2.700 ;
        RECT 14.660 2.430 15.030 2.440 ;
        RECT 15.750 1.910 16.070 2.190 ;
        RECT 15.750 0.640 16.070 0.920 ;
        RECT 12.230 0.380 12.570 0.420 ;
        RECT 12.010 0.340 12.570 0.380 ;
        RECT 14.660 0.390 15.030 0.400 ;
        RECT 12.010 0.170 12.690 0.340 ;
        RECT 12.010 0.150 12.570 0.170 ;
        RECT 12.230 0.100 12.570 0.150 ;
        RECT 14.660 0.130 15.080 0.390 ;
        RECT 14.660 0.110 15.030 0.130 ;
      LAYER via ;
        RECT 12.280 5.640 12.540 5.900 ;
        RECT 14.690 5.640 14.950 5.900 ;
        RECT 15.780 5.120 16.040 5.380 ;
        RECT 15.780 3.850 16.040 4.110 ;
        RECT 12.280 3.330 12.540 3.590 ;
        RECT 14.690 3.330 14.950 3.590 ;
        RECT 12.280 2.440 12.540 2.700 ;
        RECT 14.690 2.440 14.950 2.700 ;
        RECT 15.780 1.920 16.040 2.180 ;
        RECT 15.780 0.650 16.040 0.910 ;
        RECT 12.280 0.130 12.540 0.390 ;
        RECT 14.690 0.130 14.950 0.390 ;
      LAYER met2 ;
        RECT 12.250 5.880 12.570 5.900 ;
        RECT 14.660 5.880 14.980 5.930 ;
        RECT 12.250 5.850 14.980 5.880 ;
        RECT 10.500 5.690 14.980 5.850 ;
        RECT 10.500 5.670 12.570 5.690 ;
        RECT 12.250 5.640 12.570 5.670 ;
        RECT 14.660 5.610 14.980 5.690 ;
        RECT 12.250 3.540 12.570 3.590 ;
        RECT 14.660 3.540 14.980 3.620 ;
        RECT 12.250 3.530 14.980 3.540 ;
        RECT 10.500 3.370 14.980 3.530 ;
        RECT 12.250 3.350 14.980 3.370 ;
        RECT 12.250 3.330 12.570 3.350 ;
        RECT 14.660 3.300 14.980 3.350 ;
        RECT 12.250 0.340 12.570 0.390 ;
        RECT 14.660 0.340 14.980 0.420 ;
        RECT 12.250 0.320 14.980 0.340 ;
        RECT 10.500 0.150 14.980 0.320 ;
        RECT 12.250 0.130 12.570 0.150 ;
        RECT 14.660 0.100 14.980 0.150 ;
  END
END sky130_hilas_drainSelect01

MACRO sky130_hilas_DAC5bit01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_DAC5bit01 ;
  ORIGIN -3.820 -5.240 ;
  SIZE 16.580 BY 5.990 ;
  PIN A0
    USE ANALOG ;
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER met2 ;
        RECT 12.080 6.230 12.400 6.260 ;
        RECT 3.820 6.030 12.400 6.230 ;
        RECT 12.080 6.000 12.400 6.030 ;
    END
  END A0
  PIN A1
    USE ANALOG ;
    ANTENNAGATEAREA 0.456300 ;
    PORT
      LAYER met2 ;
        RECT 15.410 10.910 15.730 11.230 ;
        RECT 15.530 7.350 15.680 10.910 ;
        RECT 3.820 7.150 15.690 7.350 ;
        RECT 3.820 7.140 3.960 7.150 ;
    END
  END A1
  PIN A2
    USE ANALOG ;
    ANTENNAGATEAREA 0.608400 ;
    PORT
      LAYER met2 ;
        RECT 13.800 10.930 14.120 11.230 ;
        RECT 13.800 10.910 14.130 10.930 ;
        RECT 13.930 8.330 14.130 10.910 ;
        RECT 3.820 8.120 14.130 8.330 ;
    END
  END A2
  PIN A3
    USE ANALOG ;
    ANTENNAGATEAREA 2.281500 ;
    PORT
      LAYER met2 ;
        RECT 12.190 10.900 12.510 11.220 ;
        RECT 7.310 10.660 7.630 10.810 ;
        RECT 7.300 10.490 7.630 10.660 ;
        RECT 3.820 10.200 5.880 10.260 ;
        RECT 7.300 10.200 7.520 10.490 ;
        RECT 12.220 10.210 12.470 10.900 ;
        RECT 12.220 10.200 12.500 10.210 ;
        RECT 3.820 10.050 12.500 10.200 ;
        RECT 4.080 9.870 4.280 10.050 ;
        RECT 5.720 9.900 12.500 10.050 ;
        RECT 4.030 9.550 4.350 9.870 ;
    END
  END A3
  PIN A4
    USE ANALOG ;
    ANTENNAGATEAREA 3.650400 ;
    PORT
      LAYER met2 ;
        RECT 5.760 11.210 6.080 11.220 ;
        RECT 8.960 11.210 9.280 11.220 ;
        RECT 10.570 11.210 10.890 11.230 ;
        RECT 3.820 11.020 10.890 11.210 ;
        RECT 3.820 11.000 4.370 11.020 ;
        RECT 4.050 10.860 4.370 11.000 ;
        RECT 5.760 10.900 6.080 11.020 ;
        RECT 8.960 10.900 9.280 11.020 ;
        RECT 10.570 10.910 10.890 11.020 ;
    END
  END A4
  PIN VPWR
    USE ANALOG ;
    ANTENNADIFFAREA 3.264300 ;
    PORT
      LAYER met2 ;
        RECT 16.530 10.930 17.690 11.210 ;
        RECT 16.650 10.750 16.960 10.930 ;
        RECT 17.280 10.920 17.690 10.930 ;
        RECT 17.320 10.750 17.630 10.920 ;
    END
  END VPWR
  PIN OUT
    USE ANALOG ;
    ANTENNADIFFAREA 3.264300 ;
    PORT
      LAYER met1 ;
        RECT 6.830 5.480 7.060 5.530 ;
        RECT 8.450 5.480 8.680 5.530 ;
        RECT 10.050 5.480 10.280 5.530 ;
        RECT 11.670 5.480 11.900 5.530 ;
        RECT 13.270 5.480 13.500 5.530 ;
        RECT 14.890 5.480 15.120 5.530 ;
        RECT 16.490 5.480 16.720 5.530 ;
        RECT 18.100 5.480 18.330 5.530 ;
        RECT 6.830 5.250 20.400 5.480 ;
        RECT 6.830 5.240 7.060 5.250 ;
        RECT 8.450 5.240 8.680 5.250 ;
        RECT 10.050 5.240 10.280 5.250 ;
        RECT 11.670 5.240 11.900 5.250 ;
        RECT 13.270 5.240 13.500 5.250 ;
        RECT 14.890 5.240 15.120 5.250 ;
        RECT 16.490 5.240 16.720 5.250 ;
        RECT 18.100 5.240 18.330 5.250 ;
    END
  END OUT
  OBS
      LAYER nwell ;
        RECT 4.190 5.270 20.290 10.920 ;
      LAYER li1 ;
        RECT 4.100 10.710 4.310 11.140 ;
        RECT 5.810 10.750 6.020 11.180 ;
        RECT 5.830 10.730 6.000 10.750 ;
        RECT 7.160 10.740 7.590 10.760 ;
        RECT 9.010 10.750 9.220 11.180 ;
        RECT 10.620 10.760 10.830 11.190 ;
        RECT 4.120 10.690 4.290 10.710 ;
        RECT 7.140 10.570 7.590 10.740 ;
        RECT 9.030 10.730 9.200 10.750 ;
        RECT 10.640 10.740 10.810 10.760 ;
        RECT 12.240 10.750 12.450 11.180 ;
        RECT 13.850 10.760 14.060 11.190 ;
        RECT 15.460 10.760 15.670 11.190 ;
        RECT 16.770 11.040 16.980 11.050 ;
        RECT 16.660 11.000 16.980 11.040 ;
        RECT 17.330 11.000 17.650 11.040 ;
        RECT 16.660 10.810 16.990 11.000 ;
        RECT 17.330 10.810 17.660 11.000 ;
        RECT 16.660 10.780 16.980 10.810 ;
        RECT 17.330 10.780 17.650 10.810 ;
        RECT 12.260 10.730 12.430 10.750 ;
        RECT 13.870 10.740 14.040 10.760 ;
        RECT 15.480 10.740 15.650 10.760 ;
        RECT 7.160 10.550 7.590 10.570 ;
        RECT 7.800 10.270 7.970 10.280 ;
        RECT 16.770 10.270 16.980 10.780 ;
        RECT 17.440 10.270 17.610 10.780 ;
        RECT 6.190 10.040 17.620 10.270 ;
        RECT 4.080 9.400 4.290 9.830 ;
        RECT 6.190 9.700 6.360 10.040 ;
        RECT 4.100 9.380 4.270 9.400 ;
        RECT 6.180 9.370 6.360 9.700 ;
        RECT 4.100 8.450 4.310 8.880 ;
        RECT 6.190 8.740 6.360 9.370 ;
        RECT 4.120 8.430 4.290 8.450 ;
        RECT 6.180 8.410 6.360 8.740 ;
        RECT 4.100 7.510 4.310 7.940 ;
        RECT 6.190 7.780 6.360 8.410 ;
        RECT 4.120 7.490 4.290 7.510 ;
        RECT 6.180 7.450 6.360 7.780 ;
        RECT 6.190 6.820 6.360 7.450 ;
        RECT 6.180 6.490 6.360 6.820 ;
        RECT 6.190 6.480 6.360 6.490 ;
        RECT 6.850 9.700 7.020 9.710 ;
        RECT 7.800 9.700 7.970 10.040 ;
        RECT 9.390 9.700 9.560 10.040 ;
        RECT 6.850 9.370 7.030 9.700 ;
        RECT 7.790 9.370 7.970 9.700 ;
        RECT 8.470 9.670 8.640 9.700 ;
        RECT 8.470 9.370 8.650 9.670 ;
        RECT 6.850 8.740 7.020 9.370 ;
        RECT 7.800 8.740 7.970 9.370 ;
        RECT 8.480 8.740 8.650 9.370 ;
        RECT 6.850 8.410 7.030 8.740 ;
        RECT 7.790 8.410 7.970 8.740 ;
        RECT 8.470 8.410 8.650 8.740 ;
        RECT 6.850 7.780 7.020 8.410 ;
        RECT 7.800 7.780 7.970 8.410 ;
        RECT 8.480 7.780 8.650 8.410 ;
        RECT 6.850 7.450 7.030 7.780 ;
        RECT 7.790 7.450 7.970 7.780 ;
        RECT 8.470 7.450 8.650 7.780 ;
        RECT 6.850 6.820 7.020 7.450 ;
        RECT 7.800 6.820 7.970 7.450 ;
        RECT 8.480 6.820 8.650 7.450 ;
        RECT 6.850 6.490 7.030 6.820 ;
        RECT 7.790 6.490 7.970 6.820 ;
        RECT 8.470 6.490 8.650 6.820 ;
        RECT 6.850 5.500 7.020 6.490 ;
        RECT 7.800 6.480 7.970 6.490 ;
        RECT 8.480 5.500 8.650 6.490 ;
        RECT 9.390 9.370 9.570 9.700 ;
        RECT 9.390 8.740 9.560 9.370 ;
        RECT 9.390 8.410 9.570 8.740 ;
        RECT 9.390 7.780 9.560 8.410 ;
        RECT 9.390 7.450 9.570 7.780 ;
        RECT 9.390 6.820 9.560 7.450 ;
        RECT 9.390 6.490 9.570 6.820 ;
        RECT 9.390 6.480 9.560 6.490 ;
        RECT 10.080 5.500 10.250 9.750 ;
        RECT 10.540 8.460 10.750 8.890 ;
        RECT 10.560 8.440 10.730 8.460 ;
        RECT 11.010 6.480 11.180 10.040 ;
        RECT 12.630 9.700 12.800 10.040 ;
        RECT 11.690 9.370 11.870 9.700 ;
        RECT 12.620 9.370 12.800 9.700 ;
        RECT 11.700 8.740 11.870 9.370 ;
        RECT 12.630 8.740 12.800 9.370 ;
        RECT 11.690 8.410 11.870 8.740 ;
        RECT 12.620 8.410 12.800 8.740 ;
        RECT 11.700 7.780 11.870 8.410 ;
        RECT 12.140 7.980 12.310 8.000 ;
        RECT 11.690 7.450 11.870 7.780 ;
        RECT 12.120 7.550 12.330 7.980 ;
        RECT 11.700 6.820 11.870 7.450 ;
        RECT 12.630 6.820 12.800 8.410 ;
        RECT 11.690 6.490 11.870 6.820 ;
        RECT 12.620 6.500 12.800 6.820 ;
        RECT 12.620 6.490 12.790 6.500 ;
        RECT 11.700 5.500 11.870 6.490 ;
        RECT 13.300 5.500 13.470 9.750 ;
        RECT 13.760 6.550 13.970 6.980 ;
        RECT 13.780 6.530 13.950 6.550 ;
        RECT 14.230 6.490 14.400 10.040 ;
        RECT 14.920 9.700 15.090 9.750 ;
        RECT 14.910 9.370 15.090 9.700 ;
        RECT 14.920 8.740 15.090 9.370 ;
        RECT 14.910 8.410 15.090 8.740 ;
        RECT 14.920 7.780 15.090 8.410 ;
        RECT 14.910 7.450 15.090 7.780 ;
        RECT 14.920 6.820 15.090 7.450 ;
        RECT 14.910 6.490 15.090 6.820 ;
        RECT 15.840 6.490 16.010 10.040 ;
        RECT 14.920 5.500 15.090 6.490 ;
        RECT 16.520 5.500 16.690 9.730 ;
        RECT 17.450 6.470 17.620 10.040 ;
        RECT 18.130 5.500 18.300 9.910 ;
        RECT 6.850 5.270 7.040 5.500 ;
        RECT 8.470 5.270 8.660 5.500 ;
        RECT 10.070 5.270 10.260 5.500 ;
        RECT 11.690 5.270 11.880 5.500 ;
        RECT 13.290 5.270 13.480 5.500 ;
        RECT 14.910 5.270 15.100 5.500 ;
        RECT 16.510 5.270 16.700 5.500 ;
        RECT 18.120 5.270 18.310 5.500 ;
        RECT 6.850 5.250 7.020 5.270 ;
        RECT 8.480 5.250 8.650 5.270 ;
        RECT 10.080 5.250 10.250 5.270 ;
        RECT 11.700 5.250 11.870 5.270 ;
        RECT 13.300 5.250 13.470 5.270 ;
        RECT 14.920 5.250 15.090 5.270 ;
        RECT 16.520 5.250 16.690 5.270 ;
        RECT 18.130 5.250 18.300 5.270 ;
      LAYER mcon ;
        RECT 16.720 10.820 16.890 10.990 ;
        RECT 17.390 10.820 17.560 10.990 ;
        RECT 12.140 7.830 12.310 8.000 ;
        RECT 6.860 5.300 7.030 5.470 ;
        RECT 8.480 5.300 8.650 5.470 ;
        RECT 10.080 5.300 10.250 5.470 ;
        RECT 11.700 5.300 11.870 5.470 ;
        RECT 13.300 5.300 13.470 5.470 ;
        RECT 14.920 5.300 15.090 5.470 ;
        RECT 16.520 5.300 16.690 5.470 ;
        RECT 18.130 5.300 18.300 5.470 ;
      LAYER met1 ;
        RECT 4.050 10.860 4.370 11.180 ;
        RECT 5.760 10.900 6.080 11.220 ;
        RECT 8.960 10.900 9.280 11.220 ;
        RECT 10.570 10.910 10.890 11.230 ;
        RECT 4.090 10.630 4.320 10.860 ;
        RECT 5.800 10.670 6.030 10.900 ;
        RECT 7.310 10.770 7.630 10.810 ;
        RECT 7.080 10.540 7.630 10.770 ;
        RECT 9.000 10.670 9.230 10.900 ;
        RECT 10.610 10.680 10.840 10.910 ;
        RECT 12.190 10.900 12.510 11.220 ;
        RECT 13.800 10.910 14.120 11.230 ;
        RECT 15.410 10.910 15.730 11.230 ;
        RECT 12.230 10.670 12.460 10.900 ;
        RECT 13.840 10.680 14.070 10.910 ;
        RECT 15.450 10.680 15.680 10.910 ;
        RECT 16.650 10.750 16.970 11.070 ;
        RECT 17.320 10.750 17.640 11.070 ;
        RECT 7.310 10.490 7.630 10.540 ;
        RECT 4.030 9.550 4.350 9.870 ;
        RECT 4.070 9.320 4.300 9.550 ;
        RECT 4.050 8.600 4.370 8.920 ;
        RECT 10.560 8.890 14.010 8.970 ;
        RECT 10.540 8.800 14.010 8.890 ;
        RECT 10.540 8.670 10.760 8.800 ;
        RECT 4.090 8.370 4.320 8.600 ;
        RECT 10.530 8.380 10.760 8.670 ;
        RECT 4.050 7.660 4.370 7.980 ;
        RECT 4.090 7.430 4.320 7.660 ;
        RECT 12.110 7.550 12.340 8.060 ;
        RECT 12.110 6.290 12.290 7.550 ;
        RECT 13.810 6.980 14.010 8.800 ;
        RECT 13.760 6.960 14.010 6.980 ;
        RECT 13.760 6.760 13.980 6.960 ;
        RECT 13.750 6.470 13.980 6.760 ;
        RECT 12.110 5.970 12.370 6.290 ;
      LAYER via ;
        RECT 4.080 10.890 4.340 11.150 ;
        RECT 5.790 10.930 6.050 11.190 ;
        RECT 8.990 10.930 9.250 11.190 ;
        RECT 10.600 10.940 10.860 11.200 ;
        RECT 12.220 10.930 12.480 11.190 ;
        RECT 7.340 10.520 7.600 10.780 ;
        RECT 13.830 10.940 14.090 11.200 ;
        RECT 15.440 10.940 15.700 11.200 ;
        RECT 16.680 10.780 16.940 11.040 ;
        RECT 17.350 10.780 17.610 11.040 ;
        RECT 4.060 9.580 4.320 9.840 ;
        RECT 4.080 8.630 4.340 8.890 ;
        RECT 4.080 7.690 4.340 7.950 ;
        RECT 12.110 6.000 12.370 6.260 ;
      LAYER met2 ;
        RECT 4.050 8.600 4.370 8.920 ;
        RECT 4.050 7.660 4.370 7.980 ;
  END
END sky130_hilas_DAC5bit01

MACRO sky130_hilas_capacitorSize04
  CLASS BLOCK ;
  FOREIGN sky130_hilas_capacitorSize04 ;
  ORIGIN -14.150 0.180 ;
  SIZE 5.780 BY 5.290 ;
  PIN CAP1TERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 19.110 3.650 19.770 4.310 ;
    END
  END CAP1TERM02
  PIN CAP2TERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 19.110 0.650 19.770 1.310 ;
    END
  END CAP2TERM02
  PIN CAP2TERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 14.270 1.050 14.930 1.310 ;
        RECT 16.710 1.050 17.160 1.060 ;
        RECT 14.270 0.650 17.210 1.050 ;
        RECT 14.720 0.640 17.210 0.650 ;
        RECT 16.690 0.560 17.210 0.640 ;
    END
  END CAP2TERM01
  PIN CAP1TERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 14.240 4.060 14.900 4.310 ;
        RECT 16.710 4.060 17.160 4.070 ;
        RECT 14.240 3.650 17.210 4.060 ;
        RECT 16.690 3.570 17.210 3.650 ;
    END
  END CAP1TERM01
  OBS
      LAYER met2 ;
        RECT 14.170 4.800 19.920 4.980 ;
        RECT 14.170 4.370 19.920 4.550 ;
        RECT 14.370 4.130 14.740 4.190 ;
        RECT 14.170 3.850 14.740 4.130 ;
        RECT 14.370 3.790 14.740 3.850 ;
        RECT 19.240 4.130 19.610 4.190 ;
        RECT 19.240 3.850 19.920 4.130 ;
        RECT 19.240 3.790 19.610 3.850 ;
        RECT 14.170 3.370 19.920 3.550 ;
        RECT 14.170 2.940 19.920 3.120 ;
        RECT 14.170 1.790 19.920 1.960 ;
        RECT 14.170 1.370 19.920 1.540 ;
        RECT 14.400 1.130 14.770 1.190 ;
        RECT 14.170 0.850 14.770 1.130 ;
        RECT 14.400 0.790 14.770 0.850 ;
        RECT 19.240 1.130 19.610 1.190 ;
        RECT 19.240 0.850 19.930 1.130 ;
        RECT 19.240 0.790 19.610 0.850 ;
        RECT 14.170 0.390 19.920 0.560 ;
        RECT 14.170 -0.050 19.920 0.120 ;
      LAYER via2 ;
        RECT 14.420 3.850 14.700 4.130 ;
        RECT 19.290 3.850 19.570 4.130 ;
        RECT 14.450 0.850 14.730 1.130 ;
        RECT 19.290 0.850 19.570 1.130 ;
      LAYER met3 ;
        RECT 15.860 4.340 18.160 5.110 ;
        RECT 14.150 3.590 14.940 4.340 ;
        RECT 15.860 3.590 19.810 4.340 ;
        RECT 15.860 2.830 18.160 3.590 ;
        RECT 14.180 0.590 14.970 1.340 ;
        RECT 15.860 1.330 18.160 2.100 ;
        RECT 19.020 1.330 19.810 1.340 ;
        RECT 15.860 0.600 19.810 1.330 ;
        RECT 15.860 -0.180 18.160 0.600 ;
        RECT 19.020 0.590 19.810 0.600 ;
      LAYER via3 ;
        RECT 14.340 3.740 14.770 4.220 ;
        RECT 19.210 3.740 19.640 4.220 ;
        RECT 14.370 0.740 14.800 1.220 ;
        RECT 19.210 0.740 19.640 1.220 ;
  END
END sky130_hilas_capacitorSize04

MACRO sky130_hilas_capacitorArray01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_capacitorArray01 ;
  ORIGIN 13.040 0.790 ;
  SIZE 36.700 BY 6.500 ;
  PIN CAPTERM2
    USE ANALOG ;
    PORT
      LAYER met3 ;
        RECT 22.190 1.630 23.340 3.270 ;
        RECT 22.640 1.620 23.340 1.630 ;
    END
  END CAPTERM2
  PIN CAPTERM1
    USE ANALOG ;
    ANTENNAGATEAREA 0.720000 ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met3 ;
        RECT -1.790 5.170 -1.410 5.460 ;
        RECT -1.870 3.920 -1.330 5.170 ;
    END
  END CAPTERM1
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -5.520 5.480 -2.960 5.710 ;
        RECT -5.520 -0.560 22.380 5.480 ;
        RECT -5.520 -0.790 -2.960 -0.560 ;
        RECT -1.040 -0.570 22.380 -0.560 ;
      LAYER met1 ;
        RECT -3.480 5.000 -3.320 5.700 ;
        RECT -3.590 4.450 -3.320 5.000 ;
        RECT -3.590 4.400 -3.310 4.450 ;
        RECT -3.480 4.310 -3.310 4.400 ;
        RECT -3.480 3.840 -3.320 4.310 ;
        RECT -3.480 3.750 -3.310 3.840 ;
        RECT -3.590 3.700 -3.310 3.750 ;
        RECT -3.590 3.150 -3.320 3.700 ;
        RECT -3.480 1.760 -3.320 3.150 ;
        RECT -3.590 1.210 -3.320 1.760 ;
        RECT -3.590 1.160 -3.310 1.210 ;
        RECT -3.480 1.070 -3.310 1.160 ;
        RECT -3.480 0.610 -3.320 1.070 ;
        RECT -3.480 0.520 -3.310 0.610 ;
        RECT -3.590 0.470 -3.310 0.520 ;
        RECT -3.590 -0.080 -3.320 0.470 ;
        RECT -3.480 -0.780 -3.320 -0.080 ;
    END
  END VINJ
  PIN GATESELECT
    ANTENNAGATEAREA 0.720000 ;
    ANTENNADIFFAREA 0.417600 ;
    PORT
      LAYER met2 ;
        RECT -2.300 5.450 -1.790 5.480 ;
        RECT -4.370 5.360 -4.050 5.430 ;
        RECT -2.300 5.360 -1.370 5.450 ;
        RECT -4.370 5.170 -1.370 5.360 ;
        RECT -1.870 5.150 -1.370 5.170 ;
      LAYER via2 ;
        RECT -1.740 5.150 -1.460 5.430 ;
    END
  END GATESELECT
  PIN VTUN
    ANTENNADIFFAREA 2.237600 ;
    PORT
      LAYER nwell ;
        RECT -13.030 3.120 -11.300 5.700 ;
        RECT -13.040 2.940 -11.300 3.120 ;
        RECT -13.030 -0.790 -11.300 2.940 ;
      LAYER met1 ;
        RECT -12.680 -0.790 -12.280 5.710 ;
    END
  END VTUN
  PIN GATE
    USE ANALOG ;
    ANTENNADIFFAREA 3.253900 ;
    PORT
      LAYER nwell ;
        RECT -9.280 -0.790 -7.050 5.700 ;
      LAYER met1 ;
        RECT -8.630 3.560 -8.250 5.710 ;
        RECT -8.640 1.700 -8.250 3.560 ;
        RECT -8.630 -0.420 -8.250 1.700 ;
        RECT -8.640 -0.570 -8.250 -0.420 ;
        RECT -8.630 -0.790 -8.250 -0.570 ;
    END
  END GATE
  PIN DRAIN2
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT -5.430 3.180 -5.120 3.190 ;
        RECT -13.030 3.120 -2.960 3.180 ;
        RECT 22.650 3.120 23.660 3.130 ;
        RECT -13.040 3.000 23.660 3.120 ;
        RECT -13.040 2.940 -12.920 3.000 ;
        RECT -5.430 2.860 -5.120 3.000 ;
        RECT -4.100 2.940 23.660 3.000 ;
    END
  END DRAIN2
  PIN DRAIN1
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT -5.430 5.150 -5.120 5.290 ;
        RECT -13.030 4.980 -2.960 5.150 ;
        RECT -13.030 4.970 23.660 4.980 ;
        RECT -13.030 4.800 -12.920 4.970 ;
        RECT -5.430 4.960 -5.120 4.970 ;
        RECT -4.060 4.800 23.660 4.970 ;
    END
  END DRAIN1
  PIN DRAIN4
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT -13.020 -0.050 -12.920 0.120 ;
        RECT -5.430 -0.050 -5.120 -0.040 ;
        RECT -4.230 -0.050 23.660 0.120 ;
        RECT -13.030 -0.220 -2.960 -0.050 ;
        RECT -5.430 -0.230 -2.960 -0.220 ;
        RECT -5.430 -0.370 -5.120 -0.230 ;
    END
  END DRAIN4
  PIN DRAIN3
    ANTENNADIFFAREA 0.115200 ;
    PORT
      LAYER met2 ;
        RECT -13.020 1.910 -12.920 1.960 ;
        RECT -5.430 1.910 -5.120 2.050 ;
        RECT -4.270 1.910 23.660 1.960 ;
        RECT -13.030 1.790 23.660 1.910 ;
        RECT -13.030 1.730 -2.960 1.790 ;
        RECT -5.430 1.720 -5.120 1.730 ;
    END
  END DRAIN3
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT -10.280 0.990 -9.960 1.000 ;
        RECT -6.350 0.990 -6.030 1.050 ;
        RECT -10.280 0.810 -6.030 0.990 ;
        RECT -10.280 0.740 -9.960 0.810 ;
        RECT -6.350 0.760 -6.030 0.810 ;
    END
    PORT
      LAYER met1 ;
        RECT -6.310 4.320 -6.070 5.710 ;
        RECT -6.330 3.660 -6.060 4.320 ;
        RECT -6.310 1.070 -6.070 3.660 ;
        RECT -6.320 0.750 -6.060 1.070 ;
        RECT -6.310 -0.790 -6.070 0.750 ;
      LAYER via ;
        RECT -6.320 0.780 -6.060 1.040 ;
    END
    PORT
      LAYER met1 ;
        RECT -10.240 4.300 -10.000 5.710 ;
        RECT -10.250 3.640 -9.990 4.300 ;
        RECT -10.240 1.030 -10.000 3.640 ;
        RECT -10.250 0.710 -9.990 1.030 ;
        RECT -10.240 -0.790 -10.000 0.710 ;
      LAYER via ;
        RECT -10.250 0.740 -9.990 1.000 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT -5.420 5.240 -5.100 5.250 ;
        RECT -5.420 5.070 -4.840 5.240 ;
        RECT -5.420 5.020 -5.090 5.070 ;
        RECT -5.420 4.990 -5.100 5.020 ;
        RECT -3.560 4.970 -3.360 5.320 ;
        RECT -5.420 4.660 -5.100 4.700 ;
        RECT -5.420 4.620 -5.090 4.660 ;
        RECT -5.420 4.450 -4.840 4.620 ;
        RECT -5.420 4.440 -5.100 4.450 ;
        RECT -4.290 4.350 -4.090 4.950 ;
        RECT -3.560 4.940 -3.350 4.970 ;
        RECT -3.570 4.350 -3.350 4.940 ;
        RECT -10.210 3.730 -10.040 4.260 ;
        RECT -6.270 3.720 -6.100 4.250 ;
        RECT -5.420 3.700 -5.100 3.710 ;
        RECT -5.420 3.530 -4.840 3.700 ;
        RECT -5.420 3.490 -5.090 3.530 ;
        RECT -5.420 3.450 -5.100 3.490 ;
        RECT -4.290 3.200 -4.090 3.800 ;
        RECT -3.570 3.210 -3.350 3.800 ;
        RECT -3.560 3.180 -3.350 3.210 ;
        RECT -5.420 3.130 -5.100 3.160 ;
        RECT -5.420 3.080 -5.090 3.130 ;
        RECT -12.610 2.230 -12.060 2.660 ;
        RECT -10.200 2.020 -10.030 3.030 ;
        RECT -5.420 2.910 -4.840 3.080 ;
        RECT -5.420 2.900 -5.100 2.910 ;
        RECT -8.580 2.160 -8.030 2.590 ;
        RECT -6.270 1.880 -6.100 2.890 ;
        RECT -3.560 2.830 -3.360 3.180 ;
        RECT -4.170 2.370 -3.730 2.540 ;
        RECT -5.420 2.000 -5.100 2.010 ;
        RECT -5.420 1.830 -4.840 2.000 ;
        RECT -5.420 1.780 -5.090 1.830 ;
        RECT -5.420 1.750 -5.100 1.780 ;
        RECT -3.560 1.730 -3.360 2.080 ;
        RECT -5.420 1.420 -5.100 1.460 ;
        RECT -5.420 1.380 -5.090 1.420 ;
        RECT -5.420 1.210 -4.840 1.380 ;
        RECT -5.420 1.200 -5.100 1.210 ;
        RECT -4.290 1.110 -4.090 1.710 ;
        RECT -3.560 1.700 -3.350 1.730 ;
        RECT -3.570 1.110 -3.350 1.700 ;
        RECT -5.420 0.470 -5.100 0.480 ;
        RECT -5.420 0.300 -4.840 0.470 ;
        RECT -5.420 0.260 -5.090 0.300 ;
        RECT -5.420 0.220 -5.100 0.260 ;
        RECT -4.290 -0.030 -4.090 0.570 ;
        RECT -3.570 -0.020 -3.350 0.570 ;
        RECT -3.560 -0.050 -3.350 -0.020 ;
        RECT -5.420 -0.100 -5.100 -0.070 ;
        RECT -5.420 -0.150 -5.090 -0.100 ;
        RECT -5.420 -0.320 -4.840 -0.150 ;
        RECT -5.420 -0.330 -5.100 -0.320 ;
        RECT -3.560 -0.400 -3.360 -0.050 ;
      LAYER mcon ;
        RECT -5.360 5.030 -5.190 5.200 ;
        RECT -4.280 4.740 -4.110 4.910 ;
        RECT -5.360 4.480 -5.190 4.650 ;
        RECT -3.550 4.770 -3.380 4.940 ;
        RECT -10.210 4.090 -10.040 4.260 ;
        RECT -6.270 4.080 -6.100 4.250 ;
        RECT -5.360 3.500 -5.190 3.670 ;
        RECT -4.280 3.240 -4.110 3.410 ;
        RECT -3.550 3.210 -3.380 3.380 ;
        RECT -5.360 2.950 -5.190 3.120 ;
        RECT -12.610 2.310 -12.340 2.580 ;
        RECT -10.200 2.630 -10.030 2.800 ;
        RECT -10.200 2.270 -10.030 2.440 ;
        RECT -8.580 2.240 -8.310 2.510 ;
        RECT -6.270 2.490 -6.100 2.660 ;
        RECT -3.910 2.370 -3.730 2.540 ;
        RECT -6.270 2.130 -6.100 2.300 ;
        RECT -5.360 1.790 -5.190 1.960 ;
        RECT -4.280 1.500 -4.110 1.670 ;
        RECT -5.360 1.240 -5.190 1.410 ;
        RECT -3.550 1.530 -3.380 1.700 ;
        RECT -5.360 0.270 -5.190 0.440 ;
        RECT -4.280 0.010 -4.110 0.180 ;
        RECT -3.550 -0.020 -3.380 0.150 ;
        RECT -5.360 -0.280 -5.190 -0.110 ;
      LAYER met1 ;
        RECT -4.290 5.460 -4.130 5.700 ;
        RECT -5.430 4.960 -5.110 5.280 ;
        RECT -4.340 5.140 -4.080 5.460 ;
        RECT -4.290 4.970 -4.130 5.140 ;
        RECT -4.290 4.950 -4.090 4.970 ;
        RECT -5.430 4.410 -5.110 4.730 ;
        RECT -4.310 4.710 -4.080 4.950 ;
        RECT -4.290 4.660 -4.080 4.710 ;
        RECT -3.920 4.660 -3.730 5.650 ;
        RECT -5.430 3.420 -5.110 3.740 ;
        RECT -4.290 3.490 -4.130 4.660 ;
        RECT -3.900 4.540 -3.730 4.660 ;
        RECT -3.890 3.610 -3.730 4.540 ;
        RECT -3.900 3.490 -3.730 3.610 ;
        RECT -4.290 3.440 -4.080 3.490 ;
        RECT -4.310 3.200 -4.080 3.440 ;
        RECT -5.430 2.870 -5.110 3.190 ;
        RECT -4.290 3.180 -4.090 3.200 ;
        RECT -4.290 2.550 -4.130 3.180 ;
        RECT -3.920 2.570 -3.730 3.490 ;
        RECT -3.940 2.550 -3.700 2.570 ;
        RECT -4.290 2.360 -3.700 2.550 ;
        RECT -5.430 1.720 -5.110 2.040 ;
        RECT -4.290 1.730 -4.130 2.360 ;
        RECT -3.940 2.340 -3.700 2.360 ;
        RECT -4.290 1.710 -4.090 1.730 ;
        RECT -5.430 1.170 -5.110 1.490 ;
        RECT -4.310 1.470 -4.080 1.710 ;
        RECT -4.290 1.420 -4.080 1.470 ;
        RECT -3.920 1.420 -3.730 2.340 ;
        RECT -5.430 0.190 -5.110 0.510 ;
        RECT -4.290 0.260 -4.130 1.420 ;
        RECT -3.900 1.300 -3.730 1.420 ;
        RECT -3.890 0.380 -3.730 1.300 ;
        RECT -3.900 0.260 -3.730 0.380 ;
        RECT -4.290 0.210 -4.080 0.260 ;
        RECT -4.310 -0.030 -4.080 0.210 ;
        RECT -5.430 -0.360 -5.110 -0.040 ;
        RECT -4.290 -0.050 -4.090 -0.030 ;
        RECT -4.290 -0.780 -4.130 -0.050 ;
        RECT -3.920 -0.730 -3.730 0.260 ;
      LAYER via ;
        RECT -5.400 4.990 -5.140 5.250 ;
        RECT -4.340 5.170 -4.080 5.430 ;
        RECT -5.400 4.440 -5.140 4.700 ;
        RECT -5.400 3.450 -5.140 3.710 ;
        RECT -5.400 2.900 -5.140 3.160 ;
        RECT -5.400 1.750 -5.140 2.010 ;
        RECT -5.400 1.200 -5.140 1.460 ;
        RECT -5.400 0.220 -5.140 0.480 ;
        RECT -5.400 -0.330 -5.140 -0.070 ;
      LAYER met2 ;
        RECT -5.430 4.720 -5.120 4.740 ;
        RECT -5.520 4.710 -2.960 4.720 ;
        RECT -13.030 4.550 -2.960 4.710 ;
        RECT -13.030 4.540 23.660 4.550 ;
        RECT -13.030 4.530 -5.120 4.540 ;
        RECT -5.430 4.410 -5.120 4.530 ;
        RECT -4.120 4.370 23.660 4.540 ;
        RECT -5.430 3.610 -5.120 3.740 ;
        RECT -3.160 3.610 -2.790 3.720 ;
        RECT -13.030 3.550 -2.790 3.610 ;
        RECT -13.030 3.430 23.660 3.550 ;
        RECT -5.430 3.410 -5.120 3.430 ;
        RECT -4.060 3.370 23.660 3.430 ;
        RECT -3.160 3.320 -2.790 3.370 ;
        RECT 22.970 2.220 23.660 2.630 ;
        RECT -3.200 1.540 -2.830 1.630 ;
        RECT -5.430 1.480 -5.120 1.500 ;
        RECT -4.170 1.480 23.660 1.540 ;
        RECT -13.030 1.370 23.660 1.480 ;
        RECT -13.030 1.300 -2.830 1.370 ;
        RECT -5.430 1.170 -5.120 1.300 ;
        RECT -3.200 1.230 -2.830 1.300 ;
        RECT -2.110 0.560 -1.740 0.760 ;
        RECT -5.430 0.380 -5.120 0.510 ;
        RECT -4.190 0.390 23.660 0.560 ;
        RECT -13.030 0.200 -2.960 0.380 ;
        RECT -2.110 0.360 -1.740 0.390 ;
        RECT -5.430 0.180 -5.120 0.200 ;
      LAYER via2 ;
        RECT -3.110 3.380 -2.830 3.660 ;
        RECT 23.040 2.280 23.330 2.560 ;
        RECT -3.150 1.290 -2.870 1.570 ;
        RECT -2.060 0.420 -1.780 0.700 ;
      LAYER met3 ;
        RECT -3.380 3.120 -2.590 3.870 ;
        RECT -3.420 1.730 -2.630 1.780 ;
        RECT -3.420 1.430 -2.490 1.730 ;
        RECT -3.420 1.030 -2.630 1.430 ;
        RECT -2.330 0.520 -1.540 0.910 ;
        RECT -2.330 0.220 -1.400 0.520 ;
        RECT -2.330 0.160 -1.540 0.220 ;
      LAYER via3 ;
        RECT -3.190 3.270 -2.760 3.750 ;
        RECT -3.230 1.180 -2.800 1.660 ;
        RECT -2.140 0.310 -1.710 0.790 ;
      LAYER met4 ;
        RECT -0.250 4.810 3.850 5.110 ;
        RECT -1.940 4.200 0.760 4.310 ;
        RECT -1.940 3.900 0.970 4.200 ;
        RECT -3.290 3.480 -2.630 3.840 ;
        RECT 0.460 3.560 0.970 3.900 ;
        RECT 3.470 3.610 3.850 4.810 ;
        RECT 6.310 3.640 9.590 3.940 ;
        RECT -3.290 3.180 -1.270 3.480 ;
        RECT -1.570 2.620 -1.270 3.180 ;
        RECT 6.310 2.620 6.610 3.640 ;
        RECT 9.290 2.620 9.590 3.640 ;
        RECT -1.570 2.320 9.590 2.620 ;
        RECT 11.990 3.620 20.880 3.920 ;
        RECT -3.330 1.730 -2.670 1.750 ;
        RECT 0.670 1.730 3.860 1.760 ;
        RECT 6.310 1.730 6.610 1.760 ;
        RECT -3.330 1.430 9.530 1.730 ;
        RECT -3.330 1.090 -2.670 1.430 ;
        RECT 0.670 1.060 0.970 1.430 ;
        RECT 3.560 1.090 3.860 1.430 ;
        RECT 6.310 1.090 6.610 1.430 ;
        RECT 3.560 1.060 6.610 1.090 ;
        RECT 9.230 1.060 9.530 1.430 ;
        RECT -2.240 0.520 -1.580 0.880 ;
        RECT 0.670 0.760 9.530 1.060 ;
        RECT 11.990 1.100 12.290 3.620 ;
        RECT 14.820 3.590 17.930 3.620 ;
        RECT 14.820 1.100 15.120 3.590 ;
        RECT 17.630 1.100 17.930 3.590 ;
        RECT 20.580 1.100 20.880 3.620 ;
        RECT 11.990 0.800 20.940 1.100 ;
        RECT 17.630 0.790 20.940 0.800 ;
        RECT -2.240 0.220 -1.190 0.520 ;
        RECT -1.490 -0.020 -1.190 0.220 ;
        RECT 20.640 -0.020 20.940 0.790 ;
        RECT -1.490 -0.320 20.940 -0.020 ;
  END
END sky130_hilas_capacitorArray01

MACRO sky130_hilas_pFETmed
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pFETmed ;
  ORIGIN -1.470 0.220 ;
  SIZE 1.190 BY 2.870 ;
  OBS
      LAYER nwell ;
        RECT 1.470 -0.220 2.660 2.650 ;
      LAYER li1 ;
        RECT 1.710 -0.070 1.880 2.420 ;
        RECT 2.260 -0.080 2.430 2.420 ;
  END
END sky130_hilas_pFETmed

MACRO sky130_hilas_swc4x1cellOverlap2
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc4x1cellOverlap2 ;
  ORIGIN 1.910 3.870 ;
  SIZE 9.350 BY 6.160 ;
  OBS
      LAYER nwell ;
        RECT 4.880 2.230 7.440 2.290 ;
        RECT 0.880 -3.820 7.440 2.230 ;
        RECT 4.880 -3.870 7.440 -3.820 ;
      LAYER li1 ;
        RECT -0.850 1.020 -0.680 1.910 ;
        RECT 1.230 0.920 4.540 1.900 ;
        RECT 4.980 1.820 5.300 1.830 ;
        RECT 4.980 1.650 5.560 1.820 ;
        RECT 4.980 1.600 5.310 1.650 ;
        RECT 4.980 1.570 5.300 1.600 ;
        RECT 6.840 1.550 7.040 1.900 ;
        RECT 4.980 1.240 5.300 1.280 ;
        RECT 4.980 1.200 5.310 1.240 ;
        RECT 4.980 1.030 5.560 1.200 ;
        RECT 4.980 1.020 5.300 1.030 ;
        RECT 6.110 0.930 6.310 1.530 ;
        RECT 6.840 1.520 7.050 1.550 ;
        RECT 6.830 0.930 7.050 1.520 ;
        RECT -0.850 -0.500 -0.680 0.390 ;
        RECT 1.230 -0.550 4.540 0.430 ;
        RECT 4.980 0.390 5.300 0.400 ;
        RECT 4.980 0.220 5.560 0.390 ;
        RECT 4.980 0.180 5.310 0.220 ;
        RECT 4.980 0.140 5.300 0.180 ;
        RECT 6.110 -0.110 6.310 0.490 ;
        RECT 6.830 -0.100 7.050 0.490 ;
        RECT 6.840 -0.130 7.050 -0.100 ;
        RECT 4.980 -0.180 5.300 -0.150 ;
        RECT 4.980 -0.230 5.310 -0.180 ;
        RECT 4.980 -0.400 5.560 -0.230 ;
        RECT 4.980 -0.410 5.300 -0.400 ;
        RECT 6.840 -0.480 7.040 -0.130 ;
        RECT 6.230 -0.880 6.670 -0.710 ;
        RECT -0.850 -1.950 -0.680 -1.060 ;
        RECT 1.230 -2.020 4.540 -1.040 ;
        RECT 4.980 -1.190 5.300 -1.180 ;
        RECT 4.980 -1.360 5.560 -1.190 ;
        RECT 4.980 -1.410 5.310 -1.360 ;
        RECT 4.980 -1.440 5.300 -1.410 ;
        RECT 6.840 -1.460 7.040 -1.110 ;
        RECT 4.980 -1.770 5.300 -1.730 ;
        RECT 4.980 -1.810 5.310 -1.770 ;
        RECT 4.980 -1.980 5.560 -1.810 ;
        RECT 4.980 -1.990 5.300 -1.980 ;
        RECT 6.110 -2.080 6.310 -1.480 ;
        RECT 6.840 -1.490 7.050 -1.460 ;
        RECT 6.830 -2.080 7.050 -1.490 ;
        RECT -0.850 -3.490 -0.680 -2.600 ;
        RECT 1.230 -3.490 4.540 -2.510 ;
        RECT 4.980 -2.610 5.300 -2.600 ;
        RECT 4.980 -2.780 5.560 -2.610 ;
        RECT 4.980 -2.820 5.310 -2.780 ;
        RECT 4.980 -2.860 5.300 -2.820 ;
        RECT 6.110 -3.110 6.310 -2.510 ;
        RECT 6.830 -3.100 7.050 -2.510 ;
        RECT 6.840 -3.130 7.050 -3.100 ;
        RECT 4.980 -3.180 5.300 -3.150 ;
        RECT 4.980 -3.230 5.310 -3.180 ;
        RECT 4.980 -3.400 5.560 -3.230 ;
        RECT 4.980 -3.410 5.300 -3.400 ;
        RECT 6.840 -3.480 7.040 -3.130 ;
      LAYER mcon ;
        RECT -0.850 1.710 -0.680 1.880 ;
        RECT 2.800 1.670 2.970 1.840 ;
        RECT 5.040 1.610 5.210 1.780 ;
        RECT 6.120 1.320 6.290 1.490 ;
        RECT 2.800 0.980 2.970 1.150 ;
        RECT 5.040 1.060 5.210 1.230 ;
        RECT 6.850 1.350 7.020 1.520 ;
        RECT -0.850 0.190 -0.680 0.360 ;
        RECT 2.800 0.200 2.970 0.370 ;
        RECT 5.040 0.190 5.210 0.360 ;
        RECT 6.120 -0.070 6.290 0.100 ;
        RECT 6.850 -0.100 7.020 0.070 ;
        RECT 2.800 -0.490 2.970 -0.320 ;
        RECT 5.040 -0.360 5.210 -0.190 ;
        RECT 6.490 -0.880 6.670 -0.710 ;
        RECT -0.850 -1.260 -0.680 -1.090 ;
        RECT 2.800 -1.270 2.970 -1.100 ;
        RECT 5.040 -1.400 5.210 -1.230 ;
        RECT 6.120 -1.690 6.290 -1.520 ;
        RECT 2.800 -1.960 2.970 -1.790 ;
        RECT 5.040 -1.950 5.210 -1.780 ;
        RECT 6.850 -1.660 7.020 -1.490 ;
        RECT -0.850 -2.800 -0.680 -2.630 ;
        RECT 2.800 -2.740 2.970 -2.570 ;
        RECT 5.040 -2.810 5.210 -2.640 ;
        RECT 6.120 -3.070 6.290 -2.900 ;
        RECT 6.850 -3.100 7.020 -2.930 ;
        RECT 2.800 -3.430 2.970 -3.260 ;
        RECT 5.040 -3.360 5.210 -3.190 ;
      LAYER met1 ;
        RECT -0.900 -3.820 -0.630 2.230 ;
        RECT 2.760 1.260 3.000 1.900 ;
        RECT 4.970 1.540 5.290 1.860 ;
        RECT 6.110 1.550 6.270 2.280 ;
        RECT 6.110 1.530 6.310 1.550 ;
        RECT 2.770 1.000 3.000 1.260 ;
        RECT 2.770 0.780 3.010 1.000 ;
        RECT 4.970 0.990 5.290 1.310 ;
        RECT 6.090 1.290 6.320 1.530 ;
        RECT 6.110 1.240 6.320 1.290 ;
        RECT 6.480 1.240 6.670 2.230 ;
        RECT 6.920 1.580 7.080 2.280 ;
        RECT 2.760 -0.210 3.000 0.430 ;
        RECT 4.970 0.110 5.290 0.430 ;
        RECT 6.110 0.180 6.270 1.240 ;
        RECT 6.500 1.120 6.670 1.240 ;
        RECT 6.510 0.300 6.670 1.120 ;
        RECT 6.810 1.030 7.080 1.580 ;
        RECT 6.810 0.980 7.090 1.030 ;
        RECT 6.920 0.890 7.090 0.980 ;
        RECT 6.920 0.530 7.080 0.890 ;
        RECT 6.920 0.440 7.090 0.530 ;
        RECT 6.500 0.180 6.670 0.300 ;
        RECT 6.110 0.130 6.320 0.180 ;
        RECT 6.090 -0.110 6.320 0.130 ;
        RECT 2.770 -0.470 3.000 -0.210 ;
        RECT 4.970 -0.440 5.290 -0.120 ;
        RECT 6.110 -0.130 6.310 -0.110 ;
        RECT 2.770 -0.690 3.010 -0.470 ;
        RECT 2.760 -1.680 3.000 -1.040 ;
        RECT 4.970 -1.470 5.290 -1.150 ;
        RECT 6.110 -1.460 6.270 -0.130 ;
        RECT 6.480 -0.680 6.670 0.180 ;
        RECT 6.810 0.390 7.090 0.440 ;
        RECT 6.810 -0.160 7.080 0.390 ;
        RECT 6.460 -0.910 6.700 -0.680 ;
        RECT 6.110 -1.480 6.310 -1.460 ;
        RECT 2.770 -1.940 3.000 -1.680 ;
        RECT 2.770 -2.160 3.010 -1.940 ;
        RECT 4.970 -2.020 5.290 -1.700 ;
        RECT 6.090 -1.720 6.320 -1.480 ;
        RECT 6.110 -1.770 6.320 -1.720 ;
        RECT 6.480 -1.770 6.670 -0.910 ;
        RECT 6.920 -1.430 7.080 -0.160 ;
        RECT 2.760 -3.150 3.000 -2.510 ;
        RECT 4.970 -2.890 5.290 -2.570 ;
        RECT 6.110 -2.820 6.270 -1.770 ;
        RECT 6.500 -1.890 6.670 -1.770 ;
        RECT 6.510 -2.700 6.670 -1.890 ;
        RECT 6.810 -1.980 7.080 -1.430 ;
        RECT 6.810 -2.030 7.090 -1.980 ;
        RECT 6.920 -2.120 7.090 -2.030 ;
        RECT 6.920 -2.470 7.080 -2.120 ;
        RECT 6.920 -2.560 7.090 -2.470 ;
        RECT 6.500 -2.820 6.670 -2.700 ;
        RECT 6.110 -2.870 6.320 -2.820 ;
        RECT 6.090 -3.110 6.320 -2.870 ;
        RECT 2.770 -3.410 3.000 -3.150 ;
        RECT 2.770 -3.630 3.010 -3.410 ;
        RECT 4.970 -3.440 5.290 -3.120 ;
        RECT 6.110 -3.130 6.310 -3.110 ;
        RECT 6.110 -3.860 6.270 -3.130 ;
        RECT 6.480 -3.810 6.670 -2.820 ;
        RECT 6.810 -2.610 7.090 -2.560 ;
        RECT 6.810 -3.160 7.080 -2.610 ;
        RECT 6.920 -3.860 7.080 -3.160 ;
      LAYER via ;
        RECT 5.000 1.570 5.260 1.830 ;
        RECT 5.000 1.020 5.260 1.280 ;
        RECT 5.000 0.140 5.260 0.400 ;
        RECT 5.000 -0.410 5.260 -0.150 ;
        RECT 5.000 -1.440 5.260 -1.180 ;
        RECT 5.000 -1.990 5.260 -1.730 ;
        RECT 5.000 -2.860 5.260 -2.600 ;
        RECT 5.000 -3.410 5.260 -3.150 ;
      LAYER met2 ;
        RECT 4.970 1.730 5.280 1.870 ;
        RECT -1.910 1.550 7.440 1.730 ;
        RECT 4.970 1.540 5.280 1.550 ;
        RECT 4.970 1.300 5.280 1.320 ;
        RECT -1.910 1.120 7.440 1.300 ;
        RECT 4.970 0.990 5.280 1.120 ;
        RECT 4.970 0.300 5.280 0.430 ;
        RECT -1.910 0.120 7.440 0.300 ;
        RECT 4.970 0.100 5.280 0.120 ;
        RECT 4.970 -0.130 5.280 -0.120 ;
        RECT -1.910 -0.200 4.960 -0.130 ;
        RECT 4.970 -0.200 7.440 -0.130 ;
        RECT -1.910 -0.310 7.440 -0.200 ;
        RECT 4.970 -0.450 5.280 -0.310 ;
        RECT 4.970 -1.280 5.280 -1.140 ;
        RECT 4.970 -1.290 7.440 -1.280 ;
        RECT -1.910 -1.460 7.440 -1.290 ;
        RECT 4.970 -1.470 5.280 -1.460 ;
        RECT 4.970 -1.710 5.280 -1.690 ;
        RECT -1.910 -1.880 7.440 -1.710 ;
        RECT 4.880 -1.890 7.440 -1.880 ;
        RECT 4.970 -2.020 5.280 -1.890 ;
        RECT 4.970 -2.690 5.280 -2.570 ;
        RECT -1.910 -2.700 5.280 -2.690 ;
        RECT -1.910 -2.860 7.440 -2.700 ;
        RECT 4.880 -2.880 7.440 -2.860 ;
        RECT 4.970 -2.900 5.280 -2.880 ;
        RECT 4.970 -3.130 5.280 -3.120 ;
        RECT -1.910 -3.300 7.440 -3.130 ;
        RECT 4.970 -3.310 7.440 -3.300 ;
        RECT 4.970 -3.450 5.280 -3.310 ;
  END
END sky130_hilas_swc4x1cellOverlap2

MACRO sky130_hilas_TA2SignalBiasCell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TA2SignalBiasCell ;
  ORIGIN 5.690 -1.400 ;
  SIZE 8.880 BY 6.050 ;
  PIN VOUT_AMP2
    USE ANALOG ;
    ANTENNADIFFAREA 0.308800 ;
    PORT
      LAYER met2 ;
        RECT 0.270 4.970 0.580 5.030 ;
        RECT 2.570 4.970 2.880 4.990 ;
        RECT 0.270 4.740 3.190 4.970 ;
        RECT 0.270 4.700 0.580 4.740 ;
        RECT 2.570 4.660 2.880 4.740 ;
    END
  END VOUT_AMP2
  PIN VOUT_AMP1
    USE ANALOG ;
    ANTENNADIFFAREA 0.308800 ;
    PORT
      LAYER met2 ;
        RECT 0.270 4.140 0.580 4.190 ;
        RECT 2.560 4.140 2.870 4.270 ;
        RECT 0.270 3.920 3.190 4.140 ;
        RECT 0.270 3.860 0.580 3.920 ;
    END
  END VOUT_AMP1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 1.230 1.400 1.570 7.450 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -5.690 7.440 -1.650 7.450 ;
        RECT -5.690 1.410 -0.090 7.440 ;
        RECT -1.950 1.400 -0.090 1.410 ;
        RECT 1.910 1.400 3.190 7.450 ;
      LAYER met2 ;
        RECT -4.900 7.270 -4.660 7.450 ;
        RECT -4.940 6.980 -4.630 7.270 ;
        RECT -5.420 6.940 -4.630 6.980 ;
        RECT -5.420 6.630 -4.660 6.940 ;
        RECT -5.420 6.400 -0.880 6.630 ;
        RECT -5.420 6.160 -4.660 6.400 ;
        RECT -5.420 6.150 -4.970 6.160 ;
        RECT -1.110 6.040 -0.880 6.400 ;
        RECT 1.910 6.040 2.240 6.190 ;
        RECT -1.110 5.840 2.240 6.040 ;
        RECT -0.850 5.830 2.240 5.840 ;
        RECT 1.910 5.260 2.240 5.830 ;
        RECT -4.980 2.780 -4.670 3.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.900 6.190 2.170 7.450 ;
        RECT 1.900 5.260 2.250 6.190 ;
        RECT 1.900 3.280 2.170 5.260 ;
        RECT 1.900 2.990 2.180 3.280 ;
        RECT 1.900 1.400 2.170 2.990 ;
      LAYER via ;
        RECT 1.940 5.290 2.200 6.150 ;
    END
  END VPWR
  PIN VIN22
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -1.300 7.430 -1.050 7.440 ;
        RECT -0.700 7.430 -0.390 7.440 ;
        RECT -1.300 7.180 -0.390 7.430 ;
        RECT -0.700 7.110 -0.390 7.180 ;
    END
  END VIN22
  PIN VIN21
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -0.940 4.750 -0.630 4.790 ;
        RECT -1.030 4.740 -0.600 4.750 ;
        RECT -1.260 4.510 -0.160 4.740 ;
        RECT -0.940 4.460 -0.630 4.510 ;
    END
  END VIN21
  PIN VIN11
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -2.500 4.340 -2.190 4.390 ;
        RECT -2.820 4.110 -1.720 4.340 ;
        RECT -2.820 4.100 -2.160 4.110 ;
        RECT -2.500 4.060 -2.190 4.100 ;
    END
  END VIN11
  PIN VIN12
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -2.260 1.670 -1.950 1.740 ;
        RECT -2.860 1.420 -1.950 1.670 ;
        RECT -2.260 1.410 -1.950 1.420 ;
    END
  END VIN12
  PIN VBIAS2
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -4.010 1.670 -3.700 1.740 ;
        RECT -4.580 1.660 -3.700 1.670 ;
        RECT -5.640 1.430 -3.700 1.660 ;
        RECT -4.580 1.420 -3.700 1.430 ;
        RECT -4.010 1.410 -3.700 1.420 ;
    END
  END VBIAS2
  PIN VBIAS1
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -4.250 4.340 -3.940 4.390 ;
        RECT -5.680 4.110 -3.470 4.340 ;
        RECT -5.680 4.100 -3.910 4.110 ;
        RECT -5.680 4.090 -5.040 4.100 ;
        RECT -4.250 4.060 -3.940 4.100 ;
    END
  END VBIAS1
  OBS
      LAYER li1 ;
        RECT -0.960 7.400 -0.790 7.450 ;
        RECT -4.930 7.190 -4.610 7.230 ;
        RECT -4.930 7.000 -4.600 7.190 ;
        RECT -0.960 7.140 -0.400 7.400 ;
        RECT 0.510 7.150 0.710 7.190 ;
        RECT -0.960 7.120 -0.790 7.140 ;
        RECT -4.930 6.980 -4.610 7.000 ;
        RECT -5.020 6.970 -4.610 6.980 ;
        RECT -5.270 6.780 -4.670 6.970 ;
        RECT -5.440 6.240 -4.670 6.780 ;
        RECT -5.440 4.910 -5.270 6.240 ;
        RECT -5.430 1.970 -5.260 3.750 ;
        RECT -4.850 3.070 -4.670 6.240 ;
        RECT -4.040 5.950 -3.870 6.970 ;
        RECT -4.090 5.910 -3.770 5.950 ;
        RECT -4.090 5.720 -3.760 5.910 ;
        RECT -4.090 5.690 -3.770 5.720 ;
        RECT -4.040 5.190 -3.870 5.690 ;
        RECT -4.120 5.130 -3.580 5.190 ;
        RECT -4.120 5.020 -3.570 5.130 ;
        RECT -3.760 4.900 -3.570 5.020 ;
        RECT -4.290 4.600 -4.120 4.760 ;
        RECT -4.290 4.430 -4.070 4.600 ;
        RECT -4.240 4.350 -4.070 4.430 ;
        RECT -4.240 4.310 -3.920 4.350 ;
        RECT -4.240 4.120 -3.910 4.310 ;
        RECT -4.240 4.090 -3.920 4.120 ;
        RECT -4.970 3.030 -4.650 3.070 ;
        RECT -4.970 2.840 -4.640 3.030 ;
        RECT -4.970 2.810 -4.650 2.840 ;
        RECT -4.850 1.880 -4.670 2.810 ;
        RECT -4.040 2.540 -3.870 3.920 ;
        RECT -3.100 3.070 -2.920 6.980 ;
        RECT -2.290 5.190 -2.120 6.970 ;
        RECT -1.540 6.040 -1.360 6.970 ;
        RECT 0.280 6.890 0.710 7.150 ;
        RECT -0.810 6.710 -0.480 6.880 ;
        RECT 0.510 6.860 0.710 6.890 ;
        RECT -0.730 6.570 -0.480 6.710 ;
        RECT -0.730 6.310 -0.250 6.570 ;
        RECT 0.100 6.500 0.270 6.540 ;
        RECT 0.510 6.500 0.710 6.530 ;
        RECT -1.660 6.010 -1.340 6.040 ;
        RECT -1.660 5.820 -1.330 6.010 ;
        RECT -1.660 5.780 -1.340 5.820 ;
        RECT -2.370 5.130 -1.830 5.190 ;
        RECT -2.370 5.020 -1.820 5.130 ;
        RECT -2.010 4.900 -1.820 5.020 ;
        RECT -2.540 4.600 -2.370 4.760 ;
        RECT -2.540 4.430 -2.320 4.600 ;
        RECT -2.490 4.350 -2.320 4.430 ;
        RECT -2.490 4.310 -2.170 4.350 ;
        RECT -2.490 4.120 -2.160 4.310 ;
        RECT -2.490 4.090 -2.170 4.120 ;
        RECT -3.220 3.030 -2.900 3.070 ;
        RECT -3.220 2.840 -2.890 3.030 ;
        RECT -3.220 2.810 -2.900 2.840 ;
        RECT -4.040 2.280 -3.560 2.540 ;
        RECT -4.040 2.140 -3.790 2.280 ;
        RECT -4.120 1.970 -3.790 2.140 ;
        RECT -3.100 1.880 -2.920 2.810 ;
        RECT -2.290 2.540 -2.120 3.920 ;
        RECT -2.290 2.280 -1.810 2.540 ;
        RECT -2.290 2.140 -2.040 2.280 ;
        RECT -2.370 1.970 -2.040 2.140 ;
        RECT -1.540 1.870 -1.360 5.780 ;
        RECT -0.730 4.930 -0.560 6.310 ;
        RECT 0.100 6.240 0.710 6.500 ;
        RECT 0.100 6.210 0.270 6.240 ;
        RECT 0.510 6.200 0.710 6.240 ;
        RECT 1.100 6.200 1.650 7.190 ;
        RECT 2.470 7.040 3.100 7.210 ;
        RECT 2.470 6.940 2.860 7.040 ;
        RECT 2.470 6.910 2.850 6.940 ;
        RECT 2.470 6.760 2.830 6.910 ;
        RECT 2.120 6.590 2.830 6.760 ;
        RECT 0.100 5.650 0.270 5.680 ;
        RECT 0.510 5.650 0.710 5.690 ;
        RECT 0.100 5.390 0.710 5.650 ;
        RECT 0.100 5.350 0.270 5.390 ;
        RECT 0.510 5.360 0.710 5.390 ;
        RECT 0.510 5.000 0.710 5.030 ;
        RECT -0.930 4.730 -0.610 4.760 ;
        RECT 0.280 4.740 0.710 5.000 ;
        RECT -0.930 4.540 -0.600 4.730 ;
        RECT 0.510 4.700 0.710 4.740 ;
        RECT 1.100 4.700 1.650 5.690 ;
        RECT 1.960 5.270 2.820 6.150 ;
        RECT 1.960 5.260 2.170 5.270 ;
        RECT 2.580 4.910 2.900 4.950 ;
        RECT 2.580 4.850 2.910 4.910 ;
        RECT 2.110 4.720 2.910 4.850 ;
        RECT 2.110 4.690 2.900 4.720 ;
        RECT 2.110 4.670 2.810 4.690 ;
        RECT -0.930 4.500 -0.610 4.540 ;
        RECT -0.930 4.420 -0.760 4.500 ;
        RECT -0.980 4.250 -0.760 4.420 ;
        RECT -0.980 4.090 -0.810 4.250 ;
        RECT 2.570 4.190 2.890 4.230 ;
        RECT 0.510 4.150 0.710 4.190 ;
        RECT -0.450 3.830 -0.260 3.950 ;
        RECT 0.280 3.890 0.710 4.150 ;
        RECT 0.510 3.860 0.710 3.890 ;
        RECT -0.810 3.720 -0.260 3.830 ;
        RECT -0.810 3.660 -0.270 3.720 ;
        RECT -0.730 1.880 -0.560 3.660 ;
        RECT 0.100 3.500 0.270 3.540 ;
        RECT 0.510 3.500 0.710 3.530 ;
        RECT 0.100 3.240 0.710 3.500 ;
        RECT 0.100 3.210 0.270 3.240 ;
        RECT 0.510 3.200 0.710 3.240 ;
        RECT 1.100 3.200 1.650 4.190 ;
        RECT 2.110 4.010 2.900 4.190 ;
        RECT 2.570 4.000 2.900 4.010 ;
        RECT 2.570 3.970 2.890 4.000 ;
        RECT 2.120 3.250 2.820 3.590 ;
        RECT 1.970 3.020 2.820 3.250 ;
        RECT 2.120 2.710 2.820 3.020 ;
        RECT 0.100 2.650 0.270 2.680 ;
        RECT 0.510 2.650 0.710 2.690 ;
        RECT 0.100 2.390 0.710 2.650 ;
        RECT 0.100 2.350 0.270 2.390 ;
        RECT 0.510 2.360 0.710 2.390 ;
        RECT 0.510 2.000 0.710 2.030 ;
        RECT 0.280 1.740 0.710 2.000 ;
        RECT -4.270 1.710 -4.100 1.730 ;
        RECT -2.520 1.710 -2.350 1.730 ;
        RECT -4.270 1.450 -3.710 1.710 ;
        RECT -2.520 1.450 -1.960 1.710 ;
        RECT 0.510 1.700 0.710 1.740 ;
        RECT 1.100 1.700 1.650 2.690 ;
        RECT 2.120 2.100 2.830 2.270 ;
        RECT 2.470 1.820 2.830 2.100 ;
        RECT 2.470 1.650 3.100 1.820 ;
        RECT -4.270 1.400 -4.100 1.450 ;
        RECT -2.520 1.400 -2.350 1.450 ;
      LAYER mcon ;
        RECT -4.870 7.010 -4.700 7.180 ;
        RECT -0.630 7.180 -0.460 7.350 ;
        RECT -5.440 6.610 -5.270 6.780 ;
        RECT -4.850 6.560 -4.680 6.730 ;
        RECT -5.440 6.270 -5.270 6.440 ;
        RECT -5.440 5.930 -5.270 6.100 ;
        RECT -5.440 5.590 -5.270 5.760 ;
        RECT -5.440 5.250 -5.270 5.420 ;
        RECT -4.850 6.220 -4.680 6.390 ;
        RECT -5.430 3.580 -5.260 3.750 ;
        RECT -5.430 3.240 -5.260 3.410 ;
        RECT -4.030 5.730 -3.860 5.900 ;
        RECT -3.750 4.930 -3.580 5.100 ;
        RECT -4.180 4.130 -4.010 4.300 ;
        RECT -5.430 2.900 -5.260 3.070 ;
        RECT -4.910 2.850 -4.740 3.020 ;
        RECT -5.430 2.560 -5.260 2.730 ;
        RECT -5.430 2.220 -5.260 2.390 ;
        RECT 0.340 6.930 0.510 7.100 ;
        RECT 1.320 6.610 1.490 6.780 ;
        RECT 2.590 6.950 2.760 7.120 ;
        RECT -0.480 6.350 -0.310 6.520 ;
        RECT -1.600 5.830 -1.430 6.000 ;
        RECT -2.000 4.930 -1.830 5.100 ;
        RECT -2.430 4.130 -2.260 4.300 ;
        RECT -3.160 2.850 -2.990 3.020 ;
        RECT -3.790 2.330 -3.620 2.500 ;
        RECT -2.040 2.330 -1.870 2.500 ;
        RECT 0.290 6.280 0.460 6.450 ;
        RECT 1.980 5.980 2.150 6.150 ;
        RECT 0.290 5.440 0.460 5.610 ;
        RECT 1.320 5.110 1.490 5.280 ;
        RECT 1.980 5.640 2.150 5.810 ;
        RECT 1.980 5.280 2.150 5.450 ;
        RECT 0.340 4.790 0.510 4.960 ;
        RECT -0.870 4.550 -0.700 4.720 ;
        RECT 2.640 4.730 2.810 4.900 ;
        RECT -0.440 3.750 -0.270 3.920 ;
        RECT 0.340 3.930 0.510 4.100 ;
        RECT 2.630 4.010 2.800 4.180 ;
        RECT 1.320 3.610 1.490 3.780 ;
        RECT 0.290 3.280 0.460 3.450 ;
        RECT 1.980 3.050 2.150 3.220 ;
        RECT 0.290 2.440 0.460 2.610 ;
        RECT 1.320 2.110 1.490 2.280 ;
        RECT 0.340 1.790 0.510 1.960 ;
        RECT -3.940 1.500 -3.770 1.670 ;
        RECT 2.550 1.760 2.720 1.930 ;
        RECT -2.190 1.500 -2.020 1.670 ;
      LAYER met1 ;
        RECT -4.940 6.990 -4.620 7.260 ;
        RECT -0.710 7.110 -0.390 7.430 ;
        RECT -5.470 6.940 -4.620 6.990 ;
        RECT -5.470 6.670 -4.650 6.940 ;
        RECT 0.270 6.860 0.590 7.180 ;
        RECT 2.520 6.880 2.840 7.200 ;
        RECT -5.470 6.380 -4.620 6.670 ;
        RECT -5.470 6.130 -4.650 6.380 ;
        RECT -0.560 6.280 -0.240 6.600 ;
        RECT 0.220 6.210 0.540 6.530 ;
        RECT -5.470 3.100 -4.830 6.130 ;
        RECT -4.100 5.660 -3.780 5.980 ;
        RECT -1.670 5.750 -1.350 6.070 ;
        RECT -0.450 5.590 -0.240 5.700 ;
        RECT -0.470 5.270 -0.210 5.590 ;
        RECT 0.220 5.360 0.540 5.680 ;
        RECT -3.780 4.870 -3.550 5.160 ;
        RECT -2.030 4.870 -1.800 5.160 ;
        RECT -4.250 4.060 -3.930 4.380 ;
        RECT -3.760 3.580 -3.550 4.870 ;
        RECT -2.500 4.060 -2.180 4.380 ;
        RECT -2.010 3.580 -1.800 4.870 ;
        RECT -0.940 4.470 -0.620 4.790 ;
        RECT -0.450 3.980 -0.240 5.270 ;
        RECT 0.270 4.710 0.590 5.030 ;
        RECT 2.570 4.660 2.890 4.980 ;
        RECT -0.470 3.690 -0.240 3.980 ;
        RECT 0.270 3.860 0.590 4.180 ;
        RECT 2.560 3.940 2.880 4.260 ;
        RECT -3.780 3.260 -3.520 3.580 ;
        RECT -2.030 3.260 -1.770 3.580 ;
        RECT -3.760 3.150 -3.550 3.260 ;
        RECT -2.010 3.150 -1.800 3.260 ;
        RECT 0.220 3.210 0.540 3.530 ;
        RECT -5.470 2.780 -4.660 3.100 ;
        RECT -3.230 2.780 -2.910 3.100 ;
        RECT -5.470 1.950 -4.830 2.780 ;
        RECT -3.870 2.250 -3.550 2.570 ;
        RECT -2.120 2.250 -1.800 2.570 ;
        RECT 0.220 2.360 0.540 2.680 ;
        RECT -5.250 1.940 -4.830 1.950 ;
        RECT -4.020 1.420 -3.700 1.740 ;
        RECT -2.270 1.420 -1.950 1.740 ;
        RECT 0.270 1.710 0.590 2.030 ;
        RECT 2.480 1.690 2.800 2.010 ;
      LAYER via ;
        RECT -4.910 6.970 -4.650 7.230 ;
        RECT -0.680 7.140 -0.420 7.400 ;
        RECT -5.350 6.190 -4.760 6.910 ;
        RECT 0.300 6.890 0.560 7.150 ;
        RECT 2.550 6.910 2.810 7.170 ;
        RECT -0.530 6.310 -0.270 6.570 ;
        RECT 0.250 6.240 0.510 6.500 ;
        RECT -4.070 5.690 -3.810 5.950 ;
        RECT -1.640 5.780 -1.380 6.040 ;
        RECT -0.470 5.300 -0.210 5.560 ;
        RECT 0.250 5.390 0.510 5.650 ;
        RECT -4.220 4.090 -3.960 4.350 ;
        RECT -2.470 4.090 -2.210 4.350 ;
        RECT -0.910 4.500 -0.650 4.760 ;
        RECT 0.300 4.740 0.560 5.000 ;
        RECT 2.600 4.690 2.860 4.950 ;
        RECT 0.300 3.890 0.560 4.150 ;
        RECT 2.590 3.970 2.850 4.230 ;
        RECT -3.780 3.290 -3.520 3.550 ;
        RECT -2.030 3.290 -1.770 3.550 ;
        RECT 0.250 3.240 0.510 3.500 ;
        RECT -4.950 2.810 -4.690 3.070 ;
        RECT -3.200 2.810 -2.940 3.070 ;
        RECT -3.840 2.280 -3.580 2.540 ;
        RECT -2.090 2.280 -1.830 2.540 ;
        RECT 0.250 2.390 0.510 2.650 ;
        RECT 0.300 1.740 0.560 2.000 ;
        RECT -3.990 1.450 -3.730 1.710 ;
        RECT 2.510 1.720 2.770 1.980 ;
        RECT -2.240 1.450 -1.980 1.710 ;
      LAYER met2 ;
        RECT 0.270 7.110 0.580 7.190 ;
        RECT 2.520 7.110 2.830 7.210 ;
        RECT 0.270 6.880 2.830 7.110 ;
        RECT 0.270 6.860 0.580 6.880 ;
        RECT -0.550 6.570 -0.240 6.610 ;
        RECT -0.730 6.460 0.010 6.570 ;
        RECT 0.220 6.460 0.530 6.540 ;
        RECT -0.730 6.320 0.530 6.460 ;
        RECT -0.550 6.280 0.530 6.320 ;
        RECT -0.240 6.250 0.530 6.280 ;
        RECT -0.240 6.200 0.010 6.250 ;
        RECT 0.220 6.210 0.530 6.250 ;
        RECT -4.100 5.930 -3.790 5.990 ;
        RECT -1.670 5.930 -1.360 6.070 ;
        RECT -4.100 5.740 -1.360 5.930 ;
        RECT -4.100 5.710 -1.620 5.740 ;
        RECT -4.100 5.660 -3.790 5.710 ;
        RECT 0.220 5.640 0.530 5.680 ;
        RECT -0.210 5.560 0.530 5.640 ;
        RECT -0.500 5.540 0.530 5.560 ;
        RECT -0.550 5.430 0.530 5.540 ;
        RECT -0.550 5.350 0.000 5.430 ;
        RECT 0.220 5.350 0.530 5.430 ;
        RECT -0.550 5.290 -0.080 5.350 ;
        RECT -3.860 3.310 -3.390 3.560 ;
        RECT -2.110 3.470 -1.640 3.560 ;
        RECT -2.110 3.460 0.000 3.470 ;
        RECT 0.220 3.460 0.530 3.540 ;
        RECT -2.110 3.310 0.530 3.460 ;
        RECT -3.810 3.290 -3.490 3.310 ;
        RECT -2.060 3.290 0.530 3.310 ;
        RECT -1.770 3.270 0.530 3.290 ;
        RECT -0.080 3.250 0.530 3.270 ;
        RECT 0.220 3.210 0.530 3.250 ;
        RECT -3.230 3.100 -2.920 3.110 ;
        RECT -3.340 2.920 -2.920 3.100 ;
        RECT -3.360 2.910 -2.920 2.920 ;
        RECT -3.580 2.780 -2.920 2.910 ;
        RECT -3.580 2.570 -3.220 2.780 ;
        RECT -2.060 2.640 0.000 2.670 ;
        RECT 0.220 2.640 0.530 2.680 ;
        RECT -2.060 2.570 0.530 2.640 ;
        RECT -3.860 2.530 -3.220 2.570 ;
        RECT -2.110 2.530 0.530 2.570 ;
        RECT -4.040 2.290 -3.220 2.530 ;
        RECT -2.290 2.460 0.530 2.530 ;
        RECT -4.040 2.280 -3.490 2.290 ;
        RECT -2.290 2.280 -1.740 2.460 ;
        RECT -0.080 2.430 0.530 2.460 ;
        RECT 0.220 2.350 0.530 2.430 ;
        RECT -3.860 2.240 -3.550 2.280 ;
        RECT -2.110 2.240 -1.800 2.280 ;
        RECT 0.270 1.980 0.580 2.030 ;
        RECT 2.480 1.980 2.790 2.020 ;
        RECT 0.270 1.750 2.980 1.980 ;
        RECT 0.270 1.700 0.580 1.750 ;
        RECT 2.480 1.690 2.790 1.750 ;
  END
END sky130_hilas_TA2SignalBiasCell

MACRO sky130_hilas_Tgate4Single01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_Tgate4Single01 ;
  ORIGIN 0.360 1.640 ;
  SIZE 4.760 BY 6.410 ;
  PIN VPWR
    USE ANALOG ;
    ANTENNADIFFAREA 0.966800 ;
    PORT
      LAYER nwell ;
        RECT -0.240 -1.640 2.520 4.770 ;
      LAYER met1 ;
        RECT 0.380 3.850 0.580 4.770 ;
        RECT 0.370 3.560 0.600 3.850 ;
        RECT 0.380 2.770 0.580 3.560 ;
        RECT 0.370 2.480 0.600 2.770 ;
        RECT 0.380 0.650 0.580 2.480 ;
        RECT 0.370 0.360 0.600 0.650 ;
        RECT 0.380 -0.430 0.580 0.360 ;
        RECT 0.370 -0.720 0.600 -0.430 ;
        RECT 0.380 -1.640 0.580 -0.720 ;
    END
  END VPWR
  PIN INPUT1_2
    USE ANALOG ;
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT 1.280 1.930 1.590 2.050 ;
        RECT 0.510 1.920 1.630 1.930 ;
        RECT 2.850 1.920 3.160 2.050 ;
        RECT -0.360 1.720 3.160 1.920 ;
        RECT 0.510 1.710 1.630 1.720 ;
    END
  END INPUT1_2
  PIN SELECT2
    USE ANALOG ;
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT -0.070 2.900 0.250 2.990 ;
        RECT -0.360 2.700 0.250 2.900 ;
    END
  END SELECT2
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 3.890 3.850 4.080 4.770 ;
        RECT 3.870 3.560 4.100 3.850 ;
        RECT 3.890 2.770 4.080 3.560 ;
        RECT 3.870 2.480 4.100 2.770 ;
        RECT 3.890 0.650 4.080 2.480 ;
        RECT 3.870 0.360 4.100 0.650 ;
        RECT 3.890 -0.430 4.080 0.360 ;
        RECT 3.870 -0.720 4.100 -0.430 ;
        RECT 3.890 -1.640 4.080 -0.720 ;
    END
  END VGND
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.212400 ;
    PORT
      LAYER met2 ;
        RECT 2.200 2.900 2.520 2.920 ;
        RECT 3.210 2.900 3.530 2.930 ;
        RECT 2.150 2.700 4.400 2.900 ;
        RECT 2.200 2.660 2.520 2.700 ;
        RECT 3.210 2.670 3.530 2.700 ;
    END
  END OUTPUT2
  PIN OUTPUT4
    ANTENNADIFFAREA 0.212400 ;
    PORT
      LAYER met2 ;
        RECT 2.200 -0.300 2.520 -0.280 ;
        RECT 3.210 -0.300 3.530 -0.270 ;
        RECT 2.150 -0.500 4.400 -0.300 ;
        RECT 2.200 -0.540 2.520 -0.500 ;
        RECT 3.210 -0.530 3.530 -0.500 ;
    END
  END OUTPUT4
  PIN OUTPUT3
    ANTENNADIFFAREA 0.212400 ;
    PORT
      LAYER met2 ;
        RECT 2.200 0.430 2.520 0.470 ;
        RECT 3.210 0.430 3.530 0.460 ;
        RECT 2.150 0.230 4.400 0.430 ;
        RECT 2.200 0.210 2.520 0.230 ;
        RECT 3.210 0.200 3.530 0.230 ;
    END
  END OUTPUT3
  PIN OUTPUT1
    ANTENNADIFFAREA 0.212400 ;
    PORT
      LAYER met2 ;
        RECT 2.200 3.630 2.520 3.670 ;
        RECT 3.210 3.630 3.530 3.660 ;
        RECT 2.150 3.430 4.400 3.630 ;
        RECT 2.200 3.410 2.520 3.430 ;
        RECT 3.210 3.400 3.530 3.430 ;
    END
  END OUTPUT1
  PIN INPUT1_4
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT 1.280 -1.270 1.590 -1.150 ;
        RECT 0.510 -1.280 1.630 -1.270 ;
        RECT 2.850 -1.280 3.160 -1.150 ;
        RECT -0.360 -1.480 3.160 -1.280 ;
        RECT 0.510 -1.490 1.630 -1.480 ;
    END
  END INPUT1_4
  PIN SELECT4
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT -0.070 -0.300 0.250 -0.210 ;
        RECT -0.360 -0.500 0.250 -0.300 ;
    END
  END SELECT4
  PIN SELECT3
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT -0.360 0.230 0.250 0.430 ;
        RECT -0.070 0.140 0.250 0.230 ;
    END
  END SELECT3
  PIN INPUT1_3
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT 0.510 1.410 1.630 1.420 ;
        RECT -0.360 1.210 3.160 1.410 ;
        RECT 0.510 1.200 1.630 1.210 ;
        RECT 1.280 1.080 1.590 1.200 ;
        RECT 2.850 1.080 3.160 1.210 ;
    END
  END INPUT1_3
  PIN SELECT1
    ANTENNAGATEAREA 0.432000 ;
    PORT
      LAYER met2 ;
        RECT -0.360 3.430 0.250 3.630 ;
        RECT -0.070 3.340 0.250 3.430 ;
    END
  END SELECT1
  PIN INPUT1_1
    ANTENNADIFFAREA 0.208800 ;
    PORT
      LAYER met2 ;
        RECT 0.510 4.610 1.630 4.620 ;
        RECT -0.360 4.410 3.160 4.610 ;
        RECT 0.510 4.400 1.630 4.410 ;
        RECT 1.280 4.280 1.590 4.400 ;
        RECT 2.850 4.280 3.160 4.410 ;
    END
  END INPUT1_1
  OBS
      LAYER li1 ;
        RECT 1.290 4.550 1.610 4.580 ;
        RECT 2.860 4.550 3.180 4.580 ;
        RECT 0.070 4.210 0.240 4.490 ;
        RECT 1.290 4.360 1.620 4.550 ;
        RECT 2.300 4.410 2.490 4.430 ;
        RECT 1.290 4.320 1.610 4.360 ;
        RECT 0.070 4.170 0.280 4.210 ;
        RECT 0.070 4.150 0.300 4.170 ;
        RECT 1.420 4.160 1.590 4.320 ;
        RECT 2.030 4.240 2.490 4.410 ;
        RECT 2.860 4.360 3.190 4.550 ;
        RECT 3.430 4.410 3.620 4.440 ;
        RECT 2.860 4.320 3.180 4.360 ;
        RECT 2.280 4.230 2.490 4.240 ;
        RECT 2.300 4.200 2.490 4.230 ;
        RECT 2.920 4.160 3.090 4.320 ;
        RECT 3.430 4.240 3.870 4.410 ;
        RECT 3.430 4.210 3.620 4.240 ;
        RECT 0.070 4.130 0.330 4.150 ;
        RECT 0.070 4.080 0.410 4.130 ;
        RECT 0.070 4.020 0.560 4.080 ;
        RECT 0.070 3.990 0.580 4.020 ;
        RECT 0.110 3.960 0.580 3.990 ;
        RECT 0.240 3.910 0.580 3.960 ;
        RECT 0.360 3.900 0.580 3.910 ;
        RECT 0.370 3.870 0.580 3.900 ;
        RECT 0.390 3.790 0.580 3.870 ;
        RECT 1.750 3.790 2.080 3.910 ;
        RECT 4.150 3.820 4.320 4.500 ;
        RECT -0.100 3.740 0.070 3.760 ;
        RECT -0.120 3.310 0.090 3.740 ;
        RECT 0.390 3.620 0.910 3.790 ;
        RECT 0.390 3.590 0.580 3.620 ;
        RECT 1.260 3.610 3.160 3.790 ;
        RECT 3.890 3.780 4.320 3.820 ;
        RECT 3.540 3.620 4.320 3.780 ;
        RECT 3.540 3.610 4.080 3.620 ;
        RECT 3.890 3.590 4.080 3.610 ;
        RECT -0.120 2.590 0.090 3.020 ;
        RECT 0.390 2.710 0.580 2.740 ;
        RECT 3.890 2.720 4.080 2.740 ;
        RECT -0.100 2.570 0.070 2.590 ;
        RECT 0.390 2.540 0.910 2.710 ;
        RECT 1.260 2.540 3.160 2.720 ;
        RECT 3.540 2.710 4.080 2.720 ;
        RECT 3.540 2.550 4.320 2.710 ;
        RECT 0.390 2.460 0.580 2.540 ;
        RECT 0.370 2.430 0.580 2.460 ;
        RECT 0.360 2.420 0.580 2.430 ;
        RECT 1.750 2.420 2.080 2.540 ;
        RECT 3.890 2.510 4.320 2.550 ;
        RECT 0.240 2.370 0.580 2.420 ;
        RECT 0.110 2.340 0.580 2.370 ;
        RECT 0.070 2.310 0.580 2.340 ;
        RECT 0.070 2.250 0.560 2.310 ;
        RECT 0.070 2.200 0.410 2.250 ;
        RECT 0.070 2.180 0.330 2.200 ;
        RECT 0.070 2.160 0.300 2.180 ;
        RECT 0.070 2.120 0.280 2.160 ;
        RECT 0.070 1.840 0.240 2.120 ;
        RECT 1.420 2.010 1.590 2.170 ;
        RECT 2.300 2.100 2.490 2.130 ;
        RECT 2.280 2.090 2.490 2.100 ;
        RECT 1.290 1.970 1.610 2.010 ;
        RECT 1.290 1.780 1.620 1.970 ;
        RECT 2.030 1.920 2.490 2.090 ;
        RECT 2.920 2.010 3.090 2.170 ;
        RECT 3.430 2.090 3.620 2.120 ;
        RECT 2.300 1.900 2.490 1.920 ;
        RECT 2.860 1.970 3.180 2.010 ;
        RECT 2.860 1.780 3.190 1.970 ;
        RECT 3.430 1.920 3.870 2.090 ;
        RECT 3.430 1.890 3.620 1.920 ;
        RECT 4.150 1.830 4.320 2.510 ;
        RECT 1.290 1.750 1.610 1.780 ;
        RECT 2.860 1.750 3.180 1.780 ;
        RECT 1.290 1.350 1.610 1.380 ;
        RECT 2.860 1.350 3.180 1.380 ;
        RECT 0.070 1.010 0.240 1.290 ;
        RECT 1.290 1.160 1.620 1.350 ;
        RECT 2.300 1.210 2.490 1.230 ;
        RECT 1.290 1.120 1.610 1.160 ;
        RECT 0.070 0.970 0.280 1.010 ;
        RECT 0.070 0.950 0.300 0.970 ;
        RECT 1.420 0.960 1.590 1.120 ;
        RECT 2.030 1.040 2.490 1.210 ;
        RECT 2.860 1.160 3.190 1.350 ;
        RECT 3.430 1.210 3.620 1.240 ;
        RECT 2.860 1.120 3.180 1.160 ;
        RECT 2.280 1.030 2.490 1.040 ;
        RECT 2.300 1.000 2.490 1.030 ;
        RECT 2.920 0.960 3.090 1.120 ;
        RECT 3.430 1.040 3.870 1.210 ;
        RECT 3.430 1.010 3.620 1.040 ;
        RECT 0.070 0.930 0.330 0.950 ;
        RECT 0.070 0.880 0.410 0.930 ;
        RECT 0.070 0.820 0.560 0.880 ;
        RECT 0.070 0.790 0.580 0.820 ;
        RECT 0.110 0.760 0.580 0.790 ;
        RECT 0.240 0.710 0.580 0.760 ;
        RECT 0.360 0.700 0.580 0.710 ;
        RECT 0.370 0.670 0.580 0.700 ;
        RECT 0.390 0.590 0.580 0.670 ;
        RECT 1.750 0.590 2.080 0.710 ;
        RECT 4.150 0.620 4.320 1.300 ;
        RECT -0.100 0.540 0.070 0.560 ;
        RECT -0.120 0.110 0.090 0.540 ;
        RECT 0.390 0.420 0.910 0.590 ;
        RECT 0.390 0.390 0.580 0.420 ;
        RECT 1.260 0.410 3.160 0.590 ;
        RECT 3.890 0.580 4.320 0.620 ;
        RECT 3.540 0.420 4.320 0.580 ;
        RECT 3.540 0.410 4.080 0.420 ;
        RECT 3.890 0.390 4.080 0.410 ;
        RECT -0.120 -0.610 0.090 -0.180 ;
        RECT 0.390 -0.490 0.580 -0.460 ;
        RECT 3.890 -0.480 4.080 -0.460 ;
        RECT -0.100 -0.630 0.070 -0.610 ;
        RECT 0.390 -0.660 0.910 -0.490 ;
        RECT 1.260 -0.660 3.160 -0.480 ;
        RECT 3.540 -0.490 4.080 -0.480 ;
        RECT 3.540 -0.650 4.320 -0.490 ;
        RECT 0.390 -0.740 0.580 -0.660 ;
        RECT 0.370 -0.770 0.580 -0.740 ;
        RECT 0.360 -0.780 0.580 -0.770 ;
        RECT 1.750 -0.780 2.080 -0.660 ;
        RECT 3.890 -0.690 4.320 -0.650 ;
        RECT 0.240 -0.830 0.580 -0.780 ;
        RECT 0.110 -0.860 0.580 -0.830 ;
        RECT 0.070 -0.890 0.580 -0.860 ;
        RECT 0.070 -0.950 0.560 -0.890 ;
        RECT 0.070 -1.000 0.410 -0.950 ;
        RECT 0.070 -1.020 0.330 -1.000 ;
        RECT 0.070 -1.040 0.300 -1.020 ;
        RECT 0.070 -1.080 0.280 -1.040 ;
        RECT 0.070 -1.360 0.240 -1.080 ;
        RECT 1.420 -1.190 1.590 -1.030 ;
        RECT 2.300 -1.100 2.490 -1.070 ;
        RECT 2.280 -1.110 2.490 -1.100 ;
        RECT 1.290 -1.230 1.610 -1.190 ;
        RECT 1.290 -1.420 1.620 -1.230 ;
        RECT 2.030 -1.280 2.490 -1.110 ;
        RECT 2.920 -1.190 3.090 -1.030 ;
        RECT 3.430 -1.110 3.620 -1.080 ;
        RECT 2.300 -1.300 2.490 -1.280 ;
        RECT 2.860 -1.230 3.180 -1.190 ;
        RECT 2.860 -1.420 3.190 -1.230 ;
        RECT 3.430 -1.280 3.870 -1.110 ;
        RECT 3.430 -1.310 3.620 -1.280 ;
        RECT 4.150 -1.370 4.320 -0.690 ;
        RECT 1.290 -1.450 1.610 -1.420 ;
        RECT 2.860 -1.450 3.180 -1.420 ;
      LAYER mcon ;
        RECT 1.350 4.370 1.520 4.540 ;
        RECT 2.310 4.230 2.480 4.400 ;
        RECT 2.920 4.370 3.090 4.540 ;
        RECT 3.440 4.240 3.610 4.410 ;
        RECT -0.100 3.590 0.070 3.760 ;
        RECT 0.400 3.620 0.570 3.790 ;
        RECT 3.900 3.620 4.070 3.790 ;
        RECT 0.400 2.540 0.570 2.710 ;
        RECT 3.900 2.540 4.070 2.710 ;
        RECT 1.350 1.790 1.520 1.960 ;
        RECT 2.310 1.930 2.480 2.100 ;
        RECT 2.920 1.790 3.090 1.960 ;
        RECT 3.440 1.920 3.610 2.090 ;
        RECT 1.350 1.170 1.520 1.340 ;
        RECT 2.310 1.030 2.480 1.200 ;
        RECT 2.920 1.170 3.090 1.340 ;
        RECT 3.440 1.040 3.610 1.210 ;
        RECT -0.100 0.390 0.070 0.560 ;
        RECT 0.400 0.420 0.570 0.590 ;
        RECT 3.900 0.420 4.070 0.590 ;
        RECT 0.400 -0.660 0.570 -0.490 ;
        RECT 3.900 -0.660 4.070 -0.490 ;
        RECT 1.350 -1.410 1.520 -1.240 ;
        RECT 2.310 -1.270 2.480 -1.100 ;
        RECT 2.920 -1.410 3.090 -1.240 ;
        RECT 3.440 -1.280 3.610 -1.110 ;
      LAYER met1 ;
        RECT 1.280 4.290 1.600 4.610 ;
        RECT 2.280 4.170 2.510 4.460 ;
        RECT 2.850 4.290 3.170 4.610 ;
        RECT 3.410 4.180 3.640 4.470 ;
        RECT -0.130 3.630 0.100 3.820 ;
        RECT 2.300 3.700 2.490 4.170 ;
        RECT -0.130 3.530 0.220 3.630 ;
        RECT -0.120 3.310 0.220 3.530 ;
        RECT 2.230 3.380 2.490 3.700 ;
        RECT 3.410 3.690 3.600 4.180 ;
        RECT 3.230 3.440 3.600 3.690 ;
        RECT 3.230 3.370 3.500 3.440 ;
        RECT -0.120 2.800 0.220 3.020 ;
        RECT -0.130 2.700 0.220 2.800 ;
        RECT -0.130 2.510 0.100 2.700 ;
        RECT 2.230 2.630 2.490 2.950 ;
        RECT 3.230 2.890 3.500 2.960 ;
        RECT 3.230 2.640 3.600 2.890 ;
        RECT 2.300 2.160 2.490 2.630 ;
        RECT 1.280 1.720 1.600 2.040 ;
        RECT 2.280 1.870 2.510 2.160 ;
        RECT 3.410 2.150 3.600 2.640 ;
        RECT 2.850 1.720 3.170 2.040 ;
        RECT 3.410 1.860 3.640 2.150 ;
        RECT 1.280 1.090 1.600 1.410 ;
        RECT 2.280 0.970 2.510 1.260 ;
        RECT 2.850 1.090 3.170 1.410 ;
        RECT 3.410 0.980 3.640 1.270 ;
        RECT -0.130 0.430 0.100 0.620 ;
        RECT 2.300 0.500 2.490 0.970 ;
        RECT -0.130 0.330 0.220 0.430 ;
        RECT -0.120 0.110 0.220 0.330 ;
        RECT 2.230 0.180 2.490 0.500 ;
        RECT 3.410 0.490 3.600 0.980 ;
        RECT 3.230 0.240 3.600 0.490 ;
        RECT 3.230 0.170 3.500 0.240 ;
        RECT -0.120 -0.400 0.220 -0.180 ;
        RECT -0.130 -0.500 0.220 -0.400 ;
        RECT -0.130 -0.690 0.100 -0.500 ;
        RECT 2.230 -0.570 2.490 -0.250 ;
        RECT 3.230 -0.310 3.500 -0.240 ;
        RECT 3.230 -0.560 3.600 -0.310 ;
        RECT 2.300 -1.040 2.490 -0.570 ;
        RECT 1.280 -1.480 1.600 -1.160 ;
        RECT 2.280 -1.330 2.510 -1.040 ;
        RECT 3.410 -1.050 3.600 -0.560 ;
        RECT 2.850 -1.480 3.170 -1.160 ;
        RECT 3.410 -1.340 3.640 -1.050 ;
      LAYER via ;
        RECT 1.310 4.320 1.570 4.580 ;
        RECT 2.880 4.320 3.140 4.580 ;
        RECT -0.040 3.340 0.220 3.600 ;
        RECT 2.230 3.410 2.490 3.670 ;
        RECT 3.240 3.400 3.500 3.660 ;
        RECT -0.040 2.730 0.220 2.990 ;
        RECT 2.230 2.660 2.490 2.920 ;
        RECT 3.240 2.670 3.500 2.930 ;
        RECT 1.310 1.750 1.570 2.010 ;
        RECT 2.880 1.750 3.140 2.010 ;
        RECT 1.310 1.120 1.570 1.380 ;
        RECT 2.880 1.120 3.140 1.380 ;
        RECT -0.040 0.140 0.220 0.400 ;
        RECT 2.230 0.210 2.490 0.470 ;
        RECT 3.240 0.200 3.500 0.460 ;
        RECT -0.040 -0.470 0.220 -0.210 ;
        RECT 2.230 -0.540 2.490 -0.280 ;
        RECT 3.240 -0.530 3.500 -0.270 ;
        RECT 1.310 -1.450 1.570 -1.190 ;
        RECT 2.880 -1.450 3.140 -1.190 ;
  END
END sky130_hilas_Tgate4Single01

MACRO sky130_hilas_VinjDecode2to4
  CLASS BLOCK ;
  FOREIGN sky130_hilas_VinjDecode2to4 ;
  ORIGIN 6.370 -0.540 ;
  SIZE 12.950 BY 6.160 ;
  PIN OUTPUT00
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 3.200 5.550 3.570 5.630 ;
        RECT 3.200 5.540 4.230 5.550 ;
        RECT 6.110 5.540 6.420 5.700 ;
        RECT 3.200 5.370 6.580 5.540 ;
    END
  END OUTPUT00
  PIN OUTPUT01
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 3.200 4.040 3.570 4.120 ;
        RECT 3.200 4.030 4.230 4.040 ;
        RECT 6.110 4.030 6.420 4.190 ;
        RECT 3.200 3.860 6.580 4.030 ;
    END
  END OUTPUT01
  PIN OUTPUT10
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 3.200 2.530 3.570 2.610 ;
        RECT 3.200 2.520 4.230 2.530 ;
        RECT 6.110 2.520 6.420 2.680 ;
        RECT 3.200 2.350 6.580 2.520 ;
    END
  END OUTPUT10
  PIN OUTPUT11
    ANTENNADIFFAREA 0.275500 ;
    PORT
      LAYER met2 ;
        RECT 3.200 1.030 3.570 1.110 ;
        RECT 3.200 1.020 4.230 1.030 ;
        RECT 6.110 1.020 6.420 1.180 ;
        RECT 3.200 0.850 6.580 1.020 ;
    END
  END OUTPUT11
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 5.290 0.630 5.560 6.670 ;
    END
    PORT
      LAYER met1 ;
        RECT -3.190 2.130 -2.960 6.660 ;
    END
  END VGND
  PIN VINJ
    ANTENNADIFFAREA 0.914000 ;
    PORT
      LAYER nwell ;
        RECT -0.290 0.540 3.150 6.700 ;
      LAYER met1 ;
        RECT 0.320 6.320 0.540 6.660 ;
        RECT 0.320 6.060 0.550 6.320 ;
        RECT 0.320 5.660 0.540 6.060 ;
        RECT 0.320 5.350 0.570 5.660 ;
        RECT 0.320 4.810 0.540 5.350 ;
        RECT 0.320 4.550 0.550 4.810 ;
        RECT 0.320 4.150 0.540 4.550 ;
        RECT 0.320 3.840 0.570 4.150 ;
        RECT 0.320 3.300 0.540 3.840 ;
        RECT 0.320 3.040 0.550 3.300 ;
        RECT 0.320 2.640 0.540 3.040 ;
        RECT 0.320 2.330 0.570 2.640 ;
        RECT 0.320 1.800 0.540 2.330 ;
        RECT 0.320 1.540 0.550 1.800 ;
        RECT 0.320 1.140 0.540 1.540 ;
        RECT 0.320 0.830 0.570 1.140 ;
        RECT 0.320 0.630 0.540 0.830 ;
    END
    PORT
      LAYER nwell ;
        RECT -6.370 2.040 -4.390 6.700 ;
      LAYER met1 ;
        RECT -5.760 6.320 -5.540 6.660 ;
        RECT -5.760 6.060 -5.530 6.320 ;
        RECT -5.760 5.660 -5.540 6.060 ;
        RECT -5.760 5.350 -5.510 5.660 ;
        RECT -5.760 4.810 -5.540 5.350 ;
        RECT -5.760 4.550 -5.530 4.810 ;
        RECT -5.760 4.150 -5.540 4.550 ;
        RECT -5.760 3.840 -5.510 4.150 ;
        RECT -5.760 3.300 -5.540 3.840 ;
        RECT -5.760 3.040 -5.530 3.300 ;
        RECT -5.760 2.640 -5.540 3.040 ;
        RECT -5.760 2.330 -5.510 2.640 ;
        RECT -5.760 2.130 -5.540 2.330 ;
    END
  END VINJ
  PIN IN2
    ANTENNAGATEAREA 0.642800 ;
    PORT
      LAYER met2 ;
        RECT -1.810 6.060 -1.480 6.120 ;
        RECT 2.340 6.080 2.670 6.160 ;
        RECT 2.070 6.060 2.670 6.080 ;
        RECT -1.810 5.900 2.670 6.060 ;
        RECT -1.810 5.850 -1.480 5.900 ;
        RECT -6.370 4.740 -1.580 4.760 ;
        RECT -6.370 4.580 -1.530 4.740 ;
        RECT -1.800 4.550 -1.530 4.580 ;
        RECT -1.800 4.410 -1.520 4.550 ;
        RECT -1.750 4.390 -1.520 4.410 ;
        RECT -1.830 3.040 -1.500 3.100 ;
        RECT 2.340 3.060 2.670 3.140 ;
        RECT 2.070 3.040 2.670 3.060 ;
        RECT -1.830 2.880 2.670 3.040 ;
        RECT -1.830 2.830 -1.500 2.880 ;
    END
  END IN2
  PIN IN1
    ANTENNAGATEAREA 0.673600 ;
    PORT
      LAYER met2 ;
        RECT -2.660 6.500 3.740 6.510 ;
        RECT -2.680 6.350 3.740 6.500 ;
        RECT -2.680 6.340 -2.410 6.350 ;
        RECT -2.710 6.270 -2.410 6.340 ;
        RECT -6.370 6.090 -2.410 6.270 ;
        RECT 3.320 6.120 3.740 6.350 ;
        RECT -2.710 6.010 -2.440 6.090 ;
        RECT -2.740 5.170 -2.410 5.230 ;
        RECT -2.740 5.010 -1.100 5.170 ;
        RECT -2.740 4.960 -2.410 5.010 ;
        RECT -1.260 5.000 -1.100 5.010 ;
        RECT -1.260 4.840 3.740 5.000 ;
        RECT 3.320 4.610 3.740 4.840 ;
    END
  END IN1
  PIN ENABLE
    PORT
      LAYER met2 ;
        RECT -6.370 3.070 -2.760 3.250 ;
    END
  END ENABLE
  OBS
      LAYER li1 ;
        RECT -5.750 6.270 -5.580 6.410 ;
        RECT 0.330 6.270 0.500 6.410 ;
        RECT 1.060 6.290 1.230 6.370 ;
        RECT 1.870 6.290 2.040 6.370 ;
        RECT 3.410 6.330 3.580 6.450 ;
        RECT -5.750 6.100 -5.560 6.270 ;
        RECT -5.750 6.000 -5.580 6.100 ;
        RECT -6.180 5.620 -6.010 5.720 ;
        RECT -6.200 5.450 -6.010 5.620 ;
        RECT -6.180 5.390 -6.010 5.450 ;
        RECT -5.760 5.660 -5.590 5.720 ;
        RECT -5.760 5.390 -5.510 5.660 ;
        RECT -5.020 5.640 -4.770 5.720 ;
        RECT -5.020 5.470 -3.720 5.640 ;
        RECT -3.160 5.630 -2.990 6.260 ;
        RECT 0.330 6.100 0.520 6.270 ;
        RECT 0.330 6.000 0.500 6.100 ;
        RECT 1.060 5.720 1.270 6.290 ;
        RECT 1.830 6.040 2.040 6.290 ;
        RECT 2.430 6.110 2.600 6.210 ;
        RECT 3.370 6.160 3.580 6.330 ;
        RECT 5.300 6.260 5.560 6.330 ;
        RECT 6.100 6.260 6.280 6.390 ;
        RECT 3.410 6.120 3.580 6.160 ;
        RECT 1.830 5.720 2.000 6.040 ;
        RECT 2.400 5.940 2.600 6.110 ;
        RECT 2.430 5.840 2.600 5.940 ;
        RECT 3.970 6.080 4.840 6.250 ;
        RECT 5.300 6.080 6.280 6.260 ;
        RECT -5.750 5.370 -5.510 5.390 ;
        RECT -4.940 5.380 -4.770 5.470 ;
        RECT -3.240 5.460 -2.910 5.630 ;
        RECT -0.100 5.620 0.070 5.720 ;
        RECT -0.120 5.450 0.070 5.620 ;
        RECT -0.100 5.390 0.070 5.450 ;
        RECT 0.320 5.660 0.490 5.720 ;
        RECT 0.320 5.390 0.570 5.660 ;
        RECT 1.060 5.470 1.310 5.720 ;
        RECT 0.330 5.370 0.570 5.390 ;
        RECT 1.140 5.380 1.310 5.470 ;
        RECT 1.790 5.470 2.000 5.720 ;
        RECT 3.970 5.640 4.140 6.080 ;
        RECT 5.300 5.640 5.560 6.080 ;
        RECT 6.100 5.970 6.280 6.080 ;
        RECT 2.510 5.470 4.140 5.640 ;
        RECT 4.590 5.470 5.560 5.640 ;
        RECT 6.010 5.470 6.350 5.640 ;
        RECT 1.790 5.390 1.960 5.470 ;
        RECT 3.280 5.430 3.450 5.470 ;
        RECT -5.750 4.760 -5.580 4.900 ;
        RECT 0.330 4.760 0.500 4.900 ;
        RECT 1.060 4.780 1.230 4.860 ;
        RECT 1.870 4.780 2.040 4.860 ;
        RECT 3.410 4.820 3.580 4.940 ;
        RECT -5.750 4.590 -5.560 4.760 ;
        RECT -5.750 4.490 -5.580 4.590 ;
        RECT -6.180 4.110 -6.010 4.210 ;
        RECT -6.200 3.940 -6.010 4.110 ;
        RECT -6.180 3.880 -6.010 3.940 ;
        RECT -5.760 4.150 -5.590 4.210 ;
        RECT -5.760 3.880 -5.510 4.150 ;
        RECT -5.020 4.130 -4.770 4.210 ;
        RECT -5.020 3.960 -3.720 4.130 ;
        RECT -3.160 4.120 -2.990 4.750 ;
        RECT 0.330 4.590 0.520 4.760 ;
        RECT 0.330 4.490 0.500 4.590 ;
        RECT 1.060 4.210 1.270 4.780 ;
        RECT 1.830 4.530 2.040 4.780 ;
        RECT 2.430 4.600 2.600 4.700 ;
        RECT 3.370 4.650 3.580 4.820 ;
        RECT 5.300 4.750 5.560 4.820 ;
        RECT 6.100 4.750 6.280 4.880 ;
        RECT 3.410 4.610 3.580 4.650 ;
        RECT 1.830 4.210 2.000 4.530 ;
        RECT 2.400 4.430 2.600 4.600 ;
        RECT 2.430 4.330 2.600 4.430 ;
        RECT 3.970 4.570 4.840 4.740 ;
        RECT 5.300 4.570 6.280 4.750 ;
        RECT -5.750 3.860 -5.510 3.880 ;
        RECT -4.940 3.870 -4.770 3.960 ;
        RECT -3.240 3.950 -2.910 4.120 ;
        RECT -0.100 4.110 0.070 4.210 ;
        RECT -0.120 3.940 0.070 4.110 ;
        RECT -0.100 3.880 0.070 3.940 ;
        RECT 0.320 4.150 0.490 4.210 ;
        RECT 0.320 3.880 0.570 4.150 ;
        RECT 1.060 3.960 1.310 4.210 ;
        RECT 0.330 3.860 0.570 3.880 ;
        RECT 1.140 3.870 1.310 3.960 ;
        RECT 1.790 3.960 2.000 4.210 ;
        RECT 3.970 4.130 4.140 4.570 ;
        RECT 5.300 4.130 5.560 4.570 ;
        RECT 6.100 4.460 6.280 4.570 ;
        RECT 2.510 3.960 4.140 4.130 ;
        RECT 4.590 3.960 5.560 4.130 ;
        RECT 6.010 3.960 6.350 4.130 ;
        RECT 1.790 3.880 1.960 3.960 ;
        RECT 3.280 3.920 3.450 3.960 ;
        RECT -5.750 3.250 -5.580 3.390 ;
        RECT 0.330 3.250 0.500 3.390 ;
        RECT 1.060 3.270 1.230 3.350 ;
        RECT 1.870 3.270 2.040 3.350 ;
        RECT 3.410 3.310 3.580 3.430 ;
        RECT -5.750 3.080 -5.560 3.250 ;
        RECT -5.750 2.980 -5.580 3.080 ;
        RECT -6.180 2.600 -6.010 2.700 ;
        RECT -6.200 2.430 -6.010 2.600 ;
        RECT -6.180 2.370 -6.010 2.430 ;
        RECT -5.760 2.640 -5.590 2.700 ;
        RECT -5.760 2.370 -5.510 2.640 ;
        RECT -5.020 2.620 -4.770 2.700 ;
        RECT -5.020 2.450 -3.720 2.620 ;
        RECT -3.160 2.610 -2.990 3.240 ;
        RECT 0.330 3.080 0.520 3.250 ;
        RECT 0.330 2.980 0.500 3.080 ;
        RECT 1.060 2.700 1.270 3.270 ;
        RECT 1.830 3.020 2.040 3.270 ;
        RECT 2.430 3.090 2.600 3.190 ;
        RECT 3.370 3.140 3.580 3.310 ;
        RECT 5.300 3.240 5.560 3.310 ;
        RECT 6.100 3.240 6.280 3.370 ;
        RECT 3.410 3.100 3.580 3.140 ;
        RECT 1.830 2.700 2.000 3.020 ;
        RECT 2.400 2.920 2.600 3.090 ;
        RECT 2.430 2.820 2.600 2.920 ;
        RECT 3.970 3.060 4.840 3.230 ;
        RECT 5.300 3.060 6.280 3.240 ;
        RECT -5.750 2.350 -5.510 2.370 ;
        RECT -4.940 2.360 -4.770 2.450 ;
        RECT -3.240 2.440 -2.910 2.610 ;
        RECT -0.100 2.600 0.070 2.700 ;
        RECT -0.120 2.430 0.070 2.600 ;
        RECT -0.100 2.370 0.070 2.430 ;
        RECT 0.320 2.640 0.490 2.700 ;
        RECT 0.320 2.370 0.570 2.640 ;
        RECT 1.060 2.450 1.310 2.700 ;
        RECT 0.330 2.350 0.570 2.370 ;
        RECT 1.140 2.360 1.310 2.450 ;
        RECT 1.790 2.450 2.000 2.700 ;
        RECT 3.970 2.620 4.140 3.060 ;
        RECT 5.300 2.620 5.560 3.060 ;
        RECT 6.100 2.950 6.280 3.060 ;
        RECT 2.510 2.450 4.140 2.620 ;
        RECT 4.590 2.450 5.560 2.620 ;
        RECT 6.010 2.450 6.350 2.620 ;
        RECT 1.790 2.370 1.960 2.450 ;
        RECT 3.280 2.410 3.450 2.450 ;
        RECT 0.330 1.750 0.500 1.890 ;
        RECT 1.060 1.770 1.230 1.850 ;
        RECT 1.870 1.770 2.040 1.850 ;
        RECT 3.410 1.810 3.580 1.930 ;
        RECT 0.330 1.580 0.520 1.750 ;
        RECT 0.330 1.480 0.500 1.580 ;
        RECT 1.060 1.200 1.270 1.770 ;
        RECT 1.830 1.520 2.040 1.770 ;
        RECT 2.430 1.590 2.600 1.690 ;
        RECT 3.370 1.640 3.580 1.810 ;
        RECT 5.300 1.740 5.560 1.810 ;
        RECT 6.100 1.740 6.280 1.870 ;
        RECT 3.410 1.600 3.580 1.640 ;
        RECT 1.830 1.200 2.000 1.520 ;
        RECT 2.400 1.420 2.600 1.590 ;
        RECT 2.430 1.320 2.600 1.420 ;
        RECT 3.970 1.560 4.840 1.730 ;
        RECT 5.300 1.560 6.280 1.740 ;
        RECT -0.100 1.100 0.070 1.200 ;
        RECT -0.120 0.930 0.070 1.100 ;
        RECT -0.100 0.870 0.070 0.930 ;
        RECT 0.320 1.140 0.490 1.200 ;
        RECT 0.320 0.870 0.570 1.140 ;
        RECT 1.060 0.950 1.310 1.200 ;
        RECT 0.330 0.850 0.570 0.870 ;
        RECT 1.140 0.860 1.310 0.950 ;
        RECT 1.790 0.950 2.000 1.200 ;
        RECT 3.970 1.120 4.140 1.560 ;
        RECT 5.300 1.120 5.560 1.560 ;
        RECT 6.100 1.450 6.280 1.560 ;
        RECT 2.510 0.950 4.140 1.120 ;
        RECT 4.590 0.950 5.560 1.120 ;
        RECT 6.010 0.950 6.350 1.120 ;
        RECT 1.790 0.870 1.960 0.950 ;
        RECT 3.280 0.910 3.450 0.950 ;
      LAYER mcon ;
        RECT -5.730 6.100 -5.560 6.270 ;
        RECT 0.350 6.100 0.520 6.270 ;
        RECT -3.160 5.740 -2.990 5.910 ;
        RECT -5.720 5.420 -5.550 5.590 ;
        RECT -4.380 5.470 -4.210 5.640 ;
        RECT 0.360 5.420 0.530 5.590 ;
        RECT 5.330 5.760 5.510 5.940 ;
        RECT -5.730 4.590 -5.560 4.760 ;
        RECT 0.350 4.590 0.520 4.760 ;
        RECT -3.160 4.230 -2.990 4.400 ;
        RECT -5.720 3.910 -5.550 4.080 ;
        RECT -4.380 3.960 -4.210 4.130 ;
        RECT 0.360 3.910 0.530 4.080 ;
        RECT 5.330 4.250 5.510 4.430 ;
        RECT -5.730 3.080 -5.560 3.250 ;
        RECT 0.350 3.080 0.520 3.250 ;
        RECT -3.160 2.720 -2.990 2.890 ;
        RECT -5.720 2.400 -5.550 2.570 ;
        RECT -4.380 2.450 -4.210 2.620 ;
        RECT 0.360 2.400 0.530 2.570 ;
        RECT 5.330 2.740 5.510 2.920 ;
        RECT 0.350 1.580 0.520 1.750 ;
        RECT 0.360 0.900 0.530 1.070 ;
        RECT 5.330 1.240 5.510 1.420 ;
      LAYER met1 ;
        RECT -2.700 6.310 -2.430 6.600 ;
        RECT -2.740 6.040 -2.410 6.310 ;
        RECT -6.290 5.380 -5.980 5.730 ;
        RECT -4.460 5.420 -4.140 5.680 ;
        RECT -2.700 5.260 -2.430 6.040 ;
        RECT -2.710 4.930 -2.430 5.260 ;
        RECT -2.700 4.900 -2.430 4.930 ;
        RECT -6.290 3.870 -5.980 4.220 ;
        RECT -4.460 3.910 -4.140 4.170 ;
        RECT -2.240 3.580 -1.970 5.700 ;
        RECT -1.780 4.710 -1.510 6.170 ;
        RECT 2.340 5.900 2.670 6.160 ;
        RECT 3.310 6.120 3.740 6.410 ;
        RECT -0.830 5.670 -0.540 5.720 ;
        RECT -0.850 5.320 -0.540 5.670 ;
        RECT -0.210 5.380 0.100 5.730 ;
        RECT 3.180 5.370 3.570 5.640 ;
        RECT 6.110 5.380 6.420 5.700 ;
        RECT -1.830 4.440 -1.500 4.710 ;
        RECT -2.250 3.250 -1.970 3.580 ;
        RECT -6.290 2.360 -5.980 2.710 ;
        RECT -4.460 2.400 -4.140 2.660 ;
        RECT -2.240 2.080 -1.970 3.250 ;
        RECT -1.780 3.130 -1.510 4.440 ;
        RECT -1.800 2.800 -1.510 3.130 ;
        RECT -1.780 2.780 -1.510 2.800 ;
        RECT -1.310 4.170 -1.040 4.230 ;
        RECT -1.310 3.840 -1.030 4.170 ;
        RECT -2.240 1.750 -1.940 2.080 ;
        RECT -2.240 1.700 -1.970 1.750 ;
        RECT -1.310 1.630 -1.040 3.840 ;
        RECT -1.330 1.300 -1.040 1.630 ;
        RECT -1.310 1.270 -1.040 1.300 ;
        RECT -0.830 2.670 -0.540 5.320 ;
        RECT 2.340 4.390 2.670 4.650 ;
        RECT 3.310 4.610 3.740 4.900 ;
        RECT -0.210 3.870 0.100 4.220 ;
        RECT 3.180 3.860 3.570 4.130 ;
        RECT 6.110 3.870 6.420 4.190 ;
        RECT 2.340 2.880 2.670 3.140 ;
        RECT 3.310 3.100 3.740 3.390 ;
        RECT -0.830 2.320 -0.530 2.670 ;
        RECT -0.210 2.360 0.100 2.710 ;
        RECT 3.180 2.350 3.570 2.620 ;
        RECT 6.110 2.360 6.420 2.680 ;
        RECT -0.830 0.780 -0.540 2.320 ;
        RECT 2.340 1.380 2.670 1.640 ;
        RECT 3.310 1.600 3.740 1.890 ;
        RECT -0.210 0.860 0.100 1.210 ;
        RECT 3.180 0.850 3.570 1.120 ;
        RECT 6.110 0.860 6.420 1.180 ;
      LAYER via ;
        RECT -2.710 6.040 -2.440 6.310 ;
        RECT -6.260 5.410 -6.000 5.670 ;
        RECT -4.430 5.420 -4.170 5.680 ;
        RECT -1.780 5.850 -1.510 6.120 ;
        RECT 2.380 5.900 2.640 6.160 ;
        RECT 3.370 6.150 3.630 6.410 ;
        RECT -2.710 4.960 -2.440 5.230 ;
        RECT -2.240 5.360 -1.970 5.630 ;
        RECT -6.260 3.900 -6.000 4.160 ;
        RECT -4.430 3.910 -4.170 4.170 ;
        RECT -0.850 5.350 -0.560 5.640 ;
        RECT -0.180 5.410 0.080 5.670 ;
        RECT 3.240 5.370 3.500 5.630 ;
        RECT 6.140 5.410 6.400 5.670 ;
        RECT -1.800 4.440 -1.530 4.710 ;
        RECT -2.250 3.280 -1.980 3.550 ;
        RECT -6.260 2.390 -6.000 2.650 ;
        RECT -4.430 2.400 -4.170 2.660 ;
        RECT -1.800 2.830 -1.530 3.100 ;
        RECT -1.300 3.870 -1.030 4.140 ;
        RECT 2.380 4.390 2.640 4.650 ;
        RECT 3.370 4.640 3.630 4.900 ;
        RECT -0.810 3.840 -0.550 4.100 ;
        RECT -0.180 3.900 0.080 4.160 ;
        RECT 3.240 3.860 3.500 4.120 ;
        RECT 6.140 3.900 6.400 4.160 ;
        RECT -2.210 1.780 -1.940 2.050 ;
        RECT -1.330 1.330 -1.060 1.600 ;
        RECT 2.380 2.880 2.640 3.140 ;
        RECT 3.370 3.130 3.630 3.390 ;
        RECT -0.820 2.350 -0.530 2.640 ;
        RECT -0.180 2.390 0.080 2.650 ;
        RECT 3.240 2.350 3.500 2.610 ;
        RECT 6.140 2.390 6.400 2.650 ;
        RECT 2.380 1.380 2.640 1.640 ;
        RECT 3.370 1.630 3.630 1.890 ;
        RECT -0.830 0.810 -0.540 1.100 ;
        RECT -0.180 0.890 0.080 1.150 ;
        RECT 3.240 0.850 3.500 1.110 ;
        RECT 6.140 0.890 6.400 1.150 ;
      LAYER met2 ;
        RECT -6.290 5.570 -5.970 5.670 ;
        RECT -6.300 5.410 -5.970 5.570 ;
        RECT -4.460 5.600 -4.140 5.680 ;
        RECT -2.270 5.600 -1.940 5.630 ;
        RECT -4.460 5.420 -1.920 5.600 ;
        RECT -2.270 5.410 -1.920 5.420 ;
        RECT -0.880 5.570 -0.530 5.640 ;
        RECT -0.210 5.570 0.110 5.670 ;
        RECT -0.880 5.410 0.110 5.570 ;
        RECT -2.270 5.360 -1.940 5.410 ;
        RECT -0.880 5.350 -0.530 5.410 ;
        RECT 2.340 4.570 2.670 4.650 ;
        RECT 2.070 4.550 2.670 4.570 ;
        RECT -1.250 4.390 2.670 4.550 ;
        RECT -6.290 4.060 -5.970 4.160 ;
        RECT -6.300 3.900 -5.970 4.060 ;
        RECT -4.460 4.090 -4.140 4.170 ;
        RECT -1.250 4.140 -1.090 4.390 ;
        RECT -1.330 4.090 -1.000 4.140 ;
        RECT -4.460 3.910 -1.000 4.090 ;
        RECT -1.330 3.870 -1.000 3.910 ;
        RECT -0.840 4.060 -0.520 4.100 ;
        RECT -0.210 4.060 0.110 4.160 ;
        RECT -0.840 3.900 0.110 4.060 ;
        RECT -0.840 3.840 -0.520 3.900 ;
        RECT -2.280 3.490 -1.950 3.550 ;
        RECT -2.280 3.330 3.740 3.490 ;
        RECT -2.280 3.280 -1.950 3.330 ;
        RECT 3.320 3.100 3.740 3.330 ;
        RECT -6.290 2.550 -5.970 2.650 ;
        RECT -6.300 2.390 -5.970 2.550 ;
        RECT -4.460 2.580 -4.140 2.660 ;
        RECT -0.850 2.580 -0.500 2.640 ;
        RECT -4.460 2.550 -0.360 2.580 ;
        RECT -0.210 2.550 0.110 2.650 ;
        RECT -4.460 2.400 0.110 2.550 ;
        RECT -0.850 2.390 0.110 2.400 ;
        RECT -0.850 2.350 -0.500 2.390 ;
        RECT -2.240 1.990 -1.910 2.050 ;
        RECT -2.240 1.830 3.740 1.990 ;
        RECT -2.240 1.780 -1.910 1.830 ;
        RECT -1.360 1.540 -1.030 1.600 ;
        RECT 2.340 1.560 2.670 1.640 ;
        RECT 3.320 1.600 3.740 1.830 ;
        RECT 2.070 1.540 2.670 1.560 ;
        RECT -1.360 1.380 2.670 1.540 ;
        RECT -1.360 1.330 -1.030 1.380 ;
        RECT -0.860 1.050 -0.510 1.100 ;
        RECT -0.210 1.050 0.110 1.150 ;
        RECT -0.860 0.890 0.110 1.050 ;
        RECT -0.860 0.810 -0.510 0.890 ;
  END
END sky130_hilas_VinjDecode2to4

MACRO sky130_hilas_TA2Cell_1FG
  CLASS BLOCK ;
  FOREIGN sky130_hilas_TA2Cell_1FG ;
  ORIGIN 26.160 -1.350 ;
  SIZE 28.090 BY 6.150 ;
  PIN VIN12
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -16.850 2.660 -16.540 2.720 ;
        RECT -17.310 2.650 -16.540 2.660 ;
        RECT -17.310 2.640 -16.420 2.650 ;
        RECT -17.310 2.430 -14.630 2.640 ;
        RECT -17.310 2.410 -16.420 2.430 ;
        RECT -16.850 2.390 -16.540 2.410 ;
    END
  END VIN12
  PIN VIN11
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -16.880 6.370 -16.570 6.410 ;
        RECT -17.260 6.350 -16.420 6.370 ;
        RECT -17.260 6.170 -14.630 6.350 ;
        RECT -16.880 6.080 -16.570 6.170 ;
    END
  END VIN11
  PIN VIN21
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -2.200 4.750 -1.890 4.790 ;
        RECT -2.520 4.740 -1.860 4.750 ;
        RECT -2.520 4.510 -1.420 4.740 ;
        RECT -2.200 4.460 -1.890 4.510 ;
    END
  END VIN21
  PIN VIN22
    USE ANALOG ;
    ANTENNAGATEAREA 1.015000 ;
    PORT
      LAYER met2 ;
        RECT -1.960 7.430 -1.650 7.440 ;
        RECT -2.530 7.420 -1.650 7.430 ;
        RECT -2.600 7.180 -1.650 7.420 ;
        RECT -1.960 7.110 -1.650 7.180 ;
    END
  END VIN22
  PIN VPWR
    USE ANALOG ;
    ANTENNADIFFAREA 1.373600 ;
    PORT
      LAYER nwell ;
        RECT 0.650 1.400 1.930 7.450 ;
      LAYER met1 ;
        RECT 0.630 7.300 0.910 7.450 ;
        RECT 0.640 5.870 0.910 7.300 ;
        RECT 0.640 5.580 0.920 5.870 ;
        RECT 0.640 3.280 0.910 5.580 ;
        RECT 0.640 2.990 0.920 3.280 ;
        RECT 0.640 1.400 0.910 2.990 ;
    END
  END VPWR
  PIN VGND
    USE ANALOG ;
    ANTENNADIFFAREA 5.718600 ;
    PORT
      LAYER met2 ;
        RECT -17.680 4.290 -17.360 4.340 ;
        RECT -17.680 4.040 -11.660 4.290 ;
        RECT -11.980 3.970 -11.660 4.040 ;
        RECT -11.980 1.750 -11.660 1.760 ;
        RECT -1.540 1.750 -1.210 1.890 ;
        RECT -11.980 1.590 -1.210 1.750 ;
        RECT -11.980 1.580 -11.290 1.590 ;
        RECT -11.980 1.460 -11.660 1.580 ;
    END
    PORT
      LAYER met1 ;
        RECT -1.540 1.600 -1.210 1.890 ;
        RECT -0.030 1.600 0.310 7.450 ;
        RECT -1.550 1.570 -1.130 1.600 ;
        RECT -0.530 1.570 0.310 1.600 ;
        RECT -1.550 1.460 0.310 1.570 ;
        RECT -1.270 1.430 -0.370 1.460 ;
        RECT -0.030 1.400 0.310 1.460 ;
      LAYER via ;
        RECT -1.510 1.610 -1.240 1.870 ;
    END
    PORT
      LAYER met1 ;
        RECT -17.690 6.480 -17.460 7.450 ;
        RECT -17.700 6.230 -17.460 6.480 ;
        RECT -17.690 4.340 -17.460 6.230 ;
        RECT -17.690 4.040 -17.360 4.340 ;
        RECT -17.690 3.870 -17.440 4.040 ;
        RECT -17.690 1.400 -17.460 3.870 ;
      LAYER via ;
        RECT -17.650 4.060 -17.390 4.320 ;
    END
    PORT
      LAYER met1 ;
        RECT -11.900 4.290 -11.670 7.450 ;
        RECT -11.980 3.970 -11.660 4.290 ;
        RECT -11.900 1.760 -11.670 3.970 ;
        RECT -11.980 1.460 -11.660 1.760 ;
        RECT -11.900 1.400 -11.670 1.460 ;
      LAYER via ;
        RECT -11.950 4.000 -11.690 4.260 ;
        RECT -11.950 1.480 -11.690 1.740 ;
    END
  END VGND
  PIN VINJ
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -26.160 1.350 -22.850 7.500 ;
        RECT -6.510 7.450 -3.200 7.500 ;
        RECT -6.510 7.440 -1.730 7.450 ;
        RECT -6.510 1.400 -1.350 7.440 ;
        RECT -6.510 1.350 -3.200 1.400 ;
      LAYER met2 ;
        RECT -25.920 7.280 -25.600 7.400 ;
        RECT -3.720 7.280 -3.400 7.400 ;
        RECT -25.920 7.100 -3.400 7.280 ;
        RECT -4.590 4.590 -4.270 4.850 ;
        RECT -4.550 4.570 -3.370 4.590 ;
        RECT -4.550 4.310 -3.330 4.570 ;
        RECT -4.550 4.250 -3.370 4.310 ;
        RECT -4.590 4.240 -3.370 4.250 ;
        RECT -4.590 3.990 -4.270 4.240 ;
    END
    PORT
      LAYER met1 ;
        RECT -3.720 7.400 -3.440 7.450 ;
        RECT -3.720 7.100 -3.400 7.400 ;
        RECT -3.720 6.800 -3.440 7.100 ;
        RECT -3.830 6.200 -3.440 6.800 ;
        RECT -3.720 4.600 -3.440 6.200 ;
        RECT -3.720 4.280 -3.360 4.600 ;
        RECT -3.720 2.650 -3.440 4.280 ;
        RECT -3.830 2.050 -3.440 2.650 ;
        RECT -3.720 1.400 -3.440 2.050 ;
      LAYER via ;
        RECT -3.690 7.120 -3.430 7.380 ;
        RECT -3.620 4.310 -3.360 4.570 ;
    END
    PORT
      LAYER met1 ;
        RECT -25.920 7.400 -25.640 7.450 ;
        RECT -25.920 7.120 -25.600 7.400 ;
        RECT -25.920 6.800 -25.640 7.120 ;
        RECT -25.920 6.200 -25.530 6.800 ;
        RECT -25.920 2.650 -25.640 6.200 ;
        RECT -25.920 2.050 -25.530 2.650 ;
        RECT -25.920 1.400 -25.640 2.050 ;
      LAYER via ;
        RECT -25.890 7.130 -25.630 7.390 ;
    END
  END VINJ
  PIN OUTPUT1
    USE ANALOG ;
    ANTENNADIFFAREA 0.308800 ;
    PORT
      LAYER met2 ;
        RECT -0.990 4.970 -0.680 5.030 ;
        RECT 1.310 4.970 1.620 4.990 ;
        RECT -0.990 4.740 1.930 4.970 ;
        RECT -0.990 4.700 -0.680 4.740 ;
        RECT 1.310 4.660 1.620 4.740 ;
    END
  END OUTPUT1
  PIN OUTPUT2
    USE ANALOG ;
    ANTENNADIFFAREA 0.308800 ;
    PORT
      LAYER met2 ;
        RECT -0.990 4.140 -0.680 4.190 ;
        RECT 1.300 4.140 1.610 4.270 ;
        RECT -0.990 3.920 1.930 4.140 ;
        RECT -0.990 3.860 -0.680 3.920 ;
    END
  END OUTPUT2
  PIN DRAIN1
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER met2 ;
        RECT -23.990 6.950 -23.680 6.960 ;
        RECT -5.680 6.950 -5.370 6.960 ;
        RECT -26.160 6.770 -3.200 6.950 ;
        RECT -23.990 6.630 -23.680 6.770 ;
        RECT -5.680 6.630 -5.370 6.770 ;
    END
  END DRAIN1
  PIN DRAIN2
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER met2 ;
        RECT -23.990 2.080 -23.680 2.220 ;
        RECT -26.160 2.070 -23.680 2.080 ;
        RECT -5.680 2.080 -5.370 2.220 ;
        RECT -5.680 2.070 -3.200 2.080 ;
        RECT -26.160 1.920 -3.200 2.070 ;
        RECT -26.160 1.900 -23.680 1.920 ;
        RECT -23.990 1.890 -23.680 1.900 ;
        RECT -5.680 1.900 -3.200 1.920 ;
        RECT -5.680 1.890 -5.370 1.900 ;
    END
  END DRAIN2
  PIN COLSEL2
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT -25.390 5.990 -25.200 7.450 ;
        RECT -25.420 5.960 -25.200 5.990 ;
        RECT -25.430 5.690 -25.180 5.960 ;
        RECT -25.430 5.680 -25.190 5.690 ;
        RECT -25.420 5.440 -25.190 5.680 ;
        RECT -25.390 3.410 -25.230 5.440 ;
        RECT -25.420 3.170 -25.190 3.410 ;
        RECT -25.430 3.160 -25.190 3.170 ;
        RECT -25.430 2.890 -25.180 3.160 ;
        RECT -25.420 2.860 -25.200 2.890 ;
        RECT -25.390 1.400 -25.200 2.860 ;
    END
  END COLSEL2
  PIN GATE2
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT -21.120 5.060 -18.400 6.710 ;
        RECT -21.110 5.020 -18.400 5.060 ;
        RECT -21.110 3.690 -18.400 3.730 ;
        RECT -21.120 2.040 -18.400 3.690 ;
      LAYER met1 ;
        RECT -18.910 6.240 -18.680 7.450 ;
        RECT -18.940 5.450 -18.680 6.240 ;
        RECT -18.910 3.300 -18.680 5.450 ;
        RECT -18.940 2.510 -18.680 3.300 ;
        RECT -18.910 1.400 -18.680 2.510 ;
    END
  END GATE2
  PIN GATE1
    ANTENNADIFFAREA 1.718800 ;
    PORT
      LAYER nwell ;
        RECT -10.960 5.060 -8.240 6.710 ;
        RECT -10.960 5.020 -8.250 5.060 ;
        RECT -10.960 3.690 -8.250 3.730 ;
        RECT -10.960 2.040 -8.240 3.690 ;
      LAYER met1 ;
        RECT -10.680 6.240 -10.450 7.450 ;
        RECT -10.680 5.450 -10.420 6.240 ;
        RECT -10.680 3.300 -10.450 5.450 ;
        RECT -10.680 2.510 -10.420 3.300 ;
        RECT -10.680 1.400 -10.450 2.510 ;
    END
  END GATE1
  PIN COLSEL1
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT -4.160 5.990 -3.970 7.450 ;
        RECT -4.160 5.960 -3.940 5.990 ;
        RECT -4.180 5.690 -3.930 5.960 ;
        RECT -4.170 5.680 -3.930 5.690 ;
        RECT -4.170 5.440 -3.940 5.680 ;
        RECT -4.130 3.410 -3.970 5.440 ;
        RECT -4.170 3.170 -3.940 3.410 ;
        RECT -4.170 3.160 -3.930 3.170 ;
        RECT -4.180 2.890 -3.930 3.160 ;
        RECT -4.160 2.860 -3.940 2.890 ;
        RECT -4.160 1.400 -3.970 2.860 ;
    END
  END COLSEL1
  PIN VTUN
    ANTENNADIFFAREA 5.032200 ;
    PORT
      LAYER nwell ;
        RECT -16.370 6.700 -12.990 7.450 ;
        RECT -16.380 3.130 -12.980 6.700 ;
        RECT -16.370 1.410 -12.990 3.130 ;
      LAYER met1 ;
        RECT -15.400 7.290 -13.960 7.450 ;
        RECT -15.400 1.410 -14.980 7.290 ;
        RECT -14.380 1.400 -13.960 7.290 ;
    END
  END VTUN
  OBS
      LAYER li1 ;
        RECT -2.220 7.400 -2.050 7.450 ;
        RECT -25.760 6.770 -25.560 7.120 ;
        RECT -24.280 6.870 -23.750 7.040 ;
        RECT -25.770 6.740 -25.560 6.770 ;
        RECT -25.770 6.160 -25.550 6.740 ;
        RECT -25.770 6.150 -25.560 6.160 ;
        RECT -25.390 5.980 -25.200 5.990 ;
        RECT -25.400 5.690 -25.200 5.980 ;
        RECT -25.480 5.360 -25.190 5.690 ;
        RECT -25.000 4.880 -24.830 6.490 ;
        RECT -25.010 4.690 -24.830 4.880 ;
        RECT -24.170 5.960 -24.000 6.480 ;
        RECT -21.560 6.440 -16.500 7.270 ;
        RECT -2.220 7.140 -1.660 7.400 ;
        RECT -0.750 7.150 -0.550 7.190 ;
        RECT -2.220 7.120 -2.050 7.140 ;
        RECT -5.610 6.870 -5.080 7.040 ;
        RECT -3.800 6.770 -3.600 7.120 ;
        RECT -3.800 6.740 -3.590 6.770 ;
        RECT -17.050 6.360 -16.570 6.440 ;
        RECT -24.170 5.700 -23.840 5.960 ;
        RECT -24.170 4.790 -24.000 5.700 ;
        RECT -18.930 5.500 -18.700 6.190 ;
        RECT -17.050 6.110 -16.580 6.360 ;
        RECT -15.620 5.310 -15.070 5.740 ;
        RECT -14.290 5.310 -13.740 5.740 ;
        RECT -10.660 5.500 -10.430 6.190 ;
        RECT -5.360 5.960 -5.190 6.480 ;
        RECT -5.520 5.700 -5.190 5.960 ;
        RECT -17.860 4.470 -17.470 4.880 ;
        RECT -21.220 4.290 -17.470 4.470 ;
        RECT -25.010 3.970 -24.830 4.160 ;
        RECT -25.480 3.160 -25.190 3.490 ;
        RECT -25.400 2.870 -25.200 3.160 ;
        RECT -25.390 2.860 -25.200 2.870 ;
        RECT -25.770 2.690 -25.560 2.700 ;
        RECT -25.770 2.110 -25.550 2.690 ;
        RECT -25.000 2.360 -24.830 3.970 ;
        RECT -24.170 3.200 -24.000 4.060 ;
        RECT -17.860 3.870 -17.470 4.290 ;
        RECT -11.920 4.470 -11.500 4.880 ;
        RECT -5.360 4.790 -5.190 5.700 ;
        RECT -4.530 4.880 -4.360 6.490 ;
        RECT -3.810 6.160 -3.590 6.740 ;
        RECT -3.800 6.150 -3.590 6.160 ;
        RECT -2.800 6.040 -2.620 6.970 ;
        RECT -0.980 6.890 -0.550 7.150 ;
        RECT -2.070 6.710 -1.740 6.880 ;
        RECT -0.750 6.860 -0.550 6.890 ;
        RECT -1.990 6.570 -1.740 6.710 ;
        RECT -1.990 6.310 -1.510 6.570 ;
        RECT -1.160 6.500 -0.990 6.540 ;
        RECT -0.750 6.500 -0.550 6.530 ;
        RECT -2.920 6.010 -2.600 6.040 ;
        RECT -4.160 5.980 -3.970 5.990 ;
        RECT -4.160 5.690 -3.960 5.980 ;
        RECT -2.920 5.820 -2.590 6.010 ;
        RECT -2.920 5.780 -2.600 5.820 ;
        RECT -4.170 5.360 -3.880 5.690 ;
        RECT -4.530 4.690 -4.350 4.880 ;
        RECT -11.920 4.290 -8.140 4.470 ;
        RECT -15.620 3.580 -15.070 4.010 ;
        RECT -14.290 3.580 -13.740 4.010 ;
        RECT -11.920 3.870 -11.500 4.290 ;
        RECT -24.170 2.940 -23.840 3.200 ;
        RECT -24.170 2.370 -24.000 2.940 ;
        RECT -18.930 2.560 -18.700 3.290 ;
        RECT -16.890 2.430 -16.550 2.680 ;
        RECT -10.660 2.560 -10.430 3.290 ;
        RECT -5.360 3.200 -5.190 4.060 ;
        RECT -5.520 2.940 -5.190 3.200 ;
        RECT -16.890 2.350 -16.540 2.430 ;
        RECT -5.360 2.370 -5.190 2.940 ;
        RECT -4.530 3.970 -4.350 4.160 ;
        RECT -4.530 2.360 -4.360 3.970 ;
        RECT -4.170 3.160 -3.880 3.490 ;
        RECT -4.160 2.870 -3.960 3.160 ;
        RECT -4.160 2.860 -3.970 2.870 ;
        RECT -3.800 2.690 -3.590 2.700 ;
        RECT -25.770 2.080 -25.560 2.110 ;
        RECT -25.760 1.730 -25.560 2.080 ;
        RECT -24.280 1.810 -23.750 1.980 ;
        RECT -21.590 1.500 -16.540 2.350 ;
        RECT -3.810 2.110 -3.590 2.690 ;
        RECT -3.800 2.080 -3.590 2.110 ;
        RECT -5.610 1.810 -5.080 1.980 ;
        RECT -3.800 1.730 -3.600 2.080 ;
        RECT -2.800 1.870 -2.620 5.780 ;
        RECT -1.990 4.930 -1.820 6.310 ;
        RECT -1.160 6.240 -0.550 6.500 ;
        RECT -1.160 6.210 -0.990 6.240 ;
        RECT -0.750 6.200 -0.550 6.240 ;
        RECT -0.160 6.200 0.390 7.190 ;
        RECT 1.210 7.040 1.840 7.210 ;
        RECT 1.210 6.940 1.600 7.040 ;
        RECT 1.210 6.910 1.590 6.940 ;
        RECT 1.210 6.760 1.570 6.910 ;
        RECT 0.860 6.590 1.570 6.760 ;
        RECT 0.860 5.840 1.560 6.150 ;
        RECT -1.160 5.650 -0.990 5.680 ;
        RECT -0.750 5.650 -0.550 5.690 ;
        RECT -1.160 5.390 -0.550 5.650 ;
        RECT -1.160 5.350 -0.990 5.390 ;
        RECT -0.750 5.360 -0.550 5.390 ;
        RECT -0.750 5.000 -0.550 5.030 ;
        RECT -2.190 4.730 -1.870 4.760 ;
        RECT -0.980 4.740 -0.550 5.000 ;
        RECT -2.190 4.540 -1.860 4.730 ;
        RECT -0.750 4.700 -0.550 4.740 ;
        RECT -0.160 4.700 0.390 5.690 ;
        RECT 0.710 5.610 1.560 5.840 ;
        RECT 0.860 5.270 1.560 5.610 ;
        RECT 1.320 4.910 1.640 4.950 ;
        RECT 1.320 4.850 1.650 4.910 ;
        RECT 0.850 4.720 1.650 4.850 ;
        RECT 0.850 4.690 1.640 4.720 ;
        RECT 0.850 4.670 1.550 4.690 ;
        RECT -2.190 4.500 -1.870 4.540 ;
        RECT -2.190 4.420 -2.020 4.500 ;
        RECT -2.240 4.250 -2.020 4.420 ;
        RECT -2.240 4.090 -2.070 4.250 ;
        RECT 1.310 4.190 1.630 4.230 ;
        RECT -0.750 4.150 -0.550 4.190 ;
        RECT -1.710 3.830 -1.520 3.950 ;
        RECT -0.980 3.890 -0.550 4.150 ;
        RECT -0.750 3.860 -0.550 3.890 ;
        RECT -2.070 3.720 -1.520 3.830 ;
        RECT -2.070 3.660 -1.530 3.720 ;
        RECT -1.990 1.880 -1.820 3.660 ;
        RECT -1.160 3.500 -0.990 3.540 ;
        RECT -0.750 3.500 -0.550 3.530 ;
        RECT -1.160 3.240 -0.550 3.500 ;
        RECT -1.160 3.210 -0.990 3.240 ;
        RECT -0.750 3.200 -0.550 3.240 ;
        RECT -0.160 3.200 0.390 4.190 ;
        RECT 0.850 4.010 1.640 4.190 ;
        RECT 1.310 4.000 1.640 4.010 ;
        RECT 1.310 3.970 1.630 4.000 ;
        RECT 0.860 3.250 1.560 3.590 ;
        RECT 0.710 3.020 1.560 3.250 ;
        RECT 0.860 2.710 1.560 3.020 ;
        RECT -1.160 2.650 -0.990 2.680 ;
        RECT -0.750 2.650 -0.550 2.690 ;
        RECT -1.160 2.390 -0.550 2.650 ;
        RECT -1.160 2.350 -0.990 2.390 ;
        RECT -0.750 2.360 -0.550 2.390 ;
        RECT -0.750 2.000 -0.550 2.030 ;
        RECT -0.980 1.740 -0.550 2.000 ;
        RECT -0.750 1.700 -0.550 1.740 ;
        RECT -0.160 1.700 0.390 2.690 ;
        RECT 0.860 2.100 1.570 2.270 ;
        RECT 1.210 1.820 1.570 2.100 ;
        RECT 1.210 1.650 1.840 1.820 ;
      LAYER mcon ;
        RECT -23.930 6.870 -23.750 7.040 ;
        RECT -25.740 6.570 -25.570 6.740 ;
        RECT -25.390 5.730 -25.210 5.920 ;
        RECT -1.890 7.180 -1.720 7.350 ;
        RECT -3.790 6.570 -3.620 6.740 ;
        RECT -18.900 5.990 -18.730 6.160 ;
        RECT -16.810 6.150 -16.640 6.320 ;
        RECT -24.070 5.740 -23.900 5.910 ;
        RECT -10.630 5.990 -10.460 6.160 ;
        RECT -18.900 5.540 -18.730 5.710 ;
        RECT -15.340 5.390 -15.070 5.660 ;
        RECT -14.290 5.390 -14.020 5.660 ;
        RECT -10.630 5.540 -10.460 5.710 ;
        RECT -5.460 5.740 -5.290 5.910 ;
        RECT -17.660 4.640 -17.490 4.810 ;
        RECT -17.660 4.280 -17.490 4.450 ;
        RECT -25.390 2.930 -25.210 3.120 ;
        RECT -17.650 3.920 -17.480 4.090 ;
        RECT -11.870 4.640 -11.700 4.810 ;
        RECT -0.920 6.930 -0.750 7.100 ;
        RECT 0.060 6.610 0.230 6.780 ;
        RECT 1.330 6.950 1.500 7.120 ;
        RECT -1.740 6.350 -1.570 6.520 ;
        RECT -4.150 5.730 -3.970 5.920 ;
        RECT -2.860 5.830 -2.690 6.000 ;
        RECT -11.870 4.280 -11.700 4.450 ;
        RECT -15.340 3.660 -15.070 3.930 ;
        RECT -14.290 3.660 -14.020 3.930 ;
        RECT -11.870 3.920 -11.700 4.090 ;
        RECT -24.070 2.980 -23.900 3.150 ;
        RECT -18.900 3.040 -18.730 3.210 ;
        RECT -18.900 2.590 -18.730 2.760 ;
        RECT -10.630 3.040 -10.460 3.210 ;
        RECT -5.460 2.980 -5.290 3.150 ;
        RECT -16.780 2.460 -16.610 2.630 ;
        RECT -10.630 2.590 -10.460 2.760 ;
        RECT -4.150 2.930 -3.970 3.120 ;
        RECT -25.740 2.110 -25.570 2.280 ;
        RECT -23.930 1.810 -23.750 1.980 ;
        RECT -3.790 2.110 -3.620 2.280 ;
        RECT -0.970 6.280 -0.800 6.450 ;
        RECT -0.970 5.440 -0.800 5.610 ;
        RECT 0.720 5.640 0.890 5.810 ;
        RECT 0.060 5.110 0.230 5.280 ;
        RECT -0.920 4.790 -0.750 4.960 ;
        RECT -2.130 4.550 -1.960 4.720 ;
        RECT 1.380 4.730 1.550 4.900 ;
        RECT -1.700 3.750 -1.530 3.920 ;
        RECT -0.920 3.930 -0.750 4.100 ;
        RECT 1.370 4.010 1.540 4.180 ;
        RECT 0.060 3.610 0.230 3.780 ;
        RECT -0.970 3.280 -0.800 3.450 ;
        RECT 0.720 3.050 0.890 3.220 ;
        RECT -0.970 2.440 -0.800 2.610 ;
        RECT 0.060 2.110 0.230 2.280 ;
        RECT -0.920 1.790 -0.750 1.960 ;
        RECT 1.290 1.760 1.460 1.930 ;
      LAYER met1 ;
        RECT -1.970 7.110 -1.650 7.430 ;
        RECT -23.990 6.630 -23.680 7.070 ;
        RECT -5.680 6.630 -5.370 7.070 ;
        RECT -0.990 6.860 -0.670 7.180 ;
        RECT 1.260 6.880 1.580 7.200 ;
        RECT -16.890 6.080 -16.570 6.400 ;
        RECT -1.820 6.280 -1.500 6.600 ;
        RECT -1.040 6.210 -0.720 6.530 ;
        RECT -24.150 5.670 -23.830 5.990 ;
        RECT -5.530 5.670 -5.210 5.990 ;
        RECT -2.930 5.750 -2.610 6.070 ;
        RECT -1.710 5.590 -1.500 5.700 ;
        RECT -1.730 5.270 -1.470 5.590 ;
        RECT -1.040 5.360 -0.720 5.680 ;
        RECT -25.040 4.880 -24.800 5.010 ;
        RECT -25.060 4.560 -24.800 4.880 ;
        RECT -4.560 4.880 -4.320 5.010 ;
        RECT -4.560 4.560 -4.300 4.880 ;
        RECT -2.200 4.470 -1.880 4.790 ;
        RECT -25.060 3.960 -24.800 4.280 ;
        RECT -25.040 3.840 -24.800 3.960 ;
        RECT -4.560 3.960 -4.300 4.280 ;
        RECT -1.710 3.980 -1.500 5.270 ;
        RECT -0.990 4.710 -0.670 5.030 ;
        RECT 1.310 4.660 1.630 4.980 ;
        RECT -4.560 3.840 -4.320 3.960 ;
        RECT -1.730 3.690 -1.500 3.980 ;
        RECT -0.990 3.860 -0.670 4.180 ;
        RECT 1.300 3.940 1.620 4.260 ;
        RECT -24.150 2.910 -23.830 3.230 ;
        RECT -5.530 2.910 -5.210 3.230 ;
        RECT -1.040 3.210 -0.720 3.530 ;
        RECT -16.860 2.390 -16.540 2.710 ;
        RECT -1.040 2.360 -0.720 2.680 ;
        RECT -23.990 1.780 -23.680 2.220 ;
        RECT -5.680 1.780 -5.370 2.220 ;
        RECT -0.990 1.710 -0.670 2.030 ;
        RECT 1.220 1.690 1.540 2.010 ;
      LAYER via ;
        RECT -1.940 7.140 -1.680 7.400 ;
        RECT -23.970 6.660 -23.710 6.920 ;
        RECT -5.650 6.660 -5.390 6.920 ;
        RECT -0.960 6.890 -0.700 7.150 ;
        RECT 1.290 6.910 1.550 7.170 ;
        RECT -16.860 6.110 -16.600 6.370 ;
        RECT -1.790 6.310 -1.530 6.570 ;
        RECT -1.010 6.240 -0.750 6.500 ;
        RECT -24.120 5.700 -23.860 5.960 ;
        RECT -5.500 5.700 -5.240 5.960 ;
        RECT -2.900 5.780 -2.640 6.040 ;
        RECT -1.730 5.300 -1.470 5.560 ;
        RECT -1.010 5.390 -0.750 5.650 ;
        RECT -25.060 4.590 -24.800 4.850 ;
        RECT -4.560 4.590 -4.300 4.850 ;
        RECT -2.170 4.500 -1.910 4.760 ;
        RECT -25.060 3.990 -24.800 4.250 ;
        RECT -4.560 3.990 -4.300 4.250 ;
        RECT -0.960 4.740 -0.700 5.000 ;
        RECT 1.340 4.690 1.600 4.950 ;
        RECT -0.960 3.890 -0.700 4.150 ;
        RECT 1.330 3.970 1.590 4.230 ;
        RECT -1.010 3.240 -0.750 3.500 ;
        RECT -24.120 2.940 -23.860 3.200 ;
        RECT -5.500 2.940 -5.240 3.200 ;
        RECT -16.830 2.420 -16.570 2.680 ;
        RECT -1.010 2.390 -0.750 2.650 ;
        RECT -23.970 1.930 -23.710 2.190 ;
        RECT -5.650 1.930 -5.390 2.190 ;
        RECT -0.960 1.740 -0.700 2.000 ;
        RECT 1.250 1.720 1.510 1.980 ;
      LAYER met2 ;
        RECT -0.990 7.110 -0.680 7.190 ;
        RECT 1.260 7.110 1.570 7.210 ;
        RECT -0.990 6.880 1.570 7.110 ;
        RECT -0.990 6.860 -0.680 6.880 ;
        RECT -1.810 6.570 -1.500 6.610 ;
        RECT -1.990 6.460 -1.270 6.570 ;
        RECT -1.040 6.460 -0.730 6.540 ;
        RECT -1.990 6.320 -0.730 6.460 ;
        RECT -1.810 6.280 -0.730 6.320 ;
        RECT -1.540 6.250 -0.730 6.280 ;
        RECT -1.540 6.210 -1.270 6.250 ;
        RECT -1.040 6.210 -0.730 6.250 ;
        RECT -24.140 5.930 -23.830 6.000 ;
        RECT -26.160 5.920 -23.830 5.930 ;
        RECT -5.530 5.930 -5.220 6.000 ;
        RECT -2.930 5.930 -2.620 6.070 ;
        RECT -26.160 5.710 -6.670 5.920 ;
        RECT -24.850 5.700 -6.670 5.710 ;
        RECT -24.140 5.670 -23.830 5.700 ;
        RECT -25.090 4.730 -7.850 4.950 ;
        RECT -25.090 4.590 -24.770 4.730 ;
        RECT -25.070 4.250 -24.810 4.590 ;
        RECT -25.090 3.990 -24.770 4.250 ;
        RECT -24.140 3.170 -23.830 3.240 ;
        RECT -26.160 2.960 -11.150 3.170 ;
        RECT -24.850 2.950 -11.150 2.960 ;
        RECT -24.140 2.910 -23.830 2.950 ;
        RECT -11.370 2.620 -11.150 2.950 ;
        RECT -8.070 3.120 -7.850 4.730 ;
        RECT -6.890 4.500 -6.670 5.700 ;
        RECT -5.530 5.740 -2.620 5.930 ;
        RECT -5.530 5.710 -2.930 5.740 ;
        RECT -5.530 5.670 -5.220 5.710 ;
        RECT -1.470 5.640 -1.270 5.650 ;
        RECT -1.040 5.640 -0.730 5.680 ;
        RECT -1.470 5.560 -0.730 5.640 ;
        RECT -1.760 5.540 -0.730 5.560 ;
        RECT -1.810 5.430 -0.730 5.540 ;
        RECT -1.810 5.300 -1.250 5.430 ;
        RECT -1.040 5.350 -0.730 5.430 ;
        RECT -1.810 5.290 -1.340 5.300 ;
        RECT -6.920 4.460 -6.670 4.500 ;
        RECT -6.920 3.820 -6.660 4.460 ;
        RECT -6.920 3.610 -2.790 3.820 ;
        RECT -3.000 3.470 -2.790 3.610 ;
        RECT -1.040 3.470 -0.730 3.540 ;
        RECT -3.000 3.260 -0.730 3.470 ;
        RECT -1.340 3.250 -0.730 3.260 ;
        RECT -5.530 3.170 -5.220 3.240 ;
        RECT -1.040 3.210 -0.730 3.250 ;
        RECT -5.530 3.120 -3.200 3.170 ;
        RECT -8.070 2.960 -3.200 3.120 ;
        RECT -8.070 2.900 -5.220 2.960 ;
        RECT -1.040 2.670 -0.730 2.680 ;
        RECT -7.000 2.620 -0.730 2.670 ;
        RECT -11.370 2.460 -0.730 2.620 ;
        RECT -11.370 2.400 -6.610 2.460 ;
        RECT -1.340 2.430 -0.730 2.460 ;
        RECT -1.040 2.350 -0.730 2.430 ;
        RECT -0.990 1.980 -0.680 2.030 ;
        RECT 1.220 1.980 1.530 2.020 ;
        RECT -0.990 1.750 1.720 1.980 ;
        RECT -0.990 1.700 -0.680 1.750 ;
        RECT 1.220 1.690 1.530 1.750 ;
  END
END sky130_hilas_TA2Cell_1FG

MACRO sky130_hilas_swc4x1cellOverlap
  CLASS BLOCK ;
  FOREIGN sky130_hilas_swc4x1cellOverlap ;
  ORIGIN 2.640 4.130 ;
  SIZE 10.080 BY 6.710 ;
  OBS
      LAYER nwell ;
        RECT 2.230 2.290 4.950 2.520 ;
        RECT -2.630 -3.820 -0.900 2.230 ;
        RECT 2.230 -0.570 7.440 2.290 ;
        RECT 2.220 -3.870 7.440 -0.570 ;
        RECT 2.220 -4.070 4.940 -3.870 ;
      LAYER li1 ;
        RECT 2.630 0.950 4.580 2.120 ;
        RECT 4.980 1.820 5.300 1.830 ;
        RECT 4.980 1.650 5.560 1.820 ;
        RECT 4.980 1.600 5.310 1.650 ;
        RECT 4.980 1.570 5.300 1.600 ;
        RECT 6.840 1.550 7.040 1.900 ;
        RECT 4.980 1.240 5.300 1.280 ;
        RECT 4.980 1.200 5.310 1.240 ;
        RECT 4.980 1.030 5.560 1.200 ;
        RECT 4.980 1.020 5.300 1.030 ;
        RECT 6.110 0.930 6.310 1.530 ;
        RECT 6.840 1.520 7.050 1.550 ;
        RECT 6.830 0.930 7.050 1.520 ;
        RECT 2.630 -0.580 4.580 0.590 ;
        RECT 4.980 0.390 5.300 0.400 ;
        RECT 4.980 0.220 5.560 0.390 ;
        RECT 4.980 0.180 5.310 0.220 ;
        RECT 4.980 0.140 5.300 0.180 ;
        RECT 6.110 -0.110 6.310 0.490 ;
        RECT 6.830 -0.100 7.050 0.490 ;
        RECT 6.840 -0.130 7.050 -0.100 ;
        RECT 4.980 -0.180 5.300 -0.150 ;
        RECT 4.980 -0.230 5.310 -0.180 ;
        RECT 4.980 -0.400 5.560 -0.230 ;
        RECT 4.980 -0.410 5.300 -0.400 ;
        RECT 6.840 -0.480 7.040 -0.130 ;
        RECT -2.210 -1.020 -1.660 -0.590 ;
        RECT 6.230 -0.880 6.670 -0.710 ;
        RECT 2.620 -2.140 4.570 -0.970 ;
        RECT 4.980 -1.190 5.300 -1.180 ;
        RECT 4.980 -1.360 5.560 -1.190 ;
        RECT 4.980 -1.410 5.310 -1.360 ;
        RECT 4.980 -1.440 5.300 -1.410 ;
        RECT 6.840 -1.460 7.040 -1.110 ;
        RECT 4.980 -1.770 5.300 -1.730 ;
        RECT 4.980 -1.810 5.310 -1.770 ;
        RECT 4.980 -1.980 5.560 -1.810 ;
        RECT 4.980 -1.990 5.300 -1.980 ;
        RECT 6.110 -2.080 6.310 -1.480 ;
        RECT 6.840 -1.490 7.050 -1.460 ;
        RECT 6.830 -2.080 7.050 -1.490 ;
        RECT 2.620 -3.680 4.570 -2.510 ;
        RECT 4.980 -2.610 5.300 -2.600 ;
        RECT 4.980 -2.780 5.560 -2.610 ;
        RECT 4.980 -2.820 5.310 -2.780 ;
        RECT 4.980 -2.860 5.300 -2.820 ;
        RECT 6.110 -3.110 6.310 -2.510 ;
        RECT 6.830 -3.100 7.050 -2.510 ;
        RECT 6.840 -3.130 7.050 -3.100 ;
        RECT 4.980 -3.180 5.300 -3.150 ;
        RECT 4.980 -3.230 5.310 -3.180 ;
        RECT 4.980 -3.400 5.560 -3.230 ;
        RECT 4.980 -3.410 5.300 -3.400 ;
        RECT 6.840 -3.480 7.040 -3.130 ;
      LAYER mcon ;
        RECT 3.110 1.780 3.280 1.950 ;
        RECT 3.110 1.440 3.280 1.610 ;
        RECT 5.040 1.610 5.210 1.780 ;
        RECT 6.120 1.320 6.290 1.490 ;
        RECT 3.110 1.100 3.280 1.270 ;
        RECT 5.040 1.060 5.210 1.230 ;
        RECT 6.850 1.350 7.020 1.520 ;
        RECT 3.110 0.250 3.280 0.420 ;
        RECT 5.040 0.190 5.210 0.360 ;
        RECT 3.110 -0.090 3.280 0.080 ;
        RECT 6.120 -0.070 6.290 0.100 ;
        RECT 6.850 -0.100 7.020 0.070 ;
        RECT 3.110 -0.430 3.280 -0.260 ;
        RECT 5.040 -0.360 5.210 -0.190 ;
        RECT -2.210 -0.940 -1.940 -0.670 ;
        RECT 6.490 -0.880 6.670 -0.710 ;
        RECT 3.100 -1.310 3.270 -1.140 ;
        RECT 5.040 -1.400 5.210 -1.230 ;
        RECT 3.100 -1.650 3.270 -1.480 ;
        RECT 6.120 -1.690 6.290 -1.520 ;
        RECT 3.100 -1.990 3.270 -1.820 ;
        RECT 5.040 -1.950 5.210 -1.780 ;
        RECT 6.850 -1.660 7.020 -1.490 ;
        RECT 3.100 -2.850 3.270 -2.680 ;
        RECT 5.040 -2.810 5.210 -2.640 ;
        RECT 3.100 -3.190 3.270 -3.020 ;
        RECT 6.120 -3.070 6.290 -2.900 ;
        RECT 6.850 -3.100 7.020 -2.930 ;
        RECT 3.100 -3.530 3.270 -3.360 ;
        RECT 5.040 -3.360 5.210 -3.190 ;
      LAYER met1 ;
        RECT -2.280 -3.820 -1.880 2.170 ;
        RECT 3.070 1.530 3.330 2.010 ;
        RECT 4.970 1.540 5.290 1.860 ;
        RECT 6.110 1.550 6.270 2.280 ;
        RECT 6.110 1.530 6.310 1.550 ;
        RECT 3.060 1.010 3.330 1.530 ;
        RECT 3.060 0.560 3.320 1.010 ;
        RECT 4.970 0.990 5.290 1.310 ;
        RECT 6.090 1.290 6.320 1.530 ;
        RECT 6.110 1.240 6.320 1.290 ;
        RECT 6.480 1.240 6.670 2.230 ;
        RECT 6.920 1.580 7.080 2.280 ;
        RECT 3.070 0.000 3.330 0.480 ;
        RECT 4.970 0.110 5.290 0.430 ;
        RECT 6.110 0.180 6.270 1.240 ;
        RECT 6.500 1.120 6.670 1.240 ;
        RECT 6.510 0.300 6.670 1.120 ;
        RECT 6.810 1.030 7.080 1.580 ;
        RECT 6.810 0.980 7.090 1.030 ;
        RECT 6.920 0.890 7.090 0.980 ;
        RECT 6.920 0.530 7.080 0.890 ;
        RECT 6.920 0.440 7.090 0.530 ;
        RECT 6.500 0.180 6.670 0.300 ;
        RECT 6.110 0.130 6.320 0.180 ;
        RECT 3.060 -0.520 3.330 0.000 ;
        RECT 6.090 -0.110 6.320 0.130 ;
        RECT 4.970 -0.440 5.290 -0.120 ;
        RECT 6.110 -0.130 6.310 -0.110 ;
        RECT 3.060 -0.970 3.320 -0.520 ;
        RECT 3.060 -1.560 3.320 -1.080 ;
        RECT 4.970 -1.470 5.290 -1.150 ;
        RECT 6.110 -1.460 6.270 -0.130 ;
        RECT 6.480 -0.680 6.670 0.180 ;
        RECT 6.810 0.390 7.090 0.440 ;
        RECT 6.810 -0.160 7.080 0.390 ;
        RECT 6.460 -0.910 6.700 -0.680 ;
        RECT 6.110 -1.480 6.310 -1.460 ;
        RECT 3.050 -2.080 3.320 -1.560 ;
        RECT 4.970 -2.020 5.290 -1.700 ;
        RECT 6.090 -1.720 6.320 -1.480 ;
        RECT 6.110 -1.770 6.320 -1.720 ;
        RECT 6.480 -1.770 6.670 -0.910 ;
        RECT 6.920 -1.430 7.080 -0.160 ;
        RECT 3.050 -2.530 3.310 -2.080 ;
        RECT 3.060 -3.100 3.320 -2.620 ;
        RECT 4.970 -2.890 5.290 -2.570 ;
        RECT 6.110 -2.820 6.270 -1.770 ;
        RECT 6.500 -1.890 6.670 -1.770 ;
        RECT 6.510 -2.700 6.670 -1.890 ;
        RECT 6.810 -1.980 7.080 -1.430 ;
        RECT 6.810 -2.030 7.090 -1.980 ;
        RECT 6.920 -2.120 7.090 -2.030 ;
        RECT 6.920 -2.470 7.080 -2.120 ;
        RECT 6.920 -2.560 7.090 -2.470 ;
        RECT 6.500 -2.820 6.670 -2.700 ;
        RECT 6.110 -2.870 6.320 -2.820 ;
        RECT 3.050 -3.620 3.320 -3.100 ;
        RECT 6.090 -3.110 6.320 -2.870 ;
        RECT 4.970 -3.440 5.290 -3.120 ;
        RECT 6.110 -3.130 6.310 -3.110 ;
        RECT 3.050 -4.070 3.310 -3.620 ;
        RECT 6.110 -3.860 6.270 -3.130 ;
        RECT 6.480 -3.810 6.670 -2.820 ;
        RECT 6.810 -2.610 7.090 -2.560 ;
        RECT 6.810 -3.160 7.080 -2.610 ;
        RECT 6.920 -3.860 7.080 -3.160 ;
      LAYER via ;
        RECT 5.000 1.570 5.260 1.830 ;
        RECT 5.000 1.020 5.260 1.280 ;
        RECT 5.000 0.140 5.260 0.400 ;
        RECT 5.000 -0.410 5.260 -0.150 ;
        RECT 5.000 -1.440 5.260 -1.180 ;
        RECT 5.000 -1.990 5.260 -1.730 ;
        RECT 5.000 -2.860 5.260 -2.600 ;
        RECT 5.000 -3.410 5.260 -3.150 ;
      LAYER met2 ;
        RECT 4.970 1.730 5.280 1.870 ;
        RECT -2.640 1.550 7.440 1.730 ;
        RECT 4.970 1.540 5.280 1.550 ;
        RECT 4.970 1.300 5.280 1.320 ;
        RECT -2.640 1.120 7.440 1.300 ;
        RECT 4.970 0.990 5.280 1.120 ;
        RECT 4.970 0.300 5.280 0.430 ;
        RECT -2.640 0.120 7.440 0.300 ;
        RECT 4.970 0.100 5.280 0.120 ;
        RECT 4.970 -0.130 5.280 -0.120 ;
        RECT -2.640 -0.200 4.960 -0.130 ;
        RECT 4.970 -0.200 7.440 -0.130 ;
        RECT -2.640 -0.310 7.440 -0.200 ;
        RECT 4.970 -0.450 5.280 -0.310 ;
        RECT 4.970 -1.280 5.280 -1.140 ;
        RECT 4.970 -1.290 7.440 -1.280 ;
        RECT -2.620 -1.460 7.440 -1.290 ;
        RECT 4.970 -1.470 5.280 -1.460 ;
        RECT 4.970 -1.710 5.280 -1.690 ;
        RECT -2.620 -1.880 7.440 -1.710 ;
        RECT 4.880 -1.890 7.440 -1.880 ;
        RECT 4.970 -2.020 5.280 -1.890 ;
        RECT 4.970 -2.690 5.280 -2.570 ;
        RECT -2.620 -2.700 5.280 -2.690 ;
        RECT -2.620 -2.860 7.440 -2.700 ;
        RECT -1.840 -2.950 -0.300 -2.860 ;
        RECT 4.880 -2.880 7.440 -2.860 ;
        RECT 4.970 -2.900 5.280 -2.880 ;
        RECT 4.970 -3.130 5.280 -3.120 ;
        RECT -2.620 -3.300 7.440 -3.130 ;
        RECT 4.970 -3.310 7.440 -3.300 ;
        RECT 4.970 -3.450 5.280 -3.310 ;
  END
END sky130_hilas_swc4x1cellOverlap

MACRO sky130_hilas_capacitorSize02
  CLASS BLOCK ;
  FOREIGN sky130_hilas_capacitorSize02 ;
  ORIGIN -14.140 0.480 ;
  SIZE 7.970 BY 5.830 ;
  PIN CAPTERM02
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 21.370 2.140 22.030 2.800 ;
    END
  END CAPTERM02
  PIN CAPTERM01
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 14.250 2.720 14.910 2.780 ;
        RECT 15.300 2.720 16.310 2.730 ;
        RECT 14.250 2.220 17.940 2.720 ;
        RECT 14.250 2.210 15.660 2.220 ;
        RECT 14.250 2.120 14.910 2.210 ;
        RECT 17.300 1.100 17.930 2.220 ;
        RECT 17.300 1.090 19.450 1.100 ;
        RECT 15.980 0.790 19.450 1.090 ;
        RECT 15.980 0.620 18.990 0.790 ;
    END
  END CAPTERM01
  OBS
      LAYER met2 ;
        RECT 14.140 4.800 22.110 4.980 ;
        RECT 14.140 4.370 22.110 4.550 ;
        RECT 14.170 3.370 22.110 3.550 ;
        RECT 14.170 2.940 22.110 3.120 ;
        RECT 14.380 2.600 14.750 2.660 ;
        RECT 14.160 2.320 14.750 2.600 ;
        RECT 14.380 2.260 14.750 2.320 ;
        RECT 21.500 2.620 21.870 2.680 ;
        RECT 21.500 2.340 22.110 2.620 ;
        RECT 21.500 2.280 21.870 2.340 ;
        RECT 14.170 1.790 22.110 1.960 ;
        RECT 14.170 1.370 22.110 1.540 ;
        RECT 14.170 0.390 22.110 0.560 ;
        RECT 14.170 -0.050 22.110 0.120 ;
      LAYER via2 ;
        RECT 14.430 2.320 14.710 2.600 ;
        RECT 21.550 2.340 21.830 2.620 ;
      LAYER met3 ;
        RECT 15.600 5.320 17.910 5.350 ;
        RECT 15.600 2.830 19.830 5.320 ;
        RECT 14.160 2.060 14.950 2.810 ;
        RECT 15.600 2.080 22.070 2.830 ;
        RECT 15.600 -0.460 19.830 2.080 ;
        RECT 17.880 -0.480 19.830 -0.460 ;
      LAYER via3 ;
        RECT 14.350 2.210 14.780 2.690 ;
        RECT 21.470 2.230 21.900 2.710 ;
  END
END sky130_hilas_capacitorSize02

MACRO sky130_hilas_nFETLarge
  CLASS BLOCK ;
  FOREIGN sky130_hilas_nFETLarge ;
  ORIGIN -0.640 -4.200 ;
  SIZE 4.370 BY 5.830 ;
  PIN GATE
    USE ANALOG ;
    ANTENNAGATEAREA 6.396000 ;
    PORT
      LAYER met2 ;
        RECT 0.640 4.530 1.240 5.020 ;
        RECT 0.640 4.200 1.250 4.530 ;
    END
  END GATE
  PIN SOURCE
    USE ANALOG ;
    ANTENNADIFFAREA 4.231200 ;
    PORT
      LAYER met2 ;
        RECT 0.970 9.790 4.030 9.800 ;
        RECT 0.880 9.460 4.030 9.790 ;
        RECT 0.880 7.010 1.200 9.460 ;
        RECT 3.700 9.450 4.010 9.460 ;
        RECT 0.880 6.680 4.040 7.010 ;
        RECT 0.880 5.640 1.200 6.680 ;
        RECT 0.880 5.320 4.040 5.640 ;
        RECT 1.500 5.310 1.810 5.320 ;
        RECT 2.600 5.310 2.910 5.320 ;
        RECT 3.700 5.310 4.010 5.320 ;
    END
  END SOURCE
  PIN DRAIN
    USE ANALOG ;
    ANTENNADIFFAREA 4.231200 ;
    PORT
      LAYER met2 ;
        RECT 2.060 9.080 2.370 9.110 ;
        RECT 3.150 9.080 3.460 9.090 ;
        RECT 2.060 8.780 5.010 9.080 ;
        RECT 3.150 8.760 3.460 8.780 ;
        RECT 4.260 8.740 5.010 8.780 ;
        RECT 4.630 8.610 5.010 8.740 ;
        RECT 4.660 7.740 5.010 8.610 ;
        RECT 2.060 7.410 5.010 7.740 ;
        RECT 4.660 4.970 5.010 7.410 ;
        RECT 2.070 4.960 5.010 4.970 ;
        RECT 2.060 4.650 5.010 4.960 ;
        RECT 2.060 4.640 4.780 4.650 ;
        RECT 2.060 4.630 2.370 4.640 ;
        RECT 3.150 4.630 3.460 4.640 ;
    END
  END DRAIN
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.820 6.650 1.090 6.680 ;
        RECT 0.820 6.120 1.100 6.650 ;
        RECT 0.640 5.820 1.100 6.120 ;
        RECT 0.640 5.800 1.110 5.820 ;
        RECT 0.820 5.370 1.110 5.800 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.590 9.750 1.760 9.780 ;
        RECT 1.520 9.710 1.840 9.750 ;
        RECT 1.520 9.520 1.850 9.710 ;
        RECT 1.520 9.490 1.840 9.520 ;
        RECT 1.590 6.970 1.760 9.490 ;
        RECT 2.140 9.070 2.310 9.780 ;
        RECT 2.690 9.750 2.860 9.780 ;
        RECT 2.610 9.710 2.930 9.750 ;
        RECT 2.610 9.520 2.940 9.710 ;
        RECT 2.610 9.490 2.930 9.520 ;
        RECT 2.070 9.030 2.390 9.070 ;
        RECT 2.070 8.840 2.400 9.030 ;
        RECT 2.070 8.810 2.390 8.840 ;
        RECT 2.140 7.700 2.310 8.810 ;
        RECT 2.070 7.660 2.390 7.700 ;
        RECT 2.070 7.470 2.400 7.660 ;
        RECT 2.070 7.440 2.390 7.470 ;
        RECT 1.510 6.930 1.830 6.970 ;
        RECT 1.510 6.740 1.840 6.930 ;
        RECT 1.510 6.710 1.830 6.740 ;
        RECT 0.880 5.400 1.050 6.620 ;
        RECT 1.590 5.600 1.760 6.710 ;
        RECT 1.510 5.560 1.830 5.600 ;
        RECT 1.510 5.370 1.840 5.560 ;
        RECT 1.510 5.340 1.830 5.370 ;
        RECT 0.830 4.950 1.340 5.210 ;
        RECT 0.830 4.880 1.350 4.950 ;
        RECT 0.840 4.200 1.350 4.880 ;
        RECT 1.590 4.600 1.760 5.340 ;
        RECT 2.140 4.920 2.310 7.440 ;
        RECT 2.690 6.970 2.860 9.490 ;
        RECT 3.240 9.050 3.410 9.780 ;
        RECT 3.790 9.740 3.960 9.780 ;
        RECT 3.710 9.700 4.030 9.740 ;
        RECT 3.710 9.510 4.040 9.700 ;
        RECT 3.710 9.480 4.030 9.510 ;
        RECT 3.160 9.010 3.480 9.050 ;
        RECT 3.160 8.820 3.490 9.010 ;
        RECT 3.160 8.790 3.480 8.820 ;
        RECT 3.240 7.700 3.410 8.790 ;
        RECT 3.160 7.660 3.480 7.700 ;
        RECT 3.160 7.470 3.490 7.660 ;
        RECT 3.160 7.440 3.480 7.470 ;
        RECT 2.610 6.930 2.930 6.970 ;
        RECT 2.610 6.740 2.940 6.930 ;
        RECT 2.610 6.710 2.930 6.740 ;
        RECT 2.690 5.600 2.860 6.710 ;
        RECT 2.610 5.560 2.930 5.600 ;
        RECT 2.610 5.370 2.940 5.560 ;
        RECT 2.610 5.340 2.930 5.370 ;
        RECT 2.070 4.880 2.390 4.920 ;
        RECT 2.070 4.690 2.400 4.880 ;
        RECT 2.070 4.660 2.390 4.690 ;
        RECT 2.140 4.600 2.310 4.660 ;
        RECT 2.690 4.600 2.860 5.340 ;
        RECT 3.240 4.920 3.410 7.440 ;
        RECT 3.790 6.970 3.960 9.480 ;
        RECT 4.340 9.040 4.510 9.780 ;
        RECT 4.270 9.000 4.590 9.040 ;
        RECT 4.270 8.810 4.600 9.000 ;
        RECT 4.270 8.780 4.590 8.810 ;
        RECT 4.340 7.700 4.510 8.780 ;
        RECT 4.260 7.660 4.580 7.700 ;
        RECT 4.260 7.470 4.590 7.660 ;
        RECT 4.260 7.440 4.580 7.470 ;
        RECT 3.710 6.930 4.030 6.970 ;
        RECT 3.710 6.740 4.040 6.930 ;
        RECT 3.710 6.710 4.030 6.740 ;
        RECT 3.790 5.600 3.960 6.710 ;
        RECT 3.710 5.560 4.030 5.600 ;
        RECT 3.710 5.370 4.040 5.560 ;
        RECT 3.710 5.340 4.030 5.370 ;
        RECT 3.160 4.880 3.480 4.920 ;
        RECT 3.160 4.690 3.490 4.880 ;
        RECT 3.160 4.660 3.480 4.690 ;
        RECT 3.240 4.600 3.410 4.660 ;
        RECT 3.790 4.600 3.960 5.340 ;
        RECT 4.340 4.930 4.510 7.440 ;
        RECT 4.260 4.890 4.580 4.930 ;
        RECT 4.260 4.700 4.590 4.890 ;
        RECT 4.260 4.670 4.580 4.700 ;
        RECT 4.340 4.600 4.510 4.670 ;
      LAYER mcon ;
        RECT 1.580 9.530 1.750 9.700 ;
        RECT 2.670 9.530 2.840 9.700 ;
        RECT 2.130 8.850 2.300 9.020 ;
        RECT 2.130 7.480 2.300 7.650 ;
        RECT 1.570 6.750 1.740 6.920 ;
        RECT 0.880 6.450 1.050 6.620 ;
        RECT 0.880 6.090 1.050 6.260 ;
        RECT 1.570 5.380 1.740 5.550 ;
        RECT 1.000 4.740 1.170 4.910 ;
        RECT 3.770 9.520 3.940 9.690 ;
        RECT 3.220 8.830 3.390 9.000 ;
        RECT 3.220 7.480 3.390 7.650 ;
        RECT 2.670 6.750 2.840 6.920 ;
        RECT 2.670 5.380 2.840 5.550 ;
        RECT 2.130 4.700 2.300 4.870 ;
        RECT 4.330 8.820 4.500 8.990 ;
        RECT 4.320 7.480 4.490 7.650 ;
        RECT 3.770 6.750 3.940 6.920 ;
        RECT 3.770 5.380 3.940 5.550 ;
        RECT 3.220 4.700 3.390 4.870 ;
        RECT 4.320 4.710 4.490 4.880 ;
        RECT 1.010 4.270 1.180 4.440 ;
      LAYER met1 ;
        RECT 1.510 9.460 1.830 9.780 ;
        RECT 2.600 9.460 2.920 9.780 ;
        RECT 3.700 9.450 4.020 9.770 ;
        RECT 2.060 8.780 2.380 9.100 ;
        RECT 3.150 8.760 3.470 9.080 ;
        RECT 4.260 8.750 4.580 9.070 ;
        RECT 2.060 7.410 2.380 7.730 ;
        RECT 3.150 7.410 3.470 7.730 ;
        RECT 4.250 7.410 4.570 7.730 ;
        RECT 1.500 6.680 1.820 7.000 ;
        RECT 2.600 6.680 2.920 7.000 ;
        RECT 3.700 6.680 4.020 7.000 ;
        RECT 1.500 5.310 1.820 5.630 ;
        RECT 2.600 5.310 2.920 5.630 ;
        RECT 3.700 5.310 4.020 5.630 ;
        RECT 0.930 4.670 1.250 4.990 ;
        RECT 2.060 4.630 2.380 4.950 ;
        RECT 3.150 4.630 3.470 4.950 ;
        RECT 4.250 4.640 4.570 4.960 ;
        RECT 0.940 4.200 1.260 4.520 ;
      LAYER via ;
        RECT 1.540 9.490 1.800 9.750 ;
        RECT 2.630 9.490 2.890 9.750 ;
        RECT 3.730 9.480 3.990 9.740 ;
        RECT 2.090 8.810 2.350 9.070 ;
        RECT 3.180 8.790 3.440 9.050 ;
        RECT 4.290 8.780 4.550 9.040 ;
        RECT 2.090 7.440 2.350 7.700 ;
        RECT 3.180 7.440 3.440 7.700 ;
        RECT 4.280 7.440 4.540 7.700 ;
        RECT 1.530 6.710 1.790 6.970 ;
        RECT 2.630 6.710 2.890 6.970 ;
        RECT 3.730 6.710 3.990 6.970 ;
        RECT 1.530 5.340 1.790 5.600 ;
        RECT 2.630 5.340 2.890 5.600 ;
        RECT 3.730 5.340 3.990 5.600 ;
        RECT 0.960 4.700 1.220 4.960 ;
        RECT 2.090 4.660 2.350 4.920 ;
        RECT 3.180 4.660 3.440 4.920 ;
        RECT 4.280 4.670 4.540 4.930 ;
        RECT 0.970 4.230 1.230 4.490 ;
  END
END sky130_hilas_nFETLarge

END LIBRARY