VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_Trans2med
  CLASS BLOCK ;
  FOREIGN sky130_hilas_Trans2med ;
  ORIGIN 3.800 1.430 ;
  SIZE 3.530 BY 5.950 ;
  PIN nFET_Gate01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -3.800 0.610 -3.550 0.830 ;
    END
  END nFET_Gate01
  PIN pET_Gate02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -3.800 1.590 -0.820 1.800 ;
    END
  END pET_Gate02
  PIN pFET_Gate01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -3.800 2.150 -3.550 2.370 ;
    END
  END pFET_Gate01
  PIN nFET_Gate02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -3.800 1.190 -0.820 1.400 ;
    END
  END nFET_Gate02
  PIN pFET_Source1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -3.800 3.140 -3.530 3.360 ;
    END
  END pFET_Source1
  PIN pFET_Source2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -3.800 3.920 -1.900 4.140 ;
    END
  END pFET_Source2
  PIN nFET_Source2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -3.800 -1.190 -1.880 -0.970 ;
    END
  END nFET_Source2
  PIN nFET_Source1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -3.800 -0.740 -3.100 -0.530 ;
    END
  END nFET_Source1
  PIN nFET_Drain1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -2.140 -0.720 -0.270 -0.500 ;
    END
  END nFET_Drain1
  PIN nFET_Drain2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -0.970 -1.160 -0.270 -0.950 ;
    END
  END nFET_Drain2
  PIN pFET_Drain01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -2.120 3.170 -0.270 3.380 ;
    END
  END pFET_Drain01
  PIN pFET_Drain2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT -0.930 4.000 -0.270 4.210 ;
    END
  END pFET_Drain2
  OBS
      LAYER li1 ;
        RECT -3.530 -1.250 -0.330 4.290 ;
      LAYER met1 ;
        RECT -3.550 -1.230 -0.270 4.250 ;
      LAYER met2 ;
        RECT -1.620 3.720 -1.210 4.260 ;
        RECT -1.620 3.660 -0.500 3.720 ;
        RECT -3.250 2.890 -2.400 3.640 ;
        RECT -3.250 2.860 -0.500 2.890 ;
        RECT -3.580 2.650 -0.500 2.860 ;
        RECT -3.270 2.080 -0.500 2.650 ;
        RECT -0.540 0.910 -0.500 2.080 ;
        RECT -3.270 0.330 -0.500 0.910 ;
        RECT -3.580 -0.220 -0.500 0.330 ;
        RECT -3.580 -0.250 -2.420 -0.220 ;
        RECT -2.820 -0.690 -2.420 -0.250 ;
        RECT -1.600 -1.230 -1.250 -1.000 ;
  END
END sky130_hilas_Trans2med
END LIBRARY

