magic
tech sky130A
timestamp 1608384750
<< error_s >>
rect -596 499 -590 505
rect -491 499 -485 505
rect -170 489 -164 495
rect -117 489 -111 495
rect -602 435 -596 441
rect -485 435 -479 441
rect -176 439 -170 445
rect -111 439 -105 445
rect -596 382 -590 388
rect -491 382 -485 388
rect -170 380 -164 386
rect -117 380 -111 386
rect -176 330 -170 336
rect -111 330 -105 336
rect -602 318 -596 324
rect -485 318 -479 324
rect -596 197 -590 203
rect -491 197 -485 203
rect -170 191 -164 197
rect -117 191 -111 197
rect -176 141 -170 147
rect -111 141 -105 147
rect -602 133 -596 139
rect -485 133 -479 139
rect -596 81 -590 87
rect -491 81 -485 87
rect -170 74 -164 80
rect -117 74 -111 80
rect -176 24 -170 30
rect -111 24 -105 30
rect -602 17 -596 23
rect -485 17 -479 23
<< nwell >>
rect -1101 561 -805 562
rect -1101 546 -1060 561
rect -1101 545 -1042 546
rect -1101 369 -1060 545
rect -1112 254 -1060 369
rect -1101 -42 -1060 254
<< poly >>
rect 209 516 229 562
rect 209 -43 229 -18
<< locali >>
rect -1115 -22 -1097 67
<< metal1 >>
rect -1025 561 -1009 562
rect -944 561 -928 562
rect -762 399 -740 537
rect 131 516 154 562
rect 257 516 280 562
rect -1112 254 -1091 369
rect -772 122 -745 212
rect 131 -43 154 -18
rect 257 -43 280 -18
<< metal2 >>
rect -738 530 7 531
rect -751 512 7 530
rect -1100 494 -1061 512
rect -751 510 24 512
rect -14 491 24 510
rect -1112 418 -1097 469
rect -54 457 -50 466
rect -65 437 56 457
rect 170 426 296 442
rect -1112 402 -769 418
rect -1112 352 -1086 378
rect -1107 351 -1090 352
rect -55 351 66 371
rect 170 333 296 349
rect -1100 308 -1061 326
rect -791 304 -768 305
rect -791 301 -34 304
rect -791 284 -28 301
rect -791 274 -767 284
rect -1112 256 -767 274
rect -47 264 24 284
rect -1112 254 -775 256
rect -767 234 -32 236
rect -767 214 24 234
rect -1100 193 -1061 211
rect -1118 118 -1098 168
rect -56 152 44 168
rect 170 149 296 165
rect -1118 98 -763 118
rect -1119 47 -1091 74
rect -55 54 45 71
rect 172 56 296 72
rect -55 53 39 54
rect -1100 8 -1061 26
rect -32 8 23 9
rect -790 -14 23 8
rect -790 -15 -31 -14
rect -790 -16 -713 -15
rect -790 -20 -766 -16
rect -1114 -40 -766 -20
rect -1114 -41 -847 -40
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1607089160
transform 1 0 -1102 0 1 -26
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1607089160
transform 1 0 -1107 0 1 59
box -14 -15 20 18
use sky130_hilas_m12m2  sky130_hilas_m12m2_5
timestamp 1607949437
transform 1 0 -765 0 1 103
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_4
timestamp 1607949437
transform 1 0 -767 0 1 220
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_3
timestamp 1607949437
transform 1 0 -1105 0 1 359
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1607949437
transform 1 0 -1107 0 1 258
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1607949437
transform 1 0 -751 0 1 515
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_2
timestamp 1607949437
transform 1 0 -766 0 1 409
box -9 -10 23 22
use sky130_hilas_WTA4Stage01  sky130_hilas_WTA4Stage01_0
timestamp 1607370486
transform 1 0 67 0 1 -19
box -54 1 229 535
use sky130_hilas_swc4x1BiasCell  sky130_hilas_swc4x1BiasCell_0
timestamp 1608303107
transform -1 0 -317 0 1 339
box -266 -382 745 223
<< labels >>
rlabel metal2 289 426 296 442 0 OUTPUT1
port 4 nsew analog default
rlabel metal2 291 333 296 349 0 OUTPUT2
port 5 nsew analog default
rlabel metal2 291 149 296 165 0 OUTPUT3
port 6 nsew analog default
rlabel metal2 291 56 296 72 0 OUTPUT4
port 7 nsew analog default
rlabel metal1 257 556 280 562 0 VGND
port 1 nsew ground default
rlabel poly 209 556 229 562 0 COMMONNODE
port 2 nsew analog default
rlabel metal1 131 556 154 562 0 COMMONNODE
port 2 nsew analog default
rlabel metal1 131 -43 154 -37 0 COMMONMODE
port 3 nsew analog default
rlabel poly 209 -43 229 -37 0 COMMONMODE
port 3 nsew analog default
rlabel metal1 257 -43 280 -37 0 VGND
port 1 nsew ground default
rlabel metal2 -1112 449 -1097 469 0 INPUT1
port 8 nsew analog default
rlabel metal2 -1112 352 -1086 378 0 INPUT2
port 9 nsew analog default
rlabel metal2 -1118 151 -1098 168 0 INPUT3
port 10 nsew analog default
rlabel metal2 -1119 47 -1091 74 0 INPUT4
port 11 nsew analog default
<< end >>
