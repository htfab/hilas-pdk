magic
tech sky130A
timestamp 1629137174
<< error_p >>
rect 62 62 101 65
rect 62 20 101 23
<< nwell >>
rect 0 0 161 85
<< pmos >>
rect 62 23 101 62
<< pdiff >>
rect 34 23 62 62
rect 101 23 127 62
<< poly >>
rect 0 60 26 75
rect 62 62 101 75
rect 11 15 26 60
rect 62 15 101 23
rect 11 0 151 15
<< end >>
