magic
tech sky130A
timestamp 1628616957
<< checkpaint >>
rect -92 1170 1591 1417
rect -484 952 1591 1170
rect -592 916 1591 952
rect -628 -419 1591 916
rect -484 -426 1591 -419
rect -484 -673 1199 -426
<< metal2 >>
rect 0 485 797 503
rect 0 442 797 460
rect 3 342 797 360
rect 3 299 797 317
rect 2 237 29 265
rect 766 239 797 267
rect 3 184 797 201
rect 3 142 797 159
rect 3 44 797 61
rect 3 0 797 17
<< metal3 >>
rect 568 227 766 288
rect 568 226 764 227
rect 765 226 766 227
rect 568 213 766 226
<< metal4 >>
rect 116 277 217 278
rect 45 227 380 277
rect 45 226 152 227
rect 316 115 379 227
rect 316 85 531 115
rect 349 84 531 85
use sky130_hilas_CapModule03  sky130_hilas_CapModule03_0
timestamp 1628616692
transform 1 0 538 0 1 204
box 0 0 423 583
use sky130_hilas_m22m4  sky130_hilas_m22m4_1
timestamp 1628616715
transform 1 0 750 0 1 249
box 0 0 79 75
use sky130_hilas_m22m4  sky130_hilas_m22m4_0
timestamp 1628616715
transform 1 0 38 0 1 247
box 0 0 79 75
<< labels >>
rlabel metal2 2 237 9 265 0 CAPTERM01
port 2 nsew analog default
rlabel metal2 782 239 797 267 0 CAPTERM02
port 1 nsew analog default
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
