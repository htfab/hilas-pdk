magic
tech sky130A
timestamp 1629420194
<< error_s >>
rect 2364 6133 2393 6149
rect 2443 6133 2472 6149
rect 2522 6133 2551 6149
rect 2601 6133 2630 6149
rect 2364 6099 2365 6100
rect 2392 6099 2393 6100
rect 2443 6099 2444 6100
rect 2471 6099 2472 6100
rect 2522 6099 2523 6100
rect 2550 6099 2551 6100
rect 2601 6099 2602 6100
rect 2629 6099 2630 6100
rect 2314 6070 2331 6099
rect 2363 6098 2394 6099
rect 2442 6098 2473 6099
rect 2521 6098 2552 6099
rect 2600 6098 2631 6099
rect 2364 6091 2393 6098
rect 2443 6091 2472 6098
rect 2522 6091 2551 6098
rect 2601 6091 2630 6098
rect 2364 6077 2373 6091
rect 2620 6077 2630 6091
rect 2364 6071 2393 6077
rect 2443 6071 2472 6077
rect 2522 6071 2551 6077
rect 2601 6071 2630 6077
rect 2363 6070 2394 6071
rect 2442 6070 2473 6071
rect 2521 6070 2552 6071
rect 2600 6070 2631 6071
rect 2662 6070 2680 6099
rect 2364 6069 2365 6070
rect 2392 6069 2393 6070
rect 2443 6069 2444 6070
rect 2471 6069 2472 6070
rect 2522 6069 2523 6070
rect 2550 6069 2551 6070
rect 2601 6069 2602 6070
rect 2629 6069 2630 6070
rect 2364 6020 2393 6035
rect 2443 6020 2472 6035
rect 2522 6020 2551 6035
rect 2601 6020 2630 6035
rect 2364 5853 2393 5869
rect 2443 5853 2472 5869
rect 2522 5853 2551 5869
rect 2601 5853 2630 5869
rect 2364 5819 2365 5820
rect 2392 5819 2393 5820
rect 2443 5819 2444 5820
rect 2471 5819 2472 5820
rect 2522 5819 2523 5820
rect 2550 5819 2551 5820
rect 2601 5819 2602 5820
rect 2629 5819 2630 5820
rect 2314 5790 2331 5819
rect 2363 5818 2394 5819
rect 2442 5818 2473 5819
rect 2521 5818 2552 5819
rect 2600 5818 2631 5819
rect 2364 5811 2393 5818
rect 2443 5811 2472 5818
rect 2522 5811 2551 5818
rect 2601 5811 2630 5818
rect 2364 5797 2373 5811
rect 2620 5797 2630 5811
rect 2364 5791 2393 5797
rect 2443 5791 2472 5797
rect 2522 5791 2551 5797
rect 2601 5791 2630 5797
rect 2363 5790 2394 5791
rect 2442 5790 2473 5791
rect 2521 5790 2552 5791
rect 2600 5790 2631 5791
rect 2662 5790 2680 5819
rect 2364 5789 2365 5790
rect 2392 5789 2393 5790
rect 2443 5789 2444 5790
rect 2471 5789 2472 5790
rect 2522 5789 2523 5790
rect 2550 5789 2551 5790
rect 2601 5789 2602 5790
rect 2629 5789 2630 5790
rect 3460 5771 3489 5789
rect 2364 5740 2393 5755
rect 2443 5740 2472 5755
rect 2522 5740 2551 5755
rect 2601 5740 2630 5755
rect 3460 5739 3461 5740
rect 3488 5739 3489 5740
rect 2364 5698 2393 5714
rect 2443 5698 2472 5714
rect 2522 5698 2551 5714
rect 2601 5698 2630 5714
rect 3410 5710 3428 5739
rect 3459 5738 3490 5739
rect 3460 5729 3489 5738
rect 3460 5720 3470 5729
rect 3479 5720 3489 5729
rect 3460 5711 3489 5720
rect 3459 5710 3490 5711
rect 3521 5710 3539 5739
rect 3460 5709 3461 5710
rect 3488 5709 3489 5710
rect 2364 5664 2365 5665
rect 2392 5664 2393 5665
rect 2443 5664 2444 5665
rect 2471 5664 2472 5665
rect 2522 5664 2523 5665
rect 2550 5664 2551 5665
rect 2601 5664 2602 5665
rect 2629 5664 2630 5665
rect 2314 5635 2331 5664
rect 2363 5663 2394 5664
rect 2442 5663 2473 5664
rect 2521 5663 2552 5664
rect 2600 5663 2631 5664
rect 2364 5656 2393 5663
rect 2443 5656 2472 5663
rect 2522 5656 2551 5663
rect 2601 5656 2630 5663
rect 2364 5642 2373 5656
rect 2620 5642 2630 5656
rect 2364 5636 2393 5642
rect 2443 5636 2472 5642
rect 2522 5636 2551 5642
rect 2601 5636 2630 5642
rect 2363 5635 2394 5636
rect 2442 5635 2473 5636
rect 2521 5635 2552 5636
rect 2600 5635 2631 5636
rect 2662 5635 2680 5664
rect 3460 5660 3489 5678
rect 2364 5634 2365 5635
rect 2392 5634 2393 5635
rect 2443 5634 2444 5635
rect 2471 5634 2472 5635
rect 2522 5634 2523 5635
rect 2550 5634 2551 5635
rect 2601 5634 2602 5635
rect 2629 5634 2630 5635
rect 2364 5585 2393 5600
rect 2443 5585 2472 5600
rect 2522 5585 2551 5600
rect 2601 5585 2630 5600
rect 4242 5031 4270 5037
rect 4384 5030 4412 5037
rect 4519 5031 4569 5037
rect 4842 5030 4892 5036
rect 4242 4989 4270 4995
rect 4384 4988 4412 4995
rect 4519 4989 4569 4995
rect 4842 4988 4892 4994
rect 4193 4959 4221 4965
rect 4433 4959 4461 4965
rect 4590 4959 4641 4965
rect 4771 4964 4821 4970
rect 4193 4917 4221 4923
rect 4433 4917 4461 4923
rect 4590 4917 4641 4923
rect 4771 4922 4821 4928
rect 4242 4856 4270 4862
rect 4384 4855 4412 4862
rect 4519 4856 4569 4862
rect 4842 4855 4892 4861
rect 4242 4814 4270 4820
rect 4384 4813 4412 4820
rect 4519 4814 4569 4820
rect 4842 4813 4892 4819
rect 4193 4784 4221 4790
rect 4433 4784 4461 4790
rect 4590 4784 4641 4790
rect 4771 4789 4821 4795
rect 4193 4742 4221 4748
rect 4433 4742 4461 4748
rect 4590 4742 4641 4748
rect 4771 4747 4821 4753
rect 4242 4681 4270 4687
rect 4384 4680 4412 4687
rect 4519 4681 4569 4687
rect 7585 4686 7670 4764
rect 4842 4680 4892 4686
rect 7585 4681 7586 4686
rect 5686 4653 5736 4659
rect 5758 4653 5808 4659
rect 7727 4653 7777 4659
rect 7799 4653 7849 4659
rect 8187 4657 8214 4663
rect 4242 4639 4270 4645
rect 4384 4638 4412 4645
rect 4519 4639 4569 4645
rect 4842 4638 4892 4644
rect 4193 4609 4221 4615
rect 4433 4609 4461 4615
rect 4590 4609 4641 4615
rect 4771 4614 4821 4620
rect 5686 4611 5736 4617
rect 5758 4611 5808 4617
rect 7727 4611 7777 4617
rect 7799 4611 7849 4617
rect 8187 4615 8214 4621
rect 8187 4590 8214 4596
rect 4193 4567 4221 4573
rect 4433 4567 4461 4573
rect 4590 4567 4641 4573
rect 4771 4572 4821 4578
rect 4242 4506 4270 4512
rect 4384 4505 4412 4512
rect 4519 4506 4569 4512
rect 4842 4505 4892 4511
rect 5871 4509 5874 4559
rect 5913 4509 5916 4559
rect 6007 4509 6009 4559
rect 6049 4509 6051 4559
rect 8187 4548 8214 4554
rect 8187 4507 8214 4513
rect 4242 4464 4270 4470
rect 4384 4463 4412 4470
rect 4519 4464 4569 4470
rect 4842 4463 4892 4469
rect 4193 4434 4221 4440
rect 4433 4434 4461 4440
rect 4590 4434 4641 4440
rect 4771 4439 4821 4445
rect 5871 4430 5874 4480
rect 5913 4430 5916 4480
rect 6007 4430 6009 4480
rect 6049 4430 6051 4480
rect 8187 4465 8214 4471
rect 8187 4440 8214 4446
rect 4193 4392 4221 4398
rect 4433 4392 4461 4398
rect 4590 4392 4641 4398
rect 4771 4397 4821 4403
rect 8187 4398 8214 4404
rect 10945 4400 10985 4406
rect 11095 4400 11135 4406
rect 8187 4357 8214 4363
rect 10945 4358 10985 4364
rect 11095 4358 11135 4364
rect 5096 4340 5146 4345
rect 5276 4340 5326 4346
rect 5416 4340 5466 4345
rect 4193 4331 4221 4337
rect 4433 4331 4461 4337
rect 4590 4331 4641 4337
rect 10869 4334 10909 4339
rect 11095 4332 11135 4339
rect 4771 4326 4821 4332
rect 5096 4298 5146 4303
rect 5276 4298 5326 4304
rect 5416 4298 5466 4303
rect 4193 4289 4221 4295
rect 4433 4289 4461 4295
rect 4590 4289 4641 4295
rect 4771 4284 4821 4290
rect 5096 4273 5146 4279
rect 5416 4273 5466 4279
rect 5871 4277 5874 4327
rect 5913 4277 5916 4327
rect 6007 4277 6009 4327
rect 6049 4277 6051 4327
rect 8187 4315 8214 4321
rect 8187 4290 8214 4296
rect 10869 4292 10909 4297
rect 11095 4290 11135 4297
rect 4242 4259 4270 4265
rect 4384 4259 4412 4266
rect 4519 4259 4569 4265
rect 4842 4260 4892 4266
rect 8187 4248 8214 4254
rect 5096 4231 5146 4237
rect 5416 4231 5466 4237
rect 4242 4217 4270 4223
rect 4384 4217 4412 4224
rect 4519 4217 4569 4223
rect 4842 4218 4892 4224
rect 5871 4198 5874 4248
rect 5913 4198 5916 4248
rect 6007 4198 6009 4248
rect 6049 4198 6051 4248
rect 10869 4230 10909 4235
rect 11095 4230 11135 4237
rect 8187 4207 8214 4213
rect 10869 4188 10909 4193
rect 11095 4188 11135 4195
rect 5096 4170 5146 4176
rect 5416 4170 5466 4176
rect 8187 4165 8214 4171
rect 10945 4163 10985 4169
rect 11095 4163 11135 4169
rect 4193 4156 4221 4162
rect 4433 4156 4461 4162
rect 4590 4156 4641 4162
rect 4771 4151 4821 4157
rect 5686 4140 5736 4146
rect 5758 4140 5808 4146
rect 5096 4128 5146 4134
rect 5416 4128 5466 4134
rect 4193 4114 4221 4120
rect 4433 4114 4461 4120
rect 4590 4114 4641 4120
rect 4771 4109 4821 4115
rect 5096 4104 5146 4109
rect 5276 4103 5326 4109
rect 5416 4104 5466 4109
rect 5686 4098 5736 4104
rect 5758 4098 5808 4104
rect 4242 4084 4270 4090
rect 4384 4084 4412 4091
rect 4519 4084 4569 4090
rect 4842 4085 4892 4091
rect 7585 4078 7586 4161
rect 7727 4140 7777 4146
rect 7799 4140 7849 4146
rect 8187 4140 8214 4146
rect 10945 4121 10985 4127
rect 11095 4121 11135 4127
rect 7727 4098 7777 4104
rect 7799 4098 7849 4104
rect 8187 4098 8214 4104
rect 10945 4080 10985 4086
rect 11095 4080 11135 4086
rect 5096 4062 5146 4067
rect 5276 4061 5326 4067
rect 5416 4062 5466 4067
rect 5687 4050 5737 4056
rect 5759 4050 5809 4056
rect 7727 4050 7777 4056
rect 7799 4050 7849 4056
rect 8187 4054 8214 4060
rect 4242 4042 4270 4048
rect 4384 4042 4412 4049
rect 4519 4042 4569 4048
rect 4842 4043 4892 4049
rect 10945 4038 10985 4044
rect 11095 4038 11135 4044
rect 5096 4020 5146 4025
rect 5276 4020 5326 4026
rect 5416 4020 5466 4025
rect 5687 4008 5737 4014
rect 5759 4008 5809 4014
rect 7727 4008 7777 4014
rect 7799 4008 7849 4014
rect 8187 4012 8214 4018
rect 10869 4014 10909 4019
rect 11095 4012 11135 4019
rect 8187 3987 8214 3993
rect 4193 3981 4221 3987
rect 4433 3981 4461 3987
rect 4590 3981 4641 3987
rect 4771 3976 4821 3982
rect 5096 3978 5146 3983
rect 5276 3978 5326 3984
rect 5416 3978 5466 3983
rect 10869 3972 10909 3977
rect 11095 3970 11135 3977
rect 5096 3953 5146 3959
rect 5416 3953 5466 3959
rect 8187 3945 8214 3951
rect 4193 3939 4221 3945
rect 4433 3939 4461 3945
rect 4590 3939 4641 3945
rect 4771 3934 4821 3940
rect 4242 3909 4270 3915
rect 4384 3909 4412 3916
rect 4519 3909 4569 3915
rect 4842 3910 4892 3916
rect 5096 3911 5146 3917
rect 5416 3911 5466 3917
rect 10869 3910 10909 3915
rect 11095 3910 11135 3917
rect 8187 3904 8214 3910
rect 4242 3867 4270 3873
rect 4384 3867 4412 3874
rect 4519 3867 4569 3873
rect 4842 3868 4892 3874
rect 10869 3868 10909 3873
rect 11095 3868 11135 3875
rect 8187 3862 8214 3868
rect 5096 3850 5146 3856
rect 5416 3850 5466 3856
rect 10945 3843 10985 3849
rect 11095 3843 11135 3849
rect 8187 3837 8214 3843
rect 4193 3806 4221 3812
rect 4433 3806 4461 3812
rect 4590 3806 4641 3812
rect 5096 3808 5146 3814
rect 5416 3808 5466 3814
rect 4771 3801 4821 3807
rect 10945 3801 10985 3807
rect 11095 3801 11135 3807
rect 8187 3795 8214 3801
rect 5096 3784 5146 3789
rect 5276 3783 5326 3789
rect 5416 3784 5466 3789
rect 4193 3764 4221 3770
rect 4433 3764 4461 3770
rect 4590 3764 4641 3770
rect 4771 3759 4821 3765
rect 8187 3754 8214 3760
rect 5096 3742 5146 3747
rect 5276 3741 5326 3747
rect 5416 3742 5466 3747
rect 4242 3734 4270 3740
rect 4384 3734 4412 3741
rect 4519 3734 4569 3740
rect 4842 3735 4892 3741
rect 8187 3712 8214 3718
rect 4242 3692 4270 3698
rect 4384 3692 4412 3699
rect 4519 3692 4569 3698
rect 4842 3693 4892 3699
rect 8187 3687 8214 3693
rect 8187 3645 8214 3651
rect 8187 3604 8214 3610
rect 8187 3562 8214 3568
rect 5687 3537 5737 3543
rect 5759 3537 5809 3543
rect 7727 3537 7777 3543
rect 7799 3537 7849 3543
rect 8187 3537 8214 3543
rect 5687 3495 5737 3501
rect 5759 3495 5809 3501
rect 7727 3495 7777 3501
rect 7799 3495 7849 3501
rect 8187 3495 8214 3501
rect 4193 3318 4221 3324
rect 4433 3318 4461 3324
rect 4590 3318 4641 3324
rect 4771 3313 4821 3319
rect 5094 3293 5144 3298
rect 5274 3293 5324 3299
rect 5414 3293 5464 3298
rect 5828 3292 5878 3298
rect 5900 3292 5950 3298
rect 7584 3292 7634 3298
rect 7656 3292 7706 3298
rect 4193 3276 4221 3282
rect 4433 3276 4461 3282
rect 4590 3276 4641 3282
rect 4771 3271 4821 3277
rect 4242 3246 4270 3252
rect 4384 3246 4412 3253
rect 4519 3246 4569 3252
rect 4842 3247 4892 3253
rect 5094 3251 5144 3256
rect 5274 3251 5324 3257
rect 5414 3251 5464 3256
rect 5828 3250 5878 3256
rect 5900 3250 5950 3256
rect 7584 3250 7634 3256
rect 7656 3250 7706 3256
rect 5094 3226 5144 3232
rect 5414 3226 5464 3232
rect 5900 3223 5950 3229
rect 7584 3223 7634 3229
rect 4242 3204 4270 3210
rect 4384 3204 4412 3211
rect 4519 3204 4569 3210
rect 4842 3205 4892 3211
rect 5094 3184 5144 3190
rect 5414 3184 5464 3190
rect 5900 3181 5950 3187
rect 7584 3181 7634 3187
rect 4193 3143 4221 3149
rect 4433 3143 4461 3149
rect 4590 3143 4641 3149
rect 4771 3138 4821 3144
rect 5900 3138 5950 3144
rect 7584 3138 7634 3144
rect 5094 3123 5144 3129
rect 5414 3123 5464 3129
rect 4193 3101 4221 3107
rect 4433 3101 4461 3107
rect 4590 3101 4641 3107
rect 4771 3096 4821 3102
rect 5900 3096 5950 3102
rect 7584 3096 7634 3102
rect 5094 3081 5144 3087
rect 5414 3081 5464 3087
rect 4242 3071 4270 3077
rect 4384 3071 4412 3078
rect 4519 3071 4569 3077
rect 4842 3072 4892 3078
rect 5828 3069 5878 3075
rect 5900 3069 5950 3075
rect 7584 3069 7634 3075
rect 7656 3069 7706 3075
rect 5094 3057 5144 3062
rect 5274 3056 5324 3062
rect 5414 3057 5464 3062
rect 4242 3029 4270 3035
rect 4384 3029 4412 3036
rect 4519 3029 4569 3035
rect 4842 3030 4892 3036
rect 5828 3027 5878 3033
rect 5900 3027 5950 3033
rect 7584 3027 7634 3033
rect 7656 3027 7706 3033
rect 5094 3015 5144 3020
rect 5274 3014 5324 3020
rect 5414 3015 5464 3020
rect 4193 2968 4221 2974
rect 4433 2968 4461 2974
rect 4590 2968 4641 2974
rect 5094 2973 5144 2978
rect 5274 2973 5324 2979
rect 5414 2973 5464 2978
rect 4771 2963 4821 2969
rect 5828 2968 5878 2974
rect 5900 2968 5950 2974
rect 7584 2968 7634 2974
rect 7656 2968 7706 2974
rect 4193 2926 4221 2932
rect 4433 2926 4461 2932
rect 4590 2926 4641 2932
rect 5094 2931 5144 2936
rect 5274 2931 5324 2937
rect 5414 2931 5464 2936
rect 4771 2921 4821 2927
rect 5828 2926 5878 2932
rect 5900 2926 5950 2932
rect 7584 2926 7634 2932
rect 7656 2926 7706 2932
rect 5094 2906 5144 2912
rect 5414 2906 5464 2912
rect 4242 2896 4270 2902
rect 4384 2896 4412 2903
rect 4519 2896 4569 2902
rect 4842 2897 4892 2903
rect 5900 2899 5950 2905
rect 7584 2899 7634 2905
rect 5094 2864 5144 2870
rect 5414 2864 5464 2870
rect 4242 2854 4270 2860
rect 4384 2854 4412 2861
rect 4519 2854 4569 2860
rect 4842 2855 4892 2861
rect 5900 2857 5950 2863
rect 7584 2857 7634 2863
rect 5900 2815 5950 2821
rect 7584 2815 7634 2821
rect 5094 2803 5144 2809
rect 5414 2803 5464 2809
rect 4193 2793 4221 2799
rect 4433 2793 4461 2799
rect 4590 2793 4641 2799
rect 4771 2788 4821 2794
rect 5900 2773 5950 2779
rect 7584 2773 7634 2779
rect 5094 2761 5144 2767
rect 5414 2761 5464 2767
rect 4193 2751 4221 2757
rect 4433 2751 4461 2757
rect 4590 2751 4641 2757
rect 4771 2746 4821 2752
rect 5828 2746 5878 2752
rect 5900 2746 5950 2752
rect 7584 2746 7634 2752
rect 7656 2746 7706 2752
rect 5094 2737 5144 2742
rect 5274 2736 5324 2742
rect 5414 2737 5464 2742
rect 4242 2721 4270 2727
rect 4384 2721 4412 2728
rect 4519 2721 4569 2727
rect 4842 2722 4892 2728
rect 5828 2704 5878 2710
rect 5900 2704 5950 2710
rect 7584 2704 7634 2710
rect 7656 2704 7706 2710
rect 5094 2695 5144 2700
rect 5274 2694 5324 2700
rect 5414 2695 5464 2700
rect 4242 2679 4270 2685
rect 4384 2679 4412 2686
rect 4519 2679 4569 2685
rect 4842 2680 4892 2686
rect 4189 2412 4217 2418
rect 4429 2412 4457 2418
rect 4586 2412 4637 2418
rect 4767 2407 4817 2413
rect 4189 2370 4217 2376
rect 4429 2370 4457 2376
rect 4586 2370 4637 2376
rect 4767 2365 4817 2371
rect 5097 2366 5147 2371
rect 5277 2366 5327 2372
rect 5417 2366 5467 2371
rect 5831 2359 5881 2365
rect 5903 2359 5953 2365
rect 4238 2340 4266 2346
rect 4380 2340 4408 2347
rect 4515 2340 4565 2346
rect 4838 2341 4888 2347
rect 5097 2324 5147 2329
rect 5277 2324 5327 2330
rect 5417 2324 5467 2329
rect 5831 2317 5881 2323
rect 5903 2317 5953 2323
rect 4238 2298 4266 2304
rect 4380 2298 4408 2305
rect 4515 2298 4565 2304
rect 4838 2299 4888 2305
rect 5097 2299 5147 2305
rect 5417 2299 5467 2305
rect 5903 2290 5953 2296
rect 5097 2257 5147 2263
rect 5417 2257 5467 2263
rect 5903 2248 5953 2254
rect 4189 2237 4217 2243
rect 4429 2237 4457 2243
rect 4586 2237 4637 2243
rect 4767 2232 4817 2238
rect 5903 2207 5953 2213
rect 4189 2195 4217 2201
rect 4429 2195 4457 2201
rect 4586 2195 4637 2201
rect 5097 2196 5147 2202
rect 5417 2196 5467 2202
rect 4767 2190 4817 2196
rect 4238 2165 4266 2171
rect 4380 2165 4408 2172
rect 4515 2165 4565 2171
rect 4838 2166 4888 2172
rect 5903 2165 5953 2171
rect 5097 2154 5147 2160
rect 5417 2154 5467 2160
rect 5831 2138 5881 2144
rect 5903 2138 5953 2144
rect 5097 2130 5147 2135
rect 4238 2123 4266 2129
rect 4380 2123 4408 2130
rect 4515 2123 4565 2129
rect 4838 2124 4888 2130
rect 5277 2129 5327 2135
rect 5417 2130 5467 2135
rect 5831 2096 5881 2102
rect 5903 2096 5953 2102
rect 5097 2088 5147 2093
rect 5277 2087 5327 2093
rect 5417 2088 5467 2093
rect 4189 2062 4217 2068
rect 4429 2062 4457 2068
rect 4586 2062 4637 2068
rect 4767 2057 4817 2063
rect 5097 2046 5147 2051
rect 5277 2046 5327 2052
rect 5417 2046 5467 2051
rect 5831 2035 5881 2041
rect 5903 2035 5953 2041
rect 4189 2020 4217 2026
rect 4429 2020 4457 2026
rect 4586 2020 4637 2026
rect 4767 2015 4817 2021
rect 5097 2004 5147 2009
rect 5277 2004 5327 2010
rect 5417 2004 5467 2009
rect 4238 1990 4266 1996
rect 4380 1990 4408 1997
rect 4515 1990 4565 1996
rect 4838 1991 4888 1997
rect 5831 1993 5881 1999
rect 5903 1993 5953 1999
rect 5097 1979 5147 1985
rect 5417 1979 5467 1985
rect 5903 1966 5953 1972
rect 4238 1948 4266 1954
rect 4380 1948 4408 1955
rect 4515 1948 4565 1954
rect 4838 1949 4888 1955
rect 5097 1937 5147 1943
rect 5417 1937 5467 1943
rect 5903 1924 5953 1930
rect 4189 1887 4217 1893
rect 4429 1887 4457 1893
rect 4586 1887 4637 1893
rect 4767 1882 4817 1888
rect 5903 1882 5953 1888
rect 5097 1876 5147 1882
rect 5417 1876 5467 1882
rect 4189 1845 4217 1851
rect 4429 1845 4457 1851
rect 4586 1845 4637 1851
rect 4767 1840 4817 1846
rect 5903 1840 5953 1846
rect 5097 1834 5147 1840
rect 5417 1834 5467 1840
rect 4238 1815 4266 1821
rect 4380 1815 4408 1822
rect 4515 1815 4565 1821
rect 4838 1816 4888 1822
rect 5097 1810 5147 1815
rect 5277 1809 5327 1815
rect 5417 1810 5467 1815
rect 5831 1813 5881 1819
rect 5903 1813 5953 1819
rect 4238 1773 4266 1779
rect 4380 1773 4408 1780
rect 4515 1773 4565 1779
rect 4838 1774 4888 1780
rect 5097 1768 5147 1773
rect 5277 1767 5327 1773
rect 5417 1768 5467 1773
rect 5831 1771 5881 1777
rect 5903 1771 5953 1777
rect 10459 899 10462 938
rect 10501 899 10504 938
rect 10555 899 10558 938
rect 10597 899 10600 938
rect 10651 899 10654 938
rect 10693 899 10696 938
rect 10747 899 10750 938
rect 10789 899 10792 938
rect 10843 899 10846 938
rect 10885 899 10888 938
rect 10939 899 10942 938
rect 10981 899 10984 938
rect 10459 738 10462 777
rect 10501 738 10504 777
rect 10555 737 10558 776
rect 10597 737 10600 776
rect 10651 737 10654 776
rect 10693 737 10696 776
rect 10747 737 10750 776
rect 10789 737 10792 776
rect 10843 737 10846 776
rect 10885 737 10888 776
rect 10939 738 10942 777
rect 10981 738 10984 777
rect 10459 577 10462 616
rect 10501 577 10504 616
rect 10555 576 10558 615
rect 10597 576 10600 615
rect 10651 576 10654 615
rect 10693 576 10696 615
rect 10747 576 10750 615
rect 10789 576 10792 615
rect 10843 576 10846 615
rect 10885 576 10888 615
rect 10939 577 10942 616
rect 10981 577 10984 616
rect 10459 416 10462 455
rect 10501 416 10504 455
rect 10555 415 10558 454
rect 10597 415 10600 454
rect 10651 415 10654 454
rect 10693 415 10696 454
rect 10747 415 10750 454
rect 10789 415 10792 454
rect 10843 415 10846 454
rect 10885 415 10888 454
rect 10939 416 10942 455
rect 10981 416 10984 455
rect 10459 255 10462 294
rect 10501 255 10504 294
rect 10555 254 10558 293
rect 10597 254 10600 293
rect 10651 254 10654 293
rect 10693 254 10696 293
rect 10747 254 10750 293
rect 10789 254 10792 293
rect 10843 254 10846 293
rect 10885 254 10888 293
rect 10939 255 10942 294
rect 10981 255 10984 294
rect 10727 204 10731 205
rect 10459 94 10462 133
rect 10501 94 10504 133
rect 10555 93 10558 132
rect 10597 93 10600 132
rect 10651 93 10654 132
rect 10693 93 10696 132
rect 10747 93 10750 132
rect 10789 93 10792 132
rect 10843 93 10846 132
rect 10885 93 10888 132
rect 10939 94 10942 133
rect 10981 94 10984 133
rect 10459 -67 10462 -28
rect 10501 -67 10504 -28
rect 10555 -68 10558 -29
rect 10597 -68 10600 -29
rect 10651 -68 10654 -29
rect 10693 -68 10696 -29
rect 10747 -68 10750 -29
rect 10789 -68 10792 -29
rect 10843 -68 10846 -29
rect 10885 -68 10888 -29
rect 10939 -67 10942 -28
rect 10981 -67 10984 -28
rect 10459 -228 10462 -189
rect 10501 -228 10504 -189
rect 10555 -229 10558 -190
rect 10597 -229 10600 -190
rect 10651 -229 10654 -190
rect 10693 -229 10696 -190
rect 10747 -229 10750 -190
rect 10789 -229 10792 -190
rect 10843 -229 10846 -190
rect 10885 -229 10888 -190
rect 10939 -228 10942 -189
rect 10981 -228 10984 -189
rect 10459 -389 10462 -350
rect 10501 -389 10504 -350
rect 10555 -390 10558 -351
rect 10597 -390 10600 -351
rect 10651 -390 10654 -351
rect 10693 -390 10696 -351
rect 10747 -390 10750 -351
rect 10789 -390 10792 -351
rect 10843 -390 10846 -351
rect 10885 -390 10888 -351
rect 10939 -389 10942 -350
rect 10981 -389 10984 -350
rect 10459 -550 10462 -511
rect 10501 -550 10504 -511
rect 10555 -550 10558 -511
rect 10597 -550 10600 -511
rect 10651 -550 10654 -511
rect 10693 -550 10696 -511
rect 10747 -550 10750 -511
rect 10789 -550 10792 -511
rect 10843 -550 10846 -511
rect 10885 -550 10888 -511
rect 10939 -550 10942 -511
rect 10981 -550 10984 -511
<< nwell >>
rect 5619 4373 5622 4374
rect 4143 4359 4320 4370
rect 4707 4359 4957 4370
rect 5551 4343 5622 4373
rect 5551 4339 5619 4343
rect 5550 3734 5620 4339
rect 6597 4130 6598 4249
rect 6597 4125 6602 4130
rect 6597 4115 6603 4125
rect 6598 4003 6603 4115
rect 7940 4024 7996 4078
rect 5551 3714 5620 3734
rect 5550 1762 5725 2359
rect 5550 1759 5852 1762
rect 5764 1743 5852 1759
rect 5740 1046 5942 1615
rect 11004 -566 11139 981
rect 11003 -613 11139 -566
<< psubdiff >>
rect 886 5216 2688 5229
rect 886 5145 2258 5216
rect 2347 5145 2688 5216
rect 886 5138 2688 5145
rect 2597 1408 2688 5138
rect 6992 4911 8603 4916
rect 6992 4829 7005 4911
rect 7031 4910 8603 4911
rect 7031 4832 8338 4910
rect 8427 4832 8603 4910
rect 7031 4829 8603 4832
rect 6992 4825 8603 4829
rect 8512 3006 8603 4825
rect 2597 1374 2608 1408
rect 2625 1391 2642 1408
rect 2659 1391 2688 1408
rect 2676 1374 2688 1391
rect 2597 1356 2688 1374
rect 2597 1295 2611 1356
rect 2664 1295 2688 1356
rect 2031 529 2282 538
rect 2031 487 2059 529
rect 2032 177 2059 487
rect 2076 177 2095 529
rect 2112 177 2130 529
rect 2147 177 2165 529
rect 2182 177 2201 529
rect 2218 177 2236 529
rect 2253 177 2282 529
rect 2032 164 2282 177
rect 2597 245 2688 1295
rect 8263 2915 8603 3006
rect 8263 245 8354 2915
rect 2032 163 2067 164
rect 2597 154 9755 245
rect 2597 -243 2688 154
<< nsubdiff >>
rect 11045 950 11102 958
rect 11045 556 11058 950
rect 11049 496 11058 556
rect 11045 395 11058 496
rect 11049 335 11058 395
rect 11045 234 11058 335
rect 11048 174 11058 234
rect 11045 72 11058 174
rect 11049 12 11058 72
rect 11045 -89 11058 12
rect 11048 -149 11058 -89
rect 11045 -336 11058 -149
rect 11048 -545 11058 -336
rect 11075 -545 11102 950
rect 11048 -557 11102 -545
<< psubdiffcont >>
rect 2258 5145 2347 5216
rect 7005 4829 7031 4911
rect 8338 4832 8427 4910
rect 2608 1391 2625 1408
rect 2642 1391 2659 1408
rect 2608 1374 2676 1391
rect 2611 1295 2664 1356
rect 2059 177 2076 529
rect 2095 177 2112 529
rect 2130 177 2147 529
rect 2165 177 2182 529
rect 2201 177 2218 529
rect 2236 177 2253 529
<< nsubdiffcont >>
rect 11058 -545 11075 950
<< locali >>
rect 2200 5221 2352 5222
rect 2200 5219 2355 5221
rect 2200 5145 2207 5219
rect 2250 5216 2355 5219
rect 2250 5145 2258 5216
rect 2347 5145 2355 5216
rect 2200 5142 2355 5145
rect 6997 4911 7064 4913
rect 6997 4829 7005 4911
rect 7031 4829 7036 4911
rect 7062 4829 7064 4911
rect 6997 4826 7064 4829
rect 8225 4911 8435 4913
rect 8225 4832 8231 4911
rect 8263 4910 8435 4911
rect 8263 4832 8338 4910
rect 8427 4832 8435 4910
rect 8225 4828 8435 4832
rect 2600 1374 2608 1408
rect 2639 1391 2642 1408
rect 2600 1366 2676 1374
rect 2602 1356 2676 1366
rect 2602 1295 2611 1356
rect 2664 1295 2676 1356
rect 2602 1287 2676 1295
rect 11058 951 11095 958
rect 11058 950 11078 951
rect 2035 529 2274 534
rect 2035 497 2041 529
rect 2040 177 2041 497
rect 2058 177 2059 529
rect 2076 177 2077 529
rect 2094 177 2095 529
rect 2112 177 2113 529
rect 2147 177 2165 529
rect 2199 177 2201 529
rect 2235 177 2236 529
rect 2253 177 2254 529
rect 2271 177 2274 529
rect 2040 171 2274 177
rect 2040 170 2273 171
rect 11075 -544 11078 950
rect 11095 -544 11096 -529
rect 11075 -545 11096 -544
rect 11058 -554 11096 -545
<< viali >>
rect 2207 5145 2250 5219
rect 7036 4829 7062 4911
rect 8231 4832 8263 4911
rect 2622 1391 2625 1408
rect 2625 1391 2639 1408
rect 2659 1391 2676 1408
rect 2622 1374 2639 1391
rect 2659 1374 2676 1391
rect 2041 177 2058 529
rect 2077 177 2094 529
rect 2113 177 2130 529
rect 2182 177 2199 529
rect 2218 177 2235 529
rect 2254 177 2271 529
rect 11078 -544 11095 951
<< metal1 >>
rect 8233 6611 8267 6625
rect 9021 6611 9093 6785
rect 8233 6539 9093 6611
rect 3026 6294 3160 6339
rect 416 6254 466 6258
rect 416 6215 421 6254
rect 460 6215 466 6254
rect 3026 6252 4378 6294
rect 4557 6285 4876 6397
rect 3026 6238 3160 6252
rect 416 6210 466 6215
rect 426 5914 465 6210
rect 2485 6178 2762 6202
rect 2485 6137 2509 6178
rect 426 5909 473 5914
rect 426 5870 429 5909
rect 468 5870 473 5909
rect 426 5865 473 5870
rect 426 5864 471 5865
rect 426 53 465 5864
rect 567 5779 593 5782
rect 567 5750 593 5753
rect 568 5528 592 5750
rect 559 5525 601 5528
rect 559 5480 601 5483
rect 1148 5404 1177 5596
rect 1146 5401 1187 5404
rect 1146 5343 1154 5401
rect 1183 5343 1187 5401
rect 1146 5337 1187 5343
rect 2484 5268 2508 5591
rect 2479 5263 2513 5268
rect 2479 5237 2483 5263
rect 2509 5237 2513 5263
rect 2479 5234 2513 5237
rect 2204 5224 2253 5225
rect 2203 5219 2254 5224
rect 2203 5145 2207 5219
rect 2250 5145 2254 5219
rect 1811 4355 1834 4703
rect 1878 4641 1900 4703
rect 2147 4675 2169 5130
rect 2203 5109 2254 5145
rect 2738 5131 2762 6178
rect 3069 6145 3372 6172
rect 3540 6146 3566 6252
rect 3066 5228 3097 5598
rect 3058 5225 3097 5228
rect 3058 5194 3062 5225
rect 3093 5194 3097 5225
rect 3058 5191 3097 5194
rect 3345 5177 3372 6145
rect 4336 5927 4378 6252
rect 4717 6003 4759 6285
rect 4717 6000 4764 6003
rect 4717 5958 4720 6000
rect 4762 5958 4764 6000
rect 4717 5955 4764 5958
rect 4332 5924 4380 5927
rect 4332 5882 4335 5924
rect 4377 5882 4380 5924
rect 4332 5879 4380 5882
rect 4887 5765 4931 5768
rect 4887 5718 4931 5721
rect 5459 5765 5503 5768
rect 5459 5718 5503 5721
rect 5638 5762 5711 6401
rect 6153 6386 6251 6401
rect 5638 5718 5641 5762
rect 5685 5718 5711 5762
rect 4445 5663 4489 5666
rect 4445 5616 4489 5619
rect 3462 5277 3487 5592
rect 4166 5343 4198 5347
rect 4166 5342 4169 5343
rect 4157 5317 4169 5342
rect 4195 5317 4198 5343
rect 4157 5313 4198 5317
rect 3458 5274 3491 5277
rect 3458 5248 3462 5274
rect 3488 5248 3491 5274
rect 3458 5241 3491 5248
rect 3341 5175 3375 5177
rect 3341 5149 3345 5175
rect 3372 5149 3375 5175
rect 3341 5146 3375 5149
rect 2198 5106 2254 5109
rect 2198 5099 2212 5106
rect 2187 5071 2212 5099
rect 2247 5071 2254 5106
rect 2733 5128 2767 5131
rect 2733 5102 2737 5128
rect 2763 5102 2767 5128
rect 2733 5099 2767 5102
rect 2187 5059 2254 5071
rect 2187 5056 2253 5059
rect 2187 4675 2209 5056
rect 4157 4963 4181 5313
rect 4451 4956 4482 5616
rect 4894 4958 4923 5718
rect 5013 5619 5016 5663
rect 5060 5619 5063 5663
rect 2309 4886 2344 4890
rect 2309 4847 2314 4886
rect 2340 4847 2344 4886
rect 2309 4844 2344 4847
rect 3952 4874 3989 4877
rect 3952 4848 3954 4874
rect 3987 4848 3989 4874
rect 3952 4846 3989 4848
rect 2249 4808 2274 4820
rect 2246 4805 2278 4808
rect 2246 4765 2250 4805
rect 2276 4765 2278 4805
rect 2246 4762 2278 4765
rect 2249 4683 2274 4762
rect 2249 4680 2278 4683
rect 2249 4654 2252 4680
rect 2249 4651 2278 4654
rect 1875 4638 1901 4641
rect 1875 4609 1901 4612
rect 1878 4549 1900 4609
rect 1872 4546 1900 4549
rect 1898 4520 1900 4546
rect 1872 4517 1900 4520
rect 1878 4457 1900 4517
rect 1873 4454 1900 4457
rect 1899 4428 1900 4454
rect 1873 4425 1900 4428
rect 1808 4352 1834 4355
rect 1808 4323 1834 4326
rect 1811 4259 1834 4323
rect 1804 4256 1834 4259
rect 1830 4230 1834 4256
rect 1804 4227 1834 4230
rect 1811 4163 1834 4227
rect 1808 4160 1834 4163
rect 1808 4131 1834 4134
rect 1811 2656 1834 4131
rect 1878 2656 1900 4425
rect 2249 4591 2274 4651
rect 2249 4588 2278 4591
rect 2249 4562 2252 4588
rect 2249 4559 2278 4562
rect 2249 4499 2274 4559
rect 2249 4496 2275 4499
rect 2249 4467 2275 4470
rect 1800 2653 1834 2656
rect 1800 2606 1804 2653
rect 1830 2606 1834 2653
rect 1800 2603 1834 2606
rect 1866 2653 1900 2656
rect 1866 2606 1868 2653
rect 1894 2606 1900 2653
rect 1866 2603 1900 2606
rect 1669 2529 1692 2536
rect 1665 2503 1668 2529
rect 1694 2503 1697 2529
rect 1620 2492 1643 2496
rect 1616 2489 1643 2492
rect 1642 2463 1643 2489
rect 1616 2460 1643 2463
rect 685 2404 757 2406
rect 685 2338 688 2404
rect 754 2338 757 2404
rect 685 2336 757 2338
rect 686 1821 752 2336
rect 1620 2108 1643 2460
rect 1669 2256 1692 2503
rect 1811 2494 1834 2603
rect 1878 2530 1900 2603
rect 2054 2532 2081 2536
rect 1876 2527 1902 2530
rect 1876 2498 1902 2501
rect 2052 2529 2081 2532
rect 2079 2502 2081 2529
rect 2052 2499 2081 2502
rect 1810 2491 1836 2494
rect 1810 2462 1836 2465
rect 1999 2345 2028 2348
rect 1669 2219 1742 2256
rect 1620 2101 1646 2108
rect 1618 2100 1646 2101
rect 1615 2098 1647 2100
rect 1615 2072 1618 2098
rect 1644 2072 1647 2098
rect 1615 2069 1647 2072
rect 1205 1923 1248 1926
rect 1205 1886 1209 1923
rect 1246 1886 1248 1923
rect 1205 1883 1248 1886
rect 686 1818 760 1821
rect 686 1752 692 1818
rect 758 1752 760 1818
rect 686 1749 760 1752
rect 1210 1302 1247 1883
rect 1669 1469 1692 2219
rect 2054 2202 2081 2499
rect 2042 2177 2081 2202
rect 2102 2492 2126 2496
rect 2102 2489 2128 2492
rect 2102 2460 2128 2463
rect 2102 2146 2126 2460
rect 2042 2123 2126 2146
rect 1669 1446 1914 1469
rect 1882 1413 1914 1446
rect 1206 1299 1249 1302
rect 1206 1262 1208 1299
rect 1245 1262 1249 1299
rect 1206 1259 1249 1262
rect 1958 1256 1991 1259
rect 1944 1248 1962 1256
rect 1920 1224 1962 1248
rect 1958 1220 1962 1224
rect 1988 1220 1991 1256
rect 1958 1217 1991 1220
rect 1507 725 1536 728
rect 1507 693 1536 696
rect 1508 636 1534 693
rect 2102 657 2126 2123
rect 2147 2056 2169 4131
rect 2187 2317 2209 4131
rect 2249 2432 2274 4467
rect 2311 4390 2337 4844
rect 3888 4709 3927 4711
rect 3888 4676 3891 4709
rect 3924 4676 3927 4709
rect 3888 4674 3927 4676
rect 3830 4561 3869 4564
rect 3830 4528 3834 4561
rect 3867 4528 3869 4561
rect 3830 4525 3869 4528
rect 3766 4401 3805 4404
rect 2311 4387 2339 4390
rect 2311 4361 2313 4387
rect 3766 4368 3770 4401
rect 3803 4368 3805 4401
rect 3766 4366 3805 4368
rect 2311 4358 2339 4361
rect 3769 4365 3803 4366
rect 2311 4294 2337 4358
rect 3705 4346 3739 4347
rect 3704 4344 3740 4346
rect 3704 4311 3706 4344
rect 3739 4311 3740 4344
rect 3704 4307 3740 4311
rect 2311 4291 2340 4294
rect 2311 4265 2314 4291
rect 2311 4262 2340 4265
rect 2311 4198 2337 4262
rect 2311 4195 2339 4198
rect 2311 4169 2313 4195
rect 2311 4166 2339 4169
rect 3643 4187 3679 4190
rect 2249 2430 2275 2432
rect 2248 2429 2276 2430
rect 2248 2403 2249 2429
rect 2275 2403 2276 2429
rect 2248 2402 2276 2403
rect 2249 2400 2275 2402
rect 2183 2314 2215 2317
rect 2183 2288 2187 2314
rect 2213 2288 2215 2314
rect 2183 2285 2215 2288
rect 2143 2053 2171 2056
rect 2143 2027 2145 2053
rect 2143 2024 2171 2027
rect 2147 727 2169 2024
rect 2187 1503 2209 2285
rect 2187 1500 2216 1503
rect 2187 1458 2189 1500
rect 2215 1458 2216 1500
rect 2187 1455 2216 1458
rect 2187 1259 2209 1455
rect 2185 1256 2211 1259
rect 2185 1217 2211 1220
rect 2187 755 2209 1217
rect 2249 893 2274 2400
rect 2311 1999 2337 4166
rect 3643 4154 3645 4187
rect 3678 4154 3679 4187
rect 3643 4151 3679 4154
rect 3578 4034 3619 4037
rect 3578 4001 3582 4034
rect 3615 4001 3619 4034
rect 3578 3997 3619 4001
rect 3525 3877 3561 3880
rect 3525 3844 3526 3877
rect 3559 3844 3561 3877
rect 3525 3841 3561 3844
rect 3467 3335 3500 3337
rect 3461 3330 3500 3335
rect 3461 3297 3464 3330
rect 3497 3297 3500 3330
rect 3461 3293 3500 3297
rect 3404 3174 3437 3176
rect 3399 3171 3438 3174
rect 3399 3138 3401 3171
rect 3434 3138 3438 3171
rect 3399 3135 3438 3138
rect 3342 3019 3375 3020
rect 3339 3016 3375 3019
rect 3372 2983 3375 3016
rect 3339 2980 3375 2983
rect 3277 2868 3316 2872
rect 3277 2835 3279 2868
rect 3312 2835 3316 2868
rect 3277 2832 3316 2835
rect 3210 2351 3253 2355
rect 3210 2318 3215 2351
rect 3248 2318 3253 2351
rect 3210 2315 3253 2318
rect 3144 2194 3185 2198
rect 3144 2161 3148 2194
rect 3181 2161 3185 2194
rect 3144 2158 3185 2161
rect 3083 2030 3122 2034
rect 2310 1996 2341 1999
rect 2310 1970 2313 1996
rect 2339 1970 2341 1996
rect 3083 1997 3086 2030
rect 3119 1997 3122 2030
rect 3083 1994 3122 1997
rect 2310 1967 2341 1970
rect 2245 890 2275 893
rect 2245 857 2247 890
rect 2273 857 2275 890
rect 2245 853 2275 857
rect 2187 741 2211 755
rect 2143 724 2174 727
rect 2143 695 2144 724
rect 2173 695 2174 724
rect 2143 692 2174 695
rect 2188 678 2211 741
rect 2023 654 2126 657
rect 2023 594 2028 654
rect 2088 601 2126 654
rect 2187 675 2211 678
rect 2088 594 2102 601
rect 2023 590 2102 594
rect 2187 536 2209 675
rect 2034 529 2276 536
rect 2034 177 2041 529
rect 2058 177 2077 529
rect 2094 177 2113 529
rect 2130 177 2182 529
rect 2199 177 2218 529
rect 2235 177 2254 529
rect 2271 177 2276 529
rect 2034 168 2276 177
rect 2311 139 2337 1967
rect 3014 1886 3055 1889
rect 3014 1853 3018 1886
rect 3051 1853 3055 1886
rect 3014 1850 3055 1853
rect 2593 1488 2686 1500
rect 2593 1417 2614 1488
rect 2672 1417 2686 1488
rect 2593 1408 2686 1417
rect 2593 1374 2622 1408
rect 2639 1374 2659 1408
rect 2676 1374 2686 1408
rect 2593 1335 2686 1374
rect 2602 1287 2676 1335
rect 2302 135 2337 139
rect 2302 101 2306 135
rect 2332 101 2337 135
rect 2302 98 2337 101
rect 409 46 465 53
rect 409 7 415 46
rect 454 7 465 46
rect 409 1 465 7
rect 3020 -484 3053 1850
rect 3015 -485 3058 -484
rect 3012 -487 3061 -485
rect 3012 -530 3015 -487
rect 3058 -530 3061 -487
rect 3012 -531 3061 -530
rect 3015 -533 3058 -531
rect 3085 -563 3118 1994
rect 3076 -566 3125 -563
rect 3076 -609 3080 -566
rect 3123 -609 3125 -566
rect 3076 -612 3125 -609
rect 3150 -634 3183 2158
rect 3147 -637 3187 -634
rect 3147 -680 3187 -677
rect 3126 -720 3184 -718
rect 3126 -771 3130 -720
rect 3181 -729 3184 -720
rect 3217 -729 3250 2315
rect 3281 -271 3314 2832
rect 3281 -717 3313 -271
rect 3342 -656 3375 2980
rect 3404 -595 3437 3135
rect 3467 -528 3500 3293
rect 3527 -462 3560 3841
rect 3585 -405 3618 3997
rect 3646 -338 3679 4151
rect 3705 -277 3738 4307
rect 3769 -210 3802 4365
rect 3831 -145 3864 4525
rect 3891 -82 3924 4674
rect 3954 -21 3987 4846
rect 4167 4359 4191 4370
rect 4461 4359 4492 4370
rect 4894 4355 4923 4371
rect 5040 4319 5059 5619
rect 5468 4315 5493 5718
rect 5638 5714 5711 5718
rect 5654 4675 5671 5714
rect 6154 5661 6251 6386
rect 7416 6284 7735 6396
rect 6693 5924 6840 5930
rect 6693 5882 6697 5924
rect 6832 5882 6840 5924
rect 6693 5877 6840 5882
rect 6456 5663 6500 5666
rect 6152 5659 6253 5661
rect 6152 5618 6155 5659
rect 6250 5618 6253 5659
rect 6152 5614 6253 5618
rect 6456 5616 6500 5619
rect 5876 5267 5910 5270
rect 5876 5241 5881 5267
rect 5907 5241 5910 5267
rect 5881 5238 5907 5241
rect 5693 4914 5719 4917
rect 5693 4885 5719 4888
rect 5696 4662 5715 4885
rect 5883 4660 5904 5238
rect 6240 5178 6266 5179
rect 6238 5176 6268 5178
rect 6238 5150 6240 5176
rect 6266 5150 6268 5176
rect 6238 5148 6268 5150
rect 6240 5147 6266 5148
rect 5923 5074 5957 5077
rect 5923 5048 5927 5074
rect 5953 5048 5957 5074
rect 5923 5045 5957 5048
rect 5930 4662 5949 5045
rect 5967 4865 5996 4868
rect 5967 4839 5969 4865
rect 5995 4839 5996 4865
rect 5967 4836 5996 4839
rect 5971 4660 5992 4836
rect 6071 4817 6105 4820
rect 6071 4791 6075 4817
rect 6101 4791 6105 4817
rect 6071 4788 6105 4791
rect 6079 4663 6097 4788
rect 6243 4124 6263 5147
rect 6466 4658 6489 5616
rect 6556 5268 6584 5271
rect 6556 5242 6557 5268
rect 6583 5242 6584 5268
rect 6556 5239 6584 5242
rect 6512 5177 6540 5180
rect 6512 5151 6513 5177
rect 6539 5151 6540 5177
rect 6512 5148 6540 5151
rect 6241 4111 6263 4124
rect 6236 4108 6269 4111
rect 6236 4081 6239 4108
rect 6266 4081 6269 4108
rect 6236 4078 6269 4081
rect 6489 4067 6490 4083
rect 6515 3994 6537 5148
rect 6514 3987 6537 3994
rect 6513 3927 6533 3987
rect 6558 3942 6581 5239
rect 6695 4639 6737 5877
rect 6798 4639 6840 5877
rect 7036 5659 7080 5662
rect 7036 5612 7080 5615
rect 7046 4914 7069 5612
rect 7488 5087 7616 6284
rect 7864 5765 7892 5777
rect 7864 5762 7897 5765
rect 7864 5718 7869 5762
rect 7864 5715 7897 5718
rect 7488 5079 7618 5087
rect 7487 5078 7618 5079
rect 7487 5052 7491 5078
rect 7613 5052 7618 5078
rect 7487 5049 7618 5052
rect 7165 5013 7195 5016
rect 7165 4987 7167 5013
rect 7193 4987 7195 5013
rect 7165 4984 7195 4987
rect 7033 4913 7069 4914
rect 7030 4911 7069 4913
rect 7030 4829 7036 4911
rect 7062 4829 7069 4911
rect 7030 4824 7069 4829
rect 7046 4658 7069 4824
rect 7168 4658 7191 4984
rect 7796 4959 7839 4963
rect 7796 4933 7800 4959
rect 7826 4933 7839 4959
rect 7796 4929 7839 4933
rect 7820 4662 7839 4929
rect 7864 4653 7892 5715
rect 8034 5268 8060 5271
rect 8034 5239 8060 5242
rect 7945 5181 7971 5184
rect 7945 5152 7971 5155
rect 7948 4780 7967 5152
rect 8036 4780 8058 5239
rect 8233 4917 8267 6539
rect 10273 6287 10592 6399
rect 8683 6193 8720 6194
rect 8678 6189 8728 6193
rect 8678 6152 8686 6189
rect 8723 6152 8728 6189
rect 8678 6148 8728 6152
rect 8298 5340 8330 5344
rect 8298 5313 8301 5340
rect 8327 5313 8330 5340
rect 8298 5307 8330 5313
rect 8228 4911 8267 4917
rect 8228 4909 8231 4911
rect 8227 4832 8231 4909
rect 8263 4832 8267 4911
rect 8228 4825 8267 4832
rect 7931 4760 7999 4780
rect 7931 4734 7945 4760
rect 7971 4734 7999 4760
rect 7931 4711 7999 4734
rect 8035 4761 8103 4780
rect 8035 4735 8047 4761
rect 8073 4735 8103 4761
rect 8035 4711 8103 4735
rect 8233 4647 8267 4825
rect 8300 4769 8327 5307
rect 8300 4766 8368 4769
rect 8300 4723 8322 4766
rect 8365 4723 8368 4766
rect 8300 4719 8368 4723
rect 8300 4654 8327 4719
rect 6514 3924 6537 3927
rect 4157 3318 4181 3755
rect 4451 3311 4482 3762
rect 4894 3313 4923 3760
rect 5040 3364 5059 3754
rect 5171 3374 5194 3758
rect 5468 3375 5493 3760
rect 6515 3604 6537 3924
rect 6515 3595 6550 3604
rect 6515 3573 6566 3595
rect 5038 3314 5059 3364
rect 5169 3333 5194 3374
rect 5466 3333 5493 3375
rect 5644 3390 5672 3501
rect 5697 3432 5716 3492
rect 5897 3448 5936 3450
rect 5896 3445 5936 3448
rect 5896 3439 5903 3445
rect 5881 3438 5903 3439
rect 5697 3413 5857 3432
rect 5644 3362 5816 3390
rect 5796 3339 5816 3362
rect 5038 3301 5057 3314
rect 5169 3290 5192 3333
rect 5466 3296 5491 3333
rect 5797 3309 5813 3339
rect 5838 3301 5857 3413
rect 5878 3417 5903 3438
rect 5931 3417 5936 3445
rect 5878 3414 5936 3417
rect 5878 3412 5935 3414
rect 5878 3411 5897 3412
rect 5878 3327 5895 3411
rect 6345 3405 6368 3496
rect 6467 3408 6490 3496
rect 6293 3398 6368 3405
rect 6290 3382 6368 3398
rect 6465 3402 6490 3408
rect 6798 3415 6840 3515
rect 6290 3337 6331 3382
rect 5878 3300 5894 3327
rect 6290 3288 6328 3337
rect 6465 3302 6489 3402
rect 6798 3397 6841 3415
rect 6798 3358 6842 3397
rect 7046 3376 7069 3496
rect 6801 3337 6842 3358
rect 6801 3286 6841 3337
rect 7045 3302 7069 3376
rect 7168 3407 7191 3496
rect 7168 3369 7244 3407
rect 7820 3394 7839 3492
rect 7206 3323 7244 3369
rect 7637 3386 7665 3389
rect 7637 3360 7638 3386
rect 7664 3360 7665 3386
rect 7637 3357 7665 3360
rect 7680 3375 7839 3394
rect 7640 3309 7656 3357
rect 7680 3342 7699 3375
rect 7864 3356 7892 3501
rect 8683 3457 8720 6148
rect 8762 5843 8808 5846
rect 8762 5806 8768 5843
rect 8805 5806 8808 5843
rect 8762 5803 8808 5806
rect 8680 3452 8725 3457
rect 8680 3415 8687 3452
rect 8724 3415 8725 3452
rect 8680 3411 8725 3415
rect 8683 3407 8720 3411
rect 8764 3398 8801 5803
rect 8839 5372 8884 5375
rect 8839 5335 8845 5372
rect 8882 5335 8884 5372
rect 8839 5332 8884 5335
rect 7725 3355 7892 3356
rect 7677 3331 7699 3342
rect 7677 3301 7696 3331
rect 7721 3328 7892 3355
rect 8761 3393 8805 3398
rect 8761 3356 8764 3393
rect 8801 3356 8805 3393
rect 8761 3352 8805 3356
rect 8764 3347 8801 3352
rect 7721 3309 7737 3328
rect 8841 3163 8878 5332
rect 9496 5280 9554 5283
rect 9496 5230 9500 5280
rect 9550 5230 9554 5280
rect 9496 5227 9554 5230
rect 9378 5220 9434 5224
rect 9270 5173 9326 5177
rect 9175 5124 9231 5135
rect 9175 5074 9178 5124
rect 9228 5074 9231 5124
rect 9175 5070 9231 5074
rect 9270 5123 9273 5173
rect 9323 5123 9326 5173
rect 9378 5170 9381 5220
rect 9431 5170 9434 5220
rect 9378 5165 9434 5170
rect 9270 5119 9326 5123
rect 8928 4865 8971 4868
rect 8928 4828 8933 4865
rect 8970 4828 8971 4865
rect 8928 4824 8971 4828
rect 8838 3162 8878 3163
rect 8837 3160 8879 3162
rect 8837 3123 8838 3160
rect 8875 3123 8879 3160
rect 8837 3120 8879 3123
rect 8841 3119 8878 3120
rect 4157 2656 4181 2742
rect 4451 2656 4482 2749
rect 4157 2365 4191 2656
rect 4451 2365 4492 2656
rect 4894 2365 4923 2747
rect 4167 2341 4191 2365
rect 4461 2338 4492 2365
rect 5040 2338 5059 2747
rect 5171 2643 5194 2751
rect 5162 2639 5195 2643
rect 5162 2598 5166 2639
rect 5192 2598 5195 2639
rect 5162 2595 5195 2598
rect 5171 2334 5194 2595
rect 5468 2355 5493 2753
rect 5800 2349 5816 2754
rect 6075 2390 6099 2762
rect 6073 2365 6112 2390
rect 6087 2340 6112 2365
rect 6293 2327 6331 2776
rect 6468 2388 6492 2762
rect 6468 2361 6515 2388
rect 6488 2338 6515 2361
rect 6696 2325 6736 2778
rect 7048 2511 7072 2762
rect 8929 2645 8966 4824
rect 8925 2639 8974 2645
rect 8925 2598 8931 2639
rect 8968 2598 8974 2639
rect 8925 2594 8974 2598
rect 8929 2591 8966 2594
rect 7048 2487 7106 2511
rect 7082 2353 7106 2487
rect 5603 2252 5635 2256
rect 5603 2226 5606 2252
rect 5632 2226 5635 2252
rect 7594 2250 7620 2253
rect 5603 2222 5635 2226
rect 7593 2224 7594 2247
rect 4157 502 4181 1765
rect 4451 1657 4482 1772
rect 4894 1708 4923 1770
rect 4944 1739 4978 1742
rect 4944 1713 4948 1739
rect 4974 1713 4978 1739
rect 4944 1710 4978 1713
rect 4891 1705 4926 1708
rect 4891 1676 4894 1705
rect 4923 1676 4926 1705
rect 4891 1673 4926 1676
rect 4447 1656 4484 1657
rect 4447 1625 4450 1656
rect 4481 1625 4484 1656
rect 4894 1627 4923 1673
rect 4944 1649 4969 1710
rect 5040 1651 5059 1771
rect 5468 1704 5493 1777
rect 5611 1746 5632 2222
rect 7593 2221 7620 2224
rect 7542 2157 7568 2160
rect 7542 2128 7568 2131
rect 5737 2053 5776 2078
rect 5665 1974 5699 1977
rect 5665 1948 5669 1974
rect 5695 1948 5699 1974
rect 5665 1943 5699 1948
rect 5669 1941 5691 1943
rect 5608 1743 5636 1746
rect 5608 1717 5609 1743
rect 5635 1717 5636 1743
rect 5608 1714 5636 1717
rect 5669 1713 5689 1941
rect 5715 1759 5734 1795
rect 5711 1742 5739 1759
rect 5711 1716 5712 1742
rect 5738 1716 5739 1742
rect 5665 1710 5693 1713
rect 5711 1712 5739 1716
rect 5465 1702 5499 1704
rect 5465 1676 5469 1702
rect 5495 1676 5499 1702
rect 5665 1684 5666 1710
rect 5692 1684 5693 1710
rect 5665 1681 5693 1684
rect 5465 1675 5499 1676
rect 4447 1624 4484 1625
rect 4451 1503 4482 1624
rect 4837 1599 4923 1627
rect 4829 1598 4923 1599
rect 4939 1638 4969 1649
rect 5034 1648 5066 1651
rect 4829 1596 4875 1598
rect 4829 1554 4831 1596
rect 4873 1554 4875 1596
rect 4829 1551 4875 1554
rect 4446 1500 4488 1503
rect 4939 1487 4958 1638
rect 5034 1622 5037 1648
rect 5063 1622 5066 1648
rect 5034 1619 5066 1622
rect 5302 1598 5377 1617
rect 5327 1514 5377 1598
rect 5758 1590 5776 2053
rect 7495 1973 7521 1976
rect 7495 1944 7521 1947
rect 7445 1880 7471 1883
rect 7445 1851 7471 1854
rect 5890 1706 5916 1709
rect 5888 1704 5918 1706
rect 5888 1678 5890 1704
rect 5916 1678 5918 1704
rect 5888 1676 5918 1678
rect 5890 1675 5916 1676
rect 5758 1586 5806 1590
rect 5758 1560 5770 1586
rect 5766 1553 5770 1560
rect 5803 1553 5806 1586
rect 5891 1583 5913 1675
rect 6087 1662 6112 1785
rect 6488 1664 6515 1787
rect 6770 1744 6813 1747
rect 6770 1709 6774 1744
rect 6809 1709 6813 1744
rect 6770 1707 6813 1709
rect 6086 1636 6089 1662
rect 6115 1636 6118 1662
rect 6488 1660 6523 1664
rect 6488 1633 6493 1660
rect 6520 1633 6523 1660
rect 5766 1549 5806 1553
rect 5885 1580 5919 1583
rect 5885 1543 5919 1546
rect 5891 1535 5913 1543
rect 6286 1516 6380 1609
rect 6774 1564 6809 1707
rect 6956 1651 6978 1783
rect 7082 1711 7105 1783
rect 7082 1688 7403 1711
rect 7082 1687 7105 1688
rect 6774 1532 6778 1564
rect 6804 1532 6809 1564
rect 6774 1528 6809 1532
rect 6927 1627 6978 1651
rect 4446 1455 4488 1458
rect 4895 1481 4958 1487
rect 5278 1482 5302 1514
rect 5402 1482 5426 1514
rect 6259 1484 6283 1516
rect 6383 1484 6407 1516
rect 6927 1502 6950 1627
rect 7380 1591 7403 1688
rect 7375 1588 7406 1591
rect 7375 1554 7377 1588
rect 7403 1554 7406 1588
rect 7375 1551 7406 1554
rect 6916 1499 6962 1502
rect 4895 1449 4899 1481
rect 4931 1455 4958 1481
rect 6916 1461 6920 1499
rect 6958 1461 6962 1499
rect 6916 1458 6962 1461
rect 4931 1449 4939 1455
rect 4895 1445 4939 1449
rect 5278 1348 5302 1380
rect 5402 1347 5426 1379
rect 6259 1350 6283 1382
rect 6383 1349 6407 1381
rect 7380 1234 7403 1551
rect 7367 1212 7403 1234
rect 7347 1189 7403 1212
rect 7347 1188 7401 1189
rect 4916 927 4948 1102
rect 5278 1071 5302 1103
rect 5402 1070 5426 1102
rect 5302 1005 5328 1051
rect 5376 1007 5402 1051
rect 5301 1002 5329 1005
rect 5301 971 5329 974
rect 5375 1004 5403 1007
rect 5375 973 5403 976
rect 4904 917 4958 927
rect 4904 871 4909 917
rect 4955 871 4958 917
rect 4904 867 4958 871
rect 5302 830 5328 971
rect 5376 830 5402 973
rect 4117 485 4182 502
rect 5302 487 5402 830
rect 5753 825 5787 1104
rect 5747 822 5793 825
rect 5747 773 5793 776
rect 5896 736 5930 1103
rect 6259 1073 6283 1105
rect 6383 1073 6407 1105
rect 6283 1005 6309 1054
rect 6282 1002 6310 1005
rect 6282 971 6310 974
rect 6283 853 6309 971
rect 6357 853 6383 1054
rect 5887 733 5939 736
rect 5887 687 5890 733
rect 5936 687 5939 733
rect 5887 684 5939 687
rect 6283 493 6383 853
rect 6738 648 6765 1107
rect 7445 1067 7470 1851
rect 7495 1157 7520 1944
rect 7543 1248 7568 2128
rect 7593 1337 7618 2221
rect 9177 1487 9227 5070
rect 9270 2015 9320 5119
rect 9383 2538 9433 5165
rect 9496 3055 9546 5227
rect 10382 5067 10510 6287
rect 10381 5064 10510 5067
rect 10509 4936 10510 5064
rect 10381 4933 10510 4936
rect 10382 4884 10510 4933
rect 10818 4766 10838 4769
rect 10809 4763 10840 4766
rect 10809 4720 10813 4763
rect 10839 4720 10840 4763
rect 10809 4716 10840 4720
rect 10427 4634 10462 4637
rect 10427 4592 10430 4634
rect 10456 4592 10462 4634
rect 10427 4589 10462 4592
rect 10028 4312 10075 4318
rect 10028 4272 10030 4312
rect 10070 4272 10075 4312
rect 10028 4269 10075 4272
rect 9491 3052 9546 3055
rect 9541 3002 9546 3052
rect 9491 2999 9546 3002
rect 9382 2530 9434 2538
rect 9382 2483 9383 2530
rect 9433 2483 9434 2530
rect 9382 2482 9434 2483
rect 9269 2014 9321 2015
rect 9269 1964 9270 2014
rect 9320 1964 9321 2014
rect 9269 1963 9321 1964
rect 9161 1484 9227 1487
rect 9161 1434 9165 1484
rect 9215 1434 9227 1484
rect 9161 1430 9227 1434
rect 7588 1333 7625 1337
rect 7588 1283 7592 1333
rect 7618 1283 7625 1333
rect 7588 1279 7625 1283
rect 7535 1243 7572 1248
rect 7535 1193 7538 1243
rect 7564 1193 7572 1243
rect 7535 1190 7572 1193
rect 7486 1153 7523 1157
rect 7486 1103 7491 1153
rect 7517 1103 7523 1153
rect 7486 1099 7523 1103
rect 7439 1063 7474 1067
rect 6727 642 6776 648
rect 6727 596 6729 642
rect 6775 596 6776 642
rect 6727 592 6776 596
rect 6283 489 6485 493
rect 4117 373 4122 485
rect 4148 373 4182 485
rect 5254 483 5447 487
rect 4117 370 4182 373
rect 5200 481 5447 483
rect 5200 479 5333 481
rect 5200 367 5259 479
rect 5445 369 5447 481
rect 5371 367 5447 369
rect 5200 364 5447 367
rect 6235 483 6485 489
rect 6235 364 6240 483
rect 6426 364 6485 483
rect 3952 -23 3989 -21
rect 3952 -56 3954 -23
rect 3987 -56 3989 -23
rect 3952 -59 3989 -56
rect 3887 -85 3926 -82
rect 3887 -118 3892 -85
rect 3925 -118 3926 -85
rect 3887 -121 3926 -118
rect 3827 -148 3865 -145
rect 3827 -181 3829 -148
rect 3862 -181 3865 -148
rect 3827 -184 3865 -181
rect 3768 -211 3803 -210
rect 3768 -244 3769 -211
rect 3802 -244 3803 -211
rect 3768 -247 3803 -244
rect 3704 -279 3740 -277
rect 3704 -312 3705 -279
rect 3738 -312 3740 -279
rect 3704 -315 3740 -312
rect 3645 -339 3679 -338
rect 3643 -341 3681 -339
rect 3643 -374 3645 -341
rect 3678 -374 3681 -341
rect 3643 -376 3681 -374
rect 3645 -377 3678 -376
rect 3585 -441 3618 -438
rect 3527 -498 3560 -495
rect 3467 -531 3502 -528
rect 3467 -561 3469 -531
rect 3469 -567 3502 -564
rect 3404 -631 3437 -628
rect 3340 -659 3375 -656
rect 3373 -689 3375 -659
rect 3340 -696 3373 -693
rect 3181 -762 3250 -729
rect 3279 -720 3323 -717
rect 3279 -757 3282 -720
rect 3319 -757 3323 -720
rect 3279 -759 3323 -757
rect 3181 -771 3184 -762
rect 3126 -773 3184 -771
rect 5200 -785 5294 364
rect 6235 361 6485 364
rect 6396 -639 6485 361
rect 7312 46 7345 1045
rect 7439 1013 7443 1063
rect 7469 1013 7474 1063
rect 7439 1010 7474 1013
rect 9177 648 9227 1430
rect 9270 739 9320 1963
rect 9383 826 9433 2482
rect 9496 928 9546 2999
rect 9785 1736 9843 1740
rect 9785 1686 9789 1736
rect 9839 1686 9843 1736
rect 9785 1684 9843 1686
rect 9788 1683 9839 1684
rect 9496 925 9552 928
rect 9496 875 9502 925
rect 9496 872 9552 875
rect 9496 859 9546 872
rect 9383 777 9433 780
rect 9270 690 9320 693
rect 9177 599 9227 602
rect 9788 496 9838 1683
rect 9725 485 9838 496
rect 9725 373 9731 485
rect 9825 373 9838 485
rect 9725 368 9838 373
rect 7306 43 7349 46
rect 7306 10 7310 43
rect 7343 10 7349 43
rect 7306 7 7349 10
rect 10033 -66 10073 4269
rect 10125 4208 10128 4244
rect 10164 4208 10167 4244
rect 10032 -69 10079 -66
rect 10032 -109 10036 -69
rect 10076 -109 10079 -69
rect 10032 -112 10079 -109
rect 10126 -146 10165 4208
rect 10217 4010 10262 4012
rect 10217 3971 10220 4010
rect 10259 3971 10262 4010
rect 10217 3969 10262 3971
rect 10123 -150 10169 -146
rect 10123 -189 10127 -150
rect 10166 -189 10169 -150
rect 10123 -193 10169 -189
rect 10219 -228 10258 3969
rect 10303 3943 10341 3944
rect 10301 3941 10343 3943
rect 10301 3915 10303 3941
rect 10341 3915 10343 3941
rect 10301 3913 10343 3915
rect 10217 -232 10264 -228
rect 10217 -271 10220 -232
rect 10259 -271 10264 -232
rect 10217 -274 10264 -271
rect 10303 -308 10341 3913
rect 10437 1590 10460 4589
rect 10818 4391 10838 4716
rect 11169 4392 11188 6419
rect 11503 5540 11585 5543
rect 11503 5534 11508 5540
rect 11497 5469 11508 5534
rect 11579 5469 11585 5540
rect 11497 5465 11585 5469
rect 11497 3565 11568 5465
rect 11484 3561 11568 3565
rect 11484 3490 11489 3561
rect 11560 3490 11568 3561
rect 11484 3486 11568 3490
rect 11056 1736 11128 1739
rect 11056 1685 11069 1736
rect 11120 1685 11128 1736
rect 11056 1682 11128 1685
rect 10437 1567 10461 1590
rect 10437 986 10460 1567
rect 11062 981 11113 1682
rect 11048 976 11113 981
rect 11047 958 11113 976
rect 11044 957 11113 958
rect 11044 951 11104 957
rect 11044 733 11078 951
rect 11009 634 11078 733
rect 11044 556 11078 634
rect 11049 496 11078 556
rect 11045 495 11078 496
rect 11044 395 11078 495
rect 11049 335 11078 395
rect 11044 234 11078 335
rect 11048 174 11078 234
rect 11044 72 11078 174
rect 11049 12 11078 72
rect 11044 -89 11078 12
rect 11048 -149 11078 -89
rect 10300 -312 10344 -308
rect 10300 -350 10302 -312
rect 10340 -350 10344 -312
rect 11044 -336 11078 -149
rect 10300 -354 10344 -350
rect 11048 -544 11078 -336
rect 11095 920 11104 951
rect 11095 -544 11102 920
rect 11048 -557 11102 -544
rect 6396 -712 6488 -639
rect 6393 -785 6485 -712
<< via1 >>
rect 421 6215 460 6254
rect 429 5870 468 5909
rect 567 5753 593 5779
rect 559 5483 601 5525
rect 1154 5343 1183 5401
rect 2483 5237 2509 5263
rect 3062 5194 3093 5225
rect 4720 5958 4762 6000
rect 4335 5882 4377 5924
rect 4887 5721 4931 5765
rect 5459 5721 5503 5765
rect 5641 5718 5685 5762
rect 4445 5619 4489 5663
rect 4169 5317 4195 5343
rect 3462 5248 3488 5274
rect 3345 5149 3372 5175
rect 2212 5071 2247 5106
rect 2737 5102 2763 5128
rect 5016 5619 5060 5663
rect 2314 4847 2340 4886
rect 3954 4848 3987 4874
rect 2250 4765 2276 4805
rect 2252 4654 2278 4680
rect 1875 4612 1901 4638
rect 1872 4520 1898 4546
rect 1873 4428 1899 4454
rect 1808 4326 1834 4352
rect 1804 4230 1830 4256
rect 1808 4134 1834 4160
rect 2252 4562 2278 4588
rect 2249 4470 2275 4496
rect 1804 2606 1830 2653
rect 1868 2606 1894 2653
rect 1668 2503 1694 2529
rect 1616 2463 1642 2489
rect 688 2338 754 2404
rect 1876 2501 1902 2527
rect 2052 2502 2079 2529
rect 1810 2465 1836 2491
rect 1618 2072 1644 2098
rect 1209 1886 1246 1923
rect 692 1752 758 1818
rect 2102 2463 2128 2489
rect 1208 1262 1245 1299
rect 1962 1220 1988 1256
rect 1507 696 1536 725
rect 3891 4676 3924 4709
rect 3834 4528 3867 4561
rect 2313 4361 2339 4387
rect 3770 4368 3803 4401
rect 3706 4311 3739 4344
rect 2314 4265 2340 4291
rect 2313 4169 2339 4195
rect 2249 2403 2275 2429
rect 2187 2288 2213 2314
rect 2145 2027 2171 2053
rect 2189 1458 2215 1500
rect 2185 1220 2211 1256
rect 3645 4154 3678 4187
rect 3582 4001 3615 4034
rect 3526 3844 3559 3877
rect 3464 3297 3497 3330
rect 3401 3138 3434 3171
rect 3339 2983 3372 3016
rect 3279 2835 3312 2868
rect 3215 2318 3248 2351
rect 3148 2161 3181 2194
rect 2313 1970 2339 1996
rect 3086 1997 3119 2030
rect 2247 857 2273 890
rect 2144 695 2173 724
rect 2028 594 2088 654
rect 3018 1853 3051 1886
rect 2614 1417 2672 1488
rect 2306 101 2332 135
rect 415 7 454 46
rect 3015 -530 3058 -487
rect 3080 -609 3123 -566
rect 3147 -677 3187 -637
rect 3130 -771 3181 -720
rect 6697 5882 6832 5924
rect 6155 5618 6250 5659
rect 6456 5619 6500 5663
rect 5881 5241 5907 5267
rect 5693 4888 5719 4914
rect 6240 5150 6266 5176
rect 5927 5048 5953 5074
rect 5969 4839 5995 4865
rect 6075 4791 6101 4817
rect 6557 5242 6583 5268
rect 6513 5151 6539 5177
rect 6239 4081 6266 4108
rect 7036 5615 7080 5659
rect 7869 5718 7897 5762
rect 7491 5052 7613 5078
rect 7167 4987 7193 5013
rect 7800 4933 7826 4959
rect 8034 5242 8060 5268
rect 7945 5155 7971 5181
rect 8686 6152 8723 6189
rect 8301 5313 8327 5340
rect 7945 4734 7971 4760
rect 8047 4735 8073 4761
rect 8322 4723 8365 4766
rect 5903 3417 5931 3445
rect 7638 3360 7664 3386
rect 8768 5806 8805 5843
rect 8687 3415 8724 3452
rect 8845 5335 8882 5372
rect 8764 3356 8801 3393
rect 9500 5230 9550 5280
rect 9178 5074 9228 5124
rect 9273 5123 9323 5173
rect 9381 5170 9431 5220
rect 8933 4828 8970 4865
rect 8838 3123 8875 3160
rect 5166 2598 5192 2639
rect 8931 2598 8968 2639
rect 5606 2226 5632 2252
rect 7594 2224 7620 2250
rect 4948 1713 4974 1739
rect 4894 1676 4923 1705
rect 4450 1625 4481 1656
rect 7542 2131 7568 2157
rect 5669 1948 5695 1974
rect 5609 1717 5635 1743
rect 5712 1716 5738 1742
rect 5469 1676 5495 1702
rect 5666 1684 5692 1710
rect 4831 1554 4873 1596
rect 4446 1458 4488 1500
rect 5037 1622 5063 1648
rect 7495 1947 7521 1973
rect 7445 1854 7471 1880
rect 5890 1678 5916 1704
rect 5770 1553 5803 1586
rect 6774 1709 6809 1744
rect 6089 1636 6115 1662
rect 6493 1633 6520 1660
rect 5885 1546 5919 1580
rect 6778 1532 6804 1564
rect 7377 1554 7403 1588
rect 4899 1449 4931 1481
rect 6920 1461 6958 1499
rect 5301 974 5329 1002
rect 5375 976 5403 1004
rect 4909 871 4955 917
rect 5747 776 5793 822
rect 6282 974 6310 1002
rect 5890 687 5936 733
rect 10381 4936 10509 5064
rect 10813 4720 10839 4763
rect 10430 4592 10456 4634
rect 10030 4272 10070 4312
rect 9491 3002 9541 3052
rect 9383 2483 9433 2530
rect 9270 1964 9320 2014
rect 9165 1434 9215 1484
rect 7592 1283 7618 1333
rect 7538 1193 7564 1243
rect 7491 1103 7517 1153
rect 6729 596 6775 642
rect 4122 373 4148 485
rect 5333 479 5445 481
rect 5259 369 5445 479
rect 5259 367 5371 369
rect 6240 364 6426 483
rect 3954 -56 3987 -23
rect 3892 -118 3925 -85
rect 3829 -181 3862 -148
rect 3769 -244 3802 -211
rect 3705 -312 3738 -279
rect 3645 -374 3678 -341
rect 3585 -438 3618 -405
rect 3527 -495 3560 -462
rect 3469 -564 3502 -531
rect 3404 -628 3437 -595
rect 3340 -693 3373 -659
rect 3282 -757 3319 -720
rect 7443 1013 7469 1063
rect 9789 1686 9839 1736
rect 9502 875 9552 925
rect 9383 780 9433 826
rect 9270 693 9320 739
rect 9177 602 9227 648
rect 9731 373 9825 485
rect 7310 10 7343 43
rect 10128 4208 10164 4244
rect 10036 -109 10076 -69
rect 10220 3971 10259 4010
rect 10127 -189 10166 -150
rect 10303 3915 10341 3941
rect 10220 -271 10259 -232
rect 11508 5469 11579 5540
rect 11489 3490 11560 3561
rect 11069 1685 11120 1736
rect 10302 -350 10340 -312
<< metal2 >>
rect 295 6246 363 6368
rect 418 6254 463 6256
rect 418 6246 421 6254
rect 295 6223 421 6246
rect 295 6136 363 6223
rect 418 6215 421 6223
rect 460 6215 463 6254
rect 418 6213 463 6215
rect 8680 6189 8726 6191
rect 11767 6189 11853 6324
rect 8680 6152 8686 6189
rect 8723 6152 11853 6189
rect 8680 6150 8726 6152
rect 11767 6114 11853 6152
rect 280 6026 528 6027
rect 280 5987 675 6026
rect 507 5950 675 5987
rect 2273 6017 2348 6018
rect 2273 5987 2435 6017
rect 4718 6000 4763 6002
rect 4717 5994 4720 6000
rect 2273 5970 2297 5987
rect 2405 5965 2435 5987
rect 2478 5964 4720 5994
rect 4717 5958 4720 5964
rect 4762 5958 4765 6000
rect 4718 5956 4763 5958
rect 4333 5924 4378 5926
rect 6694 5924 6836 5927
rect 295 5827 363 5915
rect 428 5909 471 5913
rect 428 5870 429 5909
rect 468 5870 471 5909
rect 4332 5882 4335 5924
rect 4377 5923 4380 5924
rect 6694 5923 6697 5924
rect 4377 5883 6697 5923
rect 4377 5882 4380 5883
rect 6694 5882 6697 5883
rect 6832 5923 6836 5924
rect 6832 5883 6841 5923
rect 6832 5882 6836 5883
rect 4333 5880 4378 5882
rect 6694 5879 6836 5882
rect 428 5866 471 5870
rect 428 5865 622 5866
rect 437 5843 622 5865
rect 8763 5843 8807 5845
rect 11767 5843 11853 5911
rect 295 5795 631 5827
rect 8763 5806 8768 5843
rect 8805 5806 11853 5843
rect 8763 5804 8807 5806
rect 295 5683 363 5795
rect 564 5753 567 5779
rect 593 5756 622 5779
rect 593 5753 596 5756
rect 4884 5721 4887 5765
rect 4931 5762 4934 5765
rect 5456 5762 5459 5765
rect 4931 5721 5459 5762
rect 5503 5762 5506 5765
rect 5503 5721 5641 5762
rect 4899 5718 5641 5721
rect 5685 5718 7869 5762
rect 7897 5718 7900 5762
rect 11767 5701 11853 5806
rect 5016 5663 5060 5666
rect 495 5646 648 5662
rect 314 5613 648 5646
rect 4442 5619 4445 5663
rect 4489 5661 4492 5663
rect 4489 5619 5016 5661
rect 6453 5661 6456 5663
rect 5060 5659 6456 5661
rect 5060 5619 6155 5659
rect 4457 5618 6155 5619
rect 6250 5619 6456 5659
rect 6500 5661 6503 5663
rect 6500 5659 7093 5661
rect 6500 5619 7036 5659
rect 6250 5618 7036 5619
rect 4457 5617 7036 5618
rect 5016 5616 5060 5617
rect 7033 5615 7036 5617
rect 7080 5617 7093 5659
rect 7080 5615 7083 5617
rect 314 5606 541 5613
rect 314 5586 354 5606
rect 279 5546 354 5586
rect 11505 5525 11508 5540
rect 556 5483 559 5525
rect 601 5483 11508 5525
rect 11505 5469 11508 5483
rect 11579 5469 11582 5540
rect 250 5401 318 5468
rect 1142 5401 1189 5403
rect 250 5343 1154 5401
rect 1183 5343 1189 5401
rect 8841 5372 8883 5374
rect 11764 5372 11850 5502
rect 250 5319 322 5343
rect 1142 5341 1189 5343
rect 4167 5343 4197 5346
rect 250 5236 318 5319
rect 4167 5317 4169 5343
rect 4195 5340 4197 5343
rect 8299 5340 8329 5343
rect 4195 5317 8301 5340
rect 4167 5314 4197 5317
rect 8299 5313 8301 5317
rect 8327 5317 8336 5340
rect 8841 5335 8845 5372
rect 8882 5335 11850 5372
rect 8841 5333 8883 5335
rect 8327 5313 8329 5317
rect 8299 5309 8329 5313
rect 11764 5292 11850 5335
rect 3459 5274 3490 5276
rect 2480 5266 2512 5267
rect 3459 5266 3462 5274
rect 2480 5263 3462 5266
rect 2480 5237 2483 5263
rect 2509 5248 3462 5263
rect 3488 5266 3491 5274
rect 5877 5267 5909 5269
rect 6554 5268 6586 5269
rect 5877 5266 5881 5267
rect 3488 5248 5881 5266
rect 2509 5243 5881 5248
rect 2509 5237 2512 5243
rect 3459 5242 3490 5243
rect 5877 5241 5881 5243
rect 5907 5266 5910 5267
rect 6554 5266 6557 5268
rect 5907 5243 6557 5266
rect 5907 5241 5910 5243
rect 6554 5242 6557 5243
rect 6583 5266 6586 5268
rect 8031 5266 8034 5268
rect 6583 5243 8034 5266
rect 6583 5242 6586 5243
rect 8031 5242 8034 5243
rect 8060 5266 8063 5268
rect 9497 5266 9500 5280
rect 8060 5243 9500 5266
rect 8060 5242 8063 5243
rect 6554 5241 6586 5242
rect 2480 5235 2512 5237
rect 9497 5230 9500 5243
rect 9550 5230 9553 5280
rect 9497 5229 9553 5230
rect 3059 5225 3096 5227
rect 250 5186 301 5198
rect 3059 5194 3062 5225
rect 3093 5221 3096 5225
rect 9379 5221 9433 5223
rect 3093 5220 9433 5221
rect 3093 5198 9381 5220
rect 3093 5194 3096 5198
rect 3059 5192 3096 5194
rect 250 5157 560 5186
rect 6510 5177 6542 5178
rect 6239 5176 6267 5177
rect 301 5156 560 5157
rect 3342 5175 3373 5176
rect 6237 5175 6240 5176
rect 3342 5149 3345 5175
rect 3372 5152 6240 5175
rect 3372 5149 3375 5152
rect 6237 5150 6240 5152
rect 6266 5175 6269 5176
rect 6510 5175 6513 5177
rect 6266 5152 6513 5175
rect 6266 5150 6269 5152
rect 6510 5151 6513 5152
rect 6539 5175 6542 5177
rect 7942 5175 7945 5181
rect 6539 5155 7945 5175
rect 7971 5175 7974 5181
rect 9271 5175 9325 5176
rect 7971 5173 9325 5175
rect 7971 5155 9273 5173
rect 6539 5152 9273 5155
rect 6539 5151 6542 5152
rect 6510 5150 6542 5151
rect 6239 5149 6267 5150
rect 3342 5147 3373 5149
rect 2734 5129 2766 5130
rect 9177 5129 9230 5132
rect 2734 5128 9230 5129
rect 246 5106 297 5108
rect 2210 5106 2250 5107
rect 246 5071 2212 5106
rect 2247 5071 2250 5106
rect 2734 5102 2737 5128
rect 2763 5124 9230 5128
rect 2763 5106 9178 5124
rect 2763 5102 2766 5106
rect 2734 5100 2766 5102
rect 7489 5078 7617 5081
rect 246 5067 297 5071
rect 2210 5068 2250 5071
rect 5924 5074 5956 5075
rect 5924 5048 5927 5074
rect 5953 5071 5956 5074
rect 7489 5071 7491 5078
rect 5953 5052 7491 5071
rect 7613 5052 7617 5078
rect 9177 5074 9178 5106
rect 9228 5074 9230 5124
rect 9271 5123 9273 5152
rect 9323 5123 9325 5173
rect 9379 5170 9381 5198
rect 9431 5170 9433 5220
rect 9379 5167 9433 5170
rect 9271 5120 9325 5123
rect 9177 5071 9230 5074
rect 5953 5050 7617 5052
rect 5953 5048 5956 5050
rect 5924 5047 5956 5048
rect 218 4886 345 5032
rect 4930 5006 5215 5026
rect 7166 5013 7194 5015
rect 5195 4956 5215 5006
rect 7164 4987 7167 5013
rect 7193 5010 7196 5013
rect 10378 5010 10381 5064
rect 7193 4989 10381 5010
rect 7193 4987 7196 4989
rect 7166 4985 7194 4987
rect 7797 4959 7828 4962
rect 7797 4956 7800 4959
rect 4048 4921 4104 4938
rect 5195 4936 7800 4956
rect 7797 4933 7800 4936
rect 7826 4933 7828 4959
rect 10378 4936 10381 4989
rect 10509 4936 10512 5064
rect 7797 4930 7828 4933
rect 1353 4886 1383 4887
rect 2312 4886 2341 4888
rect 218 4847 2314 4886
rect 2340 4847 2344 4886
rect 3951 4848 3954 4874
rect 3987 4865 3990 4874
rect 4048 4865 4065 4921
rect 5690 4909 5693 4914
rect 5190 4889 5693 4909
rect 3987 4848 4066 4865
rect 5190 4851 5210 4889
rect 5690 4888 5693 4889
rect 5719 4909 5722 4914
rect 5719 4889 5727 4909
rect 5719 4888 5722 4889
rect 5966 4865 5997 4866
rect 8929 4865 8972 4867
rect 11764 4865 11850 5063
rect 5966 4862 5969 4865
rect 218 4844 345 4847
rect 2312 4845 2341 4847
rect 4930 4831 5210 4851
rect 5241 4842 5969 4862
rect 2248 4805 2277 4807
rect 1003 4765 2250 4805
rect 2276 4765 2279 4805
rect 247 4496 374 4583
rect 1003 4496 1043 4765
rect 2248 4764 2277 4765
rect 4048 4738 4104 4755
rect 3891 4711 3924 4712
rect 3889 4709 3926 4711
rect 1383 4697 1420 4698
rect 1204 4674 1420 4697
rect 2249 4675 2252 4680
rect 1204 4661 1946 4674
rect 1204 4591 1266 4661
rect 1383 4657 1946 4661
rect 2192 4658 2252 4675
rect 2249 4654 2252 4658
rect 2278 4675 2281 4680
rect 3889 4676 3891 4709
rect 3924 4701 3926 4709
rect 4048 4701 4065 4738
rect 3924 4684 4065 4701
rect 3924 4676 3926 4684
rect 4048 4683 4065 4684
rect 5241 4676 5261 4842
rect 5966 4839 5969 4842
rect 5995 4839 5998 4865
rect 5966 4838 5997 4839
rect 8929 4828 8933 4865
rect 8970 4853 11850 4865
rect 8970 4828 11839 4853
rect 8929 4825 8970 4828
rect 6072 4817 6104 4818
rect 6072 4814 6075 4817
rect 2278 4658 2287 4675
rect 3889 4673 3926 4676
rect 2278 4654 2281 4658
rect 4930 4656 5261 4676
rect 5296 4794 6075 4814
rect 1872 4612 1875 4638
rect 1901 4633 1904 4638
rect 1901 4616 1946 4633
rect 1901 4612 1904 4616
rect 1383 4591 1420 4595
rect 247 4456 1043 4496
rect 1151 4582 1420 4591
rect 2249 4583 2252 4588
rect 1151 4565 1946 4582
rect 2192 4566 2252 4583
rect 1151 4554 1420 4565
rect 2249 4562 2252 4566
rect 2278 4583 2281 4588
rect 2278 4566 2287 4583
rect 2278 4562 2281 4566
rect 4044 4565 4104 4582
rect 3831 4561 3870 4563
rect 1151 4543 1266 4554
rect 1151 4498 1262 4543
rect 1869 4520 1872 4546
rect 1898 4541 1901 4546
rect 1898 4524 1946 4541
rect 3831 4528 3834 4561
rect 3867 4553 3870 4561
rect 4044 4553 4061 4565
rect 3867 4536 4061 4553
rect 3867 4528 3870 4536
rect 3831 4526 3870 4528
rect 1898 4520 1901 4524
rect 1383 4498 1420 4502
rect 5296 4501 5316 4794
rect 6072 4791 6075 4794
rect 6101 4814 6104 4817
rect 6101 4794 6112 4814
rect 6101 4791 6104 4794
rect 6072 4790 6104 4791
rect 7936 4763 7994 4778
rect 7936 4760 7948 4763
rect 7936 4734 7945 4760
rect 7980 4734 7994 4763
rect 8038 4762 8096 4777
rect 8038 4761 8051 4762
rect 8038 4735 8047 4761
rect 7936 4731 7948 4734
rect 7980 4731 8000 4734
rect 7936 4715 8000 4731
rect 7976 4654 8000 4715
rect 8038 4730 8051 4735
rect 8083 4730 8096 4762
rect 8038 4714 8096 4730
rect 8320 4766 8367 4769
rect 8320 4723 8322 4766
rect 8365 4763 8367 4766
rect 10810 4764 10839 4765
rect 10810 4763 10840 4764
rect 11863 4763 11908 4765
rect 8365 4723 10813 4763
rect 8320 4720 10813 4723
rect 10839 4720 11909 4763
rect 10810 4719 10840 4720
rect 10810 4717 10839 4719
rect 11813 4652 11849 4653
rect 10428 4634 10458 4636
rect 11757 4634 11849 4652
rect 1151 4490 1420 4498
rect 2246 4491 2249 4496
rect 1151 4473 1946 4490
rect 2192 4474 2249 4491
rect 1151 4461 1420 4473
rect 2246 4470 2249 4474
rect 2275 4491 2278 4496
rect 2275 4474 2287 4491
rect 4926 4481 5316 4501
rect 5611 4614 5640 4632
rect 2275 4470 2278 4474
rect 1151 4457 1241 4461
rect 247 4395 374 4456
rect 290 4002 417 4090
rect 1151 4002 1188 4457
rect 1870 4428 1873 4454
rect 1899 4449 1902 4454
rect 1899 4432 1946 4449
rect 1899 4428 1902 4432
rect 3767 4401 3806 4402
rect 1299 4388 1948 4390
rect 290 3965 1188 4002
rect 1270 4371 1948 4388
rect 2310 4384 2313 4387
rect 1270 4353 1420 4371
rect 2189 4364 2313 4384
rect 2310 4361 2313 4364
rect 2339 4384 2342 4387
rect 2339 4364 2352 4384
rect 3767 4368 3770 4401
rect 3803 4393 3806 4401
rect 4061 4393 4104 4410
rect 3803 4376 4124 4393
rect 3803 4368 3806 4376
rect 4061 4374 4078 4376
rect 3767 4367 3806 4368
rect 2339 4361 2342 4364
rect 1270 4294 1336 4353
rect 1383 4349 1420 4353
rect 1805 4326 1808 4352
rect 1834 4348 1837 4352
rect 1834 4329 1948 4348
rect 3703 4344 3742 4347
rect 1834 4326 1837 4329
rect 3703 4311 3706 4344
rect 3739 4336 3742 4344
rect 3739 4319 4124 4336
rect 5611 4330 5629 4614
rect 10427 4592 10430 4634
rect 10456 4624 11849 4634
rect 10456 4592 11853 4624
rect 10428 4590 10458 4592
rect 11757 4558 11853 4592
rect 8046 4416 8106 4427
rect 8046 4382 8059 4416
rect 8093 4382 8106 4416
rect 8406 4410 8929 4433
rect 8966 4410 9881 4433
rect 11763 4415 11853 4558
rect 8046 4371 8106 4382
rect 9852 4400 9881 4410
rect 10650 4400 10764 4408
rect 9852 4388 10764 4400
rect 9852 4380 10685 4388
rect 9852 4379 9881 4380
rect 3739 4311 3742 4319
rect 5534 4313 5629 4330
rect 8407 4328 8929 4350
rect 8966 4328 9787 4350
rect 3703 4309 3742 4311
rect 1270 4275 1948 4294
rect 2311 4288 2314 4291
rect 1270 4257 1420 4275
rect 2189 4268 2314 4288
rect 2311 4265 2314 4268
rect 2340 4288 2343 4291
rect 2340 4268 2352 4288
rect 4968 4270 4988 4282
rect 2340 4265 2343 4268
rect 1270 4256 1337 4257
rect 1270 4252 1336 4256
rect 1383 4253 1420 4257
rect 290 3902 417 3965
rect 284 3526 411 3615
rect 1270 3526 1307 4252
rect 1801 4230 1804 4256
rect 1830 4252 1833 4256
rect 1830 4233 1948 4252
rect 4968 4250 5003 4270
rect 4968 4248 4988 4250
rect 1830 4230 1833 4233
rect 4930 4228 4988 4248
rect 284 3489 1307 3526
rect 1383 4179 1948 4198
rect 2310 4192 2313 4195
rect 284 3427 411 3489
rect 290 3042 417 3133
rect 1383 3042 1420 4179
rect 2189 4172 2313 4192
rect 2310 4169 2313 4172
rect 2339 4192 2342 4195
rect 2339 4172 2352 4192
rect 3642 4187 3681 4189
rect 2339 4169 2342 4172
rect 1805 4134 1808 4160
rect 1834 4156 1837 4160
rect 1834 4137 1948 4156
rect 3642 4154 3645 4187
rect 3678 4179 3681 4187
rect 3678 4162 4124 4179
rect 3678 4154 3681 4162
rect 3642 4152 3681 4154
rect 4069 4146 4104 4162
rect 1834 4134 1837 4137
rect 4963 4128 5000 4148
rect 4963 4073 4983 4128
rect 5567 4125 5640 4143
rect 9765 4140 9787 4328
rect 10027 4312 10073 4315
rect 10027 4272 10030 4312
rect 10070 4302 10073 4312
rect 10658 4302 10764 4310
rect 10070 4290 10764 4302
rect 11200 4290 11372 4310
rect 10070 4282 10685 4290
rect 11200 4282 11371 4290
rect 10070 4272 10073 4282
rect 10027 4270 10073 4272
rect 10128 4244 10164 4247
rect 11351 4237 11371 4282
rect 10164 4217 10764 4237
rect 11200 4217 11371 4237
rect 10128 4205 10164 4208
rect 9765 4139 9925 4140
rect 5567 4104 5585 4125
rect 9765 4119 10764 4139
rect 9765 4118 9925 4119
rect 11351 4112 11371 4217
rect 11760 4112 11850 4179
rect 6237 4109 6268 4110
rect 5528 4086 5585 4104
rect 6236 4108 6269 4109
rect 6236 4103 6239 4108
rect 6201 4098 6239 4103
rect 5878 4081 6239 4098
rect 6266 4081 6269 4108
rect 8484 4082 8929 4098
rect 5878 4076 6268 4081
rect 8481 4078 8929 4082
rect 8966 4088 10685 4098
rect 8966 4078 10764 4088
rect 4930 4053 4983 4073
rect 7940 4069 7996 4078
rect 3579 4034 3621 4035
rect 3579 4001 3582 4034
rect 3615 4026 3621 4034
rect 7940 4034 7952 4069
rect 7985 4034 7996 4069
rect 3615 4009 4069 4026
rect 3615 4001 3621 4009
rect 3579 4000 3621 4001
rect 4052 3991 4069 4009
rect 5577 4010 5632 4028
rect 7940 4024 7996 4034
rect 5577 4008 5595 4010
rect 5535 3992 5595 4008
rect 4052 3974 4104 3991
rect 4966 3917 4998 3961
rect 4966 3898 4986 3917
rect 4930 3878 4986 3898
rect 3523 3877 3562 3878
rect 3523 3844 3526 3877
rect 3559 3869 3562 3877
rect 3559 3852 4060 3869
rect 3559 3844 3562 3852
rect 3523 3843 3562 3844
rect 4044 3841 4060 3852
rect 4044 3811 4061 3841
rect 8481 3830 8504 4078
rect 10655 4068 10764 4078
rect 11351 4069 11850 4112
rect 10220 4011 10259 4013
rect 10219 4010 10260 4011
rect 10219 3971 10220 4010
rect 10259 4000 10260 4010
rect 11351 4000 11371 4069
rect 10259 3990 10685 4000
rect 10259 3980 10764 3990
rect 10259 3971 10260 3980
rect 10219 3970 10260 3971
rect 10662 3970 10764 3980
rect 11200 3970 11371 4000
rect 11760 3970 11850 4069
rect 10220 3968 10259 3970
rect 10302 3941 10342 3942
rect 10300 3915 10303 3941
rect 10341 3935 10344 3941
rect 11351 3935 11371 3970
rect 10341 3917 10685 3935
rect 11200 3917 11371 3935
rect 10341 3915 10764 3917
rect 10302 3914 10342 3915
rect 10650 3897 10764 3915
rect 11194 3903 11371 3917
rect 11194 3897 11370 3903
rect 4044 3794 4104 3811
rect 4959 3805 4997 3823
rect 8044 3813 8106 3822
rect 4959 3723 4977 3805
rect 5533 3760 5605 3778
rect 8044 3777 8061 3813
rect 8095 3777 8106 3813
rect 8406 3807 8504 3830
rect 8565 3817 8929 3837
rect 8966 3819 10685 3837
rect 8966 3817 10764 3819
rect 8044 3769 8106 3777
rect 4930 3703 4978 3723
rect 5587 3541 5605 3760
rect 8565 3747 8585 3817
rect 10659 3799 10764 3817
rect 8407 3732 8585 3747
rect 8407 3725 8582 3732
rect 11486 3561 11564 3564
rect 5587 3523 5641 3541
rect 11486 3490 11489 3561
rect 11560 3549 11564 3561
rect 11760 3549 11850 3641
rect 11560 3502 11850 3549
rect 11560 3490 11564 3502
rect 11486 3487 11564 3490
rect 8682 3452 8728 3454
rect 5901 3447 5933 3448
rect 8682 3447 8687 3452
rect 5901 3445 8687 3447
rect 5901 3417 5903 3445
rect 5931 3419 8687 3445
rect 5931 3417 5933 3419
rect 5901 3414 5933 3417
rect 8682 3415 8687 3419
rect 8724 3415 8728 3452
rect 11760 3432 11850 3502
rect 8682 3413 8728 3415
rect 8761 3393 8804 3395
rect 8761 3387 8764 3393
rect 7635 3386 8764 3387
rect 7635 3360 7638 3386
rect 7664 3361 8764 3386
rect 7664 3360 7667 3361
rect 8761 3356 8764 3361
rect 8801 3356 8804 3393
rect 8761 3354 8804 3356
rect 3462 3330 3499 3334
rect 3462 3297 3464 3330
rect 3497 3322 3499 3330
rect 3497 3305 4094 3322
rect 3497 3297 3499 3305
rect 3462 3294 3499 3297
rect 5579 3281 5597 3282
rect 5545 3270 5597 3281
rect 5545 3263 5780 3270
rect 5579 3252 5780 3263
rect 4937 3215 4997 3235
rect 3398 3171 3437 3172
rect 3398 3138 3401 3171
rect 3434 3163 3437 3171
rect 3434 3151 4094 3163
rect 8835 3160 8879 3162
rect 3434 3146 4104 3151
rect 8835 3150 8838 3160
rect 3434 3138 3437 3146
rect 3398 3137 3437 3138
rect 4065 3134 4104 3146
rect 8822 3132 8838 3150
rect 8834 3123 8838 3132
rect 8875 3123 8879 3160
rect 8834 3122 8879 3123
rect 8834 3116 8874 3122
rect 7751 3098 8874 3116
rect 4957 3095 4995 3096
rect 4955 3078 4995 3095
rect 4955 3060 4975 3078
rect 290 3005 1420 3042
rect 4930 3040 4975 3060
rect 5553 3057 5786 3073
rect 5531 3055 5786 3057
rect 5531 3039 5571 3055
rect 9488 3052 9548 3056
rect 290 2945 417 3005
rect 3336 2983 3339 3016
rect 3372 3008 3375 3016
rect 3372 2991 4054 3008
rect 9488 3002 9491 3052
rect 9541 3050 9548 3052
rect 11760 3050 11850 3153
rect 9541 3003 11850 3050
rect 9541 3002 9548 3003
rect 9488 2998 9548 3002
rect 3372 2983 3375 2991
rect 4039 2984 4054 2991
rect 4039 2973 4056 2984
rect 4039 2956 4104 2973
rect 5533 2960 5573 2961
rect 5533 2946 5574 2960
rect 5533 2945 5784 2946
rect 5556 2928 5784 2945
rect 11760 2944 11850 3003
rect 4950 2900 4995 2913
rect 4950 2885 4999 2900
rect 4930 2880 4999 2885
rect 3275 2868 3317 2869
rect 3275 2835 3279 2868
rect 3312 2860 3317 2868
rect 4930 2865 4985 2880
rect 3312 2843 4056 2860
rect 3312 2835 3317 2843
rect 3275 2833 3317 2835
rect 4039 2794 4056 2843
rect 4039 2777 4104 2794
rect 4954 2758 4997 2781
rect 284 2627 411 2711
rect 4954 2710 4974 2758
rect 5552 2732 5782 2750
rect 5552 2731 5594 2732
rect 5531 2713 5594 2731
rect 4930 2690 4974 2710
rect 1801 2653 1832 2655
rect 1867 2653 1898 2655
rect 284 2590 1254 2627
rect 1801 2606 1804 2653
rect 1830 2606 1868 2653
rect 1894 2606 2533 2653
rect 1801 2604 1832 2606
rect 1867 2604 1898 2606
rect 284 2523 411 2590
rect 1217 2455 1254 2590
rect 2486 2538 2533 2606
rect 5163 2639 5194 2641
rect 8927 2639 8972 2642
rect 5163 2598 5166 2639
rect 5192 2598 8931 2639
rect 8968 2598 8972 2639
rect 5163 2596 5194 2598
rect 8927 2596 8972 2598
rect 11763 2538 11853 2635
rect 1668 2529 1694 2532
rect 2486 2530 11853 2538
rect 1873 2525 1876 2527
rect 1694 2506 1876 2525
rect 1668 2500 1694 2503
rect 1873 2501 1876 2506
rect 1902 2525 1905 2527
rect 2049 2525 2052 2529
rect 1902 2506 2052 2525
rect 1902 2501 1905 2506
rect 2049 2502 2052 2506
rect 2079 2502 2082 2529
rect 2486 2491 9383 2530
rect 1613 2463 1616 2489
rect 1642 2485 1645 2489
rect 1807 2485 1810 2491
rect 1642 2466 1810 2485
rect 1642 2463 1645 2466
rect 1807 2465 1810 2466
rect 1836 2485 1839 2491
rect 2099 2485 2102 2489
rect 1836 2466 2102 2485
rect 1836 2465 1839 2466
rect 2099 2463 2102 2466
rect 2128 2463 2131 2489
rect 9379 2483 9383 2491
rect 9433 2491 11853 2530
rect 9433 2483 9436 2491
rect 9379 2479 9436 2483
rect 1217 2454 1420 2455
rect 1217 2436 1442 2454
rect 1217 2430 1582 2436
rect 1217 2418 1715 2430
rect 2247 2429 2277 2431
rect 2246 2427 2249 2429
rect 1383 2414 1715 2418
rect 1420 2408 1715 2414
rect 683 2404 760 2408
rect 683 2338 688 2404
rect 754 2389 760 2404
rect 2024 2405 2249 2427
rect 1383 2389 1422 2391
rect 754 2385 1422 2389
rect 754 2364 1714 2385
rect 754 2352 1421 2364
rect 2024 2361 2046 2405
rect 2246 2403 2249 2405
rect 2275 2403 2278 2429
rect 11763 2426 11853 2491
rect 2247 2401 2277 2403
rect 4058 2397 4100 2414
rect 4058 2387 4096 2397
rect 4058 2365 4086 2387
rect 754 2338 760 2352
rect 1383 2350 1420 2352
rect 3211 2351 3252 2353
rect 683 2334 760 2338
rect 3211 2318 3215 2351
rect 3248 2343 3252 2351
rect 4058 2343 4085 2365
rect 3248 2326 4085 2343
rect 5534 2337 5565 2355
rect 3248 2318 3252 2326
rect 4058 2325 4075 2326
rect 3211 2317 3252 2318
rect 2185 2314 2214 2316
rect 2184 2310 2187 2314
rect 290 2224 417 2301
rect 2027 2291 2187 2310
rect 2184 2288 2187 2291
rect 2213 2288 2216 2314
rect 4926 2309 4987 2329
rect 5547 2319 5782 2337
rect 4967 2305 4987 2309
rect 2185 2286 2214 2288
rect 4967 2285 5009 2305
rect 5611 2256 5728 2271
rect 5605 2252 5633 2256
rect 290 2187 889 2224
rect 4052 2221 4100 2238
rect 5605 2226 5606 2252
rect 5632 2226 5633 2252
rect 7591 2245 7594 2250
rect 7113 2229 7594 2245
rect 5605 2223 5633 2226
rect 7591 2224 7594 2229
rect 7620 2224 7623 2250
rect 290 2113 417 2187
rect 852 2021 889 2187
rect 3145 2194 3184 2197
rect 3145 2161 3148 2194
rect 3181 2186 3184 2194
rect 4052 2192 4069 2221
rect 4052 2186 4068 2192
rect 3181 2170 4068 2186
rect 3181 2169 4033 2170
rect 3181 2161 3184 2169
rect 3145 2159 3184 2161
rect 4966 2154 4998 2170
rect 4926 2134 4998 2154
rect 7539 2152 7542 2157
rect 5545 2129 5724 2142
rect 7113 2136 7542 2152
rect 7539 2131 7542 2136
rect 7568 2131 7571 2157
rect 5531 2124 5724 2129
rect 5531 2109 5563 2124
rect 5531 2101 5549 2109
rect 1616 2098 1645 2099
rect 1615 2072 1618 2098
rect 1644 2096 1647 2098
rect 1644 2074 1715 2096
rect 1644 2072 1647 2074
rect 1616 2070 1645 2072
rect 2142 2053 2174 2055
rect 2142 2050 2145 2053
rect 2025 2029 2145 2050
rect 2142 2027 2145 2029
rect 2171 2027 2174 2053
rect 4044 2040 4100 2057
rect 4044 2036 4061 2040
rect 2142 2025 2174 2027
rect 3084 2032 3121 2033
rect 4044 2032 4060 2036
rect 3084 2030 4060 2032
rect 852 2003 1447 2021
rect 852 1996 1454 2003
rect 1593 1996 1715 1997
rect 2311 1996 2340 1998
rect 3084 1997 3086 2030
rect 3119 2015 4060 2030
rect 5536 2018 5556 2034
rect 3119 1997 3121 2015
rect 852 1984 1715 1996
rect 2310 1993 2313 1996
rect 1383 1980 1715 1984
rect 1419 1975 1715 1980
rect 2025 1972 2313 1993
rect 1206 1923 1247 1925
rect 1383 1923 1582 1925
rect 290 1810 417 1892
rect 1206 1886 1209 1923
rect 1246 1919 1582 1923
rect 1246 1897 1715 1919
rect 1246 1886 1421 1897
rect 2025 1890 2046 1972
rect 2310 1970 2313 1972
rect 2339 1970 2342 1996
rect 3084 1994 3121 1997
rect 5538 2013 5556 2018
rect 9267 2014 9322 2015
rect 5538 1995 5727 2013
rect 4926 1977 4995 1979
rect 2311 1968 2340 1970
rect 4926 1959 5003 1977
rect 4974 1950 5003 1959
rect 5666 1974 5698 1976
rect 5666 1948 5669 1974
rect 5695 1972 5698 1974
rect 5695 1951 5727 1972
rect 7492 1968 7495 1973
rect 7113 1952 7495 1968
rect 5695 1948 5712 1951
rect 5666 1944 5712 1948
rect 7492 1947 7495 1952
rect 7521 1947 7524 1973
rect 9267 1964 9270 2014
rect 9320 2012 9323 2014
rect 11760 2012 11850 2127
rect 9320 1965 11850 2012
rect 9320 1964 9323 1965
rect 9267 1962 9322 1964
rect 11760 1918 11850 1965
rect 3015 1886 3054 1888
rect 1206 1884 1247 1886
rect 1383 1884 1420 1886
rect 3015 1853 3018 1886
rect 3051 1878 3054 1886
rect 4035 1878 4100 1885
rect 3051 1868 4100 1878
rect 7442 1875 7445 1880
rect 3051 1861 4064 1868
rect 4972 1862 5002 1866
rect 3051 1853 3054 1861
rect 4047 1859 4064 1861
rect 3015 1851 3054 1853
rect 4971 1838 5002 1862
rect 7113 1859 7445 1875
rect 7442 1854 7445 1859
rect 7471 1854 7474 1880
rect 683 1818 763 1824
rect 683 1810 692 1818
rect 290 1760 692 1810
rect 290 1704 417 1760
rect 683 1752 692 1760
rect 758 1752 763 1818
rect 4971 1804 4991 1838
rect 5562 1804 5725 1817
rect 4926 1784 4991 1804
rect 5531 1799 5725 1804
rect 5531 1786 5580 1799
rect 683 1747 763 1752
rect 5709 1747 5741 1763
rect 5606 1743 5638 1744
rect 4945 1713 4948 1739
rect 4974 1734 4977 1739
rect 5606 1734 5609 1743
rect 4974 1718 5609 1734
rect 4974 1713 4977 1718
rect 5606 1717 5609 1718
rect 5635 1717 5638 1743
rect 5606 1716 5638 1717
rect 5709 1742 6074 1747
rect 5709 1716 5712 1742
rect 5738 1734 6074 1742
rect 6771 1744 6812 1745
rect 6771 1734 6774 1744
rect 5738 1718 6774 1734
rect 5738 1716 5741 1718
rect 5709 1715 5741 1716
rect 6066 1711 6774 1718
rect 5665 1710 5693 1711
rect 4892 1705 4925 1707
rect 4891 1676 4894 1705
rect 4923 1697 4926 1705
rect 5466 1702 5498 1703
rect 5466 1697 5469 1702
rect 4923 1681 5469 1697
rect 4923 1676 4926 1681
rect 5466 1676 5469 1681
rect 5495 1676 5498 1702
rect 5663 1701 5666 1710
rect 5660 1685 5666 1701
rect 5663 1684 5666 1685
rect 5692 1701 5695 1710
rect 6771 1709 6774 1711
rect 6809 1709 6812 1744
rect 6771 1708 6812 1709
rect 9786 1736 9842 1738
rect 5887 1701 5890 1704
rect 5692 1685 5890 1701
rect 5692 1684 5695 1685
rect 5665 1683 5693 1684
rect 5887 1678 5890 1685
rect 5916 1678 5919 1704
rect 9786 1686 9789 1736
rect 9839 1731 9842 1736
rect 11058 1736 11126 1737
rect 11058 1731 11069 1736
rect 9839 1690 11069 1731
rect 9839 1686 9842 1690
rect 9786 1685 9842 1686
rect 11058 1685 11069 1690
rect 11120 1731 11126 1736
rect 11811 1731 11877 1795
rect 11120 1690 11877 1731
rect 11120 1685 11126 1690
rect 11058 1684 11126 1685
rect 11811 1680 11877 1690
rect 5889 1677 5917 1678
rect 4891 1674 4926 1676
rect 6088 1662 6116 1665
rect 4449 1656 4482 1659
rect 4449 1625 4450 1656
rect 4481 1635 4482 1656
rect 5035 1648 5065 1649
rect 5034 1635 5037 1648
rect 4481 1625 5037 1635
rect 4449 1622 5037 1625
rect 5063 1635 5066 1648
rect 6088 1636 6089 1662
rect 6115 1636 6116 1662
rect 6088 1635 6116 1636
rect 6491 1660 6521 1663
rect 6491 1635 6493 1660
rect 5063 1633 6493 1635
rect 6520 1633 6521 1660
rect 5063 1630 6520 1633
rect 5063 1622 6514 1630
rect 4449 1619 6514 1622
rect 4830 1597 4874 1598
rect 298 1596 4874 1597
rect 298 1555 4831 1596
rect 4145 1554 4193 1555
rect 4828 1554 4831 1555
rect 4873 1554 4876 1596
rect 5767 1586 5805 1589
rect 7375 1588 7405 1590
rect 4830 1553 4874 1554
rect 5767 1553 5770 1586
rect 5803 1553 5805 1586
rect 5767 1550 5805 1553
rect 5882 1546 5885 1580
rect 5919 1546 5922 1580
rect 6741 1564 6807 1566
rect 6741 1532 6778 1564
rect 6804 1532 6807 1564
rect 7304 1554 7377 1588
rect 7403 1554 7406 1588
rect 7375 1552 7406 1554
rect 6741 1530 6807 1532
rect 296 1458 2189 1500
rect 2215 1488 4446 1500
rect 2215 1458 2614 1488
rect 2601 1417 2614 1458
rect 2672 1458 4446 1488
rect 4488 1458 4494 1500
rect 6916 1499 6961 1501
rect 4897 1481 4935 1484
rect 2672 1417 2684 1458
rect 4897 1449 4899 1481
rect 4931 1449 4935 1481
rect 6916 1461 6920 1499
rect 6958 1461 6961 1499
rect 6916 1458 6961 1461
rect 9162 1484 9222 1487
rect 4897 1446 4935 1449
rect 9162 1434 9165 1484
rect 9215 1482 9222 1484
rect 11803 1482 12013 1576
rect 9215 1435 12013 1482
rect 9215 1434 9222 1435
rect 9162 1431 9222 1434
rect 2601 1408 2684 1417
rect 284 1299 411 1377
rect 11803 1368 12013 1435
rect 11805 1367 11882 1368
rect 1207 1299 1248 1301
rect 284 1262 1208 1299
rect 1245 1262 1248 1299
rect 7589 1283 7592 1333
rect 7618 1283 13243 1333
rect 284 1189 411 1262
rect 1207 1260 1248 1262
rect 1960 1256 1989 1258
rect 2183 1256 2214 1258
rect 1959 1220 1962 1256
rect 1988 1220 2185 1256
rect 2211 1220 2214 1256
rect 12633 1243 12834 1245
rect 1960 1218 1989 1220
rect 2183 1218 2214 1220
rect 7535 1193 7538 1243
rect 7564 1193 12834 1243
rect 7488 1103 7491 1153
rect 7517 1151 12415 1153
rect 7517 1103 12426 1151
rect 7440 1013 7443 1063
rect 7469 1062 12019 1063
rect 7469 1013 12040 1062
rect 5299 1004 6389 1005
rect 5299 1002 5375 1004
rect 5298 974 5301 1002
rect 5329 977 5375 1002
rect 5329 974 5332 977
rect 5372 976 5375 977
rect 5403 1002 6389 1004
rect 5403 977 6282 1002
rect 5403 976 5406 977
rect 6279 974 6282 977
rect 6310 977 6389 1002
rect 6310 974 6313 977
rect 1379 960 1416 961
rect 290 878 417 948
rect 1247 922 1508 960
rect 4906 923 4956 924
rect 9499 923 9502 925
rect 1247 878 1285 922
rect 1379 920 1416 922
rect 4906 917 9502 923
rect 2246 890 2274 891
rect 290 840 1285 878
rect 1887 857 2247 890
rect 2273 857 2276 890
rect 4906 871 4909 917
rect 4955 877 9502 917
rect 4955 871 4958 877
rect 9499 875 9502 877
rect 9552 875 9555 925
rect 4906 869 4956 871
rect 2246 855 2274 857
rect 290 760 417 840
rect 5737 826 9445 832
rect 5737 822 9383 826
rect 5737 786 5747 822
rect 5744 776 5747 786
rect 5793 786 9383 822
rect 5793 776 5796 786
rect 9380 780 9383 786
rect 9433 786 9445 826
rect 9433 780 9436 786
rect 5881 739 9336 741
rect 5881 734 9270 739
rect 5880 733 9270 734
rect 1504 696 1507 725
rect 1536 722 1539 725
rect 2142 724 2175 728
rect 2141 722 2144 724
rect 1536 696 2144 722
rect 1508 695 2144 696
rect 2173 722 2176 724
rect 2173 695 2507 722
rect 1508 693 2507 695
rect 2142 691 2175 693
rect 1888 654 2122 659
rect 1888 599 2028 654
rect 2025 594 2028 599
rect 2088 625 2122 654
rect 2088 601 2126 625
rect 2088 599 2122 601
rect 2088 594 2091 599
rect 2025 592 2091 594
rect 2028 591 2088 592
rect 2477 485 2506 693
rect 5880 687 5890 733
rect 5936 695 9270 733
rect 5936 687 5945 695
rect 9267 693 9270 695
rect 9320 695 9336 739
rect 9320 693 9323 695
rect 5880 682 5945 687
rect 6725 647 6777 649
rect 9174 647 9177 648
rect 6725 642 9177 647
rect 6725 596 6729 642
rect 6775 602 9177 642
rect 9227 647 9230 648
rect 9227 602 9239 647
rect 6775 601 9239 602
rect 6775 596 6778 601
rect 6725 591 6777 596
rect 4119 485 4151 487
rect 9719 485 9835 488
rect 290 355 417 446
rect 2458 373 4122 485
rect 4148 483 9731 485
rect 4148 481 6240 483
rect 4148 479 5333 481
rect 4148 373 5259 479
rect 4119 371 4151 373
rect 5256 367 5259 373
rect 5445 373 6240 481
rect 5445 369 5448 373
rect 5371 367 5448 369
rect 5256 365 5448 367
rect 6237 364 6240 373
rect 6426 373 9731 483
rect 9825 373 9835 485
rect 6426 364 6430 373
rect 9719 370 9835 373
rect 6237 362 6430 364
rect 290 317 1287 355
rect 290 258 417 317
rect 1249 232 1287 317
rect 1379 232 1416 233
rect 1249 194 1521 232
rect 1379 192 1416 194
rect 2304 135 2335 137
rect 1881 101 2306 135
rect 2332 101 2335 135
rect 2304 99 2335 101
rect 411 46 461 51
rect 411 7 415 46
rect 454 40 461 46
rect 7308 43 7347 44
rect 7307 40 7310 43
rect 454 12 7310 40
rect 454 7 461 12
rect 7307 10 7310 12
rect 7343 10 7347 43
rect 7308 9 7347 10
rect 411 4 461 7
rect 3949 -23 3991 -22
rect 3949 -56 3954 -23
rect 3987 -48 7976 -23
rect 3987 -56 7977 -48
rect 3949 -57 3991 -56
rect 7373 -58 7977 -56
rect 3889 -85 3927 -84
rect 277 -296 404 -108
rect 3889 -118 3892 -85
rect 3925 -118 7569 -85
rect 3889 -119 3927 -118
rect 6962 -119 7569 -118
rect 3825 -148 3867 -147
rect 3825 -181 3829 -148
rect 3862 -181 7161 -148
rect 3825 -182 3867 -181
rect 3766 -211 3806 -210
rect 3766 -244 3769 -211
rect 3802 -212 3806 -211
rect 3802 -244 6760 -212
rect 3766 -245 6760 -244
rect 3766 -246 3806 -245
rect 3700 -279 3741 -278
rect 3699 -312 3705 -279
rect 3738 -312 6351 -279
rect 3700 -314 3741 -312
rect 3642 -341 3683 -340
rect 3642 -374 3645 -341
rect 3678 -343 5949 -341
rect 3678 -374 5950 -343
rect 3642 -375 3683 -374
rect 3582 -438 3585 -405
rect 3618 -406 3621 -405
rect 3618 -438 5551 -406
rect 3592 -439 5551 -438
rect 3010 -487 3064 -484
rect 3010 -488 3015 -487
rect 1727 -492 3015 -488
rect 1722 -530 3015 -492
rect 3058 -530 3064 -487
rect 3524 -495 3527 -462
rect 3560 -467 3563 -462
rect 3560 -495 5160 -467
rect 3550 -500 5160 -495
rect 1722 -531 3064 -530
rect 284 -771 411 -583
rect 1722 -719 1923 -531
rect 3010 -534 3064 -531
rect 3466 -564 3469 -531
rect 3502 -564 4740 -531
rect 3075 -566 3129 -565
rect 3075 -572 3080 -566
rect 2132 -609 3080 -572
rect 3123 -609 3129 -566
rect 4127 -594 4329 -592
rect 3411 -595 4332 -594
rect 2132 -615 3129 -609
rect 2132 -716 2330 -615
rect 3401 -628 3404 -595
rect 3437 -627 4332 -595
rect 3437 -628 3440 -627
rect 3143 -637 3192 -633
rect 3143 -653 3147 -637
rect 2582 -655 3147 -653
rect 2525 -677 3147 -655
rect 3187 -677 3192 -637
rect 2525 -683 3192 -677
rect 2525 -693 3183 -683
rect 3337 -693 3340 -659
rect 3373 -693 3935 -659
rect 2525 -716 2723 -693
rect 3126 -716 3191 -715
rect 1720 -785 1923 -719
rect 2127 -782 2330 -716
rect 2523 -782 2726 -716
rect 2923 -720 3191 -716
rect 2923 -771 3130 -720
rect 3181 -771 3191 -720
rect 3276 -718 3331 -716
rect 3276 -720 3531 -718
rect 3732 -719 3936 -693
rect 3276 -757 3282 -720
rect 3319 -757 3531 -720
rect 3276 -761 3531 -757
rect 2923 -779 3191 -771
rect 2923 -782 3126 -779
rect 3328 -784 3531 -761
rect 3731 -785 3936 -719
rect 4124 -782 4332 -627
rect 4535 -694 4738 -564
rect 4535 -723 4739 -694
rect 4536 -784 4739 -723
rect 4953 -782 5156 -500
rect 5352 -710 5551 -439
rect 5351 -785 5554 -710
rect 5750 -712 5950 -374
rect 5747 -782 5950 -712
rect 6160 -719 6351 -312
rect 6564 -717 6759 -245
rect 6962 -717 7161 -181
rect 7373 -151 7569 -119
rect 7783 -108 7977 -58
rect 10035 -69 10078 -67
rect 8185 -72 8381 -69
rect 10033 -72 10036 -69
rect 8185 -107 10036 -72
rect 7373 -717 7568 -151
rect 7783 -715 7976 -108
rect 6152 -784 6355 -719
rect 6559 -782 6762 -717
rect 6962 -782 7165 -717
rect 7367 -782 7570 -717
rect 7774 -793 7977 -715
rect 8185 -717 8381 -107
rect 10033 -109 10036 -107
rect 10076 -109 10079 -69
rect 10035 -110 10078 -109
rect 10125 -150 10168 -148
rect 10124 -151 10127 -150
rect 8578 -189 10127 -151
rect 10166 -189 10169 -150
rect 8182 -782 8385 -717
rect 8578 -719 8774 -189
rect 10125 -191 10168 -189
rect 10217 -233 10220 -232
rect 8993 -271 10220 -233
rect 10259 -271 10262 -232
rect 8993 -717 9191 -271
rect 10301 -312 10343 -309
rect 9404 -350 10302 -312
rect 10340 -350 10343 -312
rect 8577 -784 8780 -719
rect 8989 -782 9192 -717
rect 9404 -720 9602 -350
rect 10301 -353 10343 -350
rect 9911 -649 10535 -629
rect 9911 -717 9931 -649
rect 10627 -670 10647 -629
rect 10404 -690 10647 -670
rect 10404 -717 10424 -690
rect 10724 -717 10745 -628
rect 9403 -785 9606 -720
rect 9802 -782 10005 -717
rect 10204 -747 10424 -717
rect 10204 -782 10407 -747
rect 10612 -782 10815 -717
rect 10917 -726 10938 -628
rect 11014 -647 11033 -630
rect 11014 -666 11514 -647
rect 11495 -712 11514 -666
rect 11030 -726 11233 -717
rect 11495 -719 11598 -712
rect 11839 -717 12040 1013
rect 10917 -747 11233 -726
rect 11030 -782 11233 -747
rect 11428 -784 11631 -719
rect 11833 -769 12040 -717
rect 12225 -717 12426 1103
rect 11833 -782 12036 -769
rect 12225 -782 12432 -717
rect 12633 -719 12834 1193
rect 13042 -717 13243 1283
rect 12225 -786 12426 -782
rect 12633 -784 12837 -719
rect 13039 -775 13243 -717
rect 13039 -782 13242 -775
rect 12633 -792 12834 -784
<< via2 >>
rect 7948 4760 7980 4763
rect 7948 4734 7971 4760
rect 7971 4734 7980 4760
rect 8051 4761 8083 4762
rect 8051 4735 8073 4761
rect 8073 4735 8083 4761
rect 7948 4731 7980 4734
rect 8051 4730 8083 4735
rect 8059 4382 8093 4416
rect 7952 4034 7985 4069
rect 8061 3777 8095 3813
<< metal3 >>
rect 7941 4763 7986 4769
rect 7941 4731 7948 4763
rect 7980 4731 7986 4763
rect 7941 4694 7986 4731
rect 8045 4762 8090 4768
rect 8045 4730 8051 4762
rect 8083 4730 8090 4762
rect 7941 4078 7978 4694
rect 8045 4693 8090 4730
rect 8053 4429 8090 4693
rect 8053 4416 8097 4429
rect 8053 4382 8059 4416
rect 8093 4382 8097 4416
rect 8053 4369 8097 4382
rect 7941 4069 7990 4078
rect 7941 4045 7952 4069
rect 7946 4034 7952 4045
rect 7985 4034 7990 4069
rect 7946 4029 7990 4034
rect 8053 3858 8090 4369
rect 8052 3813 8099 3858
rect 8052 3777 8061 3813
rect 8095 3777 8099 3813
rect 8052 3771 8099 3777
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_0
timestamp 1629420194
transform -1 0 2012 0 -1 1081
box 64 419 528 1018
use sky130_hilas_nFETLarge  sky130_hilas_nFETLarge_0
timestamp 1629420194
transform -1 0 2008 0 -1 1836
box 64 420 501 1003
use sky130_hilas_DAC5bit01  sky130_hilas_DAC5bit01_0
timestamp 1629420194
transform 0 1 9912 1 0 -1031
box 382 524 2040 1123
use sky130_hilas_Trans2med  sky130_hilas_Trans2med_0
timestamp 1629420194
transform 1 0 2073 0 -1 2311
box -380 -143 -27 452
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_3
timestamp 1629420194
transform -1 0 6602 0 -1 2371
box 1050 -28 1622 631
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_2
timestamp 1629420194
transform -1 0 6599 0 -1 3298
box 1050 -28 1622 631
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_3
timestamp 1629420194
transform -1 0 4923 0 -1 2334
box -30 -106 840 594
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_2
timestamp 1629420194
transform -1 0 4927 0 -1 3240
box -30 -106 840 594
use sky130_hilas_WTA4Stage01  sky130_hilas_WTA4Stage01_0
timestamp 1629420194
transform 1 0 6825 0 1 1804
box -1121 -61 296 589
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_1
timestamp 1629420194
transform 1 0 4824 0 1 606
box 64 419 528 1018
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_2
timestamp 1629420194
transform -1 0 5880 0 1 606
box 64 419 528 1018
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_3
timestamp 1629420194
transform 1 0 5805 0 1 609
box 64 419 528 1018
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_4
timestamp 1629420194
transform -1 0 6861 0 1 609
box 64 419 528 1018
use sky130_hilas_nFETLarge  sky130_hilas_nFETLarge_1
timestamp 1629420194
transform -1 0 7435 0 1 608
box 64 420 501 1003
use sky130_hilas_Trans4small  sky130_hilas_Trans4small_0
timestamp 1629420194
transform 1 0 1738 0 1 4259
box 191 -150 471 455
use sky130_hilas_TA2Cell_1FG_Strong  sky130_hilas_TA2Cell_1FG_Strong_0
timestamp 1629420194
transform 1 0 8236 0 1 3936
box -2617 135 193 828
use sky130_hilas_TA2Cell_1FG  sky130_hilas_TA2Cell_1FG_0
timestamp 1629420194
transform 1 0 8236 0 1 3333
box -2616 135 193 828
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_1
timestamp 1629420194
transform -1 0 6601 0 -1 4345
box 1050 -28 1622 631
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_1
timestamp 1629420194
transform -1 0 4927 0 -1 4253
box -30 -106 840 594
use sky130_hilas_swc4x2cell  sky130_hilas_swc4x2cell_0
timestamp 1629420194
transform 1 0 6765 0 1 2702
box -1004 -26 1008 624
use sky130_hilas_Tgate4Single01  sky130_hilas_Tgate4Single01_0
timestamp 1629420194
transform 1 0 10780 0 1 3947
box -36 -164 440 477
use sky130_hilas_FGcharacterization01  sky130_hilas_FGcharacterization01_0
timestamp 1629420194
transform -1 0 2682 0 1 5308
box -912 259 2083 864
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_0
timestamp 1629420194
transform -1 0 4927 0 1 4476
box -30 -106 840 594
<< labels >>
rlabel metal2 13039 -782 13242 -717 1 DIG24 
port 1 n
rlabel metal2 12634 -784 12837 -719 0 DIG23
port 2 nsew
rlabel metal2 12229 -782 12432 -717 0 DIG22
port 3 nsew
rlabel metal2 11833 -782 12036 -717 0 DIG21
port 4 nsew
rlabel metal2 11428 -784 11631 -719 0 DIG29
port 5 nsew
rlabel metal2 11030 -782 11233 -717 0 DIG28
port 6 nsew
rlabel metal2 10612 -782 10815 -717 0 DIG27
port 7 nsew
rlabel metal2 10204 -782 10407 -717 0 DIG26
port 8 nsew
rlabel metal2 9802 -782 10005 -717 0 DIG25
port 9 nsew
rlabel metal2 9403 -785 9606 -720 0 DIG20
port 10 nsew
rlabel metal2 8989 -782 9192 -717 0 DIG19
port 11 nsew
rlabel metal2 8577 -784 8780 -719 0 DIG18
port 12 nsew
rlabel metal2 8182 -782 8385 -717 0 DIG17
port 13 nsew
rlabel metal2 7774 -780 7977 -715 0 DIG16
port 14 nsew
rlabel metal2 7367 -782 7570 -717 0 DIG15
port 15 nsew
rlabel metal2 6962 -782 7165 -717 0 DIG14
port 16 nsew
rlabel metal2 6559 -782 6762 -717 0 DIG13
port 17 nsew
rlabel metal2 6152 -784 6355 -719 0 DIG12
port 18 nsew
rlabel metal2 5747 -778 5950 -712 0 DIG11
port 19 nsew
rlabel metal2 5351 -776 5554 -710 0 DIG10
port 20 nsew
rlabel metal2 4953 -782 5156 -716 0 DIG09
port 21 nsew
rlabel metal2 4536 -784 4739 -718 0 DIG08
port 22 nsew
rlabel metal2 4127 -782 4330 -716 0 DIG07
port 23 nsew
rlabel metal2 3731 -785 3934 -719 0 DIG06
port 24 nsew
rlabel metal2 3328 -784 3531 -718 0 DIG05
port 25 nsew
rlabel metal2 2923 -782 3126 -716 0 DIG04
port 26 nsew
rlabel metal2 2523 -782 2726 -716 0 DIG03
port 27 nsew
rlabel metal2 2127 -782 2330 -716 0 DIG02
port 28 nsew
rlabel metal2 1720 -785 1923 -719 0 DIG01
port 29 nsew
rlabel metal2 11805 1367 11882 1576 0 CAP2    
port 30 nsew
rlabel metal2 11760 1918 11850 2127 0 GENERALGATE01   
port 31 nsew
rlabel metal2 11763 2426 11853 2635 0 GATEANDCAP1    
port 32 nsew
rlabel metal2 11760 2944 11850 3153 0 GENERALGATE02
port 33 nsew
rlabel metal2 11760 3432 11850 3641 0 OUTPUTTA1    
port 34 nsew
rlabel metal2 11760 3970 11850 4179 0 GATENFET1   
port 35 nsew
rlabel metal2 11763 4415 11853 4624 0 DACOUTPUT  
port 36 nsew
rlabel metal2 11764 4853 11850 5063 0 DRAINOUT
port 37 nsew
rlabel metal2 11764 5292 11850 5502 0 ROWTERM2
port 38 nsew
rlabel metal2 11767 5701 11853 5911 0 COLUMN2
port 39 nsew
rlabel metal2 11767 6114 11853 6324 0 COLUMN1
port 40 nsew
rlabel metal1 10273 6287 10592 6399 0 GATE2
port 41 nsew
rlabel metal1 7416 6284 7735 6396 0 GATE1
port 61 nsew
rlabel metal1 4557 6285 4876 6397 0 DRAININJECT
port 42 nsew
rlabel metal1 3026 6238 3160 6339 0 VTUN
port 43 nsew
rlabel metal2 295 6136 363 6368 0 VREFCHAR
port 44 nsew
rlabel metal2 295 5683 363 5915 0 CHAROUTPUT
port 45 nsew
rlabel metal2 250 5236 318 5468 0 LARGECAPACITOR
port 46 nsew
rlabel metal2 1379 920 1416 961 0 DRAIN6N
port 47 nsew
rlabel metal2 1379 192 1416 233 0 DRAIN6P
port 48 nsew
rlabel metal2 1383 1884 1420 1925 0 DRAIN5P
port 49 nsew
rlabel metal2 1383 1980 1420 2021 0 DARIN4P
port 50 nsew
rlabel metal2 1383 2350 1420 2391 0 DRAIN5N
port 51 nsew
rlabel metal2 1383 2414 1420 2455 0 DRAIN4N
port 52 nsew
rlabel metal2 1383 4157 1420 4198 0 DRAIN3P
port 53 nsew
rlabel metal2 1383 4253 1420 4294 0 DRAIN2P
port 54 nsew
rlabel metal2 1383 4349 1420 4390 0 DRAIN1P
port 55 nsew
rlabel metal2 1383 4461 1420 4502 0 DRAIN3N
port 56 nsew
rlabel metal2 1383 4554 1420 4595 0 DRAIN2N
port 57 nsew
rlabel metal2 1383 4657 1420 4698 0 DRAIN1N
port 58 nsew
rlabel metal2 1353 4765 1383 4805 0 SOURCEN
port 59 nsew
rlabel metal2 1353 4847 1383 4887 0 SOURCEP
port 60 nsew
rlabel metal2 279 5546 324 5586 0 VGND
port 63 nsew
rlabel metal2 283 5987 328 6027 0 VINJ
port 62 nsew
rlabel metal2 250 5157 301 5198 0 VINJ
port 62 nsew
rlabel metal2 246 5067 297 5108 0 VGND
port 63 nsew
rlabel metal2 298 1555 361 1597 0 VINJ
port 62 nsew
rlabel metal2 296 1458 359 1500 0 VGND
port 63 nsew
rlabel metal2 11863 4720 11908 4765 0 VPWR
port 64 nsew
rlabel metal1 5638 6371 5711 6401 0 VINJ
port 62 nsew
rlabel metal1 6154 6380 6251 6401 0 VGND
port 63 nsew
rlabel metal2 11811 1680 11877 1795 0 VPWR
port 64 nsew
rlabel metal1 5200 -785 5292 -712 0 VPWR
port 64 nsew
rlabel metal1 6393 -785 6485 -712 0 VPWR
port 64 nsew
<< end >>
