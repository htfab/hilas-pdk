magic
tech sky130A
magscale 1 2
timestamp 1632256356
<< checkpaint >>
rect -1260 1300 9440 5924
rect 5842 618 9078 1300
<< error_s >>
rect 290 4334 300 4362
rect 7880 4354 7890 4362
rect 7880 4334 8008 4354
rect 7880 4323 7891 4334
rect 1156 3768 1194 3796
rect 6516 3780 7178 3946
rect 7910 3820 7922 3890
rect 7938 3820 7950 3862
rect 7752 3808 7852 3820
rect 7896 3808 7996 3820
rect 7910 3796 7922 3808
rect 6986 3778 7024 3780
rect 6986 3772 7154 3778
rect 7684 3736 7752 3780
rect 7852 3736 7896 3780
rect 7938 3768 7950 3808
rect 7996 3736 8064 3780
rect 7696 3726 7720 3728
rect 7752 3726 7852 3736
rect 7896 3726 7996 3736
rect 184 3708 284 3726
rect 328 3720 428 3726
rect 184 3704 242 3708
rect 130 3620 170 3656
rect 196 3606 242 3704
rect 328 3692 478 3720
rect 7696 3710 8066 3726
rect 330 3690 478 3692
rect 330 3688 432 3690
rect 7702 3688 8066 3710
rect 330 3674 336 3688
rect 7702 3674 7746 3688
rect 7844 3682 8066 3688
rect 7844 3674 7850 3682
rect 7938 3674 7984 3682
rect 116 3592 172 3606
rect 114 3524 172 3574
rect 274 3524 336 3674
rect 434 3544 478 3674
rect 7702 3634 7748 3674
rect 2820 3542 2824 3562
rect 7702 3544 7746 3634
rect 274 3506 330 3524
rect 2854 3512 2858 3542
rect 7844 3524 7906 3674
rect 7960 3656 8066 3674
rect 8010 3620 8066 3656
rect 7938 3572 7984 3574
rect 7930 3524 7984 3572
rect 8008 3524 8066 3574
rect 7808 3506 7906 3524
rect 180 3446 250 3506
rect 274 3438 290 3506
rect 7890 3454 7906 3506
rect 7918 3496 8008 3506
rect 7930 3462 8008 3496
rect 7930 3454 8000 3462
rect 534 3240 712 3364
rect 1198 3228 1262 3236
rect 1220 3200 1272 3208
rect 1794 3006 2190 3172
rect 3012 3016 3256 3400
rect 4924 3018 5168 3400
rect 7468 3240 8130 3454
rect 6918 3228 6982 3236
rect 6908 3200 7010 3208
rect 1794 3004 2062 3006
rect 1794 2906 1808 3004
rect 1948 2994 1986 3004
rect 3012 2988 3290 3016
rect 3488 2988 3534 3016
rect 4646 2988 4692 3016
rect 4890 2990 5168 3018
rect 6194 2990 6232 3018
rect 6386 3006 6680 3172
rect 7156 3058 7412 3138
rect 7622 3110 7666 3200
rect 7822 3196 7834 3206
rect 7788 3154 7800 3188
rect 7822 3162 7888 3196
rect 7788 3138 7806 3154
rect 7468 3072 7666 3110
rect 7440 3066 7666 3072
rect 7778 3070 7800 3098
rect 7748 3066 7800 3070
rect 7440 3064 7800 3066
rect 7440 3058 7666 3064
rect 2448 2952 2494 2974
rect 3012 2952 3256 2988
rect 1842 2936 3336 2952
rect 3012 2924 3256 2936
rect 1814 2908 3308 2924
rect 1808 2870 1962 2906
rect 2808 2880 2926 2892
rect 2836 2852 2898 2864
rect 2826 2810 2830 2838
rect 2890 2810 2898 2846
rect 196 2778 250 2806
rect 196 2756 242 2778
rect 130 2694 170 2730
rect 274 2676 336 2806
rect 2826 2804 2832 2810
rect 2860 2798 2898 2810
rect 434 2676 478 2786
rect 2860 2776 2890 2798
rect 2918 2776 2926 2818
rect 3012 2784 3256 2908
rect 4924 2784 5168 2990
rect 5686 2940 5732 2974
rect 7124 2948 7130 3034
rect 7156 3032 7666 3058
rect 7748 3050 7800 3064
rect 7778 3044 7800 3050
rect 7684 3032 7800 3044
rect 7156 3030 7800 3032
rect 7156 3010 7666 3030
rect 7684 3010 7800 3030
rect 7156 3006 7800 3010
rect 7152 2976 7208 3006
rect 7340 2989 7391 3006
rect 7400 2990 7800 3006
rect 7412 2989 7800 2990
rect 7340 2988 7800 2989
rect 7340 2970 7400 2988
rect 7440 2980 7800 2988
rect 7440 2976 7666 2980
rect 7684 2976 7800 2980
rect 7440 2970 7800 2976
rect 7452 2962 7636 2970
rect 7468 2954 7636 2962
rect 7456 2952 7636 2954
rect 7174 2944 7206 2952
rect 7280 2944 7398 2946
rect 7452 2926 7636 2952
rect 7664 2946 7800 2970
rect 7680 2942 7800 2946
rect 7684 2930 7800 2942
rect 7146 2916 7178 2924
rect 7308 2916 7370 2918
rect 7276 2900 7308 2916
rect 7390 2914 7452 2926
rect 7310 2900 7342 2910
rect 7276 2868 7342 2900
rect 7366 2902 7374 2910
rect 7366 2868 7376 2902
rect 7390 2889 7410 2914
rect 7400 2872 7410 2889
rect 7422 2872 7440 2914
rect 7444 2911 7452 2914
rect 7456 2886 7474 2926
rect 7506 2925 7636 2926
rect 7518 2888 7558 2904
rect 7568 2888 7636 2925
rect 7664 2906 7800 2930
rect 7664 2900 7680 2906
rect 7684 2900 7800 2906
rect 7506 2886 7568 2888
rect 7468 2878 7574 2886
rect 7452 2872 7574 2878
rect 7390 2868 7574 2872
rect 7276 2858 7574 2868
rect 7276 2852 7314 2858
rect 7276 2850 7308 2852
rect 7280 2830 7286 2850
rect 7340 2846 7574 2858
rect 7328 2818 7574 2846
rect 7390 2817 7574 2818
rect 7588 2817 7614 2888
rect 7664 2848 7800 2900
rect 7684 2832 7800 2848
rect 7390 2816 7614 2817
rect 2860 2770 2926 2776
rect 7340 2766 7494 2816
rect 7680 2800 7800 2832
rect 7390 2748 7444 2752
rect 7468 2748 7574 2766
rect 7340 2726 7574 2748
rect 7328 2724 7574 2726
rect 1464 2708 1516 2722
rect 1496 2704 1516 2708
rect 6664 2708 6716 2722
rect 6664 2704 6684 2708
rect 7328 2698 7614 2724
rect 7390 2696 7614 2698
rect 7340 2694 7531 2696
rect 7532 2694 7614 2696
rect 7280 2664 7286 2684
rect 7340 2664 7614 2694
rect 7684 2686 7800 2800
rect 7664 2670 7800 2686
rect 7844 2676 7906 2806
rect 7919 2795 7995 2806
rect 7930 2778 7984 2795
rect 7938 2756 7984 2778
rect 7960 2730 8066 2756
rect 8010 2694 8066 2730
rect 196 2646 242 2656
rect 184 2642 242 2646
rect 328 2642 336 2656
rect 434 2642 478 2660
rect 184 2614 284 2642
rect 328 2630 478 2642
rect 7244 2630 7264 2664
rect 7276 2662 7308 2664
rect 7276 2656 7314 2662
rect 7340 2656 7588 2664
rect 7276 2636 7588 2656
rect 7702 2642 7746 2670
rect 7802 2642 7852 2656
rect 7938 2646 7984 2656
rect 7938 2642 7996 2646
rect 7702 2636 7852 2642
rect 7276 2630 7452 2636
rect 7506 2630 7588 2636
rect 7696 2630 7852 2636
rect 328 2614 428 2630
rect 7276 2614 7342 2630
rect 116 2604 478 2614
rect 7276 2598 7308 2614
rect 7310 2604 7342 2614
rect 7366 2612 7376 2630
rect 7366 2604 7374 2612
rect 7390 2610 7410 2630
rect 7422 2610 7440 2630
rect 7456 2618 7474 2628
rect 7506 2626 7614 2630
rect 7568 2618 7636 2626
rect 7702 2622 7852 2630
rect 7696 2620 7852 2622
rect 7390 2603 7444 2610
rect 7452 2603 7636 2618
rect 7702 2614 7852 2620
rect 7896 2614 7996 2642
rect 1156 2570 1194 2598
rect 6986 2570 7024 2598
rect 7390 2590 7636 2603
rect 7684 2604 8064 2614
rect 7684 2602 7740 2604
rect 7648 2596 7754 2602
rect 7648 2590 7740 2596
rect 7390 2588 7784 2590
rect 7410 2580 7444 2588
rect 7452 2564 7614 2588
rect 7634 2586 7784 2588
rect 7634 2584 7740 2586
rect 7648 2568 7740 2584
rect 7452 2563 7568 2564
rect 7452 2562 7517 2563
rect 7588 2562 7614 2564
rect 7674 2562 7740 2568
rect 7456 2560 7528 2562
rect 7468 2544 7528 2560
rect 7340 2538 7400 2544
rect 7440 2542 7528 2544
rect 7588 2556 7660 2562
rect 7674 2558 7756 2562
rect 7440 2538 7564 2542
rect 7340 2530 7564 2538
rect 7588 2530 7614 2556
rect 7674 2544 7740 2558
rect 7684 2542 7740 2544
rect 7340 2526 8130 2530
rect 7340 2522 7440 2526
rect 7328 2516 7444 2522
rect 7328 2494 7420 2516
rect 7440 2494 7444 2516
rect 7362 2492 7386 2494
rect 7390 2492 7440 2494
rect 7452 2492 8130 2526
rect 7340 2490 7420 2492
rect 3516 2484 3528 2490
rect 4674 2484 4686 2490
rect 3488 2478 3534 2484
rect 4646 2478 4692 2484
rect 3482 2472 3540 2478
rect 3482 2466 3500 2472
rect 3494 2456 3500 2466
rect 3482 2448 3500 2456
rect 3522 2466 3540 2472
rect 4640 2472 4698 2478
rect 7340 2476 7440 2490
rect 7468 2476 8130 2492
rect 4640 2466 4658 2472
rect 3522 2456 3534 2466
rect 4652 2456 4658 2466
rect 3522 2448 3540 2456
rect 3482 2444 3540 2448
rect 4640 2448 4658 2456
rect 4680 2466 4698 2472
rect 7318 2468 7440 2476
rect 7318 2466 7444 2468
rect 4680 2456 4692 2466
rect 7340 2464 7440 2466
rect 4680 2448 4698 2456
rect 7340 2450 7390 2464
rect 7400 2458 7440 2464
rect 7400 2450 7440 2456
rect 7328 2448 7444 2450
rect 4640 2444 4698 2448
rect 3494 2442 3528 2444
rect 4652 2442 4686 2444
rect 3516 2432 3528 2442
rect 4674 2432 4686 2442
rect 7318 2438 7444 2448
rect 7328 2424 7444 2438
rect 7328 2422 7420 2424
rect 7440 2422 7444 2424
rect 7366 2420 7386 2422
rect 7400 2420 7440 2422
rect 7452 2420 7486 2464
rect 7518 2458 7558 2476
rect 7518 2422 7558 2456
rect 7340 2388 7390 2420
rect 7400 2390 7420 2420
rect 7506 2394 7568 2422
rect 7452 2388 7568 2394
rect 7340 2372 7400 2388
rect 7440 2380 7556 2388
rect 7440 2372 7588 2380
rect 7340 2370 7588 2372
rect 7362 2352 7440 2370
rect 7452 2362 7588 2370
rect 7456 2352 7494 2354
rect 7496 2352 7588 2362
rect 7390 2326 7418 2344
rect 7452 2340 7486 2352
rect 7506 2350 7588 2352
rect 7452 2326 7506 2340
rect 3496 2306 3502 2308
rect 3524 2306 3530 2308
rect 3496 2302 3530 2306
rect 3538 2302 3562 2324
rect 3496 2300 3562 2302
rect 4652 2306 4658 2316
rect 4680 2310 4686 2316
rect 4680 2306 4692 2310
rect 4652 2300 4692 2306
rect 3496 2290 3508 2300
rect 3518 2294 3562 2300
rect 3518 2288 3530 2294
rect 3534 2290 3562 2294
rect 4674 2294 4692 2300
rect 7276 2300 7308 2316
rect 7362 2310 7370 2318
rect 7390 2314 7452 2326
rect 7310 2300 7342 2310
rect 4674 2288 4686 2294
rect 7276 2268 7342 2300
rect 7362 2302 7374 2310
rect 7362 2272 7376 2302
rect 7390 2300 7418 2314
rect 7390 2289 7410 2300
rect 7400 2272 7410 2289
rect 7422 2272 7440 2314
rect 7444 2311 7452 2314
rect 7456 2286 7474 2326
rect 7506 2325 7568 2326
rect 7554 2304 7568 2325
rect 7518 2288 7568 2304
rect 7506 2278 7568 2288
rect 7452 2272 7568 2278
rect 7366 2268 7376 2272
rect 7390 2268 7568 2272
rect 7276 2258 7568 2268
rect 7276 2252 7314 2258
rect 7340 2256 7568 2258
rect 7276 2250 7308 2252
rect 7280 2230 7286 2250
rect 7340 2246 7556 2256
rect 7328 2238 7556 2246
rect 7328 2236 7530 2238
rect 7328 2218 7531 2236
rect 7390 2216 7506 2218
rect 7340 2166 7494 2216
rect 7390 2148 7444 2152
rect 7340 2126 7494 2148
rect 1794 1932 1810 2064
rect 6306 2032 6324 2060
rect 6334 2038 6336 2104
rect 7328 2098 7536 2126
rect 7336 2096 7506 2098
rect 7280 2064 7286 2084
rect 7340 2072 7494 2096
rect 7506 2078 7531 2096
rect 7506 2076 7530 2078
rect 7506 2074 7556 2076
rect 7506 2072 7564 2074
rect 7276 2062 7308 2064
rect 7276 2056 7314 2062
rect 7340 2058 7564 2072
rect 7340 2056 7390 2058
rect 7276 2046 7390 2056
rect 7276 2014 7342 2046
rect 7276 1998 7308 2014
rect 7310 2004 7342 2014
rect 7366 2012 7376 2046
rect 7400 2025 7410 2056
rect 7366 2004 7374 2012
rect 7390 2010 7410 2025
rect 7422 2010 7440 2056
rect 7452 2036 7568 2058
rect 7456 2018 7474 2028
rect 7506 2026 7568 2036
rect 7390 2003 7444 2010
rect 7452 2003 7568 2018
rect 7390 1988 7568 2003
rect 7410 1980 7444 1988
rect 7452 1964 7506 1988
rect 1794 1896 1962 1932
rect 7156 1924 7412 1964
rect 7452 1963 7568 1964
rect 7452 1962 7517 1963
rect 7456 1960 7494 1962
rect 7440 1940 7494 1944
rect 7496 1942 7528 1962
rect 7496 1940 7564 1942
rect 7440 1926 7564 1940
rect 7156 1902 7420 1924
rect 7440 1902 7444 1922
rect 7452 1902 7486 1926
rect 6362 1872 6472 1894
rect 7156 1892 7486 1902
rect 7506 1892 7568 1926
rect 6334 1844 6500 1866
rect 7156 1856 7480 1892
rect 7156 1838 7412 1856
rect 7440 1842 7506 1856
rect 7020 1834 7048 1836
rect 7154 1834 7412 1838
rect 6194 1796 6232 1824
rect 6282 1796 6338 1824
rect 7154 1796 7208 1834
rect 7622 1796 7666 2088
rect 6202 1768 6266 1792
rect 7788 1754 7806 1770
rect 7816 1754 7850 1788
rect 7788 1720 7800 1754
rect 7822 1720 7838 1736
rect 7822 1702 7834 1720
rect 6386 1652 6476 1678
rect 6118 1556 6490 1652
rect 6118 1510 6554 1556
rect 6118 1498 6490 1510
rect 6322 1478 6346 1498
rect 6356 1478 6412 1498
rect 6356 1464 6380 1478
rect 6390 1472 6412 1478
rect 6330 1450 6346 1464
rect 6302 1426 6320 1448
rect 6356 1444 6364 1464
rect 6418 1444 6440 1498
rect 6418 1394 6460 1416
rect 6434 1374 6480 1388
rect 6410 1366 6480 1374
rect 6410 1358 6460 1366
rect 6434 1342 6440 1358
rect 6434 1330 6480 1342
rect 6844 610 7216 852
<< nwell >>
rect 1794 3004 2190 3006
rect 6386 3004 6680 3006
rect 7156 2970 7412 3006
rect 1794 2870 1808 2906
rect 1794 1896 1810 1932
rect 7156 1796 7412 1834
<< locali >>
rect 3492 2478 3532 2492
rect 3492 2444 3494 2478
rect 3528 2444 3532 2478
rect 3492 2334 3532 2444
rect 3492 2300 3496 2334
rect 3530 2300 3532 2334
rect 3492 2290 3532 2300
rect 4642 2478 4700 2492
rect 4642 2444 4652 2478
rect 4686 2444 4700 2478
rect 4642 2334 4700 2444
rect 4642 2300 4652 2334
rect 4686 2300 4700 2334
rect 4642 2290 4700 2300
<< viali >>
rect 3494 2444 3528 2478
rect 3496 2300 3530 2334
rect 4652 2444 4686 2478
rect 4652 2300 4686 2334
<< metal1 >>
rect 1842 2996 1898 3006
rect 1842 2994 1906 2996
rect 1948 2994 1986 3006
rect 1842 2942 1848 2994
rect 1900 2942 1906 2994
rect 3244 2988 3290 3004
rect 3488 2988 3534 3004
rect 3946 2974 4234 3006
rect 4646 2988 4692 3006
rect 4890 2990 4936 3006
rect 6194 2990 6232 3006
rect 6282 2996 6338 3006
rect 6282 2992 6346 2996
rect 1842 2940 1906 2942
rect 6282 2940 6288 2992
rect 6340 2940 6346 2992
rect 7020 2978 7088 3006
rect 7152 2976 7208 3006
rect 6282 2936 6346 2940
rect 3494 2442 3528 2444
rect 4652 2442 4686 2444
rect 3490 2380 3554 2384
rect 3490 2302 3496 2380
rect 3548 2328 3554 2380
rect 3530 2324 3554 2328
rect 4630 2368 4694 2374
rect 3530 2302 3538 2324
rect 4630 2316 4636 2368
rect 4688 2316 4694 2368
rect 4630 2310 4652 2316
rect 3534 2290 3538 2302
rect 4686 2310 4694 2316
rect 6718 1890 6784 1894
rect 4630 1864 4694 1868
rect 4630 1812 4636 1864
rect 4688 1812 4694 1864
rect 6718 1838 6724 1890
rect 6778 1838 6784 1890
rect 6718 1836 6784 1838
rect 4630 1808 4694 1812
rect 6716 1830 6800 1836
rect 6920 1834 7020 1836
rect 6920 1830 7088 1834
rect 6716 1808 7088 1830
rect 6194 1796 6232 1806
rect 6282 1796 6338 1806
rect 6772 1802 6952 1808
rect 7020 1796 7088 1808
rect 7154 1796 7208 1838
<< via1 >>
rect 1848 2942 1900 2994
rect 6288 2940 6340 2992
rect 3496 2334 3548 2380
rect 3496 2328 3530 2334
rect 3530 2328 3548 2334
rect 4636 2334 4688 2368
rect 4636 2316 4652 2334
rect 4652 2316 4686 2334
rect 4686 2316 4688 2334
rect 4636 1812 4688 1864
rect 6724 1838 6778 1890
<< metal2 >>
rect 1842 2994 1906 2996
rect 1842 2942 1848 2994
rect 1900 2972 1906 2994
rect 6282 2992 6346 2996
rect 6282 2972 6288 2992
rect 1900 2942 6288 2972
rect 1842 2940 6288 2942
rect 6340 2940 6346 2992
rect 6506 2952 6568 3000
rect 1842 2936 6346 2940
rect 1794 2870 1808 2906
rect 6728 2826 6772 2830
rect 3574 2750 3742 2790
rect 6718 2758 6772 2826
rect 3664 2656 5692 2700
rect 6370 2658 6440 2702
rect 3654 2462 5456 2506
rect 3490 2380 3554 2384
rect 3490 2328 3496 2380
rect 3548 2374 3554 2380
rect 3548 2368 4694 2374
rect 3548 2328 4636 2368
rect 3490 2324 4636 2328
rect 4630 2316 4636 2324
rect 4688 2316 4694 2368
rect 4630 2310 4694 2316
rect 3664 2106 4796 2150
rect 3564 2046 3660 2048
rect 3564 1998 3742 2046
rect 4752 2040 4796 2106
rect 5412 2140 5456 2462
rect 5648 2416 5692 2656
rect 6732 2644 6772 2646
rect 6732 2578 6776 2644
rect 6736 2576 6776 2578
rect 6522 2418 6586 2466
rect 7390 2464 7412 2510
rect 5642 2408 5692 2416
rect 5642 2280 5694 2408
rect 7390 2300 7412 2344
rect 5642 2238 6468 2280
rect 6426 2210 6468 2238
rect 6426 2168 6830 2210
rect 5412 2096 5982 2140
rect 5626 2040 6830 2050
rect 4752 2008 6830 2040
rect 4752 1996 5704 2008
rect 1794 1896 1810 1932
rect 6718 1890 6784 1894
rect 4630 1866 4694 1868
rect 6718 1866 6724 1890
rect 4630 1864 6724 1866
rect 4630 1812 4636 1864
rect 4688 1838 6724 1864
rect 6778 1838 6784 1890
rect 4688 1834 6784 1838
rect 4688 1832 4768 1834
rect 4688 1812 4694 1832
rect 4630 1808 4694 1812
use sky130_hilas_FGBias2x1cell  sky130_hilas_FGBias2x1cell_0
timestamp 1632256332
transform 1 0 4872 0 1 2560
box 0 0 3308 2104
use sky130_hilas_FGBiasWeakGate2x1cell  sky130_hilas_FGBiasWeakGate2x1cell_0
timestamp 1632256335
transform -1 0 3308 0 1 2560
box 0 0 3308 2104
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1632256331
transform 1 0 7102 0 1 1878
box 0 0 716 1504
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1632255311
transform 1 0 6118 0 -1 2126
box 0 0 1098 2126
<< labels >>
rlabel metal2 3574 2750 3646 2788 0 VIN11
port 2 nsew analog default
rlabel metal2 3564 1998 3636 2048 0 VIN12
port 1 nsew analog default
rlabel metal1 7020 2994 7088 3006 0 VGND
port 7 nsew analog default
rlabel metal1 7152 2994 7208 3006 0 VPWR
port 6 nsew analog default
rlabel metal1 7154 1796 7208 1808 0 VPWR
port 6 nsew power default
rlabel metal1 7020 1796 7088 1808 0 VGND
port 7 nsew ground default
rlabel metal2 6522 2418 6586 2466 0 VIN21
port 3 nsew analog default
rlabel metal2 6506 2952 6568 3000 1 VIN22
port 4 n analog default
rlabel metal1 6282 2990 6338 3006 0 VINJ
port 8 nsew power default
rlabel metal1 6282 1796 6338 1806 0 VINJ
port 8 nsew power default
rlabel metal2 7390 2464 7412 2510 0 OUTPUT1
port 9 nsew analog default
rlabel metal2 7390 2300 7412 2344 0 OUTPUT2
port 10 nsew analog default
rlabel metal2 1794 2870 1808 2906 0 DRAIN1
port 11 nsew
rlabel metal2 1794 1896 1810 1932 0 DRAIN2
port 12 nsew
rlabel metal1 1842 2992 1898 3006 0 VINJ
port 8 nsew
rlabel metal1 1948 2994 1986 3006 0 COLSEL2
port 13 nsew
rlabel metal1 3244 2988 3290 3004 0 GATE2
port 14 nsew
rlabel metal1 3488 2988 3534 3004 0 VGND
port 7 nsew
rlabel metal1 4890 2990 4936 3006 0 GATE1
port 15 nsew
rlabel metal1 4646 2990 4692 3006 0 VGND
port 7 nsew
rlabel metal1 6194 2990 6232 3006 0 COLSEL1
port 16 nsew
rlabel metal1 6194 1796 6232 1806 0 COLSEL1
port 16 nsew
rlabel metal1 4030 2982 4150 3006 0 VTUN
port 17 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
