* NGSPICE file created from /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_capacitorSize01.ext - technology: sky130A

.subckt sky130_hilas_CapModule02 c1_n808_n410# $SUB m3_n886_n490#
X0 c1_n808_n410# m3_n886_n490# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=6.38e+06u
.ends

.subckt home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_capacitorSize01
+ CapTerm02 CapTerm01
Xsky130_hilas_CapModule02_0 CapTerm01 $SUB CapTerm02 sky130_hilas_CapModule02
.ends

