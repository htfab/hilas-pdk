VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_capacitorSize01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_capacitorSize01 ;
  ORIGIN -14.140 0.480 ;
  SIZE 10.420 BY 5.830 ;
  PIN CapTerm02
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 24.200 2.330 24.560 2.610 ;
    END
  END CapTerm02
  PIN CapTerm01
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 14.160 2.320 14.430 2.600 ;
    END
  END CapTerm01
  OBS
      LAYER met2 ;
        RECT 14.140 2.890 24.560 4.980 ;
        RECT 14.140 2.880 23.920 2.890 ;
        RECT 14.710 2.050 23.920 2.880 ;
        RECT 14.710 2.040 24.560 2.050 ;
        RECT 14.140 -0.050 24.560 2.040 ;
      LAYER met3 ;
        RECT 14.160 -0.480 24.440 5.350 ;
      LAYER met4 ;
        RECT 14.250 0.620 24.400 2.790 ;
  END
END sky130_hilas_capacitorSize01
END LIBRARY

