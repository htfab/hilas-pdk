magic
tech sky130A
timestamp 1628704418
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_3
timestamp 1628285143
transform 1 0 73 0 1 22
box 147 -22 266 265
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_4
timestamp 1628285143
transform 1 0 -147 0 1 22
box 147 -22 266 265
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_0
timestamp 1628285143
transform 1 0 -92 0 1 22
box 147 -22 266 265
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_1
timestamp 1628285143
transform 1 0 -37 0 1 22
box 147 -22 266 265
use sky130_hilas_pFETmed  sky130_hilas_pFETmed_2
timestamp 1628285143
transform 1 0 18 0 1 22
box 147 -22 266 265
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
