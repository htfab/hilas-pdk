magic
tech sky130A
timestamp 1632256320
<< error_s >>
rect 63 578 102 581
rect 63 536 102 539
rect 61 482 100 485
rect 61 440 100 443
rect 61 386 100 389
rect 61 344 100 347
rect 40 324 121 336
rect 61 302 100 305
rect 61 260 100 263
rect 134 245 150 255
rect 155 219 171 245
rect 0 96 161 212
rect 164 203 185 204
rect 63 62 102 65
rect 63 20 102 23
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_0
timestamp 1632251308
transform 1 0 1 0 1 480
box 0 0 172 121
use sky130_hilas_pFETdevice01b  sky130_hilas_pFETdevice01b_1
timestamp 1632255311
transform 1 0 0 0 1 192
box 0 0 188 133
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_6
timestamp 1632251433
transform 1 0 0 0 1 384
box 0 0 161 121
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_3
timestamp 1632251433
transform 1 0 0 0 1 288
box 0 0 161 121
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_0
timestamp 1632251433
transform 1 0 0 0 1 96
box 0 0 161 121
use sky130_hilas_pFETdevice01a  sky130_hilas_pFETdevice01a_0
timestamp 1632251417
transform 1 0 1 0 1 0
box 0 0 161 85
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
