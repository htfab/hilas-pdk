magic
tech sky130A
timestamp 1628616643
<< error_p >>
rect 62 98 101 101
rect 62 56 101 59
<< nwell >>
rect 0 0 161 121
<< pmos >>
rect 62 59 101 98
<< pdiff >>
rect 34 59 62 98
rect 101 59 127 98
<< poly >>
rect 0 96 26 111
rect 62 98 101 111
rect 11 51 26 96
rect 62 51 101 59
rect 11 36 151 51
rect 136 15 151 36
rect 136 0 172 15
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
