VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_horiztranscell01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_horiztranscell01 ;
  ORIGIN 4.760 -0.480 ;
  SIZE 4.430 BY 3.110 ;
  OBS
      LAYER nwell ;
        RECT -3.640 0.480 -0.330 3.590 ;
      LAYER li1 ;
        RECT -4.600 3.040 -4.260 3.210 ;
        RECT -3.240 3.040 -2.910 3.210 ;
        RECT -4.610 2.250 -4.260 2.420 ;
        RECT -3.240 2.250 -2.910 2.420 ;
        RECT -4.610 1.460 -4.260 1.630 ;
        RECT -3.240 1.460 -2.910 1.630 ;
        RECT -2.490 1.440 -2.320 3.130 ;
        RECT -1.660 3.040 -1.480 3.230 ;
        RECT -1.660 1.430 -1.490 3.040 ;
        RECT -1.300 2.230 -1.060 2.560 ;
        RECT -1.290 1.940 -1.090 2.230 ;
        RECT -1.290 1.930 -1.100 1.940 ;
        RECT -0.930 1.760 -0.720 1.770 ;
        RECT -0.940 1.180 -0.720 1.760 ;
        RECT -0.930 1.150 -0.720 1.180 ;
        RECT -2.740 0.880 -2.210 1.050 ;
        RECT -0.930 0.800 -0.730 1.150 ;
      LAYER mcon ;
        RECT -1.280 2.000 -1.100 2.190 ;
        RECT -0.920 1.180 -0.750 1.350 ;
      LAYER met1 ;
        RECT -1.690 2.910 -1.450 3.290 ;
        RECT -1.260 2.480 -1.100 3.500 ;
        RECT -1.300 2.240 -1.070 2.480 ;
        RECT -1.300 2.230 -1.060 2.240 ;
        RECT -1.310 1.960 -1.060 2.230 ;
        RECT -1.290 1.930 -1.070 1.960 ;
        RECT -2.810 0.770 -2.510 1.150 ;
        RECT -1.290 0.480 -1.100 1.930 ;
        RECT -0.850 1.810 -0.690 3.500 ;
        RECT -0.850 1.720 -0.680 1.810 ;
        RECT -0.960 1.670 -0.680 1.720 ;
        RECT -0.960 1.120 -0.690 1.670 ;
        RECT -0.850 0.480 -0.690 1.120 ;
      LAYER via ;
        RECT -2.790 0.820 -2.530 1.090 ;
      LAYER met2 ;
        RECT -2.890 0.970 -0.330 1.150 ;
        RECT -2.810 0.770 -2.510 0.970 ;
  END
END sky130_hilas_horiztranscell01
END LIBRARY

