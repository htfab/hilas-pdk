magic
tech sky130A
timestamp 1627400803
<< error_s >>
rect 783 388 784 389
<< nwell >>
rect 0 604 191 605
rect 0 44 560 604
rect 760 587 888 605
rect 0 26 43 44
rect 0 3 71 26
rect 0 1 43 3
rect 760 0 888 19
<< nsubdiff >>
rect 19 521 50 558
rect 19 504 25 521
rect 42 504 50 521
rect 19 487 50 504
rect 19 470 25 487
rect 42 470 50 487
rect 19 453 50 470
rect 19 436 25 453
rect 42 436 50 453
rect 19 419 50 436
rect 19 402 25 419
rect 42 402 50 419
rect 19 385 50 402
rect 19 368 25 385
rect 42 368 50 385
rect 19 353 50 368
rect 18 218 50 251
rect 18 201 26 218
rect 43 201 50 218
rect 18 184 50 201
rect 18 167 26 184
rect 43 167 50 184
rect 18 150 50 167
rect 18 133 26 150
rect 43 133 50 150
rect 18 116 50 133
rect 18 99 26 116
rect 43 99 50 116
rect 18 82 50 99
rect 18 65 26 82
rect 43 65 50 82
rect 18 50 50 65
<< nsubdiffcont >>
rect 25 504 42 521
rect 25 470 42 487
rect 25 436 42 453
rect 25 402 42 419
rect 25 368 42 385
rect 26 201 43 218
rect 26 167 43 184
rect 26 133 43 150
rect 26 99 43 116
rect 26 65 43 82
<< locali >>
rect 67 557 101 558
rect 42 533 101 557
rect 42 484 84 533
rect 765 458 767 475
rect 784 458 790 475
rect 765 421 790 458
rect 765 405 786 421
rect 765 388 767 405
rect 784 388 786 405
rect 765 386 786 388
rect 25 351 42 368
rect 26 57 43 65
<< viali >>
rect 25 521 42 538
rect 25 487 42 504
rect 84 516 101 533
rect 84 482 101 499
rect 25 453 42 470
rect 25 419 42 436
rect 25 385 42 402
rect 767 458 784 475
rect 767 388 784 405
rect 26 218 43 235
rect 26 184 43 201
rect 26 150 43 167
rect 26 116 43 133
rect 26 82 43 99
<< metal1 >>
rect 692 591 726 605
rect 759 590 786 605
rect 22 558 75 559
rect 22 557 101 558
rect 22 551 104 557
rect 22 538 34 551
rect 22 521 25 538
rect 93 533 104 551
rect 22 504 34 521
rect 101 527 104 533
rect 101 516 107 527
rect 22 487 25 504
rect 93 499 107 516
rect 22 479 34 487
rect 101 498 107 499
rect 101 482 104 498
rect 93 479 104 482
rect 22 473 104 479
rect 762 475 794 479
rect 22 470 86 473
rect 22 453 25 470
rect 42 453 86 470
rect 22 436 86 453
rect 22 419 25 436
rect 42 419 86 436
rect 22 402 86 419
rect 22 385 25 402
rect 42 385 86 402
rect 762 389 763 475
rect 789 389 794 475
rect 762 388 767 389
rect 784 388 794 389
rect 762 387 794 388
rect 765 386 794 387
rect 22 235 86 385
rect 22 218 26 235
rect 43 218 86 235
rect 22 201 86 218
rect 22 184 26 201
rect 43 184 86 201
rect 22 167 86 184
rect 22 150 26 167
rect 43 150 86 167
rect 22 133 86 150
rect 22 116 26 133
rect 43 116 86 133
rect 22 99 86 116
rect 22 82 26 99
rect 43 82 86 99
rect 22 55 86 82
rect 44 54 86 55
rect 692 0 726 19
rect 759 0 786 21
<< via1 >>
rect 34 538 93 551
rect 34 521 42 538
rect 42 533 93 538
rect 42 521 84 533
rect 34 516 84 521
rect 84 516 93 533
rect 34 504 93 516
rect 34 487 42 504
rect 42 499 93 504
rect 42 487 84 499
rect 34 482 84 487
rect 84 482 93 499
rect 34 479 93 482
rect 763 458 767 475
rect 767 458 784 475
rect 784 458 789 475
rect 763 405 789 458
rect 763 389 767 405
rect 767 389 784 405
rect 784 389 789 405
<< metal2 >>
rect 79 558 103 605
rect 439 578 464 604
rect 27 551 103 558
rect 27 479 34 551
rect 93 523 103 551
rect 93 500 481 523
rect 93 479 103 500
rect 27 476 103 479
rect 27 475 72 476
rect 458 464 481 500
rect 545 480 570 517
rect 760 475 793 479
rect 760 464 763 475
rect 188 431 407 453
rect 458 444 763 464
rect 484 443 763 444
rect 548 395 569 424
rect 760 389 763 443
rect 789 389 793 475
rect 760 386 793 389
rect 873 334 888 356
rect 443 311 468 334
rect 1 270 147 294
rect 287 270 315 294
rect 1 269 65 270
rect 873 252 888 274
rect 392 187 569 207
rect 235 152 251 170
rect 233 151 251 152
rect 211 138 251 151
rect 211 89 247 138
rect 363 106 569 127
rect 5 3 170 26
rect 283 2 309 27
<< rmetal2 >>
rect 72 475 103 476
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_0
timestamp 1608384750
transform 1 0 85 0 1 440
box 133 -440 320 165
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1608384750
transform 1 0 241 0 -1 165
box 133 -440 320 165
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_2
timestamp 1608384750
transform 1 0 -90 0 1 440
box 133 -440 320 165
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1607089160
transform 1 0 173 0 1 441
box -14 -15 20 18
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1608069483
transform 1 0 733 0 1 41
box -172 -22 155 550
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1607089160
transform 1 0 89 0 1 569
box -14 -15 20 18
<< labels >>
rlabel metal1 692 0 726 6 0 VGND
port 3 nsew ground default
rlabel metal1 759 0 786 6 0 VPWR
port 4 nsew power default
rlabel metal1 692 600 726 605 0 VGND
port 3 nsew ground default
rlabel metal1 759 600 786 605 0 VPWR
port 4 nsew power default
rlabel metal2 287 270 310 294 0 VIN11
port 7 nsew analog default
rlabel metal2 443 311 468 334 0 VIN21
port 6 nsew analog default
rlabel metal2 283 2 306 27 0 VIN12
port 8 nsew analog default
rlabel metal2 439 578 464 604 0 VIN22
port 5 nsew analog default
rlabel metal2 873 252 888 274 0 VOUT_AMP1
port 2 nsew analog default
rlabel metal2 873 334 888 356 0 VOUT_AMP2
port 1 nsew analog default
rlabel metal2 79 597 103 605 0 VPWR
port 4 nsew power default
rlabel metal2 43 270 50 294 0 VBIAS1
port 10 nsew analog default
rlabel metal2 43 3 50 26 0 VBIAS2
port 9 nsew analog default
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
