magic
tech sky130A
timestamp 1607186163
<< error_s >>
rect 85 -19 102 -18
rect 109 -30 110 11
rect 73 -42 77 -30
rect 109 -42 114 -30
rect 109 -58 110 -42
rect 109 -90 110 -59
rect 109 -148 110 -119
<< nwell >>
rect -61 112 158 285
<< nmos >>
rect -8 11 25 40
rect 77 11 110 40
rect -8 -119 25 -90
rect 77 -119 110 -90
<< pmos >>
rect -40 164 28 194
rect 64 164 132 194
<< ndiff >>
rect -8 64 25 68
rect -8 47 0 64
rect 17 47 25 64
rect -8 40 25 47
rect 77 64 110 68
rect 77 47 85 64
rect 102 47 110 64
rect 77 40 110 47
rect -8 4 25 11
rect -8 -13 0 4
rect 17 -13 25 4
rect -8 -19 25 -13
rect -8 -67 25 -60
rect -8 -84 0 -67
rect 17 -84 25 -67
rect -8 -90 25 -84
rect 77 4 110 11
rect 77 -13 85 4
rect 102 -13 110 4
rect 77 -19 110 -13
rect 77 -66 110 -59
rect 77 -83 85 -66
rect 102 -83 110 -66
rect 77 -90 110 -83
rect -8 -126 25 -119
rect -8 -143 -1 -126
rect 17 -143 25 -126
rect -8 -147 25 -143
rect 77 -125 110 -119
rect 77 -142 84 -125
rect 103 -142 110 -125
rect 77 -148 110 -142
<< pdiff >>
rect -40 218 28 224
rect -40 201 -32 218
rect -14 201 4 218
rect 22 201 28 218
rect -40 194 28 201
rect 64 218 132 224
rect 64 201 72 218
rect 90 201 109 218
rect 128 201 132 218
rect 64 194 132 201
rect -40 157 28 164
rect -40 140 -32 157
rect -14 140 4 157
rect 22 140 28 157
rect -40 131 28 140
rect 64 157 132 164
rect 64 140 70 157
rect 88 140 106 157
rect 124 140 132 157
rect 64 136 132 140
rect 71 131 132 136
<< ndiffc >>
rect 0 47 17 64
rect 85 47 102 64
rect 0 -13 17 4
rect 0 -84 17 -67
rect 85 -13 102 4
rect 85 -83 102 -66
rect -1 -143 17 -126
rect 84 -142 103 -125
<< pdiffc >>
rect -32 201 -14 218
rect 4 201 22 218
rect 72 201 90 218
rect 109 201 128 218
rect -32 140 -14 157
rect 4 140 22 157
rect 70 140 88 157
rect 106 140 124 157
<< psubdiff >>
rect -8 -31 25 -19
rect -8 -48 0 -31
rect 17 -48 25 -31
rect -8 -60 25 -48
rect 77 -30 110 -19
rect 77 -47 85 -30
rect 102 -47 110 -30
rect 77 -58 110 -47
rect 77 -59 109 -58
<< nsubdiff >>
rect -40 253 28 265
rect -40 236 -32 253
rect -14 236 4 253
rect 22 236 28 253
rect -40 224 28 236
rect 64 253 132 265
rect 64 236 72 253
rect 90 236 109 253
rect 128 236 132 253
rect 64 224 132 236
<< psubdiffcont >>
rect 0 -48 17 -31
rect 85 -47 102 -30
<< nsubdiffcont >>
rect -32 236 -14 253
rect 4 236 22 253
rect 72 236 90 253
rect 109 236 128 253
<< poly >>
rect -53 164 -40 194
rect 28 164 64 194
rect 132 164 145 194
rect 36 120 53 164
rect 30 112 57 120
rect 30 95 35 112
rect 52 95 57 112
rect 30 87 57 95
rect -278 23 -251 27
rect -33 11 -8 40
rect 25 11 38 40
rect 63 11 77 40
rect 110 11 133 40
rect -33 -90 -17 11
rect 117 -90 133 11
rect -33 -119 -8 -90
rect 25 -119 38 -90
rect 62 -119 77 -90
rect 110 -119 133 -90
rect -278 -123 -251 -120
rect -33 -158 -17 -119
rect -33 -166 26 -158
rect 117 -159 133 -119
rect -33 -183 -1 -166
rect 17 -183 26 -166
rect -33 -189 26 -183
rect 77 -167 133 -159
rect 77 -184 86 -167
rect 103 -184 133 -167
rect 77 -189 133 -184
<< polycont >>
rect 35 95 52 112
rect -1 -183 17 -166
rect 86 -184 103 -167
<< locali >>
rect -40 236 -32 253
rect -14 236 4 253
rect 22 236 72 253
rect 90 236 109 253
rect 128 236 136 253
rect -40 218 136 236
rect -40 201 -32 218
rect -14 201 4 218
rect 22 201 72 218
rect 90 201 109 218
rect 128 201 136 218
rect -40 140 -32 157
rect -14 140 4 157
rect 22 140 31 157
rect 62 140 70 157
rect 88 140 106 157
rect 124 140 132 157
rect -5 123 31 140
rect -5 112 60 123
rect -5 95 35 112
rect 52 95 60 112
rect -5 87 60 95
rect -5 64 22 87
rect 85 65 110 140
rect 77 64 110 65
rect -8 47 0 64
rect 17 47 25 64
rect 77 47 85 64
rect 102 47 110 64
rect -12 -13 0 4
rect 17 -13 29 4
rect -12 -20 29 -13
rect 73 -13 85 4
rect 102 -13 114 4
rect 73 -20 114 -13
rect -12 -30 114 -20
rect -12 -31 85 -30
rect -12 -48 0 -31
rect 17 -47 85 -31
rect 102 -47 114 -30
rect 17 -48 114 -47
rect -12 -58 114 -48
rect -12 -67 29 -58
rect -12 -84 0 -67
rect 17 -84 29 -67
rect 73 -66 114 -58
rect 73 -83 85 -66
rect 102 -83 114 -66
rect -9 -143 -1 -126
rect 17 -143 25 -126
rect 76 -142 84 -125
rect 103 -142 112 -125
rect 76 -143 112 -142
rect -1 -166 17 -143
rect -1 -192 17 -183
rect 84 -167 103 -143
rect 84 -184 86 -167
rect 84 -192 103 -184
use nFET03  nFET03_3
timestamp 1607185713
transform 1 0 -278 0 1 46
box -31 -19 58 42
use nFET03  nFET03_2
timestamp 1607185713
transform 1 0 -278 0 1 -19
box -31 -19 58 42
use nFET03  nFET03_1
timestamp 1607185713
transform 1 0 -278 0 1 -101
box -31 -19 58 42
use nFET03  nFET03_0
timestamp 1607185713
transform 1 0 -278 0 1 -165
box -31 -19 58 42
<< end >>
