magic
tech sky130A
timestamp 1627744303
<< locali >>
rect -13 10 19 14
rect -13 9 20 10
rect -13 -8 -7 9
rect 10 -8 20 9
rect -13 -9 20 -8
rect -13 -12 19 -9
<< viali >>
rect -7 -8 10 9
<< metal1 >>
rect -14 14 18 17
rect -14 -12 -11 14
rect 15 -12 18 14
rect -14 -15 18 -12
<< via1 >>
rect -11 9 15 14
rect -11 -8 -7 9
rect -7 -8 10 9
rect 10 -8 15 9
rect -11 -12 15 -8
<< metal2 >>
rect -14 14 17 18
rect -14 -12 -11 14
rect 15 -12 17 14
rect -14 -15 17 -12
<< end >>
