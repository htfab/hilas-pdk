magic
tech sky130A
timestamp 1628285143
<< error_s >>
rect -147 91 -97 97
rect 173 91 223 97
rect -147 49 -97 55
rect 173 49 223 55
rect -147 25 -97 30
rect -7 24 43 30
rect 173 25 223 30
rect -147 -17 -97 -12
rect -7 -18 43 -12
rect 173 -17 223 -12
<< nwell >>
rect -232 -45 110 124
<< mvnmos >>
rect 173 55 223 91
rect 173 -12 223 25
<< mvpmos >>
rect -147 55 -97 91
rect -147 -12 -97 25
rect -7 -12 43 24
<< mvndiff >>
rect 145 79 173 91
rect 145 62 150 79
rect 167 62 173 79
rect 145 55 173 62
rect 223 79 251 91
rect 223 62 229 79
rect 246 62 251 79
rect 223 55 251 62
rect 145 17 173 25
rect 145 0 150 17
rect 167 0 173 17
rect 145 -12 173 0
rect 223 17 251 25
rect 223 0 229 17
rect 246 0 251 17
rect 223 -12 251 0
<< mvpdiff >>
rect -177 78 -147 91
rect -177 61 -170 78
rect -153 61 -147 78
rect -177 55 -147 61
rect -97 79 -67 91
rect -97 62 -91 79
rect -74 62 -67 79
rect -97 55 -67 62
rect -177 18 -147 25
rect -177 1 -170 18
rect -153 1 -147 18
rect -177 -12 -147 1
rect -97 17 -67 25
rect -97 0 -91 17
rect -73 0 -67 17
rect -97 -12 -67 0
rect -37 17 -7 24
rect -37 0 -30 17
rect -13 0 -7 17
rect -37 -12 -7 0
rect 43 17 73 24
rect 43 0 49 17
rect 66 0 73 17
rect 43 -12 73 0
<< mvndiffc >>
rect 150 62 167 79
rect 229 62 246 79
rect 150 0 167 17
rect 229 0 246 17
<< mvpdiffc >>
rect -170 61 -153 78
rect -91 62 -74 79
rect -170 1 -153 18
rect -91 0 -73 17
rect -30 0 -13 17
rect 49 0 66 17
<< psubdiff >>
rect 283 22 314 34
rect 283 5 287 22
rect 304 5 314 22
rect 283 -7 314 5
<< nsubdiff >>
rect -214 56 -189 86
rect -214 39 -210 56
rect -193 39 -189 56
rect -214 22 -189 39
rect -214 5 -210 22
rect -193 5 -189 22
rect -214 -7 -189 5
<< psubdiffcont >>
rect 287 5 304 22
<< nsubdiffcont >>
rect -210 39 -193 56
rect -210 5 -193 22
<< poly >>
rect -147 99 319 114
rect -147 91 -97 99
rect 173 91 223 99
rect 283 96 319 99
rect -51 67 -11 71
rect -51 65 43 67
rect -147 25 -97 55
rect -51 48 -43 65
rect -26 48 43 65
rect 283 79 294 96
rect 311 79 319 96
rect 283 74 319 79
rect -51 43 43 48
rect -7 24 43 43
rect 173 25 223 55
rect -147 -25 -97 -12
rect -7 -25 43 -12
rect 173 -25 223 -12
<< polycont >>
rect -43 48 -26 65
rect 294 79 311 96
<< locali >>
rect 294 96 311 104
rect -170 78 -153 86
rect -210 56 -193 60
rect -210 22 -193 24
rect -100 62 -91 79
rect -74 65 150 79
rect -74 62 -43 65
rect -170 50 -153 61
rect -52 48 -43 62
rect -26 62 150 65
rect 167 62 175 79
rect 221 62 229 79
rect 246 62 258 79
rect 294 69 311 79
rect -26 48 -18 62
rect 294 52 300 69
rect 294 48 311 52
rect -52 44 -18 48
rect -170 18 -153 33
rect 287 22 304 30
rect -170 -7 -153 1
rect -100 0 -91 17
rect -73 1 -72 17
rect 199 17 223 21
rect -55 1 -30 17
rect -73 0 -30 1
rect -13 0 -4 17
rect 41 0 49 17
rect 66 0 128 17
rect 145 0 150 17
rect 167 0 175 17
rect 199 0 203 17
rect 220 0 229 17
rect 246 0 256 17
rect 199 -3 223 0
<< viali >>
rect -210 60 -193 77
rect -210 39 -193 41
rect -210 24 -193 39
rect -210 -12 -193 5
rect -170 33 -153 50
rect 300 52 317 69
rect -72 1 -55 18
rect 128 0 145 17
rect 203 0 220 17
rect 287 -12 304 5
<< metal1 >>
rect -174 89 -149 124
rect -213 77 -149 89
rect -213 60 -210 77
rect -193 60 -149 77
rect -213 50 -149 60
rect -213 41 -170 50
rect -213 24 -210 41
rect -193 33 -170 41
rect -153 33 -149 50
rect -193 24 -149 33
rect -213 5 -149 24
rect -59 22 -25 25
rect -59 21 -54 22
rect -213 -12 -210 5
rect -193 -12 -149 5
rect -81 18 -54 21
rect -81 1 -72 18
rect -55 1 -54 18
rect -81 -2 -54 1
rect -59 -4 -54 -2
rect -28 17 -25 22
rect 125 17 148 125
rect 260 31 279 125
rect 293 74 325 75
rect 293 48 296 74
rect 322 48 325 74
rect 293 47 325 48
rect -28 0 -13 17
rect 125 0 128 17
rect 145 0 148 17
rect -28 -4 -25 0
rect -59 -7 -25 -4
rect -213 -18 -149 -12
rect -174 -40 -149 -18
rect 125 -40 148 0
rect 184 22 221 23
rect 184 -4 187 22
rect 213 17 226 22
rect 220 0 226 17
rect 213 -4 226 0
rect 260 5 307 31
rect 184 -6 221 -4
rect 260 -12 287 5
rect 304 -12 307 5
rect 260 -18 307 -12
rect 260 -40 279 -18
<< via1 >>
rect -54 -4 -28 22
rect 296 69 322 74
rect 296 52 300 69
rect 300 52 317 69
rect 317 52 322 69
rect 296 48 322 52
rect 187 17 213 22
rect 187 0 203 17
rect 203 0 213 17
rect 187 -4 213 0
<< metal2 >>
rect 292 74 326 76
rect 292 48 296 74
rect 322 69 326 74
rect 322 48 336 69
rect 292 46 336 48
rect 184 22 216 25
rect -57 -4 -54 22
rect -28 17 -25 22
rect 184 17 187 22
rect -28 -2 187 17
rect -28 -4 -25 -2
rect 184 -4 187 -2
rect 213 -4 216 22
rect 184 -7 216 -4
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1628285143
transform 1 0 266 0 1 65
box -10 -8 13 21
<< end >>
