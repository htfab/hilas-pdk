magic
tech sky130A
timestamp 1632398358
<< error_s >>
rect -87 240 -60 246
rect -87 198 -60 204
rect -87 173 -60 179
rect -87 131 -60 137
rect -87 90 -60 96
rect -87 48 -60 54
rect -87 23 -60 29
rect -87 -19 -60 -13
<< metal1 >>
rect -41 -22 -7 550
rect 26 -21 53 549
<< metal2 >>
rect -136 211 155 233
rect -137 -6 134 17
use sky130_hilas_pFETmirror02  sky130_hilas_pFETmirror02_0
timestamp 1629420194
transform 1 0 88 0 1 -111
box -61 89 67 373
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_1
timestamp 1629420194
transform 1 0 -113 0 1 130
box -59 -6 125 123
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_0
timestamp 1629420194
transform 1 0 -113 0 -1 97
box -59 -6 125 123
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1629420194
transform 1 0 106 0 1 228
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1629420194
transform 1 0 98 0 1 3
box -14 -15 20 18
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1629420194
transform 1 0 41 0 1 126
box -10 -8 13 21
<< labels >>
rlabel space 144 211 155 234 0 output2
<< end >>
