magic
tech sky130A
timestamp 1628704362
<< metal1 >>
rect 1167 35561 1231 35955
rect 0 35079 81 35469
rect 1167 32703 1231 33097
rect 0 32220 81 32610
rect 1168 29842 1232 30236
rect 0 29361 81 29751
rect 1167 26984 1231 27378
rect 1 26502 82 26892
rect 1168 24126 1232 24520
rect 0 23643 81 24033
rect 1167 21267 1231 21661
rect 0 20784 81 21174
rect 1167 18408 1231 18802
rect 0 17926 81 18316
rect 1167 15548 1231 15942
rect 2 15067 83 15457
rect 1167 12689 1231 13083
rect 1 12207 82 12597
rect 1166 9832 1230 10226
rect 1 9348 82 9738
rect 1166 6972 1230 7366
rect 1 6489 82 6879
rect 1168 4112 1232 4506
rect 2 3630 83 4020
rect 1168 1255 1232 1649
rect 0 771 81 1161
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_0
timestamp 1627735001
transform 0 -1 939 1 0 745
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_1
timestamp 1627735001
transform 0 -1 939 1 0 3604
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_2
timestamp 1627735001
transform 0 -1 939 1 0 6463
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_3
timestamp 1627735001
transform 0 -1 939 1 0 9322
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_4
timestamp 1627735001
transform 0 -1 939 1 0 12181
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_6
timestamp 1627735001
transform 0 -1 939 1 0 15040
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_9
timestamp 1627735001
transform 0 -1 939 1 0 17899
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_7
timestamp 1627735001
transform 0 -1 939 1 0 20758
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_8
timestamp 1627735001
transform 0 -1 939 1 0 23617
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_5
timestamp 1627735001
transform 0 -1 939 1 0 26476
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_10
timestamp 1627735001
transform 0 -1 939 1 0 29335
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_11
timestamp 1627735001
transform 0 -1 939 1 0 32194
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_12
timestamp 1627735001
transform 0 -1 939 1 0 35053
box -745 -229 2114 858
<< labels >>
rlabel metal1 0 35079 81 35469 0 IO25
port 1 nsew
rlabel metal1 0 32220 81 32610 0 IO26
port 2 nsew
rlabel metal1 0 29361 81 29751 0 IO27
port 3 nsew
rlabel metal1 1 26502 82 26892 0 IO28
port 4 nsew
rlabel metal1 0 23643 81 24033 0 IO29
port 5 nsew
rlabel metal1 0 20784 81 21174 0 IO30
port 6 nsew
rlabel metal1 0 17926 81 18316 0 IO31
port 7 nsew
rlabel metal1 2 15067 83 15457 0 IO32
port 8 nsew
rlabel metal1 1 12207 82 12597 0 IO33
port 9 nsew
rlabel metal1 1 9348 82 9738 0 IO34
port 10 nsew
rlabel metal1 1 6489 82 6879 0 IO35
port 11 nsew
rlabel metal1 2 3630 83 4020 0 IO36
port 12 nsew
rlabel metal1 0 771 81 1161 0 IO37
port 13 nsew
rlabel metal1 1167 35561 1231 35955 0 PIN1
port 14 nsew
rlabel metal1 1167 32703 1231 33097 0 PIN2
port 15 nsew
rlabel metal1 1168 29842 1232 30236 0 PIN3
rlabel metal1 1167 26984 1231 27378 0 PIN4
port 16 nsew
rlabel metal1 1168 24126 1232 24520 0 PIN5
port 17 nsew
rlabel metal1 1167 21267 1231 21661 0 PIN6
port 18 nsew
rlabel metal1 1167 18408 1231 18802 0 PIN7
port 19 nsew
rlabel metal1 1167 15548 1231 15942 0 PIN8
port 20 nsew
rlabel metal1 1167 12689 1231 13083 0 PIN9
port 21 nsew
rlabel metal1 1166 9832 1230 10226 0 PIN10
port 22 nsew
rlabel metal1 1166 6972 1230 7366 0 PIN11
port 23 nsew
rlabel metal1 1168 4112 1232 4506 0 PIN12
port 24 nsew
rlabel metal1 1168 1255 1232 1649 0 PIN13
port 25 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
