magic
tech sky130A
timestamp 1628704268
<< metal1 >>
rect 1 18408 72 18804
rect 1156 17926 1228 18315
rect 0 15548 70 15944
rect 1156 15067 1228 15456
rect 2 12689 72 13085
rect 1156 12207 1228 12596
rect 0 9830 70 10226
rect 1156 9350 1228 9739
rect 0 6970 70 7366
rect 1155 6490 1227 6879
rect 1 4112 71 4508
rect 1156 3631 1228 4020
rect 1 1252 71 1648
rect 1156 771 1228 1160
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_9
timestamp 1627735001
transform 0 1 299 1 0 745
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_7
timestamp 1627735001
transform 0 1 299 1 0 3604
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_8
timestamp 1627735001
transform 0 1 299 1 0 6463
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_5
timestamp 1627735001
transform 0 1 299 1 0 9322
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_10
timestamp 1627735001
transform 0 1 299 1 0 12181
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_11
timestamp 1627735001
transform 0 1 299 1 0 15040
box -745 -229 2114 858
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_12
timestamp 1627735001
transform 0 1 299 1 0 17899
box -745 -229 2114 858
<< labels >>
rlabel metal1 1156 771 1228 1160 0 IO7
port 1 nsew
rlabel metal1 1156 3631 1228 4020 0 IO8
port 2 nsew
rlabel metal1 1155 6490 1227 6879 0 IO9
port 3 nsew
rlabel metal1 1156 9350 1228 9739 0 IO10
port 4 nsew
rlabel metal1 1156 12207 1228 12596 0 IO11
port 5 nsew
rlabel metal1 1156 15067 1228 15456 0 IO12
port 7 nsew
rlabel metal1 1156 17926 1228 18315 0 IO13
port 6 nsew
rlabel metal1 1 1252 71 1648 0 PIN1
port 8 nsew
rlabel metal1 1 4112 71 4508 0 PIN2
port 9 nsew
rlabel metal1 0 6970 70 7366 0 PIN3
port 10 nsew
rlabel metal1 0 9830 70 10226 0 PIN4
port 11 nsew
rlabel metal1 2 12689 72 13085 0 PIN5
port 12 nsew
rlabel metal1 0 15548 70 15944 0 PIN6
port 13 nsew
rlabel metal1 1 18408 71 18804 0 PIN7
port 14 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
