magic
tech sky130A
timestamp 1608234847
<< nwell >>
rect 401 -87 455 159
rect 383 -132 455 -87
rect 198 -150 455 -132
<< psubdiff >>
rect 397 368 439 375
rect 397 351 410 368
rect 427 351 439 368
rect 397 344 439 351
<< nsubdiff >>
rect 396 -110 437 -105
rect 396 -127 408 -110
rect 425 -127 437 -110
rect 396 -132 437 -127
<< psubdiffcont >>
rect 410 351 427 368
<< nsubdiffcont >>
rect 408 -127 425 -110
<< locali >>
rect 411 376 428 381
rect 410 373 428 376
rect 410 368 453 373
rect 427 351 453 368
rect 410 348 453 351
rect 410 342 427 348
rect 396 -127 408 -110
rect 425 -127 438 -110
<< metal1 >>
rect 409 -150 431 438
rect 449 -150 471 438
<< metal2 >>
rect 191 398 198 415
rect 389 399 471 416
rect 191 357 198 374
rect 191 306 198 323
rect 389 307 471 324
rect 191 265 198 282
rect 191 214 198 231
rect 389 215 471 232
rect 191 173 198 190
rect 191 112 198 131
rect 391 105 471 125
rect 191 70 198 89
rect 191 16 198 35
rect 391 9 471 29
rect 191 -26 198 -7
rect 191 -80 198 -61
rect 390 -87 471 -67
rect 191 -122 198 -103
use sky130_hilas_nFET03a  sky130_hilas_nFET03a_3
timestamp 1608056777
transform 1 0 309 0 1 396
box -111 -47 97 42
use sky130_hilas_nFET03a  sky130_hilas_nFET03a_1
timestamp 1608056777
transform 1 0 309 0 1 304
box -111 -47 97 42
use sky130_hilas_nFET03a  sky130_hilas_nFET03a_0
timestamp 1608056777
transform 1 0 309 0 1 212
box -111 -47 97 42
use sky130_hilas_pFETdevice01e  sky130_hilas_pFETdevice01e_2
timestamp 1608055794
transform 1 0 319 0 1 -77
box -121 -55 82 44
use sky130_hilas_pFETdevice01e  sky130_hilas_pFETdevice01e_1
timestamp 1608055794
transform 1 0 319 0 1 19
box -121 -55 82 44
use sky130_hilas_pFETdevice01e  sky130_hilas_pFETdevice01e_0
timestamp 1608055794
transform 1 0 319 0 1 115
box -121 -55 82 44
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1607179295
transform 0 1 411 -1 0 -120
box -10 -8 13 21
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1607179295
transform 1 0 458 0 1 354
box -10 -8 13 21
<< labels >>
rlabel metal1 409 -150 431 -141 0 Well
port 13 nsew power default
rlabel metal1 449 -150 471 -141 0 GND
port 14 nsew ground default
rlabel metal1 409 429 431 438 0 Well
port 13 nsew ground default
rlabel metal1 449 429 471 438 0 GND
port 14 nsew power default
rlabel metal2 191 398 198 415 0 nFET_Source1
port 1 nsew analog default
rlabel metal2 191 357 198 374 0 nFET_Gate1
port 2 nsew analog default
rlabel metal2 191 306 198 323 0 nFET_Source2
port 3 nsew analog default
rlabel metal2 191 265 198 282 0 nFET_Gate2
port 4 nsew analog default
rlabel metal2 191 214 198 231 0 nFET_Source3
port 5 nsew analog default
rlabel metal2 191 173 198 190 0 nFET_Gate3
port 6 nsew analog default
rlabel metal2 191 70 198 89 0 pFET_Gate1
port 8 nsew analog default
rlabel metal2 191 112 198 131 0 pFET_Source1
port 7 nsew analog default
rlabel metal2 191 16 198 35 0 pFET_Source2
port 9 nsew analog default
rlabel metal2 191 -26 198 -7 0 pFET_Gate2
port 10 nsew analog default
rlabel metal2 191 -80 198 -61 0 pFET_Source3
port 11 nsew analog default
rlabel metal2 191 -122 198 -103 0 pFET_Gate3
port 12 nsew analog default
rlabel metal2 465 105 471 125 0 pFET_Drain1
port 17 nsew analog default
rlabel metal2 465 9 471 29 0 pFET_Drain2
port 16 nsew analog default
rlabel metal2 465 -87 471 -67 0 pFET_Drain3
port 15 nsew analog default
rlabel metal2 466 399 471 416 0 nFET_Drain1
port 20 nsew analog default
rlabel metal2 466 307 471 324 0 nFET_Drain2
port 19 nsew analog default
rlabel metal2 466 215 471 232 0 nFET_Drain3
port 18 nsew analog default
<< end >>
