* NGSPICE file created from /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_TACoreBlock.ext - technology: sky130A

.subckt sky130_hilas_TunCap01 $SUB
X0 a_n2872_n666# w_n2902_n800# w_n2902_n800# sky130_fd_pr__cap_var w=590000u l=500000u
.ends

.subckt sky130_hilas_horizPcell01 $SUB
X0 w_n578_94# a_n300_94# a_n344_162# w_n578_94# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
X1 a_n344_286# a_n578_238# a_n502_286# w_n578_94# sky130_fd_pr__pfet_g5v0d10v5 w=300000u l=500000u
X2 a_n344_162# a_n578_238# a_n508_162# w_n578_94# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
.ends

.subckt sky130_hilas_FGVaractorCapacitor $SUB
X0 a_n1882_n672# w_n1914_n790# w_n1914_n790# sky130_fd_pr__cap_var w=1.11e+06u l=640000u
.ends


* Top level circuit /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_TACoreBlock

Xsky130_hilas_TunCap01_0 $SUB sky130_hilas_TunCap01
Xsky130_hilas_horizPcell01_0 $SUB sky130_hilas_horizPcell01
Xsky130_hilas_FGVaractorCapacitor_0 $SUB sky130_hilas_FGVaractorCapacitor
X0 a_n16_78# a_n42_20# a_n16_n38# $SUB sky130_fd_pr__nfet_01v8 w=330000u l=290000u
.end

