VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_fgtrans2x1cell
  CLASS BLOCK ;
  FOREIGN sky130_hilas_fgtrans2x1cell ;
  ORIGIN 3.950 3.820 ;
  SIZE 11.520 BY 6.050 ;
  OBS
      LAYER nwell ;
        RECT -3.370 -2.420 -2.810 0.000 ;
      LAYER li1 ;
        RECT 3.860 1.630 4.740 1.800 ;
        RECT 3.860 1.240 4.030 1.630 ;
        RECT 3.640 1.070 4.030 1.240 ;
        RECT 4.440 1.070 4.660 1.240 ;
        RECT 2.210 0.280 3.290 0.450 ;
        RECT 3.620 0.280 4.700 0.450 ;
        RECT -0.920 -0.750 -0.730 -0.340 ;
        RECT 4.640 -0.510 4.720 -0.340 ;
        RECT -0.920 -0.930 2.630 -0.750 ;
        RECT -0.920 -1.350 -0.730 -0.930 ;
        RECT 3.380 -1.080 3.550 -0.510 ;
        RECT 3.560 -1.110 3.640 -1.100 ;
        RECT 4.220 -1.110 4.270 -1.100 ;
        RECT 3.560 -1.150 4.270 -1.110 ;
        RECT 3.540 -1.190 4.270 -1.150 ;
        RECT 3.470 -1.310 4.310 -1.190 ;
        RECT 4.640 -1.250 4.690 -1.080 ;
        RECT 2.060 -2.040 3.300 -1.870 ;
        RECT 3.620 -2.040 4.700 -1.870 ;
        RECT 2.800 -2.360 2.970 -2.300 ;
        RECT 2.780 -2.570 2.990 -2.360 ;
        RECT 2.800 -2.640 2.970 -2.570 ;
        RECT 3.640 -2.670 4.100 -2.660 ;
        RECT 3.630 -2.820 4.100 -2.670 ;
        RECT 3.640 -2.830 4.100 -2.820 ;
        RECT 4.450 -2.830 4.660 -2.660 ;
        RECT 3.910 -3.170 4.100 -2.830 ;
        RECT 3.910 -3.350 4.870 -3.170 ;
      LAYER met1 ;
        RECT -3.610 -3.810 -3.190 2.230 ;
        RECT -1.130 -3.820 -0.900 2.230 ;
        RECT 2.790 -2.300 2.970 2.230 ;
        RECT 2.740 -2.640 3.030 -2.300 ;
        RECT 2.790 -3.820 2.970 -2.640 ;
        RECT 3.840 -3.820 4.050 2.230 ;
        RECT 4.270 -3.810 4.460 2.230 ;
        RECT 4.720 -0.560 4.930 2.220 ;
        RECT 6.210 -1.010 6.450 -0.590 ;
        RECT 4.720 -3.320 4.910 -1.070 ;
        RECT 5.220 -3.320 5.230 -3.310 ;
        RECT 4.690 -3.810 4.920 -3.320 ;
      LAYER met2 ;
        RECT 4.840 1.730 5.160 1.750 ;
        RECT -3.950 1.550 5.160 1.730 ;
        RECT -3.950 0.000 2.690 0.190 ;
        RECT -3.950 -0.730 6.210 -0.690 ;
        RECT -3.950 -0.920 6.220 -0.730 ;
        RECT -3.950 -1.860 2.700 -1.670 ;
        RECT 5.100 -3.150 5.260 -3.130 ;
        RECT -3.950 -3.200 5.260 -3.150 ;
        RECT -3.950 -3.300 5.140 -3.200 ;
  END
END sky130_hilas_fgtrans2x1cell
END LIBRARY

