* Copyright 2020 The Hilas PDK Authors
* 
* This file is part of HILAS.
* 
* HILAS is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published by
* the Free Software Foundation, version 3 of the License.
* 
* HILAS is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
* 
* You should have received a copy of the GNU Lesser General Public License
* along with HILAS.  If not, see <https://www.gnu.org/licenses/>.
* 
* Licensed under the Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
* https://www.gnu.org/licenses/lgpl-3.0.en.html
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
* SPDX-License-Identifier: LGPL-3.0
* 
* 

* NGSPICE file created from sky130_hilas_nFETLargePart1.ext - technology: sky130A

.subckt sky130_hilas_nFETmed a_84_n62# $SUB a_n24_n62#
X0 a_84_n62# a_32_n88# a_n24_n62# $SUB sky130_fd_pr__nfet_01v8 w=2.46e+06u l=260000u
.ends


* Top level circuit sky130_hilas_nFETLargePart1

Xsky130_hilas_nFETmed_0 sky130_hilas_nFETmed_0/a_84_n62# $SUB sky130_hilas_nFETmed_4/a_84_n62#
+ sky130_hilas_nFETmed
Xsky130_hilas_nFETmed_1 sky130_hilas_nFETmed_1/a_84_n62# $SUB sky130_hilas_nFETmed_0/a_84_n62#
+ sky130_hilas_nFETmed
Xsky130_hilas_nFETmed_2 sky130_hilas_nFETmed_2/a_84_n62# $SUB sky130_hilas_nFETmed_1/a_84_n62#
+ sky130_hilas_nFETmed
Xsky130_hilas_nFETmed_3 sky130_hilas_nFETmed_3/a_84_n62# $SUB sky130_hilas_nFETmed_2/a_84_n62#
+ sky130_hilas_nFETmed
Xsky130_hilas_nFETmed_4 sky130_hilas_nFETmed_4/a_84_n62# $SUB sky130_hilas_nFETmed_4/a_n24_n62#
+ sky130_hilas_nFETmed
.end

