magic
tech sky130A
magscale 1 2
timestamp 1632256360
<< error_s >>
rect 2014 876 2182 910
rect 2216 890 2370 1034
rect 2780 1000 2792 1288
rect 2960 1272 2971 1279
rect 2914 1268 2971 1272
rect 3004 1268 3102 1294
rect 3313 1268 3324 1279
rect 2914 1260 3324 1268
rect 2914 1240 3004 1260
rect 3102 1246 3324 1260
rect 3406 1240 3446 1272
rect 2914 1172 2915 1173
rect 2960 1172 3004 1240
rect 3102 1172 3324 1240
rect 3445 1172 3446 1173
rect 2814 1114 2850 1172
rect 2913 1171 3004 1172
rect 2914 1156 3004 1171
rect 2914 1128 2934 1156
rect 2960 1128 3004 1156
rect 3072 1146 3324 1172
rect 3388 1171 3447 1172
rect 3388 1156 3446 1171
rect 3388 1146 3406 1156
rect 3102 1128 3324 1146
rect 3428 1128 3446 1156
rect 2914 1116 3004 1128
rect 2914 1115 2960 1116
rect 3072 1115 3324 1128
rect 3388 1115 3446 1128
rect 2913 1114 2960 1115
rect 2972 1114 2973 1115
rect 3071 1114 3324 1115
rect 3387 1114 3447 1115
rect 3512 1114 3546 1172
rect 5616 1154 5650 1186
rect 5616 1144 5670 1154
rect 5600 1138 5670 1144
rect 5600 1114 5634 1138
rect 5738 1116 5754 1164
rect 5766 1132 5782 1184
rect 5896 1152 5934 1186
rect 5896 1144 5946 1152
rect 5874 1138 5946 1144
rect 5874 1116 5908 1138
rect 2914 1113 2915 1114
rect 2971 1113 2972 1114
rect 3072 1113 3073 1114
rect 3102 1096 3324 1114
rect 3388 1113 3389 1114
rect 3445 1113 3446 1114
rect 5592 1104 5634 1114
rect 5872 1104 5914 1116
rect 2960 1058 3324 1096
rect 2960 1044 3004 1058
rect 3102 1044 3324 1058
rect 2914 1016 3004 1044
rect 2914 1014 2972 1016
rect 2960 1005 2971 1014
rect 2993 1005 3004 1016
rect 3072 1014 3102 1044
rect 3388 1014 3446 1044
rect 2780 978 3580 1000
rect 5270 984 5322 986
rect 2416 910 2452 912
rect 2498 910 2558 930
rect 2416 890 2466 904
rect 2216 876 2538 890
rect 2072 746 2538 876
rect 2558 782 2568 834
rect 2894 828 3438 978
rect 5144 960 5196 984
rect 5228 950 5298 952
rect 5228 938 5326 950
rect 5228 928 5322 938
rect 5228 920 5246 928
rect 5256 904 5320 924
rect 5256 892 5274 904
rect 5302 884 5320 904
rect 5256 860 5320 884
rect 5244 832 5298 856
rect 5302 814 5310 860
rect 5330 832 5348 952
rect 5366 928 5390 1052
rect 5486 928 5550 946
rect 5634 938 5696 946
rect 5522 922 5544 928
rect 5634 924 5698 938
rect 5768 926 5832 946
rect 5804 920 5826 926
rect 5458 900 5578 918
rect 5606 910 5724 918
rect 5522 894 5572 900
rect 5606 896 5726 910
rect 5740 898 5860 918
rect 5804 894 5816 898
rect 5804 892 5826 894
rect 5330 786 5338 832
rect 5602 828 5734 848
rect 5816 830 5826 838
rect 5636 806 5700 814
rect 5636 794 5702 806
rect 5816 802 5826 810
rect 2072 640 2548 746
rect 2698 680 2742 754
rect 2072 638 2182 640
rect 2014 600 2182 638
rect 2324 638 2548 640
rect 2780 638 2792 746
rect 2914 680 2972 712
rect 3072 680 3130 712
rect 3230 680 3288 712
rect 3388 680 3446 712
rect 5144 698 5208 716
rect 5242 698 5270 716
rect 2324 636 2538 638
rect 2326 600 2370 636
rect 2380 604 2538 636
rect 2850 612 2894 680
rect 5144 676 5196 698
rect 5283 683 5322 698
rect 5270 666 5296 668
rect 5298 666 5322 683
rect 5208 652 5253 666
rect 5270 642 5322 666
rect 2914 612 2915 613
rect 2971 612 2972 613
rect 3072 612 3073 613
rect 3129 612 3130 613
rect 3230 612 3231 613
rect 3287 612 3288 613
rect 3388 612 3389 613
rect 3445 612 3446 613
rect 2380 600 2494 604
rect 2116 598 2182 600
rect 2814 554 2894 612
rect 2913 611 2973 612
rect 3071 611 3131 612
rect 3229 611 3289 612
rect 3387 611 3447 612
rect 2914 596 2972 611
rect 3072 596 3130 611
rect 3230 596 3288 611
rect 3388 596 3446 611
rect 2914 568 2934 596
rect 3428 568 3446 596
rect 2914 555 2972 568
rect 3072 555 3130 568
rect 3230 555 3288 568
rect 3388 555 3446 568
rect 2913 554 2973 555
rect 3071 554 3131 555
rect 3229 554 3289 555
rect 3387 554 3447 555
rect 3512 554 3546 612
rect 5332 554 5354 570
rect 278 494 336 530
rect 278 430 279 431
rect 335 430 336 431
rect 178 372 214 430
rect 277 429 337 430
rect 278 410 336 429
rect 278 392 298 410
rect 316 392 336 410
rect 278 373 336 392
rect 277 372 337 373
rect 400 372 436 430
rect 950 424 994 504
rect 278 371 279 372
rect 335 371 336 372
rect 884 358 1060 424
rect 2698 370 2742 486
rect 2850 484 2894 554
rect 2914 553 2915 554
rect 2971 553 2972 554
rect 3072 553 3073 554
rect 3129 553 3130 554
rect 3230 553 3231 554
rect 3287 553 3288 554
rect 3388 553 3389 554
rect 3445 553 3446 554
rect 5740 552 5860 562
rect 5768 524 5832 534
rect 2914 454 2972 484
rect 3072 454 3130 484
rect 3230 454 3288 484
rect 3388 454 3446 484
rect 2914 370 2972 402
rect 3072 370 3130 402
rect 3230 370 3288 402
rect 3388 370 3446 402
rect 5256 398 5272 432
rect 5292 428 5306 434
rect 5290 390 5306 428
rect 5292 382 5306 390
rect 5360 376 5378 384
rect 884 336 1118 358
rect 278 272 336 308
rect 884 270 1060 336
rect 2850 302 2894 370
rect 5586 354 5608 388
rect 5620 384 5642 422
rect 5610 362 5664 384
rect 2914 302 2915 303
rect 2971 302 2972 303
rect 3072 302 3073 303
rect 3129 302 3130 303
rect 3230 302 3231 303
rect 3287 302 3288 303
rect 3388 302 3389 303
rect 3445 302 3446 303
rect 2814 244 2894 302
rect 2913 301 2973 302
rect 3071 301 3131 302
rect 3229 301 3289 302
rect 3387 301 3447 302
rect 2914 286 2972 301
rect 3072 286 3130 301
rect 3230 286 3288 301
rect 3388 286 3446 301
rect 2914 258 2934 286
rect 3428 258 3446 286
rect 2914 245 2972 258
rect 3072 245 3130 258
rect 3230 245 3288 258
rect 3388 245 3446 258
rect 2913 244 2973 245
rect 3071 244 3131 245
rect 3229 244 3289 245
rect 3387 244 3447 245
rect 3512 244 3546 302
rect 2850 174 2894 244
rect 2914 243 2915 244
rect 2971 243 2972 244
rect 3072 243 3073 244
rect 3129 243 3130 244
rect 3230 243 3231 244
rect 3287 243 3288 244
rect 3388 243 3389 244
rect 3445 243 3446 244
rect 5352 200 5414 218
rect 5638 196 5700 218
rect 2914 144 2972 174
rect 3072 144 3130 174
rect 3230 144 3288 174
rect 3388 144 3446 174
rect 5324 172 5442 190
rect 5610 168 5728 190
rect 5156 124 5158 134
rect 5388 92 5390 120
rect 5536 92 5538 120
rect 5676 92 5678 120
rect 5180 78 5206 84
rect 5322 80 5380 84
rect 5388 58 5424 86
rect 5536 58 5572 86
rect 5676 58 5712 86
rect 5152 50 5206 56
rect 5294 52 5352 56
<< nwell >>
rect 1776 876 2006 910
rect 2014 876 2116 910
rect 1738 640 2538 876
rect 1738 638 2116 640
rect 2380 638 2538 640
rect 1776 600 2006 638
rect 2014 598 2116 638
rect 2326 600 2380 636
rect 5366 500 5914 1200
rect 950 336 994 358
<< mvnmos >>
rect 5144 1010 5270 1110
rect 5144 566 5270 666
rect 5144 232 5268 386
rect 5434 232 5562 342
rect 5718 232 5846 342
<< mvpmos >>
rect 5440 958 5560 1068
rect 5720 958 5840 1068
rect 5440 624 5560 734
rect 5720 624 5840 734
<< mvndiff >>
rect 5144 1156 5270 1164
rect 5144 1122 5156 1156
rect 5190 1122 5224 1156
rect 5258 1122 5270 1156
rect 5144 1110 5270 1122
rect 5144 984 5270 1010
rect 5144 666 5270 676
rect 5144 554 5270 566
rect 5144 520 5154 554
rect 5188 520 5222 554
rect 5256 520 5270 554
rect 5144 508 5270 520
rect 5144 432 5268 448
rect 5144 398 5154 432
rect 5188 398 5222 432
rect 5256 398 5268 432
rect 5144 386 5268 398
rect 5434 388 5562 402
rect 5434 354 5448 388
rect 5482 354 5516 388
rect 5550 354 5562 388
rect 5434 342 5562 354
rect 5718 388 5846 400
rect 5718 354 5730 388
rect 5764 354 5798 388
rect 5832 354 5846 388
rect 5718 342 5846 354
rect 5144 220 5268 232
rect 5144 186 5152 220
rect 5186 186 5220 220
rect 5254 186 5268 220
rect 5144 172 5268 186
rect 5434 220 5562 232
rect 5434 186 5448 220
rect 5482 186 5516 220
rect 5550 186 5562 220
rect 5434 172 5562 186
rect 5718 220 5846 232
rect 5718 186 5730 220
rect 5764 186 5798 220
rect 5832 186 5846 220
rect 5718 174 5846 186
<< mvpdiff >>
rect 5440 1114 5560 1126
rect 5440 1080 5448 1114
rect 5482 1080 5516 1114
rect 5550 1080 5560 1114
rect 5440 1068 5560 1080
rect 5720 1114 5840 1126
rect 5720 1080 5730 1114
rect 5764 1080 5798 1114
rect 5832 1080 5840 1114
rect 5720 1068 5840 1080
rect 5440 944 5560 958
rect 5440 910 5448 944
rect 5482 910 5516 944
rect 5550 910 5560 944
rect 5440 876 5560 910
rect 5440 780 5560 816
rect 5440 746 5448 780
rect 5482 746 5516 780
rect 5550 746 5560 780
rect 5440 734 5560 746
rect 5720 944 5840 958
rect 5720 910 5730 944
rect 5764 910 5798 944
rect 5832 910 5840 944
rect 5720 876 5840 910
rect 5720 780 5840 816
rect 5720 746 5730 780
rect 5764 746 5798 780
rect 5832 746 5840 780
rect 5720 734 5840 746
rect 5440 612 5560 624
rect 5440 578 5448 612
rect 5482 578 5516 612
rect 5550 578 5560 612
rect 5440 566 5560 578
rect 5720 612 5840 624
rect 5720 578 5730 612
rect 5764 578 5798 612
rect 5832 578 5840 612
rect 5720 566 5840 578
<< mvndiffc >>
rect 5156 1122 5190 1156
rect 5224 1122 5258 1156
rect 5154 520 5188 554
rect 5222 520 5256 554
rect 5154 398 5188 432
rect 5222 398 5256 432
rect 5448 354 5482 388
rect 5516 354 5550 388
rect 5730 354 5764 388
rect 5798 354 5832 388
rect 5152 186 5186 220
rect 5220 186 5254 220
rect 5448 186 5482 220
rect 5516 186 5550 220
rect 5730 186 5764 220
rect 5798 186 5832 220
<< mvpdiffc >>
rect 5448 1080 5482 1114
rect 5516 1080 5550 1114
rect 5730 1080 5764 1114
rect 5798 1080 5832 1114
rect 5448 910 5482 944
rect 5516 910 5550 944
rect 5448 746 5482 780
rect 5516 746 5550 780
rect 5730 910 5764 944
rect 5798 910 5832 944
rect 5730 746 5764 780
rect 5798 746 5832 780
rect 5448 578 5482 612
rect 5516 578 5550 612
rect 5730 578 5764 612
rect 5798 578 5832 612
<< psubdiff >>
rect 702 756 1370 766
rect 702 722 782 756
rect 816 722 850 756
rect 884 722 918 756
rect 952 722 986 756
rect 1020 722 1054 756
rect 1088 722 1122 756
rect 1156 722 1190 756
rect 1224 722 1258 756
rect 1292 722 1370 756
rect 702 714 1370 722
rect 702 676 760 714
rect 702 642 714 676
rect 748 642 760 676
rect 702 618 760 642
rect 470 608 760 618
rect 470 592 714 608
rect 470 558 510 592
rect 544 558 578 592
rect 612 558 646 592
rect 680 574 714 592
rect 748 574 760 608
rect 680 558 760 574
rect 470 542 760 558
rect 702 540 760 542
rect 702 506 714 540
rect 748 506 760 540
rect 702 472 760 506
rect 702 438 714 472
rect 748 438 760 472
rect 702 404 760 438
rect 702 370 714 404
rect 748 370 760 404
rect 702 336 760 370
rect 2664 688 2742 754
rect 2664 654 2688 688
rect 2722 654 2742 688
rect 2664 596 2742 654
rect 2664 562 2688 596
rect 2722 562 2742 596
rect 2664 520 2742 562
rect 2664 486 2688 520
rect 2722 486 2742 520
rect 2664 434 2742 486
rect 2664 400 2688 434
rect 2722 400 2742 434
rect 702 302 714 336
rect 748 302 760 336
rect 702 268 760 302
rect 702 234 714 268
rect 748 234 760 268
rect 702 200 760 234
rect 702 166 714 200
rect 748 166 760 200
rect 2664 324 2742 400
rect 2664 290 2688 324
rect 2722 290 2742 324
rect 2664 244 2742 290
rect 2664 210 2688 244
rect 2722 210 2742 244
rect 702 142 760 166
rect 2664 172 2742 210
rect 2664 138 2688 172
rect 2722 138 2742 172
rect 2664 96 2742 138
rect 2664 62 2686 96
rect 2720 62 2742 96
rect 2664 30 2742 62
<< mvpsubdiff >>
rect 5146 86 5854 98
rect 5146 84 5306 86
rect 5146 50 5170 84
rect 5204 50 5238 84
rect 5272 52 5306 84
rect 5340 52 5378 86
rect 5412 52 5450 86
rect 5484 52 5518 86
rect 5552 52 5586 86
rect 5620 52 5654 86
rect 5688 52 5722 86
rect 5756 52 5790 86
rect 5824 52 5854 86
rect 5272 50 5854 52
rect 5146 38 5854 50
<< mvnsubdiff >>
rect 2390 858 2472 874
rect 2390 832 2414 858
rect 2362 824 2414 832
rect 2448 824 2472 858
rect 2362 790 2472 824
rect 2362 756 2414 790
rect 2448 756 2472 790
rect 2362 754 2472 756
rect 2390 722 2472 754
rect 2390 688 2414 722
rect 2448 688 2472 722
rect 2390 678 2472 688
rect 2392 670 2472 678
rect 5440 862 5560 876
rect 5440 828 5482 862
rect 5516 828 5560 862
rect 5440 816 5560 828
rect 5720 862 5840 876
rect 5720 828 5762 862
rect 5796 828 5840 862
rect 5720 816 5840 828
rect 950 336 994 358
<< psubdiffcont >>
rect 782 722 816 756
rect 850 722 884 756
rect 918 722 952 756
rect 986 722 1020 756
rect 1054 722 1088 756
rect 1122 722 1156 756
rect 1190 722 1224 756
rect 1258 722 1292 756
rect 714 642 748 676
rect 510 558 544 592
rect 578 558 612 592
rect 646 558 680 592
rect 714 574 748 608
rect 714 506 748 540
rect 714 438 748 472
rect 714 370 748 404
rect 2688 654 2722 688
rect 2688 562 2722 596
rect 2688 486 2722 520
rect 2688 400 2722 434
rect 714 302 748 336
rect 714 234 748 268
rect 714 166 748 200
rect 2688 290 2722 324
rect 2688 210 2722 244
rect 2688 138 2722 172
rect 2686 62 2720 96
<< mvpsubdiffcont >>
rect 5170 50 5204 84
rect 5238 50 5272 84
rect 5306 52 5340 86
rect 5378 52 5412 86
rect 5450 52 5484 86
rect 5518 52 5552 86
rect 5586 52 5620 86
rect 5654 52 5688 86
rect 5722 52 5756 86
rect 5790 52 5824 86
<< mvnsubdiffcont >>
rect 2414 824 2448 858
rect 2414 756 2448 790
rect 2414 688 2448 722
rect 5482 828 5516 862
rect 5762 828 5796 862
<< poly >>
rect 352 974 408 1074
rect 358 840 408 974
rect 1396 914 1494 1088
rect 4722 1084 5144 1110
rect 1396 910 1784 914
rect 2350 910 2452 912
rect 2498 910 2890 1084
rect 4720 1010 5144 1084
rect 5270 1010 5296 1110
rect 5592 1112 5608 1144
rect 5592 1068 5632 1112
rect 5874 1110 5892 1144
rect 5868 1068 5904 1110
rect 4720 982 4828 1010
rect 5412 958 5440 1068
rect 5560 958 5632 1068
rect 5688 958 5720 1068
rect 5840 958 5904 1068
rect 1396 840 2088 910
rect 134 792 2088 840
rect 134 434 210 792
rect 1396 600 2088 792
rect 5236 798 5330 866
rect 5298 666 5330 798
rect 5592 734 5632 958
rect 5870 734 5904 958
rect 2350 636 2452 638
rect 2326 600 2452 636
rect 1396 598 1784 600
rect 1986 598 2088 600
rect 1396 348 1494 598
rect 5114 566 5144 666
rect 5270 566 5330 666
rect 5412 624 5440 734
rect 5560 624 5632 734
rect 5692 624 5720 734
rect 5840 624 5904 734
rect 5320 472 5396 474
rect 1396 290 1974 348
rect 5284 396 5396 472
rect 5284 386 5326 396
rect 1396 180 1494 290
rect 5114 232 5144 386
rect 5268 356 5326 386
rect 5268 232 5296 356
rect 5402 232 5434 342
rect 5562 232 5718 342
rect 5846 232 5872 342
<< locali >>
rect 5140 1122 5156 1156
rect 5258 1122 5274 1156
rect 5600 1114 5616 1144
rect 5874 1116 5892 1144
rect 5714 1114 5914 1116
rect 5432 1080 5448 1114
rect 5550 1080 5634 1114
rect 5714 1080 5730 1114
rect 5832 1080 5914 1114
rect 5432 910 5448 944
rect 5550 910 5730 944
rect 5832 910 5848 944
rect 2414 858 2448 874
rect 5448 828 5482 862
rect 5550 828 5728 862
rect 5796 828 5812 862
rect 2414 804 2448 824
rect 2414 790 2534 804
rect 714 756 748 760
rect 2448 756 2534 790
rect 714 722 782 756
rect 816 722 850 756
rect 884 722 918 756
rect 952 722 986 756
rect 1020 722 1054 756
rect 1088 722 1122 756
rect 1156 722 1190 756
rect 1224 722 1258 756
rect 1292 722 1326 756
rect 2414 752 2534 756
rect 2414 722 2448 752
rect 5432 746 5448 780
rect 5550 746 5730 780
rect 5832 746 5848 780
rect 714 676 748 722
rect 2414 672 2448 688
rect 2688 688 2722 710
rect 714 608 748 642
rect 494 558 510 592
rect 544 558 578 592
rect 612 558 646 592
rect 680 574 714 592
rect 680 558 748 574
rect 714 540 748 558
rect 714 472 748 506
rect 714 404 748 438
rect 714 336 748 370
rect 714 268 748 302
rect 714 200 748 234
rect 2688 596 2722 654
rect 5432 578 5448 612
rect 5550 578 5568 612
rect 5714 578 5730 612
rect 5832 578 5848 612
rect 2688 520 2722 562
rect 5138 520 5154 554
rect 5188 520 5222 554
rect 5256 520 5366 554
rect 2688 434 2722 486
rect 2688 324 2722 400
rect 5138 398 5154 432
rect 5256 398 5272 432
rect 5432 354 5448 388
rect 5550 354 5608 388
rect 5714 354 5730 388
rect 5832 354 5848 388
rect 2688 244 2722 290
rect 2688 180 2722 210
rect 5134 186 5152 220
rect 5186 186 5220 220
rect 5254 186 5448 220
rect 5482 186 5516 220
rect 5550 186 5730 220
rect 5764 186 5798 220
rect 5832 186 5850 220
rect 714 76 748 166
rect 2686 172 2722 180
rect 2686 138 2688 172
rect 2686 96 2722 138
rect 2720 62 2722 96
rect 5188 86 5324 96
rect 5188 84 5306 86
rect 2686 34 2722 62
rect 5154 50 5170 84
rect 5204 50 5238 84
rect 5272 52 5306 84
rect 5340 52 5378 86
rect 5412 52 5450 86
rect 5484 52 5518 86
rect 5552 52 5586 86
rect 5620 52 5654 86
rect 5688 52 5722 86
rect 5756 52 5790 86
rect 5824 52 5840 86
rect 5272 50 5324 52
<< viali >>
rect 5190 1122 5224 1156
rect 5482 1080 5516 1114
rect 5764 1080 5798 1114
rect 5482 910 5516 944
rect 5764 910 5798 944
rect 5516 828 5550 862
rect 5728 828 5762 862
rect 5482 746 5516 780
rect 5764 746 5798 780
rect 5482 578 5516 612
rect 5764 578 5798 612
rect 5188 398 5222 432
rect 5482 354 5516 388
rect 5764 354 5798 388
<< metal1 >>
rect 0 1032 52 1210
rect 940 960 994 1210
rect 2114 1128 2162 1210
rect 5178 1156 5236 1162
rect 5178 1122 5190 1156
rect 5224 1122 5236 1156
rect 5178 1116 5236 1122
rect 5330 1114 5536 1130
rect 5330 1080 5482 1114
rect 5516 1080 5536 1114
rect 5330 1068 5536 1080
rect 5742 1114 5818 1130
rect 5742 1080 5764 1114
rect 5798 1080 5818 1114
rect 5742 1068 5818 1080
rect 5180 978 5234 1004
rect 5162 960 5234 978
rect 5162 920 5246 960
rect 5162 732 5208 920
rect 5162 696 5234 732
rect 158 36 208 410
rect 156 0 208 36
rect 938 0 1000 518
rect 5180 438 5234 696
rect 5330 514 5378 1068
rect 5476 944 5522 956
rect 5476 910 5482 944
rect 5516 910 5522 944
rect 5756 944 5804 956
rect 5756 910 5764 944
rect 5798 910 5804 944
rect 5466 862 5816 910
rect 5466 828 5516 862
rect 5550 828 5728 862
rect 5762 828 5816 862
rect 5466 780 5816 828
rect 5466 778 5482 780
rect 5476 746 5482 778
rect 5516 778 5764 780
rect 5516 746 5522 778
rect 5476 734 5522 746
rect 5756 746 5764 778
rect 5798 778 5816 780
rect 5798 746 5804 778
rect 5756 734 5804 746
rect 5476 612 5522 624
rect 5476 578 5482 612
rect 5516 578 5522 612
rect 5168 432 5234 438
rect 5168 398 5188 432
rect 5222 398 5234 432
rect 5168 392 5234 398
rect 5476 388 5522 578
rect 2116 0 2164 376
rect 5476 354 5482 388
rect 5516 354 5522 388
rect 5476 342 5522 354
rect 5758 612 5804 624
rect 5758 578 5764 612
rect 5798 578 5804 612
rect 5758 388 5804 578
rect 5758 354 5764 388
rect 5798 354 5804 388
rect 5758 342 5804 354
rect 4778 0 4836 212
<< metal2 >>
rect 5176 1116 5754 1164
rect 2470 918 5400 944
rect 2470 902 5934 918
rect 2116 762 2176 854
rect 2262 764 2322 856
rect 2538 768 2586 902
rect 5372 868 5934 902
rect 5244 600 5298 856
rect 5400 766 5934 868
rect 5244 598 5802 600
rect 5244 554 5934 598
rect 5348 552 5934 554
rect 5810 456 5934 520
rect 5328 378 5934 424
rect 5158 124 5934 190
rect 5156 106 5934 124
rect 5158 92 5934 106
rect 5206 56 5294 92
rect 706 14 5352 56
use sky130_hilas_pFETdevice01w1  sky130_hilas_pFETdevice01w1_0
timestamp 1632251336
transform 1 0 2216 0 1 792
box 0 0 322 242
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_0
timestamp 1632251362
transform 1 0 178 0 1 272
box 0 0 258 258
use sky130_hilas_li2m2  sky130_hilas_li2m2_14
timestamp 1632251356
transform 1 0 728 0 1 48
box 0 0 68 66
use sky130_hilas_li2m2  sky130_hilas_li2m2_13
timestamp 1632251356
transform 1 0 2146 0 1 790
box 0 0 68 66
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_2
timestamp 1632251432
transform 1 0 2894 0 1 1030
box 0 0 544 338
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_0
timestamp 1632251432
transform 1 0 2894 0 1 828
box 0 0 544 338
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_0
timestamp 1632251342
transform 1 0 2780 0 1 978
box 0 0 800 328
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_2
timestamp 1632251342
transform 1 0 2780 0 1 108
box 0 0 800 328
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_1
timestamp 1632251342
transform 1 0 2780 0 1 418
box 0 0 800 328
use sky130_hilas_li2m2  sky130_hilas_li2m2_11
timestamp 1632251356
transform 1 0 2556 0 1 776
box 0 0 68 66
use sky130_hilas_li2m2  sky130_hilas_li2m2_12
timestamp 1632251356
transform 1 0 2284 0 1 792
box 0 0 68 66
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1632251356
transform 1 0 2700 0 1 44
box 0 0 68 66
use sky130_hilas_li2m2  sky130_hilas_li2m2_9
timestamp 1632251356
transform 1 0 5180 0 1 78
box 0 0 68 66
use sky130_hilas_li2m2  sky130_hilas_li2m2_6
timestamp 1632251356
transform 1 0 5470 0 1 80
box 0 0 68 66
use sky130_hilas_li2m2  sky130_hilas_li2m2_5
timestamp 1632251356
transform 1 0 5322 0 1 80
box 0 0 68 66
use sky130_hilas_li2m2  sky130_hilas_li2m2_4
timestamp 1632251356
transform 1 0 5352 0 1 200
box 0 0 68 66
use sky130_hilas_li2m2  sky130_hilas_li2m2_8
timestamp 1632251356
transform 1 0 5796 0 1 80
box 0 0 68 66
use sky130_hilas_li2m2  sky130_hilas_li2m2_7
timestamp 1632251356
transform 1 0 5610 0 1 80
box 0 0 68 66
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1632251356
transform 1 0 5638 0 1 196
box 0 0 68 66
use sky130_hilas_nDiffThOxContact  sky130_hilas_nDiffThOxContact_3
timestamp 1632251312
transform 1 0 5192 0 1 642
box 0 0 134 58
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1632251332
transform 1 0 5350 0 1 530
box 0 0 46 58
use sky130_hilas_li2m2  sky130_hilas_li2m2_10
timestamp 1632251356
transform -1 0 5358 0 -1 440
box 0 0 68 66
use sky130_hilas_poly2li  sky130_hilas_poly2li_5
timestamp 1632251374
transform -1 0 5378 0 -1 442
box 0 0 54 66
use sky130_hilas_m12m2  sky130_hilas_m12m2_9
timestamp 1632251372
transform 1 0 5768 0 1 476
box 0 0 64 64
use sky130_hilas_poly2li  sky130_hilas_poly2li_3
timestamp 1632251374
transform 1 0 5610 0 1 362
box 0 0 54 66
use sky130_hilas_nDiffThOxContact  sky130_hilas_nDiffThOxContact_0
timestamp 1632251312
transform 1 0 5192 0 1 928
box 0 0 134 58
use sky130_hilas_m12m2  sky130_hilas_m12m2_6
timestamp 1632251372
transform 1 0 5486 0 1 922
box 0 0 64 64
use sky130_hilas_m12m2  sky130_hilas_m12m2_4
timestamp 1632251372
transform 1 0 5482 0 1 750
box 0 0 64 64
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1632251372
transform 1 0 5486 0 1 834
box 0 0 64 64
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_0
timestamp 1632251409
transform 1 0 5254 0 1 814
box 0 0 66 110
use sky130_hilas_m12m2  sky130_hilas_m12m2_3
timestamp 1632251372
transform 1 0 5768 0 1 746
box 0 0 64 64
use sky130_hilas_m12m2  sky130_hilas_m12m2_2
timestamp 1632251372
transform 1 0 5768 0 1 920
box 0 0 64 64
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1632251372
transform 1 0 5768 0 1 830
box 0 0 64 64
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1632251356
transform 1 0 5634 0 1 924
box 0 0 68 66
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1632251356
transform 1 0 5634 0 1 756
box 0 0 68 66
use sky130_hilas_m12m2  sky130_hilas_m12m2_10
timestamp 1632251372
transform 1 0 5194 0 1 1136
box 0 0 64 64
use sky130_hilas_m12m2  sky130_hilas_m12m2_7
timestamp 1632251372
transform 1 0 5766 0 1 1126
box 0 0 64 64
use sky130_hilas_poly2li  sky130_hilas_poly2li_1
timestamp 1632251374
transform 1 0 5616 0 1 1138
box 0 0 54 66
use sky130_hilas_poly2li  sky130_hilas_poly2li_4
timestamp 1632251374
transform 1 0 5896 0 1 1138
box 0 0 54 66
use sky130_hilas_FGVaractorTunnelCap01  sky130_hilas_FGVaractorTunnelCap01_0
timestamp 1632251358
transform 1 0 1954 0 1 1618
box 0 0 444 338
use sky130_hilas_FGHugeVaractorCapacitor01  sky130_hilas_FGHugeVaractorCapacitor01_0
timestamp 1632251344
transform 1 0 3966 0 1 1636
box 0 0 2058 1198
use sky130_hilas_FGVaractorCapacitor02  sky130_hilas_FGVaractorCapacitor02_1
timestamp 1632251432
transform 1 0 2894 0 1 1628
box 0 0 544 338
<< labels >>
rlabel metal2 5922 92 5934 190 0 VGND
port 8 nsew ground default
rlabel metal2 5922 456 5934 520 0 OUTPUT
port 10 nsew analog default
rlabel metal2 5920 766 5934 918 0 VINJ
port 9 nsew power default
rlabel metal2 5922 378 5934 424 0 VBIAS
port 12 nsew analog default
rlabel metal2 5922 552 5934 598 0 VREF
port 11 nsew analog default
rlabel metal1 4778 4 4836 14 0 LARGECAPACITOR
port 7 nsew analog default
rlabel metal1 2114 1198 2162 1210 0 GATE3
port 3 nsew analog default
rlabel metal1 2116 0 2164 14 0 GATE4
port 6 nsew analog default
rlabel metal1 938 0 1000 14 0 GATE2
port 5 nsew analog default
rlabel metal1 940 1192 994 1210 0 GATE1
port 2 nsew analog default
rlabel metal1 156 0 208 20 0 VTUNOVERLAP01
port 4 nsew analog default
rlabel metal1 0 1196 52 1210 0 VTUN
port 1 nsew analog default
rlabel metal2 2116 832 2176 854 0 DRAIN1
port 13 nsew
rlabel metal2 2262 834 2320 856 0 SOURCE1
port 14 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
