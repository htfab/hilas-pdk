magic
tech sky130A
timestamp 1628178864
<< nwell >>
rect -1005 -215 -734 -211
rect -1005 -380 -733 -215
<< mvvaractor >>
rect -901 -322 -790 -272
<< mvnsubdiff >>
rect -972 -265 -790 -246
rect -972 -287 -950 -265
rect -901 -272 -790 -265
rect -954 -304 -950 -287
rect -972 -337 -950 -304
rect -901 -347 -790 -322
<< mvnsubdiffcont >>
rect -972 -304 -954 -287
<< poly >>
rect -941 -322 -901 -272
rect -790 -322 -749 -272
<< locali >>
rect -975 -263 -952 -259
rect -975 -280 -972 -263
rect -955 -280 -952 -263
rect -975 -287 -952 -280
rect -975 -304 -972 -287
rect -954 -304 -952 -287
rect -975 -308 -952 -304
rect -975 -325 -972 -308
rect -955 -325 -952 -308
rect -975 -328 -952 -325
<< viali >>
rect -972 -280 -955 -263
rect -972 -325 -955 -308
<< metal1 >>
rect -977 -263 -951 -254
rect -977 -280 -972 -263
rect -955 -280 -951 -263
rect -977 -308 -951 -280
rect -977 -325 -972 -308
rect -955 -325 -951 -308
rect -977 -333 -951 -325
<< end >>
