VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_m12m2
  CLASS BLOCK ;
  FOREIGN /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_m12m2 ;
  ORIGIN 0.090 0.100 ;
  SIZE 0.320 BY 0.320 ;
  OBS
      LAYER met1 ;
        RECT -0.060 -0.100 0.200 0.220 ;
      LAYER met2 ;
        RECT -0.090 -0.070 0.230 0.190 ;
  END
END /home/bjmuld/work/hilas/fastlane/PDKs/sky130A_hilas/libs.ref/sky130_hilas_sc/mag/sky130_hilas_m12m2
END LIBRARY

