magic
tech sky130A
timestamp 1627759106
<< error_s >>
rect -2550 711 -2500 722
rect -2478 711 -2428 722
rect -509 711 -459 722
rect -437 711 -387 722
rect -49 717 -22 724
rect 154 704 171 709
rect -2428 680 -2394 681
rect -543 680 -509 681
rect -2550 669 -2500 680
rect -2478 669 -2428 680
rect -509 669 -459 680
rect -437 669 -387 680
rect -49 675 -22 682
rect -49 651 -22 658
rect -2486 648 -2477 650
rect -2426 648 -2394 650
rect -2362 648 -2323 650
rect -2227 648 -2187 650
rect -750 648 -710 650
rect -614 648 -575 650
rect -543 648 -511 650
rect -460 648 -451 650
rect -2505 544 -2500 585
rect -2365 573 -2362 623
rect -2323 573 -2320 623
rect -2229 573 -2227 623
rect -2187 573 -2185 623
rect -752 573 -750 623
rect -710 573 -708 623
rect -617 573 -614 623
rect -575 573 -572 623
rect -49 609 -22 616
rect -437 561 -432 585
rect -49 569 -22 576
rect -413 544 -408 561
rect -2365 494 -2362 544
rect -2323 494 -2320 544
rect -2229 494 -2227 544
rect -2187 494 -2185 544
rect -752 494 -750 544
rect -710 494 -708 544
rect -617 494 -614 544
rect -575 494 -572 544
rect -49 527 -22 534
rect -49 503 -22 510
rect -49 461 -22 468
rect -49 421 -22 428
rect -2505 324 -2500 365
rect -2365 341 -2362 391
rect -2323 341 -2320 391
rect -2229 341 -2227 391
rect -2187 341 -2185 391
rect -752 341 -750 391
rect -710 341 -708 391
rect -617 341 -614 391
rect -575 341 -572 391
rect -49 379 -22 386
rect -437 341 -432 365
rect -49 355 -22 362
rect -413 324 -408 341
rect -49 313 -22 320
rect -2365 262 -2362 312
rect -2323 262 -2320 312
rect -2229 262 -2227 312
rect -2187 262 -2185 312
rect -752 262 -750 312
rect -710 262 -708 312
rect -617 262 -614 312
rect -575 262 -572 312
rect -49 273 -22 280
rect -2486 235 -2477 237
rect -2426 235 -2394 237
rect -2362 235 -2323 237
rect -2227 235 -2187 237
rect -750 235 -710 237
rect -614 235 -575 237
rect -543 235 -511 237
rect -460 235 -451 237
rect -49 231 -22 238
rect -2550 205 -2500 216
rect -2478 205 -2428 216
rect -509 205 -459 216
rect -437 205 -387 216
rect -49 207 -22 214
rect -2428 204 -2394 205
rect -543 204 -509 205
rect 130 201 154 206
rect -2550 163 -2500 174
rect -2478 163 -2428 174
rect -509 163 -459 174
rect -437 163 -387 174
rect -49 165 -22 172
<< nwell >>
rect -2617 744 -2286 745
rect -320 744 -186 745
rect -2597 713 -2565 743
rect -370 713 -338 743
rect 65 727 193 745
rect 65 140 193 159
<< metal1 >>
rect -2581 743 -2565 745
rect -2597 741 -2565 743
rect -2597 715 -2594 741
rect -2568 715 -2565 741
rect -2540 739 -2521 745
rect -2353 734 -2332 745
rect -2306 737 -2287 745
rect -2265 739 -2244 745
rect -2157 738 -2139 745
rect -1541 730 -1499 745
rect -1438 730 -1396 745
rect -1068 737 -1045 745
rect -416 737 -397 745
rect -372 743 -344 745
rect -372 741 -338 743
rect -372 737 -367 741
rect -1541 716 -1396 730
rect -2597 713 -2565 715
rect -370 715 -367 737
rect -341 715 -338 741
rect -3 731 31 745
rect 63 730 91 745
rect -370 713 -338 715
rect -156 188 -124 190
rect -1775 173 -1743 175
rect -2352 141 -2329 153
rect -1775 147 -1772 173
rect -1746 147 -1743 173
rect -1775 145 -1743 147
rect -1195 173 -1163 175
rect -1195 147 -1192 173
rect -1166 147 -1163 173
rect -156 162 -153 188
rect -127 162 -124 188
rect -156 160 -124 162
rect -156 159 -2 160
rect -156 154 31 159
rect -1195 145 -1163 147
rect -151 146 31 154
rect -416 140 -397 145
rect -372 140 -344 145
rect -3 140 31 146
rect 64 140 91 161
<< via1 >>
rect -2594 715 -2568 741
rect -367 715 -341 741
rect -1772 147 -1746 173
rect -1192 147 -1166 173
rect -153 162 -127 188
<< metal2 >>
rect -2597 741 -2565 743
rect -2597 715 -2594 741
rect -2568 731 -2565 741
rect -370 741 -338 743
rect -370 731 -367 741
rect -2568 715 -367 731
rect -341 715 -338 741
rect -260 718 -229 742
rect -2597 713 -338 715
rect -2617 677 -2609 695
rect -149 655 -127 657
rect -154 621 -127 655
rect -328 571 -293 593
rect -147 564 -127 565
rect -1466 522 -667 542
rect -147 531 -125 564
rect -145 530 -125 531
rect -807 454 -785 455
rect -1465 429 -782 454
rect -689 450 -667 522
rect -252 451 -220 475
rect 182 474 193 497
rect -1465 337 -1114 356
rect -1137 277 -1114 337
rect -811 312 -782 429
rect -692 446 -667 450
rect -692 382 -666 446
rect 182 392 193 414
rect -692 361 -279 382
rect -300 347 -279 361
rect -300 326 -113 347
rect -811 290 -522 312
rect -811 289 -782 290
rect -1137 262 -1115 277
rect -700 262 -113 267
rect -1137 246 -113 262
rect -1137 240 -661 246
rect -2617 190 -2609 208
rect -156 188 -124 190
rect -156 175 -153 188
rect -1775 173 -153 175
rect -1775 147 -1772 173
rect -1746 160 -1192 173
rect -1746 147 -1743 160
rect -1775 145 -1743 147
rect -1195 147 -1192 160
rect -1166 162 -153 173
rect -127 162 -124 188
rect -1166 160 -124 162
rect -1166 147 -1163 160
rect -1195 145 -1163 147
use sky130_hilas_DualTACore01  sky130_hilas_DualTACore01_0
timestamp 1627744303
transform 1 0 38 0 1 181
box -172 -22 155 550
use sky130_hilas_pTransistorPair  sky130_hilas_pTransistorPair_1
timestamp 1627744303
transform 1 0 -454 0 -1 305
box 133 -440 320 165
use sky130_hilas_FGBias2x1cell  sky130_hilas_FGBias2x1cell_0
timestamp 1627759106
transform 1 0 -1077 0 1 522
box -396 -382 757 223
use sky130_hilas_FGtrans2x1cell  sky130_hilas_FGtrans2x1cell_0
timestamp 1627744303
transform -1 0 -1860 0 1 522
box -395 -382 757 223
<< labels >>
rlabel metal1 -3 739 31 745 0 VGND
port 11 nsew
rlabel metal1 63 739 91 745 0 VPWR
port 10 nsew
rlabel metal1 64 140 91 146 0 VPWR
port 10 nsew
rlabel metal1 -3 140 31 146 0 VGND
port 11 nsew
rlabel metal2 -252 451 -220 475 0 VIN21
port 9 nsew
rlabel metal2 -260 718 -229 742 1 VIN22
port 8 n
rlabel metal1 -2352 141 -2329 153 0 VIN12
port 18 nsew
rlabel metal1 -2353 734 -2332 745 0 VIN11
port 5 nsew
rlabel metal1 -1438 738 -1396 745 0 VTUN
port 1 nsew
rlabel metal1 -1541 738 -1499 745 0 VTUN
rlabel metal1 -2265 739 -2244 745 0 PROG
port 3 nsew
rlabel metal1 -2581 739 -2565 745 0 VINJ
port 6 nsew
rlabel metal1 -372 737 -344 745 0 VINJ
port 6 nsew
rlabel metal2 182 474 193 497 0 OUTPUT1
port 13 nsew
rlabel metal2 182 392 193 414 0 OUTPUT2
port 12 nsew
rlabel metal1 -2540 739 -2521 745 0 GATESEL1
port 14 nsew
rlabel metal1 -416 140 -397 145 0 GATESEL2
port 15 nsew
rlabel metal1 -372 140 -344 145 0 VINJ
port 6 nsew
rlabel metal1 -416 737 -397 745 0 GATESEL2
port 15 nsew
rlabel metal2 -2617 677 -2609 695 0 DRAIN1
port 16 nsew
rlabel metal2 -2617 190 -2609 208 0 DRAIN2
port 17 nsew
rlabel metal1 -1068 737 -1045 745 0 GATE1
port 4 nsew
rlabel metal1 -2306 737 -2287 745 0 GATE2
port 19 nsew
rlabel metal1 -2157 738 -2139 745 0 RUN
port 20 nsew
<< end >>
