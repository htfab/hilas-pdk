magic
tech sky130A
timestamp 1627255200
<< nwell >>
rect 133 -140 319 -133
rect 267 -169 312 -146
<< poly >>
rect 225 -104 248 -100
rect 227 -407 248 -406
<< locali >>
rect 279 -70 301 -61
rect 279 -78 287 -70
rect 174 -192 192 -86
rect 247 -133 252 -120
rect 235 -146 252 -133
rect 272 -352 279 -350
rect 272 -366 280 -352
rect 249 -435 256 -409
<< metal1 >>
rect 283 -265 304 -88
<< metal2 >>
rect 225 -169 312 -146
rect 225 -170 268 -169
rect 273 -249 320 -224
rect 255 -352 310 -327
rect 201 -438 289 -413
use sky130_hilas_pTransistorVert01  sky130_hilas_pTransistorVert01_1
timestamp 1627255200
transform 1 0 496 0 1 5
box -363 -444 -177 -145
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1627255200
transform 1 0 175 0 1 -287
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1627255200
transform -1 0 275 0 -1 -421
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1627255200
transform 1 0 248 0 1 -159
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1627255200
transform -1 0 290 0 -1 -338
box -14 -15 20 18
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1627255200
transform 1 0 287 0 1 -244
box -9 -10 23 22
use sky130_hilas_poly2li  sky130_hilas_poly2li_1
timestamp 1627255200
transform 1 0 236 0 1 -426
box -9 -14 18 19
use sky130_hilas_pTransistorVert01  sky130_hilas_pTransistorVert01_0
timestamp 1627255200
transform 1 0 496 0 1 310
box -363 -444 -177 -145
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1627255200
transform 1 0 291 0 1 -85
box -10 -8 13 21
use sky130_hilas_poly2li  sky130_hilas_poly2li_0
timestamp 1627255200
transform 1 0 234 0 1 -123
box -9 -14 18 19
<< end >>
