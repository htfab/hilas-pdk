magic
tech sky130A
timestamp 1607268356
<< error_s >>
rect 78 67 101 73
rect 78 50 81 67
rect 78 44 101 50
<< psubdiff >>
rect 84 100 125 109
rect 84 83 96 100
rect 113 83 125 100
rect 84 74 125 83
rect 84 34 125 43
rect 84 17 96 34
rect 113 17 125 34
rect 84 8 125 17
<< psubdiffcont >>
rect 96 83 113 100
rect 96 17 113 34
<< poly >>
rect -46 56 53 66
rect -46 51 26 56
rect -46 43 -19 51
<< locali >>
rect 79 100 114 108
rect 79 83 96 100
rect 113 83 114 100
rect 59 75 78 76
rect 79 75 114 83
rect 59 42 114 75
rect 79 34 114 42
rect 79 17 96 34
rect 113 17 114 34
rect 79 9 114 17
<< metal2 >>
rect -59 14 -26 35
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1607179295
transform 1 0 88 0 1 52
box -10 -8 13 21
use sky130_hilas_nFET03  sky130_hilas_nFET03_0
timestamp 1607185713
transform 1 0 26 0 1 14
box -31 -19 58 42
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1607089160
transform 1 0 -15 0 1 25
box -14 -15 20 18
use sky130_hilas_poly2li  sky130_hilas_poly2li_0
timestamp 1607178257
transform 1 0 -37 0 1 24
box -9 -14 18 19
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1607089160
transform 1 0 -10 0 1 90
box -14 -15 20 18
use sky130_hilas_nFET03  sky130_hilas_nFET03_1
timestamp 1607185713
transform 1 0 26 0 1 80
box -31 -19 58 42
<< end >>
