magic
tech sky130A
timestamp 1608079637
<< error_s >>
rect -539 538 -533 544
rect -434 538 -428 544
rect 432 538 438 544
rect 537 538 543 544
rect -113 528 -107 534
rect -60 528 -54 534
rect 58 528 64 534
rect 111 528 117 534
rect -545 474 -539 480
rect -428 474 -422 480
rect -119 478 -113 484
rect -54 478 -48 484
rect 52 478 58 484
rect 117 478 123 484
rect 426 474 432 480
rect 543 474 549 480
rect -539 421 -533 427
rect -434 421 -428 427
rect -113 419 -107 425
rect -60 419 -54 425
rect 58 419 64 425
rect 111 419 117 425
rect 432 421 438 427
rect 537 421 543 427
rect -119 369 -113 375
rect -54 369 -48 375
rect 52 369 58 375
rect 117 369 123 375
rect -545 357 -539 363
rect -428 357 -422 363
rect 426 357 432 363
rect 543 357 549 363
rect -539 236 -533 242
rect -434 236 -428 242
rect 432 236 438 242
rect 537 236 543 242
rect -113 230 -107 236
rect -60 230 -54 236
rect 58 230 64 236
rect 111 230 117 236
rect -119 180 -113 186
rect -54 180 -48 186
rect 52 180 58 186
rect 117 180 123 186
rect -545 172 -539 178
rect -428 172 -422 178
rect 426 172 432 178
rect 543 172 549 178
rect -539 120 -533 126
rect -434 120 -428 126
rect 432 120 438 126
rect 537 120 543 126
rect -113 113 -107 119
rect -60 113 -54 119
rect 58 113 64 119
rect 111 113 117 119
rect -119 63 -113 69
rect -54 63 -48 69
rect 52 63 58 69
rect 117 63 123 69
rect -545 56 -539 62
rect -428 56 -422 62
rect 426 56 432 62
rect 543 56 549 62
<< metal1 >>
rect -968 596 -952 601
rect -475 591 -437 601
rect -72 588 -32 601
rect 36 591 76 601
rect 441 591 479 601
rect 875 596 891 601
rect 912 596 931 601
rect 956 596 972 601
rect -968 -4 -952 2
rect -475 -4 -437 5
rect -72 -4 -32 8
rect 36 -4 76 8
rect 441 -4 479 11
rect 956 -3 972 3
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_1
timestamp 1608069483
transform -1 0 -260 0 1 378
box -264 -382 744 223
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_0
timestamp 1608069483
transform 1 0 264 0 1 378
box -264 -382 744 223
<< labels >>
rlabel metal1 441 591 479 601 0 Gate2
port 1 nsew analog default
rlabel metal1 -72 -4 -32 8 0 Vtun
port 2 nsew power default
rlabel metal1 36 -4 76 8 0 Vtun
port 2 nsew power default
rlabel metal1 36 591 76 601 0 Vtun
port 2 nsew power default
rlabel metal1 -72 588 -32 601 0 Vtun
port 2 nsew power default
rlabel metal1 -475 591 -437 601 0 Gate1
port 3 nsew analog default
rlabel metal1 -475 -4 -437 5 0 Gate1
port 3 nsew analog default
rlabel metal1 -968 -4 -952 2 0 Vdd
port 4 nsew power default
rlabel metal1 -968 596 -952 601 0 Vdd
port 4 nsew power default
rlabel metal1 956 -3 972 3 0 Vdd
port 4 nsew power default
rlabel metal1 441 -4 479 11 0 Gate2
port 1 nsew analog default
rlabel metal1 875 596 891 601 0 Horiz2
port 5 nsew analog default
rlabel metal1 912 596 931 601 0 SelectGate2
rlabel metal1 956 596 972 601 0 Vinj
port 6 nsew power default
<< end >>
