VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO FGtrans2x1cell
  CLASS BLOCK ;
  FOREIGN FGtrans2x1cell ;
  ORIGIN 3.960 3.820 ;
  SIZE 11.530 BY 6.050 ;
  OBS
      LAYER li1 ;
        RECT 5.160 1.650 5.690 1.820 ;
        RECT 6.970 1.550 7.170 1.900 ;
        RECT 6.970 1.520 7.180 1.550 ;
        RECT 3.290 1.070 3.640 1.240 ;
        RECT 4.660 1.070 4.990 1.240 ;
        RECT -3.520 0.090 -2.970 0.520 ;
        RECT 0.110 0.280 0.340 0.970 ;
        RECT 3.290 0.280 3.640 0.450 ;
        RECT 4.660 0.280 4.990 0.450 ;
        RECT 3.300 -0.510 3.640 -0.340 ;
        RECT 4.660 -0.510 4.990 -0.340 ;
        RECT 5.410 -0.430 5.580 1.260 ;
        RECT 6.240 -0.340 6.410 1.270 ;
        RECT 6.960 0.940 7.180 1.520 ;
        RECT 6.970 0.930 7.180 0.940 ;
        RECT 6.610 0.760 6.800 0.770 ;
        RECT 6.610 0.470 6.810 0.760 ;
        RECT 6.600 0.140 6.840 0.470 ;
        RECT 6.240 -0.530 6.420 -0.340 ;
        RECT -3.520 -1.640 -2.970 -1.210 ;
        RECT 3.300 -1.250 3.640 -1.080 ;
        RECT 4.660 -1.250 4.990 -1.080 ;
        RECT 0.110 -2.660 0.340 -1.970 ;
        RECT 3.290 -2.040 3.640 -1.870 ;
        RECT 4.660 -2.040 4.990 -1.870 ;
        RECT 3.290 -2.830 3.640 -2.660 ;
        RECT 4.660 -2.830 4.990 -2.660 ;
        RECT 5.410 -2.850 5.580 -1.160 ;
        RECT 6.240 -1.250 6.420 -1.060 ;
        RECT 6.240 -2.860 6.410 -1.250 ;
        RECT 6.600 -2.060 6.840 -1.730 ;
        RECT 6.610 -2.350 6.810 -2.060 ;
        RECT 6.610 -2.360 6.800 -2.350 ;
        RECT 6.970 -2.530 7.180 -2.520 ;
        RECT 6.960 -3.110 7.180 -2.530 ;
        RECT 6.970 -3.140 7.180 -3.110 ;
        RECT 5.160 -3.410 5.690 -3.240 ;
        RECT 6.970 -3.490 7.170 -3.140 ;
      LAYER mcon ;
        RECT 6.980 1.350 7.150 1.520 ;
        RECT 0.140 0.770 0.310 0.940 ;
        RECT -3.520 0.170 -3.250 0.440 ;
        RECT 0.140 0.320 0.310 0.490 ;
        RECT 6.620 0.510 6.800 0.700 ;
        RECT -3.520 -1.560 -3.250 -1.290 ;
        RECT 0.140 -2.180 0.310 -2.010 ;
        RECT 0.140 -2.630 0.310 -2.460 ;
        RECT 6.620 -2.290 6.800 -2.100 ;
        RECT 6.980 -3.110 7.150 -2.940 ;
      LAYER met1 ;
        RECT -3.610 -3.820 -3.190 2.230 ;
        RECT 5.090 1.550 5.390 1.930 ;
        RECT 0.090 0.230 0.350 1.020 ;
        RECT 6.610 0.770 6.800 2.230 ;
        RECT 7.050 1.580 7.210 2.230 ;
        RECT 6.940 1.030 7.210 1.580 ;
        RECT 6.940 0.980 7.220 1.030 ;
        RECT 7.050 0.890 7.220 0.980 ;
        RECT 6.610 0.740 6.830 0.770 ;
        RECT 6.590 0.470 6.840 0.740 ;
        RECT 6.600 0.460 6.840 0.470 ;
        RECT 6.600 0.220 6.830 0.460 ;
        RECT 6.210 -0.590 6.450 -0.210 ;
        RECT 6.210 -1.380 6.450 -1.000 ;
        RECT 6.640 -1.810 6.800 0.220 ;
        RECT 0.090 -2.710 0.350 -1.920 ;
        RECT 6.600 -2.050 6.830 -1.810 ;
        RECT 6.600 -2.060 6.840 -2.050 ;
        RECT 6.590 -2.330 6.840 -2.060 ;
        RECT 6.610 -2.360 6.830 -2.330 ;
        RECT 5.090 -3.520 5.390 -3.140 ;
        RECT 6.610 -3.820 6.800 -2.360 ;
        RECT 7.050 -2.480 7.210 0.890 ;
        RECT 7.050 -2.570 7.220 -2.480 ;
        RECT 6.940 -2.620 7.220 -2.570 ;
        RECT 6.940 -3.170 7.210 -2.620 ;
        RECT 7.050 -3.820 7.210 -3.170 ;
      LAYER via ;
        RECT 5.110 1.610 5.370 1.880 ;
        RECT 5.110 -3.470 5.370 -3.200 ;
      LAYER met2 ;
        RECT 5.090 1.750 5.390 1.930 ;
        RECT 4.840 1.730 5.390 1.750 ;
        RECT -3.960 1.550 7.570 1.730 ;
        RECT 5.100 -3.140 5.140 -3.130 ;
        RECT 5.010 -3.150 7.570 -3.140 ;
        RECT -3.940 -3.300 7.570 -3.150 ;
        RECT 5.010 -3.320 7.570 -3.300 ;
        RECT 5.090 -3.520 5.390 -3.320 ;
  END
END FGtrans2x1cell
END LIBRARY

