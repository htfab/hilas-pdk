magic
tech sky130A
timestamp 1632256337
<< error_p >>
rect 0 575 7 641
rect 57 575 116 606
rect 0 566 116 575
rect 0 557 149 566
rect 24 489 149 557
rect 398 483 410 572
rect 57 246 116 278
rect 24 161 149 246
rect 398 159 410 252
<< error_s >>
rect 1481 1023 1499 1051
rect 1508 1023 1526 1053
rect 1508 1017 1540 1023
rect 1508 967 1529 1017
rect 1508 959 1540 967
rect 1481 938 1499 959
rect 1388 934 1499 938
rect 1508 949 1526 959
rect 1508 933 1567 949
rect 1388 907 1499 911
rect 1481 886 1499 907
rect 1508 906 1567 922
rect 1508 886 1526 906
rect 1466 883 1499 886
rect 1107 698 1157 704
rect 1179 698 1229 704
rect 874 664 890 678
rect 911 663 930 677
rect 955 663 971 677
rect 1078 662 1108 664
rect 1078 658 1157 662
rect 1107 656 1157 658
rect 1179 656 1229 662
rect 1064 646 1094 650
rect 1066 644 1094 646
rect 431 572 542 600
rect 410 483 575 572
rect 1040 541 1296 641
rect 1332 614 1423 859
rect 1508 848 1529 883
rect 1502 844 1540 848
rect 1492 819 1499 844
rect 1475 794 1499 819
rect 1502 836 1567 844
rect 1502 819 1540 836
rect 1502 774 1526 819
rect 1481 698 1499 726
rect 1508 698 1526 733
rect 1508 697 1540 698
rect 1508 647 1529 697
rect 1508 634 1540 647
rect 1481 614 1499 634
rect 1332 609 1499 614
rect 1508 621 1526 634
rect 1508 613 1567 621
rect 1332 587 1423 609
rect 1332 582 1499 587
rect 828 374 1013 457
rect 828 373 912 374
rect 930 373 1013 374
rect 887 369 1013 373
rect 887 366 900 369
rect 895 362 900 366
rect 907 362 1013 369
rect 895 357 1013 362
rect 1040 357 1057 501
rect 1107 462 1157 468
rect 1332 436 1423 582
rect 1481 559 1499 582
rect 1508 586 1567 594
rect 1508 559 1526 586
rect 1508 558 1540 559
rect 1508 508 1529 558
rect 1508 495 1540 508
rect 1481 470 1499 495
rect 1508 474 1526 495
rect 1107 420 1157 426
rect 1066 409 1094 411
rect 1064 405 1094 409
rect 1078 391 1108 397
rect 1066 378 1092 380
rect 1066 370 1108 378
rect 1236 370 1256 378
rect 904 352 917 357
rect 904 349 912 352
rect 930 350 933 354
rect 1066 351 1092 370
rect 1097 353 1108 361
rect 1078 334 1108 340
rect 1064 322 1094 326
rect 1066 320 1094 322
rect 431 252 542 276
rect 410 159 575 252
rect 1040 217 1296 318
rect 1107 139 1157 145
rect 1040 99 1054 117
rect 1107 97 1157 103
rect 1066 86 1094 88
rect 1064 82 1094 86
rect 1107 74 1157 76
rect 1078 70 1157 74
rect 1179 70 1229 76
rect 1078 68 1108 70
rect 1107 28 1157 34
rect 1179 28 1229 34
<< nwell >>
rect 0 557 7 575
rect 57 522 116 533
rect 431 516 542 539
rect 895 373 930 374
rect 895 357 912 373
rect 929 357 930 373
rect 57 194 116 213
rect 431 192 542 219
<< psubdiff >>
rect 278 527 304 550
rect 278 510 282 527
rect 299 510 304 527
rect 670 526 697 552
rect 278 484 304 510
rect 670 509 676 526
rect 693 509 697 526
rect 670 486 697 509
rect 279 415 304 442
rect 279 398 283 415
rect 300 398 304 415
rect 279 381 304 398
rect 279 364 283 381
rect 300 364 304 381
rect 279 347 304 364
rect 279 330 283 347
rect 300 330 304 347
rect 279 302 304 330
rect 672 401 697 428
rect 672 384 676 401
rect 693 384 697 401
rect 672 367 697 384
rect 672 350 676 367
rect 693 350 697 367
rect 672 333 697 350
rect 672 316 676 333
rect 693 316 697 333
rect 672 303 697 316
<< mvnsubdiff >>
rect 57 522 116 533
rect 431 516 542 539
rect 57 194 116 213
rect 431 192 542 219
<< psubdiffcont >>
rect 282 510 299 527
rect 676 509 693 526
rect 283 398 300 415
rect 283 364 300 381
rect 283 330 300 347
rect 676 384 693 401
rect 676 350 693 367
rect 676 316 693 333
<< poly >>
rect 583 596 751 613
rect 156 559 393 583
rect 156 450 391 474
rect 582 442 751 459
rect 912 373 930 374
rect 928 357 930 373
rect 156 270 393 294
rect 640 289 660 295
rect 583 272 751 289
rect 158 120 391 144
rect 583 120 752 136
<< polycont >>
rect 895 357 912 374
<< locali >>
rect 282 527 299 529
rect 676 526 693 528
rect 283 415 300 423
rect 283 381 300 383
rect 283 322 300 330
rect 676 401 693 409
rect 676 367 693 369
rect 886 357 895 374
rect 676 308 693 316
<< viali >>
rect 282 529 299 546
rect 282 493 299 510
rect 676 528 693 545
rect 676 492 693 509
rect 283 398 300 400
rect 283 383 300 398
rect 283 347 300 364
rect 676 384 693 386
rect 676 369 693 384
rect 912 357 930 374
rect 676 333 693 350
<< metal1 >>
rect 35 41 75 691
rect 279 550 303 691
rect 440 658 478 691
rect 672 552 696 691
rect 874 664 890 668
rect 911 663 930 668
rect 955 663 971 668
rect 278 546 304 550
rect 278 529 282 546
rect 299 529 304 546
rect 278 510 304 529
rect 278 493 282 510
rect 299 493 304 510
rect 278 484 304 493
rect 670 545 697 552
rect 670 528 676 545
rect 693 528 697 545
rect 670 509 697 528
rect 670 492 676 509
rect 693 492 697 509
rect 670 486 697 492
rect 279 400 303 484
rect 279 383 283 400
rect 300 383 303 400
rect 279 364 303 383
rect 279 347 283 364
rect 300 347 303 364
rect 279 223 303 347
rect 672 386 696 486
rect 672 369 676 386
rect 693 369 696 386
rect 917 377 930 379
rect 909 375 933 377
rect 672 350 696 369
rect 889 374 933 375
rect 889 357 912 374
rect 930 357 933 374
rect 889 356 933 357
rect 909 354 933 356
rect 919 350 930 354
rect 672 333 676 350
rect 693 333 696 350
rect 672 227 696 333
rect 671 224 697 227
rect 278 220 304 223
rect 671 195 697 198
rect 278 191 304 194
rect 279 41 303 191
rect 440 41 478 101
rect 672 41 696 195
<< via1 >>
rect 278 194 304 220
rect 671 198 697 224
<< metal2 >>
rect 0 617 763 635
rect 0 573 763 591
rect 0 463 763 481
rect 0 420 763 438
rect 0 293 762 311
rect 0 250 763 268
rect 668 224 700 225
rect 275 194 278 220
rect 304 219 307 220
rect 668 219 671 224
rect 304 201 671 219
rect 304 194 307 201
rect 668 198 671 201
rect 697 198 700 224
rect 668 196 700 198
rect 0 140 762 158
rect 0 98 760 115
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_1
timestamp 1632255311
transform 1 0 1040 0 1 0
box 0 0 256 191
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_2
timestamp 1632255311
transform 1 0 1040 0 -1 408
box 0 0 256 191
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_3
timestamp 1632255311
transform 1 0 1040 0 -1 732
box 0 0 256 191
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_0
timestamp 1632255311
transform 1 0 1040 0 1 323
box 0 0 256 191
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_0
timestamp 1632251397
transform 1 0 1332 0 1 436
box 0 0 223 186
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_1
timestamp 1632251302
transform 1 0 1451 0 1 441
box 0 0 173 190
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_1
timestamp 1632251397
transform 1 0 1332 0 1 575
box 0 0 223 186
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_2
timestamp 1632251397
transform 1 0 1332 0 1 760
box 0 0 223 186
use sky130_hilas_wellContact  sky130_hilas_wellContact_1
timestamp 1632251355
transform 1 0 1448 0 1 738
box 0 0 173 186
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_2
timestamp 1632251302
transform 1 0 1451 0 1 769
box 0 0 173 190
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_0
timestamp 1632251302
transform 1 0 1451 0 1 580
box 0 0 173 190
use sky130_hilas_wellContact  sky130_hilas_wellContact_0
timestamp 1632251355
transform 1 0 1851 0 1 731
box 0 0 173 186
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_3
timestamp 1632251397
transform 1 0 1332 0 1 900
box 0 0 223 186
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_3
timestamp 1632251302
transform 1 0 1451 0 1 900
box 0 0 173 190
<< labels >>
rlabel metal1 35 656 75 668 0 VTUN
port 1 nsew
rlabel metal1 955 663 971 668 0 VINJ
port 2 nsew
rlabel metal1 911 663 930 668 0 COLSEL1
port 3 nsew
rlabel metal1 874 664 890 668 0 COL1
port 4 nsew
rlabel metal1 440 658 478 668 0 GATE1
port 5 nsew
rlabel poly 642 279 659 294 0 FG3
rlabel metal1 279 663 303 668 0 VGND
port 14 nsew
rlabel metal1 672 663 696 668 0 VGND
port 14 nsew
rlabel metal1 672 63 696 69 0 VGND
port 14 nsew
rlabel metal1 279 63 303 69 0 VGND
port 14 nsew
rlabel metal1 440 63 478 72 0 GATE1
port 5 nsew
rlabel metal2 0 98 8 115 0 DRAIN4
port 15 nsew
rlabel metal2 0 140 6 158 0 ROW4
port 11 nsew
rlabel metal2 0 617 6 635 0 DRAIN1
port 16 nsew
rlabel metal2 0 573 6 591 0 ROW1
port 17 nsew
rlabel metal2 0 250 6 268 0 ROW3
port 18 nsew
rlabel metal2 0 293 6 311 0 DRAIN3
port 19 nsew
rlabel metal2 0 420 6 438 0 DRAIN2
port 20 nsew
rlabel metal2 0 463 6 481 0 ROW2
port 21 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
