magic
tech sky130A
timestamp 1632251410
<< checkpaint >>
rect -41 952 1939 1417
rect -592 -383 1939 952
rect -41 -426 1939 -383
<< metal2 >>
rect 0 485 1042 503
rect 0 442 1042 460
rect 3 342 1042 360
rect 851 317 1042 318
rect 3 299 1042 317
rect 2 237 29 265
rect 1006 238 1042 266
rect 3 184 1042 201
rect 3 142 1042 159
rect 3 44 1042 61
rect 3 0 1042 17
<< metal3 >>
rect 823 212 1019 287
<< metal4 >>
rect 116 277 217 278
rect 45 227 380 277
rect 45 226 152 227
rect 316 115 379 227
rect 316 85 531 115
rect 349 84 531 85
use sky130_hilas_CapModule02  sky130_hilas_CapModule02_0
timestamp 1632251385
transform 1 0 589 0 1 204
box 0 0 720 583
use sky130_hilas_m22m4  sky130_hilas_m22m4_0
timestamp 1632251386
transform 1 0 38 0 1 247
box 0 0 79 75
use sky130_hilas_m22m4  sky130_hilas_m22m4_1
timestamp 1632251386
transform 1 0 987 0 1 248
box 0 0 79 75
<< labels >>
rlabel metal2 2 237 9 265 0 CAPTERM01
port 2 nsew analog default
rlabel metal2 1030 238 1042 266 0 CAPTERM02
port 1 nsew analog default
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
