magic
tech sky130A
timestamp 1632492731
<< metal1 >>
rect -887 596 -871 601
rect -693 592 -669 601
rect -475 591 -437 601
rect -300 595 -276 601
rect -72 588 -32 601
rect 36 591 76 601
rect 280 596 304 601
rect 441 591 479 601
rect 673 594 697 601
rect 875 596 891 601
rect -32 565 36 587
rect -887 -3 -871 3
rect -693 -4 -669 4
rect -475 -4 -437 5
rect -300 -4 -276 3
rect -72 -4 -32 8
rect 36 -4 76 8
rect 280 -4 304 3
rect 441 -4 479 11
rect 673 -4 697 2
rect 875 -3 891 3
<< metal2 >>
rect -1004 507 -997 525
rect 999 507 1008 525
rect -1004 396 -998 414
rect 1002 396 1008 414
rect -1004 183 -997 201
rect 999 183 1008 201
rect -334 134 342 152
rect -1004 73 -997 91
rect 999 73 1008 91
use sky130_hilas_cellAttempt01d3  sky130_hilas_cellAttempt01d3_1
timestamp 1632492731
transform -1 0 -260 0 1 378
box -263 -404 744 246
use sky130_hilas_cellAttempt01d3  sky130_hilas_cellAttempt01d3_0
timestamp 1632492731
transform 1 0 264 0 1 378
box -263 -404 744 246
<< labels >>
rlabel metal1 441 591 479 601 0 GATE2
port 1 nsew analog default
rlabel metal1 -72 -4 -32 8 0 VTUN
port 2 nsew power default
rlabel metal1 36 -4 76 8 0 VTUN
port 2 nsew power default
rlabel metal1 36 591 76 601 0 VTUN
port 2 nsew power default
rlabel metal1 -72 588 -32 601 0 VTUN
port 2 nsew power default
rlabel metal1 -475 591 -437 601 0 GATE1
port 3 nsew analog default
rlabel metal1 -475 -4 -437 5 0 GATE1
port 3 nsew analog default
rlabel metal1 441 -4 479 11 0 GATE2
port 1 nsew analog default
rlabel metal1 -887 596 -871 601 0 COL1
port 12 nsew analog default
rlabel metal1 -887 -3 -871 3 0 COL1
port 12 nsew analog default
rlabel metal1 875 -3 891 3 0 COL2
port 13 nsew analog default
rlabel metal1 875 596 891 601 0 COL2
port 13 nsew analog default
rlabel metal1 -693 595 -669 601 0 VGND
port 22 nsew
rlabel metal1 -693 -4 -669 4 0 VGND
port 22 nsew
rlabel metal1 -300 -4 -276 3 0 VGND
port 22 nsew
rlabel metal1 -300 595 -276 601 0 VGND
port 22 nsew
rlabel metal1 280 -4 304 3 0 VGND
port 22 nsew
rlabel metal1 673 -4 697 2 0 VGND
port 22 nsew
rlabel metal1 280 596 304 601 0 VGND
port 22 nsew
rlabel metal1 673 594 697 601 0 VGND
port 22 nsew
rlabel metal2 -1004 73 -997 91 0 ROW4
port 20 nsew
rlabel metal2 -1004 183 -997 201 0 ROW3
port 19 nsew
rlabel metal2 -1004 396 -998 414 0 ROW2
port 15 nsew
rlabel metal2 -1004 507 -997 525 0 ROW1
port 14 nsew
rlabel metal2 999 507 1008 525 0 ROW1
port 14 nsew
rlabel metal2 1002 396 1008 414 0 ROW2
port 15 nsew
rlabel metal2 999 183 1008 201 0 ROW3
port 19 nsew
rlabel metal2 999 73 1008 91 0 ROW4
port 20 nsew
<< end >>
