magic
tech sky130A
timestamp 1627744303
<< error_s >>
rect 9 -126 49 -115
rect 9 -168 49 -157
<< nwell >>
rect -18 -97 96 -38
rect -67 -181 96 -97
<< pmos >>
rect 9 -157 49 -126
<< pdiff >>
rect -20 -133 9 -126
rect -20 -150 -14 -133
rect 3 -150 9 -133
rect -20 -157 9 -150
rect 49 -133 78 -126
rect 49 -150 55 -133
rect 72 -150 78 -133
rect 49 -157 78 -150
<< pdiffc >>
rect -14 -150 3 -133
rect 55 -150 72 -133
<< poly >>
rect -18 -56 96 -40
rect 9 -126 49 -103
rect 9 -170 49 -157
<< locali >>
rect -18 -88 96 -70
rect -14 -133 3 -125
rect 47 -150 55 -133
rect 72 -150 85 -132
rect -14 -155 3 -150
<< metal1 >>
rect 74 -126 93 -67
rect 72 -155 95 -126
<< metal2 >>
rect 59 -72 96 -52
rect -67 -150 -45 -149
rect -67 -170 96 -150
rect -67 -171 -45 -170
use sky130_hilas_li2m1  sky130_hilas_li2m1_3
timestamp 1627744303
transform 1 0 82 0 1 -147
box -10 -8 13 21
use sky130_hilas_m12m2  sky130_hilas_m12m2_2
timestamp 1627744303
transform 1 0 73 0 1 -69
box -9 -10 23 22
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1627744303
transform 1 0 -14 0 1 -155
box -14 -15 20 18
<< end >>
