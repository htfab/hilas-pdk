magic
tech sky130A
timestamp 1634057761
<< nwell >>
rect 1487 191 2692 785
<< mvndiff >>
rect 187 772 1344 777
rect 187 755 193 772
rect 1338 755 1344 772
rect 187 746 1344 755
rect 187 715 218 746
rect 187 708 1344 715
rect 187 691 193 708
rect 1338 691 1344 708
rect 187 684 1344 691
rect 187 653 218 684
rect 187 646 1344 653
rect 187 629 193 646
rect 1337 629 1344 646
rect 187 623 1344 629
rect 187 593 218 623
rect 187 586 1344 593
rect 187 569 193 586
rect 1338 569 1344 586
rect 187 563 1344 569
rect 187 533 218 563
rect 187 527 1344 533
rect 187 510 193 527
rect 1338 510 1344 527
rect 187 504 1344 510
rect 187 474 218 504
rect 187 468 1344 474
rect 187 451 193 468
rect 1338 451 1344 468
rect 187 445 1344 451
rect 187 415 218 445
rect 187 409 1344 415
rect 187 392 193 409
rect 1337 392 1344 409
rect 187 385 1344 392
rect 187 354 218 385
rect 1313 384 1344 385
rect 187 348 1344 354
rect 187 331 193 348
rect 1338 331 1344 348
rect 187 324 1344 331
rect 187 293 218 324
rect 187 286 1344 293
rect 187 269 194 286
rect 1338 269 1344 286
rect 187 263 1344 269
rect 187 233 218 263
rect 186 225 1344 233
rect 186 208 193 225
rect 1337 208 1344 225
rect 186 203 1344 208
<< mvpdiff >>
rect 1579 692 2595 697
rect 1579 675 1592 692
rect 2564 675 2595 692
rect 1579 668 2595 675
rect 2564 633 2595 668
rect 1581 625 2595 633
rect 1581 608 1589 625
rect 2558 608 2595 625
rect 1581 601 2595 608
rect 2564 559 2595 601
rect 1586 552 2595 559
rect 1586 535 1594 552
rect 2569 535 2595 552
rect 1586 527 2595 535
rect 2564 490 2595 527
rect 1586 484 2595 490
rect 1586 467 1593 484
rect 2561 467 2595 484
rect 1586 458 2595 467
rect 2564 425 2595 458
rect 1582 417 2595 425
rect 1582 400 1589 417
rect 2563 400 2595 417
rect 1582 392 2595 400
rect 2564 361 2595 392
rect 1582 353 2595 361
rect 1582 336 1588 353
rect 2561 336 2595 353
rect 1582 328 2595 336
rect 2564 298 2595 328
rect 1582 291 2595 298
rect 1582 274 1590 291
rect 2561 274 2595 291
rect 1582 267 2595 274
<< mvndiffc >>
rect 193 755 1338 772
rect 193 691 1338 708
rect 193 629 1337 646
rect 193 569 1338 586
rect 193 510 1338 527
rect 193 451 1338 468
rect 193 392 1337 409
rect 193 331 1338 348
rect 194 269 1338 286
rect 193 208 1337 225
<< mvpdiffc >>
rect 1592 675 2564 692
rect 1589 608 2558 625
rect 1594 535 2569 552
rect 1593 467 2561 484
rect 1589 400 2563 417
rect 1588 336 2561 353
rect 1590 274 2561 291
<< psubdiff >>
rect 47 877 81 878
rect 47 875 99 877
rect 1447 875 2799 877
rect 47 869 2799 875
rect 47 852 124 869
rect 2711 852 2799 869
rect 47 835 2799 852
rect 47 818 124 835
rect 2711 818 2799 835
rect 47 812 2799 818
rect 47 174 55 812
rect 72 799 114 812
rect 72 190 89 799
rect 106 190 114 799
rect 1391 808 2801 812
rect 1391 799 1454 808
rect 72 174 114 190
rect 47 173 114 174
rect 1391 185 1396 799
rect 1413 797 1454 799
rect 1413 185 1430 797
rect 1391 184 1430 185
rect 1447 184 1454 797
rect 2733 806 2801 808
rect 1391 177 1454 184
rect 2733 184 2738 806
rect 2755 802 2801 806
rect 2755 184 2776 802
rect 2733 183 2776 184
rect 2793 183 2801 802
rect 2733 177 2801 183
rect 1391 173 2801 177
rect 47 167 2801 173
rect 47 150 121 167
rect 2722 150 2801 167
rect 47 133 2801 150
rect 47 122 121 133
rect 48 116 121 122
rect 2722 116 2801 133
rect 48 110 2801 116
rect 48 106 114 110
rect 1280 108 2801 110
rect 48 105 99 106
<< nsubdiff >>
rect 1518 746 2654 752
rect 1518 729 1547 746
rect 2614 729 2654 746
rect 1518 724 2654 729
rect 1518 711 1546 724
rect 1518 252 1523 711
rect 1540 252 1546 711
rect 2626 721 2654 724
rect 1518 240 1546 252
rect 2626 252 2631 721
rect 2648 252 2654 721
rect 2626 240 2654 252
rect 1512 235 2654 240
rect 1512 218 1553 235
rect 2620 218 2654 235
rect 1512 212 2654 218
<< psubdiffcont >>
rect 124 852 2711 869
rect 124 818 2711 835
rect 55 174 72 812
rect 89 190 106 799
rect 1396 185 1413 799
rect 1430 184 1447 797
rect 2738 184 2755 806
rect 2776 183 2793 802
rect 121 150 2722 167
rect 121 116 2722 133
<< nsubdiffcont >>
rect 1547 729 2614 746
rect 1523 252 1540 711
rect 2631 252 2648 721
rect 1553 218 2620 235
<< poly >>
rect 777 1025 794 1036
rect 1445 1025 1462 1036
rect 768 1019 818 1025
rect 768 1002 777 1019
rect 794 1002 818 1019
rect 768 985 818 1002
rect 768 968 777 985
rect 794 968 818 985
rect 768 951 818 968
rect 768 934 777 951
rect 794 934 818 951
rect 768 917 818 934
rect 1399 1017 1471 1025
rect 1399 1000 1445 1017
rect 1462 1000 1471 1017
rect 1399 983 1471 1000
rect 1399 966 1445 983
rect 1462 966 1471 983
rect 1399 949 1471 966
rect 1399 932 1445 949
rect 1462 932 1471 949
rect 768 900 777 917
rect 794 900 818 917
rect 768 893 818 900
rect 1399 893 1471 932
<< polycont >>
rect 777 1002 794 1019
rect 777 968 794 985
rect 777 934 794 951
rect 1445 1000 1462 1017
rect 1445 966 1462 983
rect 1445 932 1462 949
rect 777 900 794 917
<< npolyres >>
rect 818 923 1399 1025
<< locali >>
rect 773 1019 798 1039
rect 773 987 777 1019
rect 794 987 798 1019
rect 773 985 798 987
rect 773 934 777 985
rect 794 934 798 985
rect 773 931 798 934
rect 773 900 777 931
rect 794 900 798 931
rect 773 893 798 900
rect 1441 1036 1466 1038
rect 1441 1019 1445 1036
rect 1462 1019 1466 1036
rect 1441 1017 1466 1019
rect 1441 966 1445 1017
rect 1462 966 1466 1017
rect 1441 964 1466 966
rect 1441 932 1445 964
rect 1462 932 1466 964
rect 1441 928 1466 932
rect 1441 911 1445 928
rect 1462 911 1466 928
rect 777 892 794 893
rect 1441 890 1466 911
rect 55 853 124 869
rect 55 835 63 853
rect 2711 852 2793 869
rect 250 835 2399 852
rect 55 818 124 835
rect 2715 834 2793 852
rect 2711 829 2793 834
rect 2711 818 2756 829
rect 55 816 135 818
rect 55 812 67 816
rect 85 799 107 816
rect 85 626 89 799
rect 72 190 89 626
rect 106 625 107 799
rect 125 625 135 816
rect 1396 799 1447 818
rect 193 773 210 781
rect 1317 773 1340 782
rect 193 772 1340 773
rect 192 755 193 772
rect 1338 755 1340 772
rect 192 739 1340 755
rect 192 722 226 739
rect 1324 722 1340 739
rect 192 708 1340 722
rect 192 691 193 708
rect 1338 691 1340 708
rect 192 677 1340 691
rect 192 660 226 677
rect 1324 660 1340 677
rect 192 646 1340 660
rect 192 629 193 646
rect 1337 629 1340 646
rect 192 615 1340 629
rect 192 598 227 615
rect 1325 598 1340 615
rect 192 586 1340 598
rect 192 569 193 586
rect 1338 569 1340 586
rect 192 557 1340 569
rect 192 540 229 557
rect 1327 540 1340 557
rect 192 527 1340 540
rect 192 510 193 527
rect 1338 510 1340 527
rect 192 498 1340 510
rect 192 481 230 498
rect 1328 481 1340 498
rect 192 468 1340 481
rect 192 451 193 468
rect 1338 451 1340 468
rect 192 438 1340 451
rect 192 421 230 438
rect 1328 421 1340 438
rect 192 409 1340 421
rect 192 392 193 409
rect 1337 392 1340 409
rect 192 378 1340 392
rect 192 361 225 378
rect 1323 361 1340 378
rect 192 348 1340 361
rect 192 331 193 348
rect 1338 331 1340 348
rect 192 317 1340 331
rect 192 300 226 317
rect 1324 300 1340 317
rect 192 286 1340 300
rect 192 269 194 286
rect 1338 269 1340 286
rect 192 257 1340 269
rect 192 240 225 257
rect 1323 240 1340 257
rect 192 225 1340 240
rect 185 208 193 225
rect 1337 208 1340 225
rect 192 202 211 208
rect 72 174 106 190
rect 1317 184 1340 208
rect 1413 797 1447 799
rect 1413 185 1430 797
rect 1396 184 1430 185
rect 2738 806 2756 818
rect 1523 729 1547 746
rect 2614 729 2648 746
rect 1523 711 1540 729
rect 2631 721 2648 729
rect 1579 696 2590 697
rect 1579 692 2592 696
rect 1579 675 1592 692
rect 2564 675 2592 692
rect 1579 663 2592 675
rect 1579 646 1599 663
rect 2544 646 2592 663
rect 1579 625 2592 646
rect 1579 608 1589 625
rect 2558 608 2592 625
rect 1579 588 2592 608
rect 1579 571 1598 588
rect 2537 571 2592 588
rect 1579 552 2592 571
rect 1579 535 1594 552
rect 2569 535 2592 552
rect 1579 516 2592 535
rect 1579 499 1601 516
rect 2541 499 2592 516
rect 1579 484 2592 499
rect 1579 467 1593 484
rect 2561 467 2592 484
rect 1579 450 2592 467
rect 1579 433 1602 450
rect 2539 433 2592 450
rect 1579 417 2592 433
rect 1579 400 1589 417
rect 2563 400 2592 417
rect 1579 385 2592 400
rect 1579 368 1601 385
rect 2546 368 2592 385
rect 1579 353 2592 368
rect 1579 336 1588 353
rect 2561 336 2592 353
rect 1579 321 2592 336
rect 1579 304 1602 321
rect 2541 304 2592 321
rect 1579 291 2592 304
rect 1579 274 1590 291
rect 2561 274 2592 291
rect 1579 273 2592 274
rect 1579 265 2590 273
rect 1523 242 1540 252
rect 1522 235 1540 242
rect 2648 542 2692 553
rect 2648 252 2649 542
rect 2631 235 2649 252
rect 1522 218 1553 235
rect 2620 218 2649 235
rect 2638 212 2649 218
rect 2684 212 2692 542
rect 2638 207 2692 212
rect 55 167 106 174
rect 180 167 360 168
rect 1396 167 1447 184
rect 2755 736 2756 806
rect 2776 802 2793 829
rect 2755 184 2776 736
rect 2738 183 2776 184
rect 2737 167 2793 183
rect 55 150 121 167
rect 2722 150 2793 167
rect 55 133 2793 150
rect 58 116 121 133
rect 2722 116 2793 133
rect 58 114 127 116
rect 178 115 358 116
<< viali >>
rect 777 1002 794 1004
rect 777 987 794 1002
rect 777 951 794 968
rect 777 917 794 931
rect 777 914 794 917
rect 1445 1019 1462 1036
rect 1445 983 1462 1000
rect 1445 949 1462 964
rect 1445 947 1462 949
rect 1445 911 1462 928
rect 63 852 124 853
rect 124 852 249 853
rect 63 835 250 852
rect 2399 835 2715 852
rect 2399 834 2711 835
rect 2711 834 2715 835
rect 67 812 85 816
rect 67 626 72 812
rect 72 626 85 812
rect 107 625 125 816
rect 226 722 1324 739
rect 226 660 1324 677
rect 227 598 1325 615
rect 229 540 1327 557
rect 230 481 1328 498
rect 230 421 1328 438
rect 225 361 1323 378
rect 226 300 1324 317
rect 225 240 1323 257
rect 1599 646 2544 663
rect 1598 571 2537 588
rect 1601 499 2541 516
rect 1602 433 2539 450
rect 1601 368 2546 385
rect 1602 304 2541 321
rect 2649 212 2684 542
rect 2756 736 2776 829
<< metal1 >>
rect 771 1028 1161 1087
rect 1435 1036 1470 1041
rect 771 1004 800 1028
rect 1435 1025 1445 1036
rect 771 987 777 1004
rect 794 987 800 1004
rect 771 968 800 987
rect 771 951 777 968
rect 794 951 800 968
rect 771 931 800 951
rect 771 914 777 931
rect 794 914 800 931
rect 1434 1019 1445 1025
rect 1462 1025 1470 1036
rect 1462 1019 1471 1025
rect 1434 1000 1471 1019
rect 1434 983 1445 1000
rect 1462 983 1471 1000
rect 1434 964 1471 983
rect 1434 947 1445 964
rect 1462 947 1471 964
rect 1434 930 1471 947
rect 771 893 800 914
rect 1399 928 1646 930
rect 1399 911 1445 928
rect 1462 911 1646 928
rect 1399 893 1646 911
rect 44 861 281 876
rect 44 853 66 861
rect 44 835 63 853
rect 44 828 66 835
rect 269 828 281 861
rect 44 816 281 828
rect 44 813 67 816
rect 47 804 67 813
rect 85 804 107 816
rect 125 813 281 816
rect 125 804 142 813
rect 217 811 275 813
rect 47 742 60 804
rect 130 742 142 804
rect 1255 747 1646 893
rect 2378 863 2791 868
rect 2378 852 2405 863
rect 2704 852 2791 863
rect 2378 834 2399 852
rect 2715 834 2791 852
rect 2378 828 2405 834
rect 2704 829 2791 834
rect 2704 828 2756 829
rect 2378 824 2756 828
rect 2776 828 2791 829
rect 2776 824 2792 828
rect 2378 819 2748 824
rect 284 746 1646 747
rect 47 626 67 742
rect 85 626 107 742
rect 47 625 107 626
rect 125 625 142 742
rect 47 617 142 625
rect 70 50 142 617
rect 217 739 1646 746
rect 217 722 226 739
rect 1324 722 1646 739
rect 2739 748 2748 819
rect 2783 748 2792 824
rect 2739 736 2756 748
rect 2776 736 2792 748
rect 2739 729 2792 736
rect 217 690 1646 722
rect 217 677 2552 690
rect 217 660 226 677
rect 1324 663 2552 677
rect 1324 660 1599 663
rect 217 646 1599 660
rect 2544 646 2552 663
rect 217 615 2552 646
rect 217 598 227 615
rect 1325 598 2552 615
rect 217 588 2552 598
rect 217 571 1598 588
rect 2537 571 2552 588
rect 217 557 2552 571
rect 217 540 229 557
rect 1327 540 2552 557
rect 217 516 2552 540
rect 217 499 1601 516
rect 2541 499 2552 516
rect 217 498 2552 499
rect 217 481 230 498
rect 1328 481 2552 498
rect 217 450 2552 481
rect 217 438 1602 450
rect 217 421 230 438
rect 1328 433 1602 438
rect 2539 433 2552 450
rect 1328 421 2552 433
rect 217 385 2552 421
rect 217 378 1601 385
rect 217 361 225 378
rect 1323 368 1601 378
rect 2546 368 2552 385
rect 1323 361 2552 368
rect 217 321 2552 361
rect 217 317 1602 321
rect 217 300 226 317
rect 1324 304 1602 317
rect 2541 304 2552 321
rect 1324 300 2552 304
rect 217 260 2552 300
rect 2629 548 2686 549
rect 2629 542 2691 548
rect 2629 536 2649 542
rect 2684 536 2691 542
rect 217 257 1646 260
rect 217 240 225 257
rect 1323 240 1646 257
rect 217 232 1646 240
rect 1255 77 1646 232
rect 2629 219 2645 536
rect 2687 219 2691 536
rect 2629 212 2649 219
rect 2684 212 2691 219
rect 2629 206 2691 212
rect 2629 205 2686 206
rect 2546 89 2602 92
rect 1253 0 1648 77
rect 2546 42 2548 89
rect 2547 37 2548 42
rect 2600 37 2602 89
rect 2547 20 2602 37
<< via1 >>
rect 66 853 269 861
rect 66 852 249 853
rect 249 852 269 853
rect 66 835 250 852
rect 250 835 269 852
rect 66 828 269 835
rect 60 742 67 804
rect 67 742 85 804
rect 85 742 107 804
rect 107 742 125 804
rect 125 742 130 804
rect 2405 852 2704 863
rect 2405 834 2704 852
rect 2405 828 2704 834
rect 2748 748 2756 824
rect 2756 748 2776 824
rect 2776 748 2783 824
rect 2645 219 2649 536
rect 2649 219 2684 536
rect 2684 219 2687 536
rect 2548 37 2600 89
<< metal2 >>
rect 0 863 2859 878
rect 0 861 2405 863
rect 0 828 66 861
rect 269 828 2405 861
rect 2704 828 2859 863
rect 0 824 2859 828
rect 0 804 2748 824
rect 0 742 60 804
rect 130 748 2748 804
rect 2783 748 2859 824
rect 130 742 2859 748
rect 0 738 2859 742
rect 47 737 140 738
rect 72 626 89 737
rect 2634 536 2698 549
rect 2634 248 2645 536
rect 0 219 2645 248
rect 2687 248 2698 536
rect 2687 219 2859 248
rect 0 108 2859 219
rect 2544 95 2807 108
rect 2544 89 2799 95
rect 2544 37 2548 89
rect 2600 44 2799 89
rect 2600 37 2606 44
<< labels >>
rlabel metal1 1253 0 1648 77 0 OUTPUT 
port 2 nsew
rlabel space 1 737 24 878 0 VGND
port 3 nsew
rlabel metal2 2823 738 2859 878 0 VGND
port 3 nsew
rlabel metal2 1 108 22 248 0 VINJ
port 4 nsew
rlabel metal2 2829 108 2859 248 0 VINJ
port 4 nsew
rlabel metal1 771 1040 1160 1087 0 INPUT
port 5 nsew
rlabel metal2 2620 44 2799 69 0 VINJ
port 4 nsew
rlabel metal1 70 50 142 84 0 VGND
port 3 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
