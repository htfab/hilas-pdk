magic
tech sky130A
timestamp 1628704286
<< checkpaint >>
rect -629 -630 2255 1679
<< error_s >>
rect 432 564 438 570
rect 537 564 543 570
rect 58 554 64 560
rect 111 554 117 560
rect 52 504 58 510
rect 117 504 123 510
rect 426 500 432 506
rect 543 500 549 506
rect 58 445 64 451
rect 111 445 117 451
rect 432 447 438 453
rect 537 447 543 453
rect 52 395 58 401
rect 117 395 123 401
rect 426 383 432 389
rect 543 383 549 389
rect 3635 307 3637 335
rect 432 262 438 268
rect 537 262 543 268
rect 58 256 64 262
rect 111 256 117 262
rect 52 206 58 212
rect 117 206 123 212
rect 426 198 432 204
rect 543 198 549 204
rect 432 146 438 152
rect 537 146 543 152
rect 58 139 64 145
rect 111 139 117 145
rect 52 89 58 95
rect 117 89 123 95
rect 426 82 432 88
rect 543 82 549 88
<< nwell >>
rect 1007 626 3542 627
rect 1008 619 3542 626
rect 1 559 12 577
rect 0 373 12 391
rect 2 74 12 91
rect 1006 28 3542 619
rect 1007 23 3542 28
rect 1200 22 3542 23
<< metal1 >>
rect 36 613 76 627
rect 280 621 304 627
rect 442 619 479 627
rect 673 620 697 627
rect 912 622 931 627
rect 956 622 972 627
rect 441 614 479 619
rect 440 35 441 37
rect 36 22 75 34
rect 280 22 304 29
rect 440 23 479 35
rect 440 22 441 23
rect 673 22 697 29
rect 875 23 891 29
rect 912 23 931 29
rect 956 23 972 29
<< metal2 >>
rect 1074 624 1125 627
rect 1074 622 1167 624
rect 1074 615 1130 622
rect 888 596 1130 615
rect 1117 594 1130 596
rect 1158 594 1167 622
rect 1 559 12 577
rect 898 559 3670 577
rect 892 516 3670 534
rect 898 416 3670 434
rect 3569 391 3670 392
rect 0 373 12 391
rect 894 373 3670 391
rect 3601 335 3670 342
rect 3601 307 3608 335
rect 3637 307 3670 335
rect 3601 301 3670 307
rect 2 258 12 275
rect 877 258 3670 275
rect 887 216 3670 233
rect 885 118 3670 135
rect 2 74 12 91
rect 881 74 3670 91
<< via2 >>
rect 1130 594 1158 622
rect 3608 307 3637 335
<< metal3 >>
rect 1125 622 1163 625
rect 1125 596 1130 622
rect 1117 594 1130 596
rect 1158 596 1163 622
rect 1158 594 1171 596
rect 1117 471 1171 594
rect 3523 335 3638 406
rect 3523 307 3608 335
rect 3637 307 3638 335
rect 1037 222 1055 252
rect 3523 242 3638 307
rect 3568 241 3638 242
rect 1146 101 1164 131
<< metal4 >>
rect 1279 560 1689 590
rect 1110 499 1380 510
rect 1110 469 1401 499
rect 1350 435 1401 469
rect 1651 440 1689 560
rect 1935 443 2263 473
rect 1041 397 1177 427
rect 1147 341 1177 397
rect 1935 341 1965 443
rect 2233 341 2263 443
rect 1147 311 2263 341
rect 2503 441 3392 471
rect 1371 252 1690 255
rect 1935 252 1965 255
rect 1037 222 2257 252
rect 1371 185 1401 222
rect 1660 188 1690 222
rect 1935 188 1965 222
rect 1660 185 1965 188
rect 2227 185 2257 222
rect 1371 155 2257 185
rect 2503 189 2533 441
rect 2786 438 3097 441
rect 2786 189 2816 438
rect 3067 189 3097 438
rect 3362 189 3392 441
rect 2503 159 3398 189
rect 3067 158 3398 159
rect 1134 101 1185 131
rect 1155 77 1185 101
rect 3368 77 3398 158
rect 1155 47 3398 77
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_1
timestamp 1628285143
transform 1 0 264 0 1 404
box -263 -404 1361 645
use sky130_hilas_cellAttempt01  sky130_hilas_cellAttempt01_0
timestamp 1628285143
transform 1 0 264 0 1 404
box -263 -404 1361 645
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1628285143
transform 1 0 876 0 1 603
box -9 -10 23 22
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1628285143
transform 1 0 876 0 1 603
box -9 -10 23 22
use sky130_hilas_m22m4  sky130_hilas_m22m4_3
timestamp 1607701799
transform 1 0 1107 0 1 131
box -36 -36 43 39
use sky130_hilas_m22m4  sky130_hilas_m22m4_2
timestamp 1607701799
transform 1 0 998 0 1 218
box -36 -36 43 39
use sky130_hilas_m22m4  sky130_hilas_m22m4_1
timestamp 1607701799
transform 1 0 1002 0 1 427
box -36 -36 43 39
<< labels >>
rlabel metal2 3658 301 3670 342 0 CAPTERM2
port 1 nsew analog default
rlabel metal2 1074 614 1125 627 0 CAPTERM1
port 2 nsew analog default
rlabel metal1 912 622 931 627 0 GATESELECT
port 4 nsew
rlabel metal1 956 622 972 627 0 VINJ
port 3 nsew power default
rlabel metal1 442 614 479 627 0 GATE
port 6 nsew analog default
rlabel metal1 36 613 76 627 0 VTUN
port 5 nsew
rlabel metal1 36 22 75 34 0 VTUN
port 5 nsew
rlabel metal1 440 23 479 35 0 GATE
port 6 nsew
rlabel metal1 956 23 972 29 0 VINJ
rlabel metal1 875 23 891 29 0 CAPTERM1
rlabel metal1 912 23 931 29 0 GATESELECT
rlabel metal2 1 559 12 577 0 DRAIN1
port 8 nsew
rlabel metal2 0 373 12 391 0 DRAIN2
port 7 nsew
rlabel metal2 3660 74 3670 91 0 DRAIN4
port 10 nsew
rlabel metal2 3660 559 3670 577 0 DRAIN1
port 8 nsew
rlabel metal2 3659 373 3670 392 0 DRAIN2
port 7 nsew
rlabel metal2 3659 258 3670 275 0 DRAIN3
port 11 nsew
rlabel metal2 2 258 12 275 0 DRAIN3
port 11 nsew
rlabel metal2 2 74 12 91 0 DRAIN4
port 10 nsew
rlabel metal1 280 621 304 627 0 VGND
port 12 nsew
rlabel metal1 673 620 697 627 0 VGND
port 12 nsew
rlabel metal1 280 22 304 29 0 VGND
port 12 nsew
rlabel metal1 673 22 697 29 0 VGND
port 12 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
