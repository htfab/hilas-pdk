magic
tech sky130A
timestamp 1628707377
<< error_p >>
rect 31 48 58 55
rect 31 6 58 13
<< nmos >>
rect 31 13 58 48
<< ndiff >>
rect 0 39 31 48
rect 0 22 5 39
rect 25 22 31 39
rect 0 13 31 22
rect 58 39 89 48
rect 58 22 64 39
rect 84 22 89 39
rect 58 13 89 22
<< ndiffc >>
rect 5 22 25 39
rect 64 22 84 39
<< poly >>
rect 31 48 58 61
rect 31 0 58 13
<< locali >>
rect 5 39 25 47
rect 5 14 25 22
rect 64 39 84 47
rect 64 14 84 22
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
