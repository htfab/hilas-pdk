magic
tech sky130A
timestamp 1628704264
<< error_p >>
rect 0 23 23 29
rect 0 6 3 23
rect 0 0 23 6
<< locali >>
rect 2 23 21 26
rect 2 6 3 23
rect 20 6 21 23
rect 2 3 21 6
<< viali >>
rect 3 6 20 23
<< metal1 >>
rect 0 23 23 29
rect 0 6 3 23
rect 20 6 23 23
rect 0 0 23 6
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
