magic
tech sky130A
timestamp 1634057794
<< psubdiff >>
rect 12 24 634 32
rect 12 7 27 24
rect 44 7 634 24
rect 12 0 634 7
<< psubdiffcont >>
rect 27 7 44 24
<< poly >>
rect 24 69 68 82
rect 24 52 37 69
rect 54 52 68 69
rect 24 40 68 52
rect 581 71 627 82
rect 581 54 596 71
rect 613 54 630 71
rect 581 40 627 54
<< polycont >>
rect 37 52 54 69
rect 596 54 613 71
<< npolyres >>
rect 68 40 581 82
<< locali >>
rect 54 52 62 69
rect 588 54 596 71
rect 588 52 630 54
rect 16 7 27 24
<< viali >>
rect 20 52 37 69
rect 613 54 630 71
rect 44 7 61 24
<< metal1 >>
rect 0 69 57 74
rect 0 52 20 69
rect 37 52 57 69
rect 0 47 57 52
rect 596 71 649 77
rect 596 54 613 71
rect 630 54 649 71
rect 596 47 649 54
rect 41 24 67 27
rect 15 20 44 24
rect 0 7 44 20
rect 61 7 67 24
rect 0 4 67 7
<< labels >>
rlabel metal1 1 47 10 74 0 TERM1
port 1 nsew
rlabel metal1 637 47 649 77 0 TERM2
port 2 nsew
rlabel metal1 0 4 9 20 0 VGND
port 3 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
