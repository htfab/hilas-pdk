**.subckt pFETLarge Well Source1p Gate1p Drain1p
*.iopin Well
*.iopin Source1p
*.ipin Gate1p
*.iopin Drain1p
XM1 Source1p Gate1p Drain1p Well sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
**.ends
** flattened .save nodes
.end
