magic
tech sky130A
timestamp 1628704422
<< error_p >>
rect 50 180 79 208
rect 129 180 158 208
rect 208 180 237 208
rect 28 173 258 180
rect 28 158 35 173
rect 50 167 79 173
rect 129 167 158 173
rect 208 167 237 173
rect 50 158 51 159
rect 78 158 79 159
rect 129 158 130 159
rect 157 158 158 159
rect 208 158 209 159
rect 236 158 237 159
rect 251 158 258 173
rect 0 129 41 158
rect 49 157 80 158
rect 128 157 159 158
rect 207 157 238 158
rect 50 130 79 157
rect 129 130 158 157
rect 208 130 237 157
rect 49 129 80 130
rect 128 129 159 130
rect 207 129 238 130
rect 245 129 287 158
rect 28 79 35 129
rect 50 128 51 129
rect 78 128 79 129
rect 129 128 130 129
rect 157 128 158 129
rect 208 128 209 129
rect 236 128 237 129
rect 50 79 51 80
rect 78 79 79 80
rect 129 79 130 80
rect 157 79 158 80
rect 208 79 209 80
rect 236 79 237 80
rect 251 79 258 129
rect 0 50 41 79
rect 49 78 80 79
rect 128 78 159 79
rect 207 78 238 79
rect 50 51 79 78
rect 129 51 158 78
rect 208 51 237 78
rect 49 50 80 51
rect 128 50 159 51
rect 207 50 238 51
rect 245 50 287 79
rect 28 35 35 50
rect 50 49 51 50
rect 78 49 79 50
rect 129 49 130 50
rect 157 49 158 50
rect 208 49 209 50
rect 236 49 237 50
rect 50 35 79 41
rect 129 35 158 41
rect 208 35 237 41
rect 251 35 258 50
rect 28 28 258 35
rect 50 0 79 28
rect 129 0 158 28
rect 208 0 237 28
<< nwell >>
rect 6 6 278 202
<< mvpmos >>
rect 41 158 245 167
rect 41 129 50 158
rect 79 129 129 158
rect 158 129 208 158
rect 237 129 245 158
rect 41 79 245 129
rect 41 50 50 79
rect 79 50 129 79
rect 158 50 208 79
rect 237 50 245 79
rect 41 41 245 50
<< mvpdiff >>
rect 50 152 79 158
rect 50 135 56 152
rect 73 135 79 152
rect 50 129 79 135
rect 129 152 158 158
rect 129 135 135 152
rect 152 135 158 152
rect 129 129 158 135
rect 208 152 237 158
rect 208 135 214 152
rect 231 135 237 152
rect 208 129 237 135
rect 50 72 79 79
rect 50 56 56 72
rect 73 56 79 72
rect 50 50 79 56
rect 129 72 158 79
rect 129 56 135 72
rect 152 56 158 72
rect 129 50 158 56
rect 208 73 237 79
rect 208 56 214 73
rect 231 56 237 73
rect 208 50 237 56
<< mvpdiffc >>
rect 56 135 73 152
rect 135 135 152 152
rect 214 135 231 152
rect 56 56 73 72
rect 135 56 152 72
rect 214 56 231 73
<< poly >>
rect 35 167 251 173
rect 35 41 41 167
rect 245 41 251 167
rect 35 35 251 41
<< locali >>
rect 46 152 241 162
rect 46 135 56 152
rect 73 145 135 152
rect 73 135 94 145
rect 46 128 94 135
rect 111 135 135 145
rect 152 135 214 152
rect 231 135 241 152
rect 111 128 241 135
rect 46 111 241 128
rect 46 94 94 111
rect 111 94 241 111
rect 46 77 241 94
rect 46 72 94 77
rect 46 56 56 72
rect 73 60 94 72
rect 111 73 241 77
rect 111 72 214 73
rect 111 60 135 72
rect 73 56 135 60
rect 152 56 214 72
rect 231 56 241 73
rect 46 45 241 56
<< viali >>
rect 94 128 111 145
rect 94 94 111 111
rect 94 60 111 77
<< metal1 >>
rect 90 145 116 151
rect 90 128 94 145
rect 111 128 116 145
rect 90 111 116 128
rect 90 103 94 111
rect 89 94 94 103
rect 111 94 116 111
rect 89 77 116 94
rect 89 60 94 77
rect 111 60 116 77
rect 89 51 116 60
rect 89 6 115 51
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
