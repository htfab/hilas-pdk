* Copyright 2020 The Hilas PDK Authors
* 
* This file is part of HILAS.
* 
* HILAS is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published by
* the Free Software Foundation, version 3 of the License.
* 
* HILAS is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
* 
* You should have received a copy of the GNU Lesser General Public License
* along with HILAS.  If not, see <https://www.gnu.org/licenses/>.
* 
* Licensed under the Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
* https://www.gnu.org/licenses/lgpl-3.0.en.html
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
* SPDX-License-Identifier: LGPL-3.0
* 
* 

* NGSPICE file created from sky130_hilas_DAC6TransistorStack01c.ext - technology: sky130A

.subckt sky130_hilas_pFETdevice01b VSUBS w_n158_n156#
X0 a_42_n38# a_n36_n84# a_n90_n38# w_n158_n156# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends

.subckt sky130_hilas_pFETdevice01 VSUBS w_n158_n156#
X0 a_42_n38# a_n158_36# a_n90_n38# w_n158_n156# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends

.subckt sky130_hilas_pFETdevice01aa VSUBS w_n160_n156#
X0 a_42_n38# a_n160_36# a_n92_n38# w_n160_n156# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends

.subckt sky130_hilas_pFETdevice01a VSUBS w_n160_n84#
X0 a_42_n38# a_n160_36# a_n92_n38# w_n160_n84# sky130_fd_pr__pfet_01v8 w=390000u l=390000u
.ends


* Top level circuit sky130_hilas_DAC6TransistorStack01c

Xsky130_hilas_pFETdevice01b_1 VSUBS sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01b
Xsky130_hilas_pFETdevice01_0 VSUBS sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01_3 VSUBS sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01_6 VSUBS sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01
Xsky130_hilas_pFETdevice01aa_0 VSUBS sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01aa
Xsky130_hilas_pFETdevice01a_0 VSUBS sky130_hilas_pFETdevice01a_0/w_n160_n84# sky130_hilas_pFETdevice01a
.end

