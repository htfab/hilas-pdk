magic
tech sky130A
timestamp 1628698506
<< nmos >>
rect -5 0 1 3
<< pmos >>
rect 26 0 32 3
<< ndiff >>
rect -5 9 1 10
rect -5 5 -4 9
rect 0 5 1 9
rect -5 3 1 5
rect -5 -2 1 0
rect -5 -6 -4 -2
rect 0 -6 1 -2
rect -5 -7 1 -6
<< pdiff >>
rect 26 10 32 11
rect 26 6 27 10
rect 31 6 32 10
rect 26 3 32 6
rect 26 -3 32 0
rect 26 -7 27 -3
rect 31 -7 32 -3
rect 26 -8 32 -7
<< ndiffc >>
rect -4 5 0 9
rect -4 -6 0 -2
<< pdiffc >>
rect 27 6 31 10
rect 27 -7 31 -3
<< poly >>
rect -8 0 -5 3
rect 1 0 26 3
rect 32 0 34 3
rect 11 -3 14 0
rect 9 -4 15 -3
rect 9 -8 10 -4
rect 14 -8 15 -4
rect 9 -9 15 -8
<< metal1 >>
rect 10 9 14 16
rect 0 6 27 9
rect 0 5 31 6
rect -8 -6 -4 -2
rect 31 -7 34 -3
rect 10 -15 14 -8
<< via1 >>
rect -12 -6 -8 -2
rect 34 -7 38 -3
<< metal2 >>
rect -13 -2 -7 15
rect -13 -6 -12 -2
rect -8 -6 -7 -2
rect -13 -12 -7 -6
rect 33 -3 39 15
rect 33 -7 34 -3
rect 38 -7 39 -3
rect 33 -12 39 -7
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
