magic
tech sky130A
timestamp 1634057824
<< psubdiff >>
rect 34 873 5355 877
rect 34 856 72 873
rect 5335 856 5355 873
rect 34 853 5355 856
rect 34 850 58 853
rect 34 90 38 850
rect 55 90 58 850
rect 5491 851 5515 877
rect 34 74 58 90
rect 5491 142 5495 851
rect 5512 142 5515 851
rect 5491 122 5515 142
<< psubdiffcont >>
rect 72 856 5335 873
rect 38 90 55 850
rect 5495 142 5512 851
<< poly >>
rect 2107 1003 2156 1025
rect 2107 986 2117 1003
rect 2134 986 2156 1003
rect 2107 967 2156 986
rect 2107 950 2117 967
rect 2134 950 2156 967
rect 2107 931 2156 950
rect 2107 914 2117 931
rect 2134 914 2156 931
rect 2754 1020 2819 1025
rect 2754 1003 2792 1020
rect 2809 1003 2819 1020
rect 2754 986 2819 1003
rect 2754 969 2792 986
rect 2809 969 2819 986
rect 2754 952 2819 969
rect 2754 935 2792 952
rect 2809 935 2819 952
rect 2107 890 2156 914
rect 2754 918 2819 935
rect 2754 901 2792 918
rect 2809 901 2819 918
rect 2754 890 2819 901
rect 5370 869 5476 875
rect 5370 852 5379 869
rect 5467 852 5476 869
rect 5370 847 5476 852
rect 5330 845 5476 847
rect 67 829 5476 845
rect 67 803 83 829
rect 5370 828 5476 829
rect 67 787 5479 803
rect 67 761 83 762
rect 5463 761 5479 787
rect 67 745 5479 761
rect 67 722 83 745
rect 67 706 5479 722
rect 5463 681 5479 706
rect 67 665 5479 681
rect 67 643 83 665
rect 67 627 5479 643
rect 67 604 83 605
rect 5463 604 5479 627
rect 67 588 5479 604
rect 67 564 83 588
rect 67 548 5479 564
rect 67 526 83 527
rect 5463 526 5479 548
rect 67 510 5479 526
rect 67 484 83 510
rect 67 468 5479 484
rect 5463 443 5479 468
rect 67 427 5479 443
rect 67 406 82 427
rect 67 390 5479 406
rect 5463 368 5479 390
rect 67 352 5479 368
rect 67 330 83 352
rect 67 314 5479 330
rect 5463 291 5479 314
rect 67 275 5479 291
rect 67 253 83 275
rect 67 237 5479 253
rect 5463 215 5479 237
rect 69 199 5479 215
rect 69 178 85 199
rect 69 162 5480 178
rect 5464 141 5480 162
rect 72 125 5480 141
rect 72 103 88 125
rect 72 87 5479 103
rect 5463 64 5479 87
rect 2687 56 5479 64
rect 2682 39 2699 56
rect 2716 39 2733 56
rect 2750 39 2767 56
rect 2784 39 2801 56
rect 2818 39 2835 56
rect 2852 39 2869 56
rect 2886 48 5479 56
rect 2886 39 2923 48
rect 2687 30 2923 39
<< polycont >>
rect 2117 986 2134 1003
rect 2117 950 2134 967
rect 2117 914 2134 931
rect 2792 1003 2809 1020
rect 2792 969 2809 986
rect 2792 935 2809 952
rect 2792 901 2809 918
rect 5379 852 5467 869
rect 2699 39 2716 56
rect 2733 39 2750 56
rect 2767 39 2784 56
rect 2801 39 2818 56
rect 2835 39 2852 56
rect 2869 39 2886 56
<< npolyres >>
rect 2156 925 2754 1025
<< locali >>
rect 2114 1021 2136 1024
rect 2114 1004 2117 1021
rect 2134 1004 2136 1021
rect 2114 1003 2136 1004
rect 2114 986 2117 1003
rect 2134 986 2136 1003
rect 2114 985 2136 986
rect 2114 968 2117 985
rect 2134 968 2136 985
rect 2114 967 2136 968
rect 2114 950 2117 967
rect 2134 950 2136 967
rect 2114 949 2136 950
rect 2114 932 2117 949
rect 2134 932 2136 949
rect 2114 931 2136 932
rect 2114 914 2117 931
rect 2134 914 2136 931
rect 2114 913 2136 914
rect 2114 912 2117 913
rect 2109 896 2117 912
rect 2134 912 2136 913
rect 2788 1020 2812 1028
rect 2788 987 2792 1020
rect 2809 987 2812 1020
rect 2788 986 2812 987
rect 2788 969 2792 986
rect 2809 969 2812 986
rect 2788 968 2812 969
rect 2788 935 2792 968
rect 2809 935 2812 968
rect 2788 932 2812 935
rect 2134 896 2142 912
rect 2109 893 2142 896
rect 2788 901 2792 932
rect 2809 901 2812 932
rect 2788 893 2812 901
rect 38 856 72 873
rect 5335 869 5512 873
rect 5335 856 5379 869
rect 38 852 5379 856
rect 38 850 72 852
rect 55 835 72 850
rect 2462 846 3350 852
rect 2462 835 2472 846
rect 55 833 2472 835
rect 3341 835 3350 846
rect 5467 851 5512 869
rect 5467 835 5495 851
rect 3341 833 5495 835
rect 5495 125 5512 142
rect 38 73 55 90
rect 2716 39 2719 56
rect 2750 39 2756 56
rect 2784 39 2792 56
rect 2818 39 2828 56
rect 2852 39 2864 56
rect 2886 39 2901 56
<< viali >>
rect 2117 1004 2134 1021
rect 2117 968 2134 985
rect 2117 932 2134 949
rect 2117 896 2134 913
rect 2792 1003 2809 1004
rect 2792 987 2809 1003
rect 2792 952 2809 968
rect 2792 951 2809 952
rect 2792 918 2809 932
rect 2792 915 2809 918
rect 72 835 2462 852
rect 3350 835 5467 852
rect 2682 39 2699 56
rect 2719 39 2733 56
rect 2733 39 2736 56
rect 2756 39 2767 56
rect 2767 39 2773 56
rect 2792 39 2801 56
rect 2801 39 2809 56
rect 2828 39 2835 56
rect 2835 39 2845 56
rect 2864 39 2869 56
rect 2869 39 2882 56
rect 2901 39 2918 56
<< metal1 >>
rect 2106 1025 2347 1089
rect 2108 1021 2149 1025
rect 2108 1004 2117 1021
rect 2134 1004 2149 1021
rect 2108 985 2149 1004
rect 2108 968 2117 985
rect 2134 968 2149 985
rect 2108 949 2149 968
rect 2781 1004 2822 1036
rect 2781 987 2792 1004
rect 2809 987 2822 1004
rect 2781 968 2822 987
rect 2781 959 2792 968
rect 2108 932 2117 949
rect 2134 932 2149 949
rect 2108 913 2149 932
rect 2108 896 2117 913
rect 2134 896 2149 913
rect 2108 890 2149 896
rect 2754 951 2792 959
rect 2809 951 2822 968
rect 2754 932 2822 951
rect 2754 915 2792 932
rect 2809 915 2923 932
rect 2754 889 2923 915
rect 33 871 2470 873
rect 27 867 2470 871
rect 27 852 82 867
rect 27 835 72 852
rect 2462 835 2470 867
rect 27 832 2470 835
rect 27 7 68 832
rect 2687 82 2923 889
rect 3350 872 5486 873
rect 3344 867 5486 872
rect 3344 835 3350 867
rect 5436 852 5486 867
rect 5467 835 5486 852
rect 3344 833 5486 835
rect 3344 832 5470 833
rect 2675 56 2923 82
rect 2675 39 2682 56
rect 2699 39 2719 56
rect 2736 39 2756 56
rect 2773 39 2792 56
rect 2809 39 2828 56
rect 2845 39 2864 56
rect 2882 39 2901 56
rect 2918 39 2923 56
rect 2675 0 2923 39
<< via1 >>
rect 82 852 2462 867
rect 82 841 2462 852
rect 3350 852 5436 867
rect 3350 841 5436 852
<< metal2 >>
rect 0 867 5547 877
rect 0 841 82 867
rect 2462 841 3350 867
rect 5436 841 5547 867
rect 0 738 5547 841
rect 0 108 5547 248
<< labels >>
rlabel metal1 2107 1040 2345 1079 0 INPUT
port 2 nsew
rlabel metal1 2675 0 2923 27 0 OUTPUT
port 3 nsew
rlabel metal1 27 7 68 18 0 VGND
port 4 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
