magic
tech sky130A
timestamp 1628616956
<< nwell >>
rect 0 0 186 299
<< mvpmos >>
rect 65 48 115 251
<< mvpdiff >>
rect 34 244 65 251
rect 34 227 41 244
rect 58 227 65 244
rect 34 210 65 227
rect 34 193 41 210
rect 58 193 65 210
rect 34 176 65 193
rect 34 159 41 176
rect 58 159 65 176
rect 34 142 65 159
rect 34 125 41 142
rect 58 125 65 142
rect 34 108 65 125
rect 34 91 41 108
rect 58 91 65 108
rect 34 74 65 91
rect 34 57 41 74
rect 58 57 65 74
rect 34 48 65 57
rect 115 243 153 251
rect 115 226 122 243
rect 139 226 153 243
rect 115 209 153 226
rect 115 192 122 209
rect 139 192 153 209
rect 115 175 153 192
rect 115 158 122 175
rect 139 158 153 175
rect 115 141 153 158
rect 115 124 122 141
rect 139 124 153 141
rect 115 107 153 124
rect 115 90 122 107
rect 139 90 153 107
rect 115 73 153 90
rect 115 56 122 73
rect 139 56 153 73
rect 115 48 153 56
<< mvpdiffc >>
rect 41 227 58 244
rect 41 193 58 210
rect 41 159 58 176
rect 41 125 58 142
rect 41 91 58 108
rect 41 57 58 74
rect 122 226 139 243
rect 122 192 139 209
rect 122 158 139 175
rect 122 124 139 141
rect 122 90 139 107
rect 122 56 139 73
<< poly >>
rect 65 251 115 269
rect 65 33 115 48
<< locali >>
rect 41 244 59 252
rect 58 227 59 244
rect 41 210 59 227
rect 58 193 59 210
rect 41 176 59 193
rect 58 159 59 176
rect 41 142 59 159
rect 58 125 59 142
rect 41 108 59 125
rect 58 91 59 108
rect 41 74 59 91
rect 58 57 59 74
rect 122 243 139 251
rect 122 209 139 226
rect 122 175 139 192
rect 122 141 139 158
rect 122 107 139 124
rect 122 73 139 90
rect 41 47 59 57
rect 114 56 122 73
rect 139 56 147 73
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
