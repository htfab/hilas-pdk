magic
tech sky130A
magscale 1 2
timestamp 1632256364
<< error_s >>
rect 28350 2014 28384 2236
rect 28418 2014 28452 2210
rect 28614 2014 30928 2022
rect 31032 2014 31066 2210
rect 31100 2014 31134 2206
rect 31332 2060 31918 2076
rect 32082 2060 32238 2076
rect 31214 2022 31276 2048
rect 31332 2022 31890 2048
rect 32110 2022 32210 2048
rect 31276 2014 31890 2022
rect 32136 2014 32210 2022
rect 21298 1980 31864 2014
rect 31865 2006 32135 2014
rect 31879 1999 32135 2006
rect 28350 1972 28410 1980
rect 28418 1972 28452 1980
rect 28454 1972 28490 1980
rect 28614 1974 28676 1980
rect 28614 1972 28629 1973
rect 28661 1972 28676 1973
rect 31032 1972 31066 1980
rect 31100 1972 31134 1980
rect 31276 1975 31864 1980
rect 31214 1974 31864 1975
rect 31894 1996 32135 1999
rect 31276 1972 31286 1974
rect 31394 1972 31409 1973
rect 31894 1972 32106 1996
rect 27854 1967 32106 1972
rect 27854 1952 32121 1967
rect 32136 1952 32184 2014
rect 27854 1938 32088 1952
rect 32136 1938 32137 1952
rect 32184 1938 32210 1952
rect 28334 1926 28490 1938
rect 28334 1915 28345 1926
rect 28334 1874 28345 1885
rect 28374 1874 28410 1926
rect 28454 1874 28490 1926
rect 28614 1926 28676 1938
rect 28692 1932 30888 1938
rect 28614 1911 28629 1926
rect 28661 1918 28676 1926
rect 31022 1926 31148 1938
rect 28661 1911 30928 1918
rect 31022 1915 31033 1926
rect 31137 1915 31148 1926
rect 31276 1926 31332 1938
rect 31276 1915 31287 1926
rect 31321 1915 31332 1926
rect 31438 1904 33328 1938
rect 28334 1862 28490 1874
rect 28614 1874 28629 1889
rect 30913 1874 30928 1889
rect 28334 1842 28468 1862
rect 28334 1831 28345 1842
rect 28457 1831 28468 1842
rect 28614 1858 30928 1874
rect 31022 1874 31033 1885
rect 31137 1874 31148 1885
rect 28614 1842 28676 1858
rect 28614 1827 28629 1842
rect 28661 1827 28676 1842
rect 31022 1842 31148 1874
rect 31022 1831 31033 1842
rect 31137 1831 31148 1842
rect 31276 1874 31287 1885
rect 31321 1874 31332 1885
rect 32136 1878 32137 1904
rect 32184 1878 32210 1904
rect 31276 1842 31332 1874
rect 31276 1831 31287 1842
rect 31321 1831 31332 1842
rect 31402 1874 31417 1878
rect 31402 1842 32112 1874
rect 31402 1827 31417 1842
rect 32080 1829 32112 1842
rect 32065 1814 32127 1829
rect 32136 1814 32184 1878
rect 28334 1790 28345 1801
rect 28457 1790 28468 1801
rect 28334 1758 28468 1790
rect 28334 1747 28345 1758
rect 28457 1747 28468 1758
rect 28614 1790 28629 1805
rect 30913 1790 30928 1798
rect 28614 1758 30928 1790
rect 28614 1743 28629 1758
rect 30913 1743 30928 1758
rect 31022 1790 31033 1801
rect 31137 1790 31148 1801
rect 31022 1758 31148 1790
rect 31022 1747 31033 1758
rect 31137 1747 31148 1758
rect 31276 1790 31287 1801
rect 31321 1790 31332 1801
rect 31276 1758 31332 1790
rect 31276 1747 31287 1758
rect 31321 1747 31332 1758
rect 28334 1712 28345 1723
rect 28457 1712 28468 1723
rect 28334 1680 28468 1712
rect 28334 1669 28345 1680
rect 28457 1669 28468 1680
rect 28614 1712 28629 1727
rect 28661 1712 28676 1727
rect 31276 1723 31286 1747
rect 32136 1730 32137 1814
rect 32184 1730 32210 1814
rect 28614 1680 28676 1712
rect 28614 1666 28629 1680
rect 28661 1678 28676 1680
rect 31022 1712 31033 1723
rect 31137 1712 31148 1723
rect 31022 1680 31148 1712
rect 28614 1665 28626 1666
rect 28661 1665 30928 1678
rect 31022 1669 31033 1680
rect 31137 1669 31148 1680
rect 31276 1712 31287 1723
rect 31321 1712 31332 1723
rect 31276 1680 31332 1712
rect 31276 1669 31287 1680
rect 31321 1669 31332 1680
rect 31412 1712 31427 1727
rect 31412 1681 32112 1712
rect 31412 1680 32127 1681
rect 28334 1630 28345 1641
rect 28457 1630 28468 1641
rect 28334 1598 28468 1630
rect 28334 1587 28345 1598
rect 28457 1587 28468 1598
rect 28614 1630 28629 1645
rect 30913 1630 30928 1645
rect 31276 1641 31286 1669
rect 31412 1666 31427 1680
rect 32065 1666 32127 1680
rect 32136 1666 32184 1730
rect 28614 1620 30928 1630
rect 31022 1630 31033 1641
rect 31137 1630 31148 1641
rect 28614 1598 28676 1620
rect 28614 1583 28629 1598
rect 28661 1583 28676 1598
rect 31022 1598 31148 1630
rect 31022 1587 31033 1598
rect 31137 1587 31148 1598
rect 31276 1630 31287 1641
rect 31321 1630 31332 1641
rect 31276 1598 31332 1630
rect 31276 1587 31287 1598
rect 31321 1587 31332 1598
rect 32136 1592 32137 1666
rect 32184 1592 32210 1666
rect 28334 1554 28345 1565
rect 28457 1554 28468 1565
rect 28334 1522 28468 1554
rect 28334 1511 28345 1522
rect 28457 1511 28468 1522
rect 28614 1554 28629 1569
rect 31276 1565 31286 1587
rect 31412 1583 32127 1592
rect 30913 1554 30928 1560
rect 28614 1522 30928 1554
rect 28614 1507 28629 1522
rect 30913 1507 30928 1522
rect 31022 1554 31033 1565
rect 31137 1554 31148 1565
rect 31022 1522 31148 1554
rect 31022 1511 31033 1522
rect 31137 1511 31148 1522
rect 31276 1554 31287 1565
rect 31321 1554 31332 1565
rect 31276 1522 31332 1554
rect 31412 1554 31427 1569
rect 31412 1543 32112 1554
rect 31412 1528 32127 1543
rect 32136 1528 32184 1592
rect 31276 1511 31287 1522
rect 31321 1511 31332 1522
rect 28334 1476 28345 1487
rect 28457 1476 28468 1487
rect 28334 1444 28468 1476
rect 28334 1433 28345 1444
rect 28457 1433 28468 1444
rect 28614 1476 28629 1491
rect 28661 1476 28676 1491
rect 31276 1487 31286 1511
rect 28614 1444 28676 1476
rect 28614 1430 28629 1444
rect 28661 1442 28676 1444
rect 31022 1476 31033 1487
rect 31137 1476 31148 1487
rect 31022 1444 31148 1476
rect 28614 1429 28626 1430
rect 28661 1429 30928 1442
rect 31022 1433 31033 1444
rect 31137 1433 31148 1444
rect 31276 1476 31287 1487
rect 31321 1476 31332 1487
rect 31276 1444 31332 1476
rect 32136 1462 32137 1528
rect 32184 1462 32210 1528
rect 31276 1433 31287 1444
rect 31321 1433 31332 1444
rect 31404 1447 32127 1462
rect 31404 1444 32112 1447
rect 28334 1396 28345 1407
rect 28457 1396 28468 1407
rect 28334 1364 28468 1396
rect 28334 1353 28345 1364
rect 28457 1353 28468 1364
rect 28614 1396 28629 1411
rect 30913 1396 30928 1411
rect 31276 1407 31286 1433
rect 31404 1429 31419 1444
rect 28614 1382 30928 1396
rect 28614 1364 28676 1382
rect 30866 1380 30928 1382
rect 31022 1396 31033 1407
rect 31137 1396 31148 1407
rect 28614 1349 28629 1364
rect 28661 1349 28676 1364
rect 31022 1364 31148 1396
rect 31022 1353 31033 1364
rect 31137 1353 31148 1364
rect 31276 1396 31287 1407
rect 31321 1396 31332 1407
rect 31404 1396 32127 1411
rect 32136 1396 32184 1462
rect 31276 1364 31332 1396
rect 31276 1353 31287 1364
rect 31321 1353 31332 1364
rect 28334 1320 28345 1331
rect 28457 1320 28468 1331
rect 28334 1288 28468 1320
rect 28334 1277 28345 1288
rect 28457 1277 28468 1288
rect 28614 1320 28629 1335
rect 31276 1331 31286 1353
rect 32136 1334 32137 1396
rect 32184 1334 32210 1396
rect 31022 1320 31033 1331
rect 31137 1320 31148 1331
rect 28614 1288 30928 1320
rect 28614 1273 28629 1288
rect 30913 1273 30928 1288
rect 31022 1288 31148 1320
rect 31022 1277 31033 1288
rect 31137 1277 31148 1288
rect 31276 1320 31287 1331
rect 31321 1320 31332 1331
rect 31276 1288 31332 1320
rect 31276 1277 31287 1288
rect 31321 1277 31332 1288
rect 31404 1320 31419 1334
rect 32065 1320 32127 1334
rect 31404 1319 32127 1320
rect 31404 1288 32112 1319
rect 31404 1273 31419 1288
rect 32136 1268 32184 1334
rect 28334 1236 28345 1247
rect 28457 1236 28468 1247
rect 28334 1204 28468 1236
rect 28334 1193 28345 1204
rect 28457 1193 28468 1204
rect 28614 1236 28629 1251
rect 28661 1236 28676 1251
rect 28614 1204 28676 1236
rect 28614 1189 28629 1204
rect 28661 1198 28676 1204
rect 31022 1236 31033 1247
rect 31137 1236 31148 1247
rect 31022 1204 31148 1236
rect 28661 1189 30928 1198
rect 31022 1193 31033 1204
rect 31137 1193 31148 1204
rect 31276 1236 31287 1247
rect 31321 1236 31332 1247
rect 31276 1204 31332 1236
rect 32136 1208 32137 1268
rect 32184 1208 32210 1268
rect 31276 1193 31287 1204
rect 31321 1193 31332 1204
rect 31404 1204 32127 1208
rect 28334 1154 28345 1165
rect 28457 1154 28468 1165
rect 28334 1122 28468 1154
rect 28334 1111 28345 1122
rect 28457 1111 28468 1122
rect 28614 1154 28629 1169
rect 30913 1154 30928 1169
rect 31276 1165 31286 1193
rect 31404 1189 31419 1204
rect 32080 1193 32127 1204
rect 28614 1138 30928 1154
rect 31022 1154 31033 1165
rect 31137 1154 31148 1165
rect 28614 1122 28676 1138
rect 28614 1107 28629 1122
rect 28661 1107 28676 1122
rect 31022 1122 31148 1154
rect 31022 1111 31033 1122
rect 31137 1111 31148 1122
rect 31276 1154 31287 1165
rect 31321 1154 31332 1165
rect 31276 1122 31332 1154
rect 31404 1154 31419 1169
rect 32080 1161 32112 1193
rect 32080 1154 32127 1161
rect 31404 1146 32127 1154
rect 32136 1146 32184 1208
rect 31276 1111 31287 1122
rect 31321 1111 31332 1122
rect 28334 1080 28345 1091
rect 28457 1080 28468 1091
rect 28334 1048 28468 1080
rect 28614 1080 28629 1095
rect 28661 1080 28676 1095
rect 32136 1092 32144 1146
rect 32184 1092 32210 1146
rect 28614 1078 28676 1080
rect 31022 1080 31033 1091
rect 31137 1080 31148 1091
rect 28334 1037 28345 1048
rect 28457 1037 28468 1048
rect 28612 1048 30928 1078
rect 28612 1033 28627 1048
rect 30913 1033 30928 1048
rect 31022 1048 31148 1080
rect 31022 1037 31033 1048
rect 31137 1037 31148 1048
rect 31264 1080 31275 1091
rect 31264 1048 32112 1080
rect 31264 1037 31275 1048
rect 32080 1047 32112 1048
rect 32069 1036 32123 1047
rect 32136 1036 32184 1092
rect 28612 1018 30928 1019
rect 28334 1004 28345 1015
rect 28457 1004 28468 1015
rect 28334 972 28468 1004
rect 28334 961 28345 972
rect 28457 961 28468 972
rect 31022 1004 31033 1015
rect 31137 1004 31148 1015
rect 31022 972 31148 1004
rect 32136 994 32137 1036
rect 31022 961 31033 972
rect 31137 966 31148 972
rect 31137 961 32123 966
rect 32144 946 32178 1036
rect 32184 994 32210 1036
rect 28334 928 28345 939
rect 28482 928 33684 946
rect 28334 912 33684 928
rect 28334 896 32112 912
rect 28334 885 28345 896
rect 32080 878 32112 896
rect 32144 878 32178 912
rect 28334 856 28347 861
rect 28336 850 28347 856
rect 28482 850 33684 878
rect 28336 844 33684 850
rect 28336 839 32112 844
rect 28336 832 32123 839
rect 28336 824 28468 832
rect 30800 828 32123 832
rect 28336 822 28438 824
rect 32144 552 32178 844
<< metal1 >>
rect 52 2328 830 2488
rect 5770 2328 6548 2488
rect 11488 2328 12266 2488
rect 19868 2332 20646 2492
rect 28292 2328 29070 2488
rect 34010 2328 34788 2488
rect 39730 2328 40508 2488
rect 45448 2328 46226 2488
rect 51164 2328 51942 2488
rect 56882 2328 57660 2488
rect 62602 2328 63380 2488
rect 1016 0 1806 154
rect 6736 0 7526 154
rect 12452 0 13242 154
rect 21006 0 21502 154
rect 29256 2 30046 156
rect 34974 0 35764 154
rect 40692 0 41482 154
rect 46410 0 47200 154
rect 52130 0 52920 154
rect 57846 0 58636 154
rect 63564 0 64354 154
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_1
timestamp 1632251427
transform 1 0 5718 0 1 612
box 0 0 5718 2174
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_0
timestamp 1632251427
transform 1 0 0 0 1 612
box 0 0 5718 2174
use sky130_hilas_polyresistorGND  sky130_hilas_polyresistorGND_0
timestamp 1632251351
transform 1 0 21154 0 1 268
box 0 0 11094 2178
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_2
timestamp 1632251427
transform 1 0 11436 0 1 612
box 0 0 5718 2174
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_3
timestamp 1632251427
transform 1 0 28240 0 1 612
box 0 0 5718 2174
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_4
timestamp 1632251427
transform 1 0 33958 0 1 612
box 0 0 5718 2174
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_5
timestamp 1632251427
transform 1 0 39676 0 1 612
box 0 0 5718 2174
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_6
timestamp 1632251427
transform 1 0 45394 0 1 612
box 0 0 5718 2174
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_9
timestamp 1632251427
transform 1 0 51112 0 1 612
box 0 0 5718 2174
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_7
timestamp 1632251427
transform 1 0 56830 0 1 612
box 0 0 5718 2174
use sky130_hilas_VinjDiodeProtect01  sky130_hilas_VinjDiodeProtect01_8
timestamp 1632251427
transform 1 0 62548 0 1 612
box 0 0 5718 2174
<< labels >>
rlabel metal1 62602 2328 63380 2488 0 ANALOG00
port 1 nsew
rlabel metal1 56882 2328 57660 2488 0 ANALOG01
port 2 nsew
rlabel metal1 51164 2328 51942 2488 0 ANALOG02
port 3 nsew
rlabel metal1 45448 2328 46226 2488 0 ANALOG03
port 4 nsew
rlabel metal1 39730 2328 40508 2488 0 ANALOG04
port 5 nsew
rlabel metal1 34010 2328 34788 2488 0 ANALOG05
port 6 nsew
rlabel metal1 28292 2328 29070 2488 0 ANALOG06
port 7 nsew
rlabel metal1 19868 2332 20646 2492 0 ANALOG07
port 8 nsew
rlabel metal1 11488 2328 12266 2488 0 ANALOG08
port 9 nsew
rlabel metal1 5770 2328 6548 2488 0 ANALOG09
port 10 nsew
rlabel metal1 52 2328 830 2488 0 ANALOG10
port 11 nsew
rlabel metal1 63564 0 64354 154 0 PIN1
port 12 nsew
rlabel metal1 57846 0 58636 154 0 PIN2
port 13 nsew
rlabel metal1 52130 0 52920 154 0 PIN3
port 14 nsew
rlabel metal1 46410 0 47200 154 0 PIN4
port 15 nsew
rlabel metal1 40692 0 41482 154 0 PIN5
port 16 nsew
rlabel metal1 34974 0 35764 154 0 PIN6
port 17 nsew
rlabel metal1 29256 2 30046 156 0 PIN7
port 18 nsew
rlabel metal1 12452 0 13242 154 0 PIN8
port 19 nsew
rlabel metal1 6736 0 7526 154 0 PIN9
port 20 nsew
rlabel metal1 1016 0 1806 154 0 PIN10
port 21 nsew
rlabel metal1 21006 0 21502 154 0 VTUN
port 22 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
