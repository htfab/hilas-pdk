magic
tech sky130A
timestamp 1607953977
<< nwell >>
rect -251 -181 96 -29
<< nmos >>
rect 320 -94 360 -64
rect 177 -157 217 -126
rect 320 -157 360 -126
<< pmos >>
rect -138 -96 -98 -64
rect -138 -157 -98 -126
rect 9 -157 49 -126
<< ndiff >>
rect 291 -70 320 -64
rect 291 -87 296 -70
rect 313 -87 320 -70
rect 291 -94 320 -87
rect 360 -70 391 -64
rect 360 -87 367 -70
rect 384 -87 391 -70
rect 360 -94 391 -87
rect 145 -134 177 -126
rect 145 -151 151 -134
rect 168 -151 177 -134
rect 145 -157 177 -151
rect 217 -134 249 -126
rect 217 -151 225 -134
rect 242 -151 249 -134
rect 217 -157 249 -151
rect 291 -133 320 -126
rect 291 -150 297 -133
rect 314 -150 320 -133
rect 291 -157 320 -150
rect 360 -133 390 -126
rect 360 -150 366 -133
rect 383 -150 390 -133
rect 360 -157 390 -150
<< pdiff >>
rect -167 -71 -138 -64
rect -167 -88 -161 -71
rect -144 -88 -138 -71
rect -167 -96 -138 -88
rect -98 -71 -70 -64
rect -98 -88 -92 -71
rect -75 -88 -70 -71
rect -98 -96 -70 -88
rect -168 -134 -138 -126
rect -168 -151 -161 -134
rect -144 -151 -138 -134
rect -168 -157 -138 -151
rect -98 -134 -71 -126
rect -98 -151 -92 -134
rect -75 -151 -71 -134
rect -98 -157 -71 -151
rect -20 -133 9 -126
rect -20 -150 -14 -133
rect 3 -150 9 -133
rect -20 -157 9 -150
rect 49 -133 78 -126
rect 49 -150 55 -133
rect 72 -150 78 -133
rect 49 -157 78 -150
<< ndiffc >>
rect 296 -87 313 -70
rect 367 -87 384 -70
rect 151 -151 168 -134
rect 225 -151 242 -134
rect 297 -150 314 -133
rect 366 -150 383 -133
<< pdiffc >>
rect -161 -88 -144 -71
rect -92 -88 -75 -71
rect -161 -151 -144 -134
rect -92 -151 -75 -134
rect -14 -150 3 -133
rect 55 -150 72 -133
<< psubdiff >>
rect 417 -134 440 -122
rect 417 -151 420 -134
rect 437 -151 440 -134
rect 417 -163 440 -151
<< nsubdiff >>
rect -227 -130 -195 -117
rect -227 -147 -220 -130
rect -203 -147 -195 -130
rect -227 -159 -195 -147
<< psubdiffcont >>
rect 420 -151 437 -134
<< nsubdiffcont >>
rect -220 -147 -203 -130
<< poly >>
rect -234 -56 360 -40
rect -138 -64 -98 -56
rect 320 -64 360 -56
rect -52 -83 -19 -77
rect -138 -126 -98 -96
rect -52 -100 -44 -83
rect -27 -100 -19 -83
rect -52 -103 -19 -100
rect -52 -118 217 -103
rect 9 -126 49 -118
rect 177 -126 217 -118
rect 320 -126 360 -94
rect -138 -170 -98 -157
rect 9 -170 49 -157
rect 177 -170 217 -157
rect 320 -170 360 -157
<< polycont >>
rect -44 -100 -27 -83
<< locali >>
rect -101 -71 296 -70
rect -171 -83 -161 -71
rect -188 -88 -161 -83
rect -144 -88 -136 -71
rect -101 -88 -92 -71
rect -75 -83 296 -71
rect -75 -88 -44 -83
rect -188 -96 -169 -88
rect -190 -99 -169 -96
rect -191 -100 -169 -99
rect -52 -100 -44 -88
rect -27 -87 296 -83
rect 313 -87 321 -70
rect 359 -87 367 -70
rect 384 -87 394 -70
rect -27 -88 321 -87
rect -27 -100 -19 -88
rect 412 -91 437 -71
rect -203 -105 -169 -100
rect -216 -108 -169 -105
rect -220 -111 -169 -108
rect -220 -117 -171 -111
rect -220 -122 -186 -117
rect -220 -124 -194 -122
rect -92 -124 -76 -110
rect -220 -126 -197 -124
rect -220 -130 -199 -126
rect -152 -134 -134 -130
rect -220 -158 -203 -147
rect -169 -151 -161 -134
rect -144 -151 -134 -134
rect -92 -134 -75 -124
rect -92 -159 -75 -151
rect -14 -133 3 -125
rect -14 -155 3 -150
rect 55 -133 72 -124
rect 55 -159 72 -150
rect 151 -134 168 -129
rect 151 -159 168 -151
rect 225 -134 242 -122
rect 225 -160 242 -151
rect 297 -133 314 -125
rect 363 -150 366 -133
rect 383 -150 392 -133
rect 420 -134 437 -91
rect 297 -155 314 -150
rect 420 -159 437 -151
<< metal1 >>
rect -189 -181 -169 -29
rect -91 -107 -74 -80
rect 54 -105 71 -78
rect 226 -108 243 -74
rect 346 -128 365 -53
rect 394 -181 413 -29
<< metal2 >>
rect -263 -72 -202 -52
rect -93 -72 445 -52
rect -263 -122 174 -102
rect -263 -170 314 -150
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1607949437
transform 1 0 -225 0 1 -62
box -9 -10 23 22
use sky130_hilas_li2m1  sky130_hilas_li2m1_2
timestamp 1607179295
transform 1 0 -180 0 1 -86
box -10 -8 13 21
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1607089160
transform 1 0 -139 0 1 -119
box -14 -15 20 18
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1607179295
transform 1 0 -83 0 1 -127
box -10 -8 13 21
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1607949437
transform 1 0 -86 0 1 -70
box -9 -10 23 22
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1607089160
transform 1 0 -4 0 1 -156
box -14 -15 20 18
use sky130_hilas_li2m1  sky130_hilas_li2m1_3
timestamp 1607179295
transform 1 0 62 0 1 -125
box -10 -8 13 21
use sky130_hilas_m12m2  sky130_hilas_m12m2_2
timestamp 1607949437
transform 1 0 56 0 1 -69
box -9 -10 23 22
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1607089160
transform 1 0 153 0 1 -119
box -14 -15 20 18
use sky130_hilas_li2m1  sky130_hilas_li2m1_4
timestamp 1607179295
transform 1 0 233 0 1 -126
box -10 -8 13 21
use sky130_hilas_m12m2  sky130_hilas_m12m2_4
timestamp 1607949437
transform 1 0 231 0 1 -67
box -9 -10 23 22
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1607089160
transform 1 0 304 0 1 -155
box -14 -15 20 18
use sky130_hilas_li2m1  sky130_hilas_li2m1_5
timestamp 1607179295
transform 1 0 356 0 1 -148
box -10 -8 13 21
use sky130_hilas_m12m2  sky130_hilas_m12m2_3
timestamp 1607949437
transform 1 0 335 0 1 -68
box -9 -10 23 22
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1607179295
transform 1 0 402 0 1 -86
box -10 -8 13 21
use sky130_hilas_poly2m1  sky130_hilas_poly2m1_0
timestamp 1607270135
transform 1 0 -236 0 1 -65
box -9 -26 24 25
<< labels >>
rlabel metal2 439 -72 445 -52 0 output
<< end >>
