magic
tech sky130A
timestamp 1629137257
<< checkpaint >>
rect -494 2157 939 2162
rect -494 1984 1058 2157
rect -894 1803 1058 1984
rect -894 1362 1350 1803
rect -894 1278 1614 1362
rect -894 1247 1964 1278
rect -894 538 3058 1247
rect -630 97 3058 538
rect -230 -189 3058 97
rect -161 -194 3058 -189
rect 98 -547 3058 -194
rect 98 -565 1640 -547
rect 98 -630 1614 -565
<< error_s >>
rect 1084 657 1134 663
rect 1156 657 1206 663
rect 1084 615 1134 621
rect 1156 615 1206 621
rect 1156 588 1206 594
rect 1156 546 1206 552
rect 1156 505 1206 511
rect 1156 463 1206 469
rect 1084 436 1134 442
rect 1156 436 1206 442
rect 1084 394 1134 400
rect 1156 394 1206 400
rect 1084 333 1134 339
rect 1156 333 1206 339
rect 1084 291 1134 297
rect 1156 291 1206 297
rect 1156 264 1206 270
rect 1156 222 1206 228
rect 1156 180 1206 186
rect 1156 138 1206 144
rect 1084 111 1134 117
rect 1156 111 1206 117
rect 1084 69 1134 75
rect 1156 69 1206 75
<< nwell >>
rect 977 663 1273 664
rect 977 648 1018 663
rect 1546 654 1584 664
rect 1949 650 1989 664
rect 977 647 1036 648
rect 977 471 1018 647
rect 966 429 1018 471
rect 966 409 1017 429
rect 966 356 1018 409
rect 977 60 1018 356
<< poly >>
rect 2287 618 2307 664
rect 2287 59 2307 84
<< locali >>
rect 963 77 981 169
<< metal1 >>
rect 1053 657 1069 664
rect 1094 657 1113 664
rect 1134 657 1150 664
rect 1546 654 1584 664
rect 1949 636 1989 664
rect 2209 618 2232 664
rect 2335 618 2358 664
rect 1296 532 1317 606
rect 966 356 987 471
rect 1294 195 1310 345
rect 2335 229 2358 234
rect 2331 228 2359 229
rect 2331 226 2361 228
rect 2331 199 2332 226
rect 2359 199 2361 226
rect 2331 196 2361 199
rect 1546 59 1584 69
rect 2209 59 2232 84
rect 2335 59 2358 84
<< via1 >>
rect 2332 199 2359 226
<< metal2 >>
rect 962 617 1035 635
rect 1320 614 2085 633
rect 1320 612 2102 614
rect 2064 593 2102 612
rect 2013 592 2027 593
rect 966 529 981 571
rect 2013 559 2028 592
rect 2013 539 2134 559
rect 966 520 1293 529
rect 2248 528 2374 544
rect 966 514 1309 520
rect 1279 504 1309 514
rect 964 454 996 481
rect 2024 473 2144 483
rect 2023 465 2144 473
rect 2116 453 2144 465
rect 2116 451 2119 453
rect 959 422 1017 440
rect 2248 435 2374 451
rect 1287 406 1310 407
rect 1287 403 2044 406
rect 1287 386 2050 403
rect 1287 376 1311 386
rect 966 358 1311 376
rect 2031 366 2102 386
rect 966 356 1303 358
rect 1301 336 2046 338
rect 1301 316 2102 336
rect 1301 315 1333 316
rect 962 293 1017 311
rect 960 220 980 270
rect 2022 254 2122 270
rect 2248 251 2374 267
rect 2329 226 2362 227
rect 960 200 1315 220
rect 2329 218 2332 226
rect 1694 201 2332 218
rect 2329 199 2332 201
rect 2359 199 2362 226
rect 2329 198 2362 199
rect 959 149 987 176
rect 2023 156 2123 173
rect 2250 158 2374 174
rect 2023 155 2117 156
rect 960 97 1017 115
rect 2046 110 2101 111
rect 1288 88 2101 110
rect 1288 87 2047 88
rect 1288 86 1365 87
rect 964 69 998 82
rect 1288 69 1312 86
rect 964 61 1312 69
rect 975 45 1312 61
use sky130_hilas_m12m2  sky130_hilas_m12m2_5
timestamp 1629137154
transform 1 0 1287 0 1 205
box 0 0 32 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_1
timestamp 1629137154
transform 1 0 971 0 1 360
box 0 0 32 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_3
timestamp 1629137154
transform 1 0 973 0 1 461
box 0 0 32 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_2
timestamp 1629137154
transform 1 0 1300 0 1 511
box 0 0 32 32
use sky130_hilas_m12m2  sky130_hilas_m12m2_4
timestamp 1629137154
transform 1 0 1300 0 1 323
box 0 0 32 32
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1629137146
transform 1 0 976 0 1 65
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1629137146
transform 1 0 971 0 1 161
box 0 0 34 33
use sky130_hilas_WTA4stage01  sky130_hilas_WTA4stage01_0
timestamp 1629137209
transform 1 0 2145 0 1 83
box 0 0 283 534
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1629137154
transform 1 0 1302 0 1 616
box 0 0 32 32
use sky130_hilas_swc4x1BiasCell  sky130_hilas_swc4x1BiasCell_0
timestamp 1629137241
transform -1 0 1761 0 1 441
box 0 0 2025 1091
<< labels >>
rlabel metal2 2367 528 2374 544 0 OUTPUT1
port 4 nsew analog default
rlabel metal2 2369 435 2374 451 0 OUTPUT2
port 5 nsew analog default
rlabel metal2 2369 251 2374 267 0 OUTPUT3
port 6 nsew analog default
rlabel metal2 2369 158 2374 174 0 OUTPUT4
port 7 nsew analog default
rlabel metal1 2335 658 2358 664 0 VGND
port 1 nsew ground default
rlabel metal1 2335 59 2358 65 0 VGND
port 1 nsew ground default
rlabel metal2 966 551 981 571 0 INPUT1
port 8 nsew analog default
rlabel metal2 966 454 992 480 0 INPUT2
port 9 nsew analog default
rlabel metal2 960 253 980 270 0 INPUT3
port 10 nsew analog default
rlabel metal2 959 149 987 176 0 INPUT4
port 11 nsew analog default
rlabel metal1 1547 654 1583 664 0 GATE1
port 16 nsew
rlabel metal1 1949 650 1989 664 0 VTUN
port 17 nsew
rlabel metal1 2209 59 2232 65 0 WTAMIDDLENODE
port 18 nsew
rlabel metal1 2209 658 2232 664 0 WTAMIDDLENODE
port 18 nsew
rlabel metal1 1094 657 1113 664 0 COLSEL1
port 19 nsew
rlabel metal1 1053 657 1069 664 0 VINJ
port 21 nsew
rlabel metal1 1134 657 1150 664 0 VPWR
port 20 nsew
rlabel metal2 962 617 971 635 0 DRAIN1
port 12 nsew
rlabel metal2 959 422 968 440 0 DRAIN2
port 22 nsew
rlabel metal2 962 293 971 311 0 DRAIN3
port 23 nsew
rlabel metal2 960 97 969 115 0 DRAIN4
port 24 nsew
<< end >>
