magic
tech sky130A
magscale 1 2
timestamp 1632256352
<< error_s >>
rect 116 1196 166 1224
rect 714 1196 760 1224
rect 984 1200 1022 1228
rect 634 1096 734 1106
rect 914 1096 1014 1108
rect 1274 1096 1374 1106
rect 0 914 464 1080
rect 1144 1024 1156 1038
rect 634 1012 734 1022
rect 914 1012 1014 1024
rect 1274 1012 1374 1022
rect 734 962 784 1002
rect 1224 962 1274 1002
rect 734 952 794 962
rect 779 946 794 952
rect 1218 952 1274 962
rect 1374 962 1424 1002
rect 1514 968 1520 970
rect 1374 952 1430 962
rect 1218 946 1233 952
rect 1415 948 1430 952
rect 1415 946 1444 948
rect 508 918 542 946
rect 588 916 622 944
rect 728 914 1278 946
rect 1370 914 1444 946
rect 1514 946 1538 968
rect 1486 936 1506 942
rect 1464 930 1506 936
rect 1514 934 1550 946
rect 116 912 166 914
rect 508 880 542 908
rect 728 880 1278 912
rect 1370 880 1444 912
rect 1464 896 1478 930
rect 1482 896 1506 930
rect 1512 920 1580 934
rect 1516 906 1550 920
rect 1464 890 1506 896
rect 1512 892 1580 906
rect 1486 884 1506 890
rect 779 874 794 880
rect 734 864 794 874
rect 1218 874 1233 880
rect 1415 878 1444 880
rect 1514 880 1550 892
rect 1415 874 1430 878
rect 1218 864 1274 874
rect 734 824 784 864
rect 1224 824 1274 864
rect 1374 864 1430 874
rect 1374 824 1424 864
rect 1514 858 1538 880
rect 1514 856 1520 858
rect 634 804 734 814
rect 914 802 1014 814
rect 1274 804 1374 814
rect 464 664 1148 776
rect 1274 720 1374 730
rect 634 456 734 466
rect 914 456 1014 468
rect 1274 456 1374 466
rect 0 274 464 438
rect 1144 384 1156 398
rect 634 372 734 382
rect 914 372 1014 384
rect 1274 372 1374 382
rect 734 322 784 362
rect 1224 322 1274 362
rect 734 312 794 322
rect 779 306 794 312
rect 1218 312 1274 322
rect 1374 322 1424 362
rect 1514 328 1520 330
rect 1374 312 1430 322
rect 1218 306 1233 312
rect 1415 308 1430 312
rect 1415 306 1444 308
rect 508 278 542 306
rect 588 276 622 304
rect 728 274 1278 306
rect 1370 274 1444 306
rect 1514 306 1538 328
rect 1486 296 1506 302
rect 1464 290 1506 296
rect 1514 294 1550 306
rect 116 272 166 274
rect 508 240 542 268
rect 728 240 1278 272
rect 1370 240 1444 272
rect 1464 256 1478 290
rect 1482 256 1506 290
rect 1512 280 1580 294
rect 1516 266 1550 280
rect 1464 250 1506 256
rect 1512 252 1580 266
rect 1486 244 1506 250
rect 779 234 794 240
rect 734 224 794 234
rect 1218 234 1233 240
rect 1415 238 1444 240
rect 1514 240 1550 252
rect 1415 234 1430 238
rect 1218 224 1274 234
rect 734 184 784 224
rect 1224 184 1274 224
rect 1374 224 1430 234
rect 1374 184 1424 224
rect 1514 218 1538 240
rect 1514 216 1520 218
rect 634 164 734 174
rect 914 162 1014 174
rect 1274 164 1374 174
rect 1144 148 1154 162
rect 634 80 734 90
rect 914 78 1014 90
rect 1274 80 1374 90
rect 714 0 760 28
rect 984 0 1022 28
<< nwell >>
rect 0 912 684 914
rect 0 270 684 274
<< metal1 >>
rect 116 1196 166 1210
rect 714 1196 760 1210
rect 984 1200 1022 1210
rect 116 912 166 914
rect 116 272 166 274
rect 714 0 760 16
rect 984 0 1022 14
<< metal2 >>
rect 0 1124 356 1160
rect 1128 1024 1144 1070
rect 1114 756 1144 804
rect 0 664 356 696
rect 0 506 114 508
rect 0 504 254 506
rect 0 472 400 504
rect 1128 384 1144 430
rect 1126 116 1144 162
rect 0 20 356 54
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_3
timestamp 1632255311
transform 1 0 464 0 -1 522
box 0 0 1136 340
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_2
timestamp 1632255311
transform 1 0 464 0 1 24
box 0 0 1136 340
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_0
timestamp 1632255311
transform 1 0 464 0 1 664
box 0 0 1136 340
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_1
timestamp 1632255311
transform 1 0 464 0 -1 1162
box 0 0 1136 340
<< labels >>
rlabel space 114 702 124 738 0 DRAIN2
port 3 nsew analog default
rlabel metal2 114 472 124 506 0 DRAIN3
port 2 nsew
rlabel metal1 116 1196 166 1210 0 VINJ
port 9 nsew power default
rlabel metal1 714 1196 760 1210 0 DRAIN_MUX
port 10 nsew analog default
rlabel metal1 714 0 760 16 0 DRAIN_MUX
port 10 nsew analog default
rlabel metal1 984 0 1022 14 0 VGND
port 11 nsew ground default
rlabel metal1 984 1200 1022 1210 0 VGND
port 11 nsew ground default
rlabel metal2 1122 758 1144 804 0 SELECT2
port 14 nsew
rlabel metal2 1128 1024 1144 1070 0 SELECT1
port 15 nsew
rlabel metal2 1128 384 1144 430 0 SELECT3
port 16 nsew
rlabel metal2 1126 116 1144 162 0 SELECT4
port 17 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
