magic
tech sky130A
magscale 1 2
timestamp 1632255311
<< error_s >>
rect 344648 705190 344654 705268
rect 344732 705190 344738 705268
rect 344648 704868 344654 704946
rect 344732 704868 344738 704946
rect 344800 704744 345032 705360
rect 345218 705334 345235 705356
rect 345162 705330 345282 705334
rect 345180 705306 345182 705310
rect 345187 705306 345188 705318
rect 345202 705316 345266 705330
rect 345214 705306 345216 705316
rect 345162 705302 345254 705306
rect 345174 705288 345254 705302
rect 345180 705276 345182 705288
rect 345214 705286 345216 705288
rect 345104 705186 345110 705264
rect 345188 705186 345194 705264
rect 345296 705186 345302 705264
rect 345380 705186 345386 705264
rect 345488 705186 345494 705264
rect 345572 705186 345578 705264
rect 345680 705190 345686 705268
rect 345764 705190 345770 705268
rect 345064 705086 345136 705088
rect 345256 705086 345328 705088
rect 345448 705086 345520 705088
rect 345286 704962 345292 704988
rect 345302 704947 345307 704998
rect 345329 704988 345380 704998
rect 345329 704983 345410 704988
rect 345344 704970 345410 704983
rect 345448 704970 345452 705016
rect 345365 704955 345380 704970
rect 345104 704868 345110 704946
rect 345188 704868 345194 704946
rect 345296 704868 345302 704946
rect 345380 704868 345386 704946
rect 345488 704868 345494 704946
rect 345572 704868 345578 704946
rect 345680 704868 345686 704946
rect 345764 704868 345770 704946
rect 346846 664368 346862 666626
rect 346846 647396 346862 649654
<< metal1 >>
rect 273822 671750 274334 678558
rect 279428 671750 279938 683058
rect 285320 671750 285830 686874
rect 293792 671872 294186 691516
rect 302118 671750 302630 696050
rect 307716 671750 308228 700830
rect 313560 671750 314072 699328
rect 319278 671750 319790 694214
rect 324994 671750 325506 688542
rect 330552 671750 331062 684306
rect 336286 671750 336796 679802
rect 267744 665632 269422 665834
rect 267576 665102 269422 665632
rect 342952 665468 345336 665692
rect 342952 664958 345412 665468
rect 267844 659912 269422 660118
rect 267644 659384 269422 659912
rect 342952 659466 345412 659974
rect 342952 659270 345374 659466
rect 268112 654196 269422 654398
rect 267978 653666 269422 654196
rect 342952 654030 345026 654254
rect 342952 653522 346866 654030
rect 268080 648474 269422 648680
rect 267780 647948 269422 648474
rect 342952 648314 345432 648538
rect 342952 647804 345452 648314
rect 267676 642758 269422 642964
rect 267610 642230 269422 642758
rect 342952 642592 345372 642820
rect 342952 642086 346340 642592
rect 268078 637042 269422 637244
rect 267676 636512 269422 637042
rect 342952 636508 345684 637018
rect 342952 636368 345044 636508
rect 267778 630794 269422 631528
rect 342952 631160 344890 631382
rect 342952 630650 346002 631160
rect 267748 625614 269422 625810
rect 267614 625092 269422 625614
rect 340900 624628 341206 624772
rect 267310 619564 269422 620090
rect 267344 619358 269422 619564
rect 267442 613844 269422 614372
rect 267644 613640 269422 613844
rect 267676 608450 269422 608654
rect 267644 607922 269422 608450
<< metal2 >>
rect 265596 671712 266364 671730
rect 265596 670846 265610 671712
rect 266342 671378 266364 671712
rect 362332 671492 364770 671532
rect 362332 671396 362360 671492
rect 266342 670920 270008 671378
rect 342396 670964 362360 671396
rect 266342 670846 266364 670920
rect 265596 670828 266364 670846
rect 362332 670840 362360 670964
rect 364738 671396 364770 671492
rect 364738 670964 364774 671396
rect 364738 670840 364770 670964
rect 362332 670822 364770 670840
rect 270814 670358 271780 670478
rect 270814 669574 270904 670358
rect 271688 669574 271780 670358
rect 341090 670266 341842 670320
rect 341090 669752 341126 670266
rect 341792 669752 341842 670266
rect 341090 669718 341842 669752
rect 270814 669482 271780 669574
rect 339006 634310 341334 634660
rect 342376 628672 349778 628948
rect 340806 626698 392052 627292
rect 391400 623756 392052 626698
rect 389018 623746 394436 623756
rect 389018 618318 394436 618328
rect 268260 594512 270002 594792
rect 270982 593210 271262 594726
rect 290870 46538 291562 46554
rect 290870 46536 291028 46538
rect 125674 46024 291028 46536
rect 291542 46024 291562 46538
rect 125674 2884 126186 46024
rect 290870 46012 291562 46024
rect 297290 45500 297694 595892
rect 126984 45008 297694 45500
rect 126984 44988 297630 45008
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 2884
rect 126998 -800 127110 44988
rect 290914 44464 291550 44486
rect 290914 44462 290996 44464
rect 128918 43950 290996 44462
rect 291510 43950 291550 44464
rect 128918 3422 129430 43950
rect 290914 43932 291550 43950
rect 298102 43386 298506 595892
rect 130542 42874 298506 43386
rect 128918 2968 129474 3422
rect 128180 -800 128292 480
rect 129362 -800 129474 2968
rect 130544 -800 130656 42874
rect 298102 42836 298506 42874
rect 291014 42312 291704 42342
rect 291014 42310 291124 42312
rect 132422 41798 291124 42310
rect 291638 41798 291704 42312
rect 132422 2900 132934 41798
rect 291014 41782 291704 41798
rect 298896 41292 299300 595892
rect 134064 40796 299300 41292
rect 134064 40780 299276 40796
rect 132422 2468 133020 2900
rect 131726 -800 131838 480
rect 132908 -800 133020 2468
rect 134090 -800 134202 40780
rect 291072 40276 291718 40298
rect 291072 40274 291156 40276
rect 136410 39762 291156 40274
rect 291670 39762 291718 40276
rect 136410 39542 136918 39762
rect 291072 39746 291718 39762
rect 136406 2802 136918 39542
rect 299696 39208 300100 595892
rect 137622 38698 300100 39208
rect 137622 38696 299446 38698
rect 135272 -800 135384 480
rect 136454 -800 136566 2802
rect 137636 -800 137748 38696
rect 300506 32884 300910 595892
rect 141182 32430 300916 32884
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 32430
rect 301308 31980 301712 595892
rect 144714 31590 301712 31980
rect 144714 31530 301684 31590
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 31530
rect 302108 31256 302512 595892
rect 148274 31078 148386 31088
rect 302108 31078 302502 31256
rect 148274 30628 302502 31078
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 30628
rect 302926 30174 303330 595892
rect 151844 30164 303332 30174
rect 151820 29724 303332 30164
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 29724
rect 155366 29320 155478 29332
rect 303752 29320 304156 595892
rect 155366 28882 304156 29320
rect 155366 28870 303334 28882
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 28870
rect 304552 28418 304956 595892
rect 158898 27968 304982 28418
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 27968
rect 305344 27530 305748 595892
rect 162410 27080 305758 27530
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 27080
rect 305344 27032 305748 27080
rect 306154 26628 306558 595892
rect 166026 26622 306558 26628
rect 166004 26192 306558 26622
rect 166004 26178 306176 26192
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 26178
rect 169550 25724 169662 25730
rect 306972 25724 307376 595892
rect 307774 26424 308178 595892
rect 169550 25320 307376 25724
rect 169550 25274 307340 25320
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 25274
rect 307730 24804 308180 26424
rect 173088 24354 308180 24804
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 24354
rect 308582 23918 308986 595892
rect 176618 23476 308986 23918
rect 176618 23468 308892 23476
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 23468
rect 180188 23038 180300 23052
rect 309400 23038 309804 595892
rect 180168 22634 309804 23038
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 22634
rect 310210 22164 310614 595892
rect 183732 21760 310614 22164
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 21760
rect 311004 21438 311408 595892
rect 187244 21034 311408 21438
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 21034
rect 311828 20310 312232 595892
rect 190726 19906 312232 20310
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 19906
rect 312654 19292 313058 595890
rect 194400 19248 313058 19292
rect 194372 18888 313058 19248
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 18888
rect 313456 18238 313860 595892
rect 197954 18206 313860 18238
rect 197918 17834 313860 18206
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 17834
rect 201464 17218 201576 17226
rect 314258 17218 314662 595896
rect 201384 16814 314662 17218
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 16814
rect 315076 16346 315480 595892
rect 205030 16338 315480 16346
rect 205010 15942 315480 16338
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 15942
rect 315910 15400 316314 595892
rect 208584 15358 316314 15400
rect 208556 14996 316314 15358
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 14996
rect 212102 14504 212214 14552
rect 316710 14504 317114 595892
rect 317512 46524 317916 595892
rect 317446 46508 317978 46524
rect 317446 45994 317458 46508
rect 317972 45994 317978 46508
rect 317446 45982 317978 45994
rect 318304 44540 318708 595892
rect 318230 44530 318772 44540
rect 318230 44016 318250 44530
rect 318764 44016 318772 44530
rect 318230 44000 318772 44016
rect 319114 42368 319518 595892
rect 319042 42346 319580 42368
rect 319042 41832 319060 42346
rect 319574 41832 319580 42346
rect 319042 41824 319580 41832
rect 319060 41822 319574 41824
rect 319926 40324 320330 595892
rect 319856 40312 320396 40324
rect 319856 39798 319872 40312
rect 320386 39798 320396 40312
rect 319856 39788 320396 39798
rect 212062 14100 317114 14504
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 14100
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 265610 670846 266342 671712
rect 362360 670840 364738 671492
rect 270904 669574 271688 670358
rect 341126 669752 341792 670266
rect 389018 618328 394436 623746
rect 291028 46024 291542 46538
rect 290996 43950 291510 44464
rect 291124 41798 291638 42312
rect 291156 39762 291670 40276
rect 317458 45994 317972 46508
rect 318250 44016 318764 44530
rect 319060 41832 319574 42346
rect 319872 39798 320386 40312
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 703360 515394 704800
rect 520594 703360 525394 704800
rect 510594 702340 525394 703360
rect -800 683324 1700 685242
rect 18694 683324 21194 702300
rect 69238 687864 71738 702300
rect 122694 692542 125194 702300
rect 177022 698308 179522 702300
rect 229456 701902 231956 702300
rect 229456 699890 308786 701902
rect 320238 700048 322738 702300
rect 229564 699182 308786 699890
rect 177086 697114 179522 698308
rect 312730 697548 322738 700048
rect 177086 694394 303300 697114
rect 177086 694388 179522 694394
rect 414284 694110 416784 702300
rect 122600 689822 294718 692542
rect 318894 691638 416854 694110
rect 414284 691594 416784 691638
rect 466978 689538 469478 702300
rect 510596 701862 525388 702340
rect 566594 702300 571594 704800
rect 510596 692380 510888 701862
rect 525094 692380 525388 701862
rect 510596 692022 525388 692380
rect 69202 685144 286134 687864
rect 324758 687066 469738 689538
rect 568570 686634 571070 702300
rect 69238 685092 71738 685144
rect 568570 685088 570954 686634
rect -800 680824 9186 683324
rect 18672 680824 280532 683324
rect 330356 682616 570954 685088
rect 568570 682548 570954 682616
rect -800 680242 1700 680824
rect 6686 678864 9186 680824
rect 582300 680744 584800 682984
rect 6686 676392 275108 678864
rect 335804 678244 584800 680744
rect 582300 677984 584800 678244
rect 6922 676364 275108 676392
rect 264680 671744 266066 671746
rect 264680 671742 266380 671744
rect 228350 671712 266380 671742
rect 228350 671598 265610 671712
rect 228350 670910 228514 671598
rect 238740 670910 265610 671598
rect 228350 670846 265610 670910
rect 266342 670846 266380 671712
rect 228350 670812 266380 670846
rect 264994 670810 266380 670812
rect 362302 671492 382720 671588
rect 362302 670840 362360 671492
rect 364738 671336 382720 671492
rect 364738 670932 372006 671336
rect 382670 670932 382720 671336
rect 364738 670840 382720 670932
rect 362302 670780 382720 670840
rect 247894 670358 271750 670418
rect 247894 670298 270904 670358
rect 247894 669574 248104 670298
rect 254890 669574 270904 670298
rect 271688 669574 271750 670358
rect 341102 670266 360940 670296
rect 341102 669752 341126 670266
rect 341792 670202 360940 670266
rect 341792 669810 353734 670202
rect 360836 669810 360940 670202
rect 341792 669752 360940 669810
rect 341102 669734 360940 669752
rect 247894 669512 271750 669574
rect 6514 666814 8378 666828
rect 265400 666814 266130 667122
rect 6514 665212 267320 666814
rect -800 648638 1660 648642
rect -800 648300 4986 648638
rect -800 643842 1900 648300
rect 308 638642 1900 643842
rect -800 634132 1900 638642
rect 4680 634132 4986 648300
rect -800 633842 4986 634132
rect 308 633826 4986 633842
rect 286 564242 4696 564244
rect -800 564010 4696 564242
rect -800 559442 1890 564010
rect 286 554242 1890 559442
rect -800 549544 1890 554242
rect 4462 549544 4696 564010
rect -800 549442 4696 549544
rect 286 549412 4696 549442
rect 6514 511642 7976 665212
rect 344282 664640 574078 666160
rect -800 511532 7976 511642
rect 9546 660890 11082 660896
rect 9546 659288 267994 660890
rect 344282 660132 569392 660202
rect -800 511530 7960 511532
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 9546 468420 11082 659288
rect 344282 658682 570578 660132
rect 565534 655162 567136 655168
rect 12736 654544 14226 654564
rect 12736 652942 267740 654544
rect 344282 653642 567174 655162
rect 12736 652060 14226 652942
rect 12690 651470 14226 652060
rect -800 468308 11082 468420
rect 9546 468004 11082 468308
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 12736 425198 14226 651470
rect 15794 648644 268754 649216
rect 562172 648974 563774 649002
rect -800 425086 14226 425198
rect 12736 425064 14226 425086
rect 15762 647614 268754 648644
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 15762 381976 17318 647614
rect 344282 647454 563774 648974
rect 18982 643540 267994 643886
rect -800 381864 17318 381976
rect 15762 381650 17318 381864
rect 18832 642284 267994 643540
rect 558808 643474 560568 643478
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 18832 338754 20388 642284
rect 344512 641954 560568 643474
rect 22172 638278 268502 638304
rect -800 338642 20388 338754
rect 18832 338352 20388 338642
rect 21980 636702 268502 638278
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 21980 295532 23536 636702
rect 344282 636226 557126 637746
rect -800 295420 23536 295532
rect 21980 295362 23536 295420
rect 25170 631960 26726 632060
rect 25170 630358 268754 631960
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 25170 252510 26726 630358
rect 28550 625842 268502 625868
rect -800 252398 26726 252510
rect 25170 252350 26726 252398
rect 28320 624266 268502 625842
rect 337636 624754 339098 633988
rect 551362 632246 553124 632268
rect 344512 630726 553284 632246
rect 350436 629168 380732 629212
rect 381948 629168 382130 629198
rect 350436 628028 372112 629168
rect 371856 627994 372112 628028
rect 382068 627994 382130 629168
rect 371856 627932 372308 627994
rect 381948 627924 382130 627994
rect 353562 624754 361356 624858
rect 337636 624690 361356 624754
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 440 219688 7624 219778
rect -800 219146 7624 219688
rect -800 214888 2280 219146
rect 440 209688 2280 214888
rect -800 205238 2280 209688
rect 6878 205238 7624 219146
rect -800 204888 7624 205238
rect 440 204836 7624 204888
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 28320 124888 29876 624266
rect 337636 623292 353706 624690
rect 353562 622968 353706 623292
rect 361190 622968 361356 624690
rect 353562 622850 361356 622968
rect 388064 624192 394798 624400
rect 388064 624006 395168 624192
rect 31738 620738 268754 620794
rect -800 124776 29876 124888
rect 28320 124288 29876 124776
rect 31548 619192 268754 620738
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 31548 81666 33104 619192
rect 388064 618114 388772 624006
rect 394718 618114 395168 624006
rect 388064 618000 395168 618114
rect 39554 615176 268248 615210
rect -800 81554 33104 81666
rect 31548 81496 33104 81554
rect 34738 613608 268248 615176
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 34738 38444 36294 613608
rect -800 38332 36294 38444
rect 34738 38266 36294 38332
rect 37926 609374 39482 609596
rect 37926 607772 268502 609374
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 37926 17022 39482 607772
rect 228100 593970 238868 594134
rect 228100 592948 228220 593970
rect 238688 593904 238868 593970
rect 238688 593322 269202 593904
rect 388064 593616 394798 618000
rect 238688 592948 238868 593322
rect 228100 592872 238868 592948
rect 247452 592130 254918 592310
rect 247452 591498 247572 592130
rect 254828 592086 254918 592130
rect 254828 591504 271232 592086
rect 254828 591498 254918 591504
rect 247452 591318 254918 591498
rect 388064 590730 394316 593616
rect 215386 589916 394316 590730
rect 215386 582968 215548 589916
rect 219722 582968 394316 589916
rect 215386 582554 394316 582968
rect 551362 313764 553124 630726
rect 555206 313764 556966 636226
rect 558808 358986 560568 641954
rect 562172 405408 563774 647454
rect 565534 449830 567136 653642
rect 568896 494252 570578 658682
rect 572558 583674 574078 664640
rect 577036 644584 583594 644604
rect 577036 643224 584800 644584
rect 577036 630452 577726 643224
rect 582732 639784 584800 643224
rect 582732 634584 583594 639784
rect 582732 630452 584800 634584
rect 577036 629784 584800 630452
rect 577036 629762 583594 629784
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 572558 583562 584800 583674
rect 572558 583498 574078 583562
rect 582340 555072 584800 555362
rect 574216 553924 584800 555072
rect 574216 541748 575594 553924
rect 581108 550562 584800 553924
rect 581108 545362 583866 550562
rect 581108 541748 584800 545362
rect 574216 540828 584800 541748
rect 582340 540562 584800 540828
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 568896 494156 584800 494252
rect 569690 494140 584800 494156
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 565534 449718 584800 449830
rect 565534 449692 567136 449718
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 562172 405296 584800 405408
rect 562172 405264 563774 405296
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 558808 358874 584800 358986
rect 558808 358848 560568 358874
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 551362 313652 553152 313764
rect 555198 313652 584800 313764
rect 551362 269342 553124 313652
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 551362 269230 584800 269342
rect 551362 268992 553124 269230
rect 582340 240016 584800 240030
rect 577670 239570 584800 240016
rect 130618 239472 584800 239570
rect 130618 238994 578096 239472
rect 130618 226310 131182 238994
rect 141256 226310 578096 238994
rect 130618 225696 578096 226310
rect 577670 225630 578096 225696
rect 581490 235230 584800 239472
rect 581490 230030 583148 235230
rect 581490 225630 584800 230030
rect 577670 225230 584800 225630
rect 577670 225198 583148 225230
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect 582340 151592 584800 151630
rect 575734 151306 584800 151592
rect 575734 137100 575938 151306
rect 581978 146830 584800 151306
rect 581978 141630 583774 146830
rect 581978 137100 584800 141630
rect 575734 136830 584800 137100
rect 575734 136814 583774 136830
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect 290850 46552 291592 46570
rect 290850 46538 317984 46552
rect 290850 46024 291028 46538
rect 291542 46508 317984 46538
rect 291542 46038 317458 46508
rect 291542 46024 291592 46038
rect 290850 45998 291592 46024
rect 317440 45994 317458 46038
rect 317972 45994 317984 46508
rect 317440 45972 317984 45994
rect 318222 44530 318778 44550
rect 290900 44464 291570 44502
rect 290900 43950 290996 44464
rect 291510 44462 291570 44464
rect 318222 44462 318250 44530
rect 291510 44016 318250 44462
rect 318764 44016 318778 44530
rect 291510 43990 318778 44016
rect 291510 43950 318754 43990
rect 290900 43948 318754 43950
rect 290900 43920 291570 43948
rect 319024 42372 319594 42386
rect 290962 42346 319594 42372
rect 290962 42312 319060 42346
rect 290962 41858 291124 42312
rect 290966 41798 291124 41858
rect 291638 41858 319060 42312
rect 291638 41798 291750 41858
rect 319024 41832 319060 41858
rect 319574 41832 319594 42346
rect 319024 41816 319594 41832
rect 290966 41770 291750 41798
rect 319846 40314 320402 40334
rect 290962 40312 320402 40314
rect 290962 40276 319872 40312
rect 290962 39800 291156 40276
rect 290966 39762 291156 39800
rect 291670 39800 319872 40276
rect 291670 39762 291740 39800
rect 319846 39798 319872 39800
rect 320386 39798 320402 40312
rect 319846 39780 320402 39798
rect 290966 39736 291740 39762
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 39482 17022
rect 583520 16910 584800 17022
rect 37926 16766 39482 16910
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 510888 692380 525094 701862
rect 228514 670910 238740 671598
rect 372006 670932 382670 671336
rect 248104 669574 254890 670298
rect 353734 669810 360836 670202
rect 1900 634132 4680 648300
rect 1890 549544 4462 564010
rect 372112 627994 382068 629168
rect 2280 205238 6878 219146
rect 353706 622968 361190 624690
rect 388772 623746 394718 624006
rect 388772 618328 389018 623746
rect 389018 618328 394436 623746
rect 394436 618328 394718 623746
rect 388772 618114 394718 618328
rect 228220 592948 238688 593970
rect 247572 591498 254828 592130
rect 215548 582968 219722 589916
rect 577726 630452 582732 643224
rect 575594 541748 581108 553924
rect 131182 226310 141256 238994
rect 578096 225630 581490 239472
rect 575938 137100 581978 151306
<< metal4 >>
rect 510336 701862 525680 701992
rect 510336 692380 510888 701862
rect 525094 692380 525680 701862
rect 510336 690882 525680 692380
rect 227932 679440 525352 690550
rect 227932 671598 239042 679440
rect 227932 670910 228514 671598
rect 238740 670910 239042 671598
rect 1800 648300 12070 648402
rect 1800 634132 1900 648300
rect 4680 642164 12070 648300
rect 4680 634774 69488 642164
rect 4680 634132 12070 634774
rect 1800 633962 12070 634132
rect 62098 590098 69488 634774
rect 227932 594014 239042 670910
rect 247292 670298 255104 670598
rect 247292 669574 248104 670298
rect 254890 669574 255104 670298
rect 227932 593970 239192 594014
rect 227932 592948 228220 593970
rect 238688 592948 239192 593970
rect 62098 589916 220042 590098
rect 62098 582968 215548 589916
rect 219722 582968 220042 589916
rect 62098 582708 220042 582968
rect 1556 564010 8972 564778
rect 1556 549544 1890 564010
rect 4462 562936 8972 564010
rect 227932 562936 239192 592948
rect 4462 551322 239192 562936
rect 247292 592130 255104 669574
rect 247292 591498 247572 592130
rect 254828 591498 255104 592130
rect 4462 549544 8972 551322
rect 1556 549144 8972 549544
rect 130684 238994 142178 240238
rect 130684 226310 131182 238994
rect 141256 226310 142178 238994
rect 1992 219146 18372 219434
rect 1992 205238 2280 219146
rect 6878 216502 18372 219146
rect 130684 216502 142178 226310
rect 6878 205238 142178 216502
rect 1992 205008 142178 205238
rect 221812 152244 232386 551322
rect 247292 550814 255104 591498
rect 353566 670202 361378 672320
rect 353566 669810 353734 670202
rect 360836 669810 361378 670202
rect 353566 624690 361378 669810
rect 371844 671336 382954 679440
rect 371844 670932 372006 671336
rect 382670 670932 382954 671336
rect 371844 630446 382954 670932
rect 570824 643224 583248 643742
rect 570824 640780 577726 643224
rect 371756 629500 382954 630446
rect 535752 633878 577726 640780
rect 371756 629382 383090 629500
rect 371668 629168 383090 629382
rect 371668 627994 372112 629168
rect 382068 627994 383090 629168
rect 371668 627638 383090 627994
rect 371756 627338 383090 627638
rect 371756 625638 382954 627338
rect 353566 622968 353706 624690
rect 361190 622968 361378 624690
rect 371844 624602 382954 625638
rect 388602 624752 390048 624774
rect 535752 624752 542654 633878
rect 570824 630452 577726 633878
rect 582732 630452 583248 643224
rect 570824 630280 583248 630452
rect 353566 550814 361378 622968
rect 388602 624006 542654 624752
rect 388602 618114 388772 624006
rect 394718 618114 542654 624006
rect 388602 617870 542654 618114
rect 388740 617850 542654 617870
rect 567782 553924 581798 554614
rect 567782 550814 575594 553924
rect 247292 543002 575594 550814
rect 518290 454198 527212 543002
rect 567782 541748 575594 543002
rect 581108 541748 581798 553924
rect 567782 540828 581798 541748
rect 516836 445276 527212 454198
rect 518290 238370 527210 445276
rect 569176 239472 582274 240414
rect 569176 238370 578096 239472
rect 518290 229450 578096 238370
rect 569176 225630 578096 229450
rect 581490 225630 582274 239472
rect 569176 224722 582274 225630
rect 221812 152162 580060 152244
rect 221812 151306 582306 152162
rect 221812 141670 575938 151306
rect 565364 137100 575938 141670
rect 581978 137100 582306 151306
rect 565364 136324 582306 137100
rect 565364 136120 580060 136324
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use m12m3  m12m3_31
timestamp 1632251359
transform 1 0 266746 0 1 593000
box 0 0 2514 2216
use m12m3  m12m3_32
timestamp 1632251359
transform 1 0 270788 0 1 591520
box 0 0 2514 2216
use m12m3  m12m3_29
timestamp 1632251359
transform 1 0 266024 0 1 607692
box 0 0 2514 2216
use m12m3  m12m3_25
timestamp 1632251359
transform 1 0 266148 0 1 630212
box 0 0 2514 2216
use m12m3  m12m3_27
timestamp 1632251359
transform 1 0 266024 0 1 619320
box 0 0 2514 2216
use m12m3  m12m3_26
timestamp 1632251359
transform 1 0 266148 0 1 624182
box 0 0 2514 2216
use m12m3  m12m3_28
timestamp 1632251359
transform 1 0 265896 0 1 613506
box 0 0 2514 2216
use m12m3  m12m3_18
timestamp 1632251359
transform 1 0 344412 0 1 630454
box 0 0 2514 2216
use m12m3  m12m3_30
timestamp 1632251359
transform 1 0 348536 0 1 627722
box 0 0 2514 2216
use m12m3  m12m3_22
timestamp 1632251359
transform 1 0 266248 0 1 647498
box 0 0 2514 2216
use m12m3  m12m3_24
timestamp 1632251359
transform 1 0 266216 0 1 636342
box 0 0 2514 2216
use m12m3  m12m3_23
timestamp 1632251359
transform 1 0 266114 0 1 642038
box 0 0 2514 2216
use m12m3  m12m3_15
timestamp 1632251359
transform 1 0 344332 0 1 647428
box 0 0 2514 2216
use m12m3  m12m3_16
timestamp 1632251359
transform 1 0 344576 0 1 641824
box 0 0 2514 2216
use m12m3  m12m3_17
timestamp 1632251359
transform 1 0 344494 0 1 635976
box 0 0 2514 2216
use m12m3  m12m3_8
timestamp 1632251359
transform 1 0 336808 0 1 633150
box 0 0 2514 2216
use m12m3  m12m3_21
timestamp 1632251359
transform 1 0 266248 0 1 652958
box 0 0 2514 2216
use m12m3  m12m3_20
timestamp 1632251359
transform 1 0 266216 0 1 659022
box 0 0 2514 2216
use m12m3  m12m3_13
timestamp 1632251359
transform 1 0 344494 0 1 658552
box 0 0 2514 2216
use m12m3  m12m3_14
timestamp 1632251359
transform 1 0 344494 0 1 653518
box 0 0 2514 2216
use m12m3  m12m3_2
timestamp 1632251359
transform 1 0 283528 0 1 685404
box 0 0 2514 2216
use m12m3  m12m3_0
timestamp 1632251359
transform 1 0 278002 0 1 681056
box 0 0 2514 2216
use m12m3  m12m3_1
timestamp 1632251359
transform 1 0 272474 0 1 676604
box 0 0 2514 2216
use m12m3  m12m3_19
timestamp 1632251359
transform 1 0 266082 0 1 664918
box 0 0 2514 2216
use m12m3  m12m3_10
timestamp 1632251359
transform 1 0 330400 0 1 682794
box 0 0 2514 2216
use m12m3  m12m3_11
timestamp 1632251359
transform 1 0 335926 0 1 678496
box 0 0 2514 2216
use m12m3  m12m3_9
timestamp 1632251359
transform 1 0 324872 0 1 687246
box 0 0 2514 2216
use m12m3  m12m3_12
timestamp 1632251359
transform 1 0 344332 0 1 664400
box 0 0 2514 2216
use m12m3  m12m3_5
timestamp 1632251359
transform 1 0 306196 0 1 699578
box 0 0 2514 2216
use m12m3  m12m3_6
timestamp 1632251359
transform 1 0 313052 0 1 697788
box 0 0 2514 2216
use m12m3  m12m3_4
timestamp 1632251359
transform 1 0 300568 0 1 694718
box 0 0 2514 2216
use m12m3  m12m3_3
timestamp 1632251359
transform 1 0 292124 0 1 690112
box 0 0 2514 2216
use m12m3  m12m3_7
timestamp 1632251359
transform 1 0 319142 0 1 691852
box 0 0 2514 2216
use sky130_hilas_TopProtectStructure  sky130_hilas_TopProtectStructure_0
timestamp 1632255311
transform 1 0 299828 0 1 643120
box 0 0 78744 93154
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 GPIO_ANALOG\[0\]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 GPIO_ANALOG\[10\]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 GPIO_ANALOG\[11\]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 GPIO_ANALOG\[12\]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 GPIO_ANALOG\[13\]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 GPIO_ANALOG\[14\]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 GPIO_ANALOG\[15\]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 GPIO_ANALOG\[16\]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 GPIO_ANALOG\[17\]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 GPIO_ANALOG\[1\]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 GPIO_ANALOG\[2\]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 GPIO_ANALOG\[3\]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 GPIO_ANALOG\[4\]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 GPIO_ANALOG\[5\]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 GPIO_ANALOG\[6\]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 GPIO_ANALOG\[7\]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 GPIO_ANALOG\[8\]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 GPIO_ANALOG\[9\]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 GPIO_NOESD\[0\]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 GPIO_NOESD\[10\]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 GPIO_NOESD\[11\]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 GPIO_NOESD\[12\]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 GPIO_NOESD\[13\]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 GPIO_NOESD\[14\]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 GPIO_NOESD\[15\]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 GPIO_NOESD\[16\]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 GPIO_NOESD\[17\]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 GPIO_NOESD\[1\]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 GPIO_NOESD\[2\]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 GPIO_NOESD\[3\]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 GPIO_NOESD\[4\]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 GPIO_NOESD\[5\]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 GPIO_NOESD\[6\]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 GPIO_NOESD\[7\]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 GPIO_NOESD\[8\]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 GPIO_NOESD\[9\]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 IO_ANALOG\[0\]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 IO_ANALOG\[10\]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 IO_ANALOG\[1\]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 IO_ANALOG\[2\]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 IO_ANALOG\[3\]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 IO_ANALOG\[4\]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 IO_ANALOG\[5\]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 IO_ANALOG\[6\]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 IO_ANALOG\[7\]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 IO_ANALOG\[8\]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 IO_ANALOG\[9\]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 IO_ANALOG\[4\]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 IO_ANALOG\[5\]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 IO_ANALOG\[6\]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 IO_CLAMP_HIGH\[0\]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 IO_CLAMP_HIGH\[1\]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 IO_CLAMP_HIGH\[2\]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 IO_CLAMP_LOW\[0\]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 IO_CLAMP_LOW\[1\]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 IO_CLAMP_LOW\[2\]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 IO_IN\[0\]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 IO_IN\[10\]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 IO_IN\[11\]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 IO_IN\[12\]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 IO_IN\[13\]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 IO_IN\[14\]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 IO_IN\[15\]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 IO_IN\[16\]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 IO_IN\[17\]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 IO_IN\[18\]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 IO_IN\[19\]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 IO_IN\[1\]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 IO_IN\[20\]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 IO_IN\[21\]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 IO_IN\[22\]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 IO_IN\[23\]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 IO_IN\[24\]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 IO_IN\[25\]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 IO_IN\[26\]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 IO_IN\[2\]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 IO_IN\[3\]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 IO_IN\[4\]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 IO_IN\[5\]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 IO_IN\[6\]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 IO_IN\[7\]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 IO_IN\[8\]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 IO_IN\[9\]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 IO_IN_3V3\[0\]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 IO_IN_3V3\[10\]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 IO_IN_3V3\[11\]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 IO_IN_3V3\[12\]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 IO_IN_3V3\[13\]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 IO_IN_3V3\[14\]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 IO_IN_3V3\[15\]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 IO_IN_3V3\[16\]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 IO_IN_3V3\[17\]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 IO_IN_3V3\[18\]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 IO_IN_3V3\[19\]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 IO_IN_3V3\[1\]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 IO_IN_3V3\[20\]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 IO_IN_3V3\[21\]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 IO_IN_3V3\[22\]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 IO_IN_3V3\[23\]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 IO_IN_3V3\[24\]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 IO_IN_3V3\[25\]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 IO_IN_3V3\[26\]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 IO_IN_3V3\[2\]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 IO_IN_3V3\[3\]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 IO_IN_3V3\[4\]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 IO_IN_3V3\[5\]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 IO_IN_3V3\[6\]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 IO_IN_3V3\[7\]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 IO_IN_3V3\[8\]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 IO_IN_3V3\[9\]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 IO_OEB\[0\]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 IO_OEB\[10\]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 IO_OEB\[11\]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 IO_OEB\[12\]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 IO_OEB\[13\]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 IO_OEB\[14\]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 IO_OEB\[15\]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 IO_OEB\[16\]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 IO_OEB\[17\]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 IO_OEB\[18\]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 IO_OEB\[19\]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 IO_OEB\[1\]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 IO_OEB\[20\]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 IO_OEB\[21\]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 IO_OEB\[22\]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 IO_OEB\[23\]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 IO_OEB\[24\]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 IO_OEB\[25\]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 IO_OEB\[26\]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 IO_OEB\[2\]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 IO_OEB\[3\]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 IO_OEB\[4\]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 IO_OEB\[5\]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 IO_OEB\[6\]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 IO_OEB\[7\]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 IO_OEB\[8\]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 IO_OEB\[9\]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 IO_OUT\[0\]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 IO_OUT\[10\]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 IO_OUT\[11\]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 IO_OUT\[12\]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 IO_OUT\[13\]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 IO_OUT\[14\]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 IO_OUT\[15\]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 IO_OUT\[16\]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 IO_OUT\[17\]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 IO_OUT\[18\]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 IO_OUT\[19\]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 IO_OUT\[1\]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 IO_OUT\[20\]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 IO_OUT\[21\]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 IO_OUT\[22\]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 IO_OUT\[23\]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 IO_OUT\[24\]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 IO_OUT\[25\]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 IO_OUT\[26\]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 IO_OUT\[2\]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 IO_OUT\[3\]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 IO_OUT\[4\]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 IO_OUT\[5\]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 IO_OUT\[6\]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 IO_OUT\[7\]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 IO_OUT\[8\]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 IO_OUT\[9\]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[0\]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[100\]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[101\]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[102\]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[103\]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[104\]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[105\]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[106\]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[107\]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[108\]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[109\]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[10\]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[110\]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[111\]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[112\]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[113\]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[114\]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[115\]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[116\]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[117\]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[118\]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[119\]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[11\]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[120\]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[121\]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[122\]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[123\]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[124\]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[125\]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[126\]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[127\]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[12\]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[13\]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[14\]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[15\]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[16\]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[17\]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[18\]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[19\]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[1\]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[20\]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[21\]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[22\]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[23\]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[24\]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[25\]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[26\]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[27\]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[28\]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[29\]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[2\]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[30\]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[31\]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[32\]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[33\]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[34\]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[35\]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[36\]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[37\]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[38\]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[39\]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[3\]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[40\]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[41\]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[42\]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[43\]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[44\]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[45\]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[46\]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[47\]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[48\]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[49\]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[4\]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[50\]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[51\]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[52\]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[53\]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[54\]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[55\]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[56\]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[57\]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[58\]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[59\]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[5\]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[60\]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[61\]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[62\]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[63\]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[64\]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[65\]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[66\]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[67\]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[68\]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[69\]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[6\]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[70\]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[71\]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[72\]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[73\]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[74\]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[75\]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[76\]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[77\]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[78\]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[79\]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[7\]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[80\]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[81\]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[82\]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[83\]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[84\]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[85\]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[86\]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[87\]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[88\]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[89\]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[8\]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[90\]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[91\]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[92\]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[93\]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[94\]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[95\]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[96\]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[97\]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[98\]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[99\]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 LA_DATA_IN\[9\]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[0\]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[100\]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[101\]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[102\]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[103\]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[104\]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[105\]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[106\]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[107\]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[108\]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[109\]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[10\]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[110\]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[111\]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[112\]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[113\]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[114\]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[115\]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[116\]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[117\]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[118\]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[119\]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[11\]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[120\]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[121\]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[122\]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[123\]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[124\]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[125\]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[126\]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[127\]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[12\]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[13\]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[14\]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[15\]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[16\]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[17\]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[18\]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[19\]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[1\]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[20\]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[21\]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[22\]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[23\]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[24\]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[25\]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[26\]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[27\]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[28\]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[29\]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[2\]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[30\]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[31\]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[32\]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[33\]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[34\]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[35\]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[36\]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[37\]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[38\]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[39\]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[3\]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[40\]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[41\]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[42\]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[43\]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[44\]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[45\]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[46\]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[47\]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[48\]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[49\]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[4\]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[50\]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[51\]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[52\]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[53\]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[54\]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[55\]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[56\]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[57\]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[58\]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[59\]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[5\]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[60\]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[61\]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[62\]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[63\]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[64\]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[65\]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[66\]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[67\]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[68\]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[69\]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[6\]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[70\]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[71\]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[72\]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[73\]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[74\]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[75\]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[76\]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[77\]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[78\]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[79\]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[7\]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[80\]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[81\]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[82\]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[83\]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[84\]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[85\]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[86\]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[87\]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[88\]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[89\]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[8\]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[90\]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[91\]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[92\]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[93\]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[94\]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[95\]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[96\]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[97\]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[98\]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[99\]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 LA_DATA_OUT\[9\]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 LA_OENB\[0\]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 LA_OENB\[100\]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 LA_OENB\[101\]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 LA_OENB\[102\]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 LA_OENB\[103\]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 LA_OENB\[104\]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 LA_OENB\[105\]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 LA_OENB\[106\]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 LA_OENB\[107\]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 LA_OENB\[108\]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 LA_OENB\[109\]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 LA_OENB\[10\]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 LA_OENB\[110\]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 LA_OENB\[111\]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 LA_OENB\[112\]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 LA_OENB\[113\]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 LA_OENB\[114\]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 LA_OENB\[115\]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 LA_OENB\[116\]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 LA_OENB\[117\]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 LA_OENB\[118\]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 LA_OENB\[119\]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 LA_OENB\[11\]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 LA_OENB\[120\]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 LA_OENB\[121\]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 LA_OENB\[122\]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 LA_OENB\[123\]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 LA_OENB\[124\]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 LA_OENB\[125\]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 LA_OENB\[126\]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 LA_OENB\[127\]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 LA_OENB\[12\]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 LA_OENB\[13\]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 LA_OENB\[14\]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 LA_OENB\[15\]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 LA_OENB\[16\]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 LA_OENB\[17\]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 LA_OENB\[18\]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 LA_OENB\[19\]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 LA_OENB\[1\]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 LA_OENB\[20\]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 LA_OENB\[21\]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 LA_OENB\[22\]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 LA_OENB\[23\]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 LA_OENB\[24\]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 LA_OENB\[25\]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 LA_OENB\[26\]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 LA_OENB\[27\]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 LA_OENB\[28\]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 LA_OENB\[29\]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 LA_OENB\[2\]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 LA_OENB\[30\]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 LA_OENB\[31\]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 LA_OENB\[32\]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 LA_OENB\[33\]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 LA_OENB\[34\]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 LA_OENB\[35\]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 LA_OENB\[36\]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 LA_OENB\[37\]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 LA_OENB\[38\]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 LA_OENB\[39\]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 LA_OENB\[3\]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 LA_OENB\[40\]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 LA_OENB\[41\]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 LA_OENB\[42\]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 LA_OENB\[43\]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 LA_OENB\[44\]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 LA_OENB\[45\]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 LA_OENB\[46\]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 LA_OENB\[47\]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 LA_OENB\[48\]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 LA_OENB\[49\]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 LA_OENB\[4\]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 LA_OENB\[50\]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 LA_OENB\[51\]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 LA_OENB\[52\]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 LA_OENB\[53\]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 LA_OENB\[54\]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 LA_OENB\[55\]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 LA_OENB\[56\]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 LA_OENB\[57\]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 LA_OENB\[58\]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 LA_OENB\[59\]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 LA_OENB\[5\]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 LA_OENB\[60\]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 LA_OENB\[61\]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 LA_OENB\[62\]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 LA_OENB\[63\]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 LA_OENB\[64\]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 LA_OENB\[65\]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 LA_OENB\[66\]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 LA_OENB\[67\]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 LA_OENB\[68\]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 LA_OENB\[69\]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 LA_OENB\[6\]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 LA_OENB\[70\]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 LA_OENB\[71\]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 LA_OENB\[72\]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 LA_OENB\[73\]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 LA_OENB\[74\]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 LA_OENB\[75\]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 LA_OENB\[76\]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 LA_OENB\[77\]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 LA_OENB\[78\]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 LA_OENB\[79\]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 LA_OENB\[7\]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 LA_OENB\[80\]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 LA_OENB\[81\]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 LA_OENB\[82\]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 LA_OENB\[83\]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 LA_OENB\[84\]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 LA_OENB\[85\]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 LA_OENB\[86\]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 LA_OENB\[87\]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 LA_OENB\[88\]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 LA_OENB\[89\]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 LA_OENB\[8\]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 LA_OENB\[90\]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 LA_OENB\[91\]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 LA_OENB\[92\]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 LA_OENB\[93\]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 LA_OENB\[94\]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 LA_OENB\[95\]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 LA_OENB\[96\]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 LA_OENB\[97\]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 LA_OENB\[98\]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 LA_OENB\[99\]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 LA_OENB\[9\]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 USER_CLOCK2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 USER_IRQ\[0\]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 USER_IRQ\[1\]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 USER_IRQ\[2\]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 VCCD1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 VCCD1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 VCCD2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 VCCD2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 VDDA1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 VDDA1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 VDDA1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 VDDA1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 VDDA2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 VDDA2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 VSSA1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 VSSA1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 VSSA1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 VSSA1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 VSSA2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 VSSA2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 VSSD1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 VSSD1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 VSSD2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 VSSD2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 WB_CLK_I
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 WB_RST_I
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 WBS_ACK_O
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[0\]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[10\]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[11\]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[12\]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[13\]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[14\]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[15\]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[16\]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[17\]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[18\]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[19\]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[1\]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[20\]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[21\]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[22\]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[23\]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[24\]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[25\]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[26\]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[27\]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[28\]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[29\]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[2\]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[30\]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[31\]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[3\]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[4\]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[5\]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[6\]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[7\]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[8\]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 WBS_ADR_I\[9\]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 WBS_CYC_I
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[0\]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[10\]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[11\]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[12\]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[13\]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[14\]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[15\]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[16\]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[17\]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[18\]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[19\]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[1\]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[20\]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[21\]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[22\]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[23\]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[24\]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[25\]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[26\]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[27\]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[28\]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[29\]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[2\]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[30\]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[31\]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[3\]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[4\]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[5\]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[6\]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[7\]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[8\]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 WBS_DAT_I\[9\]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[0\]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[10\]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[11\]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[12\]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[13\]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[14\]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[15\]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[16\]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[17\]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[18\]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[19\]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[1\]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[20\]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[21\]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[22\]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[23\]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[24\]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[25\]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[26\]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[27\]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[28\]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[29\]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[2\]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[30\]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[31\]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[3\]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[4\]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[5\]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[6\]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[7\]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[8\]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 WBS_DAT_O\[9\]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 WBS_SEL_I\[0\]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 WBS_SEL_I\[1\]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 WBS_SEL_I\[2\]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 WBS_SEL_I\[3\]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 WBS_STB_I
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 WBS_WE_I
port 677 nsew signal input
<< properties >>
string LEFclass CORE
string LEFsite unithd
string FIXED_BBOX 0 0 584000 704000
string LEFsymmetry X Y R90
<< end >>
