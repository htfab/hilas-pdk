magic
tech sky130A
timestamp 1628704245
<< checkpaint >>
rect 822 -230 2255 1680
<< error_s >>
rect 819 616 869 622
rect 891 616 941 622
rect 819 574 869 580
rect 891 574 941 580
rect 819 547 869 553
rect 819 505 869 511
rect 819 464 869 470
rect 819 422 869 428
rect 819 395 869 401
rect 891 395 941 401
rect 819 353 869 359
rect 891 353 941 359
rect 819 292 869 298
rect 891 292 941 298
rect 819 250 869 256
rect 891 250 941 256
rect 819 223 869 229
rect 819 181 869 187
rect 819 139 869 145
rect 819 97 869 103
rect 819 70 869 76
rect 891 70 941 76
rect 819 28 869 34
rect 891 28 941 34
<< nwell >>
rect 58 477 117 493
rect 432 471 543 498
rect 752 379 761 387
rect 896 329 913 335
rect 896 328 931 329
rect 896 318 913 328
rect 930 318 931 328
rect 58 153 117 168
rect 432 151 543 170
<< psubdiff >>
rect 258 482 283 505
rect 258 465 262 482
rect 279 465 283 482
rect 660 479 685 507
rect 258 437 283 465
rect 660 462 664 479
rect 681 462 685 479
rect 660 436 685 462
rect 258 355 284 397
rect 258 338 263 355
rect 280 338 284 355
rect 258 321 284 338
rect 258 304 263 321
rect 280 304 284 321
rect 258 287 284 304
rect 258 270 263 287
rect 280 270 284 287
rect 258 259 284 270
rect 660 361 687 382
rect 660 344 665 361
rect 682 344 687 361
rect 660 327 687 344
rect 660 310 665 327
rect 682 310 687 327
rect 660 293 687 310
rect 660 276 665 293
rect 682 276 687 293
rect 263 255 280 259
rect 660 258 687 276
<< mvnsubdiff >>
rect 58 477 117 493
rect 432 471 543 498
rect 58 153 117 168
rect 432 151 543 170
<< psubdiffcont >>
rect 262 465 279 482
rect 664 462 681 479
rect 263 338 280 355
rect 263 304 280 321
rect 263 270 280 287
rect 665 344 682 361
rect 665 310 682 327
rect 665 276 682 293
<< poly >>
rect 584 555 752 572
rect 159 527 392 551
rect 157 405 392 429
rect 584 403 752 420
rect 891 325 896 326
rect 913 328 931 329
rect 929 326 931 328
rect 913 325 941 326
rect 929 318 931 325
rect 157 225 394 249
rect 584 231 752 248
rect 159 93 396 117
rect 584 78 752 95
<< polycont >>
rect 896 318 913 335
<< locali >>
rect 262 482 279 484
rect 664 479 681 481
rect 263 321 280 338
rect 263 287 280 291
rect 665 327 682 344
rect 887 318 896 335
rect 665 293 682 295
<< viali >>
rect 262 484 279 501
rect 262 448 279 465
rect 664 481 681 498
rect 664 445 681 462
rect 263 355 280 372
rect 263 304 280 308
rect 263 291 280 304
rect 263 270 280 272
rect 263 255 280 270
rect 665 361 682 378
rect 913 318 931 335
rect 665 310 682 312
rect 665 295 682 310
rect 665 259 682 276
<< metal1 >>
rect 36 0 76 650
rect 257 501 284 650
rect 441 613 479 650
rect 257 484 262 501
rect 279 484 284 501
rect 257 465 284 484
rect 257 448 262 465
rect 279 448 284 465
rect 257 372 284 448
rect 257 355 263 372
rect 280 355 284 372
rect 257 308 284 355
rect 257 291 263 308
rect 280 291 284 308
rect 257 272 284 291
rect 257 255 263 272
rect 280 255 284 272
rect 257 176 284 255
rect 660 498 685 650
rect 875 616 891 623
rect 912 616 931 623
rect 956 616 972 623
rect 660 481 664 498
rect 681 481 685 498
rect 660 462 685 481
rect 660 445 664 462
rect 681 445 685 462
rect 660 378 685 445
rect 660 361 665 378
rect 682 361 685 378
rect 660 312 685 361
rect 910 335 934 338
rect 891 326 913 335
rect 875 325 913 326
rect 891 318 913 325
rect 931 318 934 335
rect 956 325 972 326
rect 910 315 934 318
rect 660 295 665 312
rect 682 295 685 312
rect 920 305 931 315
rect 660 276 685 295
rect 660 259 665 276
rect 682 259 685 276
rect 660 179 685 259
rect 659 176 687 179
rect 255 173 286 176
rect 255 147 257 173
rect 284 147 286 173
rect 658 175 688 176
rect 658 149 660 175
rect 686 149 688 175
rect 658 148 688 149
rect 255 145 286 147
rect 659 146 687 148
rect 257 0 284 145
rect 441 0 479 28
rect 660 0 685 146
rect 875 19 891 26
rect 912 19 931 26
rect 956 19 972 26
<< via1 >>
rect 257 147 284 173
rect 660 149 686 175
<< metal2 >>
rect 999 576 1008 594
rect 1 532 762 551
rect 999 533 1008 551
rect 1 424 764 442
rect 999 424 1008 442
rect 752 380 761 383
rect 999 381 1008 399
rect 752 369 764 380
rect 749 254 764 271
rect 997 252 1008 270
rect 1 213 48 229
rect 2 212 48 213
rect 78 210 764 227
rect 997 209 1008 227
rect 657 175 689 176
rect 254 147 257 173
rect 284 170 287 173
rect 657 170 660 175
rect 284 153 660 170
rect 284 147 287 153
rect 657 149 660 153
rect 686 149 689 175
rect 657 148 689 149
rect 1 114 764 131
rect 997 99 1008 117
rect 997 56 1008 74
use sky130_hilas_wellContact  sky130_hilas_wellContact_1
timestamp 1628285143
transform 1 0 1449 0 1 693
box -1448 -441 -1275 -255
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_0
timestamp 1628285143
transform 1 0 1333 0 1 395
box -957 -395 -734 -209
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_1
timestamp 1628285143
transform 1 0 1333 0 1 530
box -957 -395 -734 -209
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_2
timestamp 1628285143
transform 1 0 1333 0 1 715
box -957 -395 -734 -209
use sky130_hilas_wellContact  sky130_hilas_wellContact_0
timestamp 1628285143
transform 1 0 1852 0 1 686
box -1448 -441 -1275 -255
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_1
timestamp 1628285143
transform 1 0 1041 0 1 -41
box -289 41 -33 232
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_2
timestamp 1628285143
transform 1 0 1041 0 -1 367
box -289 41 -33 232
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_0
timestamp 1628285143
transform 1 0 1041 0 1 284
box -289 41 -33 232
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_3
timestamp 1628285143
transform 1 0 1333 0 1 859
box -957 -395 -734 -209
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_3
timestamp 1628285143
transform 1 0 1041 0 -1 691
box -289 41 -33 232
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_0
timestamp 1628704213
transform 1 0 1452 0 1 535
box 0 0 173 190
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_1
timestamp 1628704213
transform 1 0 1452 0 1 400
box 0 0 173 190
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_3
timestamp 1628704213
transform 1 0 1452 0 1 860
box 0 0 173 190
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_2
timestamp 1628704213
transform 1 0 1452 0 1 724
box 0 0 173 190
<< labels >>
rlabel metal2 1 213 13 229 0 ROW3
port 3 nsew analog default
rlabel metal2 1 115 15 130 0 ROW4
port 4 nsew analog default
rlabel metal1 36 609 76 623 0 VTUN
port 5 nsew analog default
rlabel metal1 36 18 76 28 0 VTUN
port 5 nsew analog default
rlabel metal1 441 18 479 28 0 GATE1
port 6 nsew analog default
rlabel metal1 441 613 479 623 0 GATE1
port 6 nsew analog default
rlabel metal1 956 616 972 623 0 VINJ
port 7 nsew power default
rlabel metal1 875 616 891 623 0 VPWR
port 8 nsew power default
rlabel metal1 912 616 931 623 0 COLSEL1
rlabel metal1 956 19 972 26 0 VINJ
port 7 nsew power default
rlabel metal1 875 19 891 26 0 VPWR
port 8 nsew power default
rlabel metal1 912 19 931 26 0 COLSEL1
port 9 nsew analog default
rlabel metal1 257 615 284 623 0 VGND
port 18 nsew
rlabel metal1 660 618 685 623 0 VGND
port 18 nsew
rlabel metal1 257 18 284 25 0 VGND
port 18 nsew
rlabel metal1 660 18 685 25 0 VGND
port 18 nsew
rlabel metal2 997 209 1008 227 0 ROW3
port 3 nsew
rlabel metal2 997 252 1008 270 0 DRAIN3
port 19 nsew
rlabel metal2 997 56 1008 74 0 DRAIN4
port 20 nsew
rlabel metal2 997 99 1008 117 0 ROW4
port 4 nsew
rlabel metal2 999 576 1008 594 0 DRAIN1
port 21 nsew
rlabel metal2 999 533 1008 551 0 ROW1
port 1 nsew
rlabel metal2 999 424 1008 442 0 ROW2
port 2 nsew
rlabel metal2 999 381 1008 399 0 DRAIN2
port 22 nsew
rlabel space 0 532 12 551 0 ROW1
port 1 nsew
rlabel metal2 1 424 7 442 0 ROW2
port 2 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
