VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_drainSelect01
  CLASS BLOCK ;
  FOREIGN sky130_hilas_drainSelect01 ;
  ORIGIN -10.720 -0.050 ;
  SIZE 5.420 BY 6.050 ;
  PIN drain4
    PORT
      LAYER met2 ;
        RECT 11.070 0.570 12.280 0.740 ;
    END
  END drain4
  PIN drain3
    PORT
      LAYER met2 ;
        RECT 11.070 2.410 11.770 2.580 ;
    END
  END drain3
  PIN drain2
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 11.070 3.560 11.740 3.740 ;
    END
  END drain2
  PIN drain1
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 11.070 5.420 11.800 5.600 ;
    END
  END drain1
  PIN DrainSelect1
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 15.990 4.980 16.140 5.220 ;
    END
  END DrainSelect1
  PIN DrainSelect2
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 15.990 3.860 16.140 4.100 ;
    END
  END DrainSelect2
  PIN DrainSelect3
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 15.990 2.050 16.140 2.290 ;
    END
  END DrainSelect3
  PIN DrainSelect4
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 15.990 0.930 16.140 1.170 ;
    END
  END DrainSelect4
  PIN Vinj
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 11.080 5.370 11.330 6.100 ;
    END
  END Vinj
  PIN Drain_Mux
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 14.070 5.700 14.300 6.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 14.070 0.050 14.300 0.450 ;
    END
  END Drain_Mux
  PIN GND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 15.420 0.050 15.610 1.080 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.420 5.070 15.610 6.100 ;
    END
  END GND
  OBS
      LAYER nwell ;
        RECT 10.720 0.050 13.920 6.100 ;
      LAYER li1 ;
        RECT 11.120 0.380 15.990 5.770 ;
      LAYER met1 ;
        RECT 11.610 5.420 13.790 5.770 ;
        RECT 14.580 5.420 15.140 5.770 ;
        RECT 15.890 5.500 15.990 5.770 ;
        RECT 11.610 5.090 15.140 5.420 ;
        RECT 11.080 4.790 15.140 5.090 ;
        RECT 11.080 4.700 15.710 4.790 ;
        RECT 11.080 4.380 15.990 4.700 ;
        RECT 11.080 3.580 15.710 4.380 ;
        RECT 11.080 2.570 15.990 3.580 ;
        RECT 11.080 1.770 15.710 2.570 ;
        RECT 11.080 1.450 15.990 1.770 ;
        RECT 11.080 1.360 15.710 1.450 ;
        RECT 11.080 0.730 15.140 1.360 ;
        RECT 11.080 0.050 13.790 0.730 ;
        RECT 14.580 0.050 15.140 0.730 ;
        RECT 15.890 0.050 15.990 0.650 ;
      LAYER met2 ;
        RECT 12.080 5.140 14.980 5.770 ;
        RECT 11.740 4.020 14.980 5.140 ;
        RECT 12.020 3.280 14.980 4.020 ;
        RECT 11.740 2.860 14.980 3.280 ;
        RECT 12.050 2.130 14.980 2.860 ;
        RECT 11.740 1.020 14.980 2.130 ;
        RECT 12.560 0.380 14.980 1.020 ;
  END
END sky130_hilas_drainSelect01
END LIBRARY

