magic
tech sky130A
timestamp 1607802006
<< metal3 >>
rect -443 333 -161 336
rect -443 -245 277 333
rect -164 -247 277 -245
<< mimcap >>
rect -404 -104 234 295
rect -404 -105 -288 -104
rect -404 -118 -316 -105
rect -302 -118 -288 -105
rect -274 -118 -260 -104
rect -246 -118 -232 -104
rect -218 -118 -204 -104
rect -190 -118 -176 -104
rect -162 -118 -149 -104
rect -135 -118 -121 -104
rect -107 -118 -93 -104
rect -79 -118 234 -104
rect -404 -205 234 -118
<< mimcapcontact >>
rect -316 -118 -302 -105
rect -288 -118 -274 -104
rect -260 -118 -246 -104
rect -232 -118 -218 -104
rect -204 -118 -190 -104
rect -176 -118 -162 -104
rect -149 -118 -135 -104
rect -121 -118 -107 -104
rect -93 -118 -79 -104
<< metal4 >>
rect -354 -104 -50 -90
rect -354 -105 -288 -104
rect -354 -118 -316 -105
rect -302 -118 -288 -105
rect -274 -118 -260 -104
rect -246 -118 -232 -104
rect -218 -118 -204 -104
rect -190 -118 -176 -104
rect -162 -118 -149 -104
rect -135 -118 -121 -104
rect -107 -118 -93 -104
rect -79 -118 -50 -104
rect -354 -137 -50 -118
<< end >>
