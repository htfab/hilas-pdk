magic
tech sky130A
timestamp 1629137254
<< checkpaint >>
rect -294 7973 1995 8407
rect -294 7968 2531 7973
rect -294 7331 3001 7968
rect -795 7326 3001 7331
rect -1081 7255 3001 7326
rect -1081 7223 3889 7255
rect -1082 6933 3889 7223
rect -1082 6900 4708 6933
rect -1082 6686 4710 6900
rect -1082 6504 5339 6686
rect -1082 6471 5732 6504
rect -1082 6151 5734 6471
rect 5915 6175 8829 6504
rect 5915 6151 8907 6175
rect -1082 5769 8907 6151
rect 10233 6026 11525 6032
rect 10233 6011 11853 6026
rect -1082 5709 210 5769
rect 1107 5754 8907 5769
rect 1107 4597 2681 5754
rect 1209 4340 2681 4597
rect 3190 5174 8907 5754
rect 9932 5174 11853 6011
rect 3190 4110 11853 5174
rect 1048 3833 2407 3842
rect 935 3798 2407 3833
rect 926 3668 2407 3798
rect 3190 3757 10206 4110
rect 10233 4095 11853 4110
rect 10233 4089 11525 4095
rect 876 3620 2407 3668
rect 857 3619 2407 3620
rect 857 3565 2431 3619
rect 857 3549 2432 3565
rect 857 3547 2635 3549
rect 758 2786 2635 3547
rect 539 2102 2635 2786
rect 3186 2824 10206 3757
rect 3186 2747 7682 2824
rect 3186 2546 7683 2747
rect 539 2033 2411 2102
rect 539 2022 2316 2033
rect 539 976 2317 2022
rect 3186 1710 7740 2546
rect 9729 2501 11494 2512
rect 9633 2235 11494 2501
rect 4083 1253 7740 1710
rect 4083 1251 7739 1253
rect 4084 1207 7739 1251
rect 4084 1204 6184 1207
rect 6445 1206 7739 1207
rect 683 729 2317 976
rect 683 228 2282 729
rect 9596 -175 11494 2235
rect 9633 -369 11494 -175
rect 9833 -455 11468 -369
rect 10022 -457 11337 -455
<< error_s >>
rect 2146 6926 2175 6942
rect 2225 6926 2254 6942
rect 2304 6926 2333 6942
rect 2383 6926 2412 6942
rect 2146 6892 2147 6893
rect 2174 6892 2175 6893
rect 2225 6892 2226 6893
rect 2253 6892 2254 6893
rect 2304 6892 2305 6893
rect 2332 6892 2333 6893
rect 2383 6892 2384 6893
rect 2411 6892 2412 6893
rect 2096 6863 2113 6892
rect 2145 6891 2176 6892
rect 2224 6891 2255 6892
rect 2303 6891 2334 6892
rect 2382 6891 2413 6892
rect 2146 6884 2175 6891
rect 2225 6884 2254 6891
rect 2304 6884 2333 6891
rect 2383 6884 2412 6891
rect 2146 6870 2155 6884
rect 2402 6870 2412 6884
rect 2146 6864 2175 6870
rect 2225 6864 2254 6870
rect 2304 6864 2333 6870
rect 2383 6864 2412 6870
rect 2145 6863 2176 6864
rect 2224 6863 2255 6864
rect 2303 6863 2334 6864
rect 2382 6863 2413 6864
rect 2444 6863 2462 6892
rect 2146 6862 2147 6863
rect 2174 6862 2175 6863
rect 2225 6862 2226 6863
rect 2253 6862 2254 6863
rect 2304 6862 2305 6863
rect 2332 6862 2333 6863
rect 2383 6862 2384 6863
rect 2411 6862 2412 6863
rect 2146 6813 2175 6828
rect 2225 6813 2254 6828
rect 2304 6813 2333 6828
rect 2383 6813 2412 6828
rect 2146 6646 2175 6662
rect 2225 6646 2254 6662
rect 2304 6646 2333 6662
rect 2383 6646 2412 6662
rect 2146 6612 2147 6613
rect 2174 6612 2175 6613
rect 2225 6612 2226 6613
rect 2253 6612 2254 6613
rect 2304 6612 2305 6613
rect 2332 6612 2333 6613
rect 2383 6612 2384 6613
rect 2411 6612 2412 6613
rect 2096 6583 2113 6612
rect 2145 6611 2176 6612
rect 2224 6611 2255 6612
rect 2303 6611 2334 6612
rect 2382 6611 2413 6612
rect 2146 6604 2175 6611
rect 2225 6604 2254 6611
rect 2304 6604 2333 6611
rect 2383 6604 2412 6611
rect 2146 6590 2155 6604
rect 2402 6590 2412 6604
rect 2146 6584 2175 6590
rect 2225 6584 2254 6590
rect 2304 6584 2333 6590
rect 2383 6584 2412 6590
rect 2145 6583 2176 6584
rect 2224 6583 2255 6584
rect 2303 6583 2334 6584
rect 2382 6583 2413 6584
rect 2444 6583 2462 6612
rect 2146 6582 2147 6583
rect 2174 6582 2175 6583
rect 2225 6582 2226 6583
rect 2253 6582 2254 6583
rect 2304 6582 2305 6583
rect 2332 6582 2333 6583
rect 2383 6582 2384 6583
rect 2411 6582 2412 6583
rect 3242 6564 3271 6582
rect 2146 6533 2175 6548
rect 2225 6533 2254 6548
rect 2304 6533 2333 6548
rect 2383 6533 2412 6548
rect 3242 6532 3243 6533
rect 3270 6532 3271 6533
rect 2146 6491 2175 6507
rect 2225 6491 2254 6507
rect 2304 6491 2333 6507
rect 2383 6491 2412 6507
rect 3192 6503 3210 6532
rect 3241 6531 3272 6532
rect 3242 6522 3271 6531
rect 3242 6513 3252 6522
rect 3261 6513 3271 6522
rect 3242 6504 3271 6513
rect 3241 6503 3272 6504
rect 3303 6503 3321 6532
rect 3242 6502 3243 6503
rect 3270 6502 3271 6503
rect 2146 6457 2147 6458
rect 2174 6457 2175 6458
rect 2225 6457 2226 6458
rect 2253 6457 2254 6458
rect 2304 6457 2305 6458
rect 2332 6457 2333 6458
rect 2383 6457 2384 6458
rect 2411 6457 2412 6458
rect 2096 6428 2113 6457
rect 2145 6456 2176 6457
rect 2224 6456 2255 6457
rect 2303 6456 2334 6457
rect 2382 6456 2413 6457
rect 2146 6449 2175 6456
rect 2225 6449 2254 6456
rect 2304 6449 2333 6456
rect 2383 6449 2412 6456
rect 2146 6435 2155 6449
rect 2402 6435 2412 6449
rect 2146 6429 2175 6435
rect 2225 6429 2254 6435
rect 2304 6429 2333 6435
rect 2383 6429 2412 6435
rect 2145 6428 2176 6429
rect 2224 6428 2255 6429
rect 2303 6428 2334 6429
rect 2382 6428 2413 6429
rect 2444 6428 2462 6457
rect 3242 6453 3271 6471
rect 2146 6427 2147 6428
rect 2174 6427 2175 6428
rect 2225 6427 2226 6428
rect 2253 6427 2254 6428
rect 2304 6427 2305 6428
rect 2332 6427 2333 6428
rect 2383 6427 2384 6428
rect 2411 6427 2412 6428
rect 2146 6378 2175 6393
rect 2225 6378 2254 6393
rect 2304 6378 2333 6393
rect 2383 6378 2412 6393
rect 4024 5824 4052 5830
rect 4166 5823 4194 5830
rect 4301 5824 4351 5830
rect 4624 5823 4674 5829
rect 4024 5782 4052 5788
rect 4166 5781 4194 5788
rect 4301 5782 4351 5788
rect 4624 5781 4674 5787
rect 3975 5752 4003 5758
rect 4215 5752 4243 5758
rect 4372 5752 4423 5758
rect 4553 5757 4603 5763
rect 3975 5710 4003 5716
rect 4215 5710 4243 5716
rect 4372 5710 4423 5716
rect 4553 5715 4603 5721
rect 4024 5649 4052 5655
rect 4166 5648 4194 5655
rect 4301 5649 4351 5655
rect 4624 5648 4674 5654
rect 4024 5607 4052 5613
rect 4166 5606 4194 5613
rect 4301 5607 4351 5613
rect 4624 5606 4674 5612
rect 3975 5577 4003 5583
rect 4215 5577 4243 5583
rect 4372 5577 4423 5583
rect 4553 5582 4603 5588
rect 3975 5535 4003 5541
rect 4215 5535 4243 5541
rect 4372 5535 4423 5541
rect 4553 5540 4603 5546
rect 4024 5474 4052 5480
rect 4166 5473 4194 5480
rect 4301 5474 4351 5480
rect 4624 5473 4674 5479
rect 5468 5446 5518 5452
rect 5540 5446 5590 5452
rect 7509 5446 7559 5452
rect 7581 5446 7631 5452
rect 7969 5450 7996 5456
rect 4024 5432 4052 5438
rect 4166 5431 4194 5438
rect 4301 5432 4351 5438
rect 4624 5431 4674 5437
rect 3975 5402 4003 5408
rect 4215 5402 4243 5408
rect 4372 5402 4423 5408
rect 4553 5407 4603 5413
rect 5468 5404 5518 5410
rect 5540 5404 5590 5410
rect 7509 5404 7559 5410
rect 7581 5404 7631 5410
rect 7969 5408 7996 5414
rect 7969 5383 7996 5389
rect 3975 5360 4003 5366
rect 4215 5360 4243 5366
rect 4372 5360 4423 5366
rect 4553 5365 4603 5371
rect 4024 5299 4052 5305
rect 4166 5298 4194 5305
rect 4301 5299 4351 5305
rect 4624 5298 4674 5304
rect 5653 5302 5656 5352
rect 5695 5302 5698 5352
rect 5789 5302 5791 5352
rect 5831 5302 5833 5352
rect 7969 5341 7996 5347
rect 7969 5300 7996 5306
rect 4024 5257 4052 5263
rect 4166 5256 4194 5263
rect 4301 5257 4351 5263
rect 4624 5256 4674 5262
rect 3975 5227 4003 5233
rect 4215 5227 4243 5233
rect 4372 5227 4423 5233
rect 4553 5232 4603 5238
rect 5653 5223 5656 5273
rect 5695 5223 5698 5273
rect 5789 5223 5791 5273
rect 5831 5223 5833 5273
rect 7969 5258 7996 5264
rect 7969 5233 7996 5239
rect 3975 5185 4003 5191
rect 4215 5185 4243 5191
rect 4372 5185 4423 5191
rect 4553 5190 4603 5196
rect 7969 5191 7996 5197
rect 10727 5193 10767 5199
rect 10877 5193 10917 5199
rect 7969 5150 7996 5156
rect 10727 5151 10767 5157
rect 10877 5151 10917 5157
rect 4878 5133 4928 5138
rect 5058 5133 5108 5139
rect 5198 5133 5248 5138
rect 3975 5124 4003 5130
rect 4215 5124 4243 5130
rect 4372 5124 4423 5130
rect 10651 5127 10691 5132
rect 10877 5125 10917 5132
rect 4553 5119 4603 5125
rect 4878 5091 4928 5096
rect 5058 5091 5108 5097
rect 5198 5091 5248 5096
rect 3975 5082 4003 5088
rect 4215 5082 4243 5088
rect 4372 5082 4423 5088
rect 4553 5077 4603 5083
rect 4878 5066 4928 5072
rect 5198 5066 5248 5072
rect 5653 5070 5656 5120
rect 5695 5070 5698 5120
rect 5789 5070 5791 5120
rect 5831 5070 5833 5120
rect 7969 5108 7996 5114
rect 7969 5083 7996 5089
rect 10651 5085 10691 5090
rect 10877 5083 10917 5090
rect 4024 5052 4052 5058
rect 4166 5052 4194 5059
rect 4301 5052 4351 5058
rect 4624 5053 4674 5059
rect 7969 5041 7996 5047
rect 4878 5024 4928 5030
rect 5198 5024 5248 5030
rect 4024 5010 4052 5016
rect 4166 5010 4194 5017
rect 4301 5010 4351 5016
rect 4624 5011 4674 5017
rect 5653 4991 5656 5041
rect 5695 4991 5698 5041
rect 5789 4991 5791 5041
rect 5831 4991 5833 5041
rect 10651 5023 10691 5028
rect 10877 5023 10917 5030
rect 7969 5000 7996 5006
rect 10651 4981 10691 4986
rect 10877 4981 10917 4988
rect 4878 4963 4928 4969
rect 5198 4963 5248 4969
rect 7969 4958 7996 4964
rect 10727 4956 10767 4962
rect 10877 4956 10917 4962
rect 3975 4949 4003 4955
rect 4215 4949 4243 4955
rect 4372 4949 4423 4955
rect 4553 4944 4603 4950
rect 5468 4933 5518 4939
rect 5540 4933 5590 4939
rect 7509 4933 7559 4939
rect 7581 4933 7631 4939
rect 7969 4933 7996 4939
rect 4878 4921 4928 4927
rect 5198 4921 5248 4927
rect 10727 4914 10767 4920
rect 10877 4914 10917 4920
rect 3975 4907 4003 4913
rect 4215 4907 4243 4913
rect 4372 4907 4423 4913
rect 4553 4902 4603 4908
rect 4878 4897 4928 4902
rect 5058 4896 5108 4902
rect 5198 4897 5248 4902
rect 5468 4891 5518 4897
rect 5540 4891 5590 4897
rect 7509 4891 7559 4897
rect 7581 4891 7631 4897
rect 7969 4891 7996 4897
rect 4024 4877 4052 4883
rect 4166 4877 4194 4884
rect 4301 4877 4351 4883
rect 4624 4878 4674 4884
rect 10727 4873 10767 4879
rect 10877 4873 10917 4879
rect 4878 4855 4928 4860
rect 5058 4854 5108 4860
rect 5198 4855 5248 4860
rect 5469 4843 5519 4849
rect 5541 4843 5591 4849
rect 7509 4843 7559 4849
rect 7581 4843 7631 4849
rect 7969 4847 7996 4853
rect 4024 4835 4052 4841
rect 4166 4835 4194 4842
rect 4301 4835 4351 4841
rect 4624 4836 4674 4842
rect 10727 4831 10767 4837
rect 10877 4831 10917 4837
rect 4878 4813 4928 4818
rect 5058 4813 5108 4819
rect 5198 4813 5248 4818
rect 5469 4801 5519 4807
rect 5541 4801 5591 4807
rect 7509 4801 7559 4807
rect 7581 4801 7631 4807
rect 7969 4805 7996 4811
rect 10651 4807 10691 4812
rect 10877 4805 10917 4812
rect 7969 4780 7996 4786
rect 3975 4774 4003 4780
rect 4215 4774 4243 4780
rect 4372 4774 4423 4780
rect 4553 4769 4603 4775
rect 4878 4771 4928 4776
rect 5058 4771 5108 4777
rect 5198 4771 5248 4776
rect 10651 4765 10691 4770
rect 10877 4763 10917 4770
rect 4878 4746 4928 4752
rect 5198 4746 5248 4752
rect 7969 4738 7996 4744
rect 3975 4732 4003 4738
rect 4215 4732 4243 4738
rect 4372 4732 4423 4738
rect 4553 4727 4603 4733
rect 4024 4702 4052 4708
rect 4166 4702 4194 4709
rect 4301 4702 4351 4708
rect 4624 4703 4674 4709
rect 4878 4704 4928 4710
rect 5198 4704 5248 4710
rect 10651 4703 10691 4708
rect 10877 4703 10917 4710
rect 7969 4697 7996 4703
rect 4024 4660 4052 4666
rect 4166 4660 4194 4667
rect 4301 4660 4351 4666
rect 4624 4661 4674 4667
rect 10651 4661 10691 4666
rect 10877 4661 10917 4668
rect 7969 4655 7996 4661
rect 4878 4643 4928 4649
rect 5198 4643 5248 4649
rect 10727 4636 10767 4642
rect 10877 4636 10917 4642
rect 7969 4630 7996 4636
rect 3975 4599 4003 4605
rect 4215 4599 4243 4605
rect 4372 4599 4423 4605
rect 4878 4601 4928 4607
rect 5198 4601 5248 4607
rect 4553 4594 4603 4600
rect 10727 4594 10767 4600
rect 10877 4594 10917 4600
rect 7969 4588 7996 4594
rect 4878 4577 4928 4582
rect 5058 4576 5108 4582
rect 5198 4577 5248 4582
rect 3975 4557 4003 4563
rect 4215 4557 4243 4563
rect 4372 4557 4423 4563
rect 4553 4552 4603 4558
rect 7969 4547 7996 4553
rect 4878 4535 4928 4540
rect 5058 4534 5108 4540
rect 5198 4535 5248 4540
rect 4024 4527 4052 4533
rect 4166 4527 4194 4534
rect 4301 4527 4351 4533
rect 4624 4528 4674 4534
rect 7969 4505 7996 4511
rect 4024 4485 4052 4491
rect 4166 4485 4194 4492
rect 4301 4485 4351 4491
rect 4624 4486 4674 4492
rect 7969 4480 7996 4486
rect 7969 4438 7996 4444
rect 7969 4397 7996 4403
rect 7969 4355 7996 4361
rect 5469 4330 5519 4336
rect 5541 4330 5591 4336
rect 7509 4330 7559 4336
rect 7581 4330 7631 4336
rect 7969 4330 7996 4336
rect 5469 4288 5519 4294
rect 5541 4288 5591 4294
rect 7509 4288 7559 4294
rect 7581 4288 7631 4294
rect 7969 4288 7996 4294
rect 3975 4111 4003 4117
rect 4215 4111 4243 4117
rect 4372 4111 4423 4117
rect 4553 4106 4603 4112
rect 4876 4086 4926 4091
rect 5056 4086 5106 4092
rect 5196 4086 5246 4091
rect 5610 4085 5660 4091
rect 5682 4085 5732 4091
rect 7366 4085 7416 4091
rect 7438 4085 7488 4091
rect 3975 4069 4003 4075
rect 4215 4069 4243 4075
rect 4372 4069 4423 4075
rect 4553 4064 4603 4070
rect 4024 4039 4052 4045
rect 4166 4039 4194 4046
rect 4301 4039 4351 4045
rect 4624 4040 4674 4046
rect 4876 4044 4926 4049
rect 5056 4044 5106 4050
rect 5196 4044 5246 4049
rect 5610 4043 5660 4049
rect 5682 4043 5732 4049
rect 7366 4043 7416 4049
rect 7438 4043 7488 4049
rect 4876 4019 4926 4025
rect 5196 4019 5246 4025
rect 5682 4016 5732 4022
rect 7366 4016 7416 4022
rect 4024 3997 4052 4003
rect 4166 3997 4194 4004
rect 4301 3997 4351 4003
rect 4624 3998 4674 4004
rect 4876 3977 4926 3983
rect 5196 3977 5246 3983
rect 5682 3974 5732 3980
rect 7366 3974 7416 3980
rect 3975 3936 4003 3942
rect 4215 3936 4243 3942
rect 4372 3936 4423 3942
rect 4553 3931 4603 3937
rect 5682 3931 5732 3937
rect 7366 3931 7416 3937
rect 4876 3916 4926 3922
rect 5196 3916 5246 3922
rect 3975 3894 4003 3900
rect 4215 3894 4243 3900
rect 4372 3894 4423 3900
rect 4553 3889 4603 3895
rect 5682 3889 5732 3895
rect 7366 3889 7416 3895
rect 4876 3874 4926 3880
rect 5196 3874 5246 3880
rect 4024 3864 4052 3870
rect 4166 3864 4194 3871
rect 4301 3864 4351 3870
rect 4624 3865 4674 3871
rect 5610 3862 5660 3868
rect 5682 3862 5732 3868
rect 7366 3862 7416 3868
rect 7438 3862 7488 3868
rect 4876 3850 4926 3855
rect 5056 3849 5106 3855
rect 5196 3850 5246 3855
rect 4024 3822 4052 3828
rect 4166 3822 4194 3829
rect 4301 3822 4351 3828
rect 4624 3823 4674 3829
rect 5610 3820 5660 3826
rect 5682 3820 5732 3826
rect 7366 3820 7416 3826
rect 7438 3820 7488 3826
rect 4876 3808 4926 3813
rect 5056 3807 5106 3813
rect 5196 3808 5246 3813
rect 3975 3761 4003 3767
rect 4215 3761 4243 3767
rect 4372 3761 4423 3767
rect 4876 3766 4926 3771
rect 5056 3766 5106 3772
rect 5196 3766 5246 3771
rect 4553 3756 4603 3762
rect 5610 3761 5660 3767
rect 5682 3761 5732 3767
rect 7366 3761 7416 3767
rect 7438 3761 7488 3767
rect 3975 3719 4003 3725
rect 4215 3719 4243 3725
rect 4372 3719 4423 3725
rect 4876 3724 4926 3729
rect 5056 3724 5106 3730
rect 5196 3724 5246 3729
rect 4553 3714 4603 3720
rect 5610 3719 5660 3725
rect 5682 3719 5732 3725
rect 7366 3719 7416 3725
rect 7438 3719 7488 3725
rect 4876 3699 4926 3705
rect 5196 3699 5246 3705
rect 4024 3689 4052 3695
rect 4166 3689 4194 3696
rect 4301 3689 4351 3695
rect 4624 3690 4674 3696
rect 5682 3692 5732 3698
rect 7366 3692 7416 3698
rect 4876 3657 4926 3663
rect 5196 3657 5246 3663
rect 4024 3647 4052 3653
rect 4166 3647 4194 3654
rect 4301 3647 4351 3653
rect 4624 3648 4674 3654
rect 5682 3650 5732 3656
rect 7366 3650 7416 3656
rect 5682 3608 5732 3614
rect 7366 3608 7416 3614
rect 4876 3596 4926 3602
rect 5196 3596 5246 3602
rect 3975 3586 4003 3592
rect 4215 3586 4243 3592
rect 4372 3586 4423 3592
rect 4553 3581 4603 3587
rect 5682 3566 5732 3572
rect 7366 3566 7416 3572
rect 4876 3554 4926 3560
rect 5196 3554 5246 3560
rect 3975 3544 4003 3550
rect 4215 3544 4243 3550
rect 4372 3544 4423 3550
rect 4553 3539 4603 3545
rect 5610 3539 5660 3545
rect 5682 3539 5732 3545
rect 7366 3539 7416 3545
rect 7438 3539 7488 3545
rect 4876 3530 4926 3535
rect 5056 3529 5106 3535
rect 5196 3530 5246 3535
rect 4024 3514 4052 3520
rect 4166 3514 4194 3521
rect 4301 3514 4351 3520
rect 4624 3515 4674 3521
rect 5610 3497 5660 3503
rect 5682 3497 5732 3503
rect 7366 3497 7416 3503
rect 7438 3497 7488 3503
rect 4876 3488 4926 3493
rect 5056 3487 5106 3493
rect 5196 3488 5246 3493
rect 4024 3472 4052 3478
rect 4166 3472 4194 3479
rect 4301 3472 4351 3478
rect 4624 3473 4674 3479
rect 3971 3205 3999 3211
rect 4211 3205 4239 3211
rect 4368 3205 4419 3211
rect 4549 3200 4599 3206
rect 3971 3163 3999 3169
rect 4211 3163 4239 3169
rect 4368 3163 4419 3169
rect 4549 3158 4599 3164
rect 4879 3159 4929 3164
rect 5059 3159 5109 3165
rect 5199 3159 5249 3164
rect 5613 3152 5663 3158
rect 5685 3152 5735 3158
rect 4020 3133 4048 3139
rect 4162 3133 4190 3140
rect 4297 3133 4347 3139
rect 4620 3134 4670 3140
rect 4879 3117 4929 3122
rect 5059 3117 5109 3123
rect 5199 3117 5249 3122
rect 5613 3110 5663 3116
rect 5685 3110 5735 3116
rect 4020 3091 4048 3097
rect 4162 3091 4190 3098
rect 4297 3091 4347 3097
rect 4620 3092 4670 3098
rect 4879 3092 4929 3098
rect 5199 3092 5249 3098
rect 5685 3083 5735 3089
rect 4879 3050 4929 3056
rect 5199 3050 5249 3056
rect 5685 3041 5735 3047
rect 3971 3030 3999 3036
rect 4211 3030 4239 3036
rect 4368 3030 4419 3036
rect 4549 3025 4599 3031
rect 5685 3000 5735 3006
rect 3971 2988 3999 2994
rect 4211 2988 4239 2994
rect 4368 2988 4419 2994
rect 4879 2989 4929 2995
rect 5199 2989 5249 2995
rect 4549 2983 4599 2989
rect 4020 2958 4048 2964
rect 4162 2958 4190 2965
rect 4297 2958 4347 2964
rect 4620 2959 4670 2965
rect 5685 2958 5735 2964
rect 4879 2947 4929 2953
rect 5199 2947 5249 2953
rect 5613 2931 5663 2937
rect 5685 2931 5735 2937
rect 4879 2923 4929 2928
rect 4020 2916 4048 2922
rect 4162 2916 4190 2923
rect 4297 2916 4347 2922
rect 4620 2917 4670 2923
rect 5059 2922 5109 2928
rect 5199 2923 5249 2928
rect 5613 2889 5663 2895
rect 5685 2889 5735 2895
rect 4879 2881 4929 2886
rect 5059 2880 5109 2886
rect 5199 2881 5249 2886
rect 3971 2855 3999 2861
rect 4211 2855 4239 2861
rect 4368 2855 4419 2861
rect 4549 2850 4599 2856
rect 4879 2839 4929 2844
rect 5059 2839 5109 2845
rect 5199 2839 5249 2844
rect 5613 2828 5663 2834
rect 5685 2828 5735 2834
rect 3971 2813 3999 2819
rect 4211 2813 4239 2819
rect 4368 2813 4419 2819
rect 4549 2808 4599 2814
rect 4879 2797 4929 2802
rect 5059 2797 5109 2803
rect 5199 2797 5249 2802
rect 4020 2783 4048 2789
rect 4162 2783 4190 2790
rect 4297 2783 4347 2789
rect 4620 2784 4670 2790
rect 5613 2786 5663 2792
rect 5685 2786 5735 2792
rect 4879 2772 4929 2778
rect 5199 2772 5249 2778
rect 5685 2759 5735 2765
rect 4020 2741 4048 2747
rect 4162 2741 4190 2748
rect 4297 2741 4347 2747
rect 4620 2742 4670 2748
rect 4879 2730 4929 2736
rect 5199 2730 5249 2736
rect 5685 2717 5735 2723
rect 3971 2680 3999 2686
rect 4211 2680 4239 2686
rect 4368 2680 4419 2686
rect 4549 2675 4599 2681
rect 5685 2675 5735 2681
rect 4879 2669 4929 2675
rect 5199 2669 5249 2675
rect 3971 2638 3999 2644
rect 4211 2638 4239 2644
rect 4368 2638 4419 2644
rect 4549 2633 4599 2639
rect 5685 2633 5735 2639
rect 4879 2627 4929 2633
rect 5199 2627 5249 2633
rect 4020 2608 4048 2614
rect 4162 2608 4190 2615
rect 4297 2608 4347 2614
rect 4620 2609 4670 2615
rect 4879 2603 4929 2608
rect 5059 2602 5109 2608
rect 5199 2603 5249 2608
rect 5613 2606 5663 2612
rect 5685 2606 5735 2612
rect 4020 2566 4048 2572
rect 4162 2566 4190 2573
rect 4297 2566 4347 2572
rect 4620 2567 4670 2573
rect 4879 2561 4929 2566
rect 5059 2560 5109 2566
rect 5199 2561 5249 2566
rect 5613 2564 5663 2570
rect 5685 2564 5735 2570
rect 10241 1692 10244 1731
rect 10283 1692 10286 1731
rect 10337 1692 10340 1731
rect 10379 1692 10382 1731
rect 10433 1692 10436 1731
rect 10475 1692 10478 1731
rect 10529 1692 10532 1731
rect 10571 1692 10574 1731
rect 10625 1692 10628 1731
rect 10667 1692 10670 1731
rect 10721 1692 10724 1731
rect 10763 1692 10766 1731
rect 10241 1531 10244 1570
rect 10283 1531 10286 1570
rect 10337 1530 10340 1569
rect 10379 1530 10382 1569
rect 10433 1530 10436 1569
rect 10475 1530 10478 1569
rect 10529 1530 10532 1569
rect 10571 1530 10574 1569
rect 10625 1530 10628 1569
rect 10667 1530 10670 1569
rect 10721 1531 10724 1570
rect 10763 1531 10766 1570
rect 10241 1370 10244 1409
rect 10283 1370 10286 1409
rect 10337 1369 10340 1408
rect 10379 1369 10382 1408
rect 10433 1369 10436 1408
rect 10475 1369 10478 1408
rect 10529 1369 10532 1408
rect 10571 1369 10574 1408
rect 10625 1369 10628 1408
rect 10667 1369 10670 1408
rect 10721 1370 10724 1409
rect 10763 1370 10766 1409
rect 10241 1209 10244 1248
rect 10283 1209 10286 1248
rect 10337 1208 10340 1247
rect 10379 1208 10382 1247
rect 10433 1208 10436 1247
rect 10475 1208 10478 1247
rect 10529 1208 10532 1247
rect 10571 1208 10574 1247
rect 10625 1208 10628 1247
rect 10667 1208 10670 1247
rect 10721 1209 10724 1248
rect 10763 1209 10766 1248
rect 10241 1048 10244 1087
rect 10283 1048 10286 1087
rect 10337 1047 10340 1086
rect 10379 1047 10382 1086
rect 10433 1047 10436 1086
rect 10475 1047 10478 1086
rect 10529 1047 10532 1086
rect 10571 1047 10574 1086
rect 10625 1047 10628 1086
rect 10667 1047 10670 1086
rect 10721 1048 10724 1087
rect 10763 1048 10766 1087
rect 10509 997 10513 998
rect 10241 887 10244 926
rect 10283 887 10286 926
rect 10337 886 10340 925
rect 10379 886 10382 925
rect 10433 886 10436 925
rect 10475 886 10478 925
rect 10529 886 10532 925
rect 10571 886 10574 925
rect 10625 886 10628 925
rect 10667 886 10670 925
rect 10721 887 10724 926
rect 10763 887 10766 926
rect 10241 726 10244 765
rect 10283 726 10286 765
rect 10337 725 10340 764
rect 10379 725 10382 764
rect 10433 725 10436 764
rect 10475 725 10478 764
rect 10529 725 10532 764
rect 10571 725 10574 764
rect 10625 725 10628 764
rect 10667 725 10670 764
rect 10721 726 10724 765
rect 10763 726 10766 765
rect 10241 565 10244 604
rect 10283 565 10286 604
rect 10337 564 10340 603
rect 10379 564 10382 603
rect 10433 564 10436 603
rect 10475 564 10478 603
rect 10529 564 10532 603
rect 10571 564 10574 603
rect 10625 564 10628 603
rect 10667 564 10670 603
rect 10721 565 10724 604
rect 10763 565 10766 604
rect 10241 404 10244 443
rect 10283 404 10286 443
rect 10337 403 10340 442
rect 10379 403 10382 442
rect 10433 403 10436 442
rect 10475 403 10478 442
rect 10529 403 10532 442
rect 10571 403 10574 442
rect 10625 403 10628 442
rect 10667 403 10670 442
rect 10721 404 10724 443
rect 10763 404 10766 443
rect 10241 243 10244 282
rect 10283 243 10286 282
rect 10337 243 10340 282
rect 10379 243 10382 282
rect 10433 243 10436 282
rect 10475 243 10478 282
rect 10529 243 10532 282
rect 10571 243 10574 282
rect 10625 243 10628 282
rect 10667 243 10670 282
rect 10721 243 10724 282
rect 10763 243 10766 282
<< nwell >>
rect 5401 5166 5404 5167
rect 3925 5152 4102 5163
rect 4489 5152 4739 5163
rect 5333 5136 5404 5166
rect 5333 5132 5401 5136
rect 5332 4527 5402 5132
rect 6379 4923 6380 5042
rect 6379 4918 6384 4923
rect 6379 4908 6385 4918
rect 6380 4796 6385 4908
rect 7722 4817 7778 4871
rect 5333 4507 5402 4527
rect 5332 2555 5507 3152
rect 5332 2552 5634 2555
rect 5546 2536 5634 2552
rect 5522 1839 5724 2408
rect 10786 227 10921 1774
rect 10785 180 10921 227
<< psubdiff >>
rect 668 6009 2470 6022
rect 668 5938 2040 6009
rect 2129 5938 2470 6009
rect 668 5931 2470 5938
rect 2379 2201 2470 5931
rect 6774 5704 8385 5709
rect 6774 5622 6787 5704
rect 6813 5703 8385 5704
rect 6813 5625 8120 5703
rect 8209 5625 8385 5703
rect 6813 5622 8385 5625
rect 6774 5618 8385 5622
rect 8294 3799 8385 5618
rect 2379 2167 2390 2201
rect 2407 2184 2424 2201
rect 2441 2184 2470 2201
rect 2458 2167 2470 2184
rect 2379 2149 2470 2167
rect 2379 2088 2393 2149
rect 2446 2088 2470 2149
rect 1813 1322 2064 1331
rect 1813 1280 1841 1322
rect 1814 970 1841 1280
rect 1858 970 1877 1322
rect 1894 970 1912 1322
rect 1929 970 1947 1322
rect 1964 970 1983 1322
rect 2000 970 2018 1322
rect 2035 970 2064 1322
rect 1814 957 2064 970
rect 2379 1038 2470 2088
rect 8045 3708 8385 3799
rect 8045 1038 8136 3708
rect 1814 956 1849 957
rect 2379 947 9537 1038
rect 2379 550 2470 947
<< nsubdiff >>
rect 10827 1743 10884 1751
rect 10827 1349 10840 1743
rect 10831 1289 10840 1349
rect 10827 1188 10840 1289
rect 10831 1128 10840 1188
rect 10827 1027 10840 1128
rect 10830 967 10840 1027
rect 10827 865 10840 967
rect 10831 805 10840 865
rect 10827 704 10840 805
rect 10830 644 10840 704
rect 10827 457 10840 644
rect 10830 248 10840 457
rect 10857 248 10884 1743
rect 10830 236 10884 248
<< psubdiffcont >>
rect 2040 5938 2129 6009
rect 6787 5622 6813 5704
rect 8120 5625 8209 5703
rect 2390 2184 2407 2201
rect 2424 2184 2441 2201
rect 2390 2167 2458 2184
rect 2393 2088 2446 2149
rect 1841 970 1858 1322
rect 1877 970 1894 1322
rect 1912 970 1929 1322
rect 1947 970 1964 1322
rect 1983 970 2000 1322
rect 2018 970 2035 1322
<< nsubdiffcont >>
rect 10840 248 10857 1743
<< locali >>
rect 1982 6014 2134 6015
rect 1982 6012 2137 6014
rect 1982 5938 1989 6012
rect 2032 6009 2137 6012
rect 2032 5938 2040 6009
rect 2129 5938 2137 6009
rect 1982 5935 2137 5938
rect 6779 5704 6846 5706
rect 6779 5622 6787 5704
rect 6813 5622 6818 5704
rect 6844 5622 6846 5704
rect 6779 5619 6846 5622
rect 8007 5704 8217 5706
rect 8007 5625 8013 5704
rect 8045 5703 8217 5704
rect 8045 5625 8120 5703
rect 8209 5625 8217 5703
rect 8007 5621 8217 5625
rect 2382 2167 2390 2201
rect 2421 2184 2424 2201
rect 2382 2159 2458 2167
rect 2384 2149 2458 2159
rect 2384 2088 2393 2149
rect 2446 2088 2458 2149
rect 2384 2080 2458 2088
rect 10840 1744 10877 1751
rect 10840 1743 10860 1744
rect 1817 1322 2056 1327
rect 1817 1290 1823 1322
rect 1822 970 1823 1290
rect 1840 970 1841 1322
rect 1858 970 1859 1322
rect 1876 970 1877 1322
rect 1894 970 1895 1322
rect 1929 970 1947 1322
rect 1981 970 1983 1322
rect 2017 970 2018 1322
rect 2035 970 2036 1322
rect 2053 970 2056 1322
rect 1822 964 2056 970
rect 1822 963 2055 964
rect 10857 249 10860 1743
rect 10877 249 10878 264
rect 10857 248 10878 249
rect 10840 239 10878 248
<< viali >>
rect 1989 5938 2032 6012
rect 6818 5622 6844 5704
rect 8013 5625 8045 5704
rect 2404 2184 2407 2201
rect 2407 2184 2421 2201
rect 2441 2184 2458 2201
rect 2404 2167 2421 2184
rect 2441 2167 2458 2184
rect 1823 970 1840 1322
rect 1859 970 1876 1322
rect 1895 970 1912 1322
rect 1964 970 1981 1322
rect 2000 970 2017 1322
rect 2036 970 2053 1322
rect 10860 249 10877 1744
<< metal1 >>
rect 8015 7404 8049 7418
rect 8803 7404 8875 7578
rect 8015 7332 8875 7404
rect 2808 7087 2942 7132
rect 198 7047 248 7051
rect 198 7008 203 7047
rect 242 7008 248 7047
rect 2808 7045 4160 7087
rect 4339 7078 4658 7190
rect 2808 7031 2942 7045
rect 198 7003 248 7008
rect 208 6707 247 7003
rect 2267 6971 2544 6995
rect 2267 6930 2291 6971
rect 208 6702 255 6707
rect 208 6663 211 6702
rect 250 6663 255 6702
rect 208 6658 255 6663
rect 208 6657 253 6658
rect 208 846 247 6657
rect 349 6572 375 6575
rect 349 6543 375 6546
rect 350 6321 374 6543
rect 341 6318 383 6321
rect 341 6273 383 6276
rect 930 6197 959 6389
rect 928 6194 969 6197
rect 928 6136 936 6194
rect 965 6136 969 6194
rect 928 6130 969 6136
rect 2266 6061 2290 6384
rect 2261 6056 2295 6061
rect 2261 6030 2265 6056
rect 2291 6030 2295 6056
rect 2261 6027 2295 6030
rect 1986 6017 2035 6018
rect 1985 6012 2036 6017
rect 1985 5938 1989 6012
rect 2032 5938 2036 6012
rect 1593 5148 1616 5496
rect 1660 5434 1682 5496
rect 1929 5468 1951 5923
rect 1985 5902 2036 5938
rect 2520 5924 2544 6971
rect 2851 6938 3154 6965
rect 3322 6939 3348 7045
rect 2848 6021 2879 6391
rect 2840 6018 2879 6021
rect 2840 5987 2844 6018
rect 2875 5987 2879 6018
rect 2840 5984 2879 5987
rect 3127 5970 3154 6938
rect 4118 6720 4160 7045
rect 4499 6796 4541 7078
rect 4499 6793 4546 6796
rect 4499 6751 4502 6793
rect 4544 6751 4546 6793
rect 4499 6748 4546 6751
rect 4114 6717 4162 6720
rect 4114 6675 4117 6717
rect 4159 6675 4162 6717
rect 4114 6672 4162 6675
rect 4669 6558 4713 6561
rect 4669 6511 4713 6514
rect 5241 6558 5285 6561
rect 5241 6511 5285 6514
rect 5420 6555 5493 7194
rect 5935 7179 6033 7194
rect 5420 6511 5423 6555
rect 5467 6511 5493 6555
rect 4227 6456 4271 6459
rect 4227 6409 4271 6412
rect 3244 6070 3269 6385
rect 3948 6136 3980 6140
rect 3948 6135 3951 6136
rect 3939 6110 3951 6135
rect 3977 6110 3980 6136
rect 3939 6106 3980 6110
rect 3240 6067 3273 6070
rect 3240 6041 3244 6067
rect 3270 6041 3273 6067
rect 3240 6034 3273 6041
rect 3123 5968 3157 5970
rect 3123 5942 3127 5968
rect 3154 5942 3157 5968
rect 3123 5939 3157 5942
rect 1980 5899 2036 5902
rect 1980 5892 1994 5899
rect 1969 5864 1994 5892
rect 2029 5864 2036 5899
rect 2515 5921 2549 5924
rect 2515 5895 2519 5921
rect 2545 5895 2549 5921
rect 2515 5892 2549 5895
rect 1969 5852 2036 5864
rect 1969 5849 2035 5852
rect 1969 5468 1991 5849
rect 3939 5756 3963 6106
rect 4233 5749 4264 6409
rect 4676 5751 4705 6511
rect 4795 6412 4798 6456
rect 4842 6412 4845 6456
rect 2091 5679 2126 5683
rect 2091 5640 2096 5679
rect 2122 5640 2126 5679
rect 2091 5637 2126 5640
rect 3734 5667 3771 5670
rect 3734 5641 3736 5667
rect 3769 5641 3771 5667
rect 3734 5639 3771 5641
rect 2031 5601 2056 5613
rect 2028 5598 2060 5601
rect 2028 5558 2032 5598
rect 2058 5558 2060 5598
rect 2028 5555 2060 5558
rect 2031 5476 2056 5555
rect 2031 5473 2060 5476
rect 2031 5447 2034 5473
rect 2031 5444 2060 5447
rect 1657 5431 1683 5434
rect 1657 5402 1683 5405
rect 1660 5342 1682 5402
rect 1654 5339 1682 5342
rect 1680 5313 1682 5339
rect 1654 5310 1682 5313
rect 1660 5250 1682 5310
rect 1655 5247 1682 5250
rect 1681 5221 1682 5247
rect 1655 5218 1682 5221
rect 1590 5145 1616 5148
rect 1590 5116 1616 5119
rect 1593 5052 1616 5116
rect 1586 5049 1616 5052
rect 1612 5023 1616 5049
rect 1586 5020 1616 5023
rect 1593 4956 1616 5020
rect 1590 4953 1616 4956
rect 1590 4924 1616 4927
rect 1593 3449 1616 4924
rect 1660 3449 1682 5218
rect 2031 5384 2056 5444
rect 2031 5381 2060 5384
rect 2031 5355 2034 5381
rect 2031 5352 2060 5355
rect 2031 5292 2056 5352
rect 2031 5289 2057 5292
rect 2031 5260 2057 5263
rect 1582 3446 1616 3449
rect 1582 3399 1586 3446
rect 1612 3399 1616 3446
rect 1582 3396 1616 3399
rect 1648 3446 1682 3449
rect 1648 3399 1650 3446
rect 1676 3399 1682 3446
rect 1648 3396 1682 3399
rect 1451 3322 1474 3329
rect 1447 3296 1450 3322
rect 1476 3296 1479 3322
rect 1402 3285 1425 3289
rect 1398 3282 1425 3285
rect 1424 3256 1425 3282
rect 1398 3253 1425 3256
rect 467 3197 539 3199
rect 467 3131 470 3197
rect 536 3131 539 3197
rect 467 3129 539 3131
rect 468 2614 534 3129
rect 1402 2901 1425 3253
rect 1451 3049 1474 3296
rect 1593 3287 1616 3396
rect 1660 3323 1682 3396
rect 1836 3325 1863 3329
rect 1658 3320 1684 3323
rect 1658 3291 1684 3294
rect 1834 3322 1863 3325
rect 1861 3295 1863 3322
rect 1834 3292 1863 3295
rect 1592 3284 1618 3287
rect 1592 3255 1618 3258
rect 1781 3138 1810 3141
rect 1451 3012 1524 3049
rect 1402 2894 1428 2901
rect 1400 2893 1428 2894
rect 1397 2891 1429 2893
rect 1397 2865 1400 2891
rect 1426 2865 1429 2891
rect 1397 2862 1429 2865
rect 987 2716 1030 2719
rect 987 2679 991 2716
rect 1028 2679 1030 2716
rect 987 2676 1030 2679
rect 468 2611 542 2614
rect 468 2545 474 2611
rect 540 2545 542 2611
rect 468 2542 542 2545
rect 992 2095 1029 2676
rect 1451 2262 1474 3012
rect 1836 2995 1863 3292
rect 1824 2970 1863 2995
rect 1884 3285 1908 3289
rect 1884 3282 1910 3285
rect 1884 3253 1910 3256
rect 1884 2939 1908 3253
rect 1824 2916 1908 2939
rect 1451 2239 1696 2262
rect 1664 2206 1696 2239
rect 988 2092 1031 2095
rect 988 2055 990 2092
rect 1027 2055 1031 2092
rect 988 2052 1031 2055
rect 1740 2049 1773 2052
rect 1726 2041 1744 2049
rect 1702 2017 1744 2041
rect 1740 2013 1744 2017
rect 1770 2013 1773 2049
rect 1740 2010 1773 2013
rect 1289 1518 1318 1521
rect 1289 1486 1318 1489
rect 1290 1429 1316 1486
rect 1884 1450 1908 2916
rect 1929 2849 1951 4924
rect 1969 3110 1991 4924
rect 2031 3225 2056 5260
rect 2093 5183 2119 5637
rect 3670 5502 3709 5504
rect 3670 5469 3673 5502
rect 3706 5469 3709 5502
rect 3670 5467 3709 5469
rect 3612 5354 3651 5357
rect 3612 5321 3616 5354
rect 3649 5321 3651 5354
rect 3612 5318 3651 5321
rect 3548 5194 3587 5197
rect 2093 5180 2121 5183
rect 2093 5154 2095 5180
rect 3548 5161 3552 5194
rect 3585 5161 3587 5194
rect 3548 5159 3587 5161
rect 2093 5151 2121 5154
rect 3551 5158 3585 5159
rect 2093 5087 2119 5151
rect 3487 5139 3521 5140
rect 3486 5137 3522 5139
rect 3486 5104 3488 5137
rect 3521 5104 3522 5137
rect 3486 5100 3522 5104
rect 2093 5084 2122 5087
rect 2093 5058 2096 5084
rect 2093 5055 2122 5058
rect 2093 4991 2119 5055
rect 2093 4988 2121 4991
rect 2093 4962 2095 4988
rect 2093 4959 2121 4962
rect 3425 4980 3461 4983
rect 2031 3223 2057 3225
rect 2030 3222 2058 3223
rect 2030 3196 2031 3222
rect 2057 3196 2058 3222
rect 2030 3195 2058 3196
rect 2031 3193 2057 3195
rect 1965 3107 1997 3110
rect 1965 3081 1969 3107
rect 1995 3081 1997 3107
rect 1965 3078 1997 3081
rect 1925 2846 1953 2849
rect 1925 2820 1927 2846
rect 1925 2817 1953 2820
rect 1929 1520 1951 2817
rect 1969 2296 1991 3078
rect 1969 2293 1998 2296
rect 1969 2251 1971 2293
rect 1997 2251 1998 2293
rect 1969 2248 1998 2251
rect 1969 2052 1991 2248
rect 1967 2049 1993 2052
rect 1967 2010 1993 2013
rect 1969 1548 1991 2010
rect 2031 1686 2056 3193
rect 2093 2792 2119 4959
rect 3425 4947 3427 4980
rect 3460 4947 3461 4980
rect 3425 4944 3461 4947
rect 3360 4827 3401 4830
rect 3360 4794 3364 4827
rect 3397 4794 3401 4827
rect 3360 4790 3401 4794
rect 3307 4670 3343 4673
rect 3307 4637 3308 4670
rect 3341 4637 3343 4670
rect 3307 4634 3343 4637
rect 3249 4128 3282 4130
rect 3243 4123 3282 4128
rect 3243 4090 3246 4123
rect 3279 4090 3282 4123
rect 3243 4086 3282 4090
rect 3186 3967 3219 3969
rect 3181 3964 3220 3967
rect 3181 3931 3183 3964
rect 3216 3931 3220 3964
rect 3181 3928 3220 3931
rect 3124 3812 3157 3813
rect 3121 3809 3157 3812
rect 3154 3776 3157 3809
rect 3121 3773 3157 3776
rect 3059 3661 3098 3665
rect 3059 3628 3061 3661
rect 3094 3628 3098 3661
rect 3059 3625 3098 3628
rect 2992 3144 3035 3148
rect 2992 3111 2997 3144
rect 3030 3111 3035 3144
rect 2992 3108 3035 3111
rect 2926 2987 2967 2991
rect 2926 2954 2930 2987
rect 2963 2954 2967 2987
rect 2926 2951 2967 2954
rect 2865 2823 2904 2827
rect 2092 2789 2123 2792
rect 2092 2763 2095 2789
rect 2121 2763 2123 2789
rect 2865 2790 2868 2823
rect 2901 2790 2904 2823
rect 2865 2787 2904 2790
rect 2092 2760 2123 2763
rect 2027 1683 2057 1686
rect 2027 1650 2029 1683
rect 2055 1650 2057 1683
rect 2027 1646 2057 1650
rect 1969 1534 1993 1548
rect 1925 1517 1956 1520
rect 1925 1488 1926 1517
rect 1955 1488 1956 1517
rect 1925 1485 1956 1488
rect 1970 1471 1993 1534
rect 1805 1447 1908 1450
rect 1805 1387 1810 1447
rect 1870 1394 1908 1447
rect 1969 1468 1993 1471
rect 1870 1387 1884 1394
rect 1805 1383 1884 1387
rect 1969 1329 1991 1468
rect 1816 1322 2058 1329
rect 1816 970 1823 1322
rect 1840 970 1859 1322
rect 1876 970 1895 1322
rect 1912 970 1964 1322
rect 1981 970 2000 1322
rect 2017 970 2036 1322
rect 2053 970 2058 1322
rect 1816 961 2058 970
rect 2093 932 2119 2760
rect 2796 2679 2837 2682
rect 2796 2646 2800 2679
rect 2833 2646 2837 2679
rect 2796 2643 2837 2646
rect 2375 2281 2468 2293
rect 2375 2210 2396 2281
rect 2454 2210 2468 2281
rect 2375 2201 2468 2210
rect 2375 2167 2404 2201
rect 2421 2167 2441 2201
rect 2458 2167 2468 2201
rect 2375 2128 2468 2167
rect 2384 2080 2458 2128
rect 2084 928 2119 932
rect 2084 894 2088 928
rect 2114 894 2119 928
rect 2084 891 2119 894
rect 191 839 247 846
rect 191 800 197 839
rect 236 800 247 839
rect 191 794 247 800
rect 2802 309 2835 2643
rect 2797 308 2840 309
rect 2794 306 2843 308
rect 2794 263 2797 306
rect 2840 263 2843 306
rect 2794 262 2843 263
rect 2797 260 2840 262
rect 2867 230 2900 2787
rect 2858 227 2907 230
rect 2858 184 2862 227
rect 2905 184 2907 227
rect 2858 181 2907 184
rect 2932 159 2965 2951
rect 2929 156 2969 159
rect 2929 113 2969 116
rect 2908 73 2966 75
rect 2908 22 2912 73
rect 2963 64 2966 73
rect 2999 64 3032 3108
rect 3063 522 3096 3625
rect 3063 76 3095 522
rect 3124 137 3157 3773
rect 3186 198 3219 3928
rect 3249 265 3282 4086
rect 3309 331 3342 4634
rect 3367 388 3400 4790
rect 3428 455 3461 4944
rect 3487 516 3520 5100
rect 3551 583 3584 5158
rect 3613 648 3646 5318
rect 3673 711 3706 5467
rect 3736 772 3769 5639
rect 3949 5152 3973 5163
rect 4243 5152 4274 5163
rect 4676 5148 4705 5164
rect 4822 5112 4841 6412
rect 5250 5108 5275 6511
rect 5420 6507 5493 6511
rect 5436 5468 5453 6507
rect 5936 6454 6033 7179
rect 7198 7077 7517 7189
rect 6475 6717 6622 6723
rect 6475 6675 6479 6717
rect 6614 6675 6622 6717
rect 6475 6670 6622 6675
rect 6238 6456 6282 6459
rect 5934 6452 6035 6454
rect 5934 6411 5937 6452
rect 6032 6411 6035 6452
rect 5934 6407 6035 6411
rect 6238 6409 6282 6412
rect 5658 6060 5692 6063
rect 5658 6034 5663 6060
rect 5689 6034 5692 6060
rect 5663 6031 5689 6034
rect 5475 5707 5501 5710
rect 5475 5678 5501 5681
rect 5478 5455 5497 5678
rect 5665 5453 5686 6031
rect 6022 5971 6048 5972
rect 6020 5969 6050 5971
rect 6020 5943 6022 5969
rect 6048 5943 6050 5969
rect 6020 5941 6050 5943
rect 6022 5940 6048 5941
rect 5705 5867 5739 5870
rect 5705 5841 5709 5867
rect 5735 5841 5739 5867
rect 5705 5838 5739 5841
rect 5712 5455 5731 5838
rect 5749 5658 5778 5661
rect 5749 5632 5751 5658
rect 5777 5632 5778 5658
rect 5749 5629 5778 5632
rect 5753 5453 5774 5629
rect 5853 5610 5887 5613
rect 5853 5584 5857 5610
rect 5883 5584 5887 5610
rect 5853 5581 5887 5584
rect 5861 5456 5879 5581
rect 6025 4917 6045 5940
rect 6248 5451 6271 6409
rect 6338 6061 6366 6064
rect 6338 6035 6339 6061
rect 6365 6035 6366 6061
rect 6338 6032 6366 6035
rect 6294 5970 6322 5973
rect 6294 5944 6295 5970
rect 6321 5944 6322 5970
rect 6294 5941 6322 5944
rect 6023 4904 6045 4917
rect 6018 4901 6051 4904
rect 6018 4874 6021 4901
rect 6048 4874 6051 4901
rect 6018 4871 6051 4874
rect 6271 4860 6272 4876
rect 6297 4787 6319 5941
rect 6296 4780 6319 4787
rect 6295 4720 6315 4780
rect 6340 4735 6363 6032
rect 6477 5432 6519 6670
rect 6580 5432 6622 6670
rect 6818 6452 6862 6455
rect 6818 6405 6862 6408
rect 6828 5707 6851 6405
rect 7270 5880 7398 7077
rect 7646 6558 7674 6570
rect 7646 6555 7679 6558
rect 7646 6511 7651 6555
rect 7646 6508 7679 6511
rect 7270 5872 7400 5880
rect 7269 5871 7400 5872
rect 7269 5845 7273 5871
rect 7395 5845 7400 5871
rect 7269 5842 7400 5845
rect 6947 5806 6977 5809
rect 6947 5780 6949 5806
rect 6975 5780 6977 5806
rect 6947 5777 6977 5780
rect 6815 5706 6851 5707
rect 6812 5704 6851 5706
rect 6812 5622 6818 5704
rect 6844 5622 6851 5704
rect 6812 5617 6851 5622
rect 6828 5451 6851 5617
rect 6950 5451 6973 5777
rect 7578 5752 7621 5756
rect 7578 5726 7582 5752
rect 7608 5726 7621 5752
rect 7578 5722 7621 5726
rect 7602 5455 7621 5722
rect 7646 5446 7674 6508
rect 7816 6061 7842 6064
rect 7816 6032 7842 6035
rect 7727 5974 7753 5977
rect 7727 5945 7753 5948
rect 7730 5573 7749 5945
rect 7818 5573 7840 6032
rect 8015 5710 8049 7332
rect 10055 7080 10374 7192
rect 8465 6986 8502 6987
rect 8460 6982 8510 6986
rect 8460 6945 8468 6982
rect 8505 6945 8510 6982
rect 8460 6941 8510 6945
rect 8080 6133 8112 6137
rect 8080 6106 8083 6133
rect 8109 6106 8112 6133
rect 8080 6100 8112 6106
rect 8010 5704 8049 5710
rect 8010 5702 8013 5704
rect 8009 5625 8013 5702
rect 8045 5625 8049 5704
rect 8010 5618 8049 5625
rect 7713 5553 7781 5573
rect 7713 5527 7727 5553
rect 7753 5527 7781 5553
rect 7713 5504 7781 5527
rect 7817 5554 7885 5573
rect 7817 5528 7829 5554
rect 7855 5528 7885 5554
rect 7817 5504 7885 5528
rect 8015 5440 8049 5618
rect 8082 5562 8109 6100
rect 8082 5559 8150 5562
rect 8082 5516 8104 5559
rect 8147 5516 8150 5559
rect 8082 5512 8150 5516
rect 8082 5447 8109 5512
rect 6296 4717 6319 4720
rect 3939 4111 3963 4548
rect 4233 4104 4264 4555
rect 4676 4106 4705 4553
rect 4822 4157 4841 4547
rect 4953 4167 4976 4551
rect 5250 4168 5275 4553
rect 6297 4397 6319 4717
rect 6297 4388 6332 4397
rect 6297 4366 6348 4388
rect 4820 4107 4841 4157
rect 4951 4126 4976 4167
rect 5248 4126 5275 4168
rect 5426 4183 5454 4294
rect 5479 4225 5498 4285
rect 5679 4241 5718 4243
rect 5678 4238 5718 4241
rect 5678 4232 5685 4238
rect 5663 4231 5685 4232
rect 5479 4206 5639 4225
rect 5426 4155 5598 4183
rect 5578 4132 5598 4155
rect 4820 4094 4839 4107
rect 4951 4083 4974 4126
rect 5248 4089 5273 4126
rect 5579 4102 5595 4132
rect 5620 4094 5639 4206
rect 5660 4210 5685 4231
rect 5713 4210 5718 4238
rect 5660 4207 5718 4210
rect 5660 4205 5717 4207
rect 5660 4204 5679 4205
rect 5660 4120 5677 4204
rect 6127 4198 6150 4289
rect 6249 4201 6272 4289
rect 6075 4191 6150 4198
rect 6072 4175 6150 4191
rect 6247 4195 6272 4201
rect 6580 4208 6622 4308
rect 6072 4130 6113 4175
rect 5660 4093 5676 4120
rect 6072 4081 6110 4130
rect 6247 4095 6271 4195
rect 6580 4190 6623 4208
rect 6580 4151 6624 4190
rect 6828 4169 6851 4289
rect 6583 4130 6624 4151
rect 6583 4079 6623 4130
rect 6827 4095 6851 4169
rect 6950 4200 6973 4289
rect 6950 4162 7026 4200
rect 7602 4187 7621 4285
rect 6988 4116 7026 4162
rect 7419 4179 7447 4182
rect 7419 4153 7420 4179
rect 7446 4153 7447 4179
rect 7419 4150 7447 4153
rect 7462 4168 7621 4187
rect 7422 4102 7438 4150
rect 7462 4135 7481 4168
rect 7646 4149 7674 4294
rect 8465 4250 8502 6941
rect 8544 6636 8590 6639
rect 8544 6599 8550 6636
rect 8587 6599 8590 6636
rect 8544 6596 8590 6599
rect 8462 4245 8507 4250
rect 8462 4208 8469 4245
rect 8506 4208 8507 4245
rect 8462 4204 8507 4208
rect 8465 4200 8502 4204
rect 8546 4191 8583 6596
rect 8621 6165 8666 6168
rect 8621 6128 8627 6165
rect 8664 6128 8666 6165
rect 8621 6125 8666 6128
rect 7507 4148 7674 4149
rect 7459 4124 7481 4135
rect 7459 4094 7478 4124
rect 7503 4121 7674 4148
rect 8543 4186 8587 4191
rect 8543 4149 8546 4186
rect 8583 4149 8587 4186
rect 8543 4145 8587 4149
rect 8546 4140 8583 4145
rect 7503 4102 7519 4121
rect 8623 3956 8660 6125
rect 9278 6073 9336 6076
rect 9278 6023 9282 6073
rect 9332 6023 9336 6073
rect 9278 6020 9336 6023
rect 9160 6013 9216 6017
rect 9052 5966 9108 5970
rect 8957 5917 9013 5928
rect 8957 5867 8960 5917
rect 9010 5867 9013 5917
rect 8957 5863 9013 5867
rect 9052 5916 9055 5966
rect 9105 5916 9108 5966
rect 9160 5963 9163 6013
rect 9213 5963 9216 6013
rect 9160 5958 9216 5963
rect 9052 5912 9108 5916
rect 8710 5658 8753 5661
rect 8710 5621 8715 5658
rect 8752 5621 8753 5658
rect 8710 5617 8753 5621
rect 8620 3955 8660 3956
rect 8619 3953 8661 3955
rect 8619 3916 8620 3953
rect 8657 3916 8661 3953
rect 8619 3913 8661 3916
rect 8623 3912 8660 3913
rect 3939 3449 3963 3535
rect 4233 3449 4264 3542
rect 3939 3158 3973 3449
rect 4233 3158 4274 3449
rect 4676 3158 4705 3540
rect 3949 3134 3973 3158
rect 4243 3131 4274 3158
rect 4822 3131 4841 3540
rect 4953 3436 4976 3544
rect 4944 3432 4977 3436
rect 4944 3391 4948 3432
rect 4974 3391 4977 3432
rect 4944 3388 4977 3391
rect 4953 3127 4976 3388
rect 5250 3148 5275 3546
rect 5582 3142 5598 3547
rect 5857 3183 5881 3555
rect 5855 3158 5894 3183
rect 5869 3133 5894 3158
rect 6075 3120 6113 3569
rect 6250 3181 6274 3555
rect 6250 3154 6297 3181
rect 6270 3131 6297 3154
rect 6478 3118 6518 3571
rect 6830 3304 6854 3555
rect 8711 3438 8748 5617
rect 8707 3432 8756 3438
rect 8707 3391 8713 3432
rect 8750 3391 8756 3432
rect 8707 3387 8756 3391
rect 8711 3384 8748 3387
rect 6830 3280 6888 3304
rect 6864 3146 6888 3280
rect 5385 3045 5417 3049
rect 5385 3019 5388 3045
rect 5414 3019 5417 3045
rect 7376 3043 7402 3046
rect 5385 3015 5417 3019
rect 7375 3017 7376 3040
rect 3939 1295 3963 2558
rect 4233 2450 4264 2565
rect 4676 2501 4705 2563
rect 4726 2532 4760 2535
rect 4726 2506 4730 2532
rect 4756 2506 4760 2532
rect 4726 2503 4760 2506
rect 4673 2498 4708 2501
rect 4673 2469 4676 2498
rect 4705 2469 4708 2498
rect 4673 2466 4708 2469
rect 4229 2449 4266 2450
rect 4229 2418 4232 2449
rect 4263 2418 4266 2449
rect 4676 2420 4705 2466
rect 4726 2442 4751 2503
rect 4822 2444 4841 2564
rect 5250 2497 5275 2570
rect 5393 2539 5414 3015
rect 7375 3014 7402 3017
rect 7324 2950 7350 2953
rect 7324 2921 7350 2924
rect 5519 2846 5558 2871
rect 5447 2767 5481 2770
rect 5447 2741 5451 2767
rect 5477 2741 5481 2767
rect 5447 2736 5481 2741
rect 5451 2734 5473 2736
rect 5390 2536 5418 2539
rect 5390 2510 5391 2536
rect 5417 2510 5418 2536
rect 5390 2507 5418 2510
rect 5451 2506 5471 2734
rect 5497 2552 5516 2588
rect 5493 2535 5521 2552
rect 5493 2509 5494 2535
rect 5520 2509 5521 2535
rect 5447 2503 5475 2506
rect 5493 2505 5521 2509
rect 5247 2495 5281 2497
rect 5247 2469 5251 2495
rect 5277 2469 5281 2495
rect 5447 2477 5448 2503
rect 5474 2477 5475 2503
rect 5447 2474 5475 2477
rect 5247 2468 5281 2469
rect 4229 2417 4266 2418
rect 4233 2296 4264 2417
rect 4619 2392 4705 2420
rect 4611 2391 4705 2392
rect 4721 2431 4751 2442
rect 4816 2441 4848 2444
rect 4611 2389 4657 2391
rect 4611 2347 4613 2389
rect 4655 2347 4657 2389
rect 4611 2344 4657 2347
rect 4228 2293 4270 2296
rect 4721 2280 4740 2431
rect 4816 2415 4819 2441
rect 4845 2415 4848 2441
rect 4816 2412 4848 2415
rect 5084 2391 5159 2410
rect 5109 2307 5159 2391
rect 5540 2383 5558 2846
rect 7277 2766 7303 2769
rect 7277 2737 7303 2740
rect 7227 2673 7253 2676
rect 7227 2644 7253 2647
rect 5672 2499 5698 2502
rect 5670 2497 5700 2499
rect 5670 2471 5672 2497
rect 5698 2471 5700 2497
rect 5670 2469 5700 2471
rect 5672 2468 5698 2469
rect 5540 2379 5588 2383
rect 5540 2353 5552 2379
rect 5548 2346 5552 2353
rect 5585 2346 5588 2379
rect 5673 2376 5695 2468
rect 5869 2455 5894 2578
rect 6270 2457 6297 2580
rect 6552 2537 6595 2540
rect 6552 2502 6556 2537
rect 6591 2502 6595 2537
rect 6552 2500 6595 2502
rect 5868 2429 5871 2455
rect 5897 2429 5900 2455
rect 6270 2453 6305 2457
rect 6270 2426 6275 2453
rect 6302 2426 6305 2453
rect 5548 2342 5588 2346
rect 5667 2373 5701 2376
rect 5667 2336 5701 2339
rect 5673 2328 5695 2336
rect 6068 2309 6162 2402
rect 6556 2357 6591 2500
rect 6738 2444 6760 2576
rect 6864 2504 6887 2576
rect 6864 2481 7185 2504
rect 6864 2480 6887 2481
rect 6556 2325 6560 2357
rect 6586 2325 6591 2357
rect 6556 2321 6591 2325
rect 6709 2420 6760 2444
rect 4228 2248 4270 2251
rect 4677 2274 4740 2280
rect 5060 2275 5084 2307
rect 5184 2275 5208 2307
rect 6041 2277 6065 2309
rect 6165 2277 6189 2309
rect 6709 2295 6732 2420
rect 7162 2384 7185 2481
rect 7157 2381 7188 2384
rect 7157 2347 7159 2381
rect 7185 2347 7188 2381
rect 7157 2344 7188 2347
rect 6698 2292 6744 2295
rect 4677 2242 4681 2274
rect 4713 2248 4740 2274
rect 6698 2254 6702 2292
rect 6740 2254 6744 2292
rect 6698 2251 6744 2254
rect 4713 2242 4721 2248
rect 4677 2238 4721 2242
rect 5060 2141 5084 2173
rect 5184 2140 5208 2172
rect 6041 2143 6065 2175
rect 6165 2142 6189 2174
rect 7162 2027 7185 2344
rect 7149 2005 7185 2027
rect 7129 1982 7185 2005
rect 7129 1981 7183 1982
rect 4698 1720 4730 1895
rect 5060 1864 5084 1896
rect 5184 1863 5208 1895
rect 5084 1798 5110 1844
rect 5158 1800 5184 1844
rect 5083 1795 5111 1798
rect 5083 1764 5111 1767
rect 5157 1797 5185 1800
rect 5157 1766 5185 1769
rect 4686 1710 4740 1720
rect 4686 1664 4691 1710
rect 4737 1664 4740 1710
rect 4686 1660 4740 1664
rect 5084 1623 5110 1764
rect 5158 1623 5184 1766
rect 3899 1278 3964 1295
rect 5084 1280 5184 1623
rect 5535 1618 5569 1897
rect 5529 1615 5575 1618
rect 5529 1566 5575 1569
rect 5678 1529 5712 1896
rect 6041 1866 6065 1898
rect 6165 1866 6189 1898
rect 6065 1798 6091 1847
rect 6064 1795 6092 1798
rect 6064 1764 6092 1767
rect 6065 1646 6091 1764
rect 6139 1646 6165 1847
rect 5669 1526 5721 1529
rect 5669 1480 5672 1526
rect 5718 1480 5721 1526
rect 5669 1477 5721 1480
rect 6065 1286 6165 1646
rect 6520 1441 6547 1900
rect 7227 1860 7252 2644
rect 7277 1950 7302 2737
rect 7325 2041 7350 2921
rect 7375 2130 7400 3014
rect 8959 2280 9009 5863
rect 9052 2808 9102 5912
rect 9165 3331 9215 5958
rect 9278 3848 9328 6020
rect 10164 5860 10292 7080
rect 10163 5857 10292 5860
rect 10291 5729 10292 5857
rect 10163 5726 10292 5729
rect 10164 5677 10292 5726
rect 10600 5559 10620 5562
rect 10591 5556 10622 5559
rect 10591 5513 10595 5556
rect 10621 5513 10622 5556
rect 10591 5509 10622 5513
rect 10209 5427 10244 5430
rect 10209 5385 10212 5427
rect 10238 5385 10244 5427
rect 10209 5382 10244 5385
rect 9810 5105 9857 5111
rect 9810 5065 9812 5105
rect 9852 5065 9857 5105
rect 9810 5062 9857 5065
rect 9273 3845 9328 3848
rect 9323 3795 9328 3845
rect 9273 3792 9328 3795
rect 9164 3323 9216 3331
rect 9164 3276 9165 3323
rect 9215 3276 9216 3323
rect 9164 3275 9216 3276
rect 9051 2807 9103 2808
rect 9051 2757 9052 2807
rect 9102 2757 9103 2807
rect 9051 2756 9103 2757
rect 8943 2277 9009 2280
rect 8943 2227 8947 2277
rect 8997 2227 9009 2277
rect 8943 2223 9009 2227
rect 7370 2126 7407 2130
rect 7370 2076 7374 2126
rect 7400 2076 7407 2126
rect 7370 2072 7407 2076
rect 7317 2036 7354 2041
rect 7317 1986 7320 2036
rect 7346 1986 7354 2036
rect 7317 1983 7354 1986
rect 7268 1946 7305 1950
rect 7268 1896 7273 1946
rect 7299 1896 7305 1946
rect 7268 1892 7305 1896
rect 7221 1856 7256 1860
rect 6509 1435 6558 1441
rect 6509 1389 6511 1435
rect 6557 1389 6558 1435
rect 6509 1385 6558 1389
rect 6065 1282 6267 1286
rect 3899 1166 3904 1278
rect 3930 1166 3964 1278
rect 5036 1276 5229 1280
rect 3899 1163 3964 1166
rect 4982 1274 5229 1276
rect 4982 1272 5115 1274
rect 4982 1160 5041 1272
rect 5227 1162 5229 1274
rect 5153 1160 5229 1162
rect 4982 1157 5229 1160
rect 6017 1276 6267 1282
rect 6017 1157 6022 1276
rect 6208 1157 6267 1276
rect 3734 770 3771 772
rect 3734 737 3736 770
rect 3769 737 3771 770
rect 3734 734 3771 737
rect 3669 708 3708 711
rect 3669 675 3674 708
rect 3707 675 3708 708
rect 3669 672 3708 675
rect 3609 645 3647 648
rect 3609 612 3611 645
rect 3644 612 3647 645
rect 3609 609 3647 612
rect 3550 582 3585 583
rect 3550 549 3551 582
rect 3584 549 3585 582
rect 3550 546 3585 549
rect 3486 514 3522 516
rect 3486 481 3487 514
rect 3520 481 3522 514
rect 3486 478 3522 481
rect 3427 454 3461 455
rect 3425 452 3463 454
rect 3425 419 3427 452
rect 3460 419 3463 452
rect 3425 417 3463 419
rect 3427 416 3460 417
rect 3367 352 3400 355
rect 3309 295 3342 298
rect 3249 262 3284 265
rect 3249 232 3251 262
rect 3251 226 3284 229
rect 3186 162 3219 165
rect 3122 134 3157 137
rect 3155 104 3157 134
rect 3122 97 3155 100
rect 2963 31 3032 64
rect 3061 73 3105 76
rect 3061 36 3064 73
rect 3101 36 3105 73
rect 3061 34 3105 36
rect 2963 22 2966 31
rect 2908 20 2966 22
rect 4982 8 5076 1157
rect 6017 1154 6267 1157
rect 6178 154 6267 1154
rect 7094 839 7127 1838
rect 7221 1806 7225 1856
rect 7251 1806 7256 1856
rect 7221 1803 7256 1806
rect 8959 1441 9009 2223
rect 9052 1532 9102 2756
rect 9165 1619 9215 3275
rect 9278 1721 9328 3792
rect 9567 2529 9625 2533
rect 9567 2479 9571 2529
rect 9621 2479 9625 2529
rect 9567 2477 9625 2479
rect 9570 2476 9621 2477
rect 9278 1718 9334 1721
rect 9278 1668 9284 1718
rect 9278 1665 9334 1668
rect 9278 1652 9328 1665
rect 9165 1570 9215 1573
rect 9052 1483 9102 1486
rect 8959 1392 9009 1395
rect 9570 1289 9620 2476
rect 9507 1278 9620 1289
rect 9507 1166 9513 1278
rect 9607 1166 9620 1278
rect 9507 1161 9620 1166
rect 7088 836 7131 839
rect 7088 803 7092 836
rect 7125 803 7131 836
rect 7088 800 7131 803
rect 9815 727 9855 5062
rect 9907 5001 9910 5037
rect 9946 5001 9949 5037
rect 9814 724 9861 727
rect 9814 684 9818 724
rect 9858 684 9861 724
rect 9814 681 9861 684
rect 9908 647 9947 5001
rect 9999 4803 10044 4805
rect 9999 4764 10002 4803
rect 10041 4764 10044 4803
rect 9999 4762 10044 4764
rect 9905 643 9951 647
rect 9905 604 9909 643
rect 9948 604 9951 643
rect 9905 600 9951 604
rect 10001 565 10040 4762
rect 10085 4736 10123 4737
rect 10083 4734 10125 4736
rect 10083 4708 10085 4734
rect 10123 4708 10125 4734
rect 10083 4706 10125 4708
rect 9999 561 10046 565
rect 9999 522 10002 561
rect 10041 522 10046 561
rect 9999 519 10046 522
rect 10085 485 10123 4706
rect 10219 2383 10242 5382
rect 10600 5184 10620 5509
rect 10951 5185 10970 7212
rect 11285 6333 11367 6336
rect 11285 6327 11290 6333
rect 11279 6262 11290 6327
rect 11361 6262 11367 6333
rect 11279 6258 11367 6262
rect 11279 4358 11350 6258
rect 11266 4354 11350 4358
rect 11266 4283 11271 4354
rect 11342 4283 11350 4354
rect 11266 4279 11350 4283
rect 10838 2529 10910 2532
rect 10838 2478 10851 2529
rect 10902 2478 10910 2529
rect 10838 2475 10910 2478
rect 10219 2360 10243 2383
rect 10219 1779 10242 2360
rect 10844 1774 10895 2475
rect 10830 1769 10895 1774
rect 10829 1751 10895 1769
rect 10826 1750 10895 1751
rect 10826 1744 10886 1750
rect 10826 1526 10860 1744
rect 10791 1427 10860 1526
rect 10826 1349 10860 1427
rect 10831 1289 10860 1349
rect 10827 1288 10860 1289
rect 10826 1188 10860 1288
rect 10831 1128 10860 1188
rect 10826 1027 10860 1128
rect 10830 967 10860 1027
rect 10826 865 10860 967
rect 10831 805 10860 865
rect 10826 704 10860 805
rect 10830 644 10860 704
rect 10082 481 10126 485
rect 10082 443 10084 481
rect 10122 443 10126 481
rect 10826 457 10860 644
rect 10082 439 10126 443
rect 10830 249 10860 457
rect 10877 1713 10886 1744
rect 10877 249 10884 1713
rect 10830 236 10884 249
rect 6178 81 6270 154
rect 6175 8 6267 81
<< via1 >>
rect 203 7008 242 7047
rect 211 6663 250 6702
rect 349 6546 375 6572
rect 341 6276 383 6318
rect 936 6136 965 6194
rect 2265 6030 2291 6056
rect 2844 5987 2875 6018
rect 4502 6751 4544 6793
rect 4117 6675 4159 6717
rect 4669 6514 4713 6558
rect 5241 6514 5285 6558
rect 5423 6511 5467 6555
rect 4227 6412 4271 6456
rect 3951 6110 3977 6136
rect 3244 6041 3270 6067
rect 3127 5942 3154 5968
rect 1994 5864 2029 5899
rect 2519 5895 2545 5921
rect 4798 6412 4842 6456
rect 2096 5640 2122 5679
rect 3736 5641 3769 5667
rect 2032 5558 2058 5598
rect 2034 5447 2060 5473
rect 1657 5405 1683 5431
rect 1654 5313 1680 5339
rect 1655 5221 1681 5247
rect 1590 5119 1616 5145
rect 1586 5023 1612 5049
rect 1590 4927 1616 4953
rect 2034 5355 2060 5381
rect 2031 5263 2057 5289
rect 1586 3399 1612 3446
rect 1650 3399 1676 3446
rect 1450 3296 1476 3322
rect 1398 3256 1424 3282
rect 470 3131 536 3197
rect 1658 3294 1684 3320
rect 1834 3295 1861 3322
rect 1592 3258 1618 3284
rect 1400 2865 1426 2891
rect 991 2679 1028 2716
rect 474 2545 540 2611
rect 1884 3256 1910 3282
rect 990 2055 1027 2092
rect 1744 2013 1770 2049
rect 1289 1489 1318 1518
rect 3673 5469 3706 5502
rect 3616 5321 3649 5354
rect 2095 5154 2121 5180
rect 3552 5161 3585 5194
rect 3488 5104 3521 5137
rect 2096 5058 2122 5084
rect 2095 4962 2121 4988
rect 2031 3196 2057 3222
rect 1969 3081 1995 3107
rect 1927 2820 1953 2846
rect 1971 2251 1997 2293
rect 1967 2013 1993 2049
rect 3427 4947 3460 4980
rect 3364 4794 3397 4827
rect 3308 4637 3341 4670
rect 3246 4090 3279 4123
rect 3183 3931 3216 3964
rect 3121 3776 3154 3809
rect 3061 3628 3094 3661
rect 2997 3111 3030 3144
rect 2930 2954 2963 2987
rect 2095 2763 2121 2789
rect 2868 2790 2901 2823
rect 2029 1650 2055 1683
rect 1926 1488 1955 1517
rect 1810 1387 1870 1447
rect 2800 2646 2833 2679
rect 2396 2210 2454 2281
rect 2088 894 2114 928
rect 197 800 236 839
rect 2797 263 2840 306
rect 2862 184 2905 227
rect 2929 116 2969 156
rect 2912 22 2963 73
rect 6479 6675 6614 6717
rect 5937 6411 6032 6452
rect 6238 6412 6282 6456
rect 5663 6034 5689 6060
rect 5475 5681 5501 5707
rect 6022 5943 6048 5969
rect 5709 5841 5735 5867
rect 5751 5632 5777 5658
rect 5857 5584 5883 5610
rect 6339 6035 6365 6061
rect 6295 5944 6321 5970
rect 6021 4874 6048 4901
rect 6818 6408 6862 6452
rect 7651 6511 7679 6555
rect 7273 5845 7395 5871
rect 6949 5780 6975 5806
rect 7582 5726 7608 5752
rect 7816 6035 7842 6061
rect 7727 5948 7753 5974
rect 8468 6945 8505 6982
rect 8083 6106 8109 6133
rect 7727 5527 7753 5553
rect 7829 5528 7855 5554
rect 8104 5516 8147 5559
rect 5685 4210 5713 4238
rect 7420 4153 7446 4179
rect 8550 6599 8587 6636
rect 8469 4208 8506 4245
rect 8627 6128 8664 6165
rect 8546 4149 8583 4186
rect 9282 6023 9332 6073
rect 8960 5867 9010 5917
rect 9055 5916 9105 5966
rect 9163 5963 9213 6013
rect 8715 5621 8752 5658
rect 8620 3916 8657 3953
rect 4948 3391 4974 3432
rect 8713 3391 8750 3432
rect 5388 3019 5414 3045
rect 7376 3017 7402 3043
rect 4730 2506 4756 2532
rect 4676 2469 4705 2498
rect 4232 2418 4263 2449
rect 7324 2924 7350 2950
rect 5451 2741 5477 2767
rect 5391 2510 5417 2536
rect 5494 2509 5520 2535
rect 5251 2469 5277 2495
rect 5448 2477 5474 2503
rect 4613 2347 4655 2389
rect 4228 2251 4270 2293
rect 4819 2415 4845 2441
rect 7277 2740 7303 2766
rect 7227 2647 7253 2673
rect 5672 2471 5698 2497
rect 5552 2346 5585 2379
rect 6556 2502 6591 2537
rect 5871 2429 5897 2455
rect 6275 2426 6302 2453
rect 5667 2339 5701 2373
rect 6560 2325 6586 2357
rect 7159 2347 7185 2381
rect 4681 2242 4713 2274
rect 6702 2254 6740 2292
rect 5083 1767 5111 1795
rect 5157 1769 5185 1797
rect 4691 1664 4737 1710
rect 5529 1569 5575 1615
rect 6064 1767 6092 1795
rect 5672 1480 5718 1526
rect 10163 5729 10291 5857
rect 10595 5513 10621 5556
rect 10212 5385 10238 5427
rect 9812 5065 9852 5105
rect 9273 3795 9323 3845
rect 9165 3276 9215 3323
rect 9052 2757 9102 2807
rect 8947 2227 8997 2277
rect 7374 2076 7400 2126
rect 7320 1986 7346 2036
rect 7273 1896 7299 1946
rect 6511 1389 6557 1435
rect 3904 1166 3930 1278
rect 5115 1272 5227 1274
rect 5041 1162 5227 1272
rect 5041 1160 5153 1162
rect 6022 1157 6208 1276
rect 3736 737 3769 770
rect 3674 675 3707 708
rect 3611 612 3644 645
rect 3551 549 3584 582
rect 3487 481 3520 514
rect 3427 419 3460 452
rect 3367 355 3400 388
rect 3309 298 3342 331
rect 3251 229 3284 262
rect 3186 165 3219 198
rect 3122 100 3155 134
rect 3064 36 3101 73
rect 7225 1806 7251 1856
rect 9571 2479 9621 2529
rect 9284 1668 9334 1718
rect 9165 1573 9215 1619
rect 9052 1486 9102 1532
rect 8959 1395 9009 1441
rect 9513 1166 9607 1278
rect 7092 803 7125 836
rect 9910 5001 9946 5037
rect 9818 684 9858 724
rect 10002 4764 10041 4803
rect 9909 604 9948 643
rect 10085 4708 10123 4734
rect 10002 522 10041 561
rect 11290 6262 11361 6333
rect 11271 4283 11342 4354
rect 10851 2478 10902 2529
rect 10084 443 10122 481
<< metal2 >>
rect 77 7039 145 7161
rect 200 7047 245 7049
rect 200 7039 203 7047
rect 77 7016 203 7039
rect 77 6929 145 7016
rect 200 7008 203 7016
rect 242 7008 245 7047
rect 200 7006 245 7008
rect 8462 6982 8508 6984
rect 11549 6982 11635 7117
rect 8462 6945 8468 6982
rect 8505 6945 11635 6982
rect 8462 6943 8508 6945
rect 11549 6907 11635 6945
rect 62 6819 310 6820
rect 62 6780 457 6819
rect 289 6743 457 6780
rect 2055 6810 2130 6811
rect 2055 6780 2217 6810
rect 4500 6793 4545 6795
rect 4499 6787 4502 6793
rect 2055 6763 2079 6780
rect 2187 6758 2217 6780
rect 2260 6757 4502 6787
rect 4499 6751 4502 6757
rect 4544 6751 4547 6793
rect 4500 6749 4545 6751
rect 4115 6717 4160 6719
rect 6476 6717 6618 6720
rect 77 6620 145 6708
rect 210 6702 253 6706
rect 210 6663 211 6702
rect 250 6663 253 6702
rect 4114 6675 4117 6717
rect 4159 6716 4162 6717
rect 6476 6716 6479 6717
rect 4159 6676 6479 6716
rect 4159 6675 4162 6676
rect 6476 6675 6479 6676
rect 6614 6716 6618 6717
rect 6614 6676 6623 6716
rect 6614 6675 6618 6676
rect 4115 6673 4160 6675
rect 6476 6672 6618 6675
rect 210 6659 253 6663
rect 210 6658 404 6659
rect 219 6636 404 6658
rect 8545 6636 8589 6638
rect 11549 6636 11635 6704
rect 77 6588 413 6620
rect 8545 6599 8550 6636
rect 8587 6599 11635 6636
rect 8545 6597 8589 6599
rect 77 6476 145 6588
rect 346 6546 349 6572
rect 375 6549 404 6572
rect 375 6546 378 6549
rect 4666 6514 4669 6558
rect 4713 6555 4716 6558
rect 5238 6555 5241 6558
rect 4713 6514 5241 6555
rect 5285 6555 5288 6558
rect 5285 6514 5423 6555
rect 4681 6511 5423 6514
rect 5467 6511 7651 6555
rect 7679 6511 7682 6555
rect 11549 6494 11635 6599
rect 4798 6456 4842 6459
rect 277 6439 430 6455
rect 96 6406 430 6439
rect 4224 6412 4227 6456
rect 4271 6454 4274 6456
rect 4271 6412 4798 6454
rect 6235 6454 6238 6456
rect 4842 6452 6238 6454
rect 4842 6412 5937 6452
rect 4239 6411 5937 6412
rect 6032 6412 6238 6452
rect 6282 6454 6285 6456
rect 6282 6452 6875 6454
rect 6282 6412 6818 6452
rect 6032 6411 6818 6412
rect 4239 6410 6818 6411
rect 4798 6409 4842 6410
rect 6815 6408 6818 6410
rect 6862 6410 6875 6452
rect 6862 6408 6865 6410
rect 96 6399 323 6406
rect 96 6379 136 6399
rect 61 6339 136 6379
rect 11287 6318 11290 6333
rect 338 6276 341 6318
rect 383 6276 11290 6318
rect 11287 6262 11290 6276
rect 11361 6262 11364 6333
rect 32 6194 100 6261
rect 924 6194 971 6196
rect 32 6136 936 6194
rect 965 6136 971 6194
rect 8623 6165 8665 6167
rect 11546 6165 11632 6295
rect 32 6112 104 6136
rect 924 6134 971 6136
rect 3949 6136 3979 6139
rect 32 6029 100 6112
rect 3949 6110 3951 6136
rect 3977 6133 3979 6136
rect 8081 6133 8111 6136
rect 3977 6110 8083 6133
rect 3949 6107 3979 6110
rect 8081 6106 8083 6110
rect 8109 6110 8118 6133
rect 8623 6128 8627 6165
rect 8664 6128 11632 6165
rect 8623 6126 8665 6128
rect 8109 6106 8111 6110
rect 8081 6102 8111 6106
rect 11546 6085 11632 6128
rect 3241 6067 3272 6069
rect 2262 6059 2294 6060
rect 3241 6059 3244 6067
rect 2262 6056 3244 6059
rect 2262 6030 2265 6056
rect 2291 6041 3244 6056
rect 3270 6059 3273 6067
rect 5659 6060 5691 6062
rect 6336 6061 6368 6062
rect 5659 6059 5663 6060
rect 3270 6041 5663 6059
rect 2291 6036 5663 6041
rect 2291 6030 2294 6036
rect 3241 6035 3272 6036
rect 5659 6034 5663 6036
rect 5689 6059 5692 6060
rect 6336 6059 6339 6061
rect 5689 6036 6339 6059
rect 5689 6034 5692 6036
rect 6336 6035 6339 6036
rect 6365 6059 6368 6061
rect 7813 6059 7816 6061
rect 6365 6036 7816 6059
rect 6365 6035 6368 6036
rect 7813 6035 7816 6036
rect 7842 6059 7845 6061
rect 9279 6059 9282 6073
rect 7842 6036 9282 6059
rect 7842 6035 7845 6036
rect 6336 6034 6368 6035
rect 2262 6028 2294 6030
rect 9279 6023 9282 6036
rect 9332 6023 9335 6073
rect 9279 6022 9335 6023
rect 2841 6018 2878 6020
rect 32 5979 83 5991
rect 2841 5987 2844 6018
rect 2875 6014 2878 6018
rect 9161 6014 9215 6016
rect 2875 6013 9215 6014
rect 2875 5991 9163 6013
rect 2875 5987 2878 5991
rect 2841 5985 2878 5987
rect 32 5950 342 5979
rect 6292 5970 6324 5971
rect 6021 5969 6049 5970
rect 83 5949 342 5950
rect 3124 5968 3155 5969
rect 6019 5968 6022 5969
rect 3124 5942 3127 5968
rect 3154 5945 6022 5968
rect 3154 5942 3157 5945
rect 6019 5943 6022 5945
rect 6048 5968 6051 5969
rect 6292 5968 6295 5970
rect 6048 5945 6295 5968
rect 6048 5943 6051 5945
rect 6292 5944 6295 5945
rect 6321 5968 6324 5970
rect 7724 5968 7727 5974
rect 6321 5948 7727 5968
rect 7753 5968 7756 5974
rect 9053 5968 9107 5969
rect 7753 5966 9107 5968
rect 7753 5948 9055 5966
rect 6321 5945 9055 5948
rect 6321 5944 6324 5945
rect 6292 5943 6324 5944
rect 6021 5942 6049 5943
rect 3124 5940 3155 5942
rect 2516 5922 2548 5923
rect 8959 5922 9012 5925
rect 2516 5921 9012 5922
rect 28 5899 79 5901
rect 1992 5899 2032 5900
rect 28 5864 1994 5899
rect 2029 5864 2032 5899
rect 2516 5895 2519 5921
rect 2545 5917 9012 5921
rect 2545 5899 8960 5917
rect 2545 5895 2548 5899
rect 2516 5893 2548 5895
rect 7271 5871 7399 5874
rect 28 5860 79 5864
rect 1992 5861 2032 5864
rect 5706 5867 5738 5868
rect 5706 5841 5709 5867
rect 5735 5864 5738 5867
rect 7271 5864 7273 5871
rect 5735 5845 7273 5864
rect 7395 5845 7399 5871
rect 8959 5867 8960 5899
rect 9010 5867 9012 5917
rect 9053 5916 9055 5945
rect 9105 5916 9107 5966
rect 9161 5963 9163 5991
rect 9213 5963 9215 6013
rect 9161 5960 9215 5963
rect 9053 5913 9107 5916
rect 8959 5864 9012 5867
rect 5735 5843 7399 5845
rect 5735 5841 5738 5843
rect 5706 5840 5738 5841
rect 0 5679 127 5825
rect 4712 5799 4997 5819
rect 6948 5806 6976 5808
rect 4977 5749 4997 5799
rect 6946 5780 6949 5806
rect 6975 5803 6978 5806
rect 10160 5803 10163 5857
rect 6975 5782 10163 5803
rect 6975 5780 6978 5782
rect 6948 5778 6976 5780
rect 7579 5752 7610 5755
rect 7579 5749 7582 5752
rect 3830 5714 3886 5731
rect 4977 5729 7582 5749
rect 7579 5726 7582 5729
rect 7608 5726 7610 5752
rect 10160 5729 10163 5782
rect 10291 5729 10294 5857
rect 7579 5723 7610 5726
rect 1135 5679 1165 5680
rect 2094 5679 2123 5681
rect 0 5640 2096 5679
rect 2122 5640 2126 5679
rect 3733 5641 3736 5667
rect 3769 5658 3772 5667
rect 3830 5658 3847 5714
rect 5472 5702 5475 5707
rect 4972 5682 5475 5702
rect 3769 5641 3848 5658
rect 4972 5644 4992 5682
rect 5472 5681 5475 5682
rect 5501 5702 5504 5707
rect 5501 5682 5509 5702
rect 5501 5681 5504 5682
rect 5748 5658 5779 5659
rect 8711 5658 8754 5660
rect 11546 5658 11632 5856
rect 5748 5655 5751 5658
rect 0 5637 127 5640
rect 2094 5638 2123 5640
rect 4712 5624 4992 5644
rect 5023 5635 5751 5655
rect 2030 5598 2059 5600
rect 785 5558 2032 5598
rect 2058 5558 2061 5598
rect 29 5289 156 5376
rect 785 5289 825 5558
rect 2030 5557 2059 5558
rect 3830 5531 3886 5548
rect 3673 5504 3706 5505
rect 3671 5502 3708 5504
rect 1165 5490 1202 5491
rect 986 5467 1202 5490
rect 2031 5468 2034 5473
rect 986 5454 1728 5467
rect 986 5384 1048 5454
rect 1165 5450 1728 5454
rect 1974 5451 2034 5468
rect 2031 5447 2034 5451
rect 2060 5468 2063 5473
rect 3671 5469 3673 5502
rect 3706 5494 3708 5502
rect 3830 5494 3847 5531
rect 3706 5477 3847 5494
rect 3706 5469 3708 5477
rect 3830 5476 3847 5477
rect 5023 5469 5043 5635
rect 5748 5632 5751 5635
rect 5777 5632 5780 5658
rect 5748 5631 5779 5632
rect 8711 5621 8715 5658
rect 8752 5646 11632 5658
rect 8752 5621 11621 5646
rect 8711 5618 8752 5621
rect 5854 5610 5886 5611
rect 5854 5607 5857 5610
rect 2060 5451 2069 5468
rect 3671 5466 3708 5469
rect 2060 5447 2063 5451
rect 4712 5449 5043 5469
rect 5078 5587 5857 5607
rect 1654 5405 1657 5431
rect 1683 5426 1686 5431
rect 1683 5409 1728 5426
rect 1683 5405 1686 5409
rect 1165 5384 1202 5388
rect 29 5249 825 5289
rect 933 5375 1202 5384
rect 2031 5376 2034 5381
rect 933 5358 1728 5375
rect 1974 5359 2034 5376
rect 933 5347 1202 5358
rect 2031 5355 2034 5359
rect 2060 5376 2063 5381
rect 2060 5359 2069 5376
rect 2060 5355 2063 5359
rect 3826 5358 3886 5375
rect 3613 5354 3652 5356
rect 933 5336 1048 5347
rect 933 5291 1044 5336
rect 1651 5313 1654 5339
rect 1680 5334 1683 5339
rect 1680 5317 1728 5334
rect 3613 5321 3616 5354
rect 3649 5346 3652 5354
rect 3826 5346 3843 5358
rect 3649 5329 3843 5346
rect 3649 5321 3652 5329
rect 3613 5319 3652 5321
rect 1680 5313 1683 5317
rect 1165 5291 1202 5295
rect 5078 5294 5098 5587
rect 5854 5584 5857 5587
rect 5883 5607 5886 5610
rect 5883 5587 5894 5607
rect 5883 5584 5886 5587
rect 5854 5583 5886 5584
rect 7718 5556 7776 5571
rect 7718 5553 7730 5556
rect 7718 5527 7727 5553
rect 7762 5527 7776 5556
rect 7820 5555 7878 5570
rect 7820 5554 7833 5555
rect 7820 5528 7829 5554
rect 7718 5524 7730 5527
rect 7762 5524 7782 5527
rect 7718 5508 7782 5524
rect 7758 5447 7782 5508
rect 7820 5523 7833 5528
rect 7865 5523 7878 5555
rect 7820 5507 7878 5523
rect 8102 5559 8149 5562
rect 8102 5516 8104 5559
rect 8147 5556 8149 5559
rect 10592 5557 10621 5558
rect 10592 5556 10622 5557
rect 11645 5556 11690 5558
rect 8147 5516 10595 5556
rect 8102 5513 10595 5516
rect 10621 5513 11691 5556
rect 10592 5512 10622 5513
rect 10592 5510 10621 5512
rect 11595 5445 11631 5446
rect 10210 5427 10240 5429
rect 11539 5427 11631 5445
rect 933 5283 1202 5291
rect 2028 5284 2031 5289
rect 933 5266 1728 5283
rect 1974 5267 2031 5284
rect 933 5254 1202 5266
rect 2028 5263 2031 5267
rect 2057 5284 2060 5289
rect 2057 5267 2069 5284
rect 4708 5274 5098 5294
rect 5393 5407 5422 5425
rect 2057 5263 2060 5267
rect 933 5250 1023 5254
rect 29 5188 156 5249
rect 72 4795 199 4883
rect 933 4795 970 5250
rect 1652 5221 1655 5247
rect 1681 5242 1684 5247
rect 1681 5225 1728 5242
rect 1681 5221 1684 5225
rect 3549 5194 3588 5195
rect 1081 5181 1730 5183
rect 72 4758 970 4795
rect 1052 5164 1730 5181
rect 2092 5177 2095 5180
rect 1052 5146 1202 5164
rect 1971 5157 2095 5177
rect 2092 5154 2095 5157
rect 2121 5177 2124 5180
rect 2121 5157 2134 5177
rect 3549 5161 3552 5194
rect 3585 5186 3588 5194
rect 3843 5186 3886 5203
rect 3585 5169 3906 5186
rect 3585 5161 3588 5169
rect 3843 5167 3860 5169
rect 3549 5160 3588 5161
rect 2121 5154 2124 5157
rect 1052 5087 1118 5146
rect 1165 5142 1202 5146
rect 1587 5119 1590 5145
rect 1616 5141 1619 5145
rect 1616 5122 1730 5141
rect 3485 5137 3524 5140
rect 1616 5119 1619 5122
rect 3485 5104 3488 5137
rect 3521 5129 3524 5137
rect 3521 5112 3906 5129
rect 5393 5123 5411 5407
rect 10209 5385 10212 5427
rect 10238 5417 11631 5427
rect 10238 5385 11635 5417
rect 10210 5383 10240 5385
rect 11539 5351 11635 5385
rect 7828 5209 7888 5220
rect 7828 5175 7841 5209
rect 7875 5175 7888 5209
rect 8188 5203 8711 5226
rect 8748 5203 9663 5226
rect 11545 5208 11635 5351
rect 7828 5164 7888 5175
rect 9634 5193 9663 5203
rect 10432 5193 10546 5201
rect 9634 5181 10546 5193
rect 9634 5173 10467 5181
rect 9634 5172 9663 5173
rect 3521 5104 3524 5112
rect 5316 5106 5411 5123
rect 8189 5121 8711 5143
rect 8748 5121 9569 5143
rect 3485 5102 3524 5104
rect 1052 5068 1730 5087
rect 2093 5081 2096 5084
rect 1052 5050 1202 5068
rect 1971 5061 2096 5081
rect 2093 5058 2096 5061
rect 2122 5081 2125 5084
rect 2122 5061 2134 5081
rect 4750 5063 4770 5075
rect 2122 5058 2125 5061
rect 1052 5049 1119 5050
rect 1052 5045 1118 5049
rect 1165 5046 1202 5050
rect 72 4695 199 4758
rect 66 4319 193 4408
rect 1052 4319 1089 5045
rect 1583 5023 1586 5049
rect 1612 5045 1615 5049
rect 1612 5026 1730 5045
rect 4750 5043 4785 5063
rect 4750 5041 4770 5043
rect 1612 5023 1615 5026
rect 4712 5021 4770 5041
rect 66 4282 1089 4319
rect 1165 4972 1730 4991
rect 2092 4985 2095 4988
rect 66 4220 193 4282
rect 72 3835 199 3926
rect 1165 3835 1202 4972
rect 1971 4965 2095 4985
rect 2092 4962 2095 4965
rect 2121 4985 2124 4988
rect 2121 4965 2134 4985
rect 3424 4980 3463 4982
rect 2121 4962 2124 4965
rect 1587 4927 1590 4953
rect 1616 4949 1619 4953
rect 1616 4930 1730 4949
rect 3424 4947 3427 4980
rect 3460 4972 3463 4980
rect 3460 4955 3906 4972
rect 3460 4947 3463 4955
rect 3424 4945 3463 4947
rect 3851 4939 3886 4955
rect 1616 4927 1619 4930
rect 4745 4921 4782 4941
rect 4745 4866 4765 4921
rect 5349 4918 5422 4936
rect 9547 4933 9569 5121
rect 9809 5105 9855 5108
rect 9809 5065 9812 5105
rect 9852 5095 9855 5105
rect 10440 5095 10546 5103
rect 9852 5083 10546 5095
rect 10982 5083 11154 5103
rect 9852 5075 10467 5083
rect 10982 5075 11153 5083
rect 9852 5065 9855 5075
rect 9809 5063 9855 5065
rect 9910 5037 9946 5040
rect 11133 5030 11153 5075
rect 9946 5010 10546 5030
rect 10982 5010 11153 5030
rect 9910 4998 9946 5001
rect 9547 4932 9707 4933
rect 5349 4897 5367 4918
rect 9547 4912 10546 4932
rect 9547 4911 9707 4912
rect 11133 4905 11153 5010
rect 11542 4905 11632 4972
rect 6019 4902 6050 4903
rect 5310 4879 5367 4897
rect 6018 4901 6051 4902
rect 6018 4896 6021 4901
rect 5983 4891 6021 4896
rect 5660 4874 6021 4891
rect 6048 4874 6051 4901
rect 8266 4875 8711 4891
rect 5660 4869 6050 4874
rect 8263 4871 8711 4875
rect 8748 4881 10467 4891
rect 8748 4871 10546 4881
rect 4712 4846 4765 4866
rect 7722 4862 7778 4871
rect 3361 4827 3403 4828
rect 3361 4794 3364 4827
rect 3397 4819 3403 4827
rect 7722 4827 7734 4862
rect 7767 4827 7778 4862
rect 3397 4802 3851 4819
rect 3397 4794 3403 4802
rect 3361 4793 3403 4794
rect 3834 4784 3851 4802
rect 5359 4803 5414 4821
rect 7722 4817 7778 4827
rect 5359 4801 5377 4803
rect 5317 4785 5377 4801
rect 3834 4767 3886 4784
rect 4748 4710 4780 4754
rect 4748 4691 4768 4710
rect 4712 4671 4768 4691
rect 3305 4670 3344 4671
rect 3305 4637 3308 4670
rect 3341 4662 3344 4670
rect 3341 4645 3842 4662
rect 3341 4637 3344 4645
rect 3305 4636 3344 4637
rect 3826 4634 3842 4645
rect 3826 4604 3843 4634
rect 8263 4623 8286 4871
rect 10437 4861 10546 4871
rect 11133 4862 11632 4905
rect 10002 4804 10041 4806
rect 10001 4803 10042 4804
rect 10001 4764 10002 4803
rect 10041 4793 10042 4803
rect 11133 4793 11153 4862
rect 10041 4783 10467 4793
rect 10041 4773 10546 4783
rect 10041 4764 10042 4773
rect 10001 4763 10042 4764
rect 10444 4763 10546 4773
rect 10982 4763 11153 4793
rect 11542 4763 11632 4862
rect 10002 4761 10041 4763
rect 10084 4734 10124 4735
rect 10082 4708 10085 4734
rect 10123 4728 10126 4734
rect 11133 4728 11153 4763
rect 10123 4710 10467 4728
rect 10982 4710 11153 4728
rect 10123 4708 10546 4710
rect 10084 4707 10124 4708
rect 10432 4690 10546 4708
rect 10976 4696 11153 4710
rect 10976 4690 11152 4696
rect 3826 4587 3886 4604
rect 4741 4598 4779 4616
rect 7826 4606 7888 4615
rect 4741 4516 4759 4598
rect 5315 4553 5387 4571
rect 7826 4570 7843 4606
rect 7877 4570 7888 4606
rect 8188 4600 8286 4623
rect 8347 4610 8711 4630
rect 8748 4612 10467 4630
rect 8748 4610 10546 4612
rect 7826 4562 7888 4570
rect 4712 4496 4760 4516
rect 5369 4334 5387 4553
rect 8347 4540 8367 4610
rect 10441 4592 10546 4610
rect 8189 4525 8367 4540
rect 8189 4518 8364 4525
rect 11268 4354 11346 4357
rect 5369 4316 5423 4334
rect 11268 4283 11271 4354
rect 11342 4342 11346 4354
rect 11542 4342 11632 4434
rect 11342 4295 11632 4342
rect 11342 4283 11346 4295
rect 11268 4280 11346 4283
rect 8464 4245 8510 4247
rect 5683 4240 5715 4241
rect 8464 4240 8469 4245
rect 5683 4238 8469 4240
rect 5683 4210 5685 4238
rect 5713 4212 8469 4238
rect 5713 4210 5715 4212
rect 5683 4207 5715 4210
rect 8464 4208 8469 4212
rect 8506 4208 8510 4245
rect 11542 4225 11632 4295
rect 8464 4206 8510 4208
rect 8543 4186 8586 4188
rect 8543 4180 8546 4186
rect 7417 4179 8546 4180
rect 7417 4153 7420 4179
rect 7446 4154 8546 4179
rect 7446 4153 7449 4154
rect 8543 4149 8546 4154
rect 8583 4149 8586 4186
rect 8543 4147 8586 4149
rect 3244 4123 3281 4127
rect 3244 4090 3246 4123
rect 3279 4115 3281 4123
rect 3279 4098 3876 4115
rect 3279 4090 3281 4098
rect 3244 4087 3281 4090
rect 5361 4074 5379 4075
rect 5327 4063 5379 4074
rect 5327 4056 5562 4063
rect 5361 4045 5562 4056
rect 4719 4008 4779 4028
rect 3180 3964 3219 3965
rect 3180 3931 3183 3964
rect 3216 3956 3219 3964
rect 3216 3944 3876 3956
rect 8617 3953 8661 3955
rect 3216 3939 3886 3944
rect 8617 3943 8620 3953
rect 3216 3931 3219 3939
rect 3180 3930 3219 3931
rect 3847 3927 3886 3939
rect 8604 3925 8620 3943
rect 8616 3916 8620 3925
rect 8657 3916 8661 3953
rect 8616 3915 8661 3916
rect 8616 3909 8656 3915
rect 7533 3891 8656 3909
rect 4739 3888 4777 3889
rect 4737 3871 4777 3888
rect 4737 3853 4757 3871
rect 72 3798 1202 3835
rect 4712 3833 4757 3853
rect 5335 3850 5568 3866
rect 5313 3848 5568 3850
rect 5313 3832 5353 3848
rect 9270 3845 9330 3849
rect 72 3738 199 3798
rect 3118 3776 3121 3809
rect 3154 3801 3157 3809
rect 3154 3784 3836 3801
rect 9270 3795 9273 3845
rect 9323 3843 9330 3845
rect 11542 3843 11632 3946
rect 9323 3796 11632 3843
rect 9323 3795 9330 3796
rect 9270 3791 9330 3795
rect 3154 3776 3157 3784
rect 3821 3777 3836 3784
rect 3821 3766 3838 3777
rect 3821 3749 3886 3766
rect 5315 3753 5355 3754
rect 5315 3739 5356 3753
rect 5315 3738 5566 3739
rect 5338 3721 5566 3738
rect 11542 3737 11632 3796
rect 4732 3693 4777 3706
rect 4732 3678 4781 3693
rect 4712 3673 4781 3678
rect 3057 3661 3099 3662
rect 3057 3628 3061 3661
rect 3094 3653 3099 3661
rect 4712 3658 4767 3673
rect 3094 3636 3838 3653
rect 3094 3628 3099 3636
rect 3057 3626 3099 3628
rect 3821 3587 3838 3636
rect 3821 3570 3886 3587
rect 4736 3551 4779 3574
rect 66 3420 193 3504
rect 4736 3503 4756 3551
rect 5334 3525 5564 3543
rect 5334 3524 5354 3525
rect 5313 3506 5354 3524
rect 4712 3483 4756 3503
rect 1583 3446 1614 3448
rect 1649 3446 1680 3448
rect 66 3383 1036 3420
rect 1583 3399 1586 3446
rect 1612 3399 1650 3446
rect 1676 3399 2315 3446
rect 1583 3397 1614 3399
rect 1649 3397 1680 3399
rect 66 3316 193 3383
rect 999 3248 1036 3383
rect 2268 3331 2315 3399
rect 4945 3432 4976 3434
rect 8709 3432 8754 3435
rect 4945 3391 4948 3432
rect 4974 3391 8713 3432
rect 8750 3391 8754 3432
rect 4945 3389 4976 3391
rect 8709 3389 8754 3391
rect 11545 3331 11635 3428
rect 1450 3322 1476 3325
rect 2268 3323 11635 3331
rect 1655 3318 1658 3320
rect 1476 3299 1658 3318
rect 1450 3293 1476 3296
rect 1655 3294 1658 3299
rect 1684 3318 1687 3320
rect 1831 3318 1834 3322
rect 1684 3299 1834 3318
rect 1684 3294 1687 3299
rect 1831 3295 1834 3299
rect 1861 3295 1864 3322
rect 2268 3284 9165 3323
rect 1395 3256 1398 3282
rect 1424 3278 1427 3282
rect 1589 3278 1592 3284
rect 1424 3259 1592 3278
rect 1424 3256 1427 3259
rect 1589 3258 1592 3259
rect 1618 3278 1621 3284
rect 1881 3278 1884 3282
rect 1618 3259 1884 3278
rect 1618 3258 1621 3259
rect 1881 3256 1884 3259
rect 1910 3256 1913 3282
rect 9161 3276 9165 3284
rect 9215 3284 11635 3323
rect 9215 3276 9218 3284
rect 9161 3272 9218 3276
rect 999 3247 1202 3248
rect 999 3229 1224 3247
rect 999 3223 1364 3229
rect 999 3211 1497 3223
rect 2029 3222 2059 3224
rect 2028 3220 2031 3222
rect 1165 3207 1497 3211
rect 1202 3201 1497 3207
rect 465 3197 542 3201
rect 465 3131 470 3197
rect 536 3182 542 3197
rect 1806 3198 2031 3220
rect 1165 3182 1204 3184
rect 536 3178 1204 3182
rect 536 3157 1496 3178
rect 536 3145 1203 3157
rect 1806 3154 1828 3198
rect 2028 3196 2031 3198
rect 2057 3196 2060 3222
rect 11545 3219 11635 3284
rect 2029 3194 2059 3196
rect 3840 3190 3882 3207
rect 3840 3180 3878 3190
rect 3840 3158 3868 3180
rect 536 3131 542 3145
rect 1165 3143 1202 3145
rect 2993 3144 3034 3146
rect 465 3127 542 3131
rect 2993 3111 2997 3144
rect 3030 3136 3034 3144
rect 3840 3136 3867 3158
rect 3030 3119 3867 3136
rect 5316 3130 5347 3148
rect 3030 3111 3034 3119
rect 3840 3118 3857 3119
rect 2993 3110 3034 3111
rect 1967 3107 1996 3109
rect 1966 3103 1969 3107
rect 72 3017 199 3094
rect 1809 3084 1969 3103
rect 1966 3081 1969 3084
rect 1995 3081 1998 3107
rect 4708 3102 4769 3122
rect 5329 3112 5564 3130
rect 4749 3098 4769 3102
rect 1967 3079 1996 3081
rect 4749 3078 4791 3098
rect 5393 3049 5510 3064
rect 5387 3045 5415 3049
rect 72 2980 671 3017
rect 3834 3014 3882 3031
rect 5387 3019 5388 3045
rect 5414 3019 5415 3045
rect 7373 3038 7376 3043
rect 6895 3022 7376 3038
rect 5387 3016 5415 3019
rect 7373 3017 7376 3022
rect 7402 3017 7405 3043
rect 72 2906 199 2980
rect 634 2814 671 2980
rect 2927 2987 2966 2990
rect 2927 2954 2930 2987
rect 2963 2979 2966 2987
rect 3834 2985 3851 3014
rect 3834 2979 3850 2985
rect 2963 2963 3850 2979
rect 2963 2962 3815 2963
rect 2963 2954 2966 2962
rect 2927 2952 2966 2954
rect 4748 2947 4780 2963
rect 4708 2927 4780 2947
rect 7321 2945 7324 2950
rect 5327 2922 5506 2935
rect 6895 2929 7324 2945
rect 7321 2924 7324 2929
rect 7350 2924 7353 2950
rect 5313 2917 5506 2922
rect 5313 2902 5345 2917
rect 5313 2894 5331 2902
rect 1398 2891 1427 2892
rect 1397 2865 1400 2891
rect 1426 2889 1429 2891
rect 1426 2867 1497 2889
rect 1426 2865 1429 2867
rect 1398 2863 1427 2865
rect 1924 2846 1956 2848
rect 1924 2843 1927 2846
rect 1807 2822 1927 2843
rect 1924 2820 1927 2822
rect 1953 2820 1956 2846
rect 3826 2833 3882 2850
rect 3826 2829 3843 2833
rect 1924 2818 1956 2820
rect 2866 2825 2903 2826
rect 3826 2825 3842 2829
rect 2866 2823 3842 2825
rect 634 2796 1229 2814
rect 634 2789 1236 2796
rect 1375 2789 1497 2790
rect 2093 2789 2122 2791
rect 2866 2790 2868 2823
rect 2901 2808 3842 2823
rect 5318 2811 5338 2827
rect 2901 2790 2903 2808
rect 634 2777 1497 2789
rect 2092 2786 2095 2789
rect 1165 2773 1497 2777
rect 1201 2768 1497 2773
rect 1807 2765 2095 2786
rect 988 2716 1029 2718
rect 1165 2716 1364 2718
rect 72 2603 199 2685
rect 988 2679 991 2716
rect 1028 2712 1364 2716
rect 1028 2690 1497 2712
rect 1028 2679 1203 2690
rect 1807 2683 1828 2765
rect 2092 2763 2095 2765
rect 2121 2763 2124 2789
rect 2866 2787 2903 2790
rect 5320 2806 5338 2811
rect 9049 2807 9104 2808
rect 5320 2788 5509 2806
rect 4708 2770 4777 2772
rect 2093 2761 2122 2763
rect 4708 2752 4785 2770
rect 4756 2743 4785 2752
rect 5448 2767 5480 2769
rect 5448 2741 5451 2767
rect 5477 2765 5480 2767
rect 5477 2744 5509 2765
rect 7274 2761 7277 2766
rect 6895 2745 7277 2761
rect 5477 2741 5494 2744
rect 5448 2737 5494 2741
rect 7274 2740 7277 2745
rect 7303 2740 7306 2766
rect 9049 2757 9052 2807
rect 9102 2805 9105 2807
rect 11542 2805 11632 2920
rect 9102 2758 11632 2805
rect 9102 2757 9105 2758
rect 9049 2755 9104 2757
rect 11542 2711 11632 2758
rect 2797 2679 2836 2681
rect 988 2677 1029 2679
rect 1165 2677 1202 2679
rect 2797 2646 2800 2679
rect 2833 2671 2836 2679
rect 3817 2671 3882 2678
rect 2833 2661 3882 2671
rect 7224 2668 7227 2673
rect 2833 2654 3846 2661
rect 4754 2655 4784 2659
rect 2833 2646 2836 2654
rect 3829 2652 3846 2654
rect 2797 2644 2836 2646
rect 4753 2631 4784 2655
rect 6895 2652 7227 2668
rect 7224 2647 7227 2652
rect 7253 2647 7256 2673
rect 465 2611 545 2617
rect 465 2603 474 2611
rect 72 2553 474 2603
rect 72 2497 199 2553
rect 465 2545 474 2553
rect 540 2545 545 2611
rect 4753 2597 4773 2631
rect 5344 2597 5507 2610
rect 4708 2577 4773 2597
rect 5313 2592 5507 2597
rect 5313 2579 5362 2592
rect 465 2540 545 2545
rect 5388 2536 5420 2537
rect 4727 2506 4730 2532
rect 4756 2527 4759 2532
rect 5388 2527 5391 2536
rect 4756 2511 5391 2527
rect 4756 2506 4759 2511
rect 5388 2510 5391 2511
rect 5417 2510 5420 2536
rect 5388 2509 5420 2510
rect 5491 2535 5523 2556
rect 5491 2509 5494 2535
rect 5520 2525 5523 2535
rect 6553 2537 6594 2538
rect 6553 2527 6556 2537
rect 5856 2525 6556 2527
rect 5520 2511 6556 2525
rect 5520 2509 5523 2511
rect 5491 2508 5523 2509
rect 5848 2504 6556 2511
rect 5447 2503 5475 2504
rect 4674 2498 4707 2500
rect 4673 2469 4676 2498
rect 4705 2490 4708 2498
rect 5248 2495 5280 2496
rect 5248 2490 5251 2495
rect 4705 2474 5251 2490
rect 4705 2469 4708 2474
rect 5248 2469 5251 2474
rect 5277 2469 5280 2495
rect 5445 2494 5448 2503
rect 5442 2478 5448 2494
rect 5445 2477 5448 2478
rect 5474 2494 5477 2503
rect 6553 2502 6556 2504
rect 6591 2502 6594 2537
rect 6553 2501 6594 2502
rect 9568 2529 9624 2531
rect 5669 2494 5672 2497
rect 5474 2478 5672 2494
rect 5474 2477 5477 2478
rect 5447 2476 5475 2477
rect 5669 2471 5672 2478
rect 5698 2471 5701 2497
rect 9568 2479 9571 2529
rect 9621 2524 9624 2529
rect 10840 2529 10908 2530
rect 10840 2524 10851 2529
rect 9621 2483 10851 2524
rect 9621 2479 9624 2483
rect 9568 2478 9624 2479
rect 10840 2478 10851 2483
rect 10902 2524 10908 2529
rect 11593 2524 11659 2588
rect 10902 2483 11659 2524
rect 10902 2478 10908 2483
rect 10840 2477 10908 2478
rect 11593 2473 11659 2483
rect 5671 2470 5699 2471
rect 4673 2467 4708 2469
rect 5870 2455 5898 2458
rect 4231 2449 4264 2452
rect 4231 2418 4232 2449
rect 4263 2428 4264 2449
rect 4817 2441 4847 2442
rect 4816 2428 4819 2441
rect 4263 2418 4819 2428
rect 4231 2415 4819 2418
rect 4845 2428 4848 2441
rect 5870 2429 5871 2455
rect 5897 2429 5898 2455
rect 5870 2428 5898 2429
rect 6273 2453 6303 2456
rect 6273 2428 6275 2453
rect 4845 2426 6275 2428
rect 6302 2426 6303 2453
rect 4845 2423 6302 2426
rect 4845 2415 6296 2423
rect 4231 2412 6296 2415
rect 4612 2390 4656 2391
rect 80 2389 4656 2390
rect 80 2348 4613 2389
rect 3927 2347 3975 2348
rect 4610 2347 4613 2348
rect 4655 2347 4658 2389
rect 5549 2379 5587 2382
rect 7157 2381 7187 2383
rect 4612 2346 4656 2347
rect 5549 2346 5552 2379
rect 5585 2346 5587 2379
rect 5549 2343 5587 2346
rect 5664 2339 5667 2373
rect 5701 2339 5704 2373
rect 6523 2357 6589 2359
rect 6523 2325 6560 2357
rect 6586 2325 6589 2357
rect 7086 2347 7159 2381
rect 7185 2347 7188 2381
rect 7157 2345 7188 2347
rect 6523 2323 6589 2325
rect 78 2251 1971 2293
rect 1997 2281 4228 2293
rect 1997 2251 2396 2281
rect 2383 2210 2396 2251
rect 2454 2251 4228 2281
rect 4270 2251 4276 2293
rect 6698 2292 6743 2294
rect 4679 2274 4717 2277
rect 2454 2210 2466 2251
rect 4679 2242 4681 2274
rect 4713 2242 4717 2274
rect 6698 2254 6702 2292
rect 6740 2254 6743 2292
rect 6698 2251 6743 2254
rect 8944 2277 9004 2280
rect 4679 2239 4717 2242
rect 8944 2227 8947 2277
rect 8997 2275 9004 2277
rect 11585 2275 11795 2369
rect 8997 2228 11795 2275
rect 8997 2227 9004 2228
rect 8944 2224 9004 2227
rect 2383 2201 2466 2210
rect 66 2092 193 2170
rect 11585 2161 11795 2228
rect 11587 2160 11664 2161
rect 989 2092 1030 2094
rect 66 2055 990 2092
rect 1027 2055 1030 2092
rect 7371 2076 7374 2126
rect 7400 2076 13025 2126
rect 66 1982 193 2055
rect 989 2053 1030 2055
rect 1742 2049 1771 2051
rect 1965 2049 1996 2051
rect 1741 2013 1744 2049
rect 1770 2013 1967 2049
rect 1993 2013 1996 2049
rect 12415 2036 12616 2038
rect 1742 2011 1771 2013
rect 1965 2011 1996 2013
rect 7317 1986 7320 2036
rect 7346 1986 12616 2036
rect 7270 1896 7273 1946
rect 7299 1944 12197 1946
rect 7299 1896 12208 1944
rect 7222 1806 7225 1856
rect 7251 1855 11801 1856
rect 7251 1806 11822 1855
rect 5081 1797 6171 1798
rect 5081 1795 5157 1797
rect 5080 1767 5083 1795
rect 5111 1770 5157 1795
rect 5111 1767 5114 1770
rect 5154 1769 5157 1770
rect 5185 1795 6171 1797
rect 5185 1770 6064 1795
rect 5185 1769 5188 1770
rect 6061 1767 6064 1770
rect 6092 1770 6171 1795
rect 6092 1767 6095 1770
rect 1161 1753 1198 1754
rect 72 1671 199 1741
rect 1029 1715 1290 1753
rect 4688 1716 4738 1717
rect 9281 1716 9284 1718
rect 1029 1671 1067 1715
rect 1161 1713 1198 1715
rect 4688 1710 9284 1716
rect 2028 1683 2056 1684
rect 72 1633 1067 1671
rect 1669 1650 2029 1683
rect 2055 1650 2058 1683
rect 4688 1664 4691 1710
rect 4737 1670 9284 1710
rect 4737 1664 4740 1670
rect 9281 1668 9284 1670
rect 9334 1668 9337 1718
rect 4688 1662 4738 1664
rect 2028 1648 2056 1650
rect 72 1553 199 1633
rect 5519 1619 9227 1625
rect 5519 1615 9165 1619
rect 5519 1579 5529 1615
rect 5526 1569 5529 1579
rect 5575 1579 9165 1615
rect 5575 1569 5578 1579
rect 9162 1573 9165 1579
rect 9215 1579 9227 1619
rect 9215 1573 9218 1579
rect 5663 1532 9118 1534
rect 5663 1527 9052 1532
rect 5662 1526 9052 1527
rect 1286 1489 1289 1518
rect 1318 1515 1321 1518
rect 1924 1517 1957 1521
rect 1923 1515 1926 1517
rect 1318 1489 1926 1515
rect 1290 1488 1926 1489
rect 1955 1515 1958 1517
rect 1955 1488 2289 1515
rect 1290 1486 2289 1488
rect 1924 1484 1957 1486
rect 1670 1447 1904 1452
rect 1670 1392 1810 1447
rect 1807 1387 1810 1392
rect 1870 1418 1904 1447
rect 1870 1394 1908 1418
rect 1870 1392 1904 1394
rect 1870 1387 1873 1392
rect 1807 1385 1873 1387
rect 1810 1384 1870 1385
rect 2259 1278 2288 1486
rect 5662 1480 5672 1526
rect 5718 1488 9052 1526
rect 5718 1480 5727 1488
rect 9049 1486 9052 1488
rect 9102 1488 9118 1532
rect 9102 1486 9105 1488
rect 5662 1475 5727 1480
rect 6507 1440 6559 1442
rect 8956 1440 8959 1441
rect 6507 1435 8959 1440
rect 6507 1389 6511 1435
rect 6557 1395 8959 1435
rect 9009 1440 9012 1441
rect 9009 1395 9021 1440
rect 6557 1394 9021 1395
rect 6557 1389 6560 1394
rect 6507 1384 6559 1389
rect 3901 1278 3933 1280
rect 9501 1278 9617 1281
rect 72 1148 199 1239
rect 2240 1166 3904 1278
rect 3930 1276 9513 1278
rect 3930 1274 6022 1276
rect 3930 1272 5115 1274
rect 3930 1166 5041 1272
rect 3901 1164 3933 1166
rect 5038 1160 5041 1166
rect 5227 1166 6022 1274
rect 5227 1162 5230 1166
rect 5153 1160 5230 1162
rect 5038 1158 5230 1160
rect 6019 1157 6022 1166
rect 6208 1166 9513 1276
rect 9607 1166 9617 1278
rect 6208 1157 6212 1166
rect 9501 1163 9617 1166
rect 6019 1155 6212 1157
rect 72 1110 1069 1148
rect 72 1051 199 1110
rect 1031 1025 1069 1110
rect 1161 1025 1198 1026
rect 1031 987 1303 1025
rect 1161 985 1198 987
rect 2086 928 2117 930
rect 1663 894 2088 928
rect 2114 894 2117 928
rect 2086 892 2117 894
rect 193 839 243 844
rect 193 800 197 839
rect 236 833 243 839
rect 7090 836 7129 837
rect 7089 833 7092 836
rect 236 805 7092 833
rect 236 800 243 805
rect 7089 803 7092 805
rect 7125 803 7129 836
rect 7090 802 7129 803
rect 193 797 243 800
rect 3731 770 3773 771
rect 3731 737 3736 770
rect 3769 745 7758 770
rect 3769 737 7759 745
rect 3731 736 3773 737
rect 7155 735 7759 737
rect 3671 708 3709 709
rect 59 497 186 685
rect 3671 675 3674 708
rect 3707 675 7351 708
rect 3671 674 3709 675
rect 6744 674 7351 675
rect 3607 645 3649 646
rect 3607 612 3611 645
rect 3644 612 6943 645
rect 3607 611 3649 612
rect 3548 582 3588 583
rect 3548 549 3551 582
rect 3584 581 3588 582
rect 3584 549 6542 581
rect 3548 548 6542 549
rect 3548 547 3588 548
rect 3482 514 3523 515
rect 3481 481 3487 514
rect 3520 481 6133 514
rect 3482 479 3523 481
rect 3424 452 3465 453
rect 3424 419 3427 452
rect 3460 450 5731 452
rect 3460 419 5732 450
rect 3424 418 3465 419
rect 3364 355 3367 388
rect 3400 387 3403 388
rect 3400 355 5333 387
rect 3374 354 5333 355
rect 2792 306 2846 309
rect 2792 305 2797 306
rect 1509 301 2797 305
rect 1504 263 2797 301
rect 2840 263 2846 306
rect 3306 298 3309 331
rect 3342 326 3345 331
rect 3342 298 4942 326
rect 3332 293 4942 298
rect 1504 262 2846 263
rect 66 22 193 210
rect 1504 74 1705 262
rect 2792 259 2846 262
rect 3248 229 3251 262
rect 3284 229 4522 262
rect 2857 227 2911 228
rect 2857 221 2862 227
rect 1914 184 2862 221
rect 2905 184 2911 227
rect 3909 199 4111 201
rect 3193 198 4114 199
rect 1914 178 2911 184
rect 1914 77 2112 178
rect 3183 165 3186 198
rect 3219 166 4114 198
rect 3219 165 3222 166
rect 2925 156 2974 160
rect 2925 140 2929 156
rect 2364 138 2929 140
rect 2307 116 2929 138
rect 2969 116 2974 156
rect 2307 110 2974 116
rect 2307 100 2965 110
rect 3119 100 3122 134
rect 3155 100 3717 134
rect 2307 77 2505 100
rect 2908 77 2973 78
rect 1502 8 1705 74
rect 1909 11 2112 77
rect 2305 11 2508 77
rect 2705 73 2973 77
rect 2705 22 2912 73
rect 2963 22 2973 73
rect 3058 75 3113 77
rect 3058 73 3313 75
rect 3514 74 3718 100
rect 3058 36 3064 73
rect 3101 36 3313 73
rect 3058 32 3313 36
rect 2705 14 2973 22
rect 2705 11 2908 14
rect 3110 9 3313 32
rect 3513 8 3718 74
rect 3906 11 4114 166
rect 4317 99 4520 229
rect 4317 70 4521 99
rect 4318 9 4521 70
rect 4735 11 4938 293
rect 5134 83 5333 354
rect 5133 8 5336 83
rect 5532 81 5732 419
rect 5529 11 5732 81
rect 5942 74 6133 481
rect 6346 76 6541 548
rect 6744 76 6943 612
rect 7155 642 7351 674
rect 7565 685 7759 735
rect 9817 724 9860 726
rect 7967 721 8163 724
rect 9815 721 9818 724
rect 7967 686 9818 721
rect 7155 76 7350 642
rect 7565 78 7758 685
rect 5934 9 6137 74
rect 6341 11 6544 76
rect 6744 11 6947 76
rect 7149 11 7352 76
rect 7556 0 7759 78
rect 7967 76 8163 686
rect 9815 684 9818 686
rect 9858 684 9861 724
rect 9817 683 9860 684
rect 9907 643 9950 645
rect 9906 642 9909 643
rect 8360 604 9909 642
rect 9948 604 9951 643
rect 7964 11 8167 76
rect 8360 74 8556 604
rect 9907 602 9950 604
rect 9999 560 10002 561
rect 8775 522 10002 560
rect 10041 522 10044 561
rect 8775 76 8973 522
rect 10083 481 10125 484
rect 9186 443 10084 481
rect 10122 443 10125 481
rect 8359 9 8562 74
rect 8771 11 8974 76
rect 9186 73 9384 443
rect 10083 440 10125 443
rect 9693 144 10317 164
rect 9693 76 9713 144
rect 10409 123 10429 164
rect 10186 103 10429 123
rect 10186 76 10206 103
rect 10506 76 10527 165
rect 9185 8 9388 73
rect 9584 11 9787 76
rect 9986 46 10206 76
rect 9986 11 10189 46
rect 10394 11 10597 76
rect 10699 67 10720 165
rect 10796 146 10815 163
rect 10796 127 11296 146
rect 11277 81 11296 127
rect 10812 67 11015 76
rect 11277 74 11380 81
rect 11621 76 11822 1806
rect 10699 46 11015 67
rect 10812 11 11015 46
rect 11210 9 11413 74
rect 11615 24 11822 76
rect 12007 76 12208 1896
rect 11615 11 11818 24
rect 12007 11 12214 76
rect 12415 74 12616 1986
rect 12824 76 13025 2076
rect 12007 7 12208 11
rect 12415 9 12619 74
rect 12821 18 13025 76
rect 12821 11 13024 18
rect 12415 1 12616 9
<< via2 >>
rect 7730 5553 7762 5556
rect 7730 5527 7753 5553
rect 7753 5527 7762 5553
rect 7833 5554 7865 5555
rect 7833 5528 7855 5554
rect 7855 5528 7865 5554
rect 7730 5524 7762 5527
rect 7833 5523 7865 5528
rect 7841 5175 7875 5209
rect 7734 4827 7767 4862
rect 7843 4570 7877 4606
<< metal3 >>
rect 7723 5556 7768 5562
rect 7723 5524 7730 5556
rect 7762 5524 7768 5556
rect 7723 5487 7768 5524
rect 7827 5555 7872 5561
rect 7827 5523 7833 5555
rect 7865 5523 7872 5555
rect 7723 4871 7760 5487
rect 7827 5486 7872 5523
rect 7835 5222 7872 5486
rect 7835 5209 7879 5222
rect 7835 5175 7841 5209
rect 7875 5175 7879 5209
rect 7835 5162 7879 5175
rect 7723 4862 7772 4871
rect 7723 4838 7734 4862
rect 7728 4827 7734 4838
rect 7767 4827 7772 4862
rect 7728 4822 7772 4827
rect 7835 4651 7872 5162
rect 7834 4606 7881 4651
rect 7834 4570 7843 4606
rect 7877 4570 7881 4606
rect 7834 4564 7881 4570
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_0
timestamp 1629137236
transform -1 0 1794 0 -1 1874
box 0 0 464 599
use sky130_hilas_nFETLarge  sky130_hilas_nFETLarge_0
timestamp 1629137224
transform -1 0 1790 0 -1 2629
box 0 0 557 603
use sky130_hilas_Trans2med  sky130_hilas_Trans2med_0
timestamp 1629137246
transform 1 0 1855 0 -1 3104
box 0 0 440 593
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_2
timestamp 1629137211
transform -1 0 4709 0 -1 4033
box 0 0 889 787
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_3
timestamp 1629137211
transform -1 0 4705 0 -1 3127
box 0 0 889 787
use sky130_hilas_WTA4Stage01  sky130_hilas_WTA4Stage01_0
timestamp 1629137241
transform 1 0 6607 0 1 2597
box -2078 -102 350 989
use sky130_hilas_swc4x2cell  sky130_hilas_swc4x2cell_0
timestamp 1629137207
transform 1 0 6547 0 1 3495
box -1017 -41 3029 1049
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_1
timestamp 1629137236
transform 1 0 4606 0 1 1399
box 0 0 464 599
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_2
timestamp 1629137236
transform -1 0 5662 0 1 1399
box 0 0 464 599
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_3
timestamp 1629137236
transform 1 0 5587 0 1 1402
box 0 0 464 599
use sky130_hilas_pFETLarge  sky130_hilas_pFETLarge_4
timestamp 1629137236
transform -1 0 6643 0 1 1402
box 0 0 464 599
use sky130_hilas_nFETLarge  sky130_hilas_nFETLarge_1
timestamp 1629137224
transform -1 0 7217 0 1 1401
box 0 0 557 603
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_2
timestamp 1629137216
transform -1 0 6381 0 -1 4091
box 0 0 572 659
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_3
timestamp 1629137216
transform -1 0 6384 0 -1 3164
box 0 0 572 659
use sky130_hilas_Trans4small  sky130_hilas_Trans4small_0
timestamp 1628285143
transform 1 0 1520 0 1 5052
box 191 -150 531 496
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_1
timestamp 1629137211
transform -1 0 4709 0 -1 5046
box 0 0 889 787
use sky130_hilas_TA2Cell_1FG  sky130_hilas_TA2Cell_1FG_0
timestamp 1629137248
transform 1 0 8018 0 1 4126
box -3117 -304 259 1145
use sky130_hilas_TA2Cell_1FG_Strong  sky130_hilas_TA2Cell_1FG_Strong_0
timestamp 1629137252
transform 1 0 8018 0 1 4729
box 0 0 3352 1449
use sky130_hilas_drainSelect01  sky130_hilas_drainSelect01_1
timestamp 1629137216
transform -1 0 6383 0 -1 5138
box 0 0 572 659
use sky130_hilas_Tgate4Single01  sky130_hilas_Tgate4Single01_0
timestamp 1629137243
transform 1 0 10562 0 1 4740
box 0 0 476 641
use sky130_hilas_FGcharacterization01  sky130_hilas_FGcharacterization01_0
timestamp 1629137247
transform -1 0 2464 0 1 6101
box 0 0 3012 1417
use sky130_hilas_LevelShift4InputUp  sky130_hilas_LevelShift4InputUp_0
timestamp 1629137211
transform -1 0 4709 0 1 5269
box 0 0 889 787
use sky130_hilas_DAC5bit01  sky130_hilas_DAC5bit01_0
timestamp 1629137237
transform 0 1 9694 1 0 -238
box 382 525 2120 1170
<< labels >>
rlabel metal2 12821 11 13024 76 1 DIG24 
port 1 n
rlabel metal2 12416 9 12619 74 0 DIG23
port 2 nsew
rlabel metal2 12011 11 12214 76 0 DIG22
port 3 nsew
rlabel metal2 11615 11 11818 76 0 DIG21
port 4 nsew
rlabel metal2 11210 9 11413 74 0 DIG29
port 5 nsew
rlabel metal2 10812 11 11015 76 0 DIG28
port 6 nsew
rlabel metal2 10394 11 10597 76 0 DIG27
port 7 nsew
rlabel metal2 9986 11 10189 76 0 DIG26
port 8 nsew
rlabel metal2 9584 11 9787 76 0 DIG25
port 9 nsew
rlabel metal2 9185 8 9388 73 0 DIG20
port 10 nsew
rlabel metal2 8771 11 8974 76 0 DIG19
port 11 nsew
rlabel metal2 8359 9 8562 74 0 DIG18
port 12 nsew
rlabel metal2 7964 11 8167 76 0 DIG17
port 13 nsew
rlabel metal2 7556 13 7759 78 0 DIG16
port 14 nsew
rlabel metal2 7149 11 7352 76 0 DIG15
port 15 nsew
rlabel metal2 6744 11 6947 76 0 DIG14
port 16 nsew
rlabel metal2 6341 11 6544 76 0 DIG13
port 17 nsew
rlabel metal2 5934 9 6137 74 0 DIG12
port 18 nsew
rlabel metal2 5529 15 5732 81 0 DIG11
port 19 nsew
rlabel metal2 5133 17 5336 83 0 DIG10
port 20 nsew
rlabel metal2 4735 11 4938 77 0 DIG09
port 21 nsew
rlabel metal2 4318 9 4521 75 0 DIG08
port 22 nsew
rlabel metal2 3909 11 4112 77 0 DIG07
port 23 nsew
rlabel metal2 3513 8 3716 74 0 DIG06
port 24 nsew
rlabel metal2 3110 9 3313 75 0 DIG05
port 25 nsew
rlabel metal2 2705 11 2908 77 0 DIG04
port 26 nsew
rlabel metal2 2305 11 2508 77 0 DIG03
port 27 nsew
rlabel metal2 1909 11 2112 77 0 DIG02
port 28 nsew
rlabel metal2 1502 8 1705 74 0 DIG01
port 29 nsew
rlabel metal2 11587 2160 11664 2369 0 CAP2    
port 30 nsew
rlabel metal2 11542 2711 11632 2920 0 GENERALGATE01   
port 31 nsew
rlabel metal2 11545 3219 11635 3428 0 GATEANDCAP1    
port 32 nsew
rlabel metal2 11542 3737 11632 3946 0 GENERALGATE02
port 33 nsew
rlabel metal2 11542 4225 11632 4434 0 OUTPUTTA1    
port 34 nsew
rlabel metal2 11542 4763 11632 4972 0 GATENFET1   
port 35 nsew
rlabel metal2 11545 5208 11635 5417 0 DACOUTPUT  
port 36 nsew
rlabel metal2 11546 5646 11632 5856 0 DRAINOUT
port 37 nsew
rlabel metal2 11546 6085 11632 6295 0 ROWTERM2
port 38 nsew
rlabel metal2 11549 6494 11635 6704 0 COLUMN2
port 39 nsew
rlabel metal2 11549 6907 11635 7117 0 COLUMN1
port 40 nsew
rlabel metal1 10055 7080 10374 7192 0 GATE2
port 41 nsew
rlabel metal1 7198 7077 7517 7189 0 GATE1
port 61 nsew
rlabel metal1 4339 7078 4658 7190 0 DRAININJECT
port 42 nsew
rlabel metal1 2808 7031 2942 7132 0 VTUN
port 43 nsew
rlabel metal2 77 6929 145 7161 0 VREFCHAR
port 44 nsew
rlabel metal2 77 6476 145 6708 0 CHAROUTPUT
port 45 nsew
rlabel metal2 32 6029 100 6261 0 LARGECAPACITOR
port 46 nsew
rlabel metal2 1161 1713 1198 1754 0 DRAIN6N
port 47 nsew
rlabel metal2 1161 985 1198 1026 0 DRAIN6P
port 48 nsew
rlabel metal2 1165 2677 1202 2718 0 DRAIN5P
port 49 nsew
rlabel metal2 1165 2773 1202 2814 0 DARIN4P
port 50 nsew
rlabel metal2 1165 3143 1202 3184 0 DRAIN5N
port 51 nsew
rlabel metal2 1165 3207 1202 3248 0 DRAIN4N
port 52 nsew
rlabel metal2 1165 4950 1202 4991 0 DRAIN3P
port 53 nsew
rlabel metal2 1165 5046 1202 5087 0 DRAIN2P
port 54 nsew
rlabel metal2 1165 5142 1202 5183 0 DRAIN1P
port 55 nsew
rlabel metal2 1165 5254 1202 5295 0 DRAIN3N
port 56 nsew
rlabel metal2 1165 5347 1202 5388 0 DRAIN2N
port 57 nsew
rlabel metal2 1165 5450 1202 5491 0 DRAIN1N
port 58 nsew
rlabel metal2 1135 5558 1165 5598 0 SOURCEN
port 59 nsew
rlabel metal2 1135 5640 1165 5680 0 SOURCEP
port 60 nsew
rlabel metal2 61 6339 106 6379 0 VGND
port 63 nsew
rlabel metal2 65 6780 110 6820 0 VINJ
port 62 nsew
rlabel metal2 32 5950 83 5991 0 VINJ
port 62 nsew
rlabel metal2 28 5860 79 5901 0 VGND
port 63 nsew
rlabel metal2 80 2348 143 2390 0 VINJ
port 62 nsew
rlabel metal2 78 2251 141 2293 0 VGND
port 63 nsew
rlabel metal2 11645 5513 11690 5558 0 VPWR
port 64 nsew
rlabel metal1 5420 7164 5493 7194 0 VINJ
port 62 nsew
rlabel metal1 5936 7173 6033 7194 0 VGND
port 63 nsew
rlabel metal2 11593 2473 11659 2588 0 VPWR
port 64 nsew
rlabel metal1 4982 8 5074 81 0 VPWR
port 64 nsew
rlabel metal1 6175 8 6267 81 0 VPWR
port 64 nsew
<< end >>
