magic
tech sky130A
timestamp 1634057754
<< checkpaint >>
rect -611 1157 821 1253
rect -612 -128 821 1157
rect -612 -512 810 -128
rect -611 -608 810 -512
<< error_s >>
rect 1 522 40 525
rect 1 480 40 483
rect 0 426 39 429
rect 0 384 39 387
rect 0 330 39 333
rect 0 288 39 291
rect 0 234 39 237
rect 0 192 39 195
rect 0 138 39 141
rect 0 96 39 99
rect 1 42 40 45
rect 1 0 40 3
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_6
timestamp 1634057724
transform 1 0 18 0 1 406
box 0 0 161 121
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_3
timestamp 1634057724
transform 1 0 18 0 1 310
box 0 0 161 121
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_4
timestamp 1634057724
transform 1 0 18 0 1 214
box 0 0 161 121
use sky130_hilas_pFETdevice01  sky130_hilas_pFETdevice01_0
timestamp 1634057724
transform 1 0 18 0 1 118
box 0 0 161 121
use sky130_hilas_pFETdevice01aa  sky130_hilas_pFETdevice01aa_0
timestamp 1634057725
transform 1 0 19 0 1 502
box 0 0 172 121
use sky130_hilas_pFETdevice01a  sky130_hilas_pFETdevice01a_0
timestamp 1634057723
transform 1 0 19 0 1 22
box 0 0 161 85
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
