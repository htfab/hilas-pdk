magic
tech sky130A
timestamp 1607481960
<< error_s >>
rect 1737 475 1741 489
rect 704 359 706 360
rect 1742 -3 1797 562
rect 2075 497 3085 574
rect 3191 490 3212 562
use sky130_hilas_DAC_bit6_01  sky130_hilas_DAC_bit6_01_0
timestamp 1607481960
transform 1 0 1323 0 1 -530
box 402 524 2040 1892
use sky130_hilas_DAC5bit01  sky130_hilas_DAC5bit01_0
timestamp 1607480617
transform 1 0 -359 0 1 -530
box 382 524 2040 1121
<< end >>
