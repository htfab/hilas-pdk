magic
tech sky130A
timestamp 1628616692
<< metal3 >>
rect 0 580 231 583
rect 0 2 423 580
rect 228 0 423 2
<< mimcap >>
rect 60 143 382 542
rect 60 129 104 143
rect 118 129 132 143
rect 146 129 160 143
rect 174 129 188 143
rect 202 129 216 143
rect 230 129 243 143
rect 257 129 271 143
rect 285 129 299 143
rect 313 129 382 143
rect 60 42 382 129
<< mimcapcontact >>
rect 104 129 118 143
rect 132 129 146 143
rect 160 129 174 143
rect 188 129 202 143
rect 216 129 230 143
rect 243 129 257 143
rect 271 129 285 143
rect 299 129 313 143
<< metal4 >>
rect 38 143 339 157
rect 38 129 104 143
rect 118 129 132 143
rect 146 129 160 143
rect 174 129 188 143
rect 202 129 216 143
rect 230 129 243 143
rect 257 129 271 143
rect 285 129 299 143
rect 313 129 339 143
rect 38 110 339 129
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
