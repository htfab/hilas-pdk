magic
tech sky130A
timestamp 1628698532
<< nwell >>
rect -61 112 158 285
<< pmos >>
rect -40 164 28 194
rect 64 164 132 194
<< pdiff >>
rect -40 218 28 224
rect -40 201 -32 218
rect -14 201 4 218
rect 22 201 28 218
rect -40 194 28 201
rect 64 218 132 224
rect 64 201 72 218
rect 90 201 109 218
rect 128 201 132 218
rect 64 194 132 201
rect -40 157 28 164
rect -40 140 -32 157
rect -14 140 4 157
rect 22 140 28 157
rect -40 131 28 140
rect 64 157 132 164
rect 64 140 70 157
rect 88 140 106 157
rect 124 140 132 157
rect 64 136 132 140
rect 71 131 132 136
<< pdiffc >>
rect -32 201 -14 218
rect 4 201 22 218
rect 72 201 90 218
rect 109 201 128 218
rect -32 140 -14 157
rect 4 140 22 157
rect 70 140 88 157
rect 106 140 124 157
<< nsubdiff >>
rect -40 253 28 265
rect -40 236 -32 253
rect -14 236 4 253
rect 22 236 28 253
rect -40 224 28 236
rect 64 253 132 265
rect 64 236 72 253
rect 90 236 109 253
rect 128 236 132 253
rect 64 224 132 236
<< nsubdiffcont >>
rect -32 236 -14 253
rect 4 236 22 253
rect 72 236 90 253
rect 109 236 128 253
<< poly >>
rect -53 164 -40 194
rect 28 164 64 194
rect 132 164 145 194
rect 36 120 53 164
rect 30 112 57 120
rect 30 95 35 112
rect 52 95 57 112
rect 30 87 57 95
<< polycont >>
rect 35 95 52 112
<< locali >>
rect -40 236 -32 253
rect -14 236 4 253
rect 22 236 72 253
rect 90 236 109 253
rect 128 236 136 253
rect -40 218 136 236
rect -40 201 -32 218
rect -14 201 4 218
rect 22 201 72 218
rect 90 201 109 218
rect 128 201 136 218
rect -40 140 -32 157
rect -14 140 4 157
rect 22 140 31 157
rect 62 140 70 157
rect 88 140 106 157
rect 124 140 132 157
rect -5 123 31 140
rect -5 112 60 123
rect -5 95 35 112
rect 52 95 60 112
rect -5 87 60 95
rect -5 82 22 87
rect 85 82 110 140
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
