magic
tech sky130A
timestamp 1628704282
<< checkpaint >>
rect -630 -630 1198 1245
<< metal2 >>
rect 57 559 130 560
rect 57 543 199 559
rect 57 542 130 543
rect 57 372 124 374
rect 57 356 196 372
rect 57 257 127 258
rect 57 241 200 257
rect 57 57 203 74
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_0
timestamp 1628704264
transform 1 0 232 0 1 338
box -232 -45 336 125
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_3
timestamp 1628704264
transform 1 0 232 0 -1 277
box -232 -45 336 125
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_1
timestamp 1628704264
transform 1 0 232 0 -1 570
box -232 -45 336 125
use sky130_hilas_TgateVinj01  sky130_hilas_TgateVinj01_2
timestamp 1628704264
transform 1 0 232 0 1 45
box -232 -45 336 125
<< labels >>
rlabel metal2 57 542 62 560 0 drain1
rlabel metal2 57 356 62 374 0 drain2
rlabel metal2 57 241 62 258 0 drain3
rlabel metal2 57 57 62 74 0 drain4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
