VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_overlapcap02a
  CLASS BLOCK ;
  FOREIGN sky130_hilas_overlapcap02a ;
  ORIGIN 5.210 0.540 ;
  SIZE 4.000 BY 1.640 ;
  OBS
      LAYER nwell ;
        RECT -5.210 -0.540 -1.210 1.100 ;
      LAYER li1 ;
        RECT -4.860 -0.210 -1.550 0.770 ;
      LAYER mcon ;
        RECT -3.290 0.540 -3.120 0.710 ;
        RECT -3.290 0.190 -3.120 0.360 ;
        RECT -3.290 -0.150 -3.120 0.020 ;
      LAYER met1 ;
        RECT -3.330 0.130 -3.090 0.770 ;
        RECT -3.320 -0.130 -3.090 0.130 ;
        RECT -3.320 -0.350 -3.080 -0.130 ;
  END
END sky130_hilas_overlapcap02a
END LIBRARY

