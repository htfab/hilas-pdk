magic
tech sky130A
timestamp 1629420194
<< psubdiff >>
rect 77 642 117 896
rect 77 625 88 642
rect 105 625 117 642
rect 77 608 117 625
rect 77 591 88 608
rect 105 591 117 608
rect 77 574 117 591
rect 77 557 88 574
rect 105 557 117 574
rect 77 537 117 557
<< psubdiffcont >>
rect 88 625 105 642
rect 88 591 105 608
rect 88 557 105 574
<< poly >>
rect 126 988 428 1003
rect 126 725 145 988
rect 126 710 429 725
rect 126 523 146 710
rect 78 513 146 523
rect 78 496 83 513
rect 100 496 117 513
rect 134 496 146 513
rect 78 479 146 496
rect 78 462 84 479
rect 101 462 118 479
rect 135 462 146 479
rect 78 447 146 462
rect 78 445 428 447
rect 78 428 84 445
rect 101 428 118 445
rect 135 430 428 445
rect 135 428 161 430
rect 78 423 161 428
rect 78 420 147 423
<< polycont >>
rect 83 496 100 513
rect 117 496 134 513
rect 84 462 101 479
rect 118 462 135 479
rect 84 428 101 445
rect 118 428 135 445
<< locali >>
rect 159 700 176 738
rect 214 700 231 738
rect 269 700 286 738
rect 324 700 341 738
rect 379 700 396 738
rect 434 700 451 738
rect 88 642 105 645
rect 88 608 105 609
rect 88 574 105 591
rect 83 513 134 521
rect 100 496 117 513
rect 83 495 134 496
rect 83 488 135 495
rect 84 479 135 488
rect 101 462 118 479
rect 84 445 135 462
rect 101 428 118 445
rect 84 420 135 428
<< viali >>
rect 88 645 105 662
rect 88 625 105 626
rect 88 609 105 625
rect 88 540 105 557
<< metal1 >>
rect 82 665 109 668
rect 82 662 110 665
rect 82 645 88 662
rect 105 645 110 662
rect 82 626 110 645
rect 82 612 88 626
rect 64 609 88 612
rect 105 609 110 626
rect 64 582 110 609
rect 64 580 111 582
rect 82 557 111 580
rect 82 540 88 557
rect 105 540 111 557
rect 82 537 111 540
<< metal2 >>
rect 97 979 403 980
rect 88 946 403 979
rect 88 701 120 946
rect 207 878 501 908
rect 426 874 501 878
rect 463 861 501 874
rect 466 774 501 861
rect 206 741 501 774
rect 88 668 404 701
rect 88 564 120 668
rect 88 532 404 564
rect 64 420 124 502
rect 466 497 501 741
rect 207 465 501 497
rect 207 464 478 465
use sky130_hilas_li2m2  sky130_hilas_li2m2_10
timestamp 1629420194
transform 1 0 274 0 1 546
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_6
timestamp 1629420194
transform 1 0 384 0 1 546
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_15
timestamp 1629420194
transform 1 0 220 0 1 478
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_17
timestamp 1629420194
transform 1 0 329 0 1 478
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_19
timestamp 1629420194
transform 1 0 439 0 1 479
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_9
timestamp 1629420194
transform 1 0 164 0 1 546
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_7
timestamp 1629420194
transform 1 0 108 0 1 435
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_8
timestamp 1629420194
transform 1 0 107 0 1 482
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1629420194
transform 1 0 274 0 1 683
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1629420194
transform 1 0 384 0 1 683
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1629420194
transform 1 0 164 0 1 683
box -14 -15 20 18
use sky130_hilas_nFETLargePart1  sky130_hilas_nFETLargePart1_1
timestamp 1629420194
transform 1 0 319 0 1 473
box -165 -31 137 241
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1629420194
transform 1 0 329 0 1 756
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_4
timestamp 1629420194
transform 1 0 220 0 1 756
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_5
timestamp 1629420194
transform 1 0 439 0 1 756
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_14
timestamp 1629420194
transform 1 0 274 0 1 961
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_18
timestamp 1629420194
transform 1 0 384 0 1 960
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_11
timestamp 1629420194
transform 1 0 165 0 1 961
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_16
timestamp 1629420194
transform 1 0 220 0 1 893
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_12
timestamp 1629420194
transform 1 0 329 0 1 891
box -14 -15 20 18
use sky130_hilas_li2m2  sky130_hilas_li2m2_13
timestamp 1629420194
transform 1 0 440 0 1 890
box -14 -15 20 18
use sky130_hilas_nFETLargePart1  sky130_hilas_nFETLargePart1_0
timestamp 1629420194
transform 1 0 319 0 1 751
box -165 -31 137 241
<< labels >>
rlabel metal2 486 834 500 908 0 DRAIN
port 3 nsew analog default
rlabel metal2 88 905 102 979 0 SOURCE
port 2 nsew analog default
rlabel metal2 64 420 74 502 0 GATE
port 1 nsew analog default
rlabel metal1 64 580 71 612 0 VGND
port 4 nsew
<< end >>
