magic
tech sky130A
timestamp 1628616976
<< checkpaint >>
rect -405 1318 988 1384
rect -606 1294 988 1318
rect -665 -545 988 1294
rect -606 -569 988 -545
rect -405 -638 988 -569
<< error_s >>
rect 50 651 77 657
rect 50 609 77 615
rect 50 584 77 590
rect 50 542 77 548
rect 50 501 77 507
rect 50 459 77 465
rect 50 434 77 440
rect 50 392 77 398
rect 50 351 77 357
rect 50 309 77 315
rect 50 284 77 290
rect 50 242 77 248
rect 50 201 77 207
rect 50 159 77 165
rect 50 134 77 140
rect 50 92 77 98
<< metal1 >>
rect 96 89 130 661
rect 163 90 190 660
<< metal2 >>
rect 1 618 255 641
rect 27 404 292 427
rect 1 322 292 344
rect 0 105 271 128
use sky130_hilas_li2m2  sky130_hilas_li2m2_3
timestamp 1628616688
transform 1 0 235 0 1 114
box 0 0 34 33
use sky130_hilas_pFETmirror02  sky130_hilas_pFETmirror02_0
timestamp 1628616729
transform 1 0 225 0 1 0
box 0 0 133 292
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_0
timestamp 1628616972
transform 1 0 24 0 -1 208
box 0 0 184 147
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_1
timestamp 1628616972
transform 1 0 24 0 1 241
box 0 0 184 147
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1628616972
transform 1 0 178 0 1 237
box 0 0 23 29
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1628616688
transform 1 0 244 0 1 411
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1628616688
transform 1 0 243 0 1 339
box 0 0 34 33
use sky130_hilas_pFETmirror02  sky130_hilas_pFETmirror02_1
timestamp 1628616729
transform 1 0 225 0 -1 746
box 0 0 133 292
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_2
timestamp 1628616972
transform 1 0 24 0 1 541
box 0 0 184 147
use sky130_hilas_nMirror03  sky130_hilas_nMirror03_3
timestamp 1628616972
transform 1 0 24 0 -1 508
box 0 0 184 147
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1628616972
transform 1 0 178 0 1 496
box 0 0 23 29
use sky130_hilas_li2m2  sky130_hilas_li2m2_2
timestamp 1628616688
transform 1 0 239 0 1 633
box 0 0 34 33
<< labels >>
rlabel metal2 281 404 292 427 0 output1
rlabel space 281 322 292 345 0 output2
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
