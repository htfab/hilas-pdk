* Copyright 2020 The Hilas PDK Authors
* 
* This file is part of HILAS.
* 
* HILAS is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published by
* the Free Software Foundation, version 3 of the License.
* 
* HILAS is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
* 
* You should have received a copy of the GNU Lesser General Public License
* along with HILAS.  If not, see <https://www.gnu.org/licenses/>.
* 
* Licensed under the Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
* https://www.gnu.org/licenses/lgpl-3.0.en.html
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
* SPDX-License-Identifier: LGPL-3.0
* 
* 

* NGSPICE file created from sky130_hilas_TA2Cell_1FG_Strong.ext - technology: sky130A

.subckt sky130_hilas_nFET03 a_n62_n12# SUB a_54_n12# a_0_n38#
X0 a_54_n12# a_0_n38# a_n62_n12# SUB sky130_fd_pr__nfet_01v8 w=350000u l=270000u
.ends

.subckt sky130_hilas_nMirror03 sky130_hilas_nFET03_1/a_n62_n12# a_n92_86# sky130_hilas_li2m2_1/SUB
Xsky130_hilas_nFET03_0 a_n92_86# sky130_hilas_li2m2_1/SUB sky130_hilas_li2m2_1/SUB
+ a_n92_86# sky130_hilas_nFET03
Xsky130_hilas_nFET03_1 sky130_hilas_nFET03_1/a_n62_n12# sky130_hilas_li2m2_1/SUB sky130_hilas_li2m2_1/SUB
+ a_n92_86# sky130_hilas_nFET03
.ends

.subckt sky130_hilas_pFETmirror02 w_n122_178# SUB a_n80_650# a_n80_262#
X0 a_n80_650# a_n80_262# w_n122_178# w_n122_178# sky130_fd_pr__pfet_01v8 w=680000u l=300000u
X1 w_n122_178# a_n80_262# a_n80_262# w_n122_178# sky130_fd_pr__pfet_01v8 w=680000u l=300000u
.ends

.subckt sky130_hilas_DualTACore01 sky130_hilas_nMirror03_3/a_n92_86# sky130_hilas_nMirror03_2/a_n92_86#
+ sky130_hilas_nMirror03_1/a_n92_86# sky130_hilas_nMirror03_0/a_n92_86# SUB m1_52_n42#
Xsky130_hilas_nMirror03_3 output1 sky130_hilas_nMirror03_3/a_n92_86# SUB sky130_hilas_nMirror03
Xsky130_hilas_pFETmirror02_0 m1_52_n42# SUB m2_n272_422# m2_n274_n12# sky130_hilas_pFETmirror02
Xsky130_hilas_pFETmirror02_1 m1_52_n42# SUB output1 m2_n272_1014# sky130_hilas_pFETmirror02
Xsky130_hilas_nMirror03_0 m2_n274_n12# sky130_hilas_nMirror03_0/a_n92_86# SUB sky130_hilas_nMirror03
Xsky130_hilas_nMirror03_2 m2_n272_1014# sky130_hilas_nMirror03_2/a_n92_86# SUB sky130_hilas_nMirror03
Xsky130_hilas_nMirror03_1 m2_n272_422# sky130_hilas_nMirror03_1/a_n92_86# SUB sky130_hilas_nMirror03
.ends

.subckt sky130_hilas_TunCap01 SUB a_n2872_n666# w_n2902_n800#
X0 a_n2872_n666# w_n2902_n800# w_n2902_n800# sky130_fd_pr__cap_var w=590000u l=500000u
.ends

.subckt sky130_hilas_horizTransCell01 a_n512_284# a_n952_238# SUB a_n346_284# a_n654_284#
+ a_n926_284# a_n952_338# a_n952_496# a_n654_438# a_n926_438# a_n300_130# a_n512_162#
+ w_n728_96# a_n654_596# a_n926_596#
X0 w_n728_96# a_n300_130# a_n344_162# w_n728_96# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
X1 a_n346_284# a_n952_238# a_n512_284# w_n728_96# sky130_fd_pr__pfet_g5v0d10v5 w=1.84e+06u l=510000u
X2 a_n654_438# a_n952_338# a_n654_284# w_n728_96# sky130_fd_pr__pfet_g5v0d10v5 w=390000u l=500000u
X3 a_n654_596# a_n952_496# a_n654_438# w_n728_96# sky130_fd_pr__pfet_g5v0d10v5 w=390000u l=500000u
X4 a_n926_438# a_n952_338# a_n926_284# SUB sky130_fd_pr__nfet_g5v0d10v5 w=400000u l=500000u
X5 a_n926_596# a_n952_496# a_n926_438# SUB sky130_fd_pr__nfet_g5v0d10v5 w=400000u l=500000u
X6 a_n344_162# a_n952_238# a_n512_162# w_n728_96# sky130_fd_pr__pfet_g5v0d10v5 w=310000u l=500000u
.ends

.subckt sky130_hilas_FGVaractorCapacitor02 a_n1882_n644# SUB w_n2010_n760#
X0 a_n1882_n644# w_n2010_n760# w_n2010_n760# sky130_fd_pr__cap_var w=1.11e+06u l=500000u
.ends

.subckt sky130_hilas_FGBias2x1cell VTUN VGND GATE_CONTROL DRAIN1 DRAIN4 VINJ OUTPUT1
+ OUTPUT2 GateColSelect
Xsky130_hilas_TunCap01_1 VGND a_n560_n620# VTUN sky130_hilas_TunCap01
Xsky130_hilas_horizTransCell01_0 OUTPUT2 a_n560_n620# VGND VINJ sky130_hilas_horizTransCell01_0/a_n654_284#
+ sky130_hilas_horizTransCell01_0/a_n926_284# sky130_hilas_horizTransCell01_0/a_n952_338#
+ sky130_hilas_horizTransCell01_0/a_n952_496# li_934_n408# sky130_hilas_horizTransCell01_0/a_n926_438#
+ GateColSelect DRAIN4 VINJ li_948_n216# sky130_hilas_horizTransCell01_0/a_n926_596#
+ sky130_hilas_horizTransCell01
Xsky130_hilas_TunCap01_3 VGND a_n474_252# VTUN sky130_hilas_TunCap01
Xsky130_hilas_horizTransCell01_1 OUTPUT1 a_n474_252# VGND VINJ sky130_hilas_horizTransCell01_1/a_n654_284#
+ sky130_hilas_horizTransCell01_1/a_n926_284# sky130_hilas_horizTransCell01_1/a_n952_338#
+ sky130_hilas_horizTransCell01_1/a_n952_496# li_934_56# sky130_hilas_horizTransCell01_1/a_n926_438#
+ GateColSelect DRAIN1 VINJ li_948_n216# sky130_hilas_horizTransCell01_1/a_n926_596#
+ sky130_hilas_horizTransCell01
Xsky130_hilas_FGVaractorCapacitor02_0 a_n560_n620# VGND GATE_CONTROL sky130_hilas_FGVaractorCapacitor02
Xsky130_hilas_FGVaractorCapacitor02_2 a_n474_252# VGND GATE_CONTROL sky130_hilas_FGVaractorCapacitor02
.ends

.subckt sky130_hilas_pTransistorVert01 a_n658_n792# a_n596_n822# SUB a_n496_n792#
+ w_n726_n888#
X0 a_n496_n792# a_n596_n822# a_n658_n792# w_n726_n888# sky130_fd_pr__pfet_g5v0d10v5 w=2.03e+06u l=500000u
.ends

.subckt sky130_hilas_pTransistorPair m2_510_n704# w_534_n338# li_348_n384# SUB a_454_n814#
+ a_450_n208# m2_546_n498#
Xsky130_hilas_pTransistorVert01_0 li_348_n384# a_450_n208# SUB m2_546_n498# w_534_n338#
+ sky130_hilas_pTransistorVert01
Xsky130_hilas_pTransistorVert01_1 li_348_n384# a_454_n814# SUB m2_510_n704# w_534_n338#
+ sky130_hilas_pTransistorVert01
.ends

.subckt sky130_hilas_FGtrans2x1cell GATESELECT VINJ DRAIN1 DRAIN4 PROG RUN GATE1 GATE2
+ PROGGATE VGND VTUN DRAIN VS
Xsky130_hilas_TunCap01_1 VGND a_n560_n620# VTUN sky130_hilas_TunCap01
Xsky130_hilas_horizTransCell01_0 DRAIN a_n560_n620# VGND VS PROGGATE GATE1 RUN PROG
+ li_724_n408# li_724_n408# GATESELECT DRAIN4 VINJ GATE1 PROGGATE sky130_hilas_horizTransCell01
Xsky130_hilas_TunCap01_3 VGND a_n474_252# VTUN sky130_hilas_TunCap01
Xsky130_hilas_horizTransCell01_1 DRAIN1 a_n474_252# VGND VS PROGGATE GATE2 RUN PROG
+ li_724_56# li_724_56# GATESELECT DRAIN1 VINJ GATE2 PROGGATE sky130_hilas_horizTransCell01
Xsky130_hilas_FGVaractorCapacitor02_0 a_n560_n620# VGND li_724_n408# sky130_hilas_FGVaractorCapacitor02
Xsky130_hilas_FGVaractorCapacitor02_2 a_n474_252# VGND li_724_56# sky130_hilas_FGVaractorCapacitor02
.ends

.subckt sky130_hilas_TA2Cell_1FG_Strong VTUN VGATE2 PROG VGATE1 VINP_AMP1
Xsky130_hilas_DualTACore01_0 m2_n294_1062# m2_n308_1242# sky130_hilas_FGBias2x1cell_0/DRAIN1
+ sky130_hilas_FGtrans2x1cell_0/DRAIN SUB Vdd sky130_hilas_DualTACore01
Xsky130_hilas_FGBias2x1cell_0 VTUN SUB VGATE2 sky130_hilas_FGBias2x1cell_0/DRAIN1
+ sky130_hilas_FGBias2x1cell_0/DRAIN4 Vdd sky130_hilas_FGBias2x1cell_0/OUTPUT1 sky130_hilas_FGtrans2x1cell_0/VS
+ GateColSelect sky130_hilas_FGBias2x1cell
Xsky130_hilas_pTransistorPair_1 m2_n308_1242# Vdd sky130_hilas_FGBias2x1cell_0/OUTPUT1
+ SUB Vin-_Amp2 Vin+_Amp2 m2_n294_1062# sky130_hilas_pTransistorPair
Xsky130_hilas_FGtrans2x1cell_0 sky130_hilas_FGtrans2x1cell_0/GATESELECT sky130_hilas_FGtrans2x1cell_0/VINJ
+ sky130_hilas_FGBias2x1cell_0/DRAIN1 sky130_hilas_FGBias2x1cell_0/DRAIN4 PROG PROG
+ Vin-_Amp1 VINP_AMP1 VGATE1 SUB VTUN sky130_hilas_FGtrans2x1cell_0/DRAIN sky130_hilas_FGtrans2x1cell_0/VS
+ sky130_hilas_FGtrans2x1cell
.ends

